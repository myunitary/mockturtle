module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 ;
  assign n22 = x5 & x13 ;
  assign n23 = x6 & x14 ;
  assign n24 = n22 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n22 ^ x5 ;
  assign n28 = n27 ^ x13 ;
  assign n29 = x4 & x12 ;
  assign n30 = n29 ^ x4 ;
  assign n31 = n30 ^ x12 ;
  assign n32 = n28 & n31 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ n28 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = n26 & ~n36 ;
  assign n38 = n37 ^ n26 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ n36 ;
  assign n17 = x10 ^ x2 ;
  assign n41 = x11 ^ x3 ;
  assign n42 = ~n17 & n41 ;
  assign n43 = ~n29 & n42 ;
  assign n44 = ~n40 & n43 ;
  assign n18 = x3 & x11 ;
  assign n19 = n18 ^ x3 ;
  assign n20 = n19 ^ x11 ;
  assign n21 = ~n17 & ~n20 ;
  assign n45 = n44 ^ n21 ;
  assign n56 = x1 & x9 ;
  assign n57 = x8 & n56 ;
  assign n58 = n57 ^ n56 ;
  assign n66 = n45 & n58 ;
  assign n67 = n66 ^ n58 ;
  assign n47 = x7 & x15 ;
  assign n46 = x14 ^ x6 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = x13 ^ x5 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = ~n49 & n50 ;
  assign n52 = n51 ^ n46 ;
  assign n53 = n48 & ~n52 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = n54 ^ n47 ;
  assign n59 = x12 ^ x4 ;
  assign n60 = n41 & n59 ;
  assign n61 = n58 & n60 ;
  assign n62 = n61 ^ n60 ;
  assign n63 = n55 & n62 ;
  assign n64 = n45 & n63 ;
  assign n65 = n64 ^ n63 ;
  assign n68 = n67 ^ n65 ;
  assign n70 = x9 ^ x1 ;
  assign n71 = x2 & x10 ;
  assign n72 = ~n70 & ~n71 ;
  assign n82 = n68 & n72 ;
  assign n83 = n82 ^ n68 ;
  assign n69 = n55 & n60 ;
  assign n73 = ~x0 & x8 ;
  assign n74 = ~n56 & n73 ;
  assign n75 = n74 ^ x8 ;
  assign n76 = n75 ^ n56 ;
  assign n77 = n72 & ~n76 ;
  assign n78 = n77 ^ n72 ;
  assign n79 = n78 ^ n76 ;
  assign n80 = n69 & n79 ;
  assign n81 = n68 & n80 ;
  assign n84 = n83 ^ n81 ;
  assign n85 = n18 & n29 ;
  assign n86 = n85 ^ n18 ;
  assign n87 = n86 ^ n29 ;
  assign n88 = n71 ^ x2 ;
  assign n89 = n88 ^ x10 ;
  assign n90 = ~n20 & ~n89 ;
  assign n91 = n90 ^ n20 ;
  assign n92 = n91 ^ n89 ;
  assign n93 = n87 & ~n92 ;
  assign n94 = n93 ^ n92 ;
  assign n95 = ~n40 & ~n94 ;
  assign n96 = n95 ^ n92 ;
  assign n97 = ~x0 & ~x8 ;
  assign n98 = ~n56 & ~n71 ;
  assign n99 = ~n97 & n98 ;
  assign n100 = ~n96 & n99 ;
  assign n101 = n100 ^ n99 ;
  assign n110 = x2 & n41 ;
  assign n111 = ~n29 & n110 ;
  assign n112 = ~n40 & n111 ;
  assign n108 = x2 & ~n20 ;
  assign n109 = n108 ^ x2 ;
  assign n113 = n112 ^ n109 ;
  assign n114 = ~x0 & x1 ;
  assign n115 = ~x8 & x9 ;
  assign n116 = n114 & n115 ;
  assign n117 = x10 & n116 ;
  assign n118 = n113 & n117 ;
  assign n102 = n56 ^ x1 ;
  assign n103 = n102 ^ x9 ;
  assign n104 = n103 ^ x8 ;
  assign n105 = n103 ^ x0 ;
  assign n106 = ~n104 & ~n105 ;
  assign n107 = n106 ^ n103 ;
  assign n119 = n118 ^ n107 ;
  assign n120 = n101 & ~n119 ;
  assign n121 = n120 ^ n101 ;
  assign n122 = n121 ^ n119 ;
  assign n123 = n84 & n122 ;
  assign n124 = n123 ^ n84 ;
  assign n125 = n124 ^ n122 ;
  assign n126 = n113 ^ n70 ;
  assign n127 = n20 & ~n87 ;
  assign n128 = ~n40 & n127 ;
  assign n129 = n128 ^ n17 ;
  assign n130 = n129 ^ n20 ;
  assign n131 = n126 & n130 ;
  assign n134 = x8 ^ x0 ;
  assign n137 = n134 ^ n56 ;
  assign n138 = n137 ^ n69 ;
  assign n139 = n131 & n138 ;
  assign n132 = n70 & ~n89 ;
  assign n133 = n103 & ~n132 ;
  assign n135 = n134 ^ n133 ;
  assign n136 = ~n131 & n135 ;
  assign n140 = n139 ^ n136 ;
  assign n142 = n126 ^ n69 ;
  assign n141 = n89 ^ n70 ;
  assign n143 = n142 ^ n141 ;
  assign n144 = ~n130 & ~n143 ;
  assign n145 = n144 ^ n143 ;
  assign n146 = n145 ^ n130 ;
  assign n147 = n146 ^ n141 ;
  assign n148 = n130 ^ n69 ;
  assign n149 = n46 & n47 ;
  assign n150 = ~n26 & ~n149 ;
  assign n151 = n28 & ~n150 ;
  assign n152 = ~n29 & ~n151 ;
  assign n153 = n31 & ~n152 ;
  assign n154 = n153 ^ n41 ;
  assign n155 = ~n23 & ~n55 ;
  assign n156 = n49 & ~n155 ;
  assign n157 = ~n22 & ~n156 ;
  assign n158 = n157 ^ n59 ;
  assign n159 = ~n23 & ~n149 ;
  assign n160 = n159 ^ n49 ;
  assign y0 = ~n125 ;
  assign y1 = n140 ;
  assign y2 = ~n147 ;
  assign y3 = n148 ;
  assign y4 = n154 ;
  assign y5 = ~n158 ;
  assign y6 = ~n160 ;
  assign y7 = n48 ;
endmodule
