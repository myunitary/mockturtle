module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 ;
  assign n152 = x26 ^ x18 ;
  assign n178 = x19 & x27 ;
  assign n179 = n178 ^ x19 ;
  assign n180 = n152 & n179 ;
  assign n181 = n180 ^ n179 ;
  assign n177 = x18 & ~x26 ;
  assign n182 = n181 ^ n177 ;
  assign n147 = x24 ^ x16 ;
  assign n148 = x25 ^ x17 ;
  assign n149 = n147 & n148 ;
  assign n150 = n149 ^ n147 ;
  assign n151 = n150 ^ n148 ;
  assign n194 = x24 & ~n151 ;
  assign n195 = n182 & n194 ;
  assign n173 = x17 & ~x25 ;
  assign n174 = ~n147 & n173 ;
  assign n172 = x16 & ~x24 ;
  assign n175 = n174 ^ n172 ;
  assign n193 = x24 & ~n175 ;
  assign n196 = n195 ^ n193 ;
  assign n153 = x27 ^ x19 ;
  assign n154 = n152 & n153 ;
  assign n155 = n154 ^ n152 ;
  assign n156 = n155 ^ n153 ;
  assign n157 = n151 & n156 ;
  assign n158 = n157 ^ n151 ;
  assign n159 = n158 ^ n156 ;
  assign n129 = x28 ^ x20 ;
  assign n133 = x29 ^ x21 ;
  assign n134 = n129 & n133 ;
  assign n135 = n134 ^ n129 ;
  assign n136 = n135 ^ n133 ;
  assign n138 = x30 ^ x22 ;
  assign n162 = x31 ^ x23 ;
  assign n163 = n138 & n162 ;
  assign n164 = n163 ^ n138 ;
  assign n165 = n164 ^ n162 ;
  assign n166 = n136 & n165 ;
  assign n167 = n166 ^ n136 ;
  assign n168 = n167 ^ n165 ;
  assign n169 = ~n159 & ~n168 ;
  assign n191 = x24 & n169 ;
  assign n192 = n191 ^ x24 ;
  assign n197 = n196 ^ n192 ;
  assign n139 = x23 & x31 ;
  assign n140 = n139 ^ x23 ;
  assign n141 = n138 & n140 ;
  assign n142 = n141 ^ n140 ;
  assign n137 = x22 & ~x30 ;
  assign n143 = n142 ^ n137 ;
  assign n144 = n136 & n143 ;
  assign n145 = n144 ^ n143 ;
  assign n130 = x21 & ~x29 ;
  assign n131 = ~n129 & n130 ;
  assign n128 = x20 & ~x28 ;
  assign n132 = n131 ^ n128 ;
  assign n146 = n145 ^ n132 ;
  assign n189 = x24 & ~n159 ;
  assign n190 = n146 & n189 ;
  assign n198 = n197 ^ n190 ;
  assign n183 = x16 & ~n151 ;
  assign n184 = n182 & n183 ;
  assign n176 = x16 & ~n175 ;
  assign n185 = n184 ^ n176 ;
  assign n170 = x16 & n169 ;
  assign n171 = n170 ^ x16 ;
  assign n186 = n185 ^ n171 ;
  assign n160 = x16 & ~n159 ;
  assign n161 = n146 & n160 ;
  assign n187 = n186 ^ n161 ;
  assign n188 = n187 ^ x16 ;
  assign n199 = n198 ^ n188 ;
  assign n54 = x10 ^ x2 ;
  assign n83 = x3 & x11 ;
  assign n84 = n83 ^ x3 ;
  assign n85 = n54 & n84 ;
  assign n86 = n85 ^ n84 ;
  assign n82 = x2 & ~x10 ;
  assign n87 = n86 ^ n82 ;
  assign n49 = x8 ^ x0 ;
  assign n50 = x9 ^ x1 ;
  assign n51 = n49 & n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n52 ^ n50 ;
  assign n122 = x0 & ~n53 ;
  assign n123 = n87 & n122 ;
  assign n90 = x1 & ~x9 ;
  assign n91 = ~n49 & n90 ;
  assign n89 = x0 & ~x8 ;
  assign n92 = n91 ^ n89 ;
  assign n121 = x0 & ~n92 ;
  assign n124 = n123 ^ n121 ;
  assign n55 = x11 ^ x3 ;
  assign n56 = n54 & n55 ;
  assign n57 = n56 ^ n54 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n53 & n58 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = n60 ^ n58 ;
  assign n63 = x12 ^ x4 ;
  assign n67 = x13 ^ x5 ;
  assign n68 = n63 & n67 ;
  assign n69 = n68 ^ n63 ;
  assign n70 = n69 ^ n67 ;
  assign n72 = x14 ^ x6 ;
  assign n95 = x15 ^ x7 ;
  assign n96 = n72 & n95 ;
  assign n97 = n96 ^ n72 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = n70 & n98 ;
  assign n100 = n99 ^ n70 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = ~n61 & ~n101 ;
  assign n119 = x0 & n102 ;
  assign n120 = n119 ^ x0 ;
  assign n125 = n124 ^ n120 ;
  assign n73 = x7 & x15 ;
  assign n74 = n73 ^ x7 ;
  assign n75 = n72 & n74 ;
  assign n76 = n75 ^ n74 ;
  assign n71 = x6 & ~x14 ;
  assign n77 = n76 ^ n71 ;
  assign n78 = n70 & n77 ;
  assign n79 = n78 ^ n77 ;
  assign n64 = x5 & ~x13 ;
  assign n65 = ~n63 & n64 ;
  assign n62 = x4 & ~x12 ;
  assign n66 = n65 ^ n62 ;
  assign n80 = n79 ^ n66 ;
  assign n117 = x0 & ~n61 ;
  assign n118 = n80 & n117 ;
  assign n126 = n125 ^ n118 ;
  assign n110 = x8 & ~n53 ;
  assign n111 = n87 & n110 ;
  assign n109 = x8 & ~n92 ;
  assign n112 = n111 ^ n109 ;
  assign n107 = x8 & n102 ;
  assign n108 = n107 ^ x8 ;
  assign n113 = n112 ^ n108 ;
  assign n105 = x8 & ~n61 ;
  assign n106 = n80 & n105 ;
  assign n114 = n113 ^ n106 ;
  assign n116 = n114 ^ x8 ;
  assign n127 = n126 ^ n116 ;
  assign n201 = n199 ^ n127 ;
  assign n218 = x25 & ~n151 ;
  assign n219 = n182 & n218 ;
  assign n217 = x25 & ~n175 ;
  assign n220 = n219 ^ n217 ;
  assign n215 = x25 & n169 ;
  assign n216 = n215 ^ x25 ;
  assign n221 = n220 ^ n216 ;
  assign n213 = x25 & ~n159 ;
  assign n214 = n146 & n213 ;
  assign n222 = n221 ^ n214 ;
  assign n207 = x17 & ~n151 ;
  assign n208 = n182 & n207 ;
  assign n206 = x17 & ~n175 ;
  assign n209 = n208 ^ n206 ;
  assign n204 = x17 & n169 ;
  assign n205 = n204 ^ x17 ;
  assign n210 = n209 ^ n205 ;
  assign n202 = x17 & ~n159 ;
  assign n203 = n146 & n202 ;
  assign n211 = n210 ^ n203 ;
  assign n212 = n211 ^ x17 ;
  assign n223 = n222 ^ n212 ;
  assign n240 = x1 & ~n53 ;
  assign n241 = n87 & n240 ;
  assign n239 = x1 & ~n92 ;
  assign n242 = n241 ^ n239 ;
  assign n237 = x1 & n102 ;
  assign n238 = n237 ^ x1 ;
  assign n243 = n242 ^ n238 ;
  assign n235 = x1 & ~n61 ;
  assign n236 = n80 & n235 ;
  assign n244 = n243 ^ n236 ;
  assign n229 = x9 & ~n53 ;
  assign n230 = n87 & n229 ;
  assign n228 = x9 & ~n92 ;
  assign n231 = n230 ^ n228 ;
  assign n226 = x9 & n102 ;
  assign n227 = n226 ^ x9 ;
  assign n232 = n231 ^ n227 ;
  assign n224 = x9 & ~n61 ;
  assign n225 = n80 & n224 ;
  assign n233 = n232 ^ n225 ;
  assign n234 = n233 ^ x9 ;
  assign n245 = n244 ^ n234 ;
  assign n246 = ~n223 & n245 ;
  assign n247 = ~n201 & n246 ;
  assign n200 = n127 & ~n199 ;
  assign n248 = n247 ^ n200 ;
  assign n266 = x2 & ~n53 ;
  assign n267 = n87 & n266 ;
  assign n265 = x2 & ~n92 ;
  assign n268 = n267 ^ n265 ;
  assign n263 = x2 & n102 ;
  assign n264 = n263 ^ x2 ;
  assign n269 = n268 ^ n264 ;
  assign n261 = x2 & ~n61 ;
  assign n262 = n80 & n261 ;
  assign n270 = n269 ^ n262 ;
  assign n255 = x10 & ~n53 ;
  assign n256 = n87 & n255 ;
  assign n254 = x10 & ~n92 ;
  assign n257 = n256 ^ n254 ;
  assign n252 = x10 & n102 ;
  assign n253 = n252 ^ x10 ;
  assign n258 = n257 ^ n253 ;
  assign n250 = x10 & ~n61 ;
  assign n251 = n80 & n250 ;
  assign n259 = n258 ^ n251 ;
  assign n260 = n259 ^ x10 ;
  assign n271 = n270 ^ n260 ;
  assign n1392 = ~n248 & n271 ;
  assign n288 = x26 & ~n151 ;
  assign n289 = n182 & n288 ;
  assign n287 = x26 & ~n175 ;
  assign n290 = n289 ^ n287 ;
  assign n285 = x26 & n169 ;
  assign n286 = n285 ^ x26 ;
  assign n291 = n290 ^ n286 ;
  assign n283 = x26 & ~n159 ;
  assign n284 = n146 & n283 ;
  assign n292 = n291 ^ n284 ;
  assign n277 = x18 & ~n151 ;
  assign n278 = n182 & n277 ;
  assign n276 = x18 & ~n175 ;
  assign n279 = n278 ^ n276 ;
  assign n274 = x18 & n169 ;
  assign n275 = n274 ^ x18 ;
  assign n280 = n279 ^ n275 ;
  assign n272 = x18 & ~n159 ;
  assign n273 = n146 & n272 ;
  assign n281 = n280 ^ n273 ;
  assign n282 = n281 ^ x18 ;
  assign n293 = n292 ^ n282 ;
  assign n295 = n293 ^ n271 ;
  assign n312 = x3 & ~n53 ;
  assign n313 = n87 & n312 ;
  assign n311 = x3 & ~n92 ;
  assign n314 = n313 ^ n311 ;
  assign n309 = x3 & n102 ;
  assign n310 = n309 ^ x3 ;
  assign n315 = n314 ^ n310 ;
  assign n307 = x3 & ~n61 ;
  assign n308 = n80 & n307 ;
  assign n316 = n315 ^ n308 ;
  assign n301 = x11 & ~n53 ;
  assign n302 = n87 & n301 ;
  assign n300 = x11 & ~n92 ;
  assign n303 = n302 ^ n300 ;
  assign n298 = x11 & n102 ;
  assign n299 = n298 ^ x11 ;
  assign n304 = n303 ^ n299 ;
  assign n296 = x11 & ~n61 ;
  assign n297 = n80 & n296 ;
  assign n305 = n304 ^ n297 ;
  assign n306 = n305 ^ x11 ;
  assign n317 = n316 ^ n306 ;
  assign n334 = x27 & ~n151 ;
  assign n335 = n182 & n334 ;
  assign n333 = x27 & ~n175 ;
  assign n336 = n335 ^ n333 ;
  assign n331 = x27 & n169 ;
  assign n332 = n331 ^ x27 ;
  assign n337 = n336 ^ n332 ;
  assign n329 = x27 & ~n159 ;
  assign n330 = n146 & n329 ;
  assign n338 = n337 ^ n330 ;
  assign n323 = x19 & ~n151 ;
  assign n324 = n182 & n323 ;
  assign n322 = x19 & ~n175 ;
  assign n325 = n324 ^ n322 ;
  assign n320 = x19 & n169 ;
  assign n321 = n320 ^ x19 ;
  assign n326 = n325 ^ n321 ;
  assign n318 = x19 & ~n159 ;
  assign n319 = n146 & n318 ;
  assign n327 = n326 ^ n319 ;
  assign n328 = n327 ^ x19 ;
  assign n339 = n338 ^ n328 ;
  assign n340 = n317 & n339 ;
  assign n341 = n340 ^ n317 ;
  assign n342 = n295 & n341 ;
  assign n343 = n342 ^ n341 ;
  assign n294 = n271 & ~n293 ;
  assign n344 = n343 ^ n294 ;
  assign n345 = n245 ^ n223 ;
  assign n346 = n201 & n345 ;
  assign n347 = n346 ^ n201 ;
  assign n348 = n347 ^ n345 ;
  assign n617 = n271 & ~n348 ;
  assign n618 = n344 & n617 ;
  assign n1393 = n1392 ^ n618 ;
  assign n352 = n339 ^ n317 ;
  assign n353 = n295 & n352 ;
  assign n354 = n353 ^ n295 ;
  assign n355 = n354 ^ n352 ;
  assign n356 = n348 & n355 ;
  assign n357 = n356 ^ n348 ;
  assign n358 = n357 ^ n355 ;
  assign n397 = x28 & ~n151 ;
  assign n398 = n182 & n397 ;
  assign n396 = x28 & ~n175 ;
  assign n399 = n398 ^ n396 ;
  assign n394 = x28 & n169 ;
  assign n395 = n394 ^ x28 ;
  assign n400 = n399 ^ n395 ;
  assign n392 = x28 & ~n159 ;
  assign n393 = n146 & n392 ;
  assign n401 = n400 ^ n393 ;
  assign n386 = x20 & ~n151 ;
  assign n387 = n182 & n386 ;
  assign n385 = x20 & ~n175 ;
  assign n388 = n387 ^ n385 ;
  assign n383 = x20 & n169 ;
  assign n384 = n383 ^ x20 ;
  assign n389 = n388 ^ n384 ;
  assign n381 = x20 & ~n159 ;
  assign n382 = n146 & n381 ;
  assign n390 = n389 ^ n382 ;
  assign n391 = n390 ^ x20 ;
  assign n402 = n401 ^ n391 ;
  assign n375 = x4 & ~n53 ;
  assign n376 = n87 & n375 ;
  assign n374 = x4 & ~n92 ;
  assign n377 = n376 ^ n374 ;
  assign n372 = x4 & n102 ;
  assign n373 = n372 ^ x4 ;
  assign n378 = n377 ^ n373 ;
  assign n370 = x4 & ~n61 ;
  assign n371 = n80 & n370 ;
  assign n379 = n378 ^ n371 ;
  assign n364 = x12 & ~n53 ;
  assign n365 = n87 & n364 ;
  assign n363 = x12 & ~n92 ;
  assign n366 = n365 ^ n363 ;
  assign n361 = x12 & n102 ;
  assign n362 = n361 ^ x12 ;
  assign n367 = n366 ^ n362 ;
  assign n359 = x12 & ~n61 ;
  assign n360 = n80 & n359 ;
  assign n368 = n367 ^ n360 ;
  assign n369 = n368 ^ x12 ;
  assign n380 = n379 ^ n369 ;
  assign n403 = n402 ^ n380 ;
  assign n442 = x29 & ~n151 ;
  assign n443 = n182 & n442 ;
  assign n441 = x29 & ~n175 ;
  assign n444 = n443 ^ n441 ;
  assign n439 = x29 & n169 ;
  assign n440 = n439 ^ x29 ;
  assign n445 = n444 ^ n440 ;
  assign n437 = x29 & ~n159 ;
  assign n438 = n146 & n437 ;
  assign n446 = n445 ^ n438 ;
  assign n431 = x21 & ~n151 ;
  assign n432 = n182 & n431 ;
  assign n430 = x21 & ~n175 ;
  assign n433 = n432 ^ n430 ;
  assign n428 = x21 & n169 ;
  assign n429 = n428 ^ x21 ;
  assign n434 = n433 ^ n429 ;
  assign n426 = x21 & ~n159 ;
  assign n427 = n146 & n426 ;
  assign n435 = n434 ^ n427 ;
  assign n436 = n435 ^ x21 ;
  assign n447 = n446 ^ n436 ;
  assign n420 = x5 & ~n53 ;
  assign n421 = n87 & n420 ;
  assign n419 = x5 & ~n92 ;
  assign n422 = n421 ^ n419 ;
  assign n417 = x5 & n102 ;
  assign n418 = n417 ^ x5 ;
  assign n423 = n422 ^ n418 ;
  assign n415 = x5 & ~n61 ;
  assign n416 = n80 & n415 ;
  assign n424 = n423 ^ n416 ;
  assign n409 = x13 & ~n53 ;
  assign n410 = n87 & n409 ;
  assign n408 = x13 & ~n92 ;
  assign n411 = n410 ^ n408 ;
  assign n406 = x13 & n102 ;
  assign n407 = n406 ^ x13 ;
  assign n412 = n411 ^ n407 ;
  assign n404 = x13 & ~n61 ;
  assign n405 = n80 & n404 ;
  assign n413 = n412 ^ n405 ;
  assign n414 = n413 ^ x13 ;
  assign n425 = n424 ^ n414 ;
  assign n448 = n447 ^ n425 ;
  assign n449 = n403 & n448 ;
  assign n450 = n449 ^ n403 ;
  assign n451 = n450 ^ n448 ;
  assign n490 = x30 & ~n151 ;
  assign n491 = n182 & n490 ;
  assign n489 = x30 & ~n175 ;
  assign n492 = n491 ^ n489 ;
  assign n487 = x30 & n169 ;
  assign n488 = n487 ^ x30 ;
  assign n493 = n492 ^ n488 ;
  assign n485 = x30 & ~n159 ;
  assign n486 = n146 & n485 ;
  assign n494 = n493 ^ n486 ;
  assign n479 = x22 & ~n151 ;
  assign n480 = n182 & n479 ;
  assign n478 = x22 & ~n175 ;
  assign n481 = n480 ^ n478 ;
  assign n476 = x22 & n169 ;
  assign n477 = n476 ^ x22 ;
  assign n482 = n481 ^ n477 ;
  assign n474 = x22 & ~n159 ;
  assign n475 = n146 & n474 ;
  assign n483 = n482 ^ n475 ;
  assign n484 = n483 ^ x22 ;
  assign n495 = n494 ^ n484 ;
  assign n468 = x6 & ~n53 ;
  assign n469 = n87 & n468 ;
  assign n467 = x6 & ~n92 ;
  assign n470 = n469 ^ n467 ;
  assign n465 = x6 & n102 ;
  assign n466 = n465 ^ x6 ;
  assign n471 = n470 ^ n466 ;
  assign n463 = x6 & ~n61 ;
  assign n464 = n80 & n463 ;
  assign n472 = n471 ^ n464 ;
  assign n457 = x14 & ~n53 ;
  assign n458 = n87 & n457 ;
  assign n456 = x14 & ~n92 ;
  assign n459 = n458 ^ n456 ;
  assign n454 = x14 & n102 ;
  assign n455 = n454 ^ x14 ;
  assign n460 = n459 ^ n455 ;
  assign n452 = x14 & ~n61 ;
  assign n453 = n80 & n452 ;
  assign n461 = n460 ^ n453 ;
  assign n462 = n461 ^ x14 ;
  assign n473 = n472 ^ n462 ;
  assign n496 = n495 ^ n473 ;
  assign n534 = x7 & ~n53 ;
  assign n535 = n87 & n534 ;
  assign n533 = x7 & n92 ;
  assign n536 = n535 ^ n533 ;
  assign n537 = n536 ^ x7 ;
  assign n531 = x7 & n102 ;
  assign n532 = n531 ^ x7 ;
  assign n538 = n537 ^ n532 ;
  assign n529 = x7 & ~n61 ;
  assign n530 = n80 & n529 ;
  assign n539 = n538 ^ n530 ;
  assign n524 = x15 & ~n53 ;
  assign n525 = n87 & n524 ;
  assign n523 = x15 & n92 ;
  assign n526 = n525 ^ n523 ;
  assign n521 = x15 & n102 ;
  assign n522 = n521 ^ x15 ;
  assign n527 = n526 ^ n522 ;
  assign n519 = x15 & ~n61 ;
  assign n520 = n80 & n519 ;
  assign n528 = n527 ^ n520 ;
  assign n540 = n539 ^ n528 ;
  assign n515 = x31 & ~n159 ;
  assign n516 = n146 & n515 ;
  assign n512 = x31 & n169 ;
  assign n513 = n512 ^ x31 ;
  assign n508 = x31 & ~n151 ;
  assign n509 = n182 & n508 ;
  assign n507 = x31 & n175 ;
  assign n510 = n509 ^ n507 ;
  assign n511 = n510 ^ x31 ;
  assign n514 = n513 ^ n511 ;
  assign n517 = n516 ^ n514 ;
  assign n504 = x23 & ~n159 ;
  assign n505 = n146 & n504 ;
  assign n500 = x23 & ~n151 ;
  assign n501 = n182 & n500 ;
  assign n499 = x23 & n175 ;
  assign n502 = n501 ^ n499 ;
  assign n497 = x23 & n169 ;
  assign n498 = n497 ^ x23 ;
  assign n503 = n502 ^ n498 ;
  assign n506 = n505 ^ n503 ;
  assign n518 = n517 ^ n506 ;
  assign n541 = n540 ^ n518 ;
  assign n542 = n496 & n541 ;
  assign n543 = n542 ^ n496 ;
  assign n544 = n543 ^ n541 ;
  assign n545 = n451 & n544 ;
  assign n546 = n545 ^ n451 ;
  assign n547 = n546 ^ n544 ;
  assign n548 = ~n358 & ~n547 ;
  assign n620 = n271 & n548 ;
  assign n621 = n620 ^ n271 ;
  assign n1394 = n1393 ^ n621 ;
  assign n560 = n518 & n540 ;
  assign n561 = n560 ^ n540 ;
  assign n562 = n496 & n561 ;
  assign n563 = n562 ^ n561 ;
  assign n558 = n473 & n495 ;
  assign n559 = n558 ^ n473 ;
  assign n564 = n563 ^ n559 ;
  assign n565 = n451 & n564 ;
  assign n566 = n565 ^ n564 ;
  assign n553 = n425 & n447 ;
  assign n554 = n553 ^ n425 ;
  assign n555 = n403 & n554 ;
  assign n556 = n555 ^ n554 ;
  assign n552 = n380 & ~n402 ;
  assign n557 = n556 ^ n552 ;
  assign n567 = n566 ^ n557 ;
  assign n623 = n271 & ~n358 ;
  assign n624 = n567 & n623 ;
  assign n1395 = n1394 ^ n624 ;
  assign n1388 = n248 & n293 ;
  assign n627 = n293 & ~n348 ;
  assign n628 = n344 & n627 ;
  assign n1389 = n1388 ^ n628 ;
  assign n630 = n293 & n548 ;
  assign n631 = n630 ^ n293 ;
  assign n1390 = n1389 ^ n631 ;
  assign n633 = n293 & ~n358 ;
  assign n634 = n567 & n633 ;
  assign n1391 = n1390 ^ n634 ;
  assign n1396 = n1395 ^ n1391 ;
  assign n902 = x42 ^ x34 ;
  assign n928 = x35 & x43 ;
  assign n929 = n928 ^ x35 ;
  assign n930 = n902 & n929 ;
  assign n931 = n930 ^ n929 ;
  assign n927 = x34 & ~x42 ;
  assign n932 = n931 ^ n927 ;
  assign n897 = x40 ^ x32 ;
  assign n898 = x41 ^ x33 ;
  assign n899 = n897 & n898 ;
  assign n900 = n899 ^ n897 ;
  assign n901 = n900 ^ n898 ;
  assign n1119 = x42 & ~n901 ;
  assign n1120 = n932 & n1119 ;
  assign n923 = x33 & ~x41 ;
  assign n924 = ~n897 & n923 ;
  assign n922 = x32 & ~x40 ;
  assign n925 = n924 ^ n922 ;
  assign n1118 = x42 & ~n925 ;
  assign n1121 = n1120 ^ n1118 ;
  assign n903 = x43 ^ x35 ;
  assign n904 = n902 & n903 ;
  assign n905 = n904 ^ n902 ;
  assign n906 = n905 ^ n903 ;
  assign n907 = n901 & n906 ;
  assign n908 = n907 ^ n901 ;
  assign n909 = n908 ^ n906 ;
  assign n879 = x44 ^ x36 ;
  assign n883 = x45 ^ x37 ;
  assign n884 = n879 & n883 ;
  assign n885 = n884 ^ n879 ;
  assign n886 = n885 ^ n883 ;
  assign n888 = x46 ^ x38 ;
  assign n912 = x47 ^ x39 ;
  assign n913 = n888 & n912 ;
  assign n914 = n913 ^ n888 ;
  assign n915 = n914 ^ n912 ;
  assign n916 = n886 & n915 ;
  assign n917 = n916 ^ n886 ;
  assign n918 = n917 ^ n915 ;
  assign n919 = ~n909 & ~n918 ;
  assign n1116 = x42 & n919 ;
  assign n1117 = n1116 ^ x42 ;
  assign n1122 = n1121 ^ n1117 ;
  assign n889 = x39 & x47 ;
  assign n890 = n889 ^ x39 ;
  assign n891 = n888 & n890 ;
  assign n892 = n891 ^ n890 ;
  assign n887 = x38 & ~x46 ;
  assign n893 = n892 ^ n887 ;
  assign n894 = n886 & n893 ;
  assign n895 = n894 ^ n893 ;
  assign n880 = x37 & ~x45 ;
  assign n881 = ~n879 & n880 ;
  assign n878 = x36 & ~x44 ;
  assign n882 = n881 ^ n878 ;
  assign n896 = n895 ^ n882 ;
  assign n1114 = x42 & ~n909 ;
  assign n1115 = n896 & n1114 ;
  assign n1123 = n1122 ^ n1115 ;
  assign n1108 = x34 & ~n901 ;
  assign n1109 = n932 & n1108 ;
  assign n1107 = x34 & ~n925 ;
  assign n1110 = n1109 ^ n1107 ;
  assign n1105 = x34 & n919 ;
  assign n1106 = n1105 ^ x34 ;
  assign n1111 = n1110 ^ n1106 ;
  assign n1103 = x34 & ~n909 ;
  assign n1104 = n896 & n1103 ;
  assign n1112 = n1111 ^ n1104 ;
  assign n1113 = n1112 ^ x34 ;
  assign n1124 = n1123 ^ n1113 ;
  assign n1101 = n292 ^ x26 ;
  assign n1102 = n1101 ^ n281 ;
  assign n1125 = n1124 ^ n1102 ;
  assign n1126 = n338 ^ x27 ;
  assign n1127 = n1126 ^ n327 ;
  assign n1144 = x43 & ~n901 ;
  assign n1145 = n932 & n1144 ;
  assign n1143 = x43 & ~n925 ;
  assign n1146 = n1145 ^ n1143 ;
  assign n1141 = x43 & n919 ;
  assign n1142 = n1141 ^ x43 ;
  assign n1147 = n1146 ^ n1142 ;
  assign n1139 = x43 & ~n909 ;
  assign n1140 = n896 & n1139 ;
  assign n1148 = n1147 ^ n1140 ;
  assign n1133 = x35 & ~n901 ;
  assign n1134 = n932 & n1133 ;
  assign n1132 = x35 & ~n925 ;
  assign n1135 = n1134 ^ n1132 ;
  assign n1130 = x35 & n919 ;
  assign n1131 = n1130 ^ x35 ;
  assign n1136 = n1135 ^ n1131 ;
  assign n1128 = x35 & ~n909 ;
  assign n1129 = n896 & n1128 ;
  assign n1137 = n1136 ^ n1129 ;
  assign n1138 = n1137 ^ x35 ;
  assign n1149 = n1148 ^ n1138 ;
  assign n1175 = n1127 & n1149 ;
  assign n1176 = n1175 ^ n1127 ;
  assign n1177 = n1125 & n1176 ;
  assign n1178 = n1177 ^ n1176 ;
  assign n1174 = n1102 & ~n1124 ;
  assign n1179 = n1178 ^ n1174 ;
  assign n1066 = x40 & ~n901 ;
  assign n1067 = n932 & n1066 ;
  assign n1065 = x40 & ~n925 ;
  assign n1068 = n1067 ^ n1065 ;
  assign n1063 = x40 & n919 ;
  assign n1064 = n1063 ^ x40 ;
  assign n1069 = n1068 ^ n1064 ;
  assign n1061 = x40 & ~n909 ;
  assign n1062 = n896 & n1061 ;
  assign n1070 = n1069 ^ n1062 ;
  assign n1055 = x32 & ~n901 ;
  assign n1056 = n932 & n1055 ;
  assign n1054 = x32 & ~n925 ;
  assign n1057 = n1056 ^ n1054 ;
  assign n1052 = x32 & n919 ;
  assign n1053 = n1052 ^ x32 ;
  assign n1058 = n1057 ^ n1053 ;
  assign n1050 = x32 & ~n909 ;
  assign n1051 = n896 & n1050 ;
  assign n1059 = n1058 ^ n1051 ;
  assign n1060 = n1059 ^ x32 ;
  assign n1071 = n1070 ^ n1060 ;
  assign n1048 = n198 ^ x24 ;
  assign n1049 = n1048 ^ n187 ;
  assign n1072 = n1071 ^ n1049 ;
  assign n1091 = x41 & ~n901 ;
  assign n1092 = n932 & n1091 ;
  assign n1090 = x41 & ~n925 ;
  assign n1093 = n1092 ^ n1090 ;
  assign n1088 = x41 & n919 ;
  assign n1089 = n1088 ^ x41 ;
  assign n1094 = n1093 ^ n1089 ;
  assign n1086 = x41 & ~n909 ;
  assign n1087 = n896 & n1086 ;
  assign n1095 = n1094 ^ n1087 ;
  assign n1080 = x33 & ~n901 ;
  assign n1081 = n932 & n1080 ;
  assign n1079 = x33 & ~n925 ;
  assign n1082 = n1081 ^ n1079 ;
  assign n1077 = x33 & n919 ;
  assign n1078 = n1077 ^ x33 ;
  assign n1083 = n1082 ^ n1078 ;
  assign n1075 = x33 & ~n909 ;
  assign n1076 = n896 & n1075 ;
  assign n1084 = n1083 ^ n1076 ;
  assign n1085 = n1084 ^ x33 ;
  assign n1096 = n1095 ^ n1085 ;
  assign n1073 = n222 ^ x25 ;
  assign n1074 = n1073 ^ n211 ;
  assign n1097 = n1096 ^ n1074 ;
  assign n1098 = n1072 & n1097 ;
  assign n1099 = n1098 ^ n1072 ;
  assign n1100 = n1099 ^ n1097 ;
  assign n1382 = ~n1100 & n1124 ;
  assign n1383 = n1179 & n1382 ;
  assign n1170 = n1074 & ~n1096 ;
  assign n1171 = ~n1072 & n1170 ;
  assign n1169 = n1049 & ~n1071 ;
  assign n1172 = n1171 ^ n1169 ;
  assign n1381 = n1124 & ~n1172 ;
  assign n1384 = n1383 ^ n1381 ;
  assign n1150 = n1149 ^ n1127 ;
  assign n1151 = n1125 & n1150 ;
  assign n1152 = n1151 ^ n1125 ;
  assign n1153 = n1152 ^ n1150 ;
  assign n1154 = n1100 & n1153 ;
  assign n1155 = n1154 ^ n1100 ;
  assign n1156 = n1155 ^ n1153 ;
  assign n944 = x44 & ~n901 ;
  assign n945 = n932 & n944 ;
  assign n943 = x44 & ~n925 ;
  assign n946 = n945 ^ n943 ;
  assign n941 = x44 & n919 ;
  assign n942 = n941 ^ x44 ;
  assign n947 = n946 ^ n942 ;
  assign n939 = x44 & ~n909 ;
  assign n940 = n896 & n939 ;
  assign n948 = n947 ^ n940 ;
  assign n933 = x36 & ~n901 ;
  assign n934 = n932 & n933 ;
  assign n926 = x36 & ~n925 ;
  assign n935 = n934 ^ n926 ;
  assign n920 = x36 & n919 ;
  assign n921 = n920 ^ x36 ;
  assign n936 = n935 ^ n921 ;
  assign n910 = x36 & ~n909 ;
  assign n911 = n896 & n910 ;
  assign n937 = n936 ^ n911 ;
  assign n938 = n937 ^ x36 ;
  assign n949 = n948 ^ n938 ;
  assign n876 = n401 ^ x28 ;
  assign n877 = n876 ^ n390 ;
  assign n951 = n949 ^ n877 ;
  assign n970 = x45 & ~n901 ;
  assign n971 = n932 & n970 ;
  assign n969 = x45 & ~n925 ;
  assign n972 = n971 ^ n969 ;
  assign n967 = x45 & n919 ;
  assign n968 = n967 ^ x45 ;
  assign n973 = n972 ^ n968 ;
  assign n965 = x45 & ~n909 ;
  assign n966 = n896 & n965 ;
  assign n974 = n973 ^ n966 ;
  assign n959 = x37 & ~n901 ;
  assign n960 = n932 & n959 ;
  assign n958 = x37 & ~n925 ;
  assign n961 = n960 ^ n958 ;
  assign n956 = x37 & n919 ;
  assign n957 = n956 ^ x37 ;
  assign n962 = n961 ^ n957 ;
  assign n954 = x37 & ~n909 ;
  assign n955 = n896 & n954 ;
  assign n963 = n962 ^ n955 ;
  assign n964 = n963 ^ x37 ;
  assign n975 = n974 ^ n964 ;
  assign n952 = n446 ^ x29 ;
  assign n953 = n952 ^ n435 ;
  assign n981 = n975 ^ n953 ;
  assign n982 = n951 & n981 ;
  assign n983 = n982 ^ n951 ;
  assign n984 = n983 ^ n981 ;
  assign n1003 = x46 & ~n901 ;
  assign n1004 = n932 & n1003 ;
  assign n1002 = x46 & ~n925 ;
  assign n1005 = n1004 ^ n1002 ;
  assign n1000 = x46 & n919 ;
  assign n1001 = n1000 ^ x46 ;
  assign n1006 = n1005 ^ n1001 ;
  assign n998 = x46 & ~n909 ;
  assign n999 = n896 & n998 ;
  assign n1007 = n1006 ^ n999 ;
  assign n992 = x38 & ~n901 ;
  assign n993 = n932 & n992 ;
  assign n991 = x38 & ~n925 ;
  assign n994 = n993 ^ n991 ;
  assign n989 = x38 & n919 ;
  assign n990 = n989 ^ x38 ;
  assign n995 = n994 ^ n990 ;
  assign n987 = x38 & ~n909 ;
  assign n988 = n896 & n987 ;
  assign n996 = n995 ^ n988 ;
  assign n997 = n996 ^ x38 ;
  assign n1008 = n1007 ^ n997 ;
  assign n985 = n494 ^ x30 ;
  assign n986 = n985 ^ n483 ;
  assign n1011 = n1008 ^ n986 ;
  assign n1033 = x47 & ~n901 ;
  assign n1034 = n932 & n1033 ;
  assign n1032 = x47 & n925 ;
  assign n1035 = n1034 ^ n1032 ;
  assign n1036 = n1035 ^ x47 ;
  assign n1030 = x47 & n919 ;
  assign n1031 = n1030 ^ x47 ;
  assign n1037 = n1036 ^ n1031 ;
  assign n1028 = x47 & ~n909 ;
  assign n1029 = n896 & n1028 ;
  assign n1038 = n1037 ^ n1029 ;
  assign n1023 = x39 & ~n901 ;
  assign n1024 = n932 & n1023 ;
  assign n1022 = x39 & n925 ;
  assign n1025 = n1024 ^ n1022 ;
  assign n1020 = x39 & n919 ;
  assign n1021 = n1020 ^ x39 ;
  assign n1026 = n1025 ^ n1021 ;
  assign n1018 = x39 & ~n909 ;
  assign n1019 = n896 & n1018 ;
  assign n1027 = n1026 ^ n1019 ;
  assign n1039 = n1038 ^ n1027 ;
  assign n1014 = n502 ^ x23 ;
  assign n1015 = n1014 ^ n498 ;
  assign n1016 = n1015 ^ n505 ;
  assign n1012 = n513 ^ n510 ;
  assign n1013 = n1012 ^ n516 ;
  assign n1017 = n1016 ^ n1013 ;
  assign n1159 = n1039 ^ n1017 ;
  assign n1160 = n1011 & n1159 ;
  assign n1161 = n1160 ^ n1011 ;
  assign n1162 = n1161 ^ n1159 ;
  assign n1163 = n984 & n1162 ;
  assign n1164 = n1163 ^ n984 ;
  assign n1165 = n1164 ^ n1162 ;
  assign n1166 = ~n1156 & ~n1165 ;
  assign n1379 = n1124 & n1166 ;
  assign n1380 = n1379 ^ n1124 ;
  assign n1385 = n1384 ^ n1380 ;
  assign n1040 = n1017 & n1039 ;
  assign n1041 = n1040 ^ n1017 ;
  assign n1042 = n1011 & n1041 ;
  assign n1043 = n1042 ^ n1041 ;
  assign n1009 = n986 & n1008 ;
  assign n1010 = n1009 ^ n986 ;
  assign n1044 = n1043 ^ n1010 ;
  assign n1045 = n984 & n1044 ;
  assign n1046 = n1045 ^ n1044 ;
  assign n976 = n953 & n975 ;
  assign n977 = n976 ^ n953 ;
  assign n978 = n951 & n977 ;
  assign n979 = n978 ^ n977 ;
  assign n950 = n877 & ~n949 ;
  assign n980 = n979 ^ n950 ;
  assign n1047 = n1046 ^ n980 ;
  assign n1377 = n1124 & ~n1156 ;
  assign n1378 = n1047 & n1377 ;
  assign n1386 = n1385 ^ n1378 ;
  assign n1372 = ~n1100 & n1102 ;
  assign n1373 = n1179 & n1372 ;
  assign n1371 = n1102 & n1172 ;
  assign n1374 = n1373 ^ n1371 ;
  assign n1369 = n1102 & n1166 ;
  assign n1370 = n1369 ^ n1102 ;
  assign n1375 = n1374 ^ n1370 ;
  assign n1367 = n1102 & ~n1156 ;
  assign n1368 = n1047 & n1367 ;
  assign n1376 = n1375 ^ n1368 ;
  assign n1387 = n1386 ^ n1376 ;
  assign n1397 = n1396 ^ n1387 ;
  assign n1402 = ~n248 & n317 ;
  assign n642 = n317 & ~n348 ;
  assign n643 = n344 & n642 ;
  assign n1403 = n1402 ^ n643 ;
  assign n645 = n317 & n548 ;
  assign n646 = n645 ^ n317 ;
  assign n1404 = n1403 ^ n646 ;
  assign n648 = n317 & ~n358 ;
  assign n649 = n567 & n648 ;
  assign n1405 = n1404 ^ n649 ;
  assign n1398 = n248 & n339 ;
  assign n652 = n339 & ~n348 ;
  assign n653 = n344 & n652 ;
  assign n1399 = n1398 ^ n653 ;
  assign n655 = n339 & n548 ;
  assign n656 = n655 ^ n339 ;
  assign n1400 = n1399 ^ n656 ;
  assign n658 = n339 & ~n358 ;
  assign n659 = n567 & n658 ;
  assign n1401 = n1400 ^ n659 ;
  assign n1406 = n1405 ^ n1401 ;
  assign n1422 = ~n1100 & n1149 ;
  assign n1423 = n1179 & n1422 ;
  assign n1421 = n1149 & ~n1172 ;
  assign n1424 = n1423 ^ n1421 ;
  assign n1419 = n1149 & n1166 ;
  assign n1420 = n1419 ^ n1149 ;
  assign n1425 = n1424 ^ n1420 ;
  assign n1417 = n1149 & ~n1156 ;
  assign n1418 = n1047 & n1417 ;
  assign n1426 = n1425 ^ n1418 ;
  assign n1412 = ~n1100 & n1127 ;
  assign n1413 = n1179 & n1412 ;
  assign n1411 = n1127 & n1172 ;
  assign n1414 = n1413 ^ n1411 ;
  assign n1409 = n1127 & n1166 ;
  assign n1410 = n1409 ^ n1127 ;
  assign n1415 = n1414 ^ n1410 ;
  assign n1407 = n1127 & ~n1156 ;
  assign n1408 = n1047 & n1407 ;
  assign n1416 = n1415 ^ n1408 ;
  assign n1427 = n1426 ^ n1416 ;
  assign n1449 = n1406 & n1427 ;
  assign n1450 = n1449 ^ n1406 ;
  assign n1451 = n1397 & n1450 ;
  assign n1452 = n1451 ^ n1450 ;
  assign n1448 = ~n1387 & n1396 ;
  assign n1453 = n1452 ^ n1448 ;
  assign n1326 = n1071 & ~n1100 ;
  assign n1327 = n1179 & n1326 ;
  assign n1325 = n1071 & ~n1172 ;
  assign n1328 = n1327 ^ n1325 ;
  assign n1323 = n1071 & n1166 ;
  assign n1324 = n1323 ^ n1071 ;
  assign n1329 = n1328 ^ n1324 ;
  assign n1321 = n1071 & ~n1156 ;
  assign n1322 = n1047 & n1321 ;
  assign n1330 = n1329 ^ n1322 ;
  assign n1316 = n1049 & ~n1100 ;
  assign n1317 = n1179 & n1316 ;
  assign n1315 = n1049 & n1172 ;
  assign n1318 = n1317 ^ n1315 ;
  assign n1313 = n1049 & n1166 ;
  assign n1314 = n1313 ^ n1049 ;
  assign n1319 = n1318 ^ n1314 ;
  assign n1311 = n1049 & ~n1156 ;
  assign n1312 = n1047 & n1311 ;
  assign n1320 = n1319 ^ n1312 ;
  assign n1331 = n1330 ^ n1320 ;
  assign n1306 = n127 & ~n248 ;
  assign n349 = n127 & ~n348 ;
  assign n350 = n344 & n349 ;
  assign n1307 = n1306 ^ n350 ;
  assign n549 = n127 & n548 ;
  assign n550 = n549 ^ n127 ;
  assign n1308 = n1307 ^ n550 ;
  assign n568 = n127 & ~n358 ;
  assign n569 = n567 & n568 ;
  assign n1309 = n1308 ^ n569 ;
  assign n1302 = n199 & n248 ;
  assign n572 = n199 & ~n348 ;
  assign n573 = n344 & n572 ;
  assign n1303 = n1302 ^ n573 ;
  assign n575 = n199 & n548 ;
  assign n576 = n575 ^ n199 ;
  assign n1304 = n1303 ^ n576 ;
  assign n578 = n199 & ~n358 ;
  assign n579 = n567 & n578 ;
  assign n1305 = n1304 ^ n579 ;
  assign n1310 = n1309 ^ n1305 ;
  assign n1332 = n1331 ^ n1310 ;
  assign n1358 = n245 & ~n248 ;
  assign n585 = n245 & ~n348 ;
  assign n586 = n344 & n585 ;
  assign n1359 = n1358 ^ n586 ;
  assign n588 = n245 & n548 ;
  assign n589 = n588 ^ n245 ;
  assign n1360 = n1359 ^ n589 ;
  assign n591 = n245 & ~n358 ;
  assign n592 = n567 & n591 ;
  assign n1361 = n1360 ^ n592 ;
  assign n1354 = n223 & n248 ;
  assign n595 = n223 & ~n348 ;
  assign n596 = n344 & n595 ;
  assign n1355 = n1354 ^ n596 ;
  assign n598 = n223 & n548 ;
  assign n599 = n598 ^ n223 ;
  assign n1356 = n1355 ^ n599 ;
  assign n601 = n223 & ~n358 ;
  assign n602 = n567 & n601 ;
  assign n1357 = n1356 ^ n602 ;
  assign n1362 = n1361 ^ n1357 ;
  assign n1348 = n1096 & ~n1100 ;
  assign n1349 = n1179 & n1348 ;
  assign n1347 = n1096 & ~n1172 ;
  assign n1350 = n1349 ^ n1347 ;
  assign n1345 = n1096 & n1166 ;
  assign n1346 = n1345 ^ n1096 ;
  assign n1351 = n1350 ^ n1346 ;
  assign n1343 = n1096 & ~n1156 ;
  assign n1344 = n1047 & n1343 ;
  assign n1352 = n1351 ^ n1344 ;
  assign n1338 = n1074 & ~n1100 ;
  assign n1339 = n1179 & n1338 ;
  assign n1337 = n1074 & n1172 ;
  assign n1340 = n1339 ^ n1337 ;
  assign n1335 = n1074 & n1166 ;
  assign n1336 = n1335 ^ n1074 ;
  assign n1341 = n1340 ^ n1336 ;
  assign n1333 = n1074 & ~n1156 ;
  assign n1334 = n1047 & n1333 ;
  assign n1342 = n1341 ^ n1334 ;
  assign n1353 = n1352 ^ n1342 ;
  assign n1363 = n1362 ^ n1353 ;
  assign n1364 = n1332 & n1363 ;
  assign n1365 = n1364 ^ n1332 ;
  assign n1366 = n1365 ^ n1363 ;
  assign n1585 = n1331 & ~n1366 ;
  assign n1586 = n1453 & n1585 ;
  assign n1444 = ~n1353 & n1362 ;
  assign n1445 = ~n1332 & n1444 ;
  assign n1443 = n1310 & ~n1331 ;
  assign n1446 = n1445 ^ n1443 ;
  assign n1584 = n1331 & n1446 ;
  assign n1587 = n1586 ^ n1584 ;
  assign n1588 = n1587 ^ n1331 ;
  assign n1428 = n1427 ^ n1406 ;
  assign n1429 = n1397 & n1428 ;
  assign n1430 = n1429 ^ n1397 ;
  assign n1431 = n1430 ^ n1428 ;
  assign n1432 = ~n1366 & ~n1431 ;
  assign n1190 = n949 & ~n1100 ;
  assign n1191 = n1179 & n1190 ;
  assign n1189 = n949 & ~n1172 ;
  assign n1192 = n1191 ^ n1189 ;
  assign n1187 = n949 & n1166 ;
  assign n1188 = n1187 ^ n949 ;
  assign n1193 = n1192 ^ n1188 ;
  assign n1185 = n949 & ~n1156 ;
  assign n1186 = n1047 & n1185 ;
  assign n1194 = n1193 ^ n1186 ;
  assign n1180 = n877 & ~n1100 ;
  assign n1181 = n1179 & n1180 ;
  assign n1173 = n877 & n1172 ;
  assign n1182 = n1181 ^ n1173 ;
  assign n1167 = n877 & n1166 ;
  assign n1168 = n1167 ^ n877 ;
  assign n1183 = n1182 ^ n1168 ;
  assign n1157 = n877 & ~n1156 ;
  assign n1158 = n1047 & n1157 ;
  assign n1184 = n1183 ^ n1158 ;
  assign n1195 = n1194 ^ n1184 ;
  assign n871 = ~n248 & n380 ;
  assign n677 = ~n348 & n380 ;
  assign n678 = n344 & n677 ;
  assign n872 = n871 ^ n678 ;
  assign n680 = n380 & n548 ;
  assign n681 = n680 ^ n380 ;
  assign n873 = n872 ^ n681 ;
  assign n683 = ~n358 & n380 ;
  assign n684 = n567 & n683 ;
  assign n874 = n873 ^ n684 ;
  assign n867 = n248 & n402 ;
  assign n687 = ~n348 & n402 ;
  assign n688 = n344 & n687 ;
  assign n868 = n867 ^ n688 ;
  assign n690 = n402 & n548 ;
  assign n691 = n690 ^ n402 ;
  assign n869 = n868 ^ n691 ;
  assign n693 = ~n358 & n402 ;
  assign n694 = n567 & n693 ;
  assign n870 = n869 ^ n694 ;
  assign n875 = n874 ^ n870 ;
  assign n1197 = n1195 ^ n875 ;
  assign n1222 = n975 & ~n1100 ;
  assign n1223 = n1179 & n1222 ;
  assign n1221 = n975 & ~n1172 ;
  assign n1224 = n1223 ^ n1221 ;
  assign n1219 = n975 & n1166 ;
  assign n1220 = n1219 ^ n975 ;
  assign n1225 = n1224 ^ n1220 ;
  assign n1217 = n975 & ~n1156 ;
  assign n1218 = n1047 & n1217 ;
  assign n1226 = n1225 ^ n1218 ;
  assign n1212 = n953 & ~n1100 ;
  assign n1213 = n1179 & n1212 ;
  assign n1211 = n953 & n1172 ;
  assign n1214 = n1213 ^ n1211 ;
  assign n1209 = n953 & n1166 ;
  assign n1210 = n1209 ^ n953 ;
  assign n1215 = n1214 ^ n1210 ;
  assign n1207 = n953 & ~n1156 ;
  assign n1208 = n1047 & n1207 ;
  assign n1216 = n1215 ^ n1208 ;
  assign n1227 = n1226 ^ n1216 ;
  assign n1202 = ~n248 & n425 ;
  assign n702 = ~n348 & n425 ;
  assign n703 = n344 & n702 ;
  assign n1203 = n1202 ^ n703 ;
  assign n705 = n425 & n548 ;
  assign n706 = n705 ^ n425 ;
  assign n1204 = n1203 ^ n706 ;
  assign n708 = ~n358 & n425 ;
  assign n709 = n567 & n708 ;
  assign n1205 = n1204 ^ n709 ;
  assign n1198 = n248 & n447 ;
  assign n712 = ~n348 & n447 ;
  assign n713 = n344 & n712 ;
  assign n1199 = n1198 ^ n713 ;
  assign n715 = n447 & n548 ;
  assign n716 = n715 ^ n447 ;
  assign n1200 = n1199 ^ n716 ;
  assign n718 = ~n358 & n447 ;
  assign n719 = n567 & n718 ;
  assign n1201 = n1200 ^ n719 ;
  assign n1206 = n1205 ^ n1201 ;
  assign n1231 = n1227 ^ n1206 ;
  assign n1232 = n1197 & n1231 ;
  assign n1233 = n1232 ^ n1197 ;
  assign n1234 = n1233 ^ n1231 ;
  assign n1259 = n1008 & ~n1100 ;
  assign n1260 = n1179 & n1259 ;
  assign n1258 = n1008 & ~n1172 ;
  assign n1261 = n1260 ^ n1258 ;
  assign n1256 = n1008 & n1166 ;
  assign n1257 = n1256 ^ n1008 ;
  assign n1262 = n1261 ^ n1257 ;
  assign n1254 = n1008 & ~n1156 ;
  assign n1255 = n1047 & n1254 ;
  assign n1263 = n1262 ^ n1255 ;
  assign n1249 = n986 & ~n1100 ;
  assign n1250 = n1179 & n1249 ;
  assign n1248 = n986 & n1172 ;
  assign n1251 = n1250 ^ n1248 ;
  assign n1246 = n986 & n1166 ;
  assign n1247 = n1246 ^ n986 ;
  assign n1252 = n1251 ^ n1247 ;
  assign n1244 = n986 & ~n1156 ;
  assign n1245 = n1047 & n1244 ;
  assign n1253 = n1252 ^ n1245 ;
  assign n1264 = n1263 ^ n1253 ;
  assign n1239 = ~n248 & n473 ;
  assign n817 = ~n348 & n473 ;
  assign n818 = n344 & n817 ;
  assign n1240 = n1239 ^ n818 ;
  assign n778 = n473 & n548 ;
  assign n779 = n778 ^ n473 ;
  assign n1241 = n1240 ^ n779 ;
  assign n775 = ~n358 & n473 ;
  assign n821 = n567 & n775 ;
  assign n1242 = n1241 ^ n821 ;
  assign n1235 = n248 & n495 ;
  assign n824 = ~n348 & n495 ;
  assign n825 = n344 & n824 ;
  assign n1236 = n1235 ^ n825 ;
  assign n791 = n495 & n548 ;
  assign n792 = n791 ^ n495 ;
  assign n1237 = n1236 ^ n792 ;
  assign n788 = ~n358 & n495 ;
  assign n828 = n567 & n788 ;
  assign n1238 = n1237 ^ n828 ;
  assign n1243 = n1242 ^ n1238 ;
  assign n1266 = n1264 ^ n1243 ;
  assign n1289 = n1039 & ~n1100 ;
  assign n1290 = n1179 & n1289 ;
  assign n1288 = n1039 & ~n1172 ;
  assign n1291 = n1290 ^ n1288 ;
  assign n1286 = n1039 & n1166 ;
  assign n1287 = n1286 ^ n1039 ;
  assign n1292 = n1291 ^ n1287 ;
  assign n1284 = n1039 & ~n1156 ;
  assign n1285 = n1047 & n1284 ;
  assign n1293 = n1292 ^ n1285 ;
  assign n1278 = n1017 & ~n1100 ;
  assign n1279 = n1179 & n1278 ;
  assign n1277 = n1017 & ~n1172 ;
  assign n1280 = n1279 ^ n1277 ;
  assign n1275 = n1017 & n1166 ;
  assign n1276 = n1275 ^ n1017 ;
  assign n1281 = n1280 ^ n1276 ;
  assign n1273 = n1017 & ~n1156 ;
  assign n1274 = n1047 & n1273 ;
  assign n1282 = n1281 ^ n1274 ;
  assign n1283 = n1282 ^ n1017 ;
  assign n1294 = n1293 ^ n1283 ;
  assign n1268 = ~n248 & n540 ;
  assign n833 = ~n348 & n540 ;
  assign n834 = n344 & n833 ;
  assign n1269 = n1268 ^ n834 ;
  assign n836 = n540 & n548 ;
  assign n837 = n836 ^ n540 ;
  assign n1270 = n1269 ^ n837 ;
  assign n839 = ~n358 & n540 ;
  assign n840 = n567 & n839 ;
  assign n1271 = n1270 ^ n840 ;
  assign n847 = ~n348 & n518 ;
  assign n848 = n344 & n847 ;
  assign n846 = ~n248 & n518 ;
  assign n849 = n848 ^ n846 ;
  assign n844 = n518 & n548 ;
  assign n845 = n844 ^ n518 ;
  assign n850 = n849 ^ n845 ;
  assign n842 = ~n358 & n518 ;
  assign n843 = n567 & n842 ;
  assign n851 = n850 ^ n843 ;
  assign n1267 = n851 ^ n518 ;
  assign n1272 = n1271 ^ n1267 ;
  assign n1435 = n1294 ^ n1272 ;
  assign n1436 = n1266 & n1435 ;
  assign n1437 = n1436 ^ n1266 ;
  assign n1438 = n1437 ^ n1435 ;
  assign n1439 = ~n1234 & ~n1438 ;
  assign n1440 = n1432 & n1439 ;
  assign n1582 = n1331 & n1440 ;
  assign n1583 = n1582 ^ n1331 ;
  assign n1589 = n1588 ^ n1583 ;
  assign n1295 = n1272 & n1294 ;
  assign n1296 = n1295 ^ n1272 ;
  assign n1297 = n1266 & n1296 ;
  assign n1298 = n1297 ^ n1296 ;
  assign n1265 = n1243 & ~n1264 ;
  assign n1299 = n1298 ^ n1265 ;
  assign n1300 = ~n1234 & n1299 ;
  assign n1228 = n1206 & ~n1227 ;
  assign n1229 = ~n1197 & n1228 ;
  assign n1196 = n875 & ~n1195 ;
  assign n1230 = n1229 ^ n1196 ;
  assign n1301 = n1300 ^ n1230 ;
  assign n1580 = n1331 & n1432 ;
  assign n1581 = n1301 & n1580 ;
  assign n1590 = n1589 ^ n1581 ;
  assign n1575 = n1310 & ~n1366 ;
  assign n1576 = n1453 & n1575 ;
  assign n1574 = n1310 & n1446 ;
  assign n1577 = n1576 ^ n1574 ;
  assign n1572 = n1310 & n1440 ;
  assign n1573 = n1572 ^ n1310 ;
  assign n1578 = n1577 ^ n1573 ;
  assign n1570 = n1310 & n1432 ;
  assign n1571 = n1301 & n1570 ;
  assign n1579 = n1578 ^ n1571 ;
  assign n1591 = n1590 ^ n1579 ;
  assign n88 = ~n53 & n87 ;
  assign n93 = n92 ^ n88 ;
  assign n81 = ~n61 & n80 ;
  assign n94 = n93 ^ n81 ;
  assign n103 = n102 ^ n94 ;
  assign n104 = x0 & ~n103 ;
  assign n115 = n114 ^ n104 ;
  assign n571 = n199 & ~n248 ;
  assign n574 = n573 ^ n571 ;
  assign n577 = n576 ^ n574 ;
  assign n580 = n579 ^ n577 ;
  assign n249 = n127 & n248 ;
  assign n351 = n350 ^ n249 ;
  assign n551 = n550 ^ n351 ;
  assign n570 = n569 ^ n551 ;
  assign n581 = n580 ^ n570 ;
  assign n583 = n581 ^ n115 ;
  assign n605 = x1 & ~n103 ;
  assign n606 = n605 ^ n233 ;
  assign n594 = n223 & ~n248 ;
  assign n597 = n596 ^ n594 ;
  assign n600 = n599 ^ n597 ;
  assign n603 = n602 ^ n600 ;
  assign n584 = n245 & n248 ;
  assign n587 = n586 ^ n584 ;
  assign n590 = n589 ^ n587 ;
  assign n593 = n592 ^ n590 ;
  assign n604 = n603 ^ n593 ;
  assign n610 = n606 ^ n604 ;
  assign n611 = n583 & n610 ;
  assign n612 = n611 ^ n583 ;
  assign n613 = n612 ^ n610 ;
  assign n626 = ~n248 & n293 ;
  assign n629 = n628 ^ n626 ;
  assign n632 = n631 ^ n629 ;
  assign n635 = n634 ^ n632 ;
  assign n616 = n248 & n271 ;
  assign n619 = n618 ^ n616 ;
  assign n622 = n621 ^ n619 ;
  assign n625 = n624 ^ n622 ;
  assign n636 = n635 ^ n625 ;
  assign n614 = x2 & ~n103 ;
  assign n615 = n614 ^ n259 ;
  assign n638 = n636 ^ n615 ;
  assign n651 = ~n248 & n339 ;
  assign n654 = n653 ^ n651 ;
  assign n657 = n656 ^ n654 ;
  assign n660 = n659 ^ n657 ;
  assign n641 = n248 & n317 ;
  assign n644 = n643 ^ n641 ;
  assign n647 = n646 ^ n644 ;
  assign n650 = n649 ^ n647 ;
  assign n661 = n660 ^ n650 ;
  assign n639 = x3 & ~n103 ;
  assign n640 = n639 ^ n305 ;
  assign n669 = n661 ^ n640 ;
  assign n670 = n638 & n669 ;
  assign n671 = n670 ^ n638 ;
  assign n672 = n671 ^ n669 ;
  assign n673 = ~n613 & ~n672 ;
  assign n686 = ~n248 & n402 ;
  assign n689 = n688 ^ n686 ;
  assign n692 = n691 ^ n689 ;
  assign n695 = n694 ^ n692 ;
  assign n676 = n248 & n380 ;
  assign n679 = n678 ^ n676 ;
  assign n682 = n681 ^ n679 ;
  assign n685 = n684 ^ n682 ;
  assign n696 = n695 ^ n685 ;
  assign n674 = x4 & ~n103 ;
  assign n675 = n674 ^ n368 ;
  assign n698 = n696 ^ n675 ;
  assign n711 = ~n248 & n447 ;
  assign n714 = n713 ^ n711 ;
  assign n717 = n716 ^ n714 ;
  assign n720 = n719 ^ n717 ;
  assign n701 = n248 & n425 ;
  assign n704 = n703 ^ n701 ;
  assign n707 = n706 ^ n704 ;
  assign n710 = n709 ^ n707 ;
  assign n721 = n720 ^ n710 ;
  assign n699 = x5 & ~n103 ;
  assign n700 = n699 ^ n413 ;
  assign n727 = n721 ^ n700 ;
  assign n728 = n698 & n727 ;
  assign n729 = n728 ^ n698 ;
  assign n730 = n729 ^ n727 ;
  assign n823 = ~n248 & n495 ;
  assign n826 = n825 ^ n823 ;
  assign n827 = n826 ^ n792 ;
  assign n829 = n828 ^ n827 ;
  assign n816 = n248 & n473 ;
  assign n819 = n818 ^ n816 ;
  assign n820 = n819 ^ n779 ;
  assign n822 = n821 ^ n820 ;
  assign n830 = n829 ^ n822 ;
  assign n731 = x6 & ~n103 ;
  assign n732 = n731 ^ n461 ;
  assign n831 = n830 ^ n732 ;
  assign n832 = n248 & n540 ;
  assign n835 = n834 ^ n832 ;
  assign n838 = n837 ^ n835 ;
  assign n841 = n840 ^ n838 ;
  assign n852 = n851 ^ n841 ;
  assign n747 = x15 & ~n93 ;
  assign n746 = x15 & ~n102 ;
  assign n748 = n747 ^ n746 ;
  assign n749 = n748 ^ n520 ;
  assign n743 = x7 & n93 ;
  assign n742 = x7 & ~n102 ;
  assign n744 = n743 ^ n742 ;
  assign n745 = n744 ^ n530 ;
  assign n750 = n749 ^ n745 ;
  assign n853 = n852 ^ n750 ;
  assign n854 = n831 & n853 ;
  assign n855 = n854 ^ n831 ;
  assign n856 = n855 ^ n853 ;
  assign n857 = ~n730 & ~n856 ;
  assign n858 = n673 & n857 ;
  assign n736 = n344 & ~n348 ;
  assign n737 = n736 ^ n248 ;
  assign n803 = ~n495 & n732 ;
  assign n807 = ~n737 & n803 ;
  assign n806 = ~n548 & n803 ;
  assign n808 = n807 ^ n806 ;
  assign n804 = ~n358 & n803 ;
  assign n805 = n567 & n804 ;
  assign n809 = n808 ^ n805 ;
  assign n762 = ~n540 & n750 ;
  assign n768 = ~n348 & n762 ;
  assign n769 = n344 & n768 ;
  assign n767 = n248 & n762 ;
  assign n770 = n769 ^ n767 ;
  assign n765 = n548 & n762 ;
  assign n766 = n765 ^ n762 ;
  assign n771 = n770 ^ n766 ;
  assign n763 = ~n358 & n762 ;
  assign n764 = n567 & n763 ;
  assign n772 = n771 ^ n764 ;
  assign n751 = ~n518 & n750 ;
  assign n757 = ~n348 & n751 ;
  assign n758 = n344 & n757 ;
  assign n756 = ~n248 & n751 ;
  assign n759 = n758 ^ n756 ;
  assign n754 = n548 & n751 ;
  assign n755 = n754 ^ n751 ;
  assign n760 = n759 ^ n755 ;
  assign n752 = ~n358 & n751 ;
  assign n753 = n567 & n752 ;
  assign n761 = n760 ^ n753 ;
  assign n773 = n772 ^ n761 ;
  assign n795 = ~n348 & ~n495 ;
  assign n796 = n344 & n795 ;
  assign n794 = ~n248 & ~n495 ;
  assign n797 = n796 ^ n794 ;
  assign n793 = n792 ^ n548 ;
  assign n798 = n797 ^ n793 ;
  assign n789 = n788 ^ n358 ;
  assign n790 = n567 & ~n789 ;
  assign n799 = n798 ^ n790 ;
  assign n800 = n773 & ~n799 ;
  assign n782 = ~n348 & ~n473 ;
  assign n783 = n344 & n782 ;
  assign n781 = n248 & ~n473 ;
  assign n784 = n783 ^ n781 ;
  assign n780 = n779 ^ n548 ;
  assign n785 = n784 ^ n780 ;
  assign n776 = n775 ^ n358 ;
  assign n777 = n567 & ~n776 ;
  assign n786 = n785 ^ n777 ;
  assign n787 = n773 & ~n786 ;
  assign n801 = n800 ^ n787 ;
  assign n774 = n732 & n773 ;
  assign n802 = n801 ^ n774 ;
  assign n810 = n809 ^ n802 ;
  assign n733 = ~n473 & n732 ;
  assign n739 = n548 & n733 ;
  assign n738 = n733 & ~n737 ;
  assign n740 = n739 ^ n738 ;
  assign n734 = ~n358 & n733 ;
  assign n735 = n567 & n734 ;
  assign n741 = n740 ^ n735 ;
  assign n811 = n810 ^ n741 ;
  assign n812 = ~n730 & n811 ;
  assign n722 = n700 & n721 ;
  assign n723 = n722 ^ n700 ;
  assign n724 = n698 & n723 ;
  assign n725 = n724 ^ n723 ;
  assign n697 = n675 & ~n696 ;
  assign n726 = n725 ^ n697 ;
  assign n813 = n812 ^ n726 ;
  assign n814 = n673 & n813 ;
  assign n662 = n640 & n661 ;
  assign n663 = n662 ^ n640 ;
  assign n664 = n638 & n663 ;
  assign n665 = n664 ^ n663 ;
  assign n637 = n615 & ~n636 ;
  assign n666 = n665 ^ n637 ;
  assign n667 = ~n613 & n666 ;
  assign n607 = ~n604 & n606 ;
  assign n608 = ~n583 & n607 ;
  assign n582 = n115 & ~n581 ;
  assign n609 = n608 ^ n582 ;
  assign n668 = n667 ^ n609 ;
  assign n815 = n814 ^ n668 ;
  assign n859 = n858 ^ n815 ;
  assign n1568 = n115 & n859 ;
  assign n861 = n581 & n859 ;
  assign n1567 = n861 ^ n581 ;
  assign n1569 = n1568 ^ n1567 ;
  assign n1592 = n1591 ^ n1569 ;
  assign n1617 = n606 & n859 ;
  assign n1615 = n604 & n859 ;
  assign n1616 = n1615 ^ n604 ;
  assign n1618 = n1617 ^ n1616 ;
  assign n1608 = n1353 & ~n1366 ;
  assign n1609 = n1453 & n1608 ;
  assign n1607 = n1353 & n1446 ;
  assign n1610 = n1609 ^ n1607 ;
  assign n1611 = n1610 ^ n1353 ;
  assign n1605 = n1353 & n1440 ;
  assign n1606 = n1605 ^ n1353 ;
  assign n1612 = n1611 ^ n1606 ;
  assign n1603 = n1353 & n1432 ;
  assign n1604 = n1301 & n1603 ;
  assign n1613 = n1612 ^ n1604 ;
  assign n1598 = n1362 & ~n1366 ;
  assign n1599 = n1453 & n1598 ;
  assign n1597 = n1362 & n1446 ;
  assign n1600 = n1599 ^ n1597 ;
  assign n1595 = n1362 & n1440 ;
  assign n1596 = n1595 ^ n1362 ;
  assign n1601 = n1600 ^ n1596 ;
  assign n1593 = n1362 & n1432 ;
  assign n1594 = n1301 & n1593 ;
  assign n1602 = n1601 ^ n1594 ;
  assign n1614 = n1613 ^ n1602 ;
  assign n1619 = n1618 ^ n1614 ;
  assign n1620 = n1592 & n1619 ;
  assign n1621 = n1620 ^ n1592 ;
  assign n1622 = n1621 ^ n1619 ;
  assign n1647 = n615 & n859 ;
  assign n1645 = n636 & n859 ;
  assign n1646 = n1645 ^ n636 ;
  assign n1648 = n1647 ^ n1646 ;
  assign n1638 = ~n1366 & n1387 ;
  assign n1639 = n1453 & n1638 ;
  assign n1637 = n1387 & n1446 ;
  assign n1640 = n1639 ^ n1637 ;
  assign n1641 = n1640 ^ n1387 ;
  assign n1635 = n1387 & n1440 ;
  assign n1636 = n1635 ^ n1387 ;
  assign n1642 = n1641 ^ n1636 ;
  assign n1633 = n1387 & n1432 ;
  assign n1634 = n1301 & n1633 ;
  assign n1643 = n1642 ^ n1634 ;
  assign n1628 = ~n1366 & n1396 ;
  assign n1629 = n1453 & n1628 ;
  assign n1627 = n1396 & n1446 ;
  assign n1630 = n1629 ^ n1627 ;
  assign n1625 = n1396 & n1440 ;
  assign n1626 = n1625 ^ n1396 ;
  assign n1631 = n1630 ^ n1626 ;
  assign n1623 = n1396 & n1432 ;
  assign n1624 = n1301 & n1623 ;
  assign n1632 = n1631 ^ n1624 ;
  assign n1644 = n1643 ^ n1632 ;
  assign n1649 = n1648 ^ n1644 ;
  assign n1652 = n640 & n859 ;
  assign n1650 = n661 & n859 ;
  assign n1651 = n1650 ^ n661 ;
  assign n1653 = n1652 ^ n1651 ;
  assign n1669 = ~n1366 & n1427 ;
  assign n1670 = n1453 & n1669 ;
  assign n1668 = n1427 & n1446 ;
  assign n1671 = n1670 ^ n1668 ;
  assign n1672 = n1671 ^ n1427 ;
  assign n1666 = n1427 & n1440 ;
  assign n1667 = n1666 ^ n1427 ;
  assign n1673 = n1672 ^ n1667 ;
  assign n1664 = n1427 & n1432 ;
  assign n1665 = n1301 & n1664 ;
  assign n1674 = n1673 ^ n1665 ;
  assign n1659 = ~n1366 & n1406 ;
  assign n1660 = n1453 & n1659 ;
  assign n1658 = n1406 & n1446 ;
  assign n1661 = n1660 ^ n1658 ;
  assign n1656 = n1406 & n1440 ;
  assign n1657 = n1656 ^ n1406 ;
  assign n1662 = n1661 ^ n1657 ;
  assign n1654 = n1406 & n1432 ;
  assign n1655 = n1301 & n1654 ;
  assign n1663 = n1662 ^ n1655 ;
  assign n1675 = n1674 ^ n1663 ;
  assign n1695 = n1653 & n1675 ;
  assign n1696 = n1695 ^ n1653 ;
  assign n1697 = n1649 & n1696 ;
  assign n1698 = n1697 ^ n1696 ;
  assign n1694 = ~n1644 & n1648 ;
  assign n1699 = n1698 ^ n1694 ;
  assign n1700 = ~n1622 & n1699 ;
  assign n1691 = ~n1614 & n1618 ;
  assign n1692 = ~n1592 & n1691 ;
  assign n1690 = n1569 & ~n1591 ;
  assign n1693 = n1692 ^ n1690 ;
  assign n1701 = n1700 ^ n1693 ;
  assign n1709 = n1591 & ~n1701 ;
  assign n1676 = n1675 ^ n1653 ;
  assign n1677 = n1649 & n1676 ;
  assign n1678 = n1677 ^ n1649 ;
  assign n1679 = n1678 ^ n1676 ;
  assign n1680 = ~n1622 & ~n1679 ;
  assign n1464 = n1195 & ~n1366 ;
  assign n1465 = n1453 & n1464 ;
  assign n1463 = n1195 & n1446 ;
  assign n1466 = n1465 ^ n1463 ;
  assign n1467 = n1466 ^ n1195 ;
  assign n1461 = n1195 & n1440 ;
  assign n1462 = n1461 ^ n1195 ;
  assign n1468 = n1467 ^ n1462 ;
  assign n1459 = n1195 & n1432 ;
  assign n1460 = n1301 & n1459 ;
  assign n1469 = n1468 ^ n1460 ;
  assign n1454 = n875 & ~n1366 ;
  assign n1455 = n1453 & n1454 ;
  assign n1447 = n875 & n1446 ;
  assign n1456 = n1455 ^ n1447 ;
  assign n1441 = n875 & n1440 ;
  assign n1442 = n1441 ^ n875 ;
  assign n1457 = n1456 ^ n1442 ;
  assign n1433 = n875 & n1432 ;
  assign n1434 = n1301 & n1433 ;
  assign n1458 = n1457 ^ n1434 ;
  assign n1470 = n1469 ^ n1458 ;
  assign n865 = n675 & n859 ;
  assign n863 = n696 & n859 ;
  assign n864 = n863 ^ n696 ;
  assign n866 = n865 ^ n864 ;
  assign n1472 = n1470 ^ n866 ;
  assign n1492 = n1227 & ~n1366 ;
  assign n1493 = n1453 & n1492 ;
  assign n1491 = n1227 & n1446 ;
  assign n1494 = n1493 ^ n1491 ;
  assign n1495 = n1494 ^ n1227 ;
  assign n1489 = n1227 & n1440 ;
  assign n1490 = n1489 ^ n1227 ;
  assign n1496 = n1495 ^ n1490 ;
  assign n1487 = n1227 & n1432 ;
  assign n1488 = n1301 & n1487 ;
  assign n1497 = n1496 ^ n1488 ;
  assign n1482 = n1206 & ~n1366 ;
  assign n1483 = n1453 & n1482 ;
  assign n1481 = n1206 & n1446 ;
  assign n1484 = n1483 ^ n1481 ;
  assign n1479 = n1206 & n1440 ;
  assign n1480 = n1479 ^ n1206 ;
  assign n1485 = n1484 ^ n1480 ;
  assign n1477 = n1206 & n1432 ;
  assign n1478 = n1301 & n1477 ;
  assign n1486 = n1485 ^ n1478 ;
  assign n1498 = n1497 ^ n1486 ;
  assign n1475 = n700 & n859 ;
  assign n1473 = n721 & n859 ;
  assign n1474 = n1473 ^ n721 ;
  assign n1476 = n1475 ^ n1474 ;
  assign n1502 = n1498 ^ n1476 ;
  assign n1503 = n1472 & n1502 ;
  assign n1504 = n1503 ^ n1472 ;
  assign n1505 = n1504 ^ n1502 ;
  assign n1525 = n1264 & ~n1366 ;
  assign n1526 = n1453 & n1525 ;
  assign n1524 = n1264 & n1446 ;
  assign n1527 = n1526 ^ n1524 ;
  assign n1528 = n1527 ^ n1264 ;
  assign n1522 = n1264 & n1440 ;
  assign n1523 = n1522 ^ n1264 ;
  assign n1529 = n1528 ^ n1523 ;
  assign n1520 = n1264 & n1432 ;
  assign n1521 = n1301 & n1520 ;
  assign n1530 = n1529 ^ n1521 ;
  assign n1515 = n1243 & ~n1366 ;
  assign n1516 = n1453 & n1515 ;
  assign n1514 = n1243 & n1446 ;
  assign n1517 = n1516 ^ n1514 ;
  assign n1512 = n1243 & n1440 ;
  assign n1513 = n1512 ^ n1243 ;
  assign n1518 = n1517 ^ n1513 ;
  assign n1510 = n1243 & n1432 ;
  assign n1511 = n1301 & n1510 ;
  assign n1519 = n1518 ^ n1511 ;
  assign n1531 = n1530 ^ n1519 ;
  assign n1508 = n732 & n859 ;
  assign n1506 = n830 & n859 ;
  assign n1507 = n1506 ^ n830 ;
  assign n1509 = n1508 ^ n1507 ;
  assign n1533 = n1531 ^ n1509 ;
  assign n1554 = n1294 & ~n1366 ;
  assign n1555 = n1453 & n1554 ;
  assign n1553 = n1294 & ~n1446 ;
  assign n1556 = n1555 ^ n1553 ;
  assign n1551 = n1294 & n1440 ;
  assign n1552 = n1551 ^ n1294 ;
  assign n1557 = n1556 ^ n1552 ;
  assign n1549 = n1294 & n1432 ;
  assign n1550 = n1301 & n1549 ;
  assign n1558 = n1557 ^ n1550 ;
  assign n1543 = n1272 & ~n1366 ;
  assign n1544 = n1453 & n1543 ;
  assign n1542 = n1272 & ~n1446 ;
  assign n1545 = n1544 ^ n1542 ;
  assign n1540 = n1272 & n1440 ;
  assign n1541 = n1540 ^ n1272 ;
  assign n1546 = n1545 ^ n1541 ;
  assign n1538 = n1272 & n1432 ;
  assign n1539 = n1301 & n1538 ;
  assign n1547 = n1546 ^ n1539 ;
  assign n1548 = n1547 ^ n1272 ;
  assign n1559 = n1558 ^ n1548 ;
  assign n1536 = n750 & n859 ;
  assign n1534 = n852 & n859 ;
  assign n1535 = n1534 ^ n852 ;
  assign n1537 = n1536 ^ n1535 ;
  assign n1683 = n1559 ^ n1537 ;
  assign n1684 = n1533 & n1683 ;
  assign n1685 = n1684 ^ n1533 ;
  assign n1686 = n1685 ^ n1683 ;
  assign n1687 = ~n1505 & ~n1686 ;
  assign n1688 = n1680 & n1687 ;
  assign n1708 = n1591 & ~n1688 ;
  assign n1710 = n1709 ^ n1708 ;
  assign n1560 = n1537 & n1559 ;
  assign n1561 = n1560 ^ n1537 ;
  assign n1562 = n1533 & n1561 ;
  assign n1563 = n1562 ^ n1561 ;
  assign n1532 = n1509 & ~n1531 ;
  assign n1564 = n1563 ^ n1532 ;
  assign n1565 = ~n1505 & n1564 ;
  assign n1499 = n1476 & ~n1498 ;
  assign n1500 = ~n1472 & n1499 ;
  assign n1471 = n866 & ~n1470 ;
  assign n1501 = n1500 ^ n1471 ;
  assign n1566 = n1565 ^ n1501 ;
  assign n1706 = n1591 & n1680 ;
  assign n1707 = n1566 & n1706 ;
  assign n1711 = n1710 ^ n1707 ;
  assign n1702 = n1569 & ~n1701 ;
  assign n1689 = n1569 & ~n1688 ;
  assign n1703 = n1702 ^ n1689 ;
  assign n1681 = n1569 & n1680 ;
  assign n1682 = n1566 & n1681 ;
  assign n1704 = n1703 ^ n1682 ;
  assign n1705 = n1704 ^ n1569 ;
  assign n1712 = n1711 ^ n1705 ;
  assign n860 = n115 & ~n859 ;
  assign n862 = n861 ^ n860 ;
  assign n1714 = n1712 ^ n862 ;
  assign n1727 = n1614 & ~n1701 ;
  assign n1726 = n1614 & ~n1688 ;
  assign n1728 = n1727 ^ n1726 ;
  assign n1724 = n1614 & n1680 ;
  assign n1725 = n1566 & n1724 ;
  assign n1729 = n1728 ^ n1725 ;
  assign n1720 = n1618 & ~n1701 ;
  assign n1719 = n1618 & ~n1688 ;
  assign n1721 = n1720 ^ n1719 ;
  assign n1717 = n1618 & n1680 ;
  assign n1718 = n1566 & n1717 ;
  assign n1722 = n1721 ^ n1718 ;
  assign n1723 = n1722 ^ n1618 ;
  assign n1730 = n1729 ^ n1723 ;
  assign n1715 = n606 & ~n859 ;
  assign n1716 = n1715 ^ n1615 ;
  assign n1734 = n1730 ^ n1716 ;
  assign n1735 = n1714 & n1734 ;
  assign n1736 = n1735 ^ n1714 ;
  assign n1737 = n1736 ^ n1734 ;
  assign n1750 = n1644 & ~n1701 ;
  assign n1749 = n1644 & ~n1688 ;
  assign n1751 = n1750 ^ n1749 ;
  assign n1747 = n1644 & n1680 ;
  assign n1748 = n1566 & n1747 ;
  assign n1752 = n1751 ^ n1748 ;
  assign n1743 = n1648 & ~n1701 ;
  assign n1742 = n1648 & ~n1688 ;
  assign n1744 = n1743 ^ n1742 ;
  assign n1740 = n1648 & n1680 ;
  assign n1741 = n1566 & n1740 ;
  assign n1745 = n1744 ^ n1741 ;
  assign n1746 = n1745 ^ n1648 ;
  assign n1753 = n1752 ^ n1746 ;
  assign n1738 = n615 & ~n859 ;
  assign n1739 = n1738 ^ n1645 ;
  assign n1755 = n1753 ^ n1739 ;
  assign n1768 = n1675 & ~n1701 ;
  assign n1767 = n1675 & ~n1688 ;
  assign n1769 = n1768 ^ n1767 ;
  assign n1765 = n1675 & n1680 ;
  assign n1766 = n1566 & n1765 ;
  assign n1770 = n1769 ^ n1766 ;
  assign n1761 = n1653 & ~n1701 ;
  assign n1760 = n1653 & ~n1688 ;
  assign n1762 = n1761 ^ n1760 ;
  assign n1758 = n1653 & n1680 ;
  assign n1759 = n1566 & n1758 ;
  assign n1763 = n1762 ^ n1759 ;
  assign n1764 = n1763 ^ n1653 ;
  assign n1771 = n1770 ^ n1764 ;
  assign n1756 = n640 & ~n859 ;
  assign n1757 = n1756 ^ n1650 ;
  assign n1779 = n1771 ^ n1757 ;
  assign n1780 = n1755 & n1779 ;
  assign n1781 = n1780 ^ n1755 ;
  assign n1782 = n1781 ^ n1779 ;
  assign n1783 = ~n1737 & ~n1782 ;
  assign n1796 = n1470 & ~n1701 ;
  assign n1795 = n1470 & ~n1688 ;
  assign n1797 = n1796 ^ n1795 ;
  assign n1793 = n1470 & n1680 ;
  assign n1794 = n1566 & n1793 ;
  assign n1798 = n1797 ^ n1794 ;
  assign n1789 = n866 & ~n1701 ;
  assign n1788 = n866 & ~n1688 ;
  assign n1790 = n1789 ^ n1788 ;
  assign n1786 = n866 & n1680 ;
  assign n1787 = n1566 & n1786 ;
  assign n1791 = n1790 ^ n1787 ;
  assign n1792 = n1791 ^ n866 ;
  assign n1799 = n1798 ^ n1792 ;
  assign n1784 = n675 & ~n859 ;
  assign n1785 = n1784 ^ n863 ;
  assign n1801 = n1799 ^ n1785 ;
  assign n1814 = n1498 & ~n1701 ;
  assign n1813 = n1498 & ~n1688 ;
  assign n1815 = n1814 ^ n1813 ;
  assign n1811 = n1498 & n1680 ;
  assign n1812 = n1566 & n1811 ;
  assign n1816 = n1815 ^ n1812 ;
  assign n1807 = n1476 & ~n1701 ;
  assign n1806 = n1476 & ~n1688 ;
  assign n1808 = n1807 ^ n1806 ;
  assign n1804 = n1476 & n1680 ;
  assign n1805 = n1566 & n1804 ;
  assign n1809 = n1808 ^ n1805 ;
  assign n1810 = n1809 ^ n1476 ;
  assign n1817 = n1816 ^ n1810 ;
  assign n1802 = n700 & ~n859 ;
  assign n1803 = n1802 ^ n1473 ;
  assign n1823 = n1817 ^ n1803 ;
  assign n1824 = n1801 & n1823 ;
  assign n1825 = n1824 ^ n1801 ;
  assign n1826 = n1825 ^ n1823 ;
  assign n1865 = n1531 & ~n1701 ;
  assign n1864 = n1531 & ~n1688 ;
  assign n1866 = n1865 ^ n1864 ;
  assign n1862 = n1531 & n1680 ;
  assign n1863 = n1566 & n1862 ;
  assign n1867 = n1866 ^ n1863 ;
  assign n1856 = n1509 & ~n1701 ;
  assign n1855 = n1509 & ~n1688 ;
  assign n1857 = n1856 ^ n1855 ;
  assign n1853 = n1509 & n1680 ;
  assign n1854 = n1566 & n1853 ;
  assign n1858 = n1857 ^ n1854 ;
  assign n1859 = n1858 ^ n1509 ;
  assign n1880 = n1867 ^ n1859 ;
  assign n1830 = n732 & ~n859 ;
  assign n1831 = n1830 ^ n1506 ;
  assign n1881 = n1880 ^ n1831 ;
  assign n1894 = n1559 & ~n1622 ;
  assign n1895 = n1699 & n1894 ;
  assign n1893 = n1559 & n1693 ;
  assign n1896 = n1895 ^ n1893 ;
  assign n1897 = n1896 ^ n1559 ;
  assign n1891 = n1559 & n1688 ;
  assign n1892 = n1891 ^ n1559 ;
  assign n1898 = n1897 ^ n1892 ;
  assign n1889 = n1559 & n1680 ;
  assign n1890 = n1566 & n1889 ;
  assign n1899 = n1898 ^ n1890 ;
  assign n1885 = n1537 & ~n1701 ;
  assign n1884 = n1537 & ~n1688 ;
  assign n1886 = n1885 ^ n1884 ;
  assign n1882 = n1537 & n1680 ;
  assign n1883 = n1566 & n1882 ;
  assign n1887 = n1886 ^ n1883 ;
  assign n1888 = n1887 ^ n1537 ;
  assign n1900 = n1899 ^ n1888 ;
  assign n1834 = n750 & ~n859 ;
  assign n1835 = n1834 ^ n1534 ;
  assign n1901 = n1900 ^ n1835 ;
  assign n1902 = n1881 & n1901 ;
  assign n1903 = n1902 ^ n1881 ;
  assign n1904 = n1903 ^ n1901 ;
  assign n1905 = ~n1826 & ~n1904 ;
  assign n1906 = n1783 & n1905 ;
  assign n1827 = n1566 & n1680 ;
  assign n1828 = n1827 ^ n1701 ;
  assign n1829 = n1828 ^ n1688 ;
  assign n1872 = ~n1531 & n1831 ;
  assign n1873 = n1829 & n1872 ;
  assign n1844 = ~n1559 & n1835 ;
  assign n1848 = ~n1701 & n1844 ;
  assign n1847 = ~n1688 & n1844 ;
  assign n1849 = n1848 ^ n1847 ;
  assign n1845 = n1680 & n1844 ;
  assign n1846 = n1566 & n1845 ;
  assign n1850 = n1849 ^ n1846 ;
  assign n1836 = ~n1537 & n1835 ;
  assign n1840 = ~n1701 & n1836 ;
  assign n1839 = ~n1688 & n1836 ;
  assign n1841 = n1840 ^ n1839 ;
  assign n1837 = n1680 & n1836 ;
  assign n1838 = n1566 & n1837 ;
  assign n1842 = n1841 ^ n1838 ;
  assign n1843 = n1842 ^ n1836 ;
  assign n1851 = n1850 ^ n1843 ;
  assign n1868 = n1867 ^ n1829 ;
  assign n1869 = n1851 & n1868 ;
  assign n1860 = n1859 ^ n1829 ;
  assign n1861 = n1851 & ~n1860 ;
  assign n1870 = n1869 ^ n1861 ;
  assign n1852 = n1831 & n1851 ;
  assign n1871 = n1870 ^ n1852 ;
  assign n1874 = n1873 ^ n1871 ;
  assign n1832 = ~n1509 & n1831 ;
  assign n1833 = ~n1829 & n1832 ;
  assign n1875 = n1874 ^ n1833 ;
  assign n1876 = ~n1826 & n1875 ;
  assign n1818 = n1803 & n1817 ;
  assign n1819 = n1818 ^ n1803 ;
  assign n1820 = n1801 & n1819 ;
  assign n1821 = n1820 ^ n1819 ;
  assign n1800 = n1785 & ~n1799 ;
  assign n1822 = n1821 ^ n1800 ;
  assign n1877 = n1876 ^ n1822 ;
  assign n1878 = n1783 & n1877 ;
  assign n1772 = n1757 & n1771 ;
  assign n1773 = n1772 ^ n1757 ;
  assign n1774 = n1755 & n1773 ;
  assign n1775 = n1774 ^ n1773 ;
  assign n1754 = n1739 & ~n1753 ;
  assign n1776 = n1775 ^ n1754 ;
  assign n1777 = ~n1737 & n1776 ;
  assign n1731 = n1716 & ~n1730 ;
  assign n1732 = ~n1714 & n1731 ;
  assign n1713 = n862 & ~n1712 ;
  assign n1733 = n1732 ^ n1713 ;
  assign n1778 = n1777 ^ n1733 ;
  assign n1879 = n1878 ^ n1778 ;
  assign n1907 = n1906 ^ n1879 ;
  assign n1910 = n1712 & n1907 ;
  assign n1908 = n862 & n1907 ;
  assign n1909 = n1908 ^ n862 ;
  assign n1911 = n1910 ^ n1909 ;
  assign n1914 = n1730 & n1907 ;
  assign n1912 = n1716 & n1907 ;
  assign n1913 = n1912 ^ n1716 ;
  assign n1915 = n1914 ^ n1913 ;
  assign n1918 = n1753 & n1907 ;
  assign n1916 = n1739 & n1907 ;
  assign n1917 = n1916 ^ n1739 ;
  assign n1919 = n1918 ^ n1917 ;
  assign n1922 = n1771 & n1907 ;
  assign n1920 = n1757 & n1907 ;
  assign n1921 = n1920 ^ n1757 ;
  assign n1923 = n1922 ^ n1921 ;
  assign n1926 = n1799 & n1907 ;
  assign n1924 = n1785 & n1907 ;
  assign n1925 = n1924 ^ n1785 ;
  assign n1927 = n1926 ^ n1925 ;
  assign n1930 = n1817 & n1907 ;
  assign n1928 = n1803 & n1907 ;
  assign n1929 = n1928 ^ n1803 ;
  assign n1931 = n1930 ^ n1929 ;
  assign n1934 = n1880 & n1907 ;
  assign n1932 = n1831 & n1907 ;
  assign n1933 = n1932 ^ n1831 ;
  assign n1935 = n1934 ^ n1933 ;
  assign n1938 = n1900 & n1907 ;
  assign n1936 = n1835 & n1907 ;
  assign n1937 = n1936 ^ n1835 ;
  assign n1939 = n1938 ^ n1937 ;
  assign n1940 = n1910 ^ n1712 ;
  assign n1941 = n1940 ^ n1908 ;
  assign n1942 = n1914 ^ n1730 ;
  assign n1943 = n1942 ^ n1912 ;
  assign n1944 = n1918 ^ n1753 ;
  assign n1945 = n1944 ^ n1916 ;
  assign n1946 = n1922 ^ n1771 ;
  assign n1947 = n1946 ^ n1920 ;
  assign n1948 = n1926 ^ n1799 ;
  assign n1949 = n1948 ^ n1924 ;
  assign n1950 = n1930 ^ n1817 ;
  assign n1951 = n1950 ^ n1928 ;
  assign n1952 = n1934 ^ n1880 ;
  assign n1953 = n1952 ^ n1932 ;
  assign n1954 = n1938 ^ n1900 ;
  assign n1955 = n1954 ^ n1936 ;
  assign n1975 = n896 & ~n909 ;
  assign n1973 = ~n901 & n932 ;
  assign n1974 = n1973 ^ n925 ;
  assign n1976 = n1975 ^ n1974 ;
  assign n1977 = n1976 ^ n919 ;
  assign n1978 = x40 & ~n1977 ;
  assign n1979 = n1978 ^ n1059 ;
  assign n1984 = n1049 & ~n1172 ;
  assign n1985 = n1984 ^ n1317 ;
  assign n1986 = n1985 ^ n1314 ;
  assign n1987 = n1986 ^ n1312 ;
  assign n1980 = n1071 & n1172 ;
  assign n1981 = n1980 ^ n1327 ;
  assign n1982 = n1981 ^ n1324 ;
  assign n1983 = n1982 ^ n1322 ;
  assign n1988 = n1987 ^ n1983 ;
  assign n1990 = n1988 ^ n1979 ;
  assign n2000 = x41 & ~n1977 ;
  assign n2001 = n2000 ^ n1084 ;
  assign n1995 = n1074 & ~n1172 ;
  assign n1996 = n1995 ^ n1339 ;
  assign n1997 = n1996 ^ n1336 ;
  assign n1998 = n1997 ^ n1334 ;
  assign n1991 = n1096 & n1172 ;
  assign n1992 = n1991 ^ n1349 ;
  assign n1993 = n1992 ^ n1346 ;
  assign n1994 = n1993 ^ n1344 ;
  assign n1999 = n1998 ^ n1994 ;
  assign n2005 = n2001 ^ n1999 ;
  assign n2006 = n1990 & n2005 ;
  assign n2007 = n2006 ^ n1990 ;
  assign n2008 = n2007 ^ n2005 ;
  assign n2018 = x42 & ~n1977 ;
  assign n2019 = n2018 ^ n1112 ;
  assign n2013 = n1102 & ~n1172 ;
  assign n2014 = n2013 ^ n1373 ;
  assign n2015 = n2014 ^ n1370 ;
  assign n2016 = n2015 ^ n1368 ;
  assign n2009 = n1124 & n1172 ;
  assign n2010 = n2009 ^ n1383 ;
  assign n2011 = n2010 ^ n1380 ;
  assign n2012 = n2011 ^ n1378 ;
  assign n2017 = n2016 ^ n2012 ;
  assign n2021 = n2019 ^ n2017 ;
  assign n2031 = x43 & ~n1977 ;
  assign n2032 = n2031 ^ n1137 ;
  assign n2026 = n1127 & ~n1172 ;
  assign n2027 = n2026 ^ n1413 ;
  assign n2028 = n2027 ^ n1410 ;
  assign n2029 = n2028 ^ n1408 ;
  assign n2022 = n1149 & n1172 ;
  assign n2023 = n2022 ^ n1423 ;
  assign n2024 = n2023 ^ n1420 ;
  assign n2025 = n2024 ^ n1418 ;
  assign n2030 = n2029 ^ n2025 ;
  assign n2040 = n2032 ^ n2030 ;
  assign n2041 = n2021 & n2040 ;
  assign n2042 = n2041 ^ n2021 ;
  assign n2043 = n2042 ^ n2040 ;
  assign n2044 = ~n2008 & ~n2043 ;
  assign n2045 = x44 & ~n1977 ;
  assign n2046 = n2045 ^ n937 ;
  assign n1968 = n877 & ~n1172 ;
  assign n1969 = n1968 ^ n1181 ;
  assign n1970 = n1969 ^ n1168 ;
  assign n1971 = n1970 ^ n1158 ;
  assign n1964 = n949 & n1172 ;
  assign n1965 = n1964 ^ n1191 ;
  assign n1966 = n1965 ^ n1188 ;
  assign n1967 = n1966 ^ n1186 ;
  assign n1972 = n1971 ^ n1967 ;
  assign n2048 = n2046 ^ n1972 ;
  assign n2058 = x45 & ~n1977 ;
  assign n2059 = n2058 ^ n963 ;
  assign n2053 = n953 & ~n1172 ;
  assign n2054 = n2053 ^ n1213 ;
  assign n2055 = n2054 ^ n1210 ;
  assign n2056 = n2055 ^ n1208 ;
  assign n2049 = n975 & n1172 ;
  assign n2050 = n2049 ^ n1223 ;
  assign n2051 = n2050 ^ n1220 ;
  assign n2052 = n2051 ^ n1218 ;
  assign n2057 = n2056 ^ n2052 ;
  assign n2065 = n2059 ^ n2057 ;
  assign n2066 = n2048 & n2065 ;
  assign n2067 = n2066 ^ n2048 ;
  assign n2068 = n2067 ^ n2065 ;
  assign n2078 = x46 & ~n1977 ;
  assign n2079 = n2078 ^ n996 ;
  assign n2073 = n986 & ~n1172 ;
  assign n2074 = n2073 ^ n1250 ;
  assign n2075 = n2074 ^ n1247 ;
  assign n2076 = n2075 ^ n1245 ;
  assign n2069 = n1008 & n1172 ;
  assign n2070 = n2069 ^ n1260 ;
  assign n2071 = n2070 ^ n1257 ;
  assign n2072 = n2071 ^ n1255 ;
  assign n2077 = n2076 ^ n2072 ;
  assign n2125 = n2079 ^ n2077 ;
  assign n2126 = n1039 & n1172 ;
  assign n2127 = n2126 ^ n1290 ;
  assign n2128 = n2127 ^ n1287 ;
  assign n2129 = n2128 ^ n1285 ;
  assign n2130 = n2129 ^ n1282 ;
  assign n2087 = x39 & ~n1974 ;
  assign n2086 = x39 & ~n919 ;
  assign n2088 = n2087 ^ n2086 ;
  assign n2089 = n2088 ^ n1019 ;
  assign n2083 = x47 & n1974 ;
  assign n2082 = x47 & ~n919 ;
  assign n2084 = n2083 ^ n2082 ;
  assign n2085 = n2084 ^ n1029 ;
  assign n2090 = n2089 ^ n2085 ;
  assign n2131 = n2130 ^ n2090 ;
  assign n2132 = n2125 & n2131 ;
  assign n2133 = n2132 ^ n2125 ;
  assign n2134 = n2133 ^ n2131 ;
  assign n2135 = ~n2068 & ~n2134 ;
  assign n2136 = n2044 & n2135 ;
  assign n2102 = n1039 & ~n2090 ;
  assign n2108 = ~n1100 & n2102 ;
  assign n2109 = n1179 & n2108 ;
  assign n2107 = n1172 & n2102 ;
  assign n2110 = n2109 ^ n2107 ;
  assign n2105 = n1166 & n2102 ;
  assign n2106 = n2105 ^ n2102 ;
  assign n2111 = n2110 ^ n2106 ;
  assign n2103 = ~n1156 & n2102 ;
  assign n2104 = n1047 & n2103 ;
  assign n2112 = n2111 ^ n2104 ;
  assign n2091 = n1017 & ~n2090 ;
  assign n2097 = ~n1100 & n2091 ;
  assign n2098 = n1179 & n2097 ;
  assign n2096 = ~n1172 & n2091 ;
  assign n2099 = n2098 ^ n2096 ;
  assign n2094 = n1166 & n2091 ;
  assign n2095 = n2094 ^ n2091 ;
  assign n2100 = n2099 ^ n2095 ;
  assign n2092 = ~n1156 & n2091 ;
  assign n2093 = n1047 & n2092 ;
  assign n2101 = n2100 ^ n2093 ;
  assign n2113 = n2112 ^ n2101 ;
  assign n2117 = n2076 & n2113 ;
  assign n2116 = n2072 & n2113 ;
  assign n2118 = n2117 ^ n2116 ;
  assign n2114 = n2079 & n2113 ;
  assign n2115 = n2114 ^ n2113 ;
  assign n2119 = n2118 ^ n2115 ;
  assign n2080 = n2077 & n2079 ;
  assign n2081 = n2080 ^ n2077 ;
  assign n2120 = n2119 ^ n2081 ;
  assign n2121 = ~n2068 & n2120 ;
  assign n2060 = n2057 & n2059 ;
  assign n2061 = n2060 ^ n2057 ;
  assign n2062 = n2048 & n2061 ;
  assign n2063 = n2062 ^ n2061 ;
  assign n2047 = n1972 & ~n2046 ;
  assign n2064 = n2063 ^ n2047 ;
  assign n2122 = n2121 ^ n2064 ;
  assign n2123 = n2044 & n2122 ;
  assign n2033 = n2030 & n2032 ;
  assign n2034 = n2033 ^ n2030 ;
  assign n2035 = n2021 & n2034 ;
  assign n2036 = n2035 ^ n2034 ;
  assign n2020 = n2017 & ~n2019 ;
  assign n2037 = n2036 ^ n2020 ;
  assign n2038 = ~n2008 & n2037 ;
  assign n2002 = n1999 & ~n2001 ;
  assign n2003 = ~n1990 & n2002 ;
  assign n1989 = ~n1979 & n1988 ;
  assign n2004 = n2003 ^ n1989 ;
  assign n2039 = n2038 ^ n2004 ;
  assign n2124 = n2123 ^ n2039 ;
  assign n2137 = n2136 ^ n2124 ;
  assign n2194 = n1979 & n2137 ;
  assign n2192 = n1988 & n2137 ;
  assign n2193 = n2192 ^ n1988 ;
  assign n2195 = n2194 ^ n2193 ;
  assign n2188 = n1577 ^ n1310 ;
  assign n2189 = n2188 ^ n1573 ;
  assign n2190 = n2189 ^ n1571 ;
  assign n2186 = n1587 ^ n1583 ;
  assign n2187 = n2186 ^ n1581 ;
  assign n2191 = n2190 ^ n2187 ;
  assign n2196 = n2195 ^ n2191 ;
  assign n2203 = n1600 ^ n1362 ;
  assign n2204 = n2203 ^ n1596 ;
  assign n2205 = n2204 ^ n1594 ;
  assign n2201 = n1610 ^ n1606 ;
  assign n2202 = n2201 ^ n1604 ;
  assign n2206 = n2205 ^ n2202 ;
  assign n2199 = n2001 & n2137 ;
  assign n2197 = n1999 & n2137 ;
  assign n2198 = n2197 ^ n1999 ;
  assign n2200 = n2199 ^ n2198 ;
  assign n2207 = n2206 ^ n2200 ;
  assign n2208 = n2196 & n2207 ;
  assign n2209 = n2208 ^ n2196 ;
  assign n2210 = n2209 ^ n2207 ;
  assign n2217 = n1630 ^ n1396 ;
  assign n2218 = n2217 ^ n1626 ;
  assign n2219 = n2218 ^ n1624 ;
  assign n2215 = n1640 ^ n1636 ;
  assign n2216 = n2215 ^ n1634 ;
  assign n2220 = n2219 ^ n2216 ;
  assign n2213 = n2019 & n2137 ;
  assign n2211 = n2017 & n2137 ;
  assign n2212 = n2211 ^ n2017 ;
  assign n2214 = n2213 ^ n2212 ;
  assign n2221 = n2220 ^ n2214 ;
  assign n2224 = n1661 ^ n1406 ;
  assign n2225 = n2224 ^ n1657 ;
  assign n2226 = n2225 ^ n1655 ;
  assign n2222 = n1671 ^ n1667 ;
  assign n2223 = n2222 ^ n1665 ;
  assign n2227 = n2226 ^ n2223 ;
  assign n2230 = n2032 & n2137 ;
  assign n2228 = n2030 & n2137 ;
  assign n2229 = n2228 ^ n2030 ;
  assign n2231 = n2230 ^ n2229 ;
  assign n2251 = n2227 & n2231 ;
  assign n2252 = n2251 ^ n2227 ;
  assign n2253 = n2221 & n2252 ;
  assign n2254 = n2253 ^ n2252 ;
  assign n2250 = ~n2214 & n2220 ;
  assign n2255 = n2254 ^ n2250 ;
  assign n2256 = ~n2210 & n2255 ;
  assign n2247 = ~n2200 & n2206 ;
  assign n2248 = ~n2196 & n2247 ;
  assign n2246 = n2191 & ~n2195 ;
  assign n2249 = n2248 ^ n2246 ;
  assign n2257 = n2256 ^ n2249 ;
  assign n2369 = n2195 & ~n2257 ;
  assign n2232 = n2231 ^ n2227 ;
  assign n2233 = n2221 & n2232 ;
  assign n2234 = n2233 ^ n2221 ;
  assign n2235 = n2234 ^ n2232 ;
  assign n2236 = ~n2210 & ~n2235 ;
  assign n2140 = n2046 & n2137 ;
  assign n2138 = n1972 & n2137 ;
  assign n2139 = n2138 ^ n1972 ;
  assign n2141 = n2140 ^ n2139 ;
  assign n1960 = n1456 ^ n875 ;
  assign n1961 = n1960 ^ n1442 ;
  assign n1962 = n1961 ^ n1434 ;
  assign n1958 = n1466 ^ n1462 ;
  assign n1959 = n1958 ^ n1460 ;
  assign n1963 = n1962 ^ n1959 ;
  assign n2143 = n2141 ^ n1963 ;
  assign n2152 = n2059 & n2137 ;
  assign n2150 = n2057 & n2137 ;
  assign n2151 = n2150 ^ n2057 ;
  assign n2153 = n2152 ^ n2151 ;
  assign n2146 = n1484 ^ n1206 ;
  assign n2147 = n2146 ^ n1480 ;
  assign n2148 = n2147 ^ n1478 ;
  assign n2144 = n1494 ^ n1490 ;
  assign n2145 = n2144 ^ n1488 ;
  assign n2149 = n2148 ^ n2145 ;
  assign n2157 = n2153 ^ n2149 ;
  assign n2158 = n2143 & n2157 ;
  assign n2159 = n2158 ^ n2143 ;
  assign n2160 = n2159 ^ n2157 ;
  assign n2169 = n2079 & n2137 ;
  assign n2167 = n2077 & n2137 ;
  assign n2168 = n2167 ^ n2077 ;
  assign n2170 = n2169 ^ n2168 ;
  assign n2163 = n1517 ^ n1243 ;
  assign n2164 = n2163 ^ n1513 ;
  assign n2165 = n2164 ^ n1511 ;
  assign n2161 = n1527 ^ n1523 ;
  assign n2162 = n2161 ^ n1521 ;
  assign n2166 = n2165 ^ n2162 ;
  assign n2172 = n2170 ^ n2166 ;
  assign n2177 = n2090 & n2137 ;
  assign n2175 = n2130 & n2137 ;
  assign n2176 = n2175 ^ n2130 ;
  assign n2178 = n2177 ^ n2176 ;
  assign n2173 = n1558 ^ n1294 ;
  assign n2174 = n2173 ^ n1547 ;
  assign n2239 = n2178 ^ n2174 ;
  assign n2240 = n2172 & n2239 ;
  assign n2241 = n2240 ^ n2172 ;
  assign n2242 = n2241 ^ n2239 ;
  assign n2243 = ~n2160 & ~n2242 ;
  assign n2244 = n2236 & n2243 ;
  assign n2368 = n2195 & ~n2244 ;
  assign n2370 = n2369 ^ n2368 ;
  assign n2179 = n2174 & n2178 ;
  assign n2180 = n2179 ^ n2174 ;
  assign n2181 = n2172 & n2180 ;
  assign n2182 = n2181 ^ n2180 ;
  assign n2171 = n2166 & ~n2170 ;
  assign n2183 = n2182 ^ n2171 ;
  assign n2184 = ~n2160 & n2183 ;
  assign n2154 = n2149 & ~n2153 ;
  assign n2155 = ~n2143 & n2154 ;
  assign n2142 = n1963 & ~n2141 ;
  assign n2156 = n2155 ^ n2142 ;
  assign n2185 = n2184 ^ n2156 ;
  assign n2366 = n2195 & n2236 ;
  assign n2367 = n2185 & n2366 ;
  assign n2371 = n2370 ^ n2367 ;
  assign n2362 = n2191 & ~n2257 ;
  assign n2361 = n2191 & ~n2244 ;
  assign n2363 = n2362 ^ n2361 ;
  assign n2359 = n2191 & n2236 ;
  assign n2360 = n2185 & n2359 ;
  assign n2364 = n2363 ^ n2360 ;
  assign n2365 = n2364 ^ n2191 ;
  assign n2372 = n2371 ^ n2365 ;
  assign n2357 = n1711 ^ n1591 ;
  assign n2358 = n2357 ^ n1704 ;
  assign n2373 = n2372 ^ n2358 ;
  assign n2388 = n1729 ^ n1614 ;
  assign n2389 = n2388 ^ n1722 ;
  assign n2384 = n2200 & ~n2257 ;
  assign n2383 = n2200 & ~n2244 ;
  assign n2385 = n2384 ^ n2383 ;
  assign n2381 = n2200 & n2236 ;
  assign n2382 = n2185 & n2381 ;
  assign n2386 = n2385 ^ n2382 ;
  assign n2377 = n2206 & ~n2257 ;
  assign n2376 = n2206 & ~n2244 ;
  assign n2378 = n2377 ^ n2376 ;
  assign n2374 = n2206 & n2236 ;
  assign n2375 = n2185 & n2374 ;
  assign n2379 = n2378 ^ n2375 ;
  assign n2380 = n2379 ^ n2206 ;
  assign n2387 = n2386 ^ n2380 ;
  assign n2390 = n2389 ^ n2387 ;
  assign n2391 = n2373 & n2390 ;
  assign n2392 = n2391 ^ n2373 ;
  assign n2393 = n2392 ^ n2390 ;
  assign n2408 = n1752 ^ n1644 ;
  assign n2409 = n2408 ^ n1745 ;
  assign n2404 = n2214 & ~n2257 ;
  assign n2403 = n2214 & ~n2244 ;
  assign n2405 = n2404 ^ n2403 ;
  assign n2401 = n2214 & n2236 ;
  assign n2402 = n2185 & n2401 ;
  assign n2406 = n2405 ^ n2402 ;
  assign n2397 = n2220 & ~n2257 ;
  assign n2396 = n2220 & ~n2244 ;
  assign n2398 = n2397 ^ n2396 ;
  assign n2394 = n2220 & n2236 ;
  assign n2395 = n2185 & n2394 ;
  assign n2399 = n2398 ^ n2395 ;
  assign n2400 = n2399 ^ n2220 ;
  assign n2407 = n2406 ^ n2400 ;
  assign n2410 = n2409 ^ n2407 ;
  assign n2411 = n1770 ^ n1675 ;
  assign n2412 = n2411 ^ n1763 ;
  assign n2423 = n2231 & ~n2257 ;
  assign n2422 = n2231 & ~n2244 ;
  assign n2424 = n2423 ^ n2422 ;
  assign n2420 = n2231 & n2236 ;
  assign n2421 = n2185 & n2420 ;
  assign n2425 = n2424 ^ n2421 ;
  assign n2416 = n2227 & ~n2257 ;
  assign n2415 = n2227 & ~n2244 ;
  assign n2417 = n2416 ^ n2415 ;
  assign n2413 = n2227 & n2236 ;
  assign n2414 = n2185 & n2413 ;
  assign n2418 = n2417 ^ n2414 ;
  assign n2419 = n2418 ^ n2227 ;
  assign n2426 = n2425 ^ n2419 ;
  assign n2446 = n2412 & n2426 ;
  assign n2447 = n2446 ^ n2412 ;
  assign n2448 = n2410 & n2447 ;
  assign n2449 = n2448 ^ n2447 ;
  assign n2445 = ~n2407 & n2409 ;
  assign n2450 = n2449 ^ n2445 ;
  assign n2451 = ~n2393 & n2450 ;
  assign n2442 = ~n2387 & n2389 ;
  assign n2443 = ~n2373 & n2442 ;
  assign n2441 = n2358 & ~n2372 ;
  assign n2444 = n2443 ^ n2441 ;
  assign n2452 = n2451 ^ n2444 ;
  assign n2460 = n2372 & ~n2452 ;
  assign n2427 = n2426 ^ n2412 ;
  assign n2428 = n2410 & n2427 ;
  assign n2429 = n2428 ^ n2410 ;
  assign n2430 = n2429 ^ n2427 ;
  assign n2431 = ~n2393 & ~n2430 ;
  assign n2265 = n2141 & ~n2257 ;
  assign n2264 = n2141 & ~n2244 ;
  assign n2266 = n2265 ^ n2264 ;
  assign n2262 = n2141 & n2236 ;
  assign n2263 = n2185 & n2262 ;
  assign n2267 = n2266 ^ n2263 ;
  assign n2258 = n1963 & ~n2257 ;
  assign n2245 = n1963 & ~n2244 ;
  assign n2259 = n2258 ^ n2245 ;
  assign n2237 = n1963 & n2236 ;
  assign n2238 = n2185 & n2237 ;
  assign n2260 = n2259 ^ n2238 ;
  assign n2261 = n2260 ^ n1963 ;
  assign n2268 = n2267 ^ n2261 ;
  assign n1956 = n1798 ^ n1470 ;
  assign n1957 = n1956 ^ n1791 ;
  assign n2270 = n2268 ^ n1957 ;
  assign n2283 = n2153 & ~n2257 ;
  assign n2282 = n2153 & ~n2244 ;
  assign n2284 = n2283 ^ n2282 ;
  assign n2280 = n2153 & n2236 ;
  assign n2281 = n2185 & n2280 ;
  assign n2285 = n2284 ^ n2281 ;
  assign n2276 = n2149 & ~n2257 ;
  assign n2275 = n2149 & ~n2244 ;
  assign n2277 = n2276 ^ n2275 ;
  assign n2273 = n2149 & n2236 ;
  assign n2274 = n2185 & n2273 ;
  assign n2278 = n2277 ^ n2274 ;
  assign n2279 = n2278 ^ n2149 ;
  assign n2286 = n2285 ^ n2279 ;
  assign n2271 = n1816 ^ n1498 ;
  assign n2272 = n2271 ^ n1809 ;
  assign n2292 = n2286 ^ n2272 ;
  assign n2293 = n2270 & n2292 ;
  assign n2294 = n2293 ^ n2270 ;
  assign n2295 = n2294 ^ n2292 ;
  assign n2308 = n2170 & ~n2257 ;
  assign n2307 = n2170 & ~n2244 ;
  assign n2309 = n2308 ^ n2307 ;
  assign n2305 = n2170 & n2236 ;
  assign n2306 = n2185 & n2305 ;
  assign n2310 = n2309 ^ n2306 ;
  assign n2301 = n2166 & ~n2257 ;
  assign n2300 = n2166 & ~n2244 ;
  assign n2302 = n2301 ^ n2300 ;
  assign n2298 = n2166 & n2236 ;
  assign n2299 = n2185 & n2298 ;
  assign n2303 = n2302 ^ n2299 ;
  assign n2304 = n2303 ^ n2166 ;
  assign n2311 = n2310 ^ n2304 ;
  assign n2296 = n1867 ^ n1531 ;
  assign n2297 = n2296 ^ n1858 ;
  assign n2314 = n2311 ^ n2297 ;
  assign n2343 = n2178 & ~n2210 ;
  assign n2344 = n2255 & n2343 ;
  assign n2342 = n2178 & n2249 ;
  assign n2345 = n2344 ^ n2342 ;
  assign n2346 = n2345 ^ n2178 ;
  assign n2340 = n2178 & n2244 ;
  assign n2341 = n2340 ^ n2178 ;
  assign n2347 = n2346 ^ n2341 ;
  assign n2338 = n2178 & n2236 ;
  assign n2339 = n2185 & n2338 ;
  assign n2348 = n2347 ^ n2339 ;
  assign n2331 = n2174 & ~n2210 ;
  assign n2332 = n2255 & n2331 ;
  assign n2330 = n2174 & n2249 ;
  assign n2333 = n2332 ^ n2330 ;
  assign n2334 = n2333 ^ n2174 ;
  assign n2328 = n2174 & n2244 ;
  assign n2329 = n2328 ^ n2174 ;
  assign n2335 = n2334 ^ n2329 ;
  assign n2326 = n2174 & n2236 ;
  assign n2327 = n2185 & n2326 ;
  assign n2336 = n2335 ^ n2327 ;
  assign n2337 = n2336 ^ n2174 ;
  assign n2349 = n2348 ^ n2337 ;
  assign n2319 = n1537 & ~n1622 ;
  assign n2320 = n1699 & n2319 ;
  assign n2318 = n1537 & n1693 ;
  assign n2321 = n2320 ^ n2318 ;
  assign n2322 = n2321 ^ n1537 ;
  assign n2316 = n1537 & n1688 ;
  assign n2317 = n2316 ^ n1537 ;
  assign n2323 = n2322 ^ n2317 ;
  assign n2324 = n2323 ^ n1883 ;
  assign n2315 = n1899 ^ n1559 ;
  assign n2325 = n2324 ^ n2315 ;
  assign n2434 = n2349 ^ n2325 ;
  assign n2435 = n2314 & n2434 ;
  assign n2436 = n2435 ^ n2314 ;
  assign n2437 = n2436 ^ n2434 ;
  assign n2438 = ~n2295 & ~n2437 ;
  assign n2439 = n2431 & n2438 ;
  assign n2459 = n2372 & ~n2439 ;
  assign n2461 = n2460 ^ n2459 ;
  assign n2350 = n2325 & n2349 ;
  assign n2351 = n2350 ^ n2325 ;
  assign n2352 = n2314 & n2351 ;
  assign n2353 = n2352 ^ n2351 ;
  assign n2312 = n2297 & n2311 ;
  assign n2313 = n2312 ^ n2297 ;
  assign n2354 = n2353 ^ n2313 ;
  assign n2355 = ~n2295 & n2354 ;
  assign n2287 = n2272 & n2286 ;
  assign n2288 = n2287 ^ n2272 ;
  assign n2289 = n2270 & n2288 ;
  assign n2290 = n2289 ^ n2288 ;
  assign n2269 = n1957 & ~n2268 ;
  assign n2291 = n2290 ^ n2269 ;
  assign n2356 = n2355 ^ n2291 ;
  assign n2457 = n2372 & n2431 ;
  assign n2458 = n2356 & n2457 ;
  assign n2462 = n2461 ^ n2458 ;
  assign n2453 = n2358 & ~n2452 ;
  assign n2440 = n2358 & ~n2439 ;
  assign n2454 = n2453 ^ n2440 ;
  assign n2432 = n2358 & n2431 ;
  assign n2433 = n2356 & n2432 ;
  assign n2455 = n2454 ^ n2433 ;
  assign n2456 = n2455 ^ n2358 ;
  assign n2463 = n2462 ^ n2456 ;
  assign n2474 = n2387 & ~n2452 ;
  assign n2473 = n2387 & ~n2439 ;
  assign n2475 = n2474 ^ n2473 ;
  assign n2471 = n2387 & n2431 ;
  assign n2472 = n2356 & n2471 ;
  assign n2476 = n2475 ^ n2472 ;
  assign n2467 = n2389 & ~n2452 ;
  assign n2466 = n2389 & ~n2439 ;
  assign n2468 = n2467 ^ n2466 ;
  assign n2464 = n2389 & n2431 ;
  assign n2465 = n2356 & n2464 ;
  assign n2469 = n2468 ^ n2465 ;
  assign n2470 = n2469 ^ n2389 ;
  assign n2477 = n2476 ^ n2470 ;
  assign n2488 = n2407 & ~n2452 ;
  assign n2487 = n2407 & ~n2439 ;
  assign n2489 = n2488 ^ n2487 ;
  assign n2485 = n2407 & n2431 ;
  assign n2486 = n2356 & n2485 ;
  assign n2490 = n2489 ^ n2486 ;
  assign n2481 = n2409 & ~n2452 ;
  assign n2480 = n2409 & ~n2439 ;
  assign n2482 = n2481 ^ n2480 ;
  assign n2478 = n2409 & n2431 ;
  assign n2479 = n2356 & n2478 ;
  assign n2483 = n2482 ^ n2479 ;
  assign n2484 = n2483 ^ n2409 ;
  assign n2491 = n2490 ^ n2484 ;
  assign n2502 = n2426 & ~n2452 ;
  assign n2501 = n2426 & ~n2439 ;
  assign n2503 = n2502 ^ n2501 ;
  assign n2499 = n2426 & n2431 ;
  assign n2500 = n2356 & n2499 ;
  assign n2504 = n2503 ^ n2500 ;
  assign n2495 = n2412 & ~n2452 ;
  assign n2494 = n2412 & ~n2439 ;
  assign n2496 = n2495 ^ n2494 ;
  assign n2492 = n2412 & n2431 ;
  assign n2493 = n2356 & n2492 ;
  assign n2497 = n2496 ^ n2493 ;
  assign n2498 = n2497 ^ n2412 ;
  assign n2505 = n2504 ^ n2498 ;
  assign n2516 = n2268 & ~n2452 ;
  assign n2515 = n2268 & ~n2439 ;
  assign n2517 = n2516 ^ n2515 ;
  assign n2513 = n2268 & n2431 ;
  assign n2514 = n2356 & n2513 ;
  assign n2518 = n2517 ^ n2514 ;
  assign n2509 = n1957 & ~n2452 ;
  assign n2508 = n1957 & ~n2439 ;
  assign n2510 = n2509 ^ n2508 ;
  assign n2506 = n1957 & n2431 ;
  assign n2507 = n2356 & n2506 ;
  assign n2511 = n2510 ^ n2507 ;
  assign n2512 = n2511 ^ n1957 ;
  assign n2519 = n2518 ^ n2512 ;
  assign n2530 = n2286 & ~n2452 ;
  assign n2529 = n2286 & ~n2439 ;
  assign n2531 = n2530 ^ n2529 ;
  assign n2527 = n2286 & n2431 ;
  assign n2528 = n2356 & n2527 ;
  assign n2532 = n2531 ^ n2528 ;
  assign n2523 = n2272 & ~n2452 ;
  assign n2522 = n2272 & ~n2439 ;
  assign n2524 = n2523 ^ n2522 ;
  assign n2520 = n2272 & n2431 ;
  assign n2521 = n2356 & n2520 ;
  assign n2525 = n2524 ^ n2521 ;
  assign n2526 = n2525 ^ n2272 ;
  assign n2533 = n2532 ^ n2526 ;
  assign n2544 = n2311 & ~n2452 ;
  assign n2543 = n2311 & ~n2439 ;
  assign n2545 = n2544 ^ n2543 ;
  assign n2541 = n2311 & n2431 ;
  assign n2542 = n2356 & n2541 ;
  assign n2546 = n2545 ^ n2542 ;
  assign n2537 = n2297 & ~n2452 ;
  assign n2536 = n2297 & ~n2439 ;
  assign n2538 = n2537 ^ n2536 ;
  assign n2534 = n2297 & n2431 ;
  assign n2535 = n2356 & n2534 ;
  assign n2539 = n2538 ^ n2535 ;
  assign n2540 = n2539 ^ n2297 ;
  assign n2547 = n2546 ^ n2540 ;
  assign n2558 = n2349 & ~n2452 ;
  assign n2557 = n2349 & ~n2439 ;
  assign n2559 = n2558 ^ n2557 ;
  assign n2555 = n2349 & n2431 ;
  assign n2556 = n2356 & n2555 ;
  assign n2560 = n2559 ^ n2556 ;
  assign n2551 = n2325 & ~n2452 ;
  assign n2550 = n2325 & ~n2439 ;
  assign n2552 = n2551 ^ n2550 ;
  assign n2548 = n2325 & n2431 ;
  assign n2549 = n2356 & n2548 ;
  assign n2553 = n2552 ^ n2549 ;
  assign n2554 = n2553 ^ n2325 ;
  assign n2561 = n2560 ^ n2554 ;
  assign n2562 = n2462 ^ n2372 ;
  assign n2563 = n2562 ^ n2455 ;
  assign n2564 = n2476 ^ n2387 ;
  assign n2565 = n2564 ^ n2469 ;
  assign n2566 = n2490 ^ n2407 ;
  assign n2567 = n2566 ^ n2483 ;
  assign n2568 = n2504 ^ n2426 ;
  assign n2569 = n2568 ^ n2497 ;
  assign n2570 = n2518 ^ n2268 ;
  assign n2571 = n2570 ^ n2511 ;
  assign n2572 = n2532 ^ n2286 ;
  assign n2573 = n2572 ^ n2525 ;
  assign n2574 = n2546 ^ n2311 ;
  assign n2575 = n2574 ^ n2539 ;
  assign n2576 = n2560 ^ n2349 ;
  assign n2577 = n2576 ^ n2553 ;
  assign n2580 = n1979 & ~n2137 ;
  assign n2581 = n2580 ^ n2192 ;
  assign n2578 = n2371 ^ n2195 ;
  assign n2579 = n2578 ^ n2364 ;
  assign n2583 = n2581 ^ n2579 ;
  assign n2586 = n2001 & ~n2137 ;
  assign n2587 = n2586 ^ n2197 ;
  assign n2584 = n2386 ^ n2200 ;
  assign n2585 = n2584 ^ n2379 ;
  assign n2591 = n2587 ^ n2585 ;
  assign n2592 = n2583 & n2591 ;
  assign n2593 = n2592 ^ n2583 ;
  assign n2594 = n2593 ^ n2591 ;
  assign n2597 = n2019 & ~n2137 ;
  assign n2598 = n2597 ^ n2211 ;
  assign n2595 = n2406 ^ n2214 ;
  assign n2596 = n2595 ^ n2399 ;
  assign n2600 = n2598 ^ n2596 ;
  assign n2603 = n2032 & ~n2137 ;
  assign n2604 = n2603 ^ n2228 ;
  assign n2601 = n2425 ^ n2231 ;
  assign n2602 = n2601 ^ n2418 ;
  assign n2612 = n2604 ^ n2602 ;
  assign n2613 = n2600 & n2612 ;
  assign n2614 = n2613 ^ n2600 ;
  assign n2615 = n2614 ^ n2612 ;
  assign n2616 = ~n2594 & ~n2615 ;
  assign n2619 = n2046 & ~n2137 ;
  assign n2620 = n2619 ^ n2138 ;
  assign n2617 = n2267 ^ n2141 ;
  assign n2618 = n2617 ^ n2260 ;
  assign n2622 = n2620 ^ n2618 ;
  assign n2625 = n2059 & ~n2137 ;
  assign n2626 = n2625 ^ n2150 ;
  assign n2623 = n2285 ^ n2153 ;
  assign n2624 = n2623 ^ n2278 ;
  assign n2632 = n2626 ^ n2624 ;
  assign n2633 = n2622 & n2632 ;
  assign n2634 = n2633 ^ n2622 ;
  assign n2635 = n2634 ^ n2632 ;
  assign n2638 = n2079 & ~n2137 ;
  assign n2639 = n2638 ^ n2167 ;
  assign n2636 = n2310 ^ n2170 ;
  assign n2637 = n2636 ^ n2303 ;
  assign n2671 = n2639 ^ n2637 ;
  assign n2673 = n2178 & ~n2257 ;
  assign n2672 = n2178 & ~n2244 ;
  assign n2674 = n2673 ^ n2672 ;
  assign n2675 = n2674 ^ n2339 ;
  assign n2676 = n2675 ^ n2178 ;
  assign n2677 = n2676 ^ n2336 ;
  assign n2642 = n2090 & ~n2137 ;
  assign n2643 = n2642 ^ n2175 ;
  assign n2678 = n2677 ^ n2643 ;
  assign n2679 = n2671 & n2678 ;
  assign n2680 = n2679 ^ n2671 ;
  assign n2681 = n2680 ^ n2678 ;
  assign n2682 = ~n2635 & ~n2681 ;
  assign n2683 = n2616 & n2682 ;
  assign n2651 = n2178 & ~n2643 ;
  assign n2655 = ~n2257 & n2651 ;
  assign n2654 = ~n2244 & n2651 ;
  assign n2656 = n2655 ^ n2654 ;
  assign n2652 = n2236 & n2651 ;
  assign n2653 = n2185 & n2652 ;
  assign n2657 = n2656 ^ n2653 ;
  assign n2658 = n2657 ^ n2651 ;
  assign n2644 = n2174 & ~n2643 ;
  assign n2648 = ~n2257 & n2644 ;
  assign n2647 = ~n2244 & n2644 ;
  assign n2649 = n2648 ^ n2647 ;
  assign n2645 = n2236 & n2644 ;
  assign n2646 = n2185 & n2645 ;
  assign n2650 = n2649 ^ n2646 ;
  assign n2659 = n2658 ^ n2650 ;
  assign n2663 = n2303 & n2659 ;
  assign n2662 = n2636 & n2659 ;
  assign n2664 = n2663 ^ n2662 ;
  assign n2660 = n2639 & n2659 ;
  assign n2661 = n2660 ^ n2659 ;
  assign n2665 = n2664 ^ n2661 ;
  assign n2640 = n2637 & n2639 ;
  assign n2641 = n2640 ^ n2637 ;
  assign n2666 = n2665 ^ n2641 ;
  assign n2667 = ~n2635 & n2666 ;
  assign n2627 = n2624 & n2626 ;
  assign n2628 = n2627 ^ n2624 ;
  assign n2629 = n2622 & n2628 ;
  assign n2630 = n2629 ^ n2628 ;
  assign n2621 = n2618 & ~n2620 ;
  assign n2631 = n2630 ^ n2621 ;
  assign n2668 = n2667 ^ n2631 ;
  assign n2669 = n2616 & n2668 ;
  assign n2605 = n2602 & n2604 ;
  assign n2606 = n2605 ^ n2602 ;
  assign n2607 = n2600 & n2606 ;
  assign n2608 = n2607 ^ n2606 ;
  assign n2599 = n2596 & ~n2598 ;
  assign n2609 = n2608 ^ n2599 ;
  assign n2610 = ~n2594 & n2609 ;
  assign n2588 = n2585 & ~n2587 ;
  assign n2589 = ~n2583 & n2588 ;
  assign n2582 = n2579 & ~n2581 ;
  assign n2590 = n2589 ^ n2582 ;
  assign n2611 = n2610 ^ n2590 ;
  assign n2670 = n2669 ^ n2611 ;
  assign n2684 = n2683 ^ n2670 ;
  assign n2687 = n2581 & n2684 ;
  assign n2685 = n2579 & n2684 ;
  assign n2686 = n2685 ^ n2579 ;
  assign n2688 = n2687 ^ n2686 ;
  assign n2691 = n2587 & n2684 ;
  assign n2689 = n2585 & n2684 ;
  assign n2690 = n2689 ^ n2585 ;
  assign n2692 = n2691 ^ n2690 ;
  assign n2695 = n2598 & n2684 ;
  assign n2693 = n2596 & n2684 ;
  assign n2694 = n2693 ^ n2596 ;
  assign n2696 = n2695 ^ n2694 ;
  assign n2699 = n2604 & n2684 ;
  assign n2697 = n2602 & n2684 ;
  assign n2698 = n2697 ^ n2602 ;
  assign n2700 = n2699 ^ n2698 ;
  assign n2703 = n2620 & n2684 ;
  assign n2701 = n2618 & n2684 ;
  assign n2702 = n2701 ^ n2618 ;
  assign n2704 = n2703 ^ n2702 ;
  assign n2707 = n2626 & n2684 ;
  assign n2705 = n2624 & n2684 ;
  assign n2706 = n2705 ^ n2624 ;
  assign n2708 = n2707 ^ n2706 ;
  assign n2711 = n2639 & n2684 ;
  assign n2709 = n2637 & n2684 ;
  assign n2710 = n2709 ^ n2637 ;
  assign n2712 = n2711 ^ n2710 ;
  assign n2715 = n2643 & n2684 ;
  assign n2713 = n2677 & n2684 ;
  assign n2714 = n2713 ^ n2677 ;
  assign n2716 = n2715 ^ n2714 ;
  assign n2717 = n2687 ^ n2581 ;
  assign n2718 = n2717 ^ n2685 ;
  assign n2719 = n2691 ^ n2587 ;
  assign n2720 = n2719 ^ n2689 ;
  assign n2721 = n2695 ^ n2598 ;
  assign n2722 = n2721 ^ n2693 ;
  assign n2723 = n2699 ^ n2604 ;
  assign n2724 = n2723 ^ n2697 ;
  assign n2725 = n2703 ^ n2620 ;
  assign n2726 = n2725 ^ n2701 ;
  assign n2727 = n2707 ^ n2626 ;
  assign n2728 = n2727 ^ n2705 ;
  assign n2729 = n2711 ^ n2639 ;
  assign n2730 = n2729 ^ n2709 ;
  assign n2731 = n2715 ^ n2643 ;
  assign n2732 = n2731 ^ n2713 ;
  assign y0 = n1911 ;
  assign y1 = n1915 ;
  assign y2 = n1919 ;
  assign y3 = n1923 ;
  assign y4 = n1927 ;
  assign y5 = n1931 ;
  assign y6 = n1935 ;
  assign y7 = n1939 ;
  assign y8 = n1941 ;
  assign y9 = n1943 ;
  assign y10 = n1945 ;
  assign y11 = n1947 ;
  assign y12 = n1949 ;
  assign y13 = n1951 ;
  assign y14 = n1953 ;
  assign y15 = n1955 ;
  assign y16 = n2463 ;
  assign y17 = n2477 ;
  assign y18 = n2491 ;
  assign y19 = n2505 ;
  assign y20 = n2519 ;
  assign y21 = n2533 ;
  assign y22 = n2547 ;
  assign y23 = n2561 ;
  assign y24 = n2563 ;
  assign y25 = n2565 ;
  assign y26 = n2567 ;
  assign y27 = n2569 ;
  assign y28 = n2571 ;
  assign y29 = n2573 ;
  assign y30 = n2575 ;
  assign y31 = n2577 ;
  assign y32 = n2688 ;
  assign y33 = n2692 ;
  assign y34 = n2696 ;
  assign y35 = n2700 ;
  assign y36 = n2704 ;
  assign y37 = n2708 ;
  assign y38 = n2712 ;
  assign y39 = n2716 ;
  assign y40 = n2718 ;
  assign y41 = n2720 ;
  assign y42 = n2722 ;
  assign y43 = n2724 ;
  assign y44 = n2726 ;
  assign y45 = n2728 ;
  assign y46 = n2730 ;
  assign y47 = n2732 ;
endmodule
