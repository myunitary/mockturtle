// Benchmark "/tmp/tmp" written by ABC on Sat Nov  8 22:35:29 2025

module mult_32bit_1cc_firstframe ( 
    n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
    n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63  );
  input  n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
    n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
    n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63;
  wire new_n65, new_n66, new_n67, new_n68, new_n69, new_n70, new_n71,
    new_n72, new_n73, new_n74, new_n75, new_n76, new_n77, new_n78, new_n79,
    new_n80, new_n81, new_n82, new_n83, new_n84, new_n85, new_n86, new_n87,
    new_n88, new_n89, new_n90, new_n91, new_n92, new_n93, new_n94, new_n95,
    new_n96, new_n97, new_n98, new_n99, new_n100, new_n101, new_n102,
    new_n103, new_n104, new_n105, new_n106, new_n107, new_n108, new_n109,
    new_n110, new_n111, new_n112, new_n113, new_n114, new_n115, new_n116,
    new_n117, new_n118, new_n119, new_n120, new_n121, new_n122, new_n123,
    new_n124, new_n125, new_n126, new_n127, new_n128, new_n129, new_n130,
    new_n131, new_n132, new_n133, new_n134, new_n135, new_n136, new_n137,
    new_n138, new_n139, new_n140, new_n141, new_n142, new_n143, new_n144,
    new_n145, new_n146, new_n147, new_n148, new_n149, new_n150, new_n151,
    new_n152, new_n153, new_n154, new_n155, new_n156, new_n157, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1456, new_n1457, new_n1458, new_n1459, new_n1460,
    new_n1461, new_n1462, new_n1463, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1469, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1474, new_n1475, new_n1476, new_n1477, new_n1478,
    new_n1479, new_n1480, new_n1481, new_n1482, new_n1483, new_n1484,
    new_n1485, new_n1486, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1557, new_n1558, new_n1559, new_n1560, new_n1561, new_n1562,
    new_n1563, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1580,
    new_n1581, new_n1582, new_n1583, new_n1584, new_n1585, new_n1586,
    new_n1587, new_n1588, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1692, new_n1693, new_n1694,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1725, new_n1726, new_n1727, new_n1728, new_n1729, new_n1730,
    new_n1731, new_n1732, new_n1733, new_n1734, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1746, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1775, new_n1776, new_n1777, new_n1778,
    new_n1779, new_n1780, new_n1781, new_n1782, new_n1783, new_n1784,
    new_n1785, new_n1786, new_n1787, new_n1788, new_n1789, new_n1790,
    new_n1791, new_n1792, new_n1793, new_n1794, new_n1795, new_n1796,
    new_n1797, new_n1798, new_n1799, new_n1800, new_n1801, new_n1802,
    new_n1803, new_n1804, new_n1805, new_n1806, new_n1807, new_n1808,
    new_n1809, new_n1810, new_n1811, new_n1812, new_n1813, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1818, new_n1819, new_n1820,
    new_n1821, new_n1822, new_n1823, new_n1824, new_n1825, new_n1826,
    new_n1827, new_n1828, new_n1829, new_n1830, new_n1831, new_n1832,
    new_n1833, new_n1834, new_n1835, new_n1836, new_n1837, new_n1838,
    new_n1839, new_n1840, new_n1841, new_n1842, new_n1843, new_n1844,
    new_n1845, new_n1846, new_n1847, new_n1848, new_n1849, new_n1850,
    new_n1851, new_n1852, new_n1853, new_n1854, new_n1855, new_n1856,
    new_n1857, new_n1858, new_n1859, new_n1860, new_n1861, new_n1862,
    new_n1863, new_n1864, new_n1865, new_n1866, new_n1867, new_n1868,
    new_n1869, new_n1870, new_n1871, new_n1872, new_n1873, new_n1874,
    new_n1875, new_n1876, new_n1877, new_n1878, new_n1879, new_n1880,
    new_n1881, new_n1882, new_n1883, new_n1884, new_n1885, new_n1886,
    new_n1887, new_n1888, new_n1889, new_n1890, new_n1891, new_n1892,
    new_n1893, new_n1894, new_n1895, new_n1896, new_n1897, new_n1898,
    new_n1899, new_n1900, new_n1901, new_n1902, new_n1903, new_n1904,
    new_n1905, new_n1906, new_n1907, new_n1908, new_n1909, new_n1910,
    new_n1911, new_n1912, new_n1913, new_n1914, new_n1915, new_n1916,
    new_n1917, new_n1918, new_n1919, new_n1920, new_n1921, new_n1922,
    new_n1923, new_n1924, new_n1925, new_n1926, new_n1927, new_n1928,
    new_n1929, new_n1930, new_n1931, new_n1932, new_n1933, new_n1934,
    new_n1935, new_n1936, new_n1937, new_n1938, new_n1939, new_n1940,
    new_n1941, new_n1942, new_n1943, new_n1944, new_n1945, new_n1946,
    new_n1947, new_n1948, new_n1949, new_n1950, new_n1951, new_n1952,
    new_n1953, new_n1954, new_n1955, new_n1956, new_n1957, new_n1958,
    new_n1959, new_n1960, new_n1961, new_n1962, new_n1963, new_n1964,
    new_n1965, new_n1966, new_n1967, new_n1968, new_n1969, new_n1970,
    new_n1971, new_n1972, new_n1973, new_n1974, new_n1975, new_n1976,
    new_n1977, new_n1978, new_n1979, new_n1980, new_n1981, new_n1982,
    new_n1983, new_n1984, new_n1985, new_n1986, new_n1987, new_n1988,
    new_n1989, new_n1990, new_n1991, new_n1992, new_n1993, new_n1994,
    new_n1995, new_n1996, new_n1997, new_n1998, new_n1999, new_n2000,
    new_n2001, new_n2002, new_n2003, new_n2004, new_n2005, new_n2006,
    new_n2007, new_n2008, new_n2009, new_n2010, new_n2011, new_n2012,
    new_n2013, new_n2014, new_n2015, new_n2016, new_n2017, new_n2018,
    new_n2019, new_n2020, new_n2021, new_n2022, new_n2023, new_n2024,
    new_n2025, new_n2026, new_n2027, new_n2028, new_n2029, new_n2030,
    new_n2031, new_n2032, new_n2033, new_n2034, new_n2035, new_n2036,
    new_n2037, new_n2038, new_n2039, new_n2040, new_n2041, new_n2042,
    new_n2043, new_n2044, new_n2045, new_n2046, new_n2047, new_n2048,
    new_n2049, new_n2050, new_n2051, new_n2052, new_n2053, new_n2054,
    new_n2055, new_n2056, new_n2057, new_n2058, new_n2059, new_n2060,
    new_n2061, new_n2062, new_n2063, new_n2064, new_n2065, new_n2066,
    new_n2067, new_n2068, new_n2069, new_n2070, new_n2071, new_n2072,
    new_n2073, new_n2074, new_n2075, new_n2076, new_n2077, new_n2078,
    new_n2079, new_n2080, new_n2081, new_n2082, new_n2083, new_n2084,
    new_n2085, new_n2086, new_n2087, new_n2088, new_n2089, new_n2090,
    new_n2091, new_n2092, new_n2093, new_n2094, new_n2095, new_n2096,
    new_n2097, new_n2098, new_n2099, new_n2100, new_n2101, new_n2102,
    new_n2103, new_n2104, new_n2105, new_n2106, new_n2107, new_n2108,
    new_n2109, new_n2110, new_n2111, new_n2112, new_n2113, new_n2114,
    new_n2115, new_n2116, new_n2117, new_n2118, new_n2119, new_n2120,
    new_n2121, new_n2122, new_n2123, new_n2124, new_n2125, new_n2126,
    new_n2127, new_n2128, new_n2129, new_n2130, new_n2131, new_n2132,
    new_n2133, new_n2134, new_n2135, new_n2136, new_n2137, new_n2138,
    new_n2139, new_n2140, new_n2141, new_n2142, new_n2143, new_n2144,
    new_n2145, new_n2146, new_n2147, new_n2148, new_n2149, new_n2150,
    new_n2151, new_n2152, new_n2153, new_n2154, new_n2155, new_n2156,
    new_n2157, new_n2158, new_n2159, new_n2160, new_n2161, new_n2162,
    new_n2163, new_n2164, new_n2165, new_n2166, new_n2167, new_n2168,
    new_n2169, new_n2170, new_n2171, new_n2172, new_n2173, new_n2174,
    new_n2175, new_n2176, new_n2177, new_n2178, new_n2179, new_n2180,
    new_n2181, new_n2182, new_n2183, new_n2184, new_n2185, new_n2186,
    new_n2187, new_n2188, new_n2189, new_n2190, new_n2191, new_n2192,
    new_n2193, new_n2194, new_n2195, new_n2196, new_n2197, new_n2198,
    new_n2199, new_n2200, new_n2201, new_n2202, new_n2203, new_n2204,
    new_n2205, new_n2206, new_n2207, new_n2208, new_n2209, new_n2210,
    new_n2211, new_n2212, new_n2213, new_n2214, new_n2215, new_n2216,
    new_n2217, new_n2218, new_n2219, new_n2220, new_n2221, new_n2222,
    new_n2223, new_n2224, new_n2225, new_n2226, new_n2227, new_n2228,
    new_n2229, new_n2230, new_n2231, new_n2232, new_n2233, new_n2234,
    new_n2235, new_n2236, new_n2237, new_n2238, new_n2239, new_n2240,
    new_n2241, new_n2242, new_n2243, new_n2244, new_n2245, new_n2246,
    new_n2247, new_n2248, new_n2249, new_n2250, new_n2251, new_n2252,
    new_n2253, new_n2254, new_n2255, new_n2256, new_n2257, new_n2258,
    new_n2259, new_n2260, new_n2261, new_n2262, new_n2263, new_n2264,
    new_n2265, new_n2266, new_n2267, new_n2268, new_n2269, new_n2270,
    new_n2271, new_n2272, new_n2273, new_n2274, new_n2275, new_n2276,
    new_n2277, new_n2278, new_n2279, new_n2280, new_n2281, new_n2282,
    new_n2283, new_n2284, new_n2285, new_n2286, new_n2287, new_n2288,
    new_n2289, new_n2290, new_n2291, new_n2292, new_n2293, new_n2294,
    new_n2295, new_n2296, new_n2297, new_n2298, new_n2299, new_n2300,
    new_n2301, new_n2302, new_n2303, new_n2304, new_n2305, new_n2306,
    new_n2307, new_n2308, new_n2309, new_n2310, new_n2311, new_n2312,
    new_n2313, new_n2314, new_n2315, new_n2316, new_n2317, new_n2318,
    new_n2319, new_n2320, new_n2321, new_n2322, new_n2323, new_n2324,
    new_n2325, new_n2326, new_n2327, new_n2328, new_n2329, new_n2330,
    new_n2331, new_n2332, new_n2333, new_n2334, new_n2335, new_n2336,
    new_n2337, new_n2338, new_n2339, new_n2340, new_n2341, new_n2342,
    new_n2343, new_n2344, new_n2345, new_n2346, new_n2347, new_n2348,
    new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2362, new_n2363, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513, new_n2514, new_n2515, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2551, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577, new_n2578, new_n2579, new_n2580, new_n2581, new_n2582,
    new_n2583, new_n2584, new_n2585, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726,
    new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732,
    new_n2733, new_n2734, new_n2735, new_n2736, new_n2737, new_n2738,
    new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802, new_n2803, new_n2804,
    new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870,
    new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2879, new_n2880, new_n2881, new_n2882,
    new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902, new_n2903, new_n2904, new_n2905, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912,
    new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918,
    new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924,
    new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930,
    new_n2931, new_n2932, new_n2933, new_n2934, new_n2935, new_n2936,
    new_n2937, new_n2938, new_n2939, new_n2940, new_n2941, new_n2942,
    new_n2943, new_n2944, new_n2945, new_n2946, new_n2947, new_n2948,
    new_n2949, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954,
    new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2960,
    new_n2961, new_n2962, new_n2963, new_n2964, new_n2965, new_n2966,
    new_n2967, new_n2968, new_n2969, new_n2970, new_n2971, new_n2972,
    new_n2973, new_n2974, new_n2975, new_n2976, new_n2977, new_n2978,
    new_n2979, new_n2980, new_n2981, new_n2982, new_n2983, new_n2984,
    new_n2985, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990,
    new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996,
    new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3002,
    new_n3003, new_n3004, new_n3005, new_n3006, new_n3007, new_n3008,
    new_n3009, new_n3010, new_n3011, new_n3012, new_n3013, new_n3014,
    new_n3015, new_n3016, new_n3017, new_n3018, new_n3019, new_n3020,
    new_n3021, new_n3022, new_n3023, new_n3024, new_n3025, new_n3026,
    new_n3027, new_n3028, new_n3029, new_n3030, new_n3031, new_n3032,
    new_n3033, new_n3034, new_n3035, new_n3036, new_n3037, new_n3038,
    new_n3039, new_n3040, new_n3041, new_n3042, new_n3043, new_n3044,
    new_n3045, new_n3046, new_n3047, new_n3048, new_n3049, new_n3050,
    new_n3051, new_n3052, new_n3053, new_n3054, new_n3055, new_n3056,
    new_n3057, new_n3058, new_n3059, new_n3060, new_n3061, new_n3062,
    new_n3063, new_n3064, new_n3065, new_n3066, new_n3067, new_n3068,
    new_n3069, new_n3070, new_n3071, new_n3072, new_n3073, new_n3074,
    new_n3075, new_n3076, new_n3077, new_n3078, new_n3079, new_n3080,
    new_n3081, new_n3082, new_n3083, new_n3084, new_n3085, new_n3086,
    new_n3087, new_n3088, new_n3089, new_n3090, new_n3091, new_n3092,
    new_n3093, new_n3094, new_n3095, new_n3096, new_n3097, new_n3098,
    new_n3099, new_n3100, new_n3101, new_n3102, new_n3103, new_n3104,
    new_n3105, new_n3106, new_n3107, new_n3108, new_n3109, new_n3110,
    new_n3111, new_n3112, new_n3113, new_n3114, new_n3115, new_n3116,
    new_n3117, new_n3118, new_n3119, new_n3120, new_n3121, new_n3122,
    new_n3123, new_n3124, new_n3125, new_n3126, new_n3127, new_n3128,
    new_n3129, new_n3130, new_n3131, new_n3132, new_n3133, new_n3134,
    new_n3135, new_n3136, new_n3137, new_n3138, new_n3139, new_n3140,
    new_n3141, new_n3142, new_n3143, new_n3144, new_n3145, new_n3146,
    new_n3147, new_n3148, new_n3149, new_n3150, new_n3151, new_n3152,
    new_n3153, new_n3154, new_n3155, new_n3156, new_n3157, new_n3158,
    new_n3159, new_n3160, new_n3161, new_n3162, new_n3163, new_n3164,
    new_n3165, new_n3166, new_n3167, new_n3168, new_n3169, new_n3170,
    new_n3171, new_n3172, new_n3173, new_n3174, new_n3175, new_n3176,
    new_n3177, new_n3178, new_n3179, new_n3180, new_n3181, new_n3182,
    new_n3183, new_n3184, new_n3185, new_n3186, new_n3187, new_n3188,
    new_n3189, new_n3190, new_n3191, new_n3192, new_n3193, new_n3194,
    new_n3195, new_n3196, new_n3197, new_n3198, new_n3199, new_n3200,
    new_n3201, new_n3202, new_n3203, new_n3204, new_n3205, new_n3206,
    new_n3207, new_n3208, new_n3209, new_n3210, new_n3211, new_n3212,
    new_n3213, new_n3214, new_n3215, new_n3216, new_n3217, new_n3218,
    new_n3219, new_n3220, new_n3221, new_n3222, new_n3223, new_n3224,
    new_n3225, new_n3226, new_n3227, new_n3228, new_n3229, new_n3230,
    new_n3231, new_n3232, new_n3233, new_n3234, new_n3235, new_n3236,
    new_n3237, new_n3238, new_n3239, new_n3240, new_n3241, new_n3242,
    new_n3243, new_n3244, new_n3245, new_n3246, new_n3247, new_n3248,
    new_n3249, new_n3250, new_n3251, new_n3252, new_n3253, new_n3254,
    new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260,
    new_n3261, new_n3262, new_n3263, new_n3264, new_n3265, new_n3266,
    new_n3267, new_n3268, new_n3269, new_n3270, new_n3271, new_n3272,
    new_n3273, new_n3274, new_n3275, new_n3276, new_n3277, new_n3278,
    new_n3279, new_n3280, new_n3281, new_n3282, new_n3283, new_n3284,
    new_n3285, new_n3286, new_n3287, new_n3288, new_n3289, new_n3290,
    new_n3291, new_n3292, new_n3293, new_n3294, new_n3295, new_n3296,
    new_n3297, new_n3298, new_n3299, new_n3300, new_n3301, new_n3302,
    new_n3303, new_n3304, new_n3305, new_n3306, new_n3307, new_n3308,
    new_n3309, new_n3310, new_n3311, new_n3312, new_n3313, new_n3314,
    new_n3315, new_n3316, new_n3317, new_n3318, new_n3319, new_n3320,
    new_n3321, new_n3322, new_n3323, new_n3324, new_n3325, new_n3326,
    new_n3327, new_n3328, new_n3329, new_n3330, new_n3331, new_n3332,
    new_n3333, new_n3334, new_n3335, new_n3336, new_n3337, new_n3338,
    new_n3339, new_n3340, new_n3341, new_n3342, new_n3343, new_n3344,
    new_n3345, new_n3346, new_n3347, new_n3348, new_n3349, new_n3350,
    new_n3351, new_n3352, new_n3353, new_n3354, new_n3355, new_n3356,
    new_n3357, new_n3358, new_n3359, new_n3360, new_n3361, new_n3362,
    new_n3363, new_n3364, new_n3365, new_n3366, new_n3367, new_n3368,
    new_n3369, new_n3370, new_n3371, new_n3372, new_n3373, new_n3374,
    new_n3375, new_n3376, new_n3377, new_n3378, new_n3379, new_n3380,
    new_n3381, new_n3382, new_n3383, new_n3384, new_n3385, new_n3386,
    new_n3387, new_n3388, new_n3389, new_n3390, new_n3391, new_n3392,
    new_n3393, new_n3394, new_n3395, new_n3396, new_n3397, new_n3398,
    new_n3399, new_n3400, new_n3401, new_n3402, new_n3403, new_n3404,
    new_n3405, new_n3406, new_n3407, new_n3408, new_n3409, new_n3410,
    new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416,
    new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425, new_n3426, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458,
    new_n3459, new_n3460, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502, new_n3503, new_n3504, new_n3505, new_n3506,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561, new_n3562, new_n3563, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616, new_n3617, new_n3618, new_n3619, new_n3620,
    new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626,
    new_n3627, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649, new_n3650,
    new_n3651, new_n3652, new_n3653, new_n3654, new_n3655, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3724, new_n3725, new_n3726, new_n3727, new_n3728,
    new_n3729, new_n3730, new_n3731, new_n3732, new_n3733, new_n3734,
    new_n3735, new_n3736, new_n3737, new_n3738, new_n3739, new_n3740,
    new_n3741, new_n3742, new_n3743, new_n3744, new_n3745, new_n3746,
    new_n3747, new_n3748, new_n3749, new_n3750, new_n3751, new_n3752,
    new_n3753, new_n3754, new_n3755, new_n3756, new_n3757, new_n3758,
    new_n3759, new_n3760, new_n3761, new_n3762, new_n3763, new_n3764,
    new_n3765, new_n3766, new_n3767, new_n3768, new_n3769, new_n3770,
    new_n3771, new_n3772, new_n3773, new_n3774, new_n3775, new_n3776,
    new_n3777, new_n3778, new_n3779, new_n3780, new_n3781, new_n3782,
    new_n3783, new_n3784, new_n3785, new_n3786, new_n3787, new_n3788,
    new_n3789, new_n3790, new_n3791, new_n3792, new_n3793, new_n3794,
    new_n3795, new_n3796, new_n3797, new_n3798, new_n3799, new_n3800,
    new_n3801, new_n3802, new_n3803, new_n3804, new_n3805, new_n3806,
    new_n3807, new_n3808, new_n3809, new_n3810, new_n3811, new_n3812,
    new_n3813, new_n3814, new_n3815, new_n3816, new_n3817, new_n3818,
    new_n3819, new_n3820, new_n3821, new_n3822, new_n3823, new_n3824,
    new_n3825, new_n3826, new_n3827, new_n3828, new_n3829, new_n3830,
    new_n3831, new_n3832, new_n3833, new_n3834, new_n3835, new_n3836,
    new_n3837, new_n3838, new_n3839, new_n3840, new_n3841, new_n3842,
    new_n3843, new_n3844, new_n3845, new_n3846, new_n3847, new_n3848,
    new_n3849, new_n3850, new_n3851, new_n3852, new_n3853, new_n3854,
    new_n3855, new_n3856, new_n3857, new_n3858, new_n3859, new_n3860,
    new_n3861, new_n3862, new_n3863, new_n3864, new_n3865, new_n3866,
    new_n3867, new_n3868, new_n3869, new_n3870, new_n3871, new_n3872,
    new_n3873, new_n3874, new_n3875, new_n3876, new_n3877, new_n3878,
    new_n3879, new_n3880, new_n3881, new_n3882, new_n3883, new_n3884,
    new_n3885, new_n3886, new_n3887, new_n3888, new_n3889, new_n3890,
    new_n3891, new_n3892, new_n3893, new_n3894, new_n3895, new_n3896,
    new_n3897, new_n3898, new_n3899, new_n3900, new_n3901, new_n3902,
    new_n3903, new_n3904, new_n3905, new_n3906, new_n3907, new_n3908,
    new_n3909, new_n3910, new_n3911, new_n3912, new_n3913, new_n3914,
    new_n3915, new_n3916, new_n3917, new_n3918, new_n3919, new_n3920,
    new_n3921, new_n3922, new_n3923, new_n3924, new_n3925, new_n3926,
    new_n3927, new_n3928, new_n3929, new_n3930, new_n3931, new_n3932,
    new_n3933, new_n3934, new_n3935, new_n3936, new_n3937, new_n3938,
    new_n3939, new_n3940, new_n3941, new_n3942, new_n3943, new_n3944,
    new_n3945, new_n3946, new_n3947, new_n3948, new_n3949, new_n3950,
    new_n3951, new_n3952, new_n3953, new_n3954, new_n3955, new_n3956,
    new_n3957, new_n3958, new_n3959, new_n3960, new_n3961, new_n3962,
    new_n3963, new_n3964, new_n3965, new_n3966, new_n3967, new_n3968,
    new_n3969, new_n3970, new_n3971, new_n3972, new_n3973, new_n3974,
    new_n3975, new_n3976, new_n3977, new_n3978, new_n3979, new_n3980,
    new_n3981, new_n3982, new_n3983, new_n3984, new_n3985, new_n3986,
    new_n3987, new_n3988, new_n3989, new_n3990, new_n3991, new_n3992,
    new_n3993, new_n3994, new_n3995, new_n3996, new_n3997, new_n3998,
    new_n3999, new_n4000, new_n4001, new_n4002, new_n4003, new_n4004,
    new_n4005, new_n4006, new_n4007, new_n4008, new_n4009, new_n4010,
    new_n4011, new_n4012, new_n4013, new_n4014, new_n4015, new_n4016,
    new_n4017, new_n4018, new_n4019, new_n4020, new_n4021, new_n4022,
    new_n4023, new_n4024, new_n4025, new_n4026, new_n4027, new_n4028,
    new_n4029, new_n4030, new_n4031, new_n4032, new_n4033, new_n4034,
    new_n4035, new_n4036, new_n4037, new_n4038, new_n4039, new_n4040,
    new_n4041, new_n4042, new_n4043, new_n4044, new_n4045, new_n4046,
    new_n4047, new_n4048, new_n4049, new_n4050, new_n4051, new_n4052,
    new_n4053, new_n4054, new_n4055, new_n4056, new_n4057, new_n4058,
    new_n4059, new_n4060, new_n4061, new_n4062, new_n4063, new_n4064,
    new_n4065, new_n4066, new_n4067, new_n4068, new_n4069, new_n4070,
    new_n4071, new_n4072, new_n4073, new_n4074, new_n4075, new_n4076,
    new_n4077, new_n4078, new_n4079, new_n4080, new_n4081, new_n4082,
    new_n4083, new_n4084, new_n4085, new_n4086, new_n4087, new_n4088,
    new_n4089, new_n4090, new_n4091, new_n4092, new_n4093, new_n4094,
    new_n4095, new_n4096, new_n4097, new_n4098, new_n4099, new_n4100,
    new_n4101, new_n4102, new_n4103, new_n4104, new_n4105, new_n4106,
    new_n4107, new_n4108, new_n4109, new_n4110, new_n4111, new_n4112,
    new_n4113, new_n4114, new_n4115, new_n4116, new_n4117, new_n4118,
    new_n4119, new_n4120, new_n4121, new_n4122, new_n4123, new_n4124,
    new_n4125, new_n4126, new_n4127, new_n4128, new_n4129, new_n4130,
    new_n4131, new_n4132, new_n4133, new_n4134, new_n4135, new_n4136,
    new_n4137, new_n4138, new_n4139, new_n4140, new_n4141, new_n4142,
    new_n4143, new_n4144, new_n4145, new_n4146, new_n4147, new_n4148,
    new_n4149, new_n4150, new_n4151, new_n4152, new_n4153, new_n4154,
    new_n4155, new_n4156, new_n4157, new_n4158, new_n4159, new_n4160,
    new_n4161, new_n4162, new_n4163, new_n4164, new_n4165, new_n4166,
    new_n4167, new_n4168, new_n4169, new_n4170, new_n4171, new_n4172,
    new_n4173, new_n4174, new_n4175, new_n4176, new_n4177, new_n4178,
    new_n4179, new_n4180, new_n4181, new_n4182, new_n4183, new_n4184,
    new_n4185, new_n4186, new_n4187, new_n4188, new_n4189, new_n4190,
    new_n4191, new_n4192, new_n4193, new_n4194, new_n4195, new_n4196,
    new_n4197, new_n4198, new_n4199, new_n4200, new_n4201, new_n4202,
    new_n4203, new_n4204, new_n4205, new_n4206, new_n4207, new_n4208,
    new_n4209, new_n4210, new_n4211, new_n4212, new_n4213, new_n4214,
    new_n4215, new_n4216, new_n4217, new_n4218, new_n4219, new_n4220,
    new_n4221, new_n4222, new_n4223, new_n4224, new_n4225, new_n4226,
    new_n4227, new_n4228, new_n4229, new_n4230, new_n4231, new_n4232,
    new_n4233, new_n4234, new_n4235, new_n4236, new_n4237, new_n4238,
    new_n4239, new_n4240, new_n4241, new_n4242, new_n4243, new_n4244,
    new_n4245, new_n4246, new_n4247, new_n4248, new_n4249, new_n4250,
    new_n4251, new_n4252, new_n4253, new_n4254, new_n4255, new_n4256,
    new_n4257, new_n4258, new_n4259, new_n4260, new_n4261, new_n4262,
    new_n4263, new_n4264, new_n4265, new_n4266, new_n4267, new_n4268,
    new_n4269, new_n4270, new_n4271, new_n4272, new_n4273, new_n4274,
    new_n4275, new_n4276, new_n4277, new_n4278, new_n4279, new_n4280,
    new_n4281, new_n4282, new_n4283, new_n4284, new_n4285, new_n4286,
    new_n4287, new_n4288, new_n4289, new_n4290, new_n4291, new_n4292,
    new_n4293, new_n4294, new_n4295, new_n4296, new_n4297, new_n4298,
    new_n4299, new_n4300, new_n4301, new_n4302, new_n4303, new_n4304,
    new_n4305, new_n4306, new_n4307, new_n4308, new_n4309, new_n4310,
    new_n4311, new_n4312, new_n4313, new_n4314, new_n4315, new_n4316,
    new_n4317, new_n4318, new_n4319, new_n4320, new_n4321, new_n4322,
    new_n4323, new_n4324, new_n4325, new_n4326, new_n4327, new_n4328,
    new_n4329, new_n4330, new_n4331, new_n4332, new_n4333, new_n4334,
    new_n4335, new_n4336, new_n4337, new_n4338, new_n4339, new_n4340,
    new_n4341, new_n4342, new_n4343, new_n4344, new_n4345, new_n4346,
    new_n4347, new_n4348, new_n4349, new_n4350, new_n4351, new_n4352,
    new_n4353, new_n4354, new_n4355, new_n4356, new_n4357, new_n4358,
    new_n4359, new_n4360, new_n4361, new_n4362, new_n4363, new_n4364,
    new_n4365, new_n4366, new_n4367, new_n4368, new_n4369, new_n4370,
    new_n4371, new_n4372, new_n4373, new_n4374, new_n4375, new_n4376,
    new_n4377, new_n4378, new_n4379, new_n4380, new_n4381, new_n4382,
    new_n4383, new_n4384, new_n4385, new_n4386, new_n4387, new_n4388,
    new_n4389, new_n4390, new_n4391, new_n4392, new_n4393, new_n4394,
    new_n4395, new_n4396, new_n4397, new_n4398, new_n4399, new_n4400,
    new_n4401, new_n4402, new_n4403, new_n4404, new_n4405, new_n4406,
    new_n4407, new_n4408, new_n4409, new_n4410, new_n4411, new_n4412,
    new_n4413, new_n4414, new_n4415, new_n4416, new_n4417, new_n4418,
    new_n4419, new_n4420, new_n4421, new_n4422, new_n4423, new_n4424,
    new_n4425, new_n4426, new_n4427, new_n4428, new_n4429, new_n4430,
    new_n4431, new_n4432, new_n4433, new_n4434, new_n4435, new_n4436,
    new_n4437, new_n4438, new_n4439, new_n4440, new_n4441, new_n4442,
    new_n4443, new_n4444, new_n4445, new_n4446, new_n4447, new_n4448,
    new_n4449, new_n4450, new_n4451, new_n4452, new_n4453, new_n4454,
    new_n4455, new_n4456, new_n4457, new_n4458, new_n4459, new_n4460,
    new_n4461, new_n4462, new_n4463, new_n4464, new_n4465, new_n4466,
    new_n4467, new_n4468, new_n4469, new_n4470, new_n4471, new_n4472,
    new_n4473, new_n4474, new_n4475, new_n4476, new_n4477, new_n4478,
    new_n4479, new_n4480, new_n4481, new_n4482, new_n4483, new_n4484,
    new_n4485, new_n4486, new_n4487, new_n4488, new_n4489, new_n4490,
    new_n4491, new_n4492, new_n4493, new_n4494, new_n4495, new_n4496,
    new_n4497, new_n4498, new_n4499, new_n4500, new_n4501, new_n4502,
    new_n4503, new_n4504, new_n4505, new_n4506, new_n4507, new_n4508,
    new_n4509, new_n4510, new_n4511, new_n4512, new_n4513, new_n4514,
    new_n4515, new_n4516, new_n4517, new_n4518, new_n4519, new_n4520,
    new_n4521, new_n4522, new_n4523, new_n4524, new_n4525, new_n4526,
    new_n4527, new_n4528, new_n4529, new_n4530, new_n4531, new_n4532,
    new_n4533, new_n4534, new_n4535, new_n4536, new_n4537, new_n4538,
    new_n4539, new_n4540, new_n4541, new_n4542, new_n4543, new_n4544,
    new_n4545, new_n4546, new_n4547, new_n4548, new_n4549, new_n4550,
    new_n4551, new_n4552, new_n4553, new_n4554, new_n4555, new_n4556,
    new_n4557, new_n4558, new_n4559, new_n4560, new_n4561, new_n4562,
    new_n4563, new_n4564, new_n4565, new_n4566, new_n4567, new_n4568,
    new_n4569, new_n4570, new_n4571, new_n4572, new_n4573, new_n4574,
    new_n4575, new_n4576, new_n4577, new_n4578, new_n4579, new_n4580,
    new_n4581, new_n4582, new_n4583, new_n4584, new_n4585, new_n4586,
    new_n4587, new_n4588, new_n4589, new_n4590, new_n4591, new_n4592,
    new_n4593, new_n4594, new_n4595, new_n4596, new_n4597, new_n4598,
    new_n4599, new_n4600, new_n4601, new_n4602, new_n4603, new_n4604,
    new_n4605, new_n4606, new_n4607, new_n4608, new_n4609, new_n4610,
    new_n4611, new_n4612, new_n4613, new_n4614, new_n4615, new_n4616,
    new_n4617, new_n4618, new_n4619, new_n4620, new_n4621, new_n4622,
    new_n4623, new_n4624, new_n4625, new_n4626, new_n4627, new_n4628,
    new_n4629, new_n4630, new_n4631, new_n4632, new_n4633, new_n4634,
    new_n4635, new_n4636, new_n4637, new_n4638, new_n4639, new_n4640,
    new_n4641, new_n4642, new_n4643, new_n4644, new_n4645, new_n4646,
    new_n4647, new_n4648, new_n4649, new_n4650, new_n4651, new_n4652,
    new_n4653, new_n4654, new_n4655, new_n4656, new_n4657, new_n4658,
    new_n4659, new_n4660, new_n4661, new_n4662, new_n4663, new_n4664,
    new_n4665, new_n4666, new_n4667, new_n4668, new_n4669, new_n4670,
    new_n4671, new_n4672, new_n4673, new_n4674, new_n4675, new_n4676,
    new_n4677, new_n4678, new_n4679, new_n4680, new_n4681, new_n4682,
    new_n4683, new_n4684, new_n4685, new_n4686, new_n4687, new_n4688,
    new_n4689, new_n4690, new_n4691, new_n4692, new_n4693, new_n4694,
    new_n4695, new_n4696, new_n4697, new_n4698, new_n4699, new_n4700,
    new_n4701, new_n4702, new_n4703, new_n4704, new_n4705, new_n4706,
    new_n4707, new_n4708, new_n4709, new_n4710, new_n4711, new_n4712,
    new_n4713, new_n4714, new_n4715, new_n4716, new_n4717, new_n4718,
    new_n4719, new_n4720, new_n4721, new_n4722, new_n4723, new_n4724,
    new_n4725, new_n4726, new_n4727, new_n4728, new_n4729, new_n4730,
    new_n4731, new_n4732, new_n4733, new_n4734, new_n4735, new_n4736,
    new_n4737, new_n4738, new_n4739, new_n4740, new_n4741, new_n4742,
    new_n4743, new_n4744, new_n4745, new_n4746, new_n4747, new_n4748,
    new_n4749, new_n4750, new_n4751, new_n4752, new_n4753, new_n4754,
    new_n4755, new_n4756, new_n4757, new_n4758, new_n4759, new_n4760,
    new_n4761, new_n4762, new_n4763, new_n4764, new_n4765, new_n4766,
    new_n4767, new_n4768, new_n4769, new_n4770, new_n4771, new_n4772,
    new_n4773, new_n4774, new_n4775, new_n4776, new_n4777, new_n4778,
    new_n4779, new_n4780, new_n4781, new_n4782, new_n4783, new_n4784,
    new_n4785, new_n4786, new_n4787, new_n4788, new_n4789, new_n4790,
    new_n4791, new_n4792, new_n4793, new_n4794, new_n4795, new_n4796,
    new_n4797, new_n4798, new_n4799, new_n4800, new_n4801, new_n4802,
    new_n4803, new_n4804, new_n4805, new_n4806, new_n4807, new_n4808,
    new_n4809, new_n4810, new_n4811, new_n4812, new_n4813, new_n4814,
    new_n4815, new_n4816, new_n4817, new_n4818, new_n4819, new_n4820,
    new_n4821, new_n4822, new_n4823, new_n4824, new_n4825, new_n4826,
    new_n4827, new_n4828, new_n4829, new_n4830, new_n4831, new_n4832,
    new_n4833, new_n4834, new_n4835, new_n4836, new_n4837, new_n4838,
    new_n4839, new_n4840, new_n4841, new_n4842, new_n4843, new_n4844,
    new_n4845, new_n4846, new_n4847, new_n4848, new_n4849, new_n4850,
    new_n4851, new_n4852, new_n4853, new_n4854, new_n4855, new_n4856,
    new_n4857, new_n4858, new_n4859, new_n4860, new_n4861, new_n4862,
    new_n4863, new_n4864, new_n4865, new_n4866, new_n4867, new_n4868,
    new_n4869, new_n4870, new_n4871, new_n4872, new_n4873, new_n4874,
    new_n4875, new_n4876, new_n4877, new_n4878, new_n4879, new_n4880,
    new_n4881, new_n4882, new_n4883, new_n4884, new_n4885, new_n4886,
    new_n4887, new_n4888, new_n4889, new_n4890, new_n4891, new_n4892,
    new_n4893, new_n4894, new_n4895, new_n4896, new_n4897, new_n4898,
    new_n4899, new_n4900, new_n4901, new_n4902, new_n4903, new_n4904,
    new_n4905, new_n4906, new_n4907, new_n4908, new_n4909, new_n4910,
    new_n4911, new_n4912, new_n4913, new_n4914, new_n4915, new_n4916,
    new_n4917, new_n4918, new_n4919, new_n4920, new_n4921, new_n4922,
    new_n4923, new_n4924, new_n4925, new_n4926, new_n4927, new_n4928,
    new_n4929, new_n4930, new_n4931, new_n4932, new_n4933, new_n4934,
    new_n4935, new_n4936, new_n4937, new_n4938, new_n4939, new_n4940,
    new_n4941, new_n4942, new_n4943, new_n4944, new_n4945, new_n4946,
    new_n4947, new_n4948, new_n4949, new_n4950, new_n4951, new_n4952,
    new_n4953, new_n4954, new_n4955, new_n4956, new_n4957, new_n4958,
    new_n4959, new_n4960, new_n4961, new_n4962, new_n4963, new_n4964,
    new_n4965, new_n4966, new_n4967, new_n4968, new_n4969, new_n4970,
    new_n4971, new_n4972, new_n4973, new_n4974, new_n4975, new_n4976,
    new_n4977, new_n4978, new_n4979, new_n4980, new_n4981, new_n4982,
    new_n4983, new_n4984, new_n4985, new_n4986, new_n4987, new_n4988,
    new_n4989, new_n4990, new_n4991, new_n4992, new_n4993, new_n4994,
    new_n4995, new_n4996, new_n4997, new_n4998, new_n4999, new_n5000,
    new_n5001, new_n5002, new_n5003, new_n5004, new_n5005, new_n5006,
    new_n5007, new_n5008, new_n5009, new_n5010, new_n5011, new_n5012,
    new_n5013, new_n5014, new_n5015, new_n5016, new_n5017, new_n5018,
    new_n5019, new_n5020, new_n5021, new_n5022, new_n5023, new_n5024,
    new_n5025, new_n5026, new_n5027, new_n5028, new_n5029, new_n5030,
    new_n5031, new_n5032, new_n5033, new_n5034, new_n5035, new_n5036,
    new_n5037, new_n5038, new_n5039, new_n5040, new_n5041, new_n5042,
    new_n5043, new_n5044, new_n5045, new_n5046, new_n5047, new_n5048,
    new_n5049, new_n5050, new_n5051, new_n5052, new_n5053, new_n5054,
    new_n5055, new_n5056, new_n5057, new_n5058, new_n5059, new_n5060,
    new_n5061, new_n5062, new_n5063, new_n5064, new_n5065, new_n5066,
    new_n5067, new_n5068, new_n5069, new_n5070, new_n5071, new_n5072,
    new_n5073, new_n5074, new_n5075, new_n5076, new_n5077, new_n5078,
    new_n5079, new_n5080, new_n5081, new_n5082, new_n5083, new_n5084,
    new_n5085, new_n5086, new_n5087, new_n5088, new_n5089, new_n5090,
    new_n5091, new_n5092, new_n5093, new_n5094, new_n5095, new_n5096,
    new_n5097, new_n5098, new_n5099, new_n5100, new_n5101, new_n5102,
    new_n5103, new_n5104, new_n5105, new_n5106, new_n5107, new_n5108,
    new_n5109, new_n5110, new_n5111, new_n5112, new_n5113, new_n5114,
    new_n5115, new_n5116, new_n5117, new_n5118, new_n5119, new_n5120,
    new_n5121, new_n5122, new_n5123, new_n5124, new_n5125, new_n5126,
    new_n5127, new_n5128, new_n5129, new_n5130, new_n5131, new_n5132,
    new_n5133, new_n5134, new_n5135, new_n5136, new_n5137, new_n5138,
    new_n5139, new_n5140, new_n5141, new_n5142, new_n5143, new_n5144,
    new_n5145, new_n5146, new_n5147, new_n5148, new_n5149, new_n5150,
    new_n5151, new_n5152, new_n5153, new_n5154, new_n5155, new_n5156,
    new_n5157, new_n5158, new_n5159, new_n5160, new_n5161, new_n5162,
    new_n5163, new_n5164, new_n5165, new_n5166, new_n5167, new_n5168,
    new_n5169, new_n5170, new_n5171, new_n5172, new_n5173, new_n5174,
    new_n5175, new_n5176, new_n5177, new_n5178, new_n5179, new_n5180,
    new_n5181, new_n5182, new_n5183, new_n5184, new_n5185, new_n5186,
    new_n5187, new_n5188, new_n5189, new_n5190, new_n5191, new_n5192,
    new_n5193, new_n5194, new_n5195, new_n5196, new_n5197, new_n5198,
    new_n5199, new_n5200, new_n5201, new_n5202, new_n5203, new_n5204,
    new_n5205, new_n5206, new_n5207, new_n5208, new_n5209, new_n5210,
    new_n5211, new_n5212, new_n5213, new_n5214, new_n5215, new_n5216,
    new_n5217, new_n5218, new_n5219, new_n5220, new_n5221, new_n5222,
    new_n5223, new_n5224, new_n5225, new_n5226, new_n5227, new_n5228,
    new_n5229, new_n5230, new_n5231, new_n5232, new_n5233, new_n5234,
    new_n5235, new_n5236, new_n5237, new_n5238, new_n5239, new_n5240,
    new_n5241, new_n5242, new_n5243, new_n5244, new_n5245, new_n5246,
    new_n5247, new_n5248, new_n5249, new_n5250, new_n5251, new_n5252,
    new_n5253, new_n5254, new_n5255, new_n5256, new_n5257, new_n5258,
    new_n5259, new_n5260, new_n5261, new_n5262, new_n5263, new_n5264,
    new_n5265, new_n5266, new_n5267, new_n5268, new_n5269, new_n5270,
    new_n5271, new_n5272, new_n5273, new_n5274, new_n5275, new_n5276,
    new_n5277, new_n5278, new_n5279, new_n5280, new_n5281, new_n5282,
    new_n5283, new_n5284, new_n5285, new_n5286, new_n5287, new_n5288,
    new_n5289, new_n5290, new_n5291, new_n5292, new_n5293, new_n5294,
    new_n5295, new_n5296, new_n5297, new_n5298, new_n5299, new_n5300,
    new_n5301, new_n5302, new_n5303, new_n5304, new_n5305, new_n5306,
    new_n5307, new_n5308, new_n5309, new_n5310, new_n5311, new_n5312,
    new_n5313, new_n5314, new_n5315, new_n5316, new_n5317, new_n5318,
    new_n5319, new_n5320, new_n5321, new_n5322, new_n5323, new_n5324,
    new_n5325, new_n5326, new_n5327, new_n5328, new_n5329, new_n5330,
    new_n5331, new_n5332, new_n5333, new_n5334, new_n5335, new_n5336,
    new_n5337, new_n5338, new_n5339, new_n5340, new_n5341, new_n5342,
    new_n5343, new_n5344, new_n5345, new_n5346, new_n5347, new_n5348,
    new_n5349, new_n5350, new_n5351, new_n5352, new_n5353, new_n5354,
    new_n5355, new_n5356, new_n5357, new_n5358, new_n5359, new_n5360,
    new_n5361, new_n5362, new_n5363, new_n5364, new_n5365, new_n5366,
    new_n5367, new_n5368, new_n5369, new_n5370, new_n5371, new_n5372,
    new_n5373, new_n5374, new_n5375, new_n5376, new_n5377, new_n5378,
    new_n5379, new_n5380, new_n5381, new_n5382, new_n5383, new_n5384,
    new_n5385, new_n5386, new_n5387, new_n5388, new_n5389, new_n5390,
    new_n5391, new_n5392, new_n5393, new_n5394, new_n5395, new_n5396,
    new_n5397, new_n5398, new_n5399, new_n5400, new_n5401, new_n5402,
    new_n5403, new_n5404, new_n5405, new_n5406, new_n5407, new_n5408,
    new_n5409, new_n5410, new_n5411, new_n5412, new_n5413, new_n5414,
    new_n5415, new_n5416, new_n5417, new_n5418, new_n5419, new_n5420,
    new_n5421, new_n5422, new_n5423, new_n5424, new_n5425, new_n5426,
    new_n5427, new_n5428, new_n5429, new_n5430, new_n5431, new_n5432,
    new_n5433, new_n5434, new_n5435, new_n5436, new_n5437, new_n5438,
    new_n5439, new_n5440, new_n5441, new_n5442, new_n5443, new_n5444,
    new_n5445, new_n5446, new_n5447, new_n5448, new_n5449, new_n5450,
    new_n5451, new_n5452, new_n5453, new_n5454, new_n5455, new_n5456,
    new_n5457, new_n5458, new_n5459, new_n5460, new_n5461, new_n5462,
    new_n5463, new_n5464, new_n5465, new_n5466, new_n5467, new_n5468,
    new_n5469, new_n5470, new_n5471, new_n5472, new_n5473, new_n5474,
    new_n5475, new_n5476, new_n5477, new_n5478, new_n5479, new_n5480,
    new_n5481, new_n5482, new_n5483, new_n5484, new_n5485, new_n5486,
    new_n5487, new_n5488, new_n5489, new_n5490, new_n5491, new_n5492,
    new_n5493, new_n5494, new_n5495, new_n5496, new_n5497, new_n5498,
    new_n5499, new_n5500, new_n5501, new_n5502, new_n5503, new_n5504,
    new_n5505, new_n5506, new_n5507, new_n5508, new_n5509, new_n5510,
    new_n5511, new_n5512, new_n5513, new_n5514, new_n5515, new_n5516,
    new_n5517, new_n5518, new_n5519, new_n5520, new_n5521, new_n5522,
    new_n5523, new_n5524, new_n5525, new_n5526, new_n5527, new_n5528,
    new_n5529, new_n5530, new_n5531, new_n5532, new_n5533, new_n5534,
    new_n5535, new_n5536, new_n5537, new_n5538, new_n5539, new_n5540,
    new_n5541, new_n5542, new_n5543, new_n5544, new_n5545, new_n5546,
    new_n5547, new_n5548, new_n5549, new_n5550, new_n5551, new_n5552,
    new_n5553, new_n5554, new_n5555, new_n5556, new_n5557, new_n5558,
    new_n5559, new_n5560, new_n5561, new_n5562, new_n5563, new_n5564,
    new_n5565, new_n5566, new_n5567, new_n5568, new_n5569, new_n5570,
    new_n5571, new_n5572, new_n5573, new_n5574, new_n5575, new_n5576,
    new_n5577, new_n5578, new_n5579, new_n5580, new_n5581, new_n5582,
    new_n5583, new_n5584, new_n5585, new_n5586, new_n5587, new_n5588,
    new_n5589, new_n5590, new_n5591, new_n5592, new_n5593, new_n5594,
    new_n5595, new_n5596, new_n5597, new_n5598, new_n5599, new_n5600,
    new_n5601, new_n5602, new_n5603, new_n5604, new_n5605, new_n5606,
    new_n5607, new_n5608, new_n5609, new_n5610, new_n5611, new_n5612,
    new_n5613, new_n5614, new_n5615, new_n5616, new_n5617, new_n5618,
    new_n5619, new_n5620, new_n5621, new_n5622, new_n5623, new_n5624,
    new_n5625, new_n5626, new_n5627, new_n5628, new_n5629, new_n5630,
    new_n5631, new_n5632, new_n5633, new_n5634, new_n5635, new_n5636,
    new_n5637, new_n5638, new_n5639, new_n5640, new_n5641, new_n5642,
    new_n5643, new_n5644, new_n5645, new_n5646, new_n5647, new_n5648,
    new_n5649, new_n5650, new_n5651, new_n5652, new_n5653, new_n5654,
    new_n5655, new_n5656, new_n5657, new_n5658, new_n5659, new_n5660,
    new_n5661, new_n5662, new_n5663, new_n5664, new_n5665, new_n5666,
    new_n5667, new_n5668, new_n5669, new_n5670, new_n5671, new_n5672,
    new_n5673, new_n5674, new_n5675, new_n5676, new_n5677, new_n5678,
    new_n5679, new_n5680, new_n5681, new_n5682, new_n5683, new_n5684,
    new_n5685, new_n5686, new_n5687, new_n5688, new_n5689, new_n5690,
    new_n5691, new_n5692, new_n5693, new_n5694, new_n5695, new_n5696,
    new_n5697, new_n5698, new_n5699, new_n5700, new_n5701, new_n5702,
    new_n5703, new_n5704, new_n5705, new_n5706, new_n5707, new_n5708,
    new_n5709, new_n5710, new_n5711, new_n5712, new_n5713, new_n5714,
    new_n5715, new_n5716, new_n5717, new_n5718, new_n5719, new_n5720,
    new_n5721, new_n5722, new_n5723, new_n5724, new_n5725, new_n5726,
    new_n5727, new_n5728, new_n5729, new_n5730, new_n5731, new_n5732,
    new_n5733, new_n5734, new_n5735, new_n5736, new_n5737, new_n5738,
    new_n5739, new_n5740, new_n5741, new_n5742, new_n5743, new_n5744,
    new_n5745, new_n5746, new_n5747, new_n5748, new_n5749, new_n5750,
    new_n5751, new_n5752, new_n5753, new_n5754, new_n5755, new_n5756,
    new_n5757, new_n5758, new_n5759, new_n5760, new_n5761, new_n5762,
    new_n5763, new_n5764, new_n5765, new_n5766, new_n5767, new_n5768,
    new_n5769, new_n5770, new_n5771, new_n5772, new_n5773, new_n5774,
    new_n5775, new_n5776, new_n5777, new_n5778, new_n5779, new_n5780,
    new_n5781, new_n5782, new_n5783, new_n5784, new_n5785, new_n5786,
    new_n5787, new_n5788, new_n5789, new_n5790, new_n5791, new_n5792,
    new_n5793, new_n5794, new_n5795, new_n5796, new_n5797, new_n5798,
    new_n5799, new_n5800, new_n5801, new_n5802, new_n5803, new_n5804,
    new_n5805, new_n5806, new_n5807, new_n5808, new_n5809, new_n5810,
    new_n5811, new_n5812, new_n5813, new_n5814, new_n5815, new_n5816,
    new_n5817, new_n5818, new_n5819, new_n5820, new_n5821, new_n5822,
    new_n5823, new_n5824, new_n5825, new_n5826, new_n5827, new_n5828,
    new_n5829, new_n5830, new_n5831, new_n5832, new_n5833, new_n5834,
    new_n5835, new_n5836, new_n5837, new_n5838, new_n5839, new_n5840,
    new_n5841, new_n5842, new_n5843, new_n5844, new_n5845, new_n5846,
    new_n5847, new_n5848, new_n5849, new_n5850, new_n5851, new_n5852,
    new_n5853, new_n5854, new_n5855, new_n5856, new_n5857, new_n5858,
    new_n5859, new_n5860, new_n5861, new_n5862, new_n5863, new_n5864,
    new_n5865, new_n5866, new_n5867, new_n5868, new_n5869, new_n5870,
    new_n5871, new_n5872, new_n5873, new_n5874, new_n5875, new_n5876,
    new_n5877, new_n5878, new_n5879, new_n5880, new_n5881, new_n5882,
    new_n5883, new_n5884, new_n5885, new_n5886, new_n5887, new_n5888,
    new_n5889, new_n5890, new_n5891, new_n5892, new_n5893, new_n5894,
    new_n5895, new_n5896, new_n5897, new_n5898, new_n5899, new_n5900,
    new_n5901, new_n5902, new_n5903, new_n5904, new_n5905, new_n5906,
    new_n5907, new_n5908, new_n5909, new_n5910, new_n5911, new_n5912,
    new_n5913, new_n5914, new_n5915, new_n5916, new_n5917, new_n5918,
    new_n5919, new_n5920, new_n5921, new_n5922, new_n5923, new_n5924,
    new_n5925, new_n5926, new_n5927, new_n5928, new_n5929, new_n5930,
    new_n5931, new_n5932, new_n5933, new_n5934, new_n5935, new_n5936,
    new_n5937, new_n5938, new_n5939, new_n5940, new_n5941, new_n5942,
    new_n5943, new_n5944, new_n5945, new_n5946, new_n5947, new_n5948,
    new_n5949, new_n5950, new_n5951, new_n5952, new_n5953, new_n5954,
    new_n5955, new_n5956, new_n5957, new_n5958, new_n5959, new_n5960,
    new_n5961, new_n5962, new_n5963, new_n5964, new_n5965, new_n5966,
    new_n5967, new_n5968, new_n5969, new_n5970, new_n5971, new_n5972,
    new_n5973, new_n5974, new_n5975, new_n5976, new_n5977, new_n5978,
    new_n5979, new_n5980, new_n5981, new_n5982, new_n5983, new_n5984,
    new_n5985, new_n5986, new_n5987, new_n5988, new_n5989, new_n5990,
    new_n5991, new_n5992, new_n5993, new_n5994, new_n5995, new_n5996,
    new_n5997, new_n5998, new_n5999, new_n6000, new_n6001, new_n6002,
    new_n6003, new_n6004, new_n6005, new_n6006, new_n6007, new_n6008,
    new_n6009, new_n6010, new_n6011, new_n6012, new_n6013, new_n6014,
    new_n6015, new_n6016, new_n6017, new_n6018, new_n6019, new_n6020,
    new_n6021, new_n6022, new_n6023, new_n6024, new_n6025, new_n6026,
    new_n6027, new_n6028, new_n6029, new_n6030, new_n6031, new_n6032,
    new_n6033, new_n6034, new_n6035, new_n6036, new_n6037, new_n6038,
    new_n6039, new_n6040, new_n6041, new_n6042, new_n6043;
  assign new_n65 = n32 & n34;
  assign new_n66 = n31 & n35;
  assign new_n67 = new_n65 & new_n66;
  assign new_n68 = n31 & n34;
  assign new_n69 = n32 & n33;
  assign new_n70 = new_n69 ^ new_n68;
  assign new_n71 = new_n70 ^ new_n67;
  assign new_n72 = n30 & n35;
  assign new_n73 = new_n72 ^ new_n67;
  assign new_n74 = ~new_n73 & new_n71;
  assign new_n75 = new_n74 ^ new_n70;
  assign new_n76 = n30 & n34;
  assign new_n77 = n31 & n33;
  assign new_n78 = ~new_n65 & new_n77;
  assign new_n79 = new_n78 ^ new_n76;
  assign new_n80 = new_n79 ^ new_n75;
  assign new_n81 = n29 & n35;
  assign new_n82 = new_n81 ^ new_n75;
  assign new_n83 = ~new_n80 & new_n82;
  assign new_n84 = new_n83 ^ new_n81;
  assign new_n85 = n29 & n34;
  assign new_n86 = n30 & n33;
  assign new_n87 = ~new_n76 & new_n78;
  assign new_n88 = new_n87 ^ new_n77;
  assign new_n89 = new_n88 ^ new_n86;
  assign new_n90 = new_n89 ^ new_n85;
  assign new_n91 = new_n90 ^ new_n84;
  assign new_n92 = n28 & n35;
  assign new_n93 = new_n92 ^ new_n84;
  assign new_n94 = ~new_n93 & new_n91;
  assign new_n95 = new_n94 ^ new_n90;
  assign new_n96 = n28 & n34;
  assign new_n97 = new_n88 ^ new_n85;
  assign new_n98 = ~new_n97 & new_n89;
  assign new_n99 = new_n98 ^ new_n86;
  assign new_n100 = n29 & n33;
  assign new_n101 = new_n100 ^ new_n99;
  assign new_n102 = new_n101 ^ new_n96;
  assign new_n103 = new_n102 ^ new_n95;
  assign new_n104 = n27 & n35;
  assign new_n105 = new_n104 ^ new_n95;
  assign new_n106 = ~new_n103 & new_n105;
  assign new_n107 = new_n106 ^ new_n104;
  assign new_n108 = n27 & n34;
  assign new_n109 = new_n100 ^ new_n96;
  assign new_n110 = ~new_n101 & new_n109;
  assign new_n111 = new_n110 ^ new_n96;
  assign new_n112 = n28 & n33;
  assign new_n113 = new_n112 ^ new_n111;
  assign new_n114 = new_n113 ^ new_n108;
  assign new_n115 = new_n114 ^ new_n107;
  assign new_n116 = n26 & n35;
  assign new_n117 = new_n116 ^ new_n107;
  assign new_n118 = ~new_n117 & new_n115;
  assign new_n119 = new_n118 ^ new_n114;
  assign new_n120 = n26 & n34;
  assign new_n121 = new_n112 ^ new_n108;
  assign new_n122 = ~new_n113 & new_n121;
  assign new_n123 = new_n122 ^ new_n108;
  assign new_n124 = n27 & n33;
  assign new_n125 = new_n124 ^ new_n123;
  assign new_n126 = new_n125 ^ new_n120;
  assign new_n127 = new_n126 ^ new_n119;
  assign new_n128 = n25 & n35;
  assign new_n129 = new_n128 ^ new_n119;
  assign new_n130 = ~new_n127 & new_n129;
  assign new_n131 = new_n130 ^ new_n128;
  assign new_n132 = n25 & n34;
  assign new_n133 = new_n124 ^ new_n120;
  assign new_n134 = ~new_n125 & new_n133;
  assign new_n135 = new_n134 ^ new_n120;
  assign new_n136 = n26 & n33;
  assign new_n137 = new_n136 ^ new_n135;
  assign new_n138 = new_n137 ^ new_n132;
  assign new_n139 = new_n138 ^ new_n131;
  assign new_n140 = n24 & n35;
  assign new_n141 = new_n140 ^ new_n131;
  assign new_n142 = ~new_n141 & new_n139;
  assign new_n143 = new_n142 ^ new_n138;
  assign new_n144 = n24 & n34;
  assign new_n145 = new_n136 ^ new_n132;
  assign new_n146 = ~new_n137 & new_n145;
  assign new_n147 = new_n146 ^ new_n132;
  assign new_n148 = n25 & n33;
  assign new_n149 = new_n148 ^ new_n147;
  assign new_n150 = new_n149 ^ new_n144;
  assign new_n151 = new_n150 ^ new_n143;
  assign new_n152 = n23 & n35;
  assign new_n153 = new_n152 ^ new_n143;
  assign new_n154 = ~new_n151 & new_n153;
  assign new_n155 = new_n154 ^ new_n152;
  assign new_n156 = n23 & n34;
  assign new_n157 = new_n148 ^ new_n144;
  assign new_n158 = ~new_n149 & new_n157;
  assign new_n159 = new_n158 ^ new_n144;
  assign new_n160 = n24 & n33;
  assign new_n161 = new_n160 ^ new_n159;
  assign new_n162 = new_n161 ^ new_n156;
  assign new_n163 = new_n162 ^ new_n155;
  assign new_n164 = n22 & n35;
  assign new_n165 = new_n164 ^ new_n155;
  assign new_n166 = ~new_n165 & new_n163;
  assign new_n167 = new_n166 ^ new_n162;
  assign new_n168 = n22 & n34;
  assign new_n169 = new_n160 ^ new_n156;
  assign new_n170 = ~new_n161 & new_n169;
  assign new_n171 = new_n170 ^ new_n156;
  assign new_n172 = n23 & n33;
  assign new_n173 = new_n172 ^ new_n171;
  assign new_n174 = new_n173 ^ new_n168;
  assign new_n175 = new_n174 ^ new_n167;
  assign new_n176 = n21 & n35;
  assign new_n177 = new_n176 ^ new_n167;
  assign new_n178 = ~new_n175 & new_n177;
  assign new_n179 = new_n178 ^ new_n176;
  assign new_n180 = n21 & n34;
  assign new_n181 = new_n172 ^ new_n168;
  assign new_n182 = ~new_n173 & new_n181;
  assign new_n183 = new_n182 ^ new_n168;
  assign new_n184 = n22 & n33;
  assign new_n185 = new_n184 ^ new_n183;
  assign new_n186 = new_n185 ^ new_n180;
  assign new_n187 = new_n186 ^ new_n179;
  assign new_n188 = n20 & n35;
  assign new_n189 = new_n188 ^ new_n179;
  assign new_n190 = ~new_n189 & new_n187;
  assign new_n191 = new_n190 ^ new_n186;
  assign new_n192 = n20 & n34;
  assign new_n193 = new_n184 ^ new_n180;
  assign new_n194 = ~new_n185 & new_n193;
  assign new_n195 = new_n194 ^ new_n180;
  assign new_n196 = n21 & n33;
  assign new_n197 = new_n196 ^ new_n195;
  assign new_n198 = new_n197 ^ new_n192;
  assign new_n199 = new_n198 ^ new_n191;
  assign new_n200 = n19 & n35;
  assign new_n201 = new_n200 ^ new_n191;
  assign new_n202 = ~new_n199 & new_n201;
  assign new_n203 = new_n202 ^ new_n200;
  assign new_n204 = n19 & n34;
  assign new_n205 = new_n196 ^ new_n192;
  assign new_n206 = ~new_n197 & new_n205;
  assign new_n207 = new_n206 ^ new_n192;
  assign new_n208 = n20 & n33;
  assign new_n209 = new_n208 ^ new_n207;
  assign new_n210 = new_n209 ^ new_n204;
  assign new_n211 = new_n210 ^ new_n203;
  assign new_n212 = n18 & n35;
  assign new_n213 = new_n212 ^ new_n203;
  assign new_n214 = ~new_n213 & new_n211;
  assign new_n215 = new_n214 ^ new_n210;
  assign new_n216 = n18 & n34;
  assign new_n217 = new_n208 ^ new_n204;
  assign new_n218 = ~new_n209 & new_n217;
  assign new_n219 = new_n218 ^ new_n204;
  assign new_n220 = n19 & n33;
  assign new_n221 = new_n220 ^ new_n219;
  assign new_n222 = new_n221 ^ new_n216;
  assign new_n223 = new_n222 ^ new_n215;
  assign new_n224 = n17 & n35;
  assign new_n225 = new_n224 ^ new_n215;
  assign new_n226 = ~new_n223 & new_n225;
  assign new_n227 = new_n226 ^ new_n224;
  assign new_n228 = n17 & n34;
  assign new_n229 = new_n220 ^ new_n216;
  assign new_n230 = ~new_n221 & new_n229;
  assign new_n231 = new_n230 ^ new_n216;
  assign new_n232 = n18 & n33;
  assign new_n233 = new_n232 ^ new_n231;
  assign new_n234 = new_n233 ^ new_n228;
  assign new_n235 = new_n234 ^ new_n227;
  assign new_n236 = n16 & n35;
  assign new_n237 = new_n236 ^ new_n227;
  assign new_n238 = ~new_n237 & new_n235;
  assign new_n239 = new_n238 ^ new_n234;
  assign new_n240 = n16 & n34;
  assign new_n241 = new_n232 ^ new_n228;
  assign new_n242 = ~new_n233 & new_n241;
  assign new_n243 = new_n242 ^ new_n228;
  assign new_n244 = n17 & n33;
  assign new_n245 = new_n244 ^ new_n243;
  assign new_n246 = new_n245 ^ new_n240;
  assign new_n247 = new_n246 ^ new_n239;
  assign new_n248 = n15 & n35;
  assign new_n249 = new_n248 ^ new_n239;
  assign new_n250 = ~new_n247 & new_n249;
  assign new_n251 = new_n250 ^ new_n248;
  assign new_n252 = n15 & n34;
  assign new_n253 = new_n244 ^ new_n240;
  assign new_n254 = ~new_n245 & new_n253;
  assign new_n255 = new_n254 ^ new_n240;
  assign new_n256 = n16 & n33;
  assign new_n257 = new_n256 ^ new_n255;
  assign new_n258 = new_n257 ^ new_n252;
  assign new_n259 = new_n258 ^ new_n251;
  assign new_n260 = n14 & n35;
  assign new_n261 = new_n260 ^ new_n251;
  assign new_n262 = ~new_n261 & new_n259;
  assign new_n263 = new_n262 ^ new_n258;
  assign new_n264 = n14 & n34;
  assign new_n265 = new_n256 ^ new_n252;
  assign new_n266 = ~new_n257 & new_n265;
  assign new_n267 = new_n266 ^ new_n252;
  assign new_n268 = n15 & n33;
  assign new_n269 = new_n268 ^ new_n267;
  assign new_n270 = new_n269 ^ new_n264;
  assign new_n271 = new_n270 ^ new_n263;
  assign new_n272 = n13 & n35;
  assign new_n273 = new_n272 ^ new_n263;
  assign new_n274 = ~new_n271 & new_n273;
  assign new_n275 = new_n274 ^ new_n272;
  assign new_n276 = n13 & n34;
  assign new_n277 = new_n268 ^ new_n264;
  assign new_n278 = ~new_n269 & new_n277;
  assign new_n279 = new_n278 ^ new_n264;
  assign new_n280 = n14 & n33;
  assign new_n281 = new_n280 ^ new_n279;
  assign new_n282 = new_n281 ^ new_n276;
  assign new_n283 = new_n282 ^ new_n275;
  assign new_n284 = n12 & n35;
  assign new_n285 = new_n284 ^ new_n282;
  assign new_n286 = ~new_n283 & new_n285;
  assign new_n287 = new_n286 ^ new_n284;
  assign new_n288 = n12 & n34;
  assign new_n289 = new_n280 ^ new_n276;
  assign new_n290 = ~new_n281 & new_n289;
  assign new_n291 = new_n290 ^ new_n276;
  assign new_n292 = n13 & n33;
  assign new_n293 = new_n292 ^ new_n291;
  assign new_n294 = new_n293 ^ new_n288;
  assign new_n295 = new_n294 ^ new_n287;
  assign new_n296 = n11 & n35;
  assign new_n297 = new_n296 ^ new_n294;
  assign new_n298 = ~new_n295 & new_n297;
  assign new_n299 = new_n298 ^ new_n296;
  assign new_n300 = n11 & n34;
  assign new_n301 = new_n292 ^ new_n288;
  assign new_n302 = ~new_n293 & new_n301;
  assign new_n303 = new_n302 ^ new_n288;
  assign new_n304 = n12 & n33;
  assign new_n305 = new_n304 ^ new_n303;
  assign new_n306 = new_n305 ^ new_n300;
  assign new_n307 = new_n306 ^ new_n299;
  assign new_n308 = n10 & n35;
  assign new_n309 = new_n308 ^ new_n306;
  assign new_n310 = ~new_n307 & new_n309;
  assign new_n311 = new_n310 ^ new_n308;
  assign new_n312 = n10 & n34;
  assign new_n313 = new_n304 ^ new_n300;
  assign new_n314 = ~new_n305 & new_n313;
  assign new_n315 = new_n314 ^ new_n300;
  assign new_n316 = n11 & n33;
  assign new_n317 = new_n316 ^ new_n315;
  assign new_n318 = new_n317 ^ new_n312;
  assign new_n319 = new_n318 ^ new_n311;
  assign new_n320 = n9 & n35;
  assign new_n321 = new_n320 ^ new_n318;
  assign new_n322 = ~new_n319 & new_n321;
  assign new_n323 = new_n322 ^ new_n320;
  assign new_n324 = n9 & n34;
  assign new_n325 = new_n316 ^ new_n312;
  assign new_n326 = ~new_n317 & new_n325;
  assign new_n327 = new_n326 ^ new_n312;
  assign new_n328 = n10 & n33;
  assign new_n329 = new_n328 ^ new_n327;
  assign new_n330 = new_n329 ^ new_n324;
  assign new_n331 = new_n330 ^ new_n323;
  assign new_n332 = n8 & n35;
  assign new_n333 = new_n332 ^ new_n330;
  assign new_n334 = ~new_n331 & new_n333;
  assign new_n335 = new_n334 ^ new_n332;
  assign new_n336 = n8 & n34;
  assign new_n337 = new_n328 ^ new_n324;
  assign new_n338 = ~new_n329 & new_n337;
  assign new_n339 = new_n338 ^ new_n324;
  assign new_n340 = n9 & n33;
  assign new_n341 = new_n340 ^ new_n339;
  assign new_n342 = new_n341 ^ new_n336;
  assign new_n343 = new_n342 ^ new_n335;
  assign new_n344 = n7 & n35;
  assign new_n345 = new_n344 ^ new_n342;
  assign new_n346 = ~new_n343 & new_n345;
  assign new_n347 = new_n346 ^ new_n344;
  assign new_n348 = n7 & n34;
  assign new_n349 = new_n340 ^ new_n336;
  assign new_n350 = ~new_n341 & new_n349;
  assign new_n351 = new_n350 ^ new_n336;
  assign new_n352 = n8 & n33;
  assign new_n353 = new_n352 ^ new_n351;
  assign new_n354 = new_n353 ^ new_n348;
  assign new_n355 = new_n354 ^ new_n347;
  assign new_n356 = n6 & n35;
  assign new_n357 = new_n356 ^ new_n354;
  assign new_n358 = ~new_n355 & new_n357;
  assign new_n359 = new_n358 ^ new_n356;
  assign new_n360 = n6 & n34;
  assign new_n361 = new_n352 ^ new_n348;
  assign new_n362 = ~new_n353 & new_n361;
  assign new_n363 = new_n362 ^ new_n348;
  assign new_n364 = n7 & n33;
  assign new_n365 = new_n364 ^ new_n363;
  assign new_n366 = new_n365 ^ new_n360;
  assign new_n367 = new_n366 ^ new_n359;
  assign new_n368 = n5 & n35;
  assign new_n369 = new_n368 ^ new_n366;
  assign new_n370 = ~new_n367 & new_n369;
  assign new_n371 = new_n370 ^ new_n368;
  assign new_n372 = n5 & n34;
  assign new_n373 = new_n364 ^ new_n360;
  assign new_n374 = ~new_n365 & new_n373;
  assign new_n375 = new_n374 ^ new_n360;
  assign new_n376 = n6 & n33;
  assign new_n377 = new_n376 ^ new_n375;
  assign new_n378 = new_n377 ^ new_n372;
  assign new_n379 = new_n378 ^ new_n371;
  assign new_n380 = n4 & n35;
  assign new_n381 = new_n380 ^ new_n378;
  assign new_n382 = ~new_n379 & new_n381;
  assign new_n383 = new_n382 ^ new_n380;
  assign new_n384 = n4 & n34;
  assign new_n385 = new_n376 ^ new_n372;
  assign new_n386 = ~new_n377 & new_n385;
  assign new_n387 = new_n386 ^ new_n372;
  assign new_n388 = n5 & n33;
  assign new_n389 = new_n388 ^ new_n387;
  assign new_n390 = new_n389 ^ new_n384;
  assign new_n391 = new_n390 ^ new_n383;
  assign new_n392 = n3 & n35;
  assign new_n393 = new_n392 ^ new_n390;
  assign new_n394 = ~new_n391 & new_n393;
  assign new_n395 = new_n394 ^ new_n392;
  assign new_n396 = n3 & n34;
  assign new_n397 = new_n388 ^ new_n384;
  assign new_n398 = ~new_n389 & new_n397;
  assign new_n399 = new_n398 ^ new_n384;
  assign new_n400 = n4 & n33;
  assign new_n401 = new_n400 ^ new_n399;
  assign new_n402 = new_n401 ^ new_n396;
  assign new_n403 = new_n402 ^ new_n395;
  assign new_n404 = n2 & n35;
  assign new_n405 = new_n404 ^ new_n402;
  assign new_n406 = ~new_n403 & new_n405;
  assign new_n407 = new_n406 ^ new_n404;
  assign new_n408 = n2 & n34;
  assign new_n409 = new_n400 ^ new_n396;
  assign new_n410 = ~new_n401 & new_n409;
  assign new_n411 = new_n410 ^ new_n396;
  assign new_n412 = n3 & n33;
  assign new_n413 = new_n412 ^ new_n411;
  assign new_n414 = new_n413 ^ new_n408;
  assign new_n415 = new_n414 ^ new_n407;
  assign new_n416 = n1 & n35;
  assign new_n417 = new_n416 ^ new_n414;
  assign new_n418 = ~new_n415 & new_n417;
  assign new_n419 = new_n418 ^ new_n416;
  assign new_n420 = n1 & n34;
  assign new_n421 = new_n412 ^ new_n408;
  assign new_n422 = ~new_n413 & new_n421;
  assign new_n423 = new_n422 ^ new_n408;
  assign new_n424 = n2 & n33;
  assign new_n425 = new_n424 ^ new_n423;
  assign new_n426 = new_n425 ^ new_n420;
  assign new_n427 = new_n419 & new_n426;
  assign new_n428 = n1 & n33;
  assign new_n429 = new_n424 ^ new_n420;
  assign new_n430 = ~new_n425 & new_n429;
  assign new_n431 = new_n430 ^ new_n420;
  assign new_n432 = new_n431 ^ new_n428;
  assign new_n433 = new_n432 ^ new_n427;
  assign new_n434 = new_n426 ^ new_n419;
  assign new_n435 = new_n416 ^ new_n415;
  assign new_n436 = new_n66 ^ new_n65;
  assign new_n437 = n32 & n35;
  assign new_n438 = n31 & n36;
  assign new_n439 = new_n437 & new_n438;
  assign new_n440 = new_n439 ^ new_n436;
  assign new_n441 = n30 & n36;
  assign new_n442 = new_n441 ^ new_n439;
  assign new_n443 = ~new_n440 & new_n442;
  assign new_n444 = new_n443 ^ new_n441;
  assign new_n445 = new_n72 ^ new_n71;
  assign new_n446 = new_n445 ^ new_n444;
  assign new_n447 = n29 & n36;
  assign new_n448 = new_n447 ^ new_n444;
  assign new_n449 = ~new_n446 & new_n448;
  assign new_n450 = new_n449 ^ new_n447;
  assign new_n451 = new_n81 ^ new_n80;
  assign new_n452 = new_n451 ^ new_n450;
  assign new_n453 = n28 & n36;
  assign new_n454 = new_n453 ^ new_n450;
  assign new_n455 = ~new_n452 & new_n454;
  assign new_n456 = new_n455 ^ new_n453;
  assign new_n457 = new_n92 ^ new_n91;
  assign new_n458 = new_n457 ^ new_n456;
  assign new_n459 = n27 & n36;
  assign new_n460 = new_n459 ^ new_n456;
  assign new_n461 = ~new_n458 & new_n460;
  assign new_n462 = new_n461 ^ new_n459;
  assign new_n463 = new_n104 ^ new_n103;
  assign new_n464 = new_n463 ^ new_n462;
  assign new_n465 = n26 & n36;
  assign new_n466 = new_n465 ^ new_n462;
  assign new_n467 = ~new_n464 & new_n466;
  assign new_n468 = new_n467 ^ new_n465;
  assign new_n469 = new_n116 ^ new_n115;
  assign new_n470 = new_n469 ^ new_n468;
  assign new_n471 = n25 & n36;
  assign new_n472 = new_n471 ^ new_n468;
  assign new_n473 = ~new_n470 & new_n472;
  assign new_n474 = new_n473 ^ new_n471;
  assign new_n475 = new_n128 ^ new_n127;
  assign new_n476 = new_n475 ^ new_n474;
  assign new_n477 = n24 & n36;
  assign new_n478 = new_n477 ^ new_n474;
  assign new_n479 = ~new_n476 & new_n478;
  assign new_n480 = new_n479 ^ new_n477;
  assign new_n481 = new_n140 ^ new_n139;
  assign new_n482 = new_n481 ^ new_n480;
  assign new_n483 = n23 & n36;
  assign new_n484 = new_n483 ^ new_n480;
  assign new_n485 = ~new_n482 & new_n484;
  assign new_n486 = new_n485 ^ new_n483;
  assign new_n487 = new_n152 ^ new_n151;
  assign new_n488 = new_n487 ^ new_n486;
  assign new_n489 = n22 & n36;
  assign new_n490 = new_n489 ^ new_n486;
  assign new_n491 = ~new_n488 & new_n490;
  assign new_n492 = new_n491 ^ new_n489;
  assign new_n493 = new_n164 ^ new_n163;
  assign new_n494 = new_n493 ^ new_n492;
  assign new_n495 = n21 & n36;
  assign new_n496 = new_n495 ^ new_n492;
  assign new_n497 = ~new_n494 & new_n496;
  assign new_n498 = new_n497 ^ new_n495;
  assign new_n499 = new_n176 ^ new_n175;
  assign new_n500 = new_n499 ^ new_n498;
  assign new_n501 = n20 & n36;
  assign new_n502 = new_n501 ^ new_n498;
  assign new_n503 = ~new_n500 & new_n502;
  assign new_n504 = new_n503 ^ new_n501;
  assign new_n505 = new_n188 ^ new_n187;
  assign new_n506 = new_n505 ^ new_n504;
  assign new_n507 = n19 & n36;
  assign new_n508 = new_n507 ^ new_n504;
  assign new_n509 = ~new_n506 & new_n508;
  assign new_n510 = new_n509 ^ new_n507;
  assign new_n511 = new_n200 ^ new_n199;
  assign new_n512 = new_n511 ^ new_n510;
  assign new_n513 = n18 & n36;
  assign new_n514 = new_n513 ^ new_n510;
  assign new_n515 = ~new_n512 & new_n514;
  assign new_n516 = new_n515 ^ new_n513;
  assign new_n517 = new_n212 ^ new_n211;
  assign new_n518 = new_n517 ^ new_n516;
  assign new_n519 = n17 & n36;
  assign new_n520 = new_n519 ^ new_n516;
  assign new_n521 = ~new_n518 & new_n520;
  assign new_n522 = new_n521 ^ new_n519;
  assign new_n523 = new_n224 ^ new_n223;
  assign new_n524 = new_n523 ^ new_n522;
  assign new_n525 = n16 & n36;
  assign new_n526 = new_n525 ^ new_n522;
  assign new_n527 = ~new_n524 & new_n526;
  assign new_n528 = new_n527 ^ new_n525;
  assign new_n529 = new_n236 ^ new_n235;
  assign new_n530 = new_n529 ^ new_n528;
  assign new_n531 = n15 & n36;
  assign new_n532 = new_n531 ^ new_n528;
  assign new_n533 = ~new_n530 & new_n532;
  assign new_n534 = new_n533 ^ new_n531;
  assign new_n535 = new_n248 ^ new_n247;
  assign new_n536 = new_n535 ^ new_n534;
  assign new_n537 = n14 & n36;
  assign new_n538 = new_n537 ^ new_n534;
  assign new_n539 = ~new_n536 & new_n538;
  assign new_n540 = new_n539 ^ new_n537;
  assign new_n541 = new_n260 ^ new_n259;
  assign new_n542 = new_n541 ^ new_n540;
  assign new_n543 = n13 & n36;
  assign new_n544 = new_n543 ^ new_n540;
  assign new_n545 = ~new_n542 & new_n544;
  assign new_n546 = new_n545 ^ new_n543;
  assign new_n547 = new_n272 ^ new_n271;
  assign new_n548 = new_n547 ^ new_n546;
  assign new_n549 = n12 & n36;
  assign new_n550 = new_n549 ^ new_n546;
  assign new_n551 = ~new_n548 & new_n550;
  assign new_n552 = new_n551 ^ new_n549;
  assign new_n553 = new_n284 ^ new_n283;
  assign new_n554 = new_n553 ^ new_n552;
  assign new_n555 = n11 & n36;
  assign new_n556 = new_n555 ^ new_n553;
  assign new_n557 = ~new_n554 & new_n556;
  assign new_n558 = new_n557 ^ new_n555;
  assign new_n559 = new_n296 ^ new_n295;
  assign new_n560 = new_n559 ^ new_n558;
  assign new_n561 = n10 & n36;
  assign new_n562 = new_n561 ^ new_n559;
  assign new_n563 = ~new_n560 & new_n562;
  assign new_n564 = new_n563 ^ new_n561;
  assign new_n565 = new_n308 ^ new_n307;
  assign new_n566 = new_n565 ^ new_n564;
  assign new_n567 = n9 & n36;
  assign new_n568 = new_n567 ^ new_n565;
  assign new_n569 = ~new_n566 & new_n568;
  assign new_n570 = new_n569 ^ new_n567;
  assign new_n571 = new_n320 ^ new_n319;
  assign new_n572 = new_n571 ^ new_n570;
  assign new_n573 = n8 & n36;
  assign new_n574 = new_n573 ^ new_n571;
  assign new_n575 = ~new_n572 & new_n574;
  assign new_n576 = new_n575 ^ new_n573;
  assign new_n577 = new_n332 ^ new_n331;
  assign new_n578 = new_n577 ^ new_n576;
  assign new_n579 = n7 & n36;
  assign new_n580 = new_n579 ^ new_n577;
  assign new_n581 = ~new_n578 & new_n580;
  assign new_n582 = new_n581 ^ new_n579;
  assign new_n583 = new_n344 ^ new_n343;
  assign new_n584 = new_n583 ^ new_n582;
  assign new_n585 = n6 & n36;
  assign new_n586 = new_n585 ^ new_n583;
  assign new_n587 = ~new_n584 & new_n586;
  assign new_n588 = new_n587 ^ new_n585;
  assign new_n589 = new_n356 ^ new_n355;
  assign new_n590 = new_n589 ^ new_n588;
  assign new_n591 = n5 & n36;
  assign new_n592 = new_n591 ^ new_n589;
  assign new_n593 = ~new_n590 & new_n592;
  assign new_n594 = new_n593 ^ new_n591;
  assign new_n595 = new_n368 ^ new_n367;
  assign new_n596 = new_n595 ^ new_n594;
  assign new_n597 = n4 & n36;
  assign new_n598 = new_n597 ^ new_n595;
  assign new_n599 = ~new_n596 & new_n598;
  assign new_n600 = new_n599 ^ new_n597;
  assign new_n601 = new_n380 ^ new_n379;
  assign new_n602 = new_n601 ^ new_n600;
  assign new_n603 = n3 & n36;
  assign new_n604 = new_n603 ^ new_n601;
  assign new_n605 = ~new_n602 & new_n604;
  assign new_n606 = new_n605 ^ new_n603;
  assign new_n607 = new_n392 ^ new_n391;
  assign new_n608 = new_n607 ^ new_n606;
  assign new_n609 = n2 & n36;
  assign new_n610 = new_n609 ^ new_n607;
  assign new_n611 = ~new_n608 & new_n610;
  assign new_n612 = new_n611 ^ new_n609;
  assign new_n613 = new_n404 ^ new_n403;
  assign new_n614 = new_n613 ^ new_n612;
  assign new_n615 = n1 & n36;
  assign new_n616 = new_n615 ^ new_n613;
  assign new_n617 = ~new_n614 & new_n616;
  assign new_n618 = new_n617 ^ new_n615;
  assign new_n619 = new_n435 & new_n618;
  assign new_n620 = new_n619 ^ new_n434;
  assign new_n621 = new_n618 ^ new_n435;
  assign new_n622 = new_n615 ^ new_n614;
  assign new_n623 = new_n438 ^ new_n437;
  assign new_n624 = n32 & n36;
  assign new_n625 = n31 & n37;
  assign new_n626 = new_n624 & new_n625;
  assign new_n627 = new_n626 ^ new_n623;
  assign new_n628 = n30 & n37;
  assign new_n629 = new_n628 ^ new_n626;
  assign new_n630 = ~new_n627 & new_n629;
  assign new_n631 = new_n630 ^ new_n628;
  assign new_n632 = new_n441 ^ new_n440;
  assign new_n633 = new_n632 ^ new_n631;
  assign new_n634 = n29 & n37;
  assign new_n635 = new_n634 ^ new_n631;
  assign new_n636 = ~new_n633 & new_n635;
  assign new_n637 = new_n636 ^ new_n634;
  assign new_n638 = new_n447 ^ new_n446;
  assign new_n639 = new_n638 ^ new_n637;
  assign new_n640 = n28 & n37;
  assign new_n641 = new_n640 ^ new_n637;
  assign new_n642 = ~new_n639 & new_n641;
  assign new_n643 = new_n642 ^ new_n640;
  assign new_n644 = new_n453 ^ new_n452;
  assign new_n645 = new_n644 ^ new_n643;
  assign new_n646 = n27 & n37;
  assign new_n647 = new_n646 ^ new_n643;
  assign new_n648 = ~new_n645 & new_n647;
  assign new_n649 = new_n648 ^ new_n646;
  assign new_n650 = new_n459 ^ new_n458;
  assign new_n651 = new_n650 ^ new_n649;
  assign new_n652 = n26 & n37;
  assign new_n653 = new_n652 ^ new_n649;
  assign new_n654 = ~new_n651 & new_n653;
  assign new_n655 = new_n654 ^ new_n652;
  assign new_n656 = new_n465 ^ new_n464;
  assign new_n657 = new_n656 ^ new_n655;
  assign new_n658 = n25 & n37;
  assign new_n659 = new_n658 ^ new_n655;
  assign new_n660 = ~new_n657 & new_n659;
  assign new_n661 = new_n660 ^ new_n658;
  assign new_n662 = new_n471 ^ new_n470;
  assign new_n663 = new_n662 ^ new_n661;
  assign new_n664 = n24 & n37;
  assign new_n665 = new_n664 ^ new_n661;
  assign new_n666 = ~new_n663 & new_n665;
  assign new_n667 = new_n666 ^ new_n664;
  assign new_n668 = new_n477 ^ new_n476;
  assign new_n669 = new_n668 ^ new_n667;
  assign new_n670 = n23 & n37;
  assign new_n671 = new_n670 ^ new_n667;
  assign new_n672 = ~new_n669 & new_n671;
  assign new_n673 = new_n672 ^ new_n670;
  assign new_n674 = new_n483 ^ new_n482;
  assign new_n675 = new_n674 ^ new_n673;
  assign new_n676 = n22 & n37;
  assign new_n677 = new_n676 ^ new_n673;
  assign new_n678 = ~new_n675 & new_n677;
  assign new_n679 = new_n678 ^ new_n676;
  assign new_n680 = new_n489 ^ new_n488;
  assign new_n681 = new_n680 ^ new_n679;
  assign new_n682 = n21 & n37;
  assign new_n683 = new_n682 ^ new_n679;
  assign new_n684 = ~new_n681 & new_n683;
  assign new_n685 = new_n684 ^ new_n682;
  assign new_n686 = new_n495 ^ new_n494;
  assign new_n687 = new_n686 ^ new_n685;
  assign new_n688 = n20 & n37;
  assign new_n689 = new_n688 ^ new_n685;
  assign new_n690 = ~new_n687 & new_n689;
  assign new_n691 = new_n690 ^ new_n688;
  assign new_n692 = new_n501 ^ new_n500;
  assign new_n693 = new_n692 ^ new_n691;
  assign new_n694 = n19 & n37;
  assign new_n695 = new_n694 ^ new_n691;
  assign new_n696 = ~new_n693 & new_n695;
  assign new_n697 = new_n696 ^ new_n694;
  assign new_n698 = new_n507 ^ new_n506;
  assign new_n699 = new_n698 ^ new_n697;
  assign new_n700 = n18 & n37;
  assign new_n701 = new_n700 ^ new_n697;
  assign new_n702 = ~new_n699 & new_n701;
  assign new_n703 = new_n702 ^ new_n700;
  assign new_n704 = new_n513 ^ new_n512;
  assign new_n705 = new_n704 ^ new_n703;
  assign new_n706 = n17 & n37;
  assign new_n707 = new_n706 ^ new_n703;
  assign new_n708 = ~new_n705 & new_n707;
  assign new_n709 = new_n708 ^ new_n706;
  assign new_n710 = new_n519 ^ new_n518;
  assign new_n711 = new_n710 ^ new_n709;
  assign new_n712 = n16 & n37;
  assign new_n713 = new_n712 ^ new_n709;
  assign new_n714 = ~new_n711 & new_n713;
  assign new_n715 = new_n714 ^ new_n712;
  assign new_n716 = new_n525 ^ new_n524;
  assign new_n717 = new_n716 ^ new_n715;
  assign new_n718 = n15 & n37;
  assign new_n719 = new_n718 ^ new_n715;
  assign new_n720 = ~new_n717 & new_n719;
  assign new_n721 = new_n720 ^ new_n718;
  assign new_n722 = new_n531 ^ new_n530;
  assign new_n723 = new_n722 ^ new_n721;
  assign new_n724 = n14 & n37;
  assign new_n725 = new_n724 ^ new_n721;
  assign new_n726 = ~new_n723 & new_n725;
  assign new_n727 = new_n726 ^ new_n724;
  assign new_n728 = new_n537 ^ new_n536;
  assign new_n729 = new_n728 ^ new_n727;
  assign new_n730 = n13 & n37;
  assign new_n731 = new_n730 ^ new_n727;
  assign new_n732 = ~new_n729 & new_n731;
  assign new_n733 = new_n732 ^ new_n730;
  assign new_n734 = new_n543 ^ new_n542;
  assign new_n735 = new_n734 ^ new_n733;
  assign new_n736 = n12 & n37;
  assign new_n737 = new_n736 ^ new_n733;
  assign new_n738 = ~new_n735 & new_n737;
  assign new_n739 = new_n738 ^ new_n736;
  assign new_n740 = new_n549 ^ new_n548;
  assign new_n741 = new_n740 ^ new_n739;
  assign new_n742 = n11 & n37;
  assign new_n743 = new_n742 ^ new_n739;
  assign new_n744 = ~new_n741 & new_n743;
  assign new_n745 = new_n744 ^ new_n742;
  assign new_n746 = new_n555 ^ new_n554;
  assign new_n747 = new_n746 ^ new_n745;
  assign new_n748 = n10 & n37;
  assign new_n749 = new_n748 ^ new_n746;
  assign new_n750 = ~new_n747 & new_n749;
  assign new_n751 = new_n750 ^ new_n748;
  assign new_n752 = new_n561 ^ new_n560;
  assign new_n753 = new_n752 ^ new_n751;
  assign new_n754 = n9 & n37;
  assign new_n755 = new_n754 ^ new_n752;
  assign new_n756 = ~new_n753 & new_n755;
  assign new_n757 = new_n756 ^ new_n754;
  assign new_n758 = new_n567 ^ new_n566;
  assign new_n759 = new_n758 ^ new_n757;
  assign new_n760 = n8 & n37;
  assign new_n761 = new_n760 ^ new_n758;
  assign new_n762 = ~new_n759 & new_n761;
  assign new_n763 = new_n762 ^ new_n760;
  assign new_n764 = new_n573 ^ new_n572;
  assign new_n765 = new_n764 ^ new_n763;
  assign new_n766 = n7 & n37;
  assign new_n767 = new_n766 ^ new_n764;
  assign new_n768 = ~new_n765 & new_n767;
  assign new_n769 = new_n768 ^ new_n766;
  assign new_n770 = new_n579 ^ new_n578;
  assign new_n771 = new_n770 ^ new_n769;
  assign new_n772 = n6 & n37;
  assign new_n773 = new_n772 ^ new_n770;
  assign new_n774 = ~new_n771 & new_n773;
  assign new_n775 = new_n774 ^ new_n772;
  assign new_n776 = new_n585 ^ new_n584;
  assign new_n777 = new_n776 ^ new_n775;
  assign new_n778 = n5 & n37;
  assign new_n779 = new_n778 ^ new_n776;
  assign new_n780 = ~new_n777 & new_n779;
  assign new_n781 = new_n780 ^ new_n778;
  assign new_n782 = new_n591 ^ new_n590;
  assign new_n783 = new_n782 ^ new_n781;
  assign new_n784 = n4 & n37;
  assign new_n785 = new_n784 ^ new_n782;
  assign new_n786 = ~new_n783 & new_n785;
  assign new_n787 = new_n786 ^ new_n784;
  assign new_n788 = new_n597 ^ new_n596;
  assign new_n789 = new_n788 ^ new_n787;
  assign new_n790 = n3 & n37;
  assign new_n791 = new_n790 ^ new_n788;
  assign new_n792 = ~new_n789 & new_n791;
  assign new_n793 = new_n792 ^ new_n790;
  assign new_n794 = new_n603 ^ new_n602;
  assign new_n795 = new_n794 ^ new_n793;
  assign new_n796 = n2 & n37;
  assign new_n797 = new_n796 ^ new_n794;
  assign new_n798 = ~new_n795 & new_n797;
  assign new_n799 = new_n798 ^ new_n796;
  assign new_n800 = new_n609 ^ new_n608;
  assign new_n801 = new_n800 ^ new_n799;
  assign new_n802 = n1 & n37;
  assign new_n803 = new_n802 ^ new_n800;
  assign new_n804 = ~new_n801 & new_n803;
  assign new_n805 = new_n804 ^ new_n802;
  assign new_n806 = new_n622 & new_n805;
  assign new_n807 = new_n806 ^ new_n621;
  assign new_n808 = new_n805 ^ new_n622;
  assign new_n809 = new_n802 ^ new_n801;
  assign new_n810 = new_n625 ^ new_n624;
  assign new_n811 = n32 & n37;
  assign new_n812 = n31 & n38;
  assign new_n813 = new_n811 & new_n812;
  assign new_n814 = new_n813 ^ new_n810;
  assign new_n815 = n30 & n38;
  assign new_n816 = new_n815 ^ new_n813;
  assign new_n817 = ~new_n814 & new_n816;
  assign new_n818 = new_n817 ^ new_n815;
  assign new_n819 = new_n628 ^ new_n627;
  assign new_n820 = new_n819 ^ new_n818;
  assign new_n821 = n29 & n38;
  assign new_n822 = new_n821 ^ new_n818;
  assign new_n823 = ~new_n820 & new_n822;
  assign new_n824 = new_n823 ^ new_n821;
  assign new_n825 = new_n634 ^ new_n633;
  assign new_n826 = new_n825 ^ new_n824;
  assign new_n827 = n28 & n38;
  assign new_n828 = new_n827 ^ new_n824;
  assign new_n829 = ~new_n826 & new_n828;
  assign new_n830 = new_n829 ^ new_n827;
  assign new_n831 = new_n640 ^ new_n639;
  assign new_n832 = new_n831 ^ new_n830;
  assign new_n833 = n27 & n38;
  assign new_n834 = new_n833 ^ new_n830;
  assign new_n835 = ~new_n832 & new_n834;
  assign new_n836 = new_n835 ^ new_n833;
  assign new_n837 = new_n646 ^ new_n645;
  assign new_n838 = new_n837 ^ new_n836;
  assign new_n839 = n26 & n38;
  assign new_n840 = new_n839 ^ new_n836;
  assign new_n841 = ~new_n838 & new_n840;
  assign new_n842 = new_n841 ^ new_n839;
  assign new_n843 = new_n652 ^ new_n651;
  assign new_n844 = new_n843 ^ new_n842;
  assign new_n845 = n25 & n38;
  assign new_n846 = new_n845 ^ new_n842;
  assign new_n847 = ~new_n844 & new_n846;
  assign new_n848 = new_n847 ^ new_n845;
  assign new_n849 = new_n658 ^ new_n657;
  assign new_n850 = new_n849 ^ new_n848;
  assign new_n851 = n24 & n38;
  assign new_n852 = new_n851 ^ new_n848;
  assign new_n853 = ~new_n850 & new_n852;
  assign new_n854 = new_n853 ^ new_n851;
  assign new_n855 = new_n664 ^ new_n663;
  assign new_n856 = new_n855 ^ new_n854;
  assign new_n857 = n23 & n38;
  assign new_n858 = new_n857 ^ new_n854;
  assign new_n859 = ~new_n856 & new_n858;
  assign new_n860 = new_n859 ^ new_n857;
  assign new_n861 = new_n670 ^ new_n669;
  assign new_n862 = new_n861 ^ new_n860;
  assign new_n863 = n22 & n38;
  assign new_n864 = new_n863 ^ new_n860;
  assign new_n865 = ~new_n862 & new_n864;
  assign new_n866 = new_n865 ^ new_n863;
  assign new_n867 = new_n676 ^ new_n675;
  assign new_n868 = new_n867 ^ new_n866;
  assign new_n869 = n21 & n38;
  assign new_n870 = new_n869 ^ new_n866;
  assign new_n871 = ~new_n868 & new_n870;
  assign new_n872 = new_n871 ^ new_n869;
  assign new_n873 = new_n682 ^ new_n681;
  assign new_n874 = new_n873 ^ new_n872;
  assign new_n875 = n20 & n38;
  assign new_n876 = new_n875 ^ new_n872;
  assign new_n877 = ~new_n874 & new_n876;
  assign new_n878 = new_n877 ^ new_n875;
  assign new_n879 = new_n688 ^ new_n687;
  assign new_n880 = new_n879 ^ new_n878;
  assign new_n881 = n19 & n38;
  assign new_n882 = new_n881 ^ new_n878;
  assign new_n883 = ~new_n880 & new_n882;
  assign new_n884 = new_n883 ^ new_n881;
  assign new_n885 = new_n694 ^ new_n693;
  assign new_n886 = new_n885 ^ new_n884;
  assign new_n887 = n18 & n38;
  assign new_n888 = new_n887 ^ new_n884;
  assign new_n889 = ~new_n886 & new_n888;
  assign new_n890 = new_n889 ^ new_n887;
  assign new_n891 = new_n700 ^ new_n699;
  assign new_n892 = new_n891 ^ new_n890;
  assign new_n893 = n17 & n38;
  assign new_n894 = new_n893 ^ new_n890;
  assign new_n895 = ~new_n892 & new_n894;
  assign new_n896 = new_n895 ^ new_n893;
  assign new_n897 = new_n706 ^ new_n705;
  assign new_n898 = new_n897 ^ new_n896;
  assign new_n899 = n16 & n38;
  assign new_n900 = new_n899 ^ new_n896;
  assign new_n901 = ~new_n898 & new_n900;
  assign new_n902 = new_n901 ^ new_n899;
  assign new_n903 = new_n712 ^ new_n711;
  assign new_n904 = new_n903 ^ new_n902;
  assign new_n905 = n15 & n38;
  assign new_n906 = new_n905 ^ new_n902;
  assign new_n907 = ~new_n904 & new_n906;
  assign new_n908 = new_n907 ^ new_n905;
  assign new_n909 = new_n718 ^ new_n717;
  assign new_n910 = new_n909 ^ new_n908;
  assign new_n911 = n14 & n38;
  assign new_n912 = new_n911 ^ new_n908;
  assign new_n913 = ~new_n910 & new_n912;
  assign new_n914 = new_n913 ^ new_n911;
  assign new_n915 = new_n724 ^ new_n723;
  assign new_n916 = new_n915 ^ new_n914;
  assign new_n917 = n13 & n38;
  assign new_n918 = new_n917 ^ new_n914;
  assign new_n919 = ~new_n916 & new_n918;
  assign new_n920 = new_n919 ^ new_n917;
  assign new_n921 = new_n730 ^ new_n729;
  assign new_n922 = new_n921 ^ new_n920;
  assign new_n923 = n12 & n38;
  assign new_n924 = new_n923 ^ new_n920;
  assign new_n925 = ~new_n922 & new_n924;
  assign new_n926 = new_n925 ^ new_n923;
  assign new_n927 = new_n736 ^ new_n735;
  assign new_n928 = new_n927 ^ new_n926;
  assign new_n929 = n11 & n38;
  assign new_n930 = new_n929 ^ new_n926;
  assign new_n931 = ~new_n928 & new_n930;
  assign new_n932 = new_n931 ^ new_n929;
  assign new_n933 = new_n742 ^ new_n741;
  assign new_n934 = new_n933 ^ new_n932;
  assign new_n935 = n10 & n38;
  assign new_n936 = new_n935 ^ new_n932;
  assign new_n937 = ~new_n934 & new_n936;
  assign new_n938 = new_n937 ^ new_n935;
  assign new_n939 = new_n748 ^ new_n747;
  assign new_n940 = new_n939 ^ new_n938;
  assign new_n941 = n9 & n38;
  assign new_n942 = new_n941 ^ new_n939;
  assign new_n943 = ~new_n940 & new_n942;
  assign new_n944 = new_n943 ^ new_n941;
  assign new_n945 = new_n754 ^ new_n753;
  assign new_n946 = new_n945 ^ new_n944;
  assign new_n947 = n8 & n38;
  assign new_n948 = new_n947 ^ new_n945;
  assign new_n949 = ~new_n946 & new_n948;
  assign new_n950 = new_n949 ^ new_n947;
  assign new_n951 = new_n760 ^ new_n759;
  assign new_n952 = new_n951 ^ new_n950;
  assign new_n953 = n7 & n38;
  assign new_n954 = new_n953 ^ new_n951;
  assign new_n955 = ~new_n952 & new_n954;
  assign new_n956 = new_n955 ^ new_n953;
  assign new_n957 = new_n766 ^ new_n765;
  assign new_n958 = new_n957 ^ new_n956;
  assign new_n959 = n6 & n38;
  assign new_n960 = new_n959 ^ new_n957;
  assign new_n961 = ~new_n958 & new_n960;
  assign new_n962 = new_n961 ^ new_n959;
  assign new_n963 = new_n772 ^ new_n771;
  assign new_n964 = new_n963 ^ new_n962;
  assign new_n965 = n5 & n38;
  assign new_n966 = new_n965 ^ new_n963;
  assign new_n967 = ~new_n964 & new_n966;
  assign new_n968 = new_n967 ^ new_n965;
  assign new_n969 = new_n778 ^ new_n777;
  assign new_n970 = new_n969 ^ new_n968;
  assign new_n971 = n4 & n38;
  assign new_n972 = new_n971 ^ new_n969;
  assign new_n973 = ~new_n970 & new_n972;
  assign new_n974 = new_n973 ^ new_n971;
  assign new_n975 = new_n784 ^ new_n783;
  assign new_n976 = new_n975 ^ new_n974;
  assign new_n977 = n3 & n38;
  assign new_n978 = new_n977 ^ new_n975;
  assign new_n979 = ~new_n976 & new_n978;
  assign new_n980 = new_n979 ^ new_n977;
  assign new_n981 = new_n790 ^ new_n789;
  assign new_n982 = new_n981 ^ new_n980;
  assign new_n983 = n2 & n38;
  assign new_n984 = new_n983 ^ new_n981;
  assign new_n985 = ~new_n982 & new_n984;
  assign new_n986 = new_n985 ^ new_n983;
  assign new_n987 = new_n796 ^ new_n795;
  assign new_n988 = new_n987 ^ new_n986;
  assign new_n989 = n1 & n38;
  assign new_n990 = new_n989 ^ new_n987;
  assign new_n991 = ~new_n988 & new_n990;
  assign new_n992 = new_n991 ^ new_n989;
  assign new_n993 = new_n809 & new_n992;
  assign new_n994 = new_n993 ^ new_n808;
  assign new_n995 = new_n992 ^ new_n809;
  assign new_n996 = new_n989 ^ new_n988;
  assign new_n997 = new_n812 ^ new_n811;
  assign new_n998 = n32 & n38;
  assign new_n999 = n31 & n39;
  assign new_n1000 = new_n998 & new_n999;
  assign new_n1001 = new_n1000 ^ new_n997;
  assign new_n1002 = n30 & n39;
  assign new_n1003 = new_n1002 ^ new_n1000;
  assign new_n1004 = ~new_n1001 & new_n1003;
  assign new_n1005 = new_n1004 ^ new_n1002;
  assign new_n1006 = new_n815 ^ new_n814;
  assign new_n1007 = new_n1006 ^ new_n1005;
  assign new_n1008 = n29 & n39;
  assign new_n1009 = new_n1008 ^ new_n1005;
  assign new_n1010 = ~new_n1007 & new_n1009;
  assign new_n1011 = new_n1010 ^ new_n1008;
  assign new_n1012 = new_n821 ^ new_n820;
  assign new_n1013 = new_n1012 ^ new_n1011;
  assign new_n1014 = n28 & n39;
  assign new_n1015 = new_n1014 ^ new_n1011;
  assign new_n1016 = ~new_n1013 & new_n1015;
  assign new_n1017 = new_n1016 ^ new_n1014;
  assign new_n1018 = new_n827 ^ new_n826;
  assign new_n1019 = new_n1018 ^ new_n1017;
  assign new_n1020 = n27 & n39;
  assign new_n1021 = new_n1020 ^ new_n1017;
  assign new_n1022 = ~new_n1019 & new_n1021;
  assign new_n1023 = new_n1022 ^ new_n1020;
  assign new_n1024 = new_n833 ^ new_n832;
  assign new_n1025 = new_n1024 ^ new_n1023;
  assign new_n1026 = n26 & n39;
  assign new_n1027 = new_n1026 ^ new_n1023;
  assign new_n1028 = ~new_n1025 & new_n1027;
  assign new_n1029 = new_n1028 ^ new_n1026;
  assign new_n1030 = new_n839 ^ new_n838;
  assign new_n1031 = new_n1030 ^ new_n1029;
  assign new_n1032 = n25 & n39;
  assign new_n1033 = new_n1032 ^ new_n1029;
  assign new_n1034 = ~new_n1031 & new_n1033;
  assign new_n1035 = new_n1034 ^ new_n1032;
  assign new_n1036 = new_n845 ^ new_n844;
  assign new_n1037 = new_n1036 ^ new_n1035;
  assign new_n1038 = n24 & n39;
  assign new_n1039 = new_n1038 ^ new_n1035;
  assign new_n1040 = ~new_n1037 & new_n1039;
  assign new_n1041 = new_n1040 ^ new_n1038;
  assign new_n1042 = new_n851 ^ new_n850;
  assign new_n1043 = new_n1042 ^ new_n1041;
  assign new_n1044 = n23 & n39;
  assign new_n1045 = new_n1044 ^ new_n1041;
  assign new_n1046 = ~new_n1043 & new_n1045;
  assign new_n1047 = new_n1046 ^ new_n1044;
  assign new_n1048 = new_n857 ^ new_n856;
  assign new_n1049 = new_n1048 ^ new_n1047;
  assign new_n1050 = n22 & n39;
  assign new_n1051 = new_n1050 ^ new_n1047;
  assign new_n1052 = ~new_n1049 & new_n1051;
  assign new_n1053 = new_n1052 ^ new_n1050;
  assign new_n1054 = new_n863 ^ new_n862;
  assign new_n1055 = new_n1054 ^ new_n1053;
  assign new_n1056 = n21 & n39;
  assign new_n1057 = new_n1056 ^ new_n1053;
  assign new_n1058 = ~new_n1055 & new_n1057;
  assign new_n1059 = new_n1058 ^ new_n1056;
  assign new_n1060 = new_n869 ^ new_n868;
  assign new_n1061 = new_n1060 ^ new_n1059;
  assign new_n1062 = n20 & n39;
  assign new_n1063 = new_n1062 ^ new_n1059;
  assign new_n1064 = ~new_n1061 & new_n1063;
  assign new_n1065 = new_n1064 ^ new_n1062;
  assign new_n1066 = new_n875 ^ new_n874;
  assign new_n1067 = new_n1066 ^ new_n1065;
  assign new_n1068 = n19 & n39;
  assign new_n1069 = new_n1068 ^ new_n1065;
  assign new_n1070 = ~new_n1067 & new_n1069;
  assign new_n1071 = new_n1070 ^ new_n1068;
  assign new_n1072 = new_n881 ^ new_n880;
  assign new_n1073 = new_n1072 ^ new_n1071;
  assign new_n1074 = n18 & n39;
  assign new_n1075 = new_n1074 ^ new_n1071;
  assign new_n1076 = ~new_n1073 & new_n1075;
  assign new_n1077 = new_n1076 ^ new_n1074;
  assign new_n1078 = new_n887 ^ new_n886;
  assign new_n1079 = new_n1078 ^ new_n1077;
  assign new_n1080 = n17 & n39;
  assign new_n1081 = new_n1080 ^ new_n1077;
  assign new_n1082 = ~new_n1079 & new_n1081;
  assign new_n1083 = new_n1082 ^ new_n1080;
  assign new_n1084 = new_n893 ^ new_n892;
  assign new_n1085 = new_n1084 ^ new_n1083;
  assign new_n1086 = n16 & n39;
  assign new_n1087 = new_n1086 ^ new_n1083;
  assign new_n1088 = ~new_n1085 & new_n1087;
  assign new_n1089 = new_n1088 ^ new_n1086;
  assign new_n1090 = new_n899 ^ new_n898;
  assign new_n1091 = new_n1090 ^ new_n1089;
  assign new_n1092 = n15 & n39;
  assign new_n1093 = new_n1092 ^ new_n1089;
  assign new_n1094 = ~new_n1091 & new_n1093;
  assign new_n1095 = new_n1094 ^ new_n1092;
  assign new_n1096 = new_n905 ^ new_n904;
  assign new_n1097 = new_n1096 ^ new_n1095;
  assign new_n1098 = n14 & n39;
  assign new_n1099 = new_n1098 ^ new_n1095;
  assign new_n1100 = ~new_n1097 & new_n1099;
  assign new_n1101 = new_n1100 ^ new_n1098;
  assign new_n1102 = new_n911 ^ new_n910;
  assign new_n1103 = new_n1102 ^ new_n1101;
  assign new_n1104 = n13 & n39;
  assign new_n1105 = new_n1104 ^ new_n1101;
  assign new_n1106 = ~new_n1103 & new_n1105;
  assign new_n1107 = new_n1106 ^ new_n1104;
  assign new_n1108 = new_n917 ^ new_n916;
  assign new_n1109 = new_n1108 ^ new_n1107;
  assign new_n1110 = n12 & n39;
  assign new_n1111 = new_n1110 ^ new_n1107;
  assign new_n1112 = ~new_n1109 & new_n1111;
  assign new_n1113 = new_n1112 ^ new_n1110;
  assign new_n1114 = new_n923 ^ new_n922;
  assign new_n1115 = new_n1114 ^ new_n1113;
  assign new_n1116 = n11 & n39;
  assign new_n1117 = new_n1116 ^ new_n1113;
  assign new_n1118 = ~new_n1115 & new_n1117;
  assign new_n1119 = new_n1118 ^ new_n1116;
  assign new_n1120 = new_n929 ^ new_n928;
  assign new_n1121 = new_n1120 ^ new_n1119;
  assign new_n1122 = n10 & n39;
  assign new_n1123 = new_n1122 ^ new_n1119;
  assign new_n1124 = ~new_n1121 & new_n1123;
  assign new_n1125 = new_n1124 ^ new_n1122;
  assign new_n1126 = new_n935 ^ new_n934;
  assign new_n1127 = new_n1126 ^ new_n1125;
  assign new_n1128 = n9 & n39;
  assign new_n1129 = new_n1128 ^ new_n1125;
  assign new_n1130 = ~new_n1127 & new_n1129;
  assign new_n1131 = new_n1130 ^ new_n1128;
  assign new_n1132 = new_n941 ^ new_n940;
  assign new_n1133 = new_n1132 ^ new_n1131;
  assign new_n1134 = n8 & n39;
  assign new_n1135 = new_n1134 ^ new_n1132;
  assign new_n1136 = ~new_n1133 & new_n1135;
  assign new_n1137 = new_n1136 ^ new_n1134;
  assign new_n1138 = new_n947 ^ new_n946;
  assign new_n1139 = new_n1138 ^ new_n1137;
  assign new_n1140 = n7 & n39;
  assign new_n1141 = new_n1140 ^ new_n1138;
  assign new_n1142 = ~new_n1139 & new_n1141;
  assign new_n1143 = new_n1142 ^ new_n1140;
  assign new_n1144 = new_n953 ^ new_n952;
  assign new_n1145 = new_n1144 ^ new_n1143;
  assign new_n1146 = n6 & n39;
  assign new_n1147 = new_n1146 ^ new_n1144;
  assign new_n1148 = ~new_n1145 & new_n1147;
  assign new_n1149 = new_n1148 ^ new_n1146;
  assign new_n1150 = new_n959 ^ new_n958;
  assign new_n1151 = new_n1150 ^ new_n1149;
  assign new_n1152 = n5 & n39;
  assign new_n1153 = new_n1152 ^ new_n1150;
  assign new_n1154 = ~new_n1151 & new_n1153;
  assign new_n1155 = new_n1154 ^ new_n1152;
  assign new_n1156 = new_n965 ^ new_n964;
  assign new_n1157 = new_n1156 ^ new_n1155;
  assign new_n1158 = n4 & n39;
  assign new_n1159 = new_n1158 ^ new_n1156;
  assign new_n1160 = ~new_n1157 & new_n1159;
  assign new_n1161 = new_n1160 ^ new_n1158;
  assign new_n1162 = new_n971 ^ new_n970;
  assign new_n1163 = new_n1162 ^ new_n1161;
  assign new_n1164 = n3 & n39;
  assign new_n1165 = new_n1164 ^ new_n1162;
  assign new_n1166 = ~new_n1163 & new_n1165;
  assign new_n1167 = new_n1166 ^ new_n1164;
  assign new_n1168 = new_n977 ^ new_n976;
  assign new_n1169 = new_n1168 ^ new_n1167;
  assign new_n1170 = n2 & n39;
  assign new_n1171 = new_n1170 ^ new_n1168;
  assign new_n1172 = ~new_n1169 & new_n1171;
  assign new_n1173 = new_n1172 ^ new_n1170;
  assign new_n1174 = new_n983 ^ new_n982;
  assign new_n1175 = new_n1174 ^ new_n1173;
  assign new_n1176 = n1 & n39;
  assign new_n1177 = new_n1176 ^ new_n1174;
  assign new_n1178 = ~new_n1175 & new_n1177;
  assign new_n1179 = new_n1178 ^ new_n1176;
  assign new_n1180 = new_n996 & new_n1179;
  assign new_n1181 = new_n1180 ^ new_n995;
  assign new_n1182 = new_n1179 ^ new_n996;
  assign new_n1183 = new_n1176 ^ new_n1175;
  assign new_n1184 = new_n999 ^ new_n998;
  assign new_n1185 = n32 & n39;
  assign new_n1186 = n31 & n40;
  assign new_n1187 = new_n1185 & new_n1186;
  assign new_n1188 = new_n1187 ^ new_n1184;
  assign new_n1189 = n30 & n40;
  assign new_n1190 = new_n1189 ^ new_n1187;
  assign new_n1191 = ~new_n1188 & new_n1190;
  assign new_n1192 = new_n1191 ^ new_n1189;
  assign new_n1193 = new_n1002 ^ new_n1001;
  assign new_n1194 = new_n1193 ^ new_n1192;
  assign new_n1195 = n29 & n40;
  assign new_n1196 = new_n1195 ^ new_n1192;
  assign new_n1197 = ~new_n1194 & new_n1196;
  assign new_n1198 = new_n1197 ^ new_n1195;
  assign new_n1199 = new_n1008 ^ new_n1007;
  assign new_n1200 = new_n1199 ^ new_n1198;
  assign new_n1201 = n28 & n40;
  assign new_n1202 = new_n1201 ^ new_n1198;
  assign new_n1203 = ~new_n1200 & new_n1202;
  assign new_n1204 = new_n1203 ^ new_n1201;
  assign new_n1205 = new_n1014 ^ new_n1013;
  assign new_n1206 = new_n1205 ^ new_n1204;
  assign new_n1207 = n27 & n40;
  assign new_n1208 = new_n1207 ^ new_n1204;
  assign new_n1209 = ~new_n1206 & new_n1208;
  assign new_n1210 = new_n1209 ^ new_n1207;
  assign new_n1211 = new_n1020 ^ new_n1019;
  assign new_n1212 = new_n1211 ^ new_n1210;
  assign new_n1213 = n26 & n40;
  assign new_n1214 = new_n1213 ^ new_n1210;
  assign new_n1215 = ~new_n1212 & new_n1214;
  assign new_n1216 = new_n1215 ^ new_n1213;
  assign new_n1217 = new_n1026 ^ new_n1025;
  assign new_n1218 = new_n1217 ^ new_n1216;
  assign new_n1219 = n25 & n40;
  assign new_n1220 = new_n1219 ^ new_n1216;
  assign new_n1221 = ~new_n1218 & new_n1220;
  assign new_n1222 = new_n1221 ^ new_n1219;
  assign new_n1223 = new_n1032 ^ new_n1031;
  assign new_n1224 = new_n1223 ^ new_n1222;
  assign new_n1225 = n24 & n40;
  assign new_n1226 = new_n1225 ^ new_n1222;
  assign new_n1227 = ~new_n1224 & new_n1226;
  assign new_n1228 = new_n1227 ^ new_n1225;
  assign new_n1229 = new_n1038 ^ new_n1037;
  assign new_n1230 = new_n1229 ^ new_n1228;
  assign new_n1231 = n23 & n40;
  assign new_n1232 = new_n1231 ^ new_n1228;
  assign new_n1233 = ~new_n1230 & new_n1232;
  assign new_n1234 = new_n1233 ^ new_n1231;
  assign new_n1235 = new_n1044 ^ new_n1043;
  assign new_n1236 = new_n1235 ^ new_n1234;
  assign new_n1237 = n22 & n40;
  assign new_n1238 = new_n1237 ^ new_n1234;
  assign new_n1239 = ~new_n1236 & new_n1238;
  assign new_n1240 = new_n1239 ^ new_n1237;
  assign new_n1241 = new_n1050 ^ new_n1049;
  assign new_n1242 = new_n1241 ^ new_n1240;
  assign new_n1243 = n21 & n40;
  assign new_n1244 = new_n1243 ^ new_n1240;
  assign new_n1245 = ~new_n1242 & new_n1244;
  assign new_n1246 = new_n1245 ^ new_n1243;
  assign new_n1247 = new_n1056 ^ new_n1055;
  assign new_n1248 = new_n1247 ^ new_n1246;
  assign new_n1249 = n20 & n40;
  assign new_n1250 = new_n1249 ^ new_n1246;
  assign new_n1251 = ~new_n1248 & new_n1250;
  assign new_n1252 = new_n1251 ^ new_n1249;
  assign new_n1253 = new_n1062 ^ new_n1061;
  assign new_n1254 = new_n1253 ^ new_n1252;
  assign new_n1255 = n19 & n40;
  assign new_n1256 = new_n1255 ^ new_n1252;
  assign new_n1257 = ~new_n1254 & new_n1256;
  assign new_n1258 = new_n1257 ^ new_n1255;
  assign new_n1259 = new_n1068 ^ new_n1067;
  assign new_n1260 = new_n1259 ^ new_n1258;
  assign new_n1261 = n18 & n40;
  assign new_n1262 = new_n1261 ^ new_n1258;
  assign new_n1263 = ~new_n1260 & new_n1262;
  assign new_n1264 = new_n1263 ^ new_n1261;
  assign new_n1265 = new_n1074 ^ new_n1073;
  assign new_n1266 = new_n1265 ^ new_n1264;
  assign new_n1267 = n17 & n40;
  assign new_n1268 = new_n1267 ^ new_n1264;
  assign new_n1269 = ~new_n1266 & new_n1268;
  assign new_n1270 = new_n1269 ^ new_n1267;
  assign new_n1271 = new_n1080 ^ new_n1079;
  assign new_n1272 = new_n1271 ^ new_n1270;
  assign new_n1273 = n16 & n40;
  assign new_n1274 = new_n1273 ^ new_n1270;
  assign new_n1275 = ~new_n1272 & new_n1274;
  assign new_n1276 = new_n1275 ^ new_n1273;
  assign new_n1277 = new_n1086 ^ new_n1085;
  assign new_n1278 = new_n1277 ^ new_n1276;
  assign new_n1279 = n15 & n40;
  assign new_n1280 = new_n1279 ^ new_n1276;
  assign new_n1281 = ~new_n1278 & new_n1280;
  assign new_n1282 = new_n1281 ^ new_n1279;
  assign new_n1283 = new_n1092 ^ new_n1091;
  assign new_n1284 = new_n1283 ^ new_n1282;
  assign new_n1285 = n14 & n40;
  assign new_n1286 = new_n1285 ^ new_n1282;
  assign new_n1287 = ~new_n1284 & new_n1286;
  assign new_n1288 = new_n1287 ^ new_n1285;
  assign new_n1289 = new_n1098 ^ new_n1097;
  assign new_n1290 = new_n1289 ^ new_n1288;
  assign new_n1291 = n13 & n40;
  assign new_n1292 = new_n1291 ^ new_n1288;
  assign new_n1293 = ~new_n1290 & new_n1292;
  assign new_n1294 = new_n1293 ^ new_n1291;
  assign new_n1295 = new_n1104 ^ new_n1103;
  assign new_n1296 = new_n1295 ^ new_n1294;
  assign new_n1297 = n12 & n40;
  assign new_n1298 = new_n1297 ^ new_n1294;
  assign new_n1299 = ~new_n1296 & new_n1298;
  assign new_n1300 = new_n1299 ^ new_n1297;
  assign new_n1301 = new_n1110 ^ new_n1109;
  assign new_n1302 = new_n1301 ^ new_n1300;
  assign new_n1303 = n11 & n40;
  assign new_n1304 = new_n1303 ^ new_n1300;
  assign new_n1305 = ~new_n1302 & new_n1304;
  assign new_n1306 = new_n1305 ^ new_n1303;
  assign new_n1307 = new_n1116 ^ new_n1115;
  assign new_n1308 = new_n1307 ^ new_n1306;
  assign new_n1309 = n10 & n40;
  assign new_n1310 = new_n1309 ^ new_n1306;
  assign new_n1311 = ~new_n1308 & new_n1310;
  assign new_n1312 = new_n1311 ^ new_n1309;
  assign new_n1313 = new_n1122 ^ new_n1121;
  assign new_n1314 = new_n1313 ^ new_n1312;
  assign new_n1315 = n9 & n40;
  assign new_n1316 = new_n1315 ^ new_n1312;
  assign new_n1317 = ~new_n1314 & new_n1316;
  assign new_n1318 = new_n1317 ^ new_n1315;
  assign new_n1319 = new_n1128 ^ new_n1127;
  assign new_n1320 = new_n1319 ^ new_n1318;
  assign new_n1321 = n8 & n40;
  assign new_n1322 = new_n1321 ^ new_n1318;
  assign new_n1323 = ~new_n1320 & new_n1322;
  assign new_n1324 = new_n1323 ^ new_n1321;
  assign new_n1325 = new_n1134 ^ new_n1133;
  assign new_n1326 = new_n1325 ^ new_n1324;
  assign new_n1327 = n7 & n40;
  assign new_n1328 = new_n1327 ^ new_n1325;
  assign new_n1329 = ~new_n1326 & new_n1328;
  assign new_n1330 = new_n1329 ^ new_n1327;
  assign new_n1331 = new_n1140 ^ new_n1139;
  assign new_n1332 = new_n1331 ^ new_n1330;
  assign new_n1333 = n6 & n40;
  assign new_n1334 = new_n1333 ^ new_n1331;
  assign new_n1335 = ~new_n1332 & new_n1334;
  assign new_n1336 = new_n1335 ^ new_n1333;
  assign new_n1337 = new_n1146 ^ new_n1145;
  assign new_n1338 = new_n1337 ^ new_n1336;
  assign new_n1339 = n5 & n40;
  assign new_n1340 = new_n1339 ^ new_n1337;
  assign new_n1341 = ~new_n1338 & new_n1340;
  assign new_n1342 = new_n1341 ^ new_n1339;
  assign new_n1343 = new_n1152 ^ new_n1151;
  assign new_n1344 = new_n1343 ^ new_n1342;
  assign new_n1345 = n4 & n40;
  assign new_n1346 = new_n1345 ^ new_n1343;
  assign new_n1347 = ~new_n1344 & new_n1346;
  assign new_n1348 = new_n1347 ^ new_n1345;
  assign new_n1349 = new_n1158 ^ new_n1157;
  assign new_n1350 = new_n1349 ^ new_n1348;
  assign new_n1351 = n3 & n40;
  assign new_n1352 = new_n1351 ^ new_n1349;
  assign new_n1353 = ~new_n1350 & new_n1352;
  assign new_n1354 = new_n1353 ^ new_n1351;
  assign new_n1355 = new_n1164 ^ new_n1163;
  assign new_n1356 = new_n1355 ^ new_n1354;
  assign new_n1357 = n2 & n40;
  assign new_n1358 = new_n1357 ^ new_n1355;
  assign new_n1359 = ~new_n1356 & new_n1358;
  assign new_n1360 = new_n1359 ^ new_n1357;
  assign new_n1361 = new_n1170 ^ new_n1169;
  assign new_n1362 = new_n1361 ^ new_n1360;
  assign new_n1363 = n1 & n40;
  assign new_n1364 = new_n1363 ^ new_n1361;
  assign new_n1365 = ~new_n1362 & new_n1364;
  assign new_n1366 = new_n1365 ^ new_n1363;
  assign new_n1367 = new_n1183 & new_n1366;
  assign new_n1368 = new_n1367 ^ new_n1182;
  assign new_n1369 = new_n1366 ^ new_n1183;
  assign new_n1370 = new_n1363 ^ new_n1362;
  assign new_n1371 = new_n1186 ^ new_n1185;
  assign new_n1372 = n32 & n40;
  assign new_n1373 = n31 & n41;
  assign new_n1374 = new_n1372 & new_n1373;
  assign new_n1375 = new_n1374 ^ new_n1371;
  assign new_n1376 = n30 & n41;
  assign new_n1377 = new_n1376 ^ new_n1374;
  assign new_n1378 = ~new_n1375 & new_n1377;
  assign new_n1379 = new_n1378 ^ new_n1376;
  assign new_n1380 = new_n1189 ^ new_n1188;
  assign new_n1381 = new_n1380 ^ new_n1379;
  assign new_n1382 = n29 & n41;
  assign new_n1383 = new_n1382 ^ new_n1379;
  assign new_n1384 = ~new_n1381 & new_n1383;
  assign new_n1385 = new_n1384 ^ new_n1382;
  assign new_n1386 = new_n1195 ^ new_n1194;
  assign new_n1387 = new_n1386 ^ new_n1385;
  assign new_n1388 = n28 & n41;
  assign new_n1389 = new_n1388 ^ new_n1385;
  assign new_n1390 = ~new_n1387 & new_n1389;
  assign new_n1391 = new_n1390 ^ new_n1388;
  assign new_n1392 = new_n1201 ^ new_n1200;
  assign new_n1393 = new_n1392 ^ new_n1391;
  assign new_n1394 = n27 & n41;
  assign new_n1395 = new_n1394 ^ new_n1391;
  assign new_n1396 = ~new_n1393 & new_n1395;
  assign new_n1397 = new_n1396 ^ new_n1394;
  assign new_n1398 = new_n1207 ^ new_n1206;
  assign new_n1399 = new_n1398 ^ new_n1397;
  assign new_n1400 = n26 & n41;
  assign new_n1401 = new_n1400 ^ new_n1397;
  assign new_n1402 = ~new_n1399 & new_n1401;
  assign new_n1403 = new_n1402 ^ new_n1400;
  assign new_n1404 = new_n1213 ^ new_n1212;
  assign new_n1405 = new_n1404 ^ new_n1403;
  assign new_n1406 = n25 & n41;
  assign new_n1407 = new_n1406 ^ new_n1403;
  assign new_n1408 = ~new_n1405 & new_n1407;
  assign new_n1409 = new_n1408 ^ new_n1406;
  assign new_n1410 = new_n1219 ^ new_n1218;
  assign new_n1411 = new_n1410 ^ new_n1409;
  assign new_n1412 = n24 & n41;
  assign new_n1413 = new_n1412 ^ new_n1409;
  assign new_n1414 = ~new_n1411 & new_n1413;
  assign new_n1415 = new_n1414 ^ new_n1412;
  assign new_n1416 = new_n1225 ^ new_n1224;
  assign new_n1417 = new_n1416 ^ new_n1415;
  assign new_n1418 = n23 & n41;
  assign new_n1419 = new_n1418 ^ new_n1415;
  assign new_n1420 = ~new_n1417 & new_n1419;
  assign new_n1421 = new_n1420 ^ new_n1418;
  assign new_n1422 = new_n1231 ^ new_n1230;
  assign new_n1423 = new_n1422 ^ new_n1421;
  assign new_n1424 = n22 & n41;
  assign new_n1425 = new_n1424 ^ new_n1421;
  assign new_n1426 = ~new_n1423 & new_n1425;
  assign new_n1427 = new_n1426 ^ new_n1424;
  assign new_n1428 = new_n1237 ^ new_n1236;
  assign new_n1429 = new_n1428 ^ new_n1427;
  assign new_n1430 = n21 & n41;
  assign new_n1431 = new_n1430 ^ new_n1427;
  assign new_n1432 = ~new_n1429 & new_n1431;
  assign new_n1433 = new_n1432 ^ new_n1430;
  assign new_n1434 = new_n1243 ^ new_n1242;
  assign new_n1435 = new_n1434 ^ new_n1433;
  assign new_n1436 = n20 & n41;
  assign new_n1437 = new_n1436 ^ new_n1433;
  assign new_n1438 = ~new_n1435 & new_n1437;
  assign new_n1439 = new_n1438 ^ new_n1436;
  assign new_n1440 = new_n1249 ^ new_n1248;
  assign new_n1441 = new_n1440 ^ new_n1439;
  assign new_n1442 = n19 & n41;
  assign new_n1443 = new_n1442 ^ new_n1439;
  assign new_n1444 = ~new_n1441 & new_n1443;
  assign new_n1445 = new_n1444 ^ new_n1442;
  assign new_n1446 = new_n1255 ^ new_n1254;
  assign new_n1447 = new_n1446 ^ new_n1445;
  assign new_n1448 = n18 & n41;
  assign new_n1449 = new_n1448 ^ new_n1445;
  assign new_n1450 = ~new_n1447 & new_n1449;
  assign new_n1451 = new_n1450 ^ new_n1448;
  assign new_n1452 = new_n1261 ^ new_n1260;
  assign new_n1453 = new_n1452 ^ new_n1451;
  assign new_n1454 = n17 & n41;
  assign new_n1455 = new_n1454 ^ new_n1451;
  assign new_n1456 = ~new_n1453 & new_n1455;
  assign new_n1457 = new_n1456 ^ new_n1454;
  assign new_n1458 = new_n1267 ^ new_n1266;
  assign new_n1459 = new_n1458 ^ new_n1457;
  assign new_n1460 = n16 & n41;
  assign new_n1461 = new_n1460 ^ new_n1457;
  assign new_n1462 = ~new_n1459 & new_n1461;
  assign new_n1463 = new_n1462 ^ new_n1460;
  assign new_n1464 = new_n1273 ^ new_n1272;
  assign new_n1465 = new_n1464 ^ new_n1463;
  assign new_n1466 = n15 & n41;
  assign new_n1467 = new_n1466 ^ new_n1463;
  assign new_n1468 = ~new_n1465 & new_n1467;
  assign new_n1469 = new_n1468 ^ new_n1466;
  assign new_n1470 = new_n1279 ^ new_n1278;
  assign new_n1471 = new_n1470 ^ new_n1469;
  assign new_n1472 = n14 & n41;
  assign new_n1473 = new_n1472 ^ new_n1469;
  assign new_n1474 = ~new_n1471 & new_n1473;
  assign new_n1475 = new_n1474 ^ new_n1472;
  assign new_n1476 = new_n1285 ^ new_n1284;
  assign new_n1477 = new_n1476 ^ new_n1475;
  assign new_n1478 = n13 & n41;
  assign new_n1479 = new_n1478 ^ new_n1475;
  assign new_n1480 = ~new_n1477 & new_n1479;
  assign new_n1481 = new_n1480 ^ new_n1478;
  assign new_n1482 = new_n1291 ^ new_n1290;
  assign new_n1483 = new_n1482 ^ new_n1481;
  assign new_n1484 = n12 & n41;
  assign new_n1485 = new_n1484 ^ new_n1481;
  assign new_n1486 = ~new_n1483 & new_n1485;
  assign new_n1487 = new_n1486 ^ new_n1484;
  assign new_n1488 = new_n1297 ^ new_n1296;
  assign new_n1489 = new_n1488 ^ new_n1487;
  assign new_n1490 = n11 & n41;
  assign new_n1491 = new_n1490 ^ new_n1487;
  assign new_n1492 = ~new_n1489 & new_n1491;
  assign new_n1493 = new_n1492 ^ new_n1490;
  assign new_n1494 = new_n1303 ^ new_n1302;
  assign new_n1495 = new_n1494 ^ new_n1493;
  assign new_n1496 = n10 & n41;
  assign new_n1497 = new_n1496 ^ new_n1493;
  assign new_n1498 = ~new_n1495 & new_n1497;
  assign new_n1499 = new_n1498 ^ new_n1496;
  assign new_n1500 = new_n1309 ^ new_n1308;
  assign new_n1501 = new_n1500 ^ new_n1499;
  assign new_n1502 = n9 & n41;
  assign new_n1503 = new_n1502 ^ new_n1499;
  assign new_n1504 = ~new_n1501 & new_n1503;
  assign new_n1505 = new_n1504 ^ new_n1502;
  assign new_n1506 = new_n1315 ^ new_n1314;
  assign new_n1507 = new_n1506 ^ new_n1505;
  assign new_n1508 = n8 & n41;
  assign new_n1509 = new_n1508 ^ new_n1505;
  assign new_n1510 = ~new_n1507 & new_n1509;
  assign new_n1511 = new_n1510 ^ new_n1508;
  assign new_n1512 = new_n1321 ^ new_n1320;
  assign new_n1513 = new_n1512 ^ new_n1511;
  assign new_n1514 = n7 & n41;
  assign new_n1515 = new_n1514 ^ new_n1511;
  assign new_n1516 = ~new_n1513 & new_n1515;
  assign new_n1517 = new_n1516 ^ new_n1514;
  assign new_n1518 = new_n1327 ^ new_n1326;
  assign new_n1519 = new_n1518 ^ new_n1517;
  assign new_n1520 = n6 & n41;
  assign new_n1521 = new_n1520 ^ new_n1518;
  assign new_n1522 = ~new_n1519 & new_n1521;
  assign new_n1523 = new_n1522 ^ new_n1520;
  assign new_n1524 = new_n1333 ^ new_n1332;
  assign new_n1525 = new_n1524 ^ new_n1523;
  assign new_n1526 = n5 & n41;
  assign new_n1527 = new_n1526 ^ new_n1524;
  assign new_n1528 = ~new_n1525 & new_n1527;
  assign new_n1529 = new_n1528 ^ new_n1526;
  assign new_n1530 = new_n1339 ^ new_n1338;
  assign new_n1531 = new_n1530 ^ new_n1529;
  assign new_n1532 = n4 & n41;
  assign new_n1533 = new_n1532 ^ new_n1530;
  assign new_n1534 = ~new_n1531 & new_n1533;
  assign new_n1535 = new_n1534 ^ new_n1532;
  assign new_n1536 = new_n1345 ^ new_n1344;
  assign new_n1537 = new_n1536 ^ new_n1535;
  assign new_n1538 = n3 & n41;
  assign new_n1539 = new_n1538 ^ new_n1536;
  assign new_n1540 = ~new_n1537 & new_n1539;
  assign new_n1541 = new_n1540 ^ new_n1538;
  assign new_n1542 = new_n1351 ^ new_n1350;
  assign new_n1543 = new_n1542 ^ new_n1541;
  assign new_n1544 = n2 & n41;
  assign new_n1545 = new_n1544 ^ new_n1542;
  assign new_n1546 = ~new_n1543 & new_n1545;
  assign new_n1547 = new_n1546 ^ new_n1544;
  assign new_n1548 = new_n1357 ^ new_n1356;
  assign new_n1549 = new_n1548 ^ new_n1547;
  assign new_n1550 = n1 & n41;
  assign new_n1551 = new_n1550 ^ new_n1548;
  assign new_n1552 = ~new_n1549 & new_n1551;
  assign new_n1553 = new_n1552 ^ new_n1550;
  assign new_n1554 = new_n1370 & new_n1553;
  assign new_n1555 = new_n1554 ^ new_n1369;
  assign new_n1556 = new_n1553 ^ new_n1370;
  assign new_n1557 = new_n1550 ^ new_n1549;
  assign new_n1558 = new_n1373 ^ new_n1372;
  assign new_n1559 = n32 & n41;
  assign new_n1560 = n31 & n42;
  assign new_n1561 = new_n1559 & new_n1560;
  assign new_n1562 = new_n1561 ^ new_n1558;
  assign new_n1563 = n30 & n42;
  assign new_n1564 = new_n1563 ^ new_n1561;
  assign new_n1565 = ~new_n1562 & new_n1564;
  assign new_n1566 = new_n1565 ^ new_n1563;
  assign new_n1567 = new_n1376 ^ new_n1375;
  assign new_n1568 = new_n1567 ^ new_n1566;
  assign new_n1569 = n29 & n42;
  assign new_n1570 = new_n1569 ^ new_n1566;
  assign new_n1571 = ~new_n1568 & new_n1570;
  assign new_n1572 = new_n1571 ^ new_n1569;
  assign new_n1573 = new_n1382 ^ new_n1381;
  assign new_n1574 = new_n1573 ^ new_n1572;
  assign new_n1575 = n28 & n42;
  assign new_n1576 = new_n1575 ^ new_n1572;
  assign new_n1577 = ~new_n1574 & new_n1576;
  assign new_n1578 = new_n1577 ^ new_n1575;
  assign new_n1579 = new_n1388 ^ new_n1387;
  assign new_n1580 = new_n1579 ^ new_n1578;
  assign new_n1581 = n27 & n42;
  assign new_n1582 = new_n1581 ^ new_n1578;
  assign new_n1583 = ~new_n1580 & new_n1582;
  assign new_n1584 = new_n1583 ^ new_n1581;
  assign new_n1585 = new_n1394 ^ new_n1393;
  assign new_n1586 = new_n1585 ^ new_n1584;
  assign new_n1587 = n26 & n42;
  assign new_n1588 = new_n1587 ^ new_n1584;
  assign new_n1589 = ~new_n1586 & new_n1588;
  assign new_n1590 = new_n1589 ^ new_n1587;
  assign new_n1591 = new_n1400 ^ new_n1399;
  assign new_n1592 = new_n1591 ^ new_n1590;
  assign new_n1593 = n25 & n42;
  assign new_n1594 = new_n1593 ^ new_n1590;
  assign new_n1595 = ~new_n1592 & new_n1594;
  assign new_n1596 = new_n1595 ^ new_n1593;
  assign new_n1597 = new_n1406 ^ new_n1405;
  assign new_n1598 = new_n1597 ^ new_n1596;
  assign new_n1599 = n24 & n42;
  assign new_n1600 = new_n1599 ^ new_n1596;
  assign new_n1601 = ~new_n1598 & new_n1600;
  assign new_n1602 = new_n1601 ^ new_n1599;
  assign new_n1603 = new_n1412 ^ new_n1411;
  assign new_n1604 = new_n1603 ^ new_n1602;
  assign new_n1605 = n23 & n42;
  assign new_n1606 = new_n1605 ^ new_n1602;
  assign new_n1607 = ~new_n1604 & new_n1606;
  assign new_n1608 = new_n1607 ^ new_n1605;
  assign new_n1609 = new_n1418 ^ new_n1417;
  assign new_n1610 = new_n1609 ^ new_n1608;
  assign new_n1611 = n22 & n42;
  assign new_n1612 = new_n1611 ^ new_n1608;
  assign new_n1613 = ~new_n1610 & new_n1612;
  assign new_n1614 = new_n1613 ^ new_n1611;
  assign new_n1615 = new_n1424 ^ new_n1423;
  assign new_n1616 = new_n1615 ^ new_n1614;
  assign new_n1617 = n21 & n42;
  assign new_n1618 = new_n1617 ^ new_n1614;
  assign new_n1619 = ~new_n1616 & new_n1618;
  assign new_n1620 = new_n1619 ^ new_n1617;
  assign new_n1621 = new_n1430 ^ new_n1429;
  assign new_n1622 = new_n1621 ^ new_n1620;
  assign new_n1623 = n20 & n42;
  assign new_n1624 = new_n1623 ^ new_n1620;
  assign new_n1625 = ~new_n1622 & new_n1624;
  assign new_n1626 = new_n1625 ^ new_n1623;
  assign new_n1627 = new_n1436 ^ new_n1435;
  assign new_n1628 = new_n1627 ^ new_n1626;
  assign new_n1629 = n19 & n42;
  assign new_n1630 = new_n1629 ^ new_n1626;
  assign new_n1631 = ~new_n1628 & new_n1630;
  assign new_n1632 = new_n1631 ^ new_n1629;
  assign new_n1633 = new_n1442 ^ new_n1441;
  assign new_n1634 = new_n1633 ^ new_n1632;
  assign new_n1635 = n18 & n42;
  assign new_n1636 = new_n1635 ^ new_n1632;
  assign new_n1637 = ~new_n1634 & new_n1636;
  assign new_n1638 = new_n1637 ^ new_n1635;
  assign new_n1639 = new_n1448 ^ new_n1447;
  assign new_n1640 = new_n1639 ^ new_n1638;
  assign new_n1641 = n17 & n42;
  assign new_n1642 = new_n1641 ^ new_n1638;
  assign new_n1643 = ~new_n1640 & new_n1642;
  assign new_n1644 = new_n1643 ^ new_n1641;
  assign new_n1645 = new_n1454 ^ new_n1453;
  assign new_n1646 = new_n1645 ^ new_n1644;
  assign new_n1647 = n16 & n42;
  assign new_n1648 = new_n1647 ^ new_n1644;
  assign new_n1649 = ~new_n1646 & new_n1648;
  assign new_n1650 = new_n1649 ^ new_n1647;
  assign new_n1651 = new_n1460 ^ new_n1459;
  assign new_n1652 = new_n1651 ^ new_n1650;
  assign new_n1653 = n15 & n42;
  assign new_n1654 = new_n1653 ^ new_n1650;
  assign new_n1655 = ~new_n1652 & new_n1654;
  assign new_n1656 = new_n1655 ^ new_n1653;
  assign new_n1657 = new_n1466 ^ new_n1465;
  assign new_n1658 = new_n1657 ^ new_n1656;
  assign new_n1659 = n14 & n42;
  assign new_n1660 = new_n1659 ^ new_n1656;
  assign new_n1661 = ~new_n1658 & new_n1660;
  assign new_n1662 = new_n1661 ^ new_n1659;
  assign new_n1663 = new_n1472 ^ new_n1471;
  assign new_n1664 = new_n1663 ^ new_n1662;
  assign new_n1665 = n13 & n42;
  assign new_n1666 = new_n1665 ^ new_n1662;
  assign new_n1667 = ~new_n1664 & new_n1666;
  assign new_n1668 = new_n1667 ^ new_n1665;
  assign new_n1669 = new_n1478 ^ new_n1477;
  assign new_n1670 = new_n1669 ^ new_n1668;
  assign new_n1671 = n12 & n42;
  assign new_n1672 = new_n1671 ^ new_n1668;
  assign new_n1673 = ~new_n1670 & new_n1672;
  assign new_n1674 = new_n1673 ^ new_n1671;
  assign new_n1675 = new_n1484 ^ new_n1483;
  assign new_n1676 = new_n1675 ^ new_n1674;
  assign new_n1677 = n11 & n42;
  assign new_n1678 = new_n1677 ^ new_n1674;
  assign new_n1679 = ~new_n1676 & new_n1678;
  assign new_n1680 = new_n1679 ^ new_n1677;
  assign new_n1681 = new_n1490 ^ new_n1489;
  assign new_n1682 = new_n1681 ^ new_n1680;
  assign new_n1683 = n10 & n42;
  assign new_n1684 = new_n1683 ^ new_n1680;
  assign new_n1685 = ~new_n1682 & new_n1684;
  assign new_n1686 = new_n1685 ^ new_n1683;
  assign new_n1687 = new_n1496 ^ new_n1495;
  assign new_n1688 = new_n1687 ^ new_n1686;
  assign new_n1689 = n9 & n42;
  assign new_n1690 = new_n1689 ^ new_n1686;
  assign new_n1691 = ~new_n1688 & new_n1690;
  assign new_n1692 = new_n1691 ^ new_n1689;
  assign new_n1693 = new_n1502 ^ new_n1501;
  assign new_n1694 = new_n1693 ^ new_n1692;
  assign new_n1695 = n8 & n42;
  assign new_n1696 = new_n1695 ^ new_n1692;
  assign new_n1697 = ~new_n1694 & new_n1696;
  assign new_n1698 = new_n1697 ^ new_n1695;
  assign new_n1699 = new_n1508 ^ new_n1507;
  assign new_n1700 = new_n1699 ^ new_n1698;
  assign new_n1701 = n7 & n42;
  assign new_n1702 = new_n1701 ^ new_n1698;
  assign new_n1703 = ~new_n1700 & new_n1702;
  assign new_n1704 = new_n1703 ^ new_n1701;
  assign new_n1705 = new_n1514 ^ new_n1513;
  assign new_n1706 = new_n1705 ^ new_n1704;
  assign new_n1707 = n6 & n42;
  assign new_n1708 = new_n1707 ^ new_n1704;
  assign new_n1709 = ~new_n1706 & new_n1708;
  assign new_n1710 = new_n1709 ^ new_n1707;
  assign new_n1711 = new_n1520 ^ new_n1519;
  assign new_n1712 = new_n1711 ^ new_n1710;
  assign new_n1713 = n5 & n42;
  assign new_n1714 = new_n1713 ^ new_n1711;
  assign new_n1715 = ~new_n1712 & new_n1714;
  assign new_n1716 = new_n1715 ^ new_n1713;
  assign new_n1717 = new_n1526 ^ new_n1525;
  assign new_n1718 = new_n1717 ^ new_n1716;
  assign new_n1719 = n4 & n42;
  assign new_n1720 = new_n1719 ^ new_n1717;
  assign new_n1721 = ~new_n1718 & new_n1720;
  assign new_n1722 = new_n1721 ^ new_n1719;
  assign new_n1723 = new_n1532 ^ new_n1531;
  assign new_n1724 = new_n1723 ^ new_n1722;
  assign new_n1725 = n3 & n42;
  assign new_n1726 = new_n1725 ^ new_n1723;
  assign new_n1727 = ~new_n1724 & new_n1726;
  assign new_n1728 = new_n1727 ^ new_n1725;
  assign new_n1729 = new_n1538 ^ new_n1537;
  assign new_n1730 = new_n1729 ^ new_n1728;
  assign new_n1731 = n2 & n42;
  assign new_n1732 = new_n1731 ^ new_n1729;
  assign new_n1733 = ~new_n1730 & new_n1732;
  assign new_n1734 = new_n1733 ^ new_n1731;
  assign new_n1735 = new_n1544 ^ new_n1543;
  assign new_n1736 = new_n1735 ^ new_n1734;
  assign new_n1737 = n1 & n42;
  assign new_n1738 = new_n1737 ^ new_n1735;
  assign new_n1739 = ~new_n1736 & new_n1738;
  assign new_n1740 = new_n1739 ^ new_n1737;
  assign new_n1741 = new_n1557 & new_n1740;
  assign new_n1742 = new_n1741 ^ new_n1556;
  assign new_n1743 = new_n1740 ^ new_n1557;
  assign new_n1744 = new_n1737 ^ new_n1736;
  assign new_n1745 = new_n1560 ^ new_n1559;
  assign new_n1746 = n32 & n42;
  assign new_n1747 = n31 & n43;
  assign new_n1748 = new_n1746 & new_n1747;
  assign new_n1749 = new_n1748 ^ new_n1745;
  assign new_n1750 = n30 & n43;
  assign new_n1751 = new_n1750 ^ new_n1748;
  assign new_n1752 = ~new_n1749 & new_n1751;
  assign new_n1753 = new_n1752 ^ new_n1750;
  assign new_n1754 = new_n1563 ^ new_n1562;
  assign new_n1755 = new_n1754 ^ new_n1753;
  assign new_n1756 = n29 & n43;
  assign new_n1757 = new_n1756 ^ new_n1753;
  assign new_n1758 = ~new_n1755 & new_n1757;
  assign new_n1759 = new_n1758 ^ new_n1756;
  assign new_n1760 = new_n1569 ^ new_n1568;
  assign new_n1761 = new_n1760 ^ new_n1759;
  assign new_n1762 = n28 & n43;
  assign new_n1763 = new_n1762 ^ new_n1759;
  assign new_n1764 = ~new_n1761 & new_n1763;
  assign new_n1765 = new_n1764 ^ new_n1762;
  assign new_n1766 = new_n1575 ^ new_n1574;
  assign new_n1767 = new_n1766 ^ new_n1765;
  assign new_n1768 = n27 & n43;
  assign new_n1769 = new_n1768 ^ new_n1765;
  assign new_n1770 = ~new_n1767 & new_n1769;
  assign new_n1771 = new_n1770 ^ new_n1768;
  assign new_n1772 = new_n1581 ^ new_n1580;
  assign new_n1773 = new_n1772 ^ new_n1771;
  assign new_n1774 = n26 & n43;
  assign new_n1775 = new_n1774 ^ new_n1771;
  assign new_n1776 = ~new_n1773 & new_n1775;
  assign new_n1777 = new_n1776 ^ new_n1774;
  assign new_n1778 = new_n1587 ^ new_n1586;
  assign new_n1779 = new_n1778 ^ new_n1777;
  assign new_n1780 = n25 & n43;
  assign new_n1781 = new_n1780 ^ new_n1777;
  assign new_n1782 = ~new_n1779 & new_n1781;
  assign new_n1783 = new_n1782 ^ new_n1780;
  assign new_n1784 = new_n1593 ^ new_n1592;
  assign new_n1785 = new_n1784 ^ new_n1783;
  assign new_n1786 = n24 & n43;
  assign new_n1787 = new_n1786 ^ new_n1783;
  assign new_n1788 = ~new_n1785 & new_n1787;
  assign new_n1789 = new_n1788 ^ new_n1786;
  assign new_n1790 = new_n1599 ^ new_n1598;
  assign new_n1791 = new_n1790 ^ new_n1789;
  assign new_n1792 = n23 & n43;
  assign new_n1793 = new_n1792 ^ new_n1789;
  assign new_n1794 = ~new_n1791 & new_n1793;
  assign new_n1795 = new_n1794 ^ new_n1792;
  assign new_n1796 = new_n1605 ^ new_n1604;
  assign new_n1797 = new_n1796 ^ new_n1795;
  assign new_n1798 = n22 & n43;
  assign new_n1799 = new_n1798 ^ new_n1795;
  assign new_n1800 = ~new_n1797 & new_n1799;
  assign new_n1801 = new_n1800 ^ new_n1798;
  assign new_n1802 = new_n1611 ^ new_n1610;
  assign new_n1803 = new_n1802 ^ new_n1801;
  assign new_n1804 = n21 & n43;
  assign new_n1805 = new_n1804 ^ new_n1801;
  assign new_n1806 = ~new_n1803 & new_n1805;
  assign new_n1807 = new_n1806 ^ new_n1804;
  assign new_n1808 = new_n1617 ^ new_n1616;
  assign new_n1809 = new_n1808 ^ new_n1807;
  assign new_n1810 = n20 & n43;
  assign new_n1811 = new_n1810 ^ new_n1807;
  assign new_n1812 = ~new_n1809 & new_n1811;
  assign new_n1813 = new_n1812 ^ new_n1810;
  assign new_n1814 = new_n1623 ^ new_n1622;
  assign new_n1815 = new_n1814 ^ new_n1813;
  assign new_n1816 = n19 & n43;
  assign new_n1817 = new_n1816 ^ new_n1813;
  assign new_n1818 = ~new_n1815 & new_n1817;
  assign new_n1819 = new_n1818 ^ new_n1816;
  assign new_n1820 = new_n1629 ^ new_n1628;
  assign new_n1821 = new_n1820 ^ new_n1819;
  assign new_n1822 = n18 & n43;
  assign new_n1823 = new_n1822 ^ new_n1819;
  assign new_n1824 = ~new_n1821 & new_n1823;
  assign new_n1825 = new_n1824 ^ new_n1822;
  assign new_n1826 = new_n1635 ^ new_n1634;
  assign new_n1827 = new_n1826 ^ new_n1825;
  assign new_n1828 = n17 & n43;
  assign new_n1829 = new_n1828 ^ new_n1825;
  assign new_n1830 = ~new_n1827 & new_n1829;
  assign new_n1831 = new_n1830 ^ new_n1828;
  assign new_n1832 = new_n1641 ^ new_n1640;
  assign new_n1833 = new_n1832 ^ new_n1831;
  assign new_n1834 = n16 & n43;
  assign new_n1835 = new_n1834 ^ new_n1831;
  assign new_n1836 = ~new_n1833 & new_n1835;
  assign new_n1837 = new_n1836 ^ new_n1834;
  assign new_n1838 = new_n1647 ^ new_n1646;
  assign new_n1839 = new_n1838 ^ new_n1837;
  assign new_n1840 = n15 & n43;
  assign new_n1841 = new_n1840 ^ new_n1837;
  assign new_n1842 = ~new_n1839 & new_n1841;
  assign new_n1843 = new_n1842 ^ new_n1840;
  assign new_n1844 = new_n1653 ^ new_n1652;
  assign new_n1845 = new_n1844 ^ new_n1843;
  assign new_n1846 = n14 & n43;
  assign new_n1847 = new_n1846 ^ new_n1843;
  assign new_n1848 = ~new_n1845 & new_n1847;
  assign new_n1849 = new_n1848 ^ new_n1846;
  assign new_n1850 = new_n1659 ^ new_n1658;
  assign new_n1851 = new_n1850 ^ new_n1849;
  assign new_n1852 = n13 & n43;
  assign new_n1853 = new_n1852 ^ new_n1849;
  assign new_n1854 = ~new_n1851 & new_n1853;
  assign new_n1855 = new_n1854 ^ new_n1852;
  assign new_n1856 = new_n1665 ^ new_n1664;
  assign new_n1857 = new_n1856 ^ new_n1855;
  assign new_n1858 = n12 & n43;
  assign new_n1859 = new_n1858 ^ new_n1855;
  assign new_n1860 = ~new_n1857 & new_n1859;
  assign new_n1861 = new_n1860 ^ new_n1858;
  assign new_n1862 = new_n1671 ^ new_n1670;
  assign new_n1863 = new_n1862 ^ new_n1861;
  assign new_n1864 = n11 & n43;
  assign new_n1865 = new_n1864 ^ new_n1861;
  assign new_n1866 = ~new_n1863 & new_n1865;
  assign new_n1867 = new_n1866 ^ new_n1864;
  assign new_n1868 = new_n1677 ^ new_n1676;
  assign new_n1869 = new_n1868 ^ new_n1867;
  assign new_n1870 = n10 & n43;
  assign new_n1871 = new_n1870 ^ new_n1867;
  assign new_n1872 = ~new_n1869 & new_n1871;
  assign new_n1873 = new_n1872 ^ new_n1870;
  assign new_n1874 = new_n1683 ^ new_n1682;
  assign new_n1875 = new_n1874 ^ new_n1873;
  assign new_n1876 = n9 & n43;
  assign new_n1877 = new_n1876 ^ new_n1873;
  assign new_n1878 = ~new_n1875 & new_n1877;
  assign new_n1879 = new_n1878 ^ new_n1876;
  assign new_n1880 = new_n1689 ^ new_n1688;
  assign new_n1881 = new_n1880 ^ new_n1879;
  assign new_n1882 = n8 & n43;
  assign new_n1883 = new_n1882 ^ new_n1879;
  assign new_n1884 = ~new_n1881 & new_n1883;
  assign new_n1885 = new_n1884 ^ new_n1882;
  assign new_n1886 = new_n1695 ^ new_n1694;
  assign new_n1887 = new_n1886 ^ new_n1885;
  assign new_n1888 = n7 & n43;
  assign new_n1889 = new_n1888 ^ new_n1885;
  assign new_n1890 = ~new_n1887 & new_n1889;
  assign new_n1891 = new_n1890 ^ new_n1888;
  assign new_n1892 = new_n1701 ^ new_n1700;
  assign new_n1893 = new_n1892 ^ new_n1891;
  assign new_n1894 = n6 & n43;
  assign new_n1895 = new_n1894 ^ new_n1891;
  assign new_n1896 = ~new_n1893 & new_n1895;
  assign new_n1897 = new_n1896 ^ new_n1894;
  assign new_n1898 = new_n1707 ^ new_n1706;
  assign new_n1899 = new_n1898 ^ new_n1897;
  assign new_n1900 = n5 & n43;
  assign new_n1901 = new_n1900 ^ new_n1897;
  assign new_n1902 = ~new_n1899 & new_n1901;
  assign new_n1903 = new_n1902 ^ new_n1900;
  assign new_n1904 = new_n1713 ^ new_n1712;
  assign new_n1905 = new_n1904 ^ new_n1903;
  assign new_n1906 = n4 & n43;
  assign new_n1907 = new_n1906 ^ new_n1904;
  assign new_n1908 = ~new_n1905 & new_n1907;
  assign new_n1909 = new_n1908 ^ new_n1906;
  assign new_n1910 = new_n1719 ^ new_n1718;
  assign new_n1911 = new_n1910 ^ new_n1909;
  assign new_n1912 = n3 & n43;
  assign new_n1913 = new_n1912 ^ new_n1910;
  assign new_n1914 = ~new_n1911 & new_n1913;
  assign new_n1915 = new_n1914 ^ new_n1912;
  assign new_n1916 = new_n1725 ^ new_n1724;
  assign new_n1917 = new_n1916 ^ new_n1915;
  assign new_n1918 = n2 & n43;
  assign new_n1919 = new_n1918 ^ new_n1916;
  assign new_n1920 = ~new_n1917 & new_n1919;
  assign new_n1921 = new_n1920 ^ new_n1918;
  assign new_n1922 = new_n1731 ^ new_n1730;
  assign new_n1923 = new_n1922 ^ new_n1921;
  assign new_n1924 = n1 & n43;
  assign new_n1925 = new_n1924 ^ new_n1922;
  assign new_n1926 = ~new_n1923 & new_n1925;
  assign new_n1927 = new_n1926 ^ new_n1924;
  assign new_n1928 = new_n1744 & new_n1927;
  assign new_n1929 = new_n1928 ^ new_n1743;
  assign new_n1930 = new_n1927 ^ new_n1744;
  assign new_n1931 = new_n1924 ^ new_n1923;
  assign new_n1932 = new_n1747 ^ new_n1746;
  assign new_n1933 = n32 & n43;
  assign new_n1934 = n31 & n44;
  assign new_n1935 = new_n1933 & new_n1934;
  assign new_n1936 = new_n1935 ^ new_n1932;
  assign new_n1937 = n30 & n44;
  assign new_n1938 = new_n1937 ^ new_n1935;
  assign new_n1939 = ~new_n1936 & new_n1938;
  assign new_n1940 = new_n1939 ^ new_n1937;
  assign new_n1941 = new_n1750 ^ new_n1749;
  assign new_n1942 = new_n1941 ^ new_n1940;
  assign new_n1943 = n29 & n44;
  assign new_n1944 = new_n1943 ^ new_n1940;
  assign new_n1945 = ~new_n1942 & new_n1944;
  assign new_n1946 = new_n1945 ^ new_n1943;
  assign new_n1947 = new_n1756 ^ new_n1755;
  assign new_n1948 = new_n1947 ^ new_n1946;
  assign new_n1949 = n28 & n44;
  assign new_n1950 = new_n1949 ^ new_n1946;
  assign new_n1951 = ~new_n1948 & new_n1950;
  assign new_n1952 = new_n1951 ^ new_n1949;
  assign new_n1953 = new_n1762 ^ new_n1761;
  assign new_n1954 = new_n1953 ^ new_n1952;
  assign new_n1955 = n27 & n44;
  assign new_n1956 = new_n1955 ^ new_n1952;
  assign new_n1957 = ~new_n1954 & new_n1956;
  assign new_n1958 = new_n1957 ^ new_n1955;
  assign new_n1959 = new_n1768 ^ new_n1767;
  assign new_n1960 = new_n1959 ^ new_n1958;
  assign new_n1961 = n26 & n44;
  assign new_n1962 = new_n1961 ^ new_n1958;
  assign new_n1963 = ~new_n1960 & new_n1962;
  assign new_n1964 = new_n1963 ^ new_n1961;
  assign new_n1965 = new_n1774 ^ new_n1773;
  assign new_n1966 = new_n1965 ^ new_n1964;
  assign new_n1967 = n25 & n44;
  assign new_n1968 = new_n1967 ^ new_n1964;
  assign new_n1969 = ~new_n1966 & new_n1968;
  assign new_n1970 = new_n1969 ^ new_n1967;
  assign new_n1971 = new_n1780 ^ new_n1779;
  assign new_n1972 = new_n1971 ^ new_n1970;
  assign new_n1973 = n24 & n44;
  assign new_n1974 = new_n1973 ^ new_n1970;
  assign new_n1975 = ~new_n1972 & new_n1974;
  assign new_n1976 = new_n1975 ^ new_n1973;
  assign new_n1977 = new_n1786 ^ new_n1785;
  assign new_n1978 = new_n1977 ^ new_n1976;
  assign new_n1979 = n23 & n44;
  assign new_n1980 = new_n1979 ^ new_n1976;
  assign new_n1981 = ~new_n1978 & new_n1980;
  assign new_n1982 = new_n1981 ^ new_n1979;
  assign new_n1983 = new_n1792 ^ new_n1791;
  assign new_n1984 = new_n1983 ^ new_n1982;
  assign new_n1985 = n22 & n44;
  assign new_n1986 = new_n1985 ^ new_n1982;
  assign new_n1987 = ~new_n1984 & new_n1986;
  assign new_n1988 = new_n1987 ^ new_n1985;
  assign new_n1989 = new_n1798 ^ new_n1797;
  assign new_n1990 = new_n1989 ^ new_n1988;
  assign new_n1991 = n21 & n44;
  assign new_n1992 = new_n1991 ^ new_n1988;
  assign new_n1993 = ~new_n1990 & new_n1992;
  assign new_n1994 = new_n1993 ^ new_n1991;
  assign new_n1995 = new_n1804 ^ new_n1803;
  assign new_n1996 = new_n1995 ^ new_n1994;
  assign new_n1997 = n20 & n44;
  assign new_n1998 = new_n1997 ^ new_n1994;
  assign new_n1999 = ~new_n1996 & new_n1998;
  assign new_n2000 = new_n1999 ^ new_n1997;
  assign new_n2001 = new_n1810 ^ new_n1809;
  assign new_n2002 = new_n2001 ^ new_n2000;
  assign new_n2003 = n19 & n44;
  assign new_n2004 = new_n2003 ^ new_n2000;
  assign new_n2005 = ~new_n2002 & new_n2004;
  assign new_n2006 = new_n2005 ^ new_n2003;
  assign new_n2007 = new_n1816 ^ new_n1815;
  assign new_n2008 = new_n2007 ^ new_n2006;
  assign new_n2009 = n18 & n44;
  assign new_n2010 = new_n2009 ^ new_n2006;
  assign new_n2011 = ~new_n2008 & new_n2010;
  assign new_n2012 = new_n2011 ^ new_n2009;
  assign new_n2013 = new_n1822 ^ new_n1821;
  assign new_n2014 = new_n2013 ^ new_n2012;
  assign new_n2015 = n17 & n44;
  assign new_n2016 = new_n2015 ^ new_n2012;
  assign new_n2017 = ~new_n2014 & new_n2016;
  assign new_n2018 = new_n2017 ^ new_n2015;
  assign new_n2019 = new_n1828 ^ new_n1827;
  assign new_n2020 = new_n2019 ^ new_n2018;
  assign new_n2021 = n16 & n44;
  assign new_n2022 = new_n2021 ^ new_n2018;
  assign new_n2023 = ~new_n2020 & new_n2022;
  assign new_n2024 = new_n2023 ^ new_n2021;
  assign new_n2025 = new_n1834 ^ new_n1833;
  assign new_n2026 = new_n2025 ^ new_n2024;
  assign new_n2027 = n15 & n44;
  assign new_n2028 = new_n2027 ^ new_n2024;
  assign new_n2029 = ~new_n2026 & new_n2028;
  assign new_n2030 = new_n2029 ^ new_n2027;
  assign new_n2031 = new_n1840 ^ new_n1839;
  assign new_n2032 = new_n2031 ^ new_n2030;
  assign new_n2033 = n14 & n44;
  assign new_n2034 = new_n2033 ^ new_n2030;
  assign new_n2035 = ~new_n2032 & new_n2034;
  assign new_n2036 = new_n2035 ^ new_n2033;
  assign new_n2037 = new_n1846 ^ new_n1845;
  assign new_n2038 = new_n2037 ^ new_n2036;
  assign new_n2039 = n13 & n44;
  assign new_n2040 = new_n2039 ^ new_n2036;
  assign new_n2041 = ~new_n2038 & new_n2040;
  assign new_n2042 = new_n2041 ^ new_n2039;
  assign new_n2043 = new_n1852 ^ new_n1851;
  assign new_n2044 = new_n2043 ^ new_n2042;
  assign new_n2045 = n12 & n44;
  assign new_n2046 = new_n2045 ^ new_n2042;
  assign new_n2047 = ~new_n2044 & new_n2046;
  assign new_n2048 = new_n2047 ^ new_n2045;
  assign new_n2049 = new_n1858 ^ new_n1857;
  assign new_n2050 = new_n2049 ^ new_n2048;
  assign new_n2051 = n11 & n44;
  assign new_n2052 = new_n2051 ^ new_n2048;
  assign new_n2053 = ~new_n2050 & new_n2052;
  assign new_n2054 = new_n2053 ^ new_n2051;
  assign new_n2055 = new_n1864 ^ new_n1863;
  assign new_n2056 = new_n2055 ^ new_n2054;
  assign new_n2057 = n10 & n44;
  assign new_n2058 = new_n2057 ^ new_n2054;
  assign new_n2059 = ~new_n2056 & new_n2058;
  assign new_n2060 = new_n2059 ^ new_n2057;
  assign new_n2061 = new_n1870 ^ new_n1869;
  assign new_n2062 = new_n2061 ^ new_n2060;
  assign new_n2063 = n9 & n44;
  assign new_n2064 = new_n2063 ^ new_n2060;
  assign new_n2065 = ~new_n2062 & new_n2064;
  assign new_n2066 = new_n2065 ^ new_n2063;
  assign new_n2067 = new_n1876 ^ new_n1875;
  assign new_n2068 = new_n2067 ^ new_n2066;
  assign new_n2069 = n8 & n44;
  assign new_n2070 = new_n2069 ^ new_n2066;
  assign new_n2071 = ~new_n2068 & new_n2070;
  assign new_n2072 = new_n2071 ^ new_n2069;
  assign new_n2073 = new_n1882 ^ new_n1881;
  assign new_n2074 = new_n2073 ^ new_n2072;
  assign new_n2075 = n7 & n44;
  assign new_n2076 = new_n2075 ^ new_n2072;
  assign new_n2077 = ~new_n2074 & new_n2076;
  assign new_n2078 = new_n2077 ^ new_n2075;
  assign new_n2079 = new_n1888 ^ new_n1887;
  assign new_n2080 = new_n2079 ^ new_n2078;
  assign new_n2081 = n6 & n44;
  assign new_n2082 = new_n2081 ^ new_n2078;
  assign new_n2083 = ~new_n2080 & new_n2082;
  assign new_n2084 = new_n2083 ^ new_n2081;
  assign new_n2085 = new_n1894 ^ new_n1893;
  assign new_n2086 = new_n2085 ^ new_n2084;
  assign new_n2087 = n5 & n44;
  assign new_n2088 = new_n2087 ^ new_n2084;
  assign new_n2089 = ~new_n2086 & new_n2088;
  assign new_n2090 = new_n2089 ^ new_n2087;
  assign new_n2091 = new_n1900 ^ new_n1899;
  assign new_n2092 = new_n2091 ^ new_n2090;
  assign new_n2093 = n4 & n44;
  assign new_n2094 = new_n2093 ^ new_n2090;
  assign new_n2095 = ~new_n2092 & new_n2094;
  assign new_n2096 = new_n2095 ^ new_n2093;
  assign new_n2097 = new_n1906 ^ new_n1905;
  assign new_n2098 = new_n2097 ^ new_n2096;
  assign new_n2099 = n3 & n44;
  assign new_n2100 = new_n2099 ^ new_n2097;
  assign new_n2101 = ~new_n2098 & new_n2100;
  assign new_n2102 = new_n2101 ^ new_n2099;
  assign new_n2103 = new_n1912 ^ new_n1911;
  assign new_n2104 = new_n2103 ^ new_n2102;
  assign new_n2105 = n2 & n44;
  assign new_n2106 = new_n2105 ^ new_n2103;
  assign new_n2107 = ~new_n2104 & new_n2106;
  assign new_n2108 = new_n2107 ^ new_n2105;
  assign new_n2109 = new_n1918 ^ new_n1917;
  assign new_n2110 = new_n2109 ^ new_n2108;
  assign new_n2111 = n1 & n44;
  assign new_n2112 = new_n2111 ^ new_n2109;
  assign new_n2113 = ~new_n2110 & new_n2112;
  assign new_n2114 = new_n2113 ^ new_n2111;
  assign new_n2115 = new_n1931 & new_n2114;
  assign new_n2116 = new_n2115 ^ new_n1930;
  assign new_n2117 = new_n2114 ^ new_n1931;
  assign new_n2118 = new_n2111 ^ new_n2110;
  assign new_n2119 = new_n1934 ^ new_n1933;
  assign new_n2120 = n32 & n44;
  assign new_n2121 = n31 & n45;
  assign new_n2122 = new_n2120 & new_n2121;
  assign new_n2123 = new_n2122 ^ new_n2119;
  assign new_n2124 = n30 & n45;
  assign new_n2125 = new_n2124 ^ new_n2122;
  assign new_n2126 = ~new_n2123 & new_n2125;
  assign new_n2127 = new_n2126 ^ new_n2124;
  assign new_n2128 = new_n1937 ^ new_n1936;
  assign new_n2129 = new_n2128 ^ new_n2127;
  assign new_n2130 = n29 & n45;
  assign new_n2131 = new_n2130 ^ new_n2127;
  assign new_n2132 = ~new_n2129 & new_n2131;
  assign new_n2133 = new_n2132 ^ new_n2130;
  assign new_n2134 = new_n1943 ^ new_n1942;
  assign new_n2135 = new_n2134 ^ new_n2133;
  assign new_n2136 = n28 & n45;
  assign new_n2137 = new_n2136 ^ new_n2133;
  assign new_n2138 = ~new_n2135 & new_n2137;
  assign new_n2139 = new_n2138 ^ new_n2136;
  assign new_n2140 = new_n1949 ^ new_n1948;
  assign new_n2141 = new_n2140 ^ new_n2139;
  assign new_n2142 = n27 & n45;
  assign new_n2143 = new_n2142 ^ new_n2139;
  assign new_n2144 = ~new_n2141 & new_n2143;
  assign new_n2145 = new_n2144 ^ new_n2142;
  assign new_n2146 = new_n1955 ^ new_n1954;
  assign new_n2147 = new_n2146 ^ new_n2145;
  assign new_n2148 = n26 & n45;
  assign new_n2149 = new_n2148 ^ new_n2145;
  assign new_n2150 = ~new_n2147 & new_n2149;
  assign new_n2151 = new_n2150 ^ new_n2148;
  assign new_n2152 = new_n1961 ^ new_n1960;
  assign new_n2153 = new_n2152 ^ new_n2151;
  assign new_n2154 = n25 & n45;
  assign new_n2155 = new_n2154 ^ new_n2151;
  assign new_n2156 = ~new_n2153 & new_n2155;
  assign new_n2157 = new_n2156 ^ new_n2154;
  assign new_n2158 = new_n1967 ^ new_n1966;
  assign new_n2159 = new_n2158 ^ new_n2157;
  assign new_n2160 = n24 & n45;
  assign new_n2161 = new_n2160 ^ new_n2157;
  assign new_n2162 = ~new_n2159 & new_n2161;
  assign new_n2163 = new_n2162 ^ new_n2160;
  assign new_n2164 = new_n1973 ^ new_n1972;
  assign new_n2165 = new_n2164 ^ new_n2163;
  assign new_n2166 = n23 & n45;
  assign new_n2167 = new_n2166 ^ new_n2163;
  assign new_n2168 = ~new_n2165 & new_n2167;
  assign new_n2169 = new_n2168 ^ new_n2166;
  assign new_n2170 = new_n1979 ^ new_n1978;
  assign new_n2171 = new_n2170 ^ new_n2169;
  assign new_n2172 = n22 & n45;
  assign new_n2173 = new_n2172 ^ new_n2169;
  assign new_n2174 = ~new_n2171 & new_n2173;
  assign new_n2175 = new_n2174 ^ new_n2172;
  assign new_n2176 = new_n1985 ^ new_n1984;
  assign new_n2177 = new_n2176 ^ new_n2175;
  assign new_n2178 = n21 & n45;
  assign new_n2179 = new_n2178 ^ new_n2175;
  assign new_n2180 = ~new_n2177 & new_n2179;
  assign new_n2181 = new_n2180 ^ new_n2178;
  assign new_n2182 = new_n1991 ^ new_n1990;
  assign new_n2183 = new_n2182 ^ new_n2181;
  assign new_n2184 = n20 & n45;
  assign new_n2185 = new_n2184 ^ new_n2181;
  assign new_n2186 = ~new_n2183 & new_n2185;
  assign new_n2187 = new_n2186 ^ new_n2184;
  assign new_n2188 = new_n1997 ^ new_n1996;
  assign new_n2189 = new_n2188 ^ new_n2187;
  assign new_n2190 = n19 & n45;
  assign new_n2191 = new_n2190 ^ new_n2187;
  assign new_n2192 = ~new_n2189 & new_n2191;
  assign new_n2193 = new_n2192 ^ new_n2190;
  assign new_n2194 = new_n2003 ^ new_n2002;
  assign new_n2195 = new_n2194 ^ new_n2193;
  assign new_n2196 = n18 & n45;
  assign new_n2197 = new_n2196 ^ new_n2193;
  assign new_n2198 = ~new_n2195 & new_n2197;
  assign new_n2199 = new_n2198 ^ new_n2196;
  assign new_n2200 = new_n2009 ^ new_n2008;
  assign new_n2201 = new_n2200 ^ new_n2199;
  assign new_n2202 = n17 & n45;
  assign new_n2203 = new_n2202 ^ new_n2199;
  assign new_n2204 = ~new_n2201 & new_n2203;
  assign new_n2205 = new_n2204 ^ new_n2202;
  assign new_n2206 = new_n2015 ^ new_n2014;
  assign new_n2207 = new_n2206 ^ new_n2205;
  assign new_n2208 = n16 & n45;
  assign new_n2209 = new_n2208 ^ new_n2205;
  assign new_n2210 = ~new_n2207 & new_n2209;
  assign new_n2211 = new_n2210 ^ new_n2208;
  assign new_n2212 = new_n2021 ^ new_n2020;
  assign new_n2213 = new_n2212 ^ new_n2211;
  assign new_n2214 = n15 & n45;
  assign new_n2215 = new_n2214 ^ new_n2211;
  assign new_n2216 = ~new_n2213 & new_n2215;
  assign new_n2217 = new_n2216 ^ new_n2214;
  assign new_n2218 = new_n2027 ^ new_n2026;
  assign new_n2219 = new_n2218 ^ new_n2217;
  assign new_n2220 = n14 & n45;
  assign new_n2221 = new_n2220 ^ new_n2217;
  assign new_n2222 = ~new_n2219 & new_n2221;
  assign new_n2223 = new_n2222 ^ new_n2220;
  assign new_n2224 = new_n2033 ^ new_n2032;
  assign new_n2225 = new_n2224 ^ new_n2223;
  assign new_n2226 = n13 & n45;
  assign new_n2227 = new_n2226 ^ new_n2223;
  assign new_n2228 = ~new_n2225 & new_n2227;
  assign new_n2229 = new_n2228 ^ new_n2226;
  assign new_n2230 = new_n2039 ^ new_n2038;
  assign new_n2231 = new_n2230 ^ new_n2229;
  assign new_n2232 = n12 & n45;
  assign new_n2233 = new_n2232 ^ new_n2229;
  assign new_n2234 = ~new_n2231 & new_n2233;
  assign new_n2235 = new_n2234 ^ new_n2232;
  assign new_n2236 = new_n2045 ^ new_n2044;
  assign new_n2237 = new_n2236 ^ new_n2235;
  assign new_n2238 = n11 & n45;
  assign new_n2239 = new_n2238 ^ new_n2235;
  assign new_n2240 = ~new_n2237 & new_n2239;
  assign new_n2241 = new_n2240 ^ new_n2238;
  assign new_n2242 = new_n2051 ^ new_n2050;
  assign new_n2243 = new_n2242 ^ new_n2241;
  assign new_n2244 = n10 & n45;
  assign new_n2245 = new_n2244 ^ new_n2241;
  assign new_n2246 = ~new_n2243 & new_n2245;
  assign new_n2247 = new_n2246 ^ new_n2244;
  assign new_n2248 = new_n2057 ^ new_n2056;
  assign new_n2249 = new_n2248 ^ new_n2247;
  assign new_n2250 = n9 & n45;
  assign new_n2251 = new_n2250 ^ new_n2247;
  assign new_n2252 = ~new_n2249 & new_n2251;
  assign new_n2253 = new_n2252 ^ new_n2250;
  assign new_n2254 = new_n2063 ^ new_n2062;
  assign new_n2255 = new_n2254 ^ new_n2253;
  assign new_n2256 = n8 & n45;
  assign new_n2257 = new_n2256 ^ new_n2253;
  assign new_n2258 = ~new_n2255 & new_n2257;
  assign new_n2259 = new_n2258 ^ new_n2256;
  assign new_n2260 = new_n2069 ^ new_n2068;
  assign new_n2261 = new_n2260 ^ new_n2259;
  assign new_n2262 = n7 & n45;
  assign new_n2263 = new_n2262 ^ new_n2259;
  assign new_n2264 = ~new_n2261 & new_n2263;
  assign new_n2265 = new_n2264 ^ new_n2262;
  assign new_n2266 = new_n2075 ^ new_n2074;
  assign new_n2267 = new_n2266 ^ new_n2265;
  assign new_n2268 = n6 & n45;
  assign new_n2269 = new_n2268 ^ new_n2265;
  assign new_n2270 = ~new_n2267 & new_n2269;
  assign new_n2271 = new_n2270 ^ new_n2268;
  assign new_n2272 = new_n2081 ^ new_n2080;
  assign new_n2273 = new_n2272 ^ new_n2271;
  assign new_n2274 = n5 & n45;
  assign new_n2275 = new_n2274 ^ new_n2271;
  assign new_n2276 = ~new_n2273 & new_n2275;
  assign new_n2277 = new_n2276 ^ new_n2274;
  assign new_n2278 = new_n2087 ^ new_n2086;
  assign new_n2279 = new_n2278 ^ new_n2277;
  assign new_n2280 = n4 & n45;
  assign new_n2281 = new_n2280 ^ new_n2277;
  assign new_n2282 = ~new_n2279 & new_n2281;
  assign new_n2283 = new_n2282 ^ new_n2280;
  assign new_n2284 = new_n2093 ^ new_n2092;
  assign new_n2285 = new_n2284 ^ new_n2283;
  assign new_n2286 = n3 & n45;
  assign new_n2287 = new_n2286 ^ new_n2283;
  assign new_n2288 = ~new_n2285 & new_n2287;
  assign new_n2289 = new_n2288 ^ new_n2286;
  assign new_n2290 = new_n2099 ^ new_n2098;
  assign new_n2291 = new_n2290 ^ new_n2289;
  assign new_n2292 = n2 & n45;
  assign new_n2293 = new_n2292 ^ new_n2290;
  assign new_n2294 = ~new_n2291 & new_n2293;
  assign new_n2295 = new_n2294 ^ new_n2292;
  assign new_n2296 = new_n2105 ^ new_n2104;
  assign new_n2297 = new_n2296 ^ new_n2295;
  assign new_n2298 = n1 & n45;
  assign new_n2299 = new_n2298 ^ new_n2296;
  assign new_n2300 = ~new_n2297 & new_n2299;
  assign new_n2301 = new_n2300 ^ new_n2298;
  assign new_n2302 = new_n2118 & new_n2301;
  assign new_n2303 = new_n2302 ^ new_n2117;
  assign new_n2304 = new_n2301 ^ new_n2118;
  assign new_n2305 = new_n2298 ^ new_n2297;
  assign new_n2306 = new_n2121 ^ new_n2120;
  assign new_n2307 = n32 & n45;
  assign new_n2308 = n31 & n46;
  assign new_n2309 = new_n2307 & new_n2308;
  assign new_n2310 = new_n2309 ^ new_n2306;
  assign new_n2311 = n30 & n46;
  assign new_n2312 = new_n2311 ^ new_n2309;
  assign new_n2313 = ~new_n2310 & new_n2312;
  assign new_n2314 = new_n2313 ^ new_n2311;
  assign new_n2315 = new_n2124 ^ new_n2123;
  assign new_n2316 = new_n2315 ^ new_n2314;
  assign new_n2317 = n29 & n46;
  assign new_n2318 = new_n2317 ^ new_n2314;
  assign new_n2319 = ~new_n2316 & new_n2318;
  assign new_n2320 = new_n2319 ^ new_n2317;
  assign new_n2321 = new_n2130 ^ new_n2129;
  assign new_n2322 = new_n2321 ^ new_n2320;
  assign new_n2323 = n28 & n46;
  assign new_n2324 = new_n2323 ^ new_n2320;
  assign new_n2325 = ~new_n2322 & new_n2324;
  assign new_n2326 = new_n2325 ^ new_n2323;
  assign new_n2327 = new_n2136 ^ new_n2135;
  assign new_n2328 = new_n2327 ^ new_n2326;
  assign new_n2329 = n27 & n46;
  assign new_n2330 = new_n2329 ^ new_n2326;
  assign new_n2331 = ~new_n2328 & new_n2330;
  assign new_n2332 = new_n2331 ^ new_n2329;
  assign new_n2333 = new_n2142 ^ new_n2141;
  assign new_n2334 = new_n2333 ^ new_n2332;
  assign new_n2335 = n26 & n46;
  assign new_n2336 = new_n2335 ^ new_n2332;
  assign new_n2337 = ~new_n2334 & new_n2336;
  assign new_n2338 = new_n2337 ^ new_n2335;
  assign new_n2339 = new_n2148 ^ new_n2147;
  assign new_n2340 = new_n2339 ^ new_n2338;
  assign new_n2341 = n25 & n46;
  assign new_n2342 = new_n2341 ^ new_n2338;
  assign new_n2343 = ~new_n2340 & new_n2342;
  assign new_n2344 = new_n2343 ^ new_n2341;
  assign new_n2345 = new_n2154 ^ new_n2153;
  assign new_n2346 = new_n2345 ^ new_n2344;
  assign new_n2347 = n24 & n46;
  assign new_n2348 = new_n2347 ^ new_n2344;
  assign new_n2349 = ~new_n2346 & new_n2348;
  assign new_n2350 = new_n2349 ^ new_n2347;
  assign new_n2351 = new_n2160 ^ new_n2159;
  assign new_n2352 = new_n2351 ^ new_n2350;
  assign new_n2353 = n23 & n46;
  assign new_n2354 = new_n2353 ^ new_n2350;
  assign new_n2355 = ~new_n2352 & new_n2354;
  assign new_n2356 = new_n2355 ^ new_n2353;
  assign new_n2357 = new_n2166 ^ new_n2165;
  assign new_n2358 = new_n2357 ^ new_n2356;
  assign new_n2359 = n22 & n46;
  assign new_n2360 = new_n2359 ^ new_n2356;
  assign new_n2361 = ~new_n2358 & new_n2360;
  assign new_n2362 = new_n2361 ^ new_n2359;
  assign new_n2363 = new_n2172 ^ new_n2171;
  assign new_n2364 = new_n2363 ^ new_n2362;
  assign new_n2365 = n21 & n46;
  assign new_n2366 = new_n2365 ^ new_n2362;
  assign new_n2367 = ~new_n2364 & new_n2366;
  assign new_n2368 = new_n2367 ^ new_n2365;
  assign new_n2369 = new_n2178 ^ new_n2177;
  assign new_n2370 = new_n2369 ^ new_n2368;
  assign new_n2371 = n20 & n46;
  assign new_n2372 = new_n2371 ^ new_n2368;
  assign new_n2373 = ~new_n2370 & new_n2372;
  assign new_n2374 = new_n2373 ^ new_n2371;
  assign new_n2375 = new_n2184 ^ new_n2183;
  assign new_n2376 = new_n2375 ^ new_n2374;
  assign new_n2377 = n19 & n46;
  assign new_n2378 = new_n2377 ^ new_n2374;
  assign new_n2379 = ~new_n2376 & new_n2378;
  assign new_n2380 = new_n2379 ^ new_n2377;
  assign new_n2381 = new_n2190 ^ new_n2189;
  assign new_n2382 = new_n2381 ^ new_n2380;
  assign new_n2383 = n18 & n46;
  assign new_n2384 = new_n2383 ^ new_n2380;
  assign new_n2385 = ~new_n2382 & new_n2384;
  assign new_n2386 = new_n2385 ^ new_n2383;
  assign new_n2387 = new_n2196 ^ new_n2195;
  assign new_n2388 = new_n2387 ^ new_n2386;
  assign new_n2389 = n17 & n46;
  assign new_n2390 = new_n2389 ^ new_n2386;
  assign new_n2391 = ~new_n2388 & new_n2390;
  assign new_n2392 = new_n2391 ^ new_n2389;
  assign new_n2393 = new_n2202 ^ new_n2201;
  assign new_n2394 = new_n2393 ^ new_n2392;
  assign new_n2395 = n16 & n46;
  assign new_n2396 = new_n2395 ^ new_n2392;
  assign new_n2397 = ~new_n2394 & new_n2396;
  assign new_n2398 = new_n2397 ^ new_n2395;
  assign new_n2399 = new_n2208 ^ new_n2207;
  assign new_n2400 = new_n2399 ^ new_n2398;
  assign new_n2401 = n15 & n46;
  assign new_n2402 = new_n2401 ^ new_n2398;
  assign new_n2403 = ~new_n2400 & new_n2402;
  assign new_n2404 = new_n2403 ^ new_n2401;
  assign new_n2405 = new_n2214 ^ new_n2213;
  assign new_n2406 = new_n2405 ^ new_n2404;
  assign new_n2407 = n14 & n46;
  assign new_n2408 = new_n2407 ^ new_n2404;
  assign new_n2409 = ~new_n2406 & new_n2408;
  assign new_n2410 = new_n2409 ^ new_n2407;
  assign new_n2411 = new_n2220 ^ new_n2219;
  assign new_n2412 = new_n2411 ^ new_n2410;
  assign new_n2413 = n13 & n46;
  assign new_n2414 = new_n2413 ^ new_n2410;
  assign new_n2415 = ~new_n2412 & new_n2414;
  assign new_n2416 = new_n2415 ^ new_n2413;
  assign new_n2417 = new_n2226 ^ new_n2225;
  assign new_n2418 = new_n2417 ^ new_n2416;
  assign new_n2419 = n12 & n46;
  assign new_n2420 = new_n2419 ^ new_n2416;
  assign new_n2421 = ~new_n2418 & new_n2420;
  assign new_n2422 = new_n2421 ^ new_n2419;
  assign new_n2423 = new_n2232 ^ new_n2231;
  assign new_n2424 = new_n2423 ^ new_n2422;
  assign new_n2425 = n11 & n46;
  assign new_n2426 = new_n2425 ^ new_n2422;
  assign new_n2427 = ~new_n2424 & new_n2426;
  assign new_n2428 = new_n2427 ^ new_n2425;
  assign new_n2429 = new_n2238 ^ new_n2237;
  assign new_n2430 = new_n2429 ^ new_n2428;
  assign new_n2431 = n10 & n46;
  assign new_n2432 = new_n2431 ^ new_n2428;
  assign new_n2433 = ~new_n2430 & new_n2432;
  assign new_n2434 = new_n2433 ^ new_n2431;
  assign new_n2435 = new_n2244 ^ new_n2243;
  assign new_n2436 = new_n2435 ^ new_n2434;
  assign new_n2437 = n9 & n46;
  assign new_n2438 = new_n2437 ^ new_n2434;
  assign new_n2439 = ~new_n2436 & new_n2438;
  assign new_n2440 = new_n2439 ^ new_n2437;
  assign new_n2441 = new_n2250 ^ new_n2249;
  assign new_n2442 = new_n2441 ^ new_n2440;
  assign new_n2443 = n8 & n46;
  assign new_n2444 = new_n2443 ^ new_n2440;
  assign new_n2445 = ~new_n2442 & new_n2444;
  assign new_n2446 = new_n2445 ^ new_n2443;
  assign new_n2447 = new_n2256 ^ new_n2255;
  assign new_n2448 = new_n2447 ^ new_n2446;
  assign new_n2449 = n7 & n46;
  assign new_n2450 = new_n2449 ^ new_n2446;
  assign new_n2451 = ~new_n2448 & new_n2450;
  assign new_n2452 = new_n2451 ^ new_n2449;
  assign new_n2453 = new_n2262 ^ new_n2261;
  assign new_n2454 = new_n2453 ^ new_n2452;
  assign new_n2455 = n6 & n46;
  assign new_n2456 = new_n2455 ^ new_n2452;
  assign new_n2457 = ~new_n2454 & new_n2456;
  assign new_n2458 = new_n2457 ^ new_n2455;
  assign new_n2459 = new_n2268 ^ new_n2267;
  assign new_n2460 = new_n2459 ^ new_n2458;
  assign new_n2461 = n5 & n46;
  assign new_n2462 = new_n2461 ^ new_n2458;
  assign new_n2463 = ~new_n2460 & new_n2462;
  assign new_n2464 = new_n2463 ^ new_n2461;
  assign new_n2465 = new_n2274 ^ new_n2273;
  assign new_n2466 = new_n2465 ^ new_n2464;
  assign new_n2467 = n4 & n46;
  assign new_n2468 = new_n2467 ^ new_n2464;
  assign new_n2469 = ~new_n2466 & new_n2468;
  assign new_n2470 = new_n2469 ^ new_n2467;
  assign new_n2471 = new_n2280 ^ new_n2279;
  assign new_n2472 = new_n2471 ^ new_n2470;
  assign new_n2473 = n3 & n46;
  assign new_n2474 = new_n2473 ^ new_n2470;
  assign new_n2475 = ~new_n2472 & new_n2474;
  assign new_n2476 = new_n2475 ^ new_n2473;
  assign new_n2477 = new_n2286 ^ new_n2285;
  assign new_n2478 = new_n2477 ^ new_n2476;
  assign new_n2479 = n2 & n46;
  assign new_n2480 = new_n2479 ^ new_n2476;
  assign new_n2481 = ~new_n2478 & new_n2480;
  assign new_n2482 = new_n2481 ^ new_n2479;
  assign new_n2483 = new_n2292 ^ new_n2291;
  assign new_n2484 = new_n2483 ^ new_n2482;
  assign new_n2485 = n1 & n46;
  assign new_n2486 = new_n2485 ^ new_n2483;
  assign new_n2487 = ~new_n2484 & new_n2486;
  assign new_n2488 = new_n2487 ^ new_n2485;
  assign new_n2489 = new_n2305 & new_n2488;
  assign new_n2490 = new_n2489 ^ new_n2304;
  assign new_n2491 = new_n2488 ^ new_n2305;
  assign new_n2492 = new_n2485 ^ new_n2484;
  assign new_n2493 = new_n2308 ^ new_n2307;
  assign new_n2494 = n32 & n46;
  assign new_n2495 = n31 & n47;
  assign new_n2496 = new_n2494 & new_n2495;
  assign new_n2497 = new_n2496 ^ new_n2493;
  assign new_n2498 = n30 & n47;
  assign new_n2499 = new_n2498 ^ new_n2496;
  assign new_n2500 = ~new_n2497 & new_n2499;
  assign new_n2501 = new_n2500 ^ new_n2498;
  assign new_n2502 = new_n2311 ^ new_n2310;
  assign new_n2503 = new_n2502 ^ new_n2501;
  assign new_n2504 = n29 & n47;
  assign new_n2505 = new_n2504 ^ new_n2501;
  assign new_n2506 = ~new_n2503 & new_n2505;
  assign new_n2507 = new_n2506 ^ new_n2504;
  assign new_n2508 = new_n2317 ^ new_n2316;
  assign new_n2509 = new_n2508 ^ new_n2507;
  assign new_n2510 = n28 & n47;
  assign new_n2511 = new_n2510 ^ new_n2507;
  assign new_n2512 = ~new_n2509 & new_n2511;
  assign new_n2513 = new_n2512 ^ new_n2510;
  assign new_n2514 = new_n2323 ^ new_n2322;
  assign new_n2515 = new_n2514 ^ new_n2513;
  assign new_n2516 = n27 & n47;
  assign new_n2517 = new_n2516 ^ new_n2513;
  assign new_n2518 = ~new_n2515 & new_n2517;
  assign new_n2519 = new_n2518 ^ new_n2516;
  assign new_n2520 = new_n2329 ^ new_n2328;
  assign new_n2521 = new_n2520 ^ new_n2519;
  assign new_n2522 = n26 & n47;
  assign new_n2523 = new_n2522 ^ new_n2519;
  assign new_n2524 = ~new_n2521 & new_n2523;
  assign new_n2525 = new_n2524 ^ new_n2522;
  assign new_n2526 = new_n2335 ^ new_n2334;
  assign new_n2527 = new_n2526 ^ new_n2525;
  assign new_n2528 = n25 & n47;
  assign new_n2529 = new_n2528 ^ new_n2525;
  assign new_n2530 = ~new_n2527 & new_n2529;
  assign new_n2531 = new_n2530 ^ new_n2528;
  assign new_n2532 = new_n2341 ^ new_n2340;
  assign new_n2533 = new_n2532 ^ new_n2531;
  assign new_n2534 = n24 & n47;
  assign new_n2535 = new_n2534 ^ new_n2531;
  assign new_n2536 = ~new_n2533 & new_n2535;
  assign new_n2537 = new_n2536 ^ new_n2534;
  assign new_n2538 = new_n2347 ^ new_n2346;
  assign new_n2539 = new_n2538 ^ new_n2537;
  assign new_n2540 = n23 & n47;
  assign new_n2541 = new_n2540 ^ new_n2537;
  assign new_n2542 = ~new_n2539 & new_n2541;
  assign new_n2543 = new_n2542 ^ new_n2540;
  assign new_n2544 = new_n2353 ^ new_n2352;
  assign new_n2545 = new_n2544 ^ new_n2543;
  assign new_n2546 = n22 & n47;
  assign new_n2547 = new_n2546 ^ new_n2543;
  assign new_n2548 = ~new_n2545 & new_n2547;
  assign new_n2549 = new_n2548 ^ new_n2546;
  assign new_n2550 = new_n2359 ^ new_n2358;
  assign new_n2551 = new_n2550 ^ new_n2549;
  assign new_n2552 = n21 & n47;
  assign new_n2553 = new_n2552 ^ new_n2549;
  assign new_n2554 = ~new_n2551 & new_n2553;
  assign new_n2555 = new_n2554 ^ new_n2552;
  assign new_n2556 = new_n2365 ^ new_n2364;
  assign new_n2557 = new_n2556 ^ new_n2555;
  assign new_n2558 = n20 & n47;
  assign new_n2559 = new_n2558 ^ new_n2555;
  assign new_n2560 = ~new_n2557 & new_n2559;
  assign new_n2561 = new_n2560 ^ new_n2558;
  assign new_n2562 = new_n2371 ^ new_n2370;
  assign new_n2563 = new_n2562 ^ new_n2561;
  assign new_n2564 = n19 & n47;
  assign new_n2565 = new_n2564 ^ new_n2561;
  assign new_n2566 = ~new_n2563 & new_n2565;
  assign new_n2567 = new_n2566 ^ new_n2564;
  assign new_n2568 = new_n2377 ^ new_n2376;
  assign new_n2569 = new_n2568 ^ new_n2567;
  assign new_n2570 = n18 & n47;
  assign new_n2571 = new_n2570 ^ new_n2567;
  assign new_n2572 = ~new_n2569 & new_n2571;
  assign new_n2573 = new_n2572 ^ new_n2570;
  assign new_n2574 = new_n2383 ^ new_n2382;
  assign new_n2575 = new_n2574 ^ new_n2573;
  assign new_n2576 = n17 & n47;
  assign new_n2577 = new_n2576 ^ new_n2573;
  assign new_n2578 = ~new_n2575 & new_n2577;
  assign new_n2579 = new_n2578 ^ new_n2576;
  assign new_n2580 = new_n2389 ^ new_n2388;
  assign new_n2581 = new_n2580 ^ new_n2579;
  assign new_n2582 = n16 & n47;
  assign new_n2583 = new_n2582 ^ new_n2579;
  assign new_n2584 = ~new_n2581 & new_n2583;
  assign new_n2585 = new_n2584 ^ new_n2582;
  assign new_n2586 = new_n2395 ^ new_n2394;
  assign new_n2587 = new_n2586 ^ new_n2585;
  assign new_n2588 = n15 & n47;
  assign new_n2589 = new_n2588 ^ new_n2585;
  assign new_n2590 = ~new_n2587 & new_n2589;
  assign new_n2591 = new_n2590 ^ new_n2588;
  assign new_n2592 = new_n2401 ^ new_n2400;
  assign new_n2593 = new_n2592 ^ new_n2591;
  assign new_n2594 = n14 & n47;
  assign new_n2595 = new_n2594 ^ new_n2591;
  assign new_n2596 = ~new_n2593 & new_n2595;
  assign new_n2597 = new_n2596 ^ new_n2594;
  assign new_n2598 = new_n2407 ^ new_n2406;
  assign new_n2599 = new_n2598 ^ new_n2597;
  assign new_n2600 = n13 & n47;
  assign new_n2601 = new_n2600 ^ new_n2597;
  assign new_n2602 = ~new_n2599 & new_n2601;
  assign new_n2603 = new_n2602 ^ new_n2600;
  assign new_n2604 = new_n2413 ^ new_n2412;
  assign new_n2605 = new_n2604 ^ new_n2603;
  assign new_n2606 = n12 & n47;
  assign new_n2607 = new_n2606 ^ new_n2603;
  assign new_n2608 = ~new_n2605 & new_n2607;
  assign new_n2609 = new_n2608 ^ new_n2606;
  assign new_n2610 = new_n2419 ^ new_n2418;
  assign new_n2611 = new_n2610 ^ new_n2609;
  assign new_n2612 = n11 & n47;
  assign new_n2613 = new_n2612 ^ new_n2609;
  assign new_n2614 = ~new_n2611 & new_n2613;
  assign new_n2615 = new_n2614 ^ new_n2612;
  assign new_n2616 = new_n2425 ^ new_n2424;
  assign new_n2617 = new_n2616 ^ new_n2615;
  assign new_n2618 = n10 & n47;
  assign new_n2619 = new_n2618 ^ new_n2615;
  assign new_n2620 = ~new_n2617 & new_n2619;
  assign new_n2621 = new_n2620 ^ new_n2618;
  assign new_n2622 = new_n2431 ^ new_n2430;
  assign new_n2623 = new_n2622 ^ new_n2621;
  assign new_n2624 = n9 & n47;
  assign new_n2625 = new_n2624 ^ new_n2621;
  assign new_n2626 = ~new_n2623 & new_n2625;
  assign new_n2627 = new_n2626 ^ new_n2624;
  assign new_n2628 = new_n2437 ^ new_n2436;
  assign new_n2629 = new_n2628 ^ new_n2627;
  assign new_n2630 = n8 & n47;
  assign new_n2631 = new_n2630 ^ new_n2627;
  assign new_n2632 = ~new_n2629 & new_n2631;
  assign new_n2633 = new_n2632 ^ new_n2630;
  assign new_n2634 = new_n2443 ^ new_n2442;
  assign new_n2635 = new_n2634 ^ new_n2633;
  assign new_n2636 = n7 & n47;
  assign new_n2637 = new_n2636 ^ new_n2633;
  assign new_n2638 = ~new_n2635 & new_n2637;
  assign new_n2639 = new_n2638 ^ new_n2636;
  assign new_n2640 = new_n2449 ^ new_n2448;
  assign new_n2641 = new_n2640 ^ new_n2639;
  assign new_n2642 = n6 & n47;
  assign new_n2643 = new_n2642 ^ new_n2639;
  assign new_n2644 = ~new_n2641 & new_n2643;
  assign new_n2645 = new_n2644 ^ new_n2642;
  assign new_n2646 = new_n2455 ^ new_n2454;
  assign new_n2647 = new_n2646 ^ new_n2645;
  assign new_n2648 = n5 & n47;
  assign new_n2649 = new_n2648 ^ new_n2645;
  assign new_n2650 = ~new_n2647 & new_n2649;
  assign new_n2651 = new_n2650 ^ new_n2648;
  assign new_n2652 = new_n2461 ^ new_n2460;
  assign new_n2653 = new_n2652 ^ new_n2651;
  assign new_n2654 = n4 & n47;
  assign new_n2655 = new_n2654 ^ new_n2651;
  assign new_n2656 = ~new_n2653 & new_n2655;
  assign new_n2657 = new_n2656 ^ new_n2654;
  assign new_n2658 = new_n2467 ^ new_n2466;
  assign new_n2659 = new_n2658 ^ new_n2657;
  assign new_n2660 = n3 & n47;
  assign new_n2661 = new_n2660 ^ new_n2657;
  assign new_n2662 = ~new_n2659 & new_n2661;
  assign new_n2663 = new_n2662 ^ new_n2660;
  assign new_n2664 = new_n2473 ^ new_n2472;
  assign new_n2665 = new_n2664 ^ new_n2663;
  assign new_n2666 = n2 & n47;
  assign new_n2667 = new_n2666 ^ new_n2663;
  assign new_n2668 = ~new_n2665 & new_n2667;
  assign new_n2669 = new_n2668 ^ new_n2666;
  assign new_n2670 = new_n2479 ^ new_n2478;
  assign new_n2671 = new_n2670 ^ new_n2669;
  assign new_n2672 = n1 & n47;
  assign new_n2673 = new_n2672 ^ new_n2669;
  assign new_n2674 = ~new_n2671 & new_n2673;
  assign new_n2675 = new_n2674 ^ new_n2672;
  assign new_n2676 = new_n2492 & new_n2675;
  assign new_n2677 = new_n2676 ^ new_n2491;
  assign new_n2678 = new_n2675 ^ new_n2492;
  assign new_n2679 = new_n2672 ^ new_n2671;
  assign new_n2680 = new_n2660 ^ new_n2659;
  assign new_n2681 = new_n2648 ^ new_n2647;
  assign new_n2682 = new_n2636 ^ new_n2635;
  assign new_n2683 = new_n2624 ^ new_n2623;
  assign new_n2684 = new_n2612 ^ new_n2611;
  assign new_n2685 = new_n2600 ^ new_n2599;
  assign new_n2686 = new_n2588 ^ new_n2587;
  assign new_n2687 = new_n2576 ^ new_n2575;
  assign new_n2688 = new_n2564 ^ new_n2563;
  assign new_n2689 = new_n2552 ^ new_n2551;
  assign new_n2690 = new_n2540 ^ new_n2539;
  assign new_n2691 = new_n2528 ^ new_n2527;
  assign new_n2692 = new_n2516 ^ new_n2515;
  assign new_n2693 = new_n2504 ^ new_n2503;
  assign new_n2694 = new_n2498 ^ new_n2497;
  assign new_n2695 = n32 & n47;
  assign new_n2696 = n31 & n48;
  assign new_n2697 = new_n2695 & new_n2696;
  assign new_n2698 = new_n2495 ^ new_n2494;
  assign new_n2699 = new_n2698 ^ new_n2697;
  assign new_n2700 = n30 & n48;
  assign new_n2701 = new_n2700 ^ new_n2697;
  assign new_n2702 = ~new_n2699 & new_n2701;
  assign new_n2703 = new_n2702 ^ new_n2700;
  assign new_n2704 = new_n2703 ^ new_n2694;
  assign new_n2705 = n29 & n48;
  assign new_n2706 = new_n2705 ^ new_n2703;
  assign new_n2707 = ~new_n2704 & new_n2706;
  assign new_n2708 = new_n2707 ^ new_n2705;
  assign new_n2709 = new_n2708 ^ new_n2693;
  assign new_n2710 = n28 & n48;
  assign new_n2711 = new_n2710 ^ new_n2708;
  assign new_n2712 = ~new_n2709 & new_n2711;
  assign new_n2713 = new_n2712 ^ new_n2710;
  assign new_n2714 = new_n2510 ^ new_n2509;
  assign new_n2715 = new_n2714 ^ new_n2713;
  assign new_n2716 = n27 & n48;
  assign new_n2717 = new_n2716 ^ new_n2713;
  assign new_n2718 = ~new_n2715 & new_n2717;
  assign new_n2719 = new_n2718 ^ new_n2716;
  assign new_n2720 = new_n2719 ^ new_n2692;
  assign new_n2721 = n26 & n48;
  assign new_n2722 = new_n2721 ^ new_n2719;
  assign new_n2723 = ~new_n2720 & new_n2722;
  assign new_n2724 = new_n2723 ^ new_n2721;
  assign new_n2725 = new_n2522 ^ new_n2521;
  assign new_n2726 = new_n2725 ^ new_n2724;
  assign new_n2727 = n25 & n48;
  assign new_n2728 = new_n2727 ^ new_n2724;
  assign new_n2729 = ~new_n2726 & new_n2728;
  assign new_n2730 = new_n2729 ^ new_n2727;
  assign new_n2731 = new_n2730 ^ new_n2691;
  assign new_n2732 = n24 & n48;
  assign new_n2733 = new_n2732 ^ new_n2730;
  assign new_n2734 = ~new_n2731 & new_n2733;
  assign new_n2735 = new_n2734 ^ new_n2732;
  assign new_n2736 = new_n2534 ^ new_n2533;
  assign new_n2737 = new_n2736 ^ new_n2735;
  assign new_n2738 = n23 & n48;
  assign new_n2739 = new_n2738 ^ new_n2735;
  assign new_n2740 = ~new_n2737 & new_n2739;
  assign new_n2741 = new_n2740 ^ new_n2738;
  assign new_n2742 = new_n2741 ^ new_n2690;
  assign new_n2743 = n22 & n48;
  assign new_n2744 = new_n2743 ^ new_n2741;
  assign new_n2745 = ~new_n2742 & new_n2744;
  assign new_n2746 = new_n2745 ^ new_n2743;
  assign new_n2747 = new_n2546 ^ new_n2545;
  assign new_n2748 = new_n2747 ^ new_n2746;
  assign new_n2749 = n21 & n48;
  assign new_n2750 = new_n2749 ^ new_n2746;
  assign new_n2751 = ~new_n2748 & new_n2750;
  assign new_n2752 = new_n2751 ^ new_n2749;
  assign new_n2753 = new_n2752 ^ new_n2689;
  assign new_n2754 = n20 & n48;
  assign new_n2755 = new_n2754 ^ new_n2752;
  assign new_n2756 = ~new_n2753 & new_n2755;
  assign new_n2757 = new_n2756 ^ new_n2754;
  assign new_n2758 = new_n2558 ^ new_n2557;
  assign new_n2759 = new_n2758 ^ new_n2757;
  assign new_n2760 = n19 & n48;
  assign new_n2761 = new_n2760 ^ new_n2757;
  assign new_n2762 = ~new_n2759 & new_n2761;
  assign new_n2763 = new_n2762 ^ new_n2760;
  assign new_n2764 = new_n2763 ^ new_n2688;
  assign new_n2765 = n18 & n48;
  assign new_n2766 = new_n2765 ^ new_n2763;
  assign new_n2767 = ~new_n2764 & new_n2766;
  assign new_n2768 = new_n2767 ^ new_n2765;
  assign new_n2769 = new_n2570 ^ new_n2569;
  assign new_n2770 = new_n2769 ^ new_n2768;
  assign new_n2771 = n17 & n48;
  assign new_n2772 = new_n2771 ^ new_n2768;
  assign new_n2773 = ~new_n2770 & new_n2772;
  assign new_n2774 = new_n2773 ^ new_n2771;
  assign new_n2775 = new_n2774 ^ new_n2687;
  assign new_n2776 = n16 & n48;
  assign new_n2777 = new_n2776 ^ new_n2774;
  assign new_n2778 = ~new_n2775 & new_n2777;
  assign new_n2779 = new_n2778 ^ new_n2776;
  assign new_n2780 = new_n2582 ^ new_n2581;
  assign new_n2781 = new_n2780 ^ new_n2779;
  assign new_n2782 = n15 & n48;
  assign new_n2783 = new_n2782 ^ new_n2779;
  assign new_n2784 = ~new_n2781 & new_n2783;
  assign new_n2785 = new_n2784 ^ new_n2782;
  assign new_n2786 = new_n2785 ^ new_n2686;
  assign new_n2787 = n14 & n48;
  assign new_n2788 = new_n2787 ^ new_n2785;
  assign new_n2789 = ~new_n2786 & new_n2788;
  assign new_n2790 = new_n2789 ^ new_n2787;
  assign new_n2791 = new_n2594 ^ new_n2593;
  assign new_n2792 = new_n2791 ^ new_n2790;
  assign new_n2793 = n13 & n48;
  assign new_n2794 = new_n2793 ^ new_n2790;
  assign new_n2795 = ~new_n2792 & new_n2794;
  assign new_n2796 = new_n2795 ^ new_n2793;
  assign new_n2797 = new_n2796 ^ new_n2685;
  assign new_n2798 = n12 & n48;
  assign new_n2799 = new_n2798 ^ new_n2796;
  assign new_n2800 = ~new_n2797 & new_n2799;
  assign new_n2801 = new_n2800 ^ new_n2798;
  assign new_n2802 = new_n2606 ^ new_n2605;
  assign new_n2803 = new_n2802 ^ new_n2801;
  assign new_n2804 = n11 & n48;
  assign new_n2805 = new_n2804 ^ new_n2801;
  assign new_n2806 = ~new_n2803 & new_n2805;
  assign new_n2807 = new_n2806 ^ new_n2804;
  assign new_n2808 = new_n2807 ^ new_n2684;
  assign new_n2809 = n10 & n48;
  assign new_n2810 = new_n2809 ^ new_n2807;
  assign new_n2811 = ~new_n2808 & new_n2810;
  assign new_n2812 = new_n2811 ^ new_n2809;
  assign new_n2813 = new_n2618 ^ new_n2617;
  assign new_n2814 = new_n2813 ^ new_n2812;
  assign new_n2815 = n9 & n48;
  assign new_n2816 = new_n2815 ^ new_n2812;
  assign new_n2817 = ~new_n2814 & new_n2816;
  assign new_n2818 = new_n2817 ^ new_n2815;
  assign new_n2819 = new_n2818 ^ new_n2683;
  assign new_n2820 = n8 & n48;
  assign new_n2821 = new_n2820 ^ new_n2818;
  assign new_n2822 = ~new_n2819 & new_n2821;
  assign new_n2823 = new_n2822 ^ new_n2820;
  assign new_n2824 = new_n2630 ^ new_n2629;
  assign new_n2825 = new_n2824 ^ new_n2823;
  assign new_n2826 = n7 & n48;
  assign new_n2827 = new_n2826 ^ new_n2823;
  assign new_n2828 = ~new_n2825 & new_n2827;
  assign new_n2829 = new_n2828 ^ new_n2826;
  assign new_n2830 = new_n2829 ^ new_n2682;
  assign new_n2831 = n6 & n48;
  assign new_n2832 = new_n2831 ^ new_n2829;
  assign new_n2833 = ~new_n2830 & new_n2832;
  assign new_n2834 = new_n2833 ^ new_n2831;
  assign new_n2835 = new_n2642 ^ new_n2641;
  assign new_n2836 = new_n2835 ^ new_n2834;
  assign new_n2837 = n5 & n48;
  assign new_n2838 = new_n2837 ^ new_n2834;
  assign new_n2839 = ~new_n2836 & new_n2838;
  assign new_n2840 = new_n2839 ^ new_n2837;
  assign new_n2841 = new_n2840 ^ new_n2681;
  assign new_n2842 = n4 & n48;
  assign new_n2843 = new_n2842 ^ new_n2840;
  assign new_n2844 = ~new_n2841 & new_n2843;
  assign new_n2845 = new_n2844 ^ new_n2842;
  assign new_n2846 = new_n2654 ^ new_n2653;
  assign new_n2847 = new_n2846 ^ new_n2845;
  assign new_n2848 = n3 & n48;
  assign new_n2849 = new_n2848 ^ new_n2845;
  assign new_n2850 = ~new_n2847 & new_n2849;
  assign new_n2851 = new_n2850 ^ new_n2848;
  assign new_n2852 = new_n2851 ^ new_n2680;
  assign new_n2853 = n2 & n48;
  assign new_n2854 = new_n2853 ^ new_n2851;
  assign new_n2855 = ~new_n2852 & new_n2854;
  assign new_n2856 = new_n2855 ^ new_n2853;
  assign new_n2857 = new_n2666 ^ new_n2665;
  assign new_n2858 = new_n2857 ^ new_n2856;
  assign new_n2859 = n1 & n48;
  assign new_n2860 = new_n2859 ^ new_n2856;
  assign new_n2861 = ~new_n2858 & new_n2860;
  assign new_n2862 = new_n2861 ^ new_n2859;
  assign new_n2863 = new_n2679 & new_n2862;
  assign new_n2864 = new_n2863 ^ new_n2678;
  assign new_n2865 = new_n2862 ^ new_n2679;
  assign new_n2866 = new_n2859 ^ new_n2858;
  assign new_n2867 = new_n2848 ^ new_n2847;
  assign new_n2868 = new_n2837 ^ new_n2836;
  assign new_n2869 = new_n2826 ^ new_n2825;
  assign new_n2870 = new_n2815 ^ new_n2814;
  assign new_n2871 = new_n2804 ^ new_n2803;
  assign new_n2872 = new_n2793 ^ new_n2792;
  assign new_n2873 = new_n2782 ^ new_n2781;
  assign new_n2874 = new_n2771 ^ new_n2770;
  assign new_n2875 = new_n2760 ^ new_n2759;
  assign new_n2876 = new_n2749 ^ new_n2748;
  assign new_n2877 = new_n2738 ^ new_n2737;
  assign new_n2878 = new_n2727 ^ new_n2726;
  assign new_n2879 = new_n2716 ^ new_n2715;
  assign new_n2880 = new_n2705 ^ new_n2704;
  assign new_n2881 = new_n2700 ^ new_n2699;
  assign new_n2882 = n32 & n48;
  assign new_n2883 = n31 & n49;
  assign new_n2884 = new_n2882 & new_n2883;
  assign new_n2885 = new_n2696 ^ new_n2695;
  assign new_n2886 = new_n2885 ^ new_n2884;
  assign new_n2887 = n30 & n49;
  assign new_n2888 = new_n2887 ^ new_n2884;
  assign new_n2889 = ~new_n2886 & new_n2888;
  assign new_n2890 = new_n2889 ^ new_n2887;
  assign new_n2891 = new_n2890 ^ new_n2881;
  assign new_n2892 = n29 & n49;
  assign new_n2893 = new_n2892 ^ new_n2890;
  assign new_n2894 = ~new_n2891 & new_n2893;
  assign new_n2895 = new_n2894 ^ new_n2892;
  assign new_n2896 = new_n2895 ^ new_n2880;
  assign new_n2897 = n28 & n49;
  assign new_n2898 = new_n2897 ^ new_n2895;
  assign new_n2899 = ~new_n2896 & new_n2898;
  assign new_n2900 = new_n2899 ^ new_n2897;
  assign new_n2901 = new_n2710 ^ new_n2709;
  assign new_n2902 = new_n2901 ^ new_n2900;
  assign new_n2903 = n27 & n49;
  assign new_n2904 = new_n2903 ^ new_n2900;
  assign new_n2905 = ~new_n2902 & new_n2904;
  assign new_n2906 = new_n2905 ^ new_n2903;
  assign new_n2907 = new_n2906 ^ new_n2879;
  assign new_n2908 = n26 & n49;
  assign new_n2909 = new_n2908 ^ new_n2906;
  assign new_n2910 = ~new_n2907 & new_n2909;
  assign new_n2911 = new_n2910 ^ new_n2908;
  assign new_n2912 = new_n2721 ^ new_n2720;
  assign new_n2913 = new_n2912 ^ new_n2911;
  assign new_n2914 = n25 & n49;
  assign new_n2915 = new_n2914 ^ new_n2911;
  assign new_n2916 = ~new_n2913 & new_n2915;
  assign new_n2917 = new_n2916 ^ new_n2914;
  assign new_n2918 = new_n2917 ^ new_n2878;
  assign new_n2919 = n24 & n49;
  assign new_n2920 = new_n2919 ^ new_n2917;
  assign new_n2921 = ~new_n2918 & new_n2920;
  assign new_n2922 = new_n2921 ^ new_n2919;
  assign new_n2923 = new_n2732 ^ new_n2731;
  assign new_n2924 = new_n2923 ^ new_n2922;
  assign new_n2925 = n23 & n49;
  assign new_n2926 = new_n2925 ^ new_n2922;
  assign new_n2927 = ~new_n2924 & new_n2926;
  assign new_n2928 = new_n2927 ^ new_n2925;
  assign new_n2929 = new_n2928 ^ new_n2877;
  assign new_n2930 = n22 & n49;
  assign new_n2931 = new_n2930 ^ new_n2928;
  assign new_n2932 = ~new_n2929 & new_n2931;
  assign new_n2933 = new_n2932 ^ new_n2930;
  assign new_n2934 = new_n2743 ^ new_n2742;
  assign new_n2935 = new_n2934 ^ new_n2933;
  assign new_n2936 = n21 & n49;
  assign new_n2937 = new_n2936 ^ new_n2933;
  assign new_n2938 = ~new_n2935 & new_n2937;
  assign new_n2939 = new_n2938 ^ new_n2936;
  assign new_n2940 = new_n2939 ^ new_n2876;
  assign new_n2941 = n20 & n49;
  assign new_n2942 = new_n2941 ^ new_n2939;
  assign new_n2943 = ~new_n2940 & new_n2942;
  assign new_n2944 = new_n2943 ^ new_n2941;
  assign new_n2945 = new_n2754 ^ new_n2753;
  assign new_n2946 = new_n2945 ^ new_n2944;
  assign new_n2947 = n19 & n49;
  assign new_n2948 = new_n2947 ^ new_n2944;
  assign new_n2949 = ~new_n2946 & new_n2948;
  assign new_n2950 = new_n2949 ^ new_n2947;
  assign new_n2951 = new_n2950 ^ new_n2875;
  assign new_n2952 = n18 & n49;
  assign new_n2953 = new_n2952 ^ new_n2950;
  assign new_n2954 = ~new_n2951 & new_n2953;
  assign new_n2955 = new_n2954 ^ new_n2952;
  assign new_n2956 = new_n2765 ^ new_n2764;
  assign new_n2957 = new_n2956 ^ new_n2955;
  assign new_n2958 = n17 & n49;
  assign new_n2959 = new_n2958 ^ new_n2955;
  assign new_n2960 = ~new_n2957 & new_n2959;
  assign new_n2961 = new_n2960 ^ new_n2958;
  assign new_n2962 = new_n2961 ^ new_n2874;
  assign new_n2963 = n16 & n49;
  assign new_n2964 = new_n2963 ^ new_n2961;
  assign new_n2965 = ~new_n2962 & new_n2964;
  assign new_n2966 = new_n2965 ^ new_n2963;
  assign new_n2967 = new_n2776 ^ new_n2775;
  assign new_n2968 = new_n2967 ^ new_n2966;
  assign new_n2969 = n15 & n49;
  assign new_n2970 = new_n2969 ^ new_n2966;
  assign new_n2971 = ~new_n2968 & new_n2970;
  assign new_n2972 = new_n2971 ^ new_n2969;
  assign new_n2973 = new_n2972 ^ new_n2873;
  assign new_n2974 = n14 & n49;
  assign new_n2975 = new_n2974 ^ new_n2972;
  assign new_n2976 = ~new_n2973 & new_n2975;
  assign new_n2977 = new_n2976 ^ new_n2974;
  assign new_n2978 = new_n2787 ^ new_n2786;
  assign new_n2979 = new_n2978 ^ new_n2977;
  assign new_n2980 = n13 & n49;
  assign new_n2981 = new_n2980 ^ new_n2977;
  assign new_n2982 = ~new_n2979 & new_n2981;
  assign new_n2983 = new_n2982 ^ new_n2980;
  assign new_n2984 = new_n2983 ^ new_n2872;
  assign new_n2985 = n12 & n49;
  assign new_n2986 = new_n2985 ^ new_n2983;
  assign new_n2987 = ~new_n2984 & new_n2986;
  assign new_n2988 = new_n2987 ^ new_n2985;
  assign new_n2989 = new_n2798 ^ new_n2797;
  assign new_n2990 = new_n2989 ^ new_n2988;
  assign new_n2991 = n11 & n49;
  assign new_n2992 = new_n2991 ^ new_n2988;
  assign new_n2993 = ~new_n2990 & new_n2992;
  assign new_n2994 = new_n2993 ^ new_n2991;
  assign new_n2995 = new_n2994 ^ new_n2871;
  assign new_n2996 = n10 & n49;
  assign new_n2997 = new_n2996 ^ new_n2994;
  assign new_n2998 = ~new_n2995 & new_n2997;
  assign new_n2999 = new_n2998 ^ new_n2996;
  assign new_n3000 = new_n2809 ^ new_n2808;
  assign new_n3001 = new_n3000 ^ new_n2999;
  assign new_n3002 = n9 & n49;
  assign new_n3003 = new_n3002 ^ new_n2999;
  assign new_n3004 = ~new_n3001 & new_n3003;
  assign new_n3005 = new_n3004 ^ new_n3002;
  assign new_n3006 = new_n3005 ^ new_n2870;
  assign new_n3007 = n8 & n49;
  assign new_n3008 = new_n3007 ^ new_n3005;
  assign new_n3009 = ~new_n3006 & new_n3008;
  assign new_n3010 = new_n3009 ^ new_n3007;
  assign new_n3011 = new_n2820 ^ new_n2819;
  assign new_n3012 = new_n3011 ^ new_n3010;
  assign new_n3013 = n7 & n49;
  assign new_n3014 = new_n3013 ^ new_n3010;
  assign new_n3015 = ~new_n3012 & new_n3014;
  assign new_n3016 = new_n3015 ^ new_n3013;
  assign new_n3017 = new_n3016 ^ new_n2869;
  assign new_n3018 = n6 & n49;
  assign new_n3019 = new_n3018 ^ new_n3016;
  assign new_n3020 = ~new_n3017 & new_n3019;
  assign new_n3021 = new_n3020 ^ new_n3018;
  assign new_n3022 = new_n2831 ^ new_n2830;
  assign new_n3023 = new_n3022 ^ new_n3021;
  assign new_n3024 = n5 & n49;
  assign new_n3025 = new_n3024 ^ new_n3021;
  assign new_n3026 = ~new_n3023 & new_n3025;
  assign new_n3027 = new_n3026 ^ new_n3024;
  assign new_n3028 = new_n3027 ^ new_n2868;
  assign new_n3029 = n4 & n49;
  assign new_n3030 = new_n3029 ^ new_n3027;
  assign new_n3031 = ~new_n3028 & new_n3030;
  assign new_n3032 = new_n3031 ^ new_n3029;
  assign new_n3033 = new_n2842 ^ new_n2841;
  assign new_n3034 = new_n3033 ^ new_n3032;
  assign new_n3035 = n3 & n49;
  assign new_n3036 = new_n3035 ^ new_n3032;
  assign new_n3037 = ~new_n3034 & new_n3036;
  assign new_n3038 = new_n3037 ^ new_n3035;
  assign new_n3039 = new_n3038 ^ new_n2867;
  assign new_n3040 = n2 & n49;
  assign new_n3041 = new_n3040 ^ new_n3038;
  assign new_n3042 = ~new_n3039 & new_n3041;
  assign new_n3043 = new_n3042 ^ new_n3040;
  assign new_n3044 = new_n2853 ^ new_n2852;
  assign new_n3045 = new_n3044 ^ new_n3043;
  assign new_n3046 = n1 & n49;
  assign new_n3047 = new_n3046 ^ new_n3043;
  assign new_n3048 = ~new_n3045 & new_n3047;
  assign new_n3049 = new_n3048 ^ new_n3046;
  assign new_n3050 = new_n2866 & new_n3049;
  assign new_n3051 = new_n3050 ^ new_n2865;
  assign new_n3052 = new_n3049 ^ new_n2866;
  assign new_n3053 = new_n3046 ^ new_n3045;
  assign new_n3054 = new_n3035 ^ new_n3034;
  assign new_n3055 = new_n3024 ^ new_n3023;
  assign new_n3056 = new_n3013 ^ new_n3012;
  assign new_n3057 = new_n3002 ^ new_n3001;
  assign new_n3058 = new_n2991 ^ new_n2990;
  assign new_n3059 = new_n2980 ^ new_n2979;
  assign new_n3060 = new_n2969 ^ new_n2968;
  assign new_n3061 = new_n2958 ^ new_n2957;
  assign new_n3062 = new_n2947 ^ new_n2946;
  assign new_n3063 = new_n2936 ^ new_n2935;
  assign new_n3064 = new_n2925 ^ new_n2924;
  assign new_n3065 = new_n2914 ^ new_n2913;
  assign new_n3066 = new_n2903 ^ new_n2902;
  assign new_n3067 = new_n2892 ^ new_n2891;
  assign new_n3068 = new_n2887 ^ new_n2886;
  assign new_n3069 = n32 & n49;
  assign new_n3070 = n31 & n50;
  assign new_n3071 = new_n3069 & new_n3070;
  assign new_n3072 = new_n2883 ^ new_n2882;
  assign new_n3073 = new_n3072 ^ new_n3071;
  assign new_n3074 = n30 & n50;
  assign new_n3075 = new_n3074 ^ new_n3071;
  assign new_n3076 = ~new_n3073 & new_n3075;
  assign new_n3077 = new_n3076 ^ new_n3074;
  assign new_n3078 = new_n3077 ^ new_n3068;
  assign new_n3079 = n29 & n50;
  assign new_n3080 = new_n3079 ^ new_n3077;
  assign new_n3081 = ~new_n3078 & new_n3080;
  assign new_n3082 = new_n3081 ^ new_n3079;
  assign new_n3083 = new_n3082 ^ new_n3067;
  assign new_n3084 = n28 & n50;
  assign new_n3085 = new_n3084 ^ new_n3082;
  assign new_n3086 = ~new_n3083 & new_n3085;
  assign new_n3087 = new_n3086 ^ new_n3084;
  assign new_n3088 = new_n2897 ^ new_n2896;
  assign new_n3089 = new_n3088 ^ new_n3087;
  assign new_n3090 = n27 & n50;
  assign new_n3091 = new_n3090 ^ new_n3087;
  assign new_n3092 = ~new_n3089 & new_n3091;
  assign new_n3093 = new_n3092 ^ new_n3090;
  assign new_n3094 = new_n3093 ^ new_n3066;
  assign new_n3095 = n26 & n50;
  assign new_n3096 = new_n3095 ^ new_n3093;
  assign new_n3097 = ~new_n3094 & new_n3096;
  assign new_n3098 = new_n3097 ^ new_n3095;
  assign new_n3099 = new_n2908 ^ new_n2907;
  assign new_n3100 = new_n3099 ^ new_n3098;
  assign new_n3101 = n25 & n50;
  assign new_n3102 = new_n3101 ^ new_n3098;
  assign new_n3103 = ~new_n3100 & new_n3102;
  assign new_n3104 = new_n3103 ^ new_n3101;
  assign new_n3105 = new_n3104 ^ new_n3065;
  assign new_n3106 = n24 & n50;
  assign new_n3107 = new_n3106 ^ new_n3104;
  assign new_n3108 = ~new_n3105 & new_n3107;
  assign new_n3109 = new_n3108 ^ new_n3106;
  assign new_n3110 = new_n2919 ^ new_n2918;
  assign new_n3111 = new_n3110 ^ new_n3109;
  assign new_n3112 = n23 & n50;
  assign new_n3113 = new_n3112 ^ new_n3109;
  assign new_n3114 = ~new_n3111 & new_n3113;
  assign new_n3115 = new_n3114 ^ new_n3112;
  assign new_n3116 = new_n3115 ^ new_n3064;
  assign new_n3117 = n22 & n50;
  assign new_n3118 = new_n3117 ^ new_n3115;
  assign new_n3119 = ~new_n3116 & new_n3118;
  assign new_n3120 = new_n3119 ^ new_n3117;
  assign new_n3121 = new_n2930 ^ new_n2929;
  assign new_n3122 = new_n3121 ^ new_n3120;
  assign new_n3123 = n21 & n50;
  assign new_n3124 = new_n3123 ^ new_n3120;
  assign new_n3125 = ~new_n3122 & new_n3124;
  assign new_n3126 = new_n3125 ^ new_n3123;
  assign new_n3127 = new_n3126 ^ new_n3063;
  assign new_n3128 = n20 & n50;
  assign new_n3129 = new_n3128 ^ new_n3126;
  assign new_n3130 = ~new_n3127 & new_n3129;
  assign new_n3131 = new_n3130 ^ new_n3128;
  assign new_n3132 = new_n2941 ^ new_n2940;
  assign new_n3133 = new_n3132 ^ new_n3131;
  assign new_n3134 = n19 & n50;
  assign new_n3135 = new_n3134 ^ new_n3131;
  assign new_n3136 = ~new_n3133 & new_n3135;
  assign new_n3137 = new_n3136 ^ new_n3134;
  assign new_n3138 = new_n3137 ^ new_n3062;
  assign new_n3139 = n18 & n50;
  assign new_n3140 = new_n3139 ^ new_n3137;
  assign new_n3141 = ~new_n3138 & new_n3140;
  assign new_n3142 = new_n3141 ^ new_n3139;
  assign new_n3143 = new_n2952 ^ new_n2951;
  assign new_n3144 = new_n3143 ^ new_n3142;
  assign new_n3145 = n17 & n50;
  assign new_n3146 = new_n3145 ^ new_n3142;
  assign new_n3147 = ~new_n3144 & new_n3146;
  assign new_n3148 = new_n3147 ^ new_n3145;
  assign new_n3149 = new_n3148 ^ new_n3061;
  assign new_n3150 = n16 & n50;
  assign new_n3151 = new_n3150 ^ new_n3148;
  assign new_n3152 = ~new_n3149 & new_n3151;
  assign new_n3153 = new_n3152 ^ new_n3150;
  assign new_n3154 = new_n2963 ^ new_n2962;
  assign new_n3155 = new_n3154 ^ new_n3153;
  assign new_n3156 = n15 & n50;
  assign new_n3157 = new_n3156 ^ new_n3153;
  assign new_n3158 = ~new_n3155 & new_n3157;
  assign new_n3159 = new_n3158 ^ new_n3156;
  assign new_n3160 = new_n3159 ^ new_n3060;
  assign new_n3161 = n14 & n50;
  assign new_n3162 = new_n3161 ^ new_n3159;
  assign new_n3163 = ~new_n3160 & new_n3162;
  assign new_n3164 = new_n3163 ^ new_n3161;
  assign new_n3165 = new_n2974 ^ new_n2973;
  assign new_n3166 = new_n3165 ^ new_n3164;
  assign new_n3167 = n13 & n50;
  assign new_n3168 = new_n3167 ^ new_n3164;
  assign new_n3169 = ~new_n3166 & new_n3168;
  assign new_n3170 = new_n3169 ^ new_n3167;
  assign new_n3171 = new_n3170 ^ new_n3059;
  assign new_n3172 = n12 & n50;
  assign new_n3173 = new_n3172 ^ new_n3170;
  assign new_n3174 = ~new_n3171 & new_n3173;
  assign new_n3175 = new_n3174 ^ new_n3172;
  assign new_n3176 = new_n2985 ^ new_n2984;
  assign new_n3177 = new_n3176 ^ new_n3175;
  assign new_n3178 = n11 & n50;
  assign new_n3179 = new_n3178 ^ new_n3175;
  assign new_n3180 = ~new_n3177 & new_n3179;
  assign new_n3181 = new_n3180 ^ new_n3178;
  assign new_n3182 = new_n3181 ^ new_n3058;
  assign new_n3183 = n10 & n50;
  assign new_n3184 = new_n3183 ^ new_n3181;
  assign new_n3185 = ~new_n3182 & new_n3184;
  assign new_n3186 = new_n3185 ^ new_n3183;
  assign new_n3187 = new_n2996 ^ new_n2995;
  assign new_n3188 = new_n3187 ^ new_n3186;
  assign new_n3189 = n9 & n50;
  assign new_n3190 = new_n3189 ^ new_n3186;
  assign new_n3191 = ~new_n3188 & new_n3190;
  assign new_n3192 = new_n3191 ^ new_n3189;
  assign new_n3193 = new_n3192 ^ new_n3057;
  assign new_n3194 = n8 & n50;
  assign new_n3195 = new_n3194 ^ new_n3192;
  assign new_n3196 = ~new_n3193 & new_n3195;
  assign new_n3197 = new_n3196 ^ new_n3194;
  assign new_n3198 = new_n3007 ^ new_n3006;
  assign new_n3199 = new_n3198 ^ new_n3197;
  assign new_n3200 = n7 & n50;
  assign new_n3201 = new_n3200 ^ new_n3197;
  assign new_n3202 = ~new_n3199 & new_n3201;
  assign new_n3203 = new_n3202 ^ new_n3200;
  assign new_n3204 = new_n3203 ^ new_n3056;
  assign new_n3205 = n6 & n50;
  assign new_n3206 = new_n3205 ^ new_n3203;
  assign new_n3207 = ~new_n3204 & new_n3206;
  assign new_n3208 = new_n3207 ^ new_n3205;
  assign new_n3209 = new_n3018 ^ new_n3017;
  assign new_n3210 = new_n3209 ^ new_n3208;
  assign new_n3211 = n5 & n50;
  assign new_n3212 = new_n3211 ^ new_n3208;
  assign new_n3213 = ~new_n3210 & new_n3212;
  assign new_n3214 = new_n3213 ^ new_n3211;
  assign new_n3215 = new_n3214 ^ new_n3055;
  assign new_n3216 = n4 & n50;
  assign new_n3217 = new_n3216 ^ new_n3214;
  assign new_n3218 = ~new_n3215 & new_n3217;
  assign new_n3219 = new_n3218 ^ new_n3216;
  assign new_n3220 = new_n3029 ^ new_n3028;
  assign new_n3221 = new_n3220 ^ new_n3219;
  assign new_n3222 = n3 & n50;
  assign new_n3223 = new_n3222 ^ new_n3219;
  assign new_n3224 = ~new_n3221 & new_n3223;
  assign new_n3225 = new_n3224 ^ new_n3222;
  assign new_n3226 = new_n3225 ^ new_n3054;
  assign new_n3227 = n2 & n50;
  assign new_n3228 = new_n3227 ^ new_n3225;
  assign new_n3229 = ~new_n3226 & new_n3228;
  assign new_n3230 = new_n3229 ^ new_n3227;
  assign new_n3231 = new_n3040 ^ new_n3039;
  assign new_n3232 = new_n3231 ^ new_n3230;
  assign new_n3233 = n1 & n50;
  assign new_n3234 = new_n3233 ^ new_n3230;
  assign new_n3235 = ~new_n3232 & new_n3234;
  assign new_n3236 = new_n3235 ^ new_n3233;
  assign new_n3237 = new_n3053 & new_n3236;
  assign new_n3238 = new_n3237 ^ new_n3052;
  assign new_n3239 = new_n3236 ^ new_n3053;
  assign new_n3240 = new_n3233 ^ new_n3232;
  assign new_n3241 = new_n3227 ^ new_n3226;
  assign new_n3242 = n2 & n51;
  assign new_n3243 = new_n3211 ^ new_n3210;
  assign new_n3244 = new_n3200 ^ new_n3199;
  assign new_n3245 = new_n3189 ^ new_n3188;
  assign new_n3246 = new_n3178 ^ new_n3177;
  assign new_n3247 = new_n3167 ^ new_n3166;
  assign new_n3248 = new_n3156 ^ new_n3155;
  assign new_n3249 = new_n3145 ^ new_n3144;
  assign new_n3250 = new_n3134 ^ new_n3133;
  assign new_n3251 = new_n3123 ^ new_n3122;
  assign new_n3252 = new_n3112 ^ new_n3111;
  assign new_n3253 = new_n3101 ^ new_n3100;
  assign new_n3254 = new_n3090 ^ new_n3089;
  assign new_n3255 = new_n3079 ^ new_n3078;
  assign new_n3256 = new_n3074 ^ new_n3073;
  assign new_n3257 = n32 & n50;
  assign new_n3258 = n31 & n51;
  assign new_n3259 = new_n3257 & new_n3258;
  assign new_n3260 = new_n3070 ^ new_n3069;
  assign new_n3261 = new_n3260 ^ new_n3259;
  assign new_n3262 = n30 & n51;
  assign new_n3263 = new_n3262 ^ new_n3259;
  assign new_n3264 = ~new_n3261 & new_n3263;
  assign new_n3265 = new_n3264 ^ new_n3262;
  assign new_n3266 = new_n3265 ^ new_n3256;
  assign new_n3267 = n29 & n51;
  assign new_n3268 = new_n3267 ^ new_n3265;
  assign new_n3269 = ~new_n3266 & new_n3268;
  assign new_n3270 = new_n3269 ^ new_n3267;
  assign new_n3271 = new_n3270 ^ new_n3255;
  assign new_n3272 = n28 & n51;
  assign new_n3273 = new_n3272 ^ new_n3270;
  assign new_n3274 = ~new_n3271 & new_n3273;
  assign new_n3275 = new_n3274 ^ new_n3272;
  assign new_n3276 = new_n3084 ^ new_n3083;
  assign new_n3277 = new_n3276 ^ new_n3275;
  assign new_n3278 = n27 & n51;
  assign new_n3279 = new_n3278 ^ new_n3275;
  assign new_n3280 = ~new_n3277 & new_n3279;
  assign new_n3281 = new_n3280 ^ new_n3278;
  assign new_n3282 = new_n3281 ^ new_n3254;
  assign new_n3283 = n26 & n51;
  assign new_n3284 = new_n3283 ^ new_n3281;
  assign new_n3285 = ~new_n3282 & new_n3284;
  assign new_n3286 = new_n3285 ^ new_n3283;
  assign new_n3287 = new_n3095 ^ new_n3094;
  assign new_n3288 = new_n3287 ^ new_n3286;
  assign new_n3289 = n25 & n51;
  assign new_n3290 = new_n3289 ^ new_n3286;
  assign new_n3291 = ~new_n3288 & new_n3290;
  assign new_n3292 = new_n3291 ^ new_n3289;
  assign new_n3293 = new_n3292 ^ new_n3253;
  assign new_n3294 = n24 & n51;
  assign new_n3295 = new_n3294 ^ new_n3292;
  assign new_n3296 = ~new_n3293 & new_n3295;
  assign new_n3297 = new_n3296 ^ new_n3294;
  assign new_n3298 = new_n3106 ^ new_n3105;
  assign new_n3299 = new_n3298 ^ new_n3297;
  assign new_n3300 = n23 & n51;
  assign new_n3301 = new_n3300 ^ new_n3297;
  assign new_n3302 = ~new_n3299 & new_n3301;
  assign new_n3303 = new_n3302 ^ new_n3300;
  assign new_n3304 = new_n3303 ^ new_n3252;
  assign new_n3305 = n22 & n51;
  assign new_n3306 = new_n3305 ^ new_n3303;
  assign new_n3307 = ~new_n3304 & new_n3306;
  assign new_n3308 = new_n3307 ^ new_n3305;
  assign new_n3309 = new_n3117 ^ new_n3116;
  assign new_n3310 = new_n3309 ^ new_n3308;
  assign new_n3311 = n21 & n51;
  assign new_n3312 = new_n3311 ^ new_n3308;
  assign new_n3313 = ~new_n3310 & new_n3312;
  assign new_n3314 = new_n3313 ^ new_n3311;
  assign new_n3315 = new_n3314 ^ new_n3251;
  assign new_n3316 = n20 & n51;
  assign new_n3317 = new_n3316 ^ new_n3314;
  assign new_n3318 = ~new_n3315 & new_n3317;
  assign new_n3319 = new_n3318 ^ new_n3316;
  assign new_n3320 = new_n3128 ^ new_n3127;
  assign new_n3321 = new_n3320 ^ new_n3319;
  assign new_n3322 = n19 & n51;
  assign new_n3323 = new_n3322 ^ new_n3319;
  assign new_n3324 = ~new_n3321 & new_n3323;
  assign new_n3325 = new_n3324 ^ new_n3322;
  assign new_n3326 = new_n3325 ^ new_n3250;
  assign new_n3327 = n18 & n51;
  assign new_n3328 = new_n3327 ^ new_n3325;
  assign new_n3329 = ~new_n3326 & new_n3328;
  assign new_n3330 = new_n3329 ^ new_n3327;
  assign new_n3331 = new_n3139 ^ new_n3138;
  assign new_n3332 = new_n3331 ^ new_n3330;
  assign new_n3333 = n17 & n51;
  assign new_n3334 = new_n3333 ^ new_n3330;
  assign new_n3335 = ~new_n3332 & new_n3334;
  assign new_n3336 = new_n3335 ^ new_n3333;
  assign new_n3337 = new_n3336 ^ new_n3249;
  assign new_n3338 = n16 & n51;
  assign new_n3339 = new_n3338 ^ new_n3336;
  assign new_n3340 = ~new_n3337 & new_n3339;
  assign new_n3341 = new_n3340 ^ new_n3338;
  assign new_n3342 = new_n3150 ^ new_n3149;
  assign new_n3343 = new_n3342 ^ new_n3341;
  assign new_n3344 = n15 & n51;
  assign new_n3345 = new_n3344 ^ new_n3341;
  assign new_n3346 = ~new_n3343 & new_n3345;
  assign new_n3347 = new_n3346 ^ new_n3344;
  assign new_n3348 = new_n3347 ^ new_n3248;
  assign new_n3349 = n14 & n51;
  assign new_n3350 = new_n3349 ^ new_n3347;
  assign new_n3351 = ~new_n3348 & new_n3350;
  assign new_n3352 = new_n3351 ^ new_n3349;
  assign new_n3353 = new_n3161 ^ new_n3160;
  assign new_n3354 = new_n3353 ^ new_n3352;
  assign new_n3355 = n13 & n51;
  assign new_n3356 = new_n3355 ^ new_n3352;
  assign new_n3357 = ~new_n3354 & new_n3356;
  assign new_n3358 = new_n3357 ^ new_n3355;
  assign new_n3359 = new_n3358 ^ new_n3247;
  assign new_n3360 = n12 & n51;
  assign new_n3361 = new_n3360 ^ new_n3358;
  assign new_n3362 = ~new_n3359 & new_n3361;
  assign new_n3363 = new_n3362 ^ new_n3360;
  assign new_n3364 = new_n3172 ^ new_n3171;
  assign new_n3365 = new_n3364 ^ new_n3363;
  assign new_n3366 = n11 & n51;
  assign new_n3367 = new_n3366 ^ new_n3363;
  assign new_n3368 = ~new_n3365 & new_n3367;
  assign new_n3369 = new_n3368 ^ new_n3366;
  assign new_n3370 = new_n3369 ^ new_n3246;
  assign new_n3371 = n10 & n51;
  assign new_n3372 = new_n3371 ^ new_n3369;
  assign new_n3373 = ~new_n3370 & new_n3372;
  assign new_n3374 = new_n3373 ^ new_n3371;
  assign new_n3375 = new_n3183 ^ new_n3182;
  assign new_n3376 = new_n3375 ^ new_n3374;
  assign new_n3377 = n9 & n51;
  assign new_n3378 = new_n3377 ^ new_n3374;
  assign new_n3379 = ~new_n3376 & new_n3378;
  assign new_n3380 = new_n3379 ^ new_n3377;
  assign new_n3381 = new_n3380 ^ new_n3245;
  assign new_n3382 = n8 & n51;
  assign new_n3383 = new_n3382 ^ new_n3380;
  assign new_n3384 = ~new_n3381 & new_n3383;
  assign new_n3385 = new_n3384 ^ new_n3382;
  assign new_n3386 = new_n3194 ^ new_n3193;
  assign new_n3387 = new_n3386 ^ new_n3385;
  assign new_n3388 = n7 & n51;
  assign new_n3389 = new_n3388 ^ new_n3385;
  assign new_n3390 = ~new_n3387 & new_n3389;
  assign new_n3391 = new_n3390 ^ new_n3388;
  assign new_n3392 = new_n3391 ^ new_n3244;
  assign new_n3393 = n6 & n51;
  assign new_n3394 = new_n3393 ^ new_n3391;
  assign new_n3395 = ~new_n3392 & new_n3394;
  assign new_n3396 = new_n3395 ^ new_n3393;
  assign new_n3397 = new_n3205 ^ new_n3204;
  assign new_n3398 = new_n3397 ^ new_n3396;
  assign new_n3399 = n5 & n51;
  assign new_n3400 = new_n3399 ^ new_n3396;
  assign new_n3401 = ~new_n3398 & new_n3400;
  assign new_n3402 = new_n3401 ^ new_n3399;
  assign new_n3403 = new_n3402 ^ new_n3243;
  assign new_n3404 = n4 & n51;
  assign new_n3405 = new_n3404 ^ new_n3402;
  assign new_n3406 = ~new_n3403 & new_n3405;
  assign new_n3407 = new_n3406 ^ new_n3404;
  assign new_n3408 = n3 & n51;
  assign new_n3409 = new_n3408 ^ new_n3407;
  assign new_n3410 = new_n3216 ^ new_n3215;
  assign new_n3411 = new_n3410 ^ new_n3408;
  assign new_n3412 = ~new_n3411 & new_n3409;
  assign new_n3413 = new_n3412 ^ new_n3407;
  assign new_n3414 = new_n3413 ^ new_n3242;
  assign new_n3415 = ~new_n3414 & new_n3242;
  assign new_n3416 = new_n3222 ^ new_n3221;
  assign new_n3417 = new_n3414 & new_n3416;
  assign new_n3418 = new_n3417 ^ new_n3415;
  assign new_n3419 = new_n3418 ^ new_n3241;
  assign new_n3420 = n1 & n51;
  assign new_n3421 = new_n3420 ^ new_n3418;
  assign new_n3422 = ~new_n3419 & new_n3421;
  assign new_n3423 = new_n3422 ^ new_n3420;
  assign new_n3424 = new_n3240 & new_n3423;
  assign new_n3425 = new_n3424 ^ new_n3239;
  assign new_n3426 = new_n3420 ^ new_n3419;
  assign new_n3427 = new_n3399 ^ new_n3398;
  assign new_n3428 = new_n3388 ^ new_n3387;
  assign new_n3429 = new_n3377 ^ new_n3376;
  assign new_n3430 = new_n3366 ^ new_n3365;
  assign new_n3431 = new_n3355 ^ new_n3354;
  assign new_n3432 = new_n3344 ^ new_n3343;
  assign new_n3433 = new_n3333 ^ new_n3332;
  assign new_n3434 = new_n3322 ^ new_n3321;
  assign new_n3435 = new_n3311 ^ new_n3310;
  assign new_n3436 = new_n3300 ^ new_n3299;
  assign new_n3437 = new_n3289 ^ new_n3288;
  assign new_n3438 = new_n3278 ^ new_n3277;
  assign new_n3439 = new_n3267 ^ new_n3266;
  assign new_n3440 = new_n3262 ^ new_n3261;
  assign new_n3441 = n32 & n51;
  assign new_n3442 = n31 & n52;
  assign new_n3443 = new_n3441 & new_n3442;
  assign new_n3444 = new_n3258 ^ new_n3257;
  assign new_n3445 = new_n3444 ^ new_n3443;
  assign new_n3446 = n30 & n52;
  assign new_n3447 = new_n3446 ^ new_n3443;
  assign new_n3448 = ~new_n3445 & new_n3447;
  assign new_n3449 = new_n3448 ^ new_n3446;
  assign new_n3450 = new_n3449 ^ new_n3440;
  assign new_n3451 = n29 & n52;
  assign new_n3452 = new_n3451 ^ new_n3449;
  assign new_n3453 = ~new_n3450 & new_n3452;
  assign new_n3454 = new_n3453 ^ new_n3451;
  assign new_n3455 = new_n3454 ^ new_n3439;
  assign new_n3456 = n28 & n52;
  assign new_n3457 = new_n3456 ^ new_n3454;
  assign new_n3458 = ~new_n3455 & new_n3457;
  assign new_n3459 = new_n3458 ^ new_n3456;
  assign new_n3460 = new_n3272 ^ new_n3271;
  assign new_n3461 = new_n3460 ^ new_n3459;
  assign new_n3462 = n27 & n52;
  assign new_n3463 = new_n3462 ^ new_n3459;
  assign new_n3464 = ~new_n3461 & new_n3463;
  assign new_n3465 = new_n3464 ^ new_n3462;
  assign new_n3466 = new_n3465 ^ new_n3438;
  assign new_n3467 = n26 & n52;
  assign new_n3468 = new_n3467 ^ new_n3465;
  assign new_n3469 = ~new_n3466 & new_n3468;
  assign new_n3470 = new_n3469 ^ new_n3467;
  assign new_n3471 = new_n3283 ^ new_n3282;
  assign new_n3472 = new_n3471 ^ new_n3470;
  assign new_n3473 = n25 & n52;
  assign new_n3474 = new_n3473 ^ new_n3470;
  assign new_n3475 = ~new_n3472 & new_n3474;
  assign new_n3476 = new_n3475 ^ new_n3473;
  assign new_n3477 = new_n3476 ^ new_n3437;
  assign new_n3478 = n24 & n52;
  assign new_n3479 = new_n3478 ^ new_n3476;
  assign new_n3480 = ~new_n3477 & new_n3479;
  assign new_n3481 = new_n3480 ^ new_n3478;
  assign new_n3482 = new_n3294 ^ new_n3293;
  assign new_n3483 = new_n3482 ^ new_n3481;
  assign new_n3484 = n23 & n52;
  assign new_n3485 = new_n3484 ^ new_n3481;
  assign new_n3486 = ~new_n3483 & new_n3485;
  assign new_n3487 = new_n3486 ^ new_n3484;
  assign new_n3488 = new_n3487 ^ new_n3436;
  assign new_n3489 = n22 & n52;
  assign new_n3490 = new_n3489 ^ new_n3487;
  assign new_n3491 = ~new_n3488 & new_n3490;
  assign new_n3492 = new_n3491 ^ new_n3489;
  assign new_n3493 = new_n3305 ^ new_n3304;
  assign new_n3494 = new_n3493 ^ new_n3492;
  assign new_n3495 = n21 & n52;
  assign new_n3496 = new_n3495 ^ new_n3492;
  assign new_n3497 = ~new_n3494 & new_n3496;
  assign new_n3498 = new_n3497 ^ new_n3495;
  assign new_n3499 = new_n3498 ^ new_n3435;
  assign new_n3500 = n20 & n52;
  assign new_n3501 = new_n3500 ^ new_n3498;
  assign new_n3502 = ~new_n3499 & new_n3501;
  assign new_n3503 = new_n3502 ^ new_n3500;
  assign new_n3504 = new_n3316 ^ new_n3315;
  assign new_n3505 = new_n3504 ^ new_n3503;
  assign new_n3506 = n19 & n52;
  assign new_n3507 = new_n3506 ^ new_n3503;
  assign new_n3508 = ~new_n3505 & new_n3507;
  assign new_n3509 = new_n3508 ^ new_n3506;
  assign new_n3510 = new_n3509 ^ new_n3434;
  assign new_n3511 = n18 & n52;
  assign new_n3512 = new_n3511 ^ new_n3509;
  assign new_n3513 = ~new_n3510 & new_n3512;
  assign new_n3514 = new_n3513 ^ new_n3511;
  assign new_n3515 = new_n3327 ^ new_n3326;
  assign new_n3516 = new_n3515 ^ new_n3514;
  assign new_n3517 = n17 & n52;
  assign new_n3518 = new_n3517 ^ new_n3514;
  assign new_n3519 = ~new_n3516 & new_n3518;
  assign new_n3520 = new_n3519 ^ new_n3517;
  assign new_n3521 = new_n3520 ^ new_n3433;
  assign new_n3522 = n16 & n52;
  assign new_n3523 = new_n3522 ^ new_n3520;
  assign new_n3524 = ~new_n3521 & new_n3523;
  assign new_n3525 = new_n3524 ^ new_n3522;
  assign new_n3526 = new_n3338 ^ new_n3337;
  assign new_n3527 = new_n3526 ^ new_n3525;
  assign new_n3528 = n15 & n52;
  assign new_n3529 = new_n3528 ^ new_n3525;
  assign new_n3530 = ~new_n3527 & new_n3529;
  assign new_n3531 = new_n3530 ^ new_n3528;
  assign new_n3532 = new_n3531 ^ new_n3432;
  assign new_n3533 = n14 & n52;
  assign new_n3534 = new_n3533 ^ new_n3531;
  assign new_n3535 = ~new_n3532 & new_n3534;
  assign new_n3536 = new_n3535 ^ new_n3533;
  assign new_n3537 = new_n3349 ^ new_n3348;
  assign new_n3538 = new_n3537 ^ new_n3536;
  assign new_n3539 = n13 & n52;
  assign new_n3540 = new_n3539 ^ new_n3536;
  assign new_n3541 = ~new_n3538 & new_n3540;
  assign new_n3542 = new_n3541 ^ new_n3539;
  assign new_n3543 = new_n3542 ^ new_n3431;
  assign new_n3544 = n12 & n52;
  assign new_n3545 = new_n3544 ^ new_n3542;
  assign new_n3546 = ~new_n3543 & new_n3545;
  assign new_n3547 = new_n3546 ^ new_n3544;
  assign new_n3548 = new_n3360 ^ new_n3359;
  assign new_n3549 = new_n3548 ^ new_n3547;
  assign new_n3550 = n11 & n52;
  assign new_n3551 = new_n3550 ^ new_n3547;
  assign new_n3552 = ~new_n3549 & new_n3551;
  assign new_n3553 = new_n3552 ^ new_n3550;
  assign new_n3554 = new_n3553 ^ new_n3430;
  assign new_n3555 = n10 & n52;
  assign new_n3556 = new_n3555 ^ new_n3553;
  assign new_n3557 = ~new_n3554 & new_n3556;
  assign new_n3558 = new_n3557 ^ new_n3555;
  assign new_n3559 = new_n3371 ^ new_n3370;
  assign new_n3560 = new_n3559 ^ new_n3558;
  assign new_n3561 = n9 & n52;
  assign new_n3562 = new_n3561 ^ new_n3558;
  assign new_n3563 = ~new_n3560 & new_n3562;
  assign new_n3564 = new_n3563 ^ new_n3561;
  assign new_n3565 = new_n3564 ^ new_n3429;
  assign new_n3566 = n8 & n52;
  assign new_n3567 = new_n3566 ^ new_n3564;
  assign new_n3568 = ~new_n3565 & new_n3567;
  assign new_n3569 = new_n3568 ^ new_n3566;
  assign new_n3570 = new_n3382 ^ new_n3381;
  assign new_n3571 = new_n3570 ^ new_n3569;
  assign new_n3572 = n7 & n52;
  assign new_n3573 = new_n3572 ^ new_n3569;
  assign new_n3574 = ~new_n3571 & new_n3573;
  assign new_n3575 = new_n3574 ^ new_n3572;
  assign new_n3576 = new_n3575 ^ new_n3428;
  assign new_n3577 = n6 & n52;
  assign new_n3578 = new_n3577 ^ new_n3575;
  assign new_n3579 = ~new_n3576 & new_n3578;
  assign new_n3580 = new_n3579 ^ new_n3577;
  assign new_n3581 = new_n3393 ^ new_n3392;
  assign new_n3582 = new_n3581 ^ new_n3580;
  assign new_n3583 = n5 & n52;
  assign new_n3584 = new_n3583 ^ new_n3580;
  assign new_n3585 = ~new_n3582 & new_n3584;
  assign new_n3586 = new_n3585 ^ new_n3583;
  assign new_n3587 = new_n3586 ^ new_n3427;
  assign new_n3588 = n4 & n52;
  assign new_n3589 = new_n3588 ^ new_n3586;
  assign new_n3590 = ~new_n3587 & new_n3589;
  assign new_n3591 = new_n3590 ^ new_n3588;
  assign new_n3592 = new_n3404 ^ new_n3403;
  assign new_n3593 = new_n3592 ^ new_n3591;
  assign new_n3594 = n3 & n52;
  assign new_n3595 = new_n3594 ^ new_n3591;
  assign new_n3596 = ~new_n3593 & new_n3595;
  assign new_n3597 = new_n3596 ^ new_n3594;
  assign new_n3598 = n2 & n52;
  assign new_n3599 = new_n3598 ^ new_n3597;
  assign new_n3600 = new_n3410 ^ new_n3409;
  assign new_n3601 = new_n3600 ^ new_n3598;
  assign new_n3602 = ~new_n3601 & new_n3599;
  assign new_n3603 = new_n3602 ^ new_n3597;
  assign new_n3604 = n1 & n52;
  assign new_n3605 = new_n3604 ^ new_n3603;
  assign new_n3606 = ~new_n3605 & new_n3603;
  assign new_n3607 = new_n3416 ^ new_n3414;
  assign new_n3608 = new_n3605 & new_n3607;
  assign new_n3609 = new_n3608 ^ new_n3606;
  assign new_n3610 = new_n3426 & new_n3609;
  assign new_n3611 = new_n3423 ^ new_n3240;
  assign new_n3612 = new_n3610 & new_n3611;
  assign new_n3613 = new_n3611 ^ new_n3610;
  assign new_n3614 = new_n3613 ^ new_n3612;
  assign new_n3615 = new_n3607 ^ new_n3605;
  assign new_n3616 = new_n3594 ^ new_n3593;
  assign new_n3617 = new_n3583 ^ new_n3582;
  assign new_n3618 = new_n3572 ^ new_n3571;
  assign new_n3619 = new_n3561 ^ new_n3560;
  assign new_n3620 = new_n3550 ^ new_n3549;
  assign new_n3621 = new_n3539 ^ new_n3538;
  assign new_n3622 = new_n3528 ^ new_n3527;
  assign new_n3623 = new_n3517 ^ new_n3516;
  assign new_n3624 = new_n3506 ^ new_n3505;
  assign new_n3625 = new_n3495 ^ new_n3494;
  assign new_n3626 = new_n3484 ^ new_n3483;
  assign new_n3627 = new_n3473 ^ new_n3472;
  assign new_n3628 = new_n3462 ^ new_n3461;
  assign new_n3629 = new_n3451 ^ new_n3450;
  assign new_n3630 = new_n3446 ^ new_n3445;
  assign new_n3631 = n32 & n52;
  assign new_n3632 = n31 & n53;
  assign new_n3633 = new_n3631 & new_n3632;
  assign new_n3634 = new_n3442 ^ new_n3441;
  assign new_n3635 = new_n3634 ^ new_n3633;
  assign new_n3636 = n30 & n53;
  assign new_n3637 = new_n3636 ^ new_n3633;
  assign new_n3638 = ~new_n3635 & new_n3637;
  assign new_n3639 = new_n3638 ^ new_n3636;
  assign new_n3640 = new_n3639 ^ new_n3630;
  assign new_n3641 = n29 & n53;
  assign new_n3642 = new_n3641 ^ new_n3639;
  assign new_n3643 = ~new_n3640 & new_n3642;
  assign new_n3644 = new_n3643 ^ new_n3641;
  assign new_n3645 = new_n3644 ^ new_n3629;
  assign new_n3646 = n28 & n53;
  assign new_n3647 = new_n3646 ^ new_n3644;
  assign new_n3648 = ~new_n3645 & new_n3647;
  assign new_n3649 = new_n3648 ^ new_n3646;
  assign new_n3650 = new_n3456 ^ new_n3455;
  assign new_n3651 = new_n3650 ^ new_n3649;
  assign new_n3652 = n27 & n53;
  assign new_n3653 = new_n3652 ^ new_n3649;
  assign new_n3654 = ~new_n3651 & new_n3653;
  assign new_n3655 = new_n3654 ^ new_n3652;
  assign new_n3656 = new_n3655 ^ new_n3628;
  assign new_n3657 = n26 & n53;
  assign new_n3658 = new_n3657 ^ new_n3655;
  assign new_n3659 = ~new_n3656 & new_n3658;
  assign new_n3660 = new_n3659 ^ new_n3657;
  assign new_n3661 = new_n3467 ^ new_n3466;
  assign new_n3662 = new_n3661 ^ new_n3660;
  assign new_n3663 = n25 & n53;
  assign new_n3664 = new_n3663 ^ new_n3660;
  assign new_n3665 = ~new_n3662 & new_n3664;
  assign new_n3666 = new_n3665 ^ new_n3663;
  assign new_n3667 = new_n3666 ^ new_n3627;
  assign new_n3668 = n24 & n53;
  assign new_n3669 = new_n3668 ^ new_n3666;
  assign new_n3670 = ~new_n3667 & new_n3669;
  assign new_n3671 = new_n3670 ^ new_n3668;
  assign new_n3672 = new_n3478 ^ new_n3477;
  assign new_n3673 = new_n3672 ^ new_n3671;
  assign new_n3674 = n23 & n53;
  assign new_n3675 = new_n3674 ^ new_n3671;
  assign new_n3676 = ~new_n3673 & new_n3675;
  assign new_n3677 = new_n3676 ^ new_n3674;
  assign new_n3678 = new_n3677 ^ new_n3626;
  assign new_n3679 = n22 & n53;
  assign new_n3680 = new_n3679 ^ new_n3677;
  assign new_n3681 = ~new_n3678 & new_n3680;
  assign new_n3682 = new_n3681 ^ new_n3679;
  assign new_n3683 = new_n3489 ^ new_n3488;
  assign new_n3684 = new_n3683 ^ new_n3682;
  assign new_n3685 = n21 & n53;
  assign new_n3686 = new_n3685 ^ new_n3682;
  assign new_n3687 = ~new_n3684 & new_n3686;
  assign new_n3688 = new_n3687 ^ new_n3685;
  assign new_n3689 = new_n3688 ^ new_n3625;
  assign new_n3690 = n20 & n53;
  assign new_n3691 = new_n3690 ^ new_n3688;
  assign new_n3692 = ~new_n3689 & new_n3691;
  assign new_n3693 = new_n3692 ^ new_n3690;
  assign new_n3694 = new_n3500 ^ new_n3499;
  assign new_n3695 = new_n3694 ^ new_n3693;
  assign new_n3696 = n19 & n53;
  assign new_n3697 = new_n3696 ^ new_n3693;
  assign new_n3698 = ~new_n3695 & new_n3697;
  assign new_n3699 = new_n3698 ^ new_n3696;
  assign new_n3700 = new_n3699 ^ new_n3624;
  assign new_n3701 = n18 & n53;
  assign new_n3702 = new_n3701 ^ new_n3699;
  assign new_n3703 = ~new_n3700 & new_n3702;
  assign new_n3704 = new_n3703 ^ new_n3701;
  assign new_n3705 = new_n3511 ^ new_n3510;
  assign new_n3706 = new_n3705 ^ new_n3704;
  assign new_n3707 = n17 & n53;
  assign new_n3708 = new_n3707 ^ new_n3704;
  assign new_n3709 = ~new_n3706 & new_n3708;
  assign new_n3710 = new_n3709 ^ new_n3707;
  assign new_n3711 = new_n3710 ^ new_n3623;
  assign new_n3712 = n16 & n53;
  assign new_n3713 = new_n3712 ^ new_n3710;
  assign new_n3714 = ~new_n3711 & new_n3713;
  assign new_n3715 = new_n3714 ^ new_n3712;
  assign new_n3716 = new_n3522 ^ new_n3521;
  assign new_n3717 = new_n3716 ^ new_n3715;
  assign new_n3718 = n15 & n53;
  assign new_n3719 = new_n3718 ^ new_n3715;
  assign new_n3720 = ~new_n3717 & new_n3719;
  assign new_n3721 = new_n3720 ^ new_n3718;
  assign new_n3722 = new_n3721 ^ new_n3622;
  assign new_n3723 = n14 & n53;
  assign new_n3724 = new_n3723 ^ new_n3721;
  assign new_n3725 = ~new_n3722 & new_n3724;
  assign new_n3726 = new_n3725 ^ new_n3723;
  assign new_n3727 = new_n3533 ^ new_n3532;
  assign new_n3728 = new_n3727 ^ new_n3726;
  assign new_n3729 = n13 & n53;
  assign new_n3730 = new_n3729 ^ new_n3726;
  assign new_n3731 = ~new_n3728 & new_n3730;
  assign new_n3732 = new_n3731 ^ new_n3729;
  assign new_n3733 = new_n3732 ^ new_n3621;
  assign new_n3734 = n12 & n53;
  assign new_n3735 = new_n3734 ^ new_n3732;
  assign new_n3736 = ~new_n3733 & new_n3735;
  assign new_n3737 = new_n3736 ^ new_n3734;
  assign new_n3738 = new_n3544 ^ new_n3543;
  assign new_n3739 = new_n3738 ^ new_n3737;
  assign new_n3740 = n11 & n53;
  assign new_n3741 = new_n3740 ^ new_n3737;
  assign new_n3742 = ~new_n3739 & new_n3741;
  assign new_n3743 = new_n3742 ^ new_n3740;
  assign new_n3744 = new_n3743 ^ new_n3620;
  assign new_n3745 = n10 & n53;
  assign new_n3746 = new_n3745 ^ new_n3743;
  assign new_n3747 = ~new_n3744 & new_n3746;
  assign new_n3748 = new_n3747 ^ new_n3745;
  assign new_n3749 = new_n3555 ^ new_n3554;
  assign new_n3750 = new_n3749 ^ new_n3748;
  assign new_n3751 = n9 & n53;
  assign new_n3752 = new_n3751 ^ new_n3748;
  assign new_n3753 = ~new_n3750 & new_n3752;
  assign new_n3754 = new_n3753 ^ new_n3751;
  assign new_n3755 = new_n3754 ^ new_n3619;
  assign new_n3756 = n8 & n53;
  assign new_n3757 = new_n3756 ^ new_n3754;
  assign new_n3758 = ~new_n3755 & new_n3757;
  assign new_n3759 = new_n3758 ^ new_n3756;
  assign new_n3760 = new_n3566 ^ new_n3565;
  assign new_n3761 = new_n3760 ^ new_n3759;
  assign new_n3762 = n7 & n53;
  assign new_n3763 = new_n3762 ^ new_n3759;
  assign new_n3764 = ~new_n3761 & new_n3763;
  assign new_n3765 = new_n3764 ^ new_n3762;
  assign new_n3766 = new_n3765 ^ new_n3618;
  assign new_n3767 = n6 & n53;
  assign new_n3768 = new_n3767 ^ new_n3765;
  assign new_n3769 = ~new_n3766 & new_n3768;
  assign new_n3770 = new_n3769 ^ new_n3767;
  assign new_n3771 = new_n3577 ^ new_n3576;
  assign new_n3772 = new_n3771 ^ new_n3770;
  assign new_n3773 = n5 & n53;
  assign new_n3774 = new_n3773 ^ new_n3770;
  assign new_n3775 = ~new_n3772 & new_n3774;
  assign new_n3776 = new_n3775 ^ new_n3773;
  assign new_n3777 = new_n3776 ^ new_n3617;
  assign new_n3778 = n4 & n53;
  assign new_n3779 = new_n3778 ^ new_n3776;
  assign new_n3780 = ~new_n3777 & new_n3779;
  assign new_n3781 = new_n3780 ^ new_n3778;
  assign new_n3782 = new_n3588 ^ new_n3587;
  assign new_n3783 = new_n3782 ^ new_n3781;
  assign new_n3784 = n3 & n53;
  assign new_n3785 = new_n3784 ^ new_n3781;
  assign new_n3786 = ~new_n3783 & new_n3785;
  assign new_n3787 = new_n3786 ^ new_n3784;
  assign new_n3788 = new_n3787 ^ new_n3616;
  assign new_n3789 = n2 & n53;
  assign new_n3790 = new_n3789 ^ new_n3787;
  assign new_n3791 = ~new_n3788 & new_n3790;
  assign new_n3792 = new_n3791 ^ new_n3789;
  assign new_n3793 = new_n3600 ^ new_n3599;
  assign new_n3794 = new_n3793 ^ new_n3792;
  assign new_n3795 = n1 & n53;
  assign new_n3796 = new_n3795 ^ new_n3792;
  assign new_n3797 = ~new_n3794 & new_n3796;
  assign new_n3798 = new_n3797 ^ new_n3795;
  assign new_n3799 = new_n3615 & new_n3798;
  assign new_n3800 = new_n3609 ^ new_n3426;
  assign new_n3801 = ~new_n3799 & ~new_n3800;
  assign new_n3802 = new_n3784 ^ new_n3783;
  assign new_n3803 = new_n3773 ^ new_n3772;
  assign new_n3804 = new_n3762 ^ new_n3761;
  assign new_n3805 = new_n3751 ^ new_n3750;
  assign new_n3806 = new_n3740 ^ new_n3739;
  assign new_n3807 = new_n3729 ^ new_n3728;
  assign new_n3808 = new_n3718 ^ new_n3717;
  assign new_n3809 = new_n3707 ^ new_n3706;
  assign new_n3810 = new_n3696 ^ new_n3695;
  assign new_n3811 = new_n3685 ^ new_n3684;
  assign new_n3812 = new_n3674 ^ new_n3673;
  assign new_n3813 = new_n3663 ^ new_n3662;
  assign new_n3814 = new_n3652 ^ new_n3651;
  assign new_n3815 = new_n3641 ^ new_n3640;
  assign new_n3816 = new_n3636 ^ new_n3635;
  assign new_n3817 = n32 & n53;
  assign new_n3818 = n31 & n54;
  assign new_n3819 = new_n3817 & new_n3818;
  assign new_n3820 = new_n3632 ^ new_n3631;
  assign new_n3821 = new_n3820 ^ new_n3819;
  assign new_n3822 = n30 & n54;
  assign new_n3823 = new_n3822 ^ new_n3819;
  assign new_n3824 = ~new_n3821 & new_n3823;
  assign new_n3825 = new_n3824 ^ new_n3822;
  assign new_n3826 = new_n3825 ^ new_n3816;
  assign new_n3827 = n29 & n54;
  assign new_n3828 = new_n3827 ^ new_n3825;
  assign new_n3829 = ~new_n3826 & new_n3828;
  assign new_n3830 = new_n3829 ^ new_n3827;
  assign new_n3831 = new_n3830 ^ new_n3815;
  assign new_n3832 = n28 & n54;
  assign new_n3833 = new_n3832 ^ new_n3830;
  assign new_n3834 = ~new_n3831 & new_n3833;
  assign new_n3835 = new_n3834 ^ new_n3832;
  assign new_n3836 = new_n3646 ^ new_n3645;
  assign new_n3837 = new_n3836 ^ new_n3835;
  assign new_n3838 = n27 & n54;
  assign new_n3839 = new_n3838 ^ new_n3835;
  assign new_n3840 = ~new_n3837 & new_n3839;
  assign new_n3841 = new_n3840 ^ new_n3838;
  assign new_n3842 = new_n3841 ^ new_n3814;
  assign new_n3843 = n26 & n54;
  assign new_n3844 = new_n3843 ^ new_n3841;
  assign new_n3845 = ~new_n3842 & new_n3844;
  assign new_n3846 = new_n3845 ^ new_n3843;
  assign new_n3847 = new_n3657 ^ new_n3656;
  assign new_n3848 = new_n3847 ^ new_n3846;
  assign new_n3849 = n25 & n54;
  assign new_n3850 = new_n3849 ^ new_n3846;
  assign new_n3851 = ~new_n3848 & new_n3850;
  assign new_n3852 = new_n3851 ^ new_n3849;
  assign new_n3853 = new_n3852 ^ new_n3813;
  assign new_n3854 = n24 & n54;
  assign new_n3855 = new_n3854 ^ new_n3852;
  assign new_n3856 = ~new_n3853 & new_n3855;
  assign new_n3857 = new_n3856 ^ new_n3854;
  assign new_n3858 = new_n3668 ^ new_n3667;
  assign new_n3859 = new_n3858 ^ new_n3857;
  assign new_n3860 = n23 & n54;
  assign new_n3861 = new_n3860 ^ new_n3857;
  assign new_n3862 = ~new_n3859 & new_n3861;
  assign new_n3863 = new_n3862 ^ new_n3860;
  assign new_n3864 = new_n3863 ^ new_n3812;
  assign new_n3865 = n22 & n54;
  assign new_n3866 = new_n3865 ^ new_n3863;
  assign new_n3867 = ~new_n3864 & new_n3866;
  assign new_n3868 = new_n3867 ^ new_n3865;
  assign new_n3869 = new_n3679 ^ new_n3678;
  assign new_n3870 = new_n3869 ^ new_n3868;
  assign new_n3871 = n21 & n54;
  assign new_n3872 = new_n3871 ^ new_n3868;
  assign new_n3873 = ~new_n3870 & new_n3872;
  assign new_n3874 = new_n3873 ^ new_n3871;
  assign new_n3875 = new_n3874 ^ new_n3811;
  assign new_n3876 = n20 & n54;
  assign new_n3877 = new_n3876 ^ new_n3874;
  assign new_n3878 = ~new_n3875 & new_n3877;
  assign new_n3879 = new_n3878 ^ new_n3876;
  assign new_n3880 = new_n3690 ^ new_n3689;
  assign new_n3881 = new_n3880 ^ new_n3879;
  assign new_n3882 = n19 & n54;
  assign new_n3883 = new_n3882 ^ new_n3879;
  assign new_n3884 = ~new_n3881 & new_n3883;
  assign new_n3885 = new_n3884 ^ new_n3882;
  assign new_n3886 = new_n3885 ^ new_n3810;
  assign new_n3887 = n18 & n54;
  assign new_n3888 = new_n3887 ^ new_n3885;
  assign new_n3889 = ~new_n3886 & new_n3888;
  assign new_n3890 = new_n3889 ^ new_n3887;
  assign new_n3891 = new_n3701 ^ new_n3700;
  assign new_n3892 = new_n3891 ^ new_n3890;
  assign new_n3893 = n17 & n54;
  assign new_n3894 = new_n3893 ^ new_n3890;
  assign new_n3895 = ~new_n3892 & new_n3894;
  assign new_n3896 = new_n3895 ^ new_n3893;
  assign new_n3897 = new_n3896 ^ new_n3809;
  assign new_n3898 = n16 & n54;
  assign new_n3899 = new_n3898 ^ new_n3896;
  assign new_n3900 = ~new_n3897 & new_n3899;
  assign new_n3901 = new_n3900 ^ new_n3898;
  assign new_n3902 = new_n3712 ^ new_n3711;
  assign new_n3903 = new_n3902 ^ new_n3901;
  assign new_n3904 = n15 & n54;
  assign new_n3905 = new_n3904 ^ new_n3901;
  assign new_n3906 = ~new_n3903 & new_n3905;
  assign new_n3907 = new_n3906 ^ new_n3904;
  assign new_n3908 = new_n3907 ^ new_n3808;
  assign new_n3909 = n14 & n54;
  assign new_n3910 = new_n3909 ^ new_n3907;
  assign new_n3911 = ~new_n3908 & new_n3910;
  assign new_n3912 = new_n3911 ^ new_n3909;
  assign new_n3913 = new_n3723 ^ new_n3722;
  assign new_n3914 = new_n3913 ^ new_n3912;
  assign new_n3915 = n13 & n54;
  assign new_n3916 = new_n3915 ^ new_n3912;
  assign new_n3917 = ~new_n3914 & new_n3916;
  assign new_n3918 = new_n3917 ^ new_n3915;
  assign new_n3919 = new_n3918 ^ new_n3807;
  assign new_n3920 = n12 & n54;
  assign new_n3921 = new_n3920 ^ new_n3918;
  assign new_n3922 = ~new_n3919 & new_n3921;
  assign new_n3923 = new_n3922 ^ new_n3920;
  assign new_n3924 = new_n3734 ^ new_n3733;
  assign new_n3925 = new_n3924 ^ new_n3923;
  assign new_n3926 = n11 & n54;
  assign new_n3927 = new_n3926 ^ new_n3923;
  assign new_n3928 = ~new_n3925 & new_n3927;
  assign new_n3929 = new_n3928 ^ new_n3926;
  assign new_n3930 = new_n3929 ^ new_n3806;
  assign new_n3931 = n10 & n54;
  assign new_n3932 = new_n3931 ^ new_n3929;
  assign new_n3933 = ~new_n3930 & new_n3932;
  assign new_n3934 = new_n3933 ^ new_n3931;
  assign new_n3935 = new_n3745 ^ new_n3744;
  assign new_n3936 = new_n3935 ^ new_n3934;
  assign new_n3937 = n9 & n54;
  assign new_n3938 = new_n3937 ^ new_n3934;
  assign new_n3939 = ~new_n3936 & new_n3938;
  assign new_n3940 = new_n3939 ^ new_n3937;
  assign new_n3941 = new_n3940 ^ new_n3805;
  assign new_n3942 = n8 & n54;
  assign new_n3943 = new_n3942 ^ new_n3940;
  assign new_n3944 = ~new_n3941 & new_n3943;
  assign new_n3945 = new_n3944 ^ new_n3942;
  assign new_n3946 = new_n3756 ^ new_n3755;
  assign new_n3947 = new_n3946 ^ new_n3945;
  assign new_n3948 = n7 & n54;
  assign new_n3949 = new_n3948 ^ new_n3945;
  assign new_n3950 = ~new_n3947 & new_n3949;
  assign new_n3951 = new_n3950 ^ new_n3948;
  assign new_n3952 = new_n3951 ^ new_n3804;
  assign new_n3953 = n6 & n54;
  assign new_n3954 = new_n3953 ^ new_n3951;
  assign new_n3955 = ~new_n3952 & new_n3954;
  assign new_n3956 = new_n3955 ^ new_n3953;
  assign new_n3957 = new_n3767 ^ new_n3766;
  assign new_n3958 = new_n3957 ^ new_n3956;
  assign new_n3959 = n5 & n54;
  assign new_n3960 = new_n3959 ^ new_n3956;
  assign new_n3961 = ~new_n3958 & new_n3960;
  assign new_n3962 = new_n3961 ^ new_n3959;
  assign new_n3963 = new_n3962 ^ new_n3803;
  assign new_n3964 = n4 & n54;
  assign new_n3965 = new_n3964 ^ new_n3962;
  assign new_n3966 = ~new_n3963 & new_n3965;
  assign new_n3967 = new_n3966 ^ new_n3964;
  assign new_n3968 = new_n3778 ^ new_n3777;
  assign new_n3969 = new_n3968 ^ new_n3967;
  assign new_n3970 = n3 & n54;
  assign new_n3971 = new_n3970 ^ new_n3967;
  assign new_n3972 = ~new_n3969 & new_n3971;
  assign new_n3973 = new_n3972 ^ new_n3970;
  assign new_n3974 = new_n3973 ^ new_n3802;
  assign new_n3975 = n2 & n54;
  assign new_n3976 = new_n3975 ^ new_n3973;
  assign new_n3977 = ~new_n3974 & new_n3976;
  assign new_n3978 = new_n3977 ^ new_n3975;
  assign new_n3979 = new_n3789 ^ new_n3788;
  assign new_n3980 = new_n3979 ^ new_n3978;
  assign new_n3981 = n1 & n54;
  assign new_n3982 = new_n3981 ^ new_n3978;
  assign new_n3983 = ~new_n3980 & new_n3982;
  assign new_n3984 = new_n3983 ^ new_n3981;
  assign new_n3985 = new_n3795 ^ new_n3794;
  assign new_n3986 = new_n3984 & new_n3985;
  assign new_n3987 = new_n3798 ^ new_n3615;
  assign new_n3988 = new_n3986 & new_n3987;
  assign new_n3989 = new_n3987 ^ new_n3986;
  assign new_n3990 = new_n3989 ^ new_n3988;
  assign new_n3991 = ~new_n3801 & new_n3990;
  assign new_n3992 = new_n3981 ^ new_n3980;
  assign new_n3993 = new_n3975 ^ new_n3974;
  assign new_n3994 = n2 & n55;
  assign new_n3995 = new_n3959 ^ new_n3958;
  assign new_n3996 = new_n3948 ^ new_n3947;
  assign new_n3997 = new_n3937 ^ new_n3936;
  assign new_n3998 = new_n3926 ^ new_n3925;
  assign new_n3999 = new_n3915 ^ new_n3914;
  assign new_n4000 = new_n3904 ^ new_n3903;
  assign new_n4001 = new_n3893 ^ new_n3892;
  assign new_n4002 = new_n3882 ^ new_n3881;
  assign new_n4003 = new_n3871 ^ new_n3870;
  assign new_n4004 = new_n3860 ^ new_n3859;
  assign new_n4005 = new_n3849 ^ new_n3848;
  assign new_n4006 = new_n3838 ^ new_n3837;
  assign new_n4007 = new_n3827 ^ new_n3826;
  assign new_n4008 = new_n3822 ^ new_n3821;
  assign new_n4009 = n32 & n54;
  assign new_n4010 = n31 & n55;
  assign new_n4011 = new_n4009 & new_n4010;
  assign new_n4012 = new_n3818 ^ new_n3817;
  assign new_n4013 = new_n4012 ^ new_n4011;
  assign new_n4014 = n30 & n55;
  assign new_n4015 = new_n4014 ^ new_n4011;
  assign new_n4016 = ~new_n4013 & new_n4015;
  assign new_n4017 = new_n4016 ^ new_n4014;
  assign new_n4018 = new_n4017 ^ new_n4008;
  assign new_n4019 = n29 & n55;
  assign new_n4020 = new_n4019 ^ new_n4017;
  assign new_n4021 = ~new_n4018 & new_n4020;
  assign new_n4022 = new_n4021 ^ new_n4019;
  assign new_n4023 = new_n4022 ^ new_n4007;
  assign new_n4024 = n28 & n55;
  assign new_n4025 = new_n4024 ^ new_n4022;
  assign new_n4026 = ~new_n4023 & new_n4025;
  assign new_n4027 = new_n4026 ^ new_n4024;
  assign new_n4028 = new_n3832 ^ new_n3831;
  assign new_n4029 = new_n4028 ^ new_n4027;
  assign new_n4030 = n27 & n55;
  assign new_n4031 = new_n4030 ^ new_n4027;
  assign new_n4032 = ~new_n4029 & new_n4031;
  assign new_n4033 = new_n4032 ^ new_n4030;
  assign new_n4034 = new_n4033 ^ new_n4006;
  assign new_n4035 = n26 & n55;
  assign new_n4036 = new_n4035 ^ new_n4033;
  assign new_n4037 = ~new_n4034 & new_n4036;
  assign new_n4038 = new_n4037 ^ new_n4035;
  assign new_n4039 = new_n3843 ^ new_n3842;
  assign new_n4040 = new_n4039 ^ new_n4038;
  assign new_n4041 = n25 & n55;
  assign new_n4042 = new_n4041 ^ new_n4038;
  assign new_n4043 = ~new_n4040 & new_n4042;
  assign new_n4044 = new_n4043 ^ new_n4041;
  assign new_n4045 = new_n4044 ^ new_n4005;
  assign new_n4046 = n24 & n55;
  assign new_n4047 = new_n4046 ^ new_n4044;
  assign new_n4048 = ~new_n4045 & new_n4047;
  assign new_n4049 = new_n4048 ^ new_n4046;
  assign new_n4050 = new_n3854 ^ new_n3853;
  assign new_n4051 = new_n4050 ^ new_n4049;
  assign new_n4052 = n23 & n55;
  assign new_n4053 = new_n4052 ^ new_n4049;
  assign new_n4054 = ~new_n4051 & new_n4053;
  assign new_n4055 = new_n4054 ^ new_n4052;
  assign new_n4056 = new_n4055 ^ new_n4004;
  assign new_n4057 = n22 & n55;
  assign new_n4058 = new_n4057 ^ new_n4055;
  assign new_n4059 = ~new_n4056 & new_n4058;
  assign new_n4060 = new_n4059 ^ new_n4057;
  assign new_n4061 = new_n3865 ^ new_n3864;
  assign new_n4062 = new_n4061 ^ new_n4060;
  assign new_n4063 = n21 & n55;
  assign new_n4064 = new_n4063 ^ new_n4060;
  assign new_n4065 = ~new_n4062 & new_n4064;
  assign new_n4066 = new_n4065 ^ new_n4063;
  assign new_n4067 = new_n4066 ^ new_n4003;
  assign new_n4068 = n20 & n55;
  assign new_n4069 = new_n4068 ^ new_n4066;
  assign new_n4070 = ~new_n4067 & new_n4069;
  assign new_n4071 = new_n4070 ^ new_n4068;
  assign new_n4072 = new_n3876 ^ new_n3875;
  assign new_n4073 = new_n4072 ^ new_n4071;
  assign new_n4074 = n19 & n55;
  assign new_n4075 = new_n4074 ^ new_n4071;
  assign new_n4076 = ~new_n4073 & new_n4075;
  assign new_n4077 = new_n4076 ^ new_n4074;
  assign new_n4078 = new_n4077 ^ new_n4002;
  assign new_n4079 = n18 & n55;
  assign new_n4080 = new_n4079 ^ new_n4077;
  assign new_n4081 = ~new_n4078 & new_n4080;
  assign new_n4082 = new_n4081 ^ new_n4079;
  assign new_n4083 = new_n3887 ^ new_n3886;
  assign new_n4084 = new_n4083 ^ new_n4082;
  assign new_n4085 = n17 & n55;
  assign new_n4086 = new_n4085 ^ new_n4082;
  assign new_n4087 = ~new_n4084 & new_n4086;
  assign new_n4088 = new_n4087 ^ new_n4085;
  assign new_n4089 = new_n4088 ^ new_n4001;
  assign new_n4090 = n16 & n55;
  assign new_n4091 = new_n4090 ^ new_n4088;
  assign new_n4092 = ~new_n4089 & new_n4091;
  assign new_n4093 = new_n4092 ^ new_n4090;
  assign new_n4094 = new_n3898 ^ new_n3897;
  assign new_n4095 = new_n4094 ^ new_n4093;
  assign new_n4096 = n15 & n55;
  assign new_n4097 = new_n4096 ^ new_n4093;
  assign new_n4098 = ~new_n4095 & new_n4097;
  assign new_n4099 = new_n4098 ^ new_n4096;
  assign new_n4100 = new_n4099 ^ new_n4000;
  assign new_n4101 = n14 & n55;
  assign new_n4102 = new_n4101 ^ new_n4099;
  assign new_n4103 = ~new_n4100 & new_n4102;
  assign new_n4104 = new_n4103 ^ new_n4101;
  assign new_n4105 = new_n3909 ^ new_n3908;
  assign new_n4106 = new_n4105 ^ new_n4104;
  assign new_n4107 = n13 & n55;
  assign new_n4108 = new_n4107 ^ new_n4104;
  assign new_n4109 = ~new_n4106 & new_n4108;
  assign new_n4110 = new_n4109 ^ new_n4107;
  assign new_n4111 = new_n4110 ^ new_n3999;
  assign new_n4112 = n12 & n55;
  assign new_n4113 = new_n4112 ^ new_n4110;
  assign new_n4114 = ~new_n4111 & new_n4113;
  assign new_n4115 = new_n4114 ^ new_n4112;
  assign new_n4116 = new_n3920 ^ new_n3919;
  assign new_n4117 = new_n4116 ^ new_n4115;
  assign new_n4118 = n11 & n55;
  assign new_n4119 = new_n4118 ^ new_n4115;
  assign new_n4120 = ~new_n4117 & new_n4119;
  assign new_n4121 = new_n4120 ^ new_n4118;
  assign new_n4122 = new_n4121 ^ new_n3998;
  assign new_n4123 = n10 & n55;
  assign new_n4124 = new_n4123 ^ new_n4121;
  assign new_n4125 = ~new_n4122 & new_n4124;
  assign new_n4126 = new_n4125 ^ new_n4123;
  assign new_n4127 = new_n3931 ^ new_n3930;
  assign new_n4128 = new_n4127 ^ new_n4126;
  assign new_n4129 = n9 & n55;
  assign new_n4130 = new_n4129 ^ new_n4126;
  assign new_n4131 = ~new_n4128 & new_n4130;
  assign new_n4132 = new_n4131 ^ new_n4129;
  assign new_n4133 = new_n4132 ^ new_n3997;
  assign new_n4134 = n8 & n55;
  assign new_n4135 = new_n4134 ^ new_n4132;
  assign new_n4136 = ~new_n4133 & new_n4135;
  assign new_n4137 = new_n4136 ^ new_n4134;
  assign new_n4138 = new_n3942 ^ new_n3941;
  assign new_n4139 = new_n4138 ^ new_n4137;
  assign new_n4140 = n7 & n55;
  assign new_n4141 = new_n4140 ^ new_n4137;
  assign new_n4142 = ~new_n4139 & new_n4141;
  assign new_n4143 = new_n4142 ^ new_n4140;
  assign new_n4144 = new_n4143 ^ new_n3996;
  assign new_n4145 = n6 & n55;
  assign new_n4146 = new_n4145 ^ new_n4143;
  assign new_n4147 = ~new_n4144 & new_n4146;
  assign new_n4148 = new_n4147 ^ new_n4145;
  assign new_n4149 = new_n3953 ^ new_n3952;
  assign new_n4150 = new_n4149 ^ new_n4148;
  assign new_n4151 = n5 & n55;
  assign new_n4152 = new_n4151 ^ new_n4148;
  assign new_n4153 = ~new_n4150 & new_n4152;
  assign new_n4154 = new_n4153 ^ new_n4151;
  assign new_n4155 = new_n4154 ^ new_n3995;
  assign new_n4156 = n4 & n55;
  assign new_n4157 = new_n4156 ^ new_n4154;
  assign new_n4158 = ~new_n4155 & new_n4157;
  assign new_n4159 = new_n4158 ^ new_n4156;
  assign new_n4160 = n3 & n55;
  assign new_n4161 = new_n4160 ^ new_n4159;
  assign new_n4162 = new_n3964 ^ new_n3963;
  assign new_n4163 = new_n4162 ^ new_n4160;
  assign new_n4164 = ~new_n4163 & new_n4161;
  assign new_n4165 = new_n4164 ^ new_n4159;
  assign new_n4166 = new_n4165 ^ new_n3994;
  assign new_n4167 = ~new_n4166 & new_n3994;
  assign new_n4168 = new_n3970 ^ new_n3969;
  assign new_n4169 = new_n4166 & new_n4168;
  assign new_n4170 = new_n4169 ^ new_n4167;
  assign new_n4171 = new_n4170 ^ new_n3993;
  assign new_n4172 = n1 & n55;
  assign new_n4173 = new_n4172 ^ new_n4170;
  assign new_n4174 = ~new_n4171 & new_n4173;
  assign new_n4175 = new_n4174 ^ new_n4172;
  assign new_n4176 = new_n3992 & new_n4175;
  assign new_n4177 = new_n3985 ^ new_n3984;
  assign new_n4178 = new_n4177 ^ new_n4176;
  assign new_n4179 = ~new_n4176 & ~new_n4177;
  assign new_n4180 = new_n4179 ^ new_n4178;
  assign new_n4181 = new_n4180 ^ new_n3988;
  assign new_n4182 = ~new_n4181 & new_n3991;
  assign new_n4183 = new_n3800 ^ new_n3799;
  assign new_n4184 = new_n4183 ^ new_n3801;
  assign new_n4185 = new_n4184 ^ new_n4182;
  assign new_n4186 = ~new_n4185 & new_n3614;
  assign new_n4187 = new_n4186 ^ new_n3612;
  assign new_n4188 = new_n4172 ^ new_n4171;
  assign new_n4189 = new_n4151 ^ new_n4150;
  assign new_n4190 = new_n4140 ^ new_n4139;
  assign new_n4191 = new_n4129 ^ new_n4128;
  assign new_n4192 = new_n4118 ^ new_n4117;
  assign new_n4193 = new_n4107 ^ new_n4106;
  assign new_n4194 = new_n4096 ^ new_n4095;
  assign new_n4195 = new_n4085 ^ new_n4084;
  assign new_n4196 = new_n4074 ^ new_n4073;
  assign new_n4197 = new_n4063 ^ new_n4062;
  assign new_n4198 = new_n4052 ^ new_n4051;
  assign new_n4199 = new_n4041 ^ new_n4040;
  assign new_n4200 = new_n4030 ^ new_n4029;
  assign new_n4201 = new_n4019 ^ new_n4018;
  assign new_n4202 = new_n4014 ^ new_n4013;
  assign new_n4203 = n32 & n55;
  assign new_n4204 = n31 & n56;
  assign new_n4205 = new_n4203 & new_n4204;
  assign new_n4206 = new_n4010 ^ new_n4009;
  assign new_n4207 = new_n4206 ^ new_n4205;
  assign new_n4208 = n30 & n56;
  assign new_n4209 = new_n4208 ^ new_n4205;
  assign new_n4210 = ~new_n4207 & new_n4209;
  assign new_n4211 = new_n4210 ^ new_n4208;
  assign new_n4212 = new_n4211 ^ new_n4202;
  assign new_n4213 = n29 & n56;
  assign new_n4214 = new_n4213 ^ new_n4211;
  assign new_n4215 = ~new_n4212 & new_n4214;
  assign new_n4216 = new_n4215 ^ new_n4213;
  assign new_n4217 = new_n4216 ^ new_n4201;
  assign new_n4218 = n28 & n56;
  assign new_n4219 = new_n4218 ^ new_n4216;
  assign new_n4220 = ~new_n4217 & new_n4219;
  assign new_n4221 = new_n4220 ^ new_n4218;
  assign new_n4222 = new_n4024 ^ new_n4023;
  assign new_n4223 = new_n4222 ^ new_n4221;
  assign new_n4224 = n27 & n56;
  assign new_n4225 = new_n4224 ^ new_n4221;
  assign new_n4226 = ~new_n4223 & new_n4225;
  assign new_n4227 = new_n4226 ^ new_n4224;
  assign new_n4228 = new_n4227 ^ new_n4200;
  assign new_n4229 = n26 & n56;
  assign new_n4230 = new_n4229 ^ new_n4227;
  assign new_n4231 = ~new_n4228 & new_n4230;
  assign new_n4232 = new_n4231 ^ new_n4229;
  assign new_n4233 = new_n4035 ^ new_n4034;
  assign new_n4234 = new_n4233 ^ new_n4232;
  assign new_n4235 = n25 & n56;
  assign new_n4236 = new_n4235 ^ new_n4232;
  assign new_n4237 = ~new_n4234 & new_n4236;
  assign new_n4238 = new_n4237 ^ new_n4235;
  assign new_n4239 = new_n4238 ^ new_n4199;
  assign new_n4240 = n24 & n56;
  assign new_n4241 = new_n4240 ^ new_n4238;
  assign new_n4242 = ~new_n4239 & new_n4241;
  assign new_n4243 = new_n4242 ^ new_n4240;
  assign new_n4244 = new_n4046 ^ new_n4045;
  assign new_n4245 = new_n4244 ^ new_n4243;
  assign new_n4246 = n23 & n56;
  assign new_n4247 = new_n4246 ^ new_n4243;
  assign new_n4248 = ~new_n4245 & new_n4247;
  assign new_n4249 = new_n4248 ^ new_n4246;
  assign new_n4250 = new_n4249 ^ new_n4198;
  assign new_n4251 = n22 & n56;
  assign new_n4252 = new_n4251 ^ new_n4249;
  assign new_n4253 = ~new_n4250 & new_n4252;
  assign new_n4254 = new_n4253 ^ new_n4251;
  assign new_n4255 = new_n4057 ^ new_n4056;
  assign new_n4256 = new_n4255 ^ new_n4254;
  assign new_n4257 = n21 & n56;
  assign new_n4258 = new_n4257 ^ new_n4254;
  assign new_n4259 = ~new_n4256 & new_n4258;
  assign new_n4260 = new_n4259 ^ new_n4257;
  assign new_n4261 = new_n4260 ^ new_n4197;
  assign new_n4262 = n20 & n56;
  assign new_n4263 = new_n4262 ^ new_n4260;
  assign new_n4264 = ~new_n4261 & new_n4263;
  assign new_n4265 = new_n4264 ^ new_n4262;
  assign new_n4266 = new_n4068 ^ new_n4067;
  assign new_n4267 = new_n4266 ^ new_n4265;
  assign new_n4268 = n19 & n56;
  assign new_n4269 = new_n4268 ^ new_n4265;
  assign new_n4270 = ~new_n4267 & new_n4269;
  assign new_n4271 = new_n4270 ^ new_n4268;
  assign new_n4272 = new_n4271 ^ new_n4196;
  assign new_n4273 = n18 & n56;
  assign new_n4274 = new_n4273 ^ new_n4271;
  assign new_n4275 = ~new_n4272 & new_n4274;
  assign new_n4276 = new_n4275 ^ new_n4273;
  assign new_n4277 = new_n4079 ^ new_n4078;
  assign new_n4278 = new_n4277 ^ new_n4276;
  assign new_n4279 = n17 & n56;
  assign new_n4280 = new_n4279 ^ new_n4276;
  assign new_n4281 = ~new_n4278 & new_n4280;
  assign new_n4282 = new_n4281 ^ new_n4279;
  assign new_n4283 = new_n4282 ^ new_n4195;
  assign new_n4284 = n16 & n56;
  assign new_n4285 = new_n4284 ^ new_n4282;
  assign new_n4286 = ~new_n4283 & new_n4285;
  assign new_n4287 = new_n4286 ^ new_n4284;
  assign new_n4288 = new_n4090 ^ new_n4089;
  assign new_n4289 = new_n4288 ^ new_n4287;
  assign new_n4290 = n15 & n56;
  assign new_n4291 = new_n4290 ^ new_n4287;
  assign new_n4292 = ~new_n4289 & new_n4291;
  assign new_n4293 = new_n4292 ^ new_n4290;
  assign new_n4294 = new_n4293 ^ new_n4194;
  assign new_n4295 = n14 & n56;
  assign new_n4296 = new_n4295 ^ new_n4293;
  assign new_n4297 = ~new_n4294 & new_n4296;
  assign new_n4298 = new_n4297 ^ new_n4295;
  assign new_n4299 = new_n4101 ^ new_n4100;
  assign new_n4300 = new_n4299 ^ new_n4298;
  assign new_n4301 = n13 & n56;
  assign new_n4302 = new_n4301 ^ new_n4298;
  assign new_n4303 = ~new_n4300 & new_n4302;
  assign new_n4304 = new_n4303 ^ new_n4301;
  assign new_n4305 = new_n4304 ^ new_n4193;
  assign new_n4306 = n12 & n56;
  assign new_n4307 = new_n4306 ^ new_n4304;
  assign new_n4308 = ~new_n4305 & new_n4307;
  assign new_n4309 = new_n4308 ^ new_n4306;
  assign new_n4310 = new_n4112 ^ new_n4111;
  assign new_n4311 = new_n4310 ^ new_n4309;
  assign new_n4312 = n11 & n56;
  assign new_n4313 = new_n4312 ^ new_n4309;
  assign new_n4314 = ~new_n4311 & new_n4313;
  assign new_n4315 = new_n4314 ^ new_n4312;
  assign new_n4316 = new_n4315 ^ new_n4192;
  assign new_n4317 = n10 & n56;
  assign new_n4318 = new_n4317 ^ new_n4315;
  assign new_n4319 = ~new_n4316 & new_n4318;
  assign new_n4320 = new_n4319 ^ new_n4317;
  assign new_n4321 = new_n4123 ^ new_n4122;
  assign new_n4322 = new_n4321 ^ new_n4320;
  assign new_n4323 = n9 & n56;
  assign new_n4324 = new_n4323 ^ new_n4320;
  assign new_n4325 = ~new_n4322 & new_n4324;
  assign new_n4326 = new_n4325 ^ new_n4323;
  assign new_n4327 = new_n4326 ^ new_n4191;
  assign new_n4328 = n8 & n56;
  assign new_n4329 = new_n4328 ^ new_n4326;
  assign new_n4330 = ~new_n4327 & new_n4329;
  assign new_n4331 = new_n4330 ^ new_n4328;
  assign new_n4332 = new_n4134 ^ new_n4133;
  assign new_n4333 = new_n4332 ^ new_n4331;
  assign new_n4334 = n7 & n56;
  assign new_n4335 = new_n4334 ^ new_n4331;
  assign new_n4336 = ~new_n4333 & new_n4335;
  assign new_n4337 = new_n4336 ^ new_n4334;
  assign new_n4338 = new_n4337 ^ new_n4190;
  assign new_n4339 = n6 & n56;
  assign new_n4340 = new_n4339 ^ new_n4337;
  assign new_n4341 = ~new_n4338 & new_n4340;
  assign new_n4342 = new_n4341 ^ new_n4339;
  assign new_n4343 = new_n4145 ^ new_n4144;
  assign new_n4344 = new_n4343 ^ new_n4342;
  assign new_n4345 = n5 & n56;
  assign new_n4346 = new_n4345 ^ new_n4342;
  assign new_n4347 = ~new_n4344 & new_n4346;
  assign new_n4348 = new_n4347 ^ new_n4345;
  assign new_n4349 = new_n4348 ^ new_n4189;
  assign new_n4350 = n4 & n56;
  assign new_n4351 = new_n4350 ^ new_n4348;
  assign new_n4352 = ~new_n4349 & new_n4351;
  assign new_n4353 = new_n4352 ^ new_n4350;
  assign new_n4354 = new_n4156 ^ new_n4155;
  assign new_n4355 = new_n4354 ^ new_n4353;
  assign new_n4356 = n3 & n56;
  assign new_n4357 = new_n4356 ^ new_n4353;
  assign new_n4358 = ~new_n4355 & new_n4357;
  assign new_n4359 = new_n4358 ^ new_n4356;
  assign new_n4360 = n2 & n56;
  assign new_n4361 = new_n4360 ^ new_n4359;
  assign new_n4362 = new_n4162 ^ new_n4161;
  assign new_n4363 = new_n4362 ^ new_n4360;
  assign new_n4364 = ~new_n4363 & new_n4361;
  assign new_n4365 = new_n4364 ^ new_n4359;
  assign new_n4366 = n1 & n56;
  assign new_n4367 = new_n4366 ^ new_n4365;
  assign new_n4368 = ~new_n4367 & new_n4365;
  assign new_n4369 = new_n4168 ^ new_n4166;
  assign new_n4370 = new_n4367 & new_n4369;
  assign new_n4371 = new_n4370 ^ new_n4368;
  assign new_n4372 = new_n4188 & new_n4371;
  assign new_n4373 = new_n4175 ^ new_n3992;
  assign new_n4374 = new_n4372 & new_n4373;
  assign new_n4375 = new_n4373 ^ new_n4372;
  assign new_n4376 = new_n4375 ^ new_n4374;
  assign new_n4377 = new_n4369 ^ new_n4367;
  assign new_n4378 = new_n4356 ^ new_n4355;
  assign new_n4379 = new_n4345 ^ new_n4344;
  assign new_n4380 = new_n4334 ^ new_n4333;
  assign new_n4381 = new_n4323 ^ new_n4322;
  assign new_n4382 = new_n4312 ^ new_n4311;
  assign new_n4383 = new_n4301 ^ new_n4300;
  assign new_n4384 = new_n4290 ^ new_n4289;
  assign new_n4385 = new_n4279 ^ new_n4278;
  assign new_n4386 = new_n4268 ^ new_n4267;
  assign new_n4387 = new_n4257 ^ new_n4256;
  assign new_n4388 = new_n4246 ^ new_n4245;
  assign new_n4389 = new_n4235 ^ new_n4234;
  assign new_n4390 = new_n4224 ^ new_n4223;
  assign new_n4391 = new_n4213 ^ new_n4212;
  assign new_n4392 = new_n4208 ^ new_n4207;
  assign new_n4393 = n32 & n56;
  assign new_n4394 = n31 & n57;
  assign new_n4395 = new_n4393 & new_n4394;
  assign new_n4396 = new_n4204 ^ new_n4203;
  assign new_n4397 = new_n4396 ^ new_n4395;
  assign new_n4398 = n30 & n57;
  assign new_n4399 = new_n4398 ^ new_n4395;
  assign new_n4400 = ~new_n4397 & new_n4399;
  assign new_n4401 = new_n4400 ^ new_n4398;
  assign new_n4402 = new_n4401 ^ new_n4392;
  assign new_n4403 = n29 & n57;
  assign new_n4404 = new_n4403 ^ new_n4401;
  assign new_n4405 = ~new_n4402 & new_n4404;
  assign new_n4406 = new_n4405 ^ new_n4403;
  assign new_n4407 = new_n4406 ^ new_n4391;
  assign new_n4408 = n28 & n57;
  assign new_n4409 = new_n4408 ^ new_n4406;
  assign new_n4410 = ~new_n4407 & new_n4409;
  assign new_n4411 = new_n4410 ^ new_n4408;
  assign new_n4412 = new_n4218 ^ new_n4217;
  assign new_n4413 = new_n4412 ^ new_n4411;
  assign new_n4414 = n27 & n57;
  assign new_n4415 = new_n4414 ^ new_n4411;
  assign new_n4416 = ~new_n4413 & new_n4415;
  assign new_n4417 = new_n4416 ^ new_n4414;
  assign new_n4418 = new_n4417 ^ new_n4390;
  assign new_n4419 = n26 & n57;
  assign new_n4420 = new_n4419 ^ new_n4417;
  assign new_n4421 = ~new_n4418 & new_n4420;
  assign new_n4422 = new_n4421 ^ new_n4419;
  assign new_n4423 = new_n4229 ^ new_n4228;
  assign new_n4424 = new_n4423 ^ new_n4422;
  assign new_n4425 = n25 & n57;
  assign new_n4426 = new_n4425 ^ new_n4422;
  assign new_n4427 = ~new_n4424 & new_n4426;
  assign new_n4428 = new_n4427 ^ new_n4425;
  assign new_n4429 = new_n4428 ^ new_n4389;
  assign new_n4430 = n24 & n57;
  assign new_n4431 = new_n4430 ^ new_n4428;
  assign new_n4432 = ~new_n4429 & new_n4431;
  assign new_n4433 = new_n4432 ^ new_n4430;
  assign new_n4434 = new_n4240 ^ new_n4239;
  assign new_n4435 = new_n4434 ^ new_n4433;
  assign new_n4436 = n23 & n57;
  assign new_n4437 = new_n4436 ^ new_n4433;
  assign new_n4438 = ~new_n4435 & new_n4437;
  assign new_n4439 = new_n4438 ^ new_n4436;
  assign new_n4440 = new_n4439 ^ new_n4388;
  assign new_n4441 = n22 & n57;
  assign new_n4442 = new_n4441 ^ new_n4439;
  assign new_n4443 = ~new_n4440 & new_n4442;
  assign new_n4444 = new_n4443 ^ new_n4441;
  assign new_n4445 = new_n4251 ^ new_n4250;
  assign new_n4446 = new_n4445 ^ new_n4444;
  assign new_n4447 = n21 & n57;
  assign new_n4448 = new_n4447 ^ new_n4444;
  assign new_n4449 = ~new_n4446 & new_n4448;
  assign new_n4450 = new_n4449 ^ new_n4447;
  assign new_n4451 = new_n4450 ^ new_n4387;
  assign new_n4452 = n20 & n57;
  assign new_n4453 = new_n4452 ^ new_n4450;
  assign new_n4454 = ~new_n4451 & new_n4453;
  assign new_n4455 = new_n4454 ^ new_n4452;
  assign new_n4456 = new_n4262 ^ new_n4261;
  assign new_n4457 = new_n4456 ^ new_n4455;
  assign new_n4458 = n19 & n57;
  assign new_n4459 = new_n4458 ^ new_n4455;
  assign new_n4460 = ~new_n4457 & new_n4459;
  assign new_n4461 = new_n4460 ^ new_n4458;
  assign new_n4462 = new_n4461 ^ new_n4386;
  assign new_n4463 = n18 & n57;
  assign new_n4464 = new_n4463 ^ new_n4461;
  assign new_n4465 = ~new_n4462 & new_n4464;
  assign new_n4466 = new_n4465 ^ new_n4463;
  assign new_n4467 = new_n4273 ^ new_n4272;
  assign new_n4468 = new_n4467 ^ new_n4466;
  assign new_n4469 = n17 & n57;
  assign new_n4470 = new_n4469 ^ new_n4466;
  assign new_n4471 = ~new_n4468 & new_n4470;
  assign new_n4472 = new_n4471 ^ new_n4469;
  assign new_n4473 = new_n4472 ^ new_n4385;
  assign new_n4474 = n16 & n57;
  assign new_n4475 = new_n4474 ^ new_n4472;
  assign new_n4476 = ~new_n4473 & new_n4475;
  assign new_n4477 = new_n4476 ^ new_n4474;
  assign new_n4478 = new_n4284 ^ new_n4283;
  assign new_n4479 = new_n4478 ^ new_n4477;
  assign new_n4480 = n15 & n57;
  assign new_n4481 = new_n4480 ^ new_n4477;
  assign new_n4482 = ~new_n4479 & new_n4481;
  assign new_n4483 = new_n4482 ^ new_n4480;
  assign new_n4484 = new_n4483 ^ new_n4384;
  assign new_n4485 = n14 & n57;
  assign new_n4486 = new_n4485 ^ new_n4483;
  assign new_n4487 = ~new_n4484 & new_n4486;
  assign new_n4488 = new_n4487 ^ new_n4485;
  assign new_n4489 = new_n4295 ^ new_n4294;
  assign new_n4490 = new_n4489 ^ new_n4488;
  assign new_n4491 = n13 & n57;
  assign new_n4492 = new_n4491 ^ new_n4488;
  assign new_n4493 = ~new_n4490 & new_n4492;
  assign new_n4494 = new_n4493 ^ new_n4491;
  assign new_n4495 = new_n4494 ^ new_n4383;
  assign new_n4496 = n12 & n57;
  assign new_n4497 = new_n4496 ^ new_n4494;
  assign new_n4498 = ~new_n4495 & new_n4497;
  assign new_n4499 = new_n4498 ^ new_n4496;
  assign new_n4500 = new_n4306 ^ new_n4305;
  assign new_n4501 = new_n4500 ^ new_n4499;
  assign new_n4502 = n11 & n57;
  assign new_n4503 = new_n4502 ^ new_n4499;
  assign new_n4504 = ~new_n4501 & new_n4503;
  assign new_n4505 = new_n4504 ^ new_n4502;
  assign new_n4506 = new_n4505 ^ new_n4382;
  assign new_n4507 = n10 & n57;
  assign new_n4508 = new_n4507 ^ new_n4505;
  assign new_n4509 = ~new_n4506 & new_n4508;
  assign new_n4510 = new_n4509 ^ new_n4507;
  assign new_n4511 = new_n4317 ^ new_n4316;
  assign new_n4512 = new_n4511 ^ new_n4510;
  assign new_n4513 = n9 & n57;
  assign new_n4514 = new_n4513 ^ new_n4510;
  assign new_n4515 = ~new_n4512 & new_n4514;
  assign new_n4516 = new_n4515 ^ new_n4513;
  assign new_n4517 = new_n4516 ^ new_n4381;
  assign new_n4518 = n8 & n57;
  assign new_n4519 = new_n4518 ^ new_n4516;
  assign new_n4520 = ~new_n4517 & new_n4519;
  assign new_n4521 = new_n4520 ^ new_n4518;
  assign new_n4522 = new_n4328 ^ new_n4327;
  assign new_n4523 = new_n4522 ^ new_n4521;
  assign new_n4524 = n7 & n57;
  assign new_n4525 = new_n4524 ^ new_n4521;
  assign new_n4526 = ~new_n4523 & new_n4525;
  assign new_n4527 = new_n4526 ^ new_n4524;
  assign new_n4528 = new_n4527 ^ new_n4380;
  assign new_n4529 = n6 & n57;
  assign new_n4530 = new_n4529 ^ new_n4527;
  assign new_n4531 = ~new_n4528 & new_n4530;
  assign new_n4532 = new_n4531 ^ new_n4529;
  assign new_n4533 = new_n4339 ^ new_n4338;
  assign new_n4534 = new_n4533 ^ new_n4532;
  assign new_n4535 = n5 & n57;
  assign new_n4536 = new_n4535 ^ new_n4532;
  assign new_n4537 = ~new_n4534 & new_n4536;
  assign new_n4538 = new_n4537 ^ new_n4535;
  assign new_n4539 = new_n4538 ^ new_n4379;
  assign new_n4540 = n4 & n57;
  assign new_n4541 = new_n4540 ^ new_n4538;
  assign new_n4542 = ~new_n4539 & new_n4541;
  assign new_n4543 = new_n4542 ^ new_n4540;
  assign new_n4544 = new_n4350 ^ new_n4349;
  assign new_n4545 = new_n4544 ^ new_n4543;
  assign new_n4546 = n3 & n57;
  assign new_n4547 = new_n4546 ^ new_n4543;
  assign new_n4548 = ~new_n4545 & new_n4547;
  assign new_n4549 = new_n4548 ^ new_n4546;
  assign new_n4550 = new_n4549 ^ new_n4378;
  assign new_n4551 = n2 & n57;
  assign new_n4552 = new_n4551 ^ new_n4549;
  assign new_n4553 = ~new_n4550 & new_n4552;
  assign new_n4554 = new_n4553 ^ new_n4551;
  assign new_n4555 = new_n4362 ^ new_n4361;
  assign new_n4556 = new_n4555 ^ new_n4554;
  assign new_n4557 = n1 & n57;
  assign new_n4558 = new_n4557 ^ new_n4554;
  assign new_n4559 = ~new_n4556 & new_n4558;
  assign new_n4560 = new_n4559 ^ new_n4557;
  assign new_n4561 = new_n4377 & new_n4560;
  assign new_n4562 = new_n4371 ^ new_n4188;
  assign new_n4563 = ~new_n4561 & ~new_n4562;
  assign new_n4564 = new_n4546 ^ new_n4545;
  assign new_n4565 = new_n4535 ^ new_n4534;
  assign new_n4566 = new_n4524 ^ new_n4523;
  assign new_n4567 = new_n4513 ^ new_n4512;
  assign new_n4568 = new_n4502 ^ new_n4501;
  assign new_n4569 = new_n4491 ^ new_n4490;
  assign new_n4570 = new_n4480 ^ new_n4479;
  assign new_n4571 = new_n4469 ^ new_n4468;
  assign new_n4572 = new_n4458 ^ new_n4457;
  assign new_n4573 = new_n4447 ^ new_n4446;
  assign new_n4574 = new_n4436 ^ new_n4435;
  assign new_n4575 = new_n4425 ^ new_n4424;
  assign new_n4576 = new_n4414 ^ new_n4413;
  assign new_n4577 = new_n4403 ^ new_n4402;
  assign new_n4578 = new_n4398 ^ new_n4397;
  assign new_n4579 = n32 & n57;
  assign new_n4580 = n31 & n58;
  assign new_n4581 = new_n4579 & new_n4580;
  assign new_n4582 = new_n4394 ^ new_n4393;
  assign new_n4583 = new_n4582 ^ new_n4581;
  assign new_n4584 = n30 & n58;
  assign new_n4585 = new_n4584 ^ new_n4581;
  assign new_n4586 = ~new_n4583 & new_n4585;
  assign new_n4587 = new_n4586 ^ new_n4584;
  assign new_n4588 = new_n4587 ^ new_n4578;
  assign new_n4589 = n29 & n58;
  assign new_n4590 = new_n4589 ^ new_n4587;
  assign new_n4591 = ~new_n4588 & new_n4590;
  assign new_n4592 = new_n4591 ^ new_n4589;
  assign new_n4593 = new_n4592 ^ new_n4577;
  assign new_n4594 = n28 & n58;
  assign new_n4595 = new_n4594 ^ new_n4592;
  assign new_n4596 = ~new_n4593 & new_n4595;
  assign new_n4597 = new_n4596 ^ new_n4594;
  assign new_n4598 = new_n4408 ^ new_n4407;
  assign new_n4599 = new_n4598 ^ new_n4597;
  assign new_n4600 = n27 & n58;
  assign new_n4601 = new_n4600 ^ new_n4597;
  assign new_n4602 = ~new_n4599 & new_n4601;
  assign new_n4603 = new_n4602 ^ new_n4600;
  assign new_n4604 = new_n4603 ^ new_n4576;
  assign new_n4605 = n26 & n58;
  assign new_n4606 = new_n4605 ^ new_n4603;
  assign new_n4607 = ~new_n4604 & new_n4606;
  assign new_n4608 = new_n4607 ^ new_n4605;
  assign new_n4609 = new_n4419 ^ new_n4418;
  assign new_n4610 = new_n4609 ^ new_n4608;
  assign new_n4611 = n25 & n58;
  assign new_n4612 = new_n4611 ^ new_n4608;
  assign new_n4613 = ~new_n4610 & new_n4612;
  assign new_n4614 = new_n4613 ^ new_n4611;
  assign new_n4615 = new_n4614 ^ new_n4575;
  assign new_n4616 = n24 & n58;
  assign new_n4617 = new_n4616 ^ new_n4614;
  assign new_n4618 = ~new_n4615 & new_n4617;
  assign new_n4619 = new_n4618 ^ new_n4616;
  assign new_n4620 = new_n4430 ^ new_n4429;
  assign new_n4621 = new_n4620 ^ new_n4619;
  assign new_n4622 = n23 & n58;
  assign new_n4623 = new_n4622 ^ new_n4619;
  assign new_n4624 = ~new_n4621 & new_n4623;
  assign new_n4625 = new_n4624 ^ new_n4622;
  assign new_n4626 = new_n4625 ^ new_n4574;
  assign new_n4627 = n22 & n58;
  assign new_n4628 = new_n4627 ^ new_n4625;
  assign new_n4629 = ~new_n4626 & new_n4628;
  assign new_n4630 = new_n4629 ^ new_n4627;
  assign new_n4631 = new_n4441 ^ new_n4440;
  assign new_n4632 = new_n4631 ^ new_n4630;
  assign new_n4633 = n21 & n58;
  assign new_n4634 = new_n4633 ^ new_n4630;
  assign new_n4635 = ~new_n4632 & new_n4634;
  assign new_n4636 = new_n4635 ^ new_n4633;
  assign new_n4637 = new_n4636 ^ new_n4573;
  assign new_n4638 = n20 & n58;
  assign new_n4639 = new_n4638 ^ new_n4636;
  assign new_n4640 = ~new_n4637 & new_n4639;
  assign new_n4641 = new_n4640 ^ new_n4638;
  assign new_n4642 = new_n4452 ^ new_n4451;
  assign new_n4643 = new_n4642 ^ new_n4641;
  assign new_n4644 = n19 & n58;
  assign new_n4645 = new_n4644 ^ new_n4641;
  assign new_n4646 = ~new_n4643 & new_n4645;
  assign new_n4647 = new_n4646 ^ new_n4644;
  assign new_n4648 = new_n4647 ^ new_n4572;
  assign new_n4649 = n18 & n58;
  assign new_n4650 = new_n4649 ^ new_n4647;
  assign new_n4651 = ~new_n4648 & new_n4650;
  assign new_n4652 = new_n4651 ^ new_n4649;
  assign new_n4653 = new_n4463 ^ new_n4462;
  assign new_n4654 = new_n4653 ^ new_n4652;
  assign new_n4655 = n17 & n58;
  assign new_n4656 = new_n4655 ^ new_n4652;
  assign new_n4657 = ~new_n4654 & new_n4656;
  assign new_n4658 = new_n4657 ^ new_n4655;
  assign new_n4659 = new_n4658 ^ new_n4571;
  assign new_n4660 = n16 & n58;
  assign new_n4661 = new_n4660 ^ new_n4658;
  assign new_n4662 = ~new_n4659 & new_n4661;
  assign new_n4663 = new_n4662 ^ new_n4660;
  assign new_n4664 = new_n4474 ^ new_n4473;
  assign new_n4665 = new_n4664 ^ new_n4663;
  assign new_n4666 = n15 & n58;
  assign new_n4667 = new_n4666 ^ new_n4663;
  assign new_n4668 = ~new_n4665 & new_n4667;
  assign new_n4669 = new_n4668 ^ new_n4666;
  assign new_n4670 = new_n4669 ^ new_n4570;
  assign new_n4671 = n14 & n58;
  assign new_n4672 = new_n4671 ^ new_n4669;
  assign new_n4673 = ~new_n4670 & new_n4672;
  assign new_n4674 = new_n4673 ^ new_n4671;
  assign new_n4675 = new_n4485 ^ new_n4484;
  assign new_n4676 = new_n4675 ^ new_n4674;
  assign new_n4677 = n13 & n58;
  assign new_n4678 = new_n4677 ^ new_n4674;
  assign new_n4679 = ~new_n4676 & new_n4678;
  assign new_n4680 = new_n4679 ^ new_n4677;
  assign new_n4681 = new_n4680 ^ new_n4569;
  assign new_n4682 = n12 & n58;
  assign new_n4683 = new_n4682 ^ new_n4680;
  assign new_n4684 = ~new_n4681 & new_n4683;
  assign new_n4685 = new_n4684 ^ new_n4682;
  assign new_n4686 = new_n4496 ^ new_n4495;
  assign new_n4687 = new_n4686 ^ new_n4685;
  assign new_n4688 = n11 & n58;
  assign new_n4689 = new_n4688 ^ new_n4685;
  assign new_n4690 = ~new_n4687 & new_n4689;
  assign new_n4691 = new_n4690 ^ new_n4688;
  assign new_n4692 = new_n4691 ^ new_n4568;
  assign new_n4693 = n10 & n58;
  assign new_n4694 = new_n4693 ^ new_n4691;
  assign new_n4695 = ~new_n4692 & new_n4694;
  assign new_n4696 = new_n4695 ^ new_n4693;
  assign new_n4697 = new_n4507 ^ new_n4506;
  assign new_n4698 = new_n4697 ^ new_n4696;
  assign new_n4699 = n9 & n58;
  assign new_n4700 = new_n4699 ^ new_n4696;
  assign new_n4701 = ~new_n4698 & new_n4700;
  assign new_n4702 = new_n4701 ^ new_n4699;
  assign new_n4703 = new_n4702 ^ new_n4567;
  assign new_n4704 = n8 & n58;
  assign new_n4705 = new_n4704 ^ new_n4702;
  assign new_n4706 = ~new_n4703 & new_n4705;
  assign new_n4707 = new_n4706 ^ new_n4704;
  assign new_n4708 = new_n4518 ^ new_n4517;
  assign new_n4709 = new_n4708 ^ new_n4707;
  assign new_n4710 = n7 & n58;
  assign new_n4711 = new_n4710 ^ new_n4707;
  assign new_n4712 = ~new_n4709 & new_n4711;
  assign new_n4713 = new_n4712 ^ new_n4710;
  assign new_n4714 = new_n4713 ^ new_n4566;
  assign new_n4715 = n6 & n58;
  assign new_n4716 = new_n4715 ^ new_n4713;
  assign new_n4717 = ~new_n4714 & new_n4716;
  assign new_n4718 = new_n4717 ^ new_n4715;
  assign new_n4719 = new_n4529 ^ new_n4528;
  assign new_n4720 = new_n4719 ^ new_n4718;
  assign new_n4721 = n5 & n58;
  assign new_n4722 = new_n4721 ^ new_n4718;
  assign new_n4723 = ~new_n4720 & new_n4722;
  assign new_n4724 = new_n4723 ^ new_n4721;
  assign new_n4725 = new_n4724 ^ new_n4565;
  assign new_n4726 = n4 & n58;
  assign new_n4727 = new_n4726 ^ new_n4724;
  assign new_n4728 = ~new_n4725 & new_n4727;
  assign new_n4729 = new_n4728 ^ new_n4726;
  assign new_n4730 = new_n4540 ^ new_n4539;
  assign new_n4731 = new_n4730 ^ new_n4729;
  assign new_n4732 = n3 & n58;
  assign new_n4733 = new_n4732 ^ new_n4729;
  assign new_n4734 = ~new_n4731 & new_n4733;
  assign new_n4735 = new_n4734 ^ new_n4732;
  assign new_n4736 = new_n4735 ^ new_n4564;
  assign new_n4737 = n2 & n58;
  assign new_n4738 = new_n4737 ^ new_n4735;
  assign new_n4739 = ~new_n4736 & new_n4738;
  assign new_n4740 = new_n4739 ^ new_n4737;
  assign new_n4741 = new_n4551 ^ new_n4550;
  assign new_n4742 = new_n4741 ^ new_n4740;
  assign new_n4743 = n1 & n58;
  assign new_n4744 = new_n4743 ^ new_n4740;
  assign new_n4745 = ~new_n4742 & new_n4744;
  assign new_n4746 = new_n4745 ^ new_n4743;
  assign new_n4747 = new_n4557 ^ new_n4556;
  assign new_n4748 = new_n4746 & new_n4747;
  assign new_n4749 = new_n4560 ^ new_n4377;
  assign new_n4750 = new_n4748 & new_n4749;
  assign new_n4751 = new_n4749 ^ new_n4748;
  assign new_n4752 = new_n4751 ^ new_n4750;
  assign new_n4753 = ~new_n4563 & new_n4752;
  assign new_n4754 = new_n4743 ^ new_n4742;
  assign new_n4755 = new_n4732 ^ new_n4731;
  assign new_n4756 = new_n4721 ^ new_n4720;
  assign new_n4757 = new_n4710 ^ new_n4709;
  assign new_n4758 = new_n4699 ^ new_n4698;
  assign new_n4759 = new_n4688 ^ new_n4687;
  assign new_n4760 = new_n4677 ^ new_n4676;
  assign new_n4761 = new_n4666 ^ new_n4665;
  assign new_n4762 = new_n4655 ^ new_n4654;
  assign new_n4763 = new_n4644 ^ new_n4643;
  assign new_n4764 = new_n4633 ^ new_n4632;
  assign new_n4765 = new_n4622 ^ new_n4621;
  assign new_n4766 = new_n4611 ^ new_n4610;
  assign new_n4767 = new_n4600 ^ new_n4599;
  assign new_n4768 = new_n4589 ^ new_n4588;
  assign new_n4769 = new_n4584 ^ new_n4583;
  assign new_n4770 = n32 & n58;
  assign new_n4771 = n31 & n59;
  assign new_n4772 = new_n4770 & new_n4771;
  assign new_n4773 = new_n4580 ^ new_n4579;
  assign new_n4774 = new_n4773 ^ new_n4772;
  assign new_n4775 = n30 & n59;
  assign new_n4776 = new_n4775 ^ new_n4772;
  assign new_n4777 = ~new_n4774 & new_n4776;
  assign new_n4778 = new_n4777 ^ new_n4775;
  assign new_n4779 = new_n4778 ^ new_n4769;
  assign new_n4780 = n29 & n59;
  assign new_n4781 = new_n4780 ^ new_n4778;
  assign new_n4782 = ~new_n4779 & new_n4781;
  assign new_n4783 = new_n4782 ^ new_n4780;
  assign new_n4784 = new_n4783 ^ new_n4768;
  assign new_n4785 = n28 & n59;
  assign new_n4786 = new_n4785 ^ new_n4783;
  assign new_n4787 = ~new_n4784 & new_n4786;
  assign new_n4788 = new_n4787 ^ new_n4785;
  assign new_n4789 = new_n4594 ^ new_n4593;
  assign new_n4790 = new_n4789 ^ new_n4788;
  assign new_n4791 = n27 & n59;
  assign new_n4792 = new_n4791 ^ new_n4788;
  assign new_n4793 = ~new_n4790 & new_n4792;
  assign new_n4794 = new_n4793 ^ new_n4791;
  assign new_n4795 = new_n4794 ^ new_n4767;
  assign new_n4796 = n26 & n59;
  assign new_n4797 = new_n4796 ^ new_n4794;
  assign new_n4798 = ~new_n4795 & new_n4797;
  assign new_n4799 = new_n4798 ^ new_n4796;
  assign new_n4800 = new_n4605 ^ new_n4604;
  assign new_n4801 = new_n4800 ^ new_n4799;
  assign new_n4802 = n25 & n59;
  assign new_n4803 = new_n4802 ^ new_n4799;
  assign new_n4804 = ~new_n4801 & new_n4803;
  assign new_n4805 = new_n4804 ^ new_n4802;
  assign new_n4806 = new_n4805 ^ new_n4766;
  assign new_n4807 = n24 & n59;
  assign new_n4808 = new_n4807 ^ new_n4805;
  assign new_n4809 = ~new_n4806 & new_n4808;
  assign new_n4810 = new_n4809 ^ new_n4807;
  assign new_n4811 = new_n4616 ^ new_n4615;
  assign new_n4812 = new_n4811 ^ new_n4810;
  assign new_n4813 = n23 & n59;
  assign new_n4814 = new_n4813 ^ new_n4810;
  assign new_n4815 = ~new_n4812 & new_n4814;
  assign new_n4816 = new_n4815 ^ new_n4813;
  assign new_n4817 = new_n4816 ^ new_n4765;
  assign new_n4818 = n22 & n59;
  assign new_n4819 = new_n4818 ^ new_n4816;
  assign new_n4820 = ~new_n4817 & new_n4819;
  assign new_n4821 = new_n4820 ^ new_n4818;
  assign new_n4822 = new_n4627 ^ new_n4626;
  assign new_n4823 = new_n4822 ^ new_n4821;
  assign new_n4824 = n21 & n59;
  assign new_n4825 = new_n4824 ^ new_n4821;
  assign new_n4826 = ~new_n4823 & new_n4825;
  assign new_n4827 = new_n4826 ^ new_n4824;
  assign new_n4828 = new_n4827 ^ new_n4764;
  assign new_n4829 = n20 & n59;
  assign new_n4830 = new_n4829 ^ new_n4827;
  assign new_n4831 = ~new_n4828 & new_n4830;
  assign new_n4832 = new_n4831 ^ new_n4829;
  assign new_n4833 = new_n4638 ^ new_n4637;
  assign new_n4834 = new_n4833 ^ new_n4832;
  assign new_n4835 = n19 & n59;
  assign new_n4836 = new_n4835 ^ new_n4832;
  assign new_n4837 = ~new_n4834 & new_n4836;
  assign new_n4838 = new_n4837 ^ new_n4835;
  assign new_n4839 = new_n4838 ^ new_n4763;
  assign new_n4840 = n18 & n59;
  assign new_n4841 = new_n4840 ^ new_n4838;
  assign new_n4842 = ~new_n4839 & new_n4841;
  assign new_n4843 = new_n4842 ^ new_n4840;
  assign new_n4844 = new_n4649 ^ new_n4648;
  assign new_n4845 = new_n4844 ^ new_n4843;
  assign new_n4846 = n17 & n59;
  assign new_n4847 = new_n4846 ^ new_n4843;
  assign new_n4848 = ~new_n4845 & new_n4847;
  assign new_n4849 = new_n4848 ^ new_n4846;
  assign new_n4850 = new_n4849 ^ new_n4762;
  assign new_n4851 = n16 & n59;
  assign new_n4852 = new_n4851 ^ new_n4849;
  assign new_n4853 = ~new_n4850 & new_n4852;
  assign new_n4854 = new_n4853 ^ new_n4851;
  assign new_n4855 = new_n4660 ^ new_n4659;
  assign new_n4856 = new_n4855 ^ new_n4854;
  assign new_n4857 = n15 & n59;
  assign new_n4858 = new_n4857 ^ new_n4854;
  assign new_n4859 = ~new_n4856 & new_n4858;
  assign new_n4860 = new_n4859 ^ new_n4857;
  assign new_n4861 = new_n4860 ^ new_n4761;
  assign new_n4862 = n14 & n59;
  assign new_n4863 = new_n4862 ^ new_n4860;
  assign new_n4864 = ~new_n4861 & new_n4863;
  assign new_n4865 = new_n4864 ^ new_n4862;
  assign new_n4866 = new_n4671 ^ new_n4670;
  assign new_n4867 = new_n4866 ^ new_n4865;
  assign new_n4868 = n13 & n59;
  assign new_n4869 = new_n4868 ^ new_n4865;
  assign new_n4870 = ~new_n4867 & new_n4869;
  assign new_n4871 = new_n4870 ^ new_n4868;
  assign new_n4872 = new_n4871 ^ new_n4760;
  assign new_n4873 = n12 & n59;
  assign new_n4874 = new_n4873 ^ new_n4871;
  assign new_n4875 = ~new_n4872 & new_n4874;
  assign new_n4876 = new_n4875 ^ new_n4873;
  assign new_n4877 = new_n4682 ^ new_n4681;
  assign new_n4878 = new_n4877 ^ new_n4876;
  assign new_n4879 = n11 & n59;
  assign new_n4880 = new_n4879 ^ new_n4876;
  assign new_n4881 = ~new_n4878 & new_n4880;
  assign new_n4882 = new_n4881 ^ new_n4879;
  assign new_n4883 = new_n4882 ^ new_n4759;
  assign new_n4884 = n10 & n59;
  assign new_n4885 = new_n4884 ^ new_n4882;
  assign new_n4886 = ~new_n4883 & new_n4885;
  assign new_n4887 = new_n4886 ^ new_n4884;
  assign new_n4888 = new_n4693 ^ new_n4692;
  assign new_n4889 = new_n4888 ^ new_n4887;
  assign new_n4890 = n9 & n59;
  assign new_n4891 = new_n4890 ^ new_n4887;
  assign new_n4892 = ~new_n4889 & new_n4891;
  assign new_n4893 = new_n4892 ^ new_n4890;
  assign new_n4894 = new_n4893 ^ new_n4758;
  assign new_n4895 = n8 & n59;
  assign new_n4896 = new_n4895 ^ new_n4893;
  assign new_n4897 = ~new_n4894 & new_n4896;
  assign new_n4898 = new_n4897 ^ new_n4895;
  assign new_n4899 = new_n4704 ^ new_n4703;
  assign new_n4900 = new_n4899 ^ new_n4898;
  assign new_n4901 = n7 & n59;
  assign new_n4902 = new_n4901 ^ new_n4898;
  assign new_n4903 = ~new_n4900 & new_n4902;
  assign new_n4904 = new_n4903 ^ new_n4901;
  assign new_n4905 = new_n4904 ^ new_n4757;
  assign new_n4906 = n6 & n59;
  assign new_n4907 = new_n4906 ^ new_n4904;
  assign new_n4908 = ~new_n4905 & new_n4907;
  assign new_n4909 = new_n4908 ^ new_n4906;
  assign new_n4910 = new_n4715 ^ new_n4714;
  assign new_n4911 = new_n4910 ^ new_n4909;
  assign new_n4912 = n5 & n59;
  assign new_n4913 = new_n4912 ^ new_n4909;
  assign new_n4914 = ~new_n4911 & new_n4913;
  assign new_n4915 = new_n4914 ^ new_n4912;
  assign new_n4916 = new_n4915 ^ new_n4756;
  assign new_n4917 = n4 & n59;
  assign new_n4918 = new_n4917 ^ new_n4915;
  assign new_n4919 = ~new_n4916 & new_n4918;
  assign new_n4920 = new_n4919 ^ new_n4917;
  assign new_n4921 = new_n4726 ^ new_n4725;
  assign new_n4922 = new_n4921 ^ new_n4920;
  assign new_n4923 = n3 & n59;
  assign new_n4924 = new_n4923 ^ new_n4920;
  assign new_n4925 = ~new_n4922 & new_n4924;
  assign new_n4926 = new_n4925 ^ new_n4923;
  assign new_n4927 = new_n4926 ^ new_n4755;
  assign new_n4928 = n2 & n59;
  assign new_n4929 = new_n4928 ^ new_n4926;
  assign new_n4930 = ~new_n4927 & new_n4929;
  assign new_n4931 = new_n4930 ^ new_n4928;
  assign new_n4932 = new_n4737 ^ new_n4736;
  assign new_n4933 = new_n4932 ^ new_n4931;
  assign new_n4934 = n1 & n59;
  assign new_n4935 = new_n4934 ^ new_n4931;
  assign new_n4936 = ~new_n4933 & new_n4935;
  assign new_n4937 = new_n4936 ^ new_n4934;
  assign new_n4938 = new_n4754 & new_n4937;
  assign new_n4939 = new_n4747 ^ new_n4746;
  assign new_n4940 = new_n4939 ^ new_n4938;
  assign new_n4941 = ~new_n4938 & ~new_n4939;
  assign new_n4942 = new_n4941 ^ new_n4940;
  assign new_n4943 = new_n4942 ^ new_n4750;
  assign new_n4944 = ~new_n4943 & new_n4753;
  assign new_n4945 = new_n4562 ^ new_n4561;
  assign new_n4946 = new_n4945 ^ new_n4563;
  assign new_n4947 = new_n4946 ^ new_n4944;
  assign new_n4948 = ~new_n4947 & new_n4376;
  assign new_n4949 = new_n4948 ^ new_n4374;
  assign new_n4950 = new_n4934 ^ new_n4933;
  assign new_n4951 = new_n4771 ^ new_n4770;
  assign new_n4952 = n31 & n60;
  assign new_n4953 = n32 & n59;
  assign new_n4954 = new_n4952 & new_n4953;
  assign new_n4955 = new_n4954 ^ new_n4951;
  assign new_n4956 = n30 & n60;
  assign new_n4957 = new_n4956 ^ new_n4954;
  assign new_n4958 = ~new_n4955 & new_n4957;
  assign new_n4959 = new_n4958 ^ new_n4956;
  assign new_n4960 = new_n4775 ^ new_n4774;
  assign new_n4961 = new_n4960 ^ new_n4959;
  assign new_n4962 = n29 & n60;
  assign new_n4963 = new_n4962 ^ new_n4960;
  assign new_n4964 = ~new_n4961 & new_n4963;
  assign new_n4965 = new_n4964 ^ new_n4962;
  assign new_n4966 = new_n4780 ^ new_n4779;
  assign new_n4967 = new_n4966 ^ new_n4965;
  assign new_n4968 = n28 & n60;
  assign new_n4969 = new_n4968 ^ new_n4965;
  assign new_n4970 = ~new_n4967 & new_n4969;
  assign new_n4971 = new_n4970 ^ new_n4968;
  assign new_n4972 = new_n4785 ^ new_n4784;
  assign new_n4973 = new_n4972 ^ new_n4971;
  assign new_n4974 = n27 & n60;
  assign new_n4975 = new_n4974 ^ new_n4972;
  assign new_n4976 = ~new_n4973 & new_n4975;
  assign new_n4977 = new_n4976 ^ new_n4974;
  assign new_n4978 = new_n4791 ^ new_n4790;
  assign new_n4979 = new_n4978 ^ new_n4977;
  assign new_n4980 = n26 & n60;
  assign new_n4981 = new_n4980 ^ new_n4977;
  assign new_n4982 = ~new_n4979 & new_n4981;
  assign new_n4983 = new_n4982 ^ new_n4980;
  assign new_n4984 = new_n4796 ^ new_n4795;
  assign new_n4985 = new_n4984 ^ new_n4983;
  assign new_n4986 = n25 & n60;
  assign new_n4987 = new_n4986 ^ new_n4984;
  assign new_n4988 = ~new_n4985 & new_n4987;
  assign new_n4989 = new_n4988 ^ new_n4986;
  assign new_n4990 = new_n4802 ^ new_n4801;
  assign new_n4991 = new_n4990 ^ new_n4989;
  assign new_n4992 = n24 & n60;
  assign new_n4993 = new_n4992 ^ new_n4989;
  assign new_n4994 = ~new_n4991 & new_n4993;
  assign new_n4995 = new_n4994 ^ new_n4992;
  assign new_n4996 = new_n4807 ^ new_n4806;
  assign new_n4997 = new_n4996 ^ new_n4995;
  assign new_n4998 = n23 & n60;
  assign new_n4999 = new_n4998 ^ new_n4996;
  assign new_n5000 = ~new_n4997 & new_n4999;
  assign new_n5001 = new_n5000 ^ new_n4998;
  assign new_n5002 = new_n4813 ^ new_n4812;
  assign new_n5003 = new_n5002 ^ new_n5001;
  assign new_n5004 = n22 & n60;
  assign new_n5005 = new_n5004 ^ new_n5001;
  assign new_n5006 = ~new_n5003 & new_n5005;
  assign new_n5007 = new_n5006 ^ new_n5004;
  assign new_n5008 = new_n4818 ^ new_n4817;
  assign new_n5009 = new_n5008 ^ new_n5007;
  assign new_n5010 = n21 & n60;
  assign new_n5011 = new_n5010 ^ new_n5008;
  assign new_n5012 = ~new_n5009 & new_n5011;
  assign new_n5013 = new_n5012 ^ new_n5010;
  assign new_n5014 = new_n4824 ^ new_n4823;
  assign new_n5015 = new_n5014 ^ new_n5013;
  assign new_n5016 = n20 & n60;
  assign new_n5017 = new_n5016 ^ new_n5013;
  assign new_n5018 = ~new_n5015 & new_n5017;
  assign new_n5019 = new_n5018 ^ new_n5016;
  assign new_n5020 = new_n4829 ^ new_n4828;
  assign new_n5021 = new_n5020 ^ new_n5019;
  assign new_n5022 = n19 & n60;
  assign new_n5023 = new_n5022 ^ new_n5020;
  assign new_n5024 = ~new_n5021 & new_n5023;
  assign new_n5025 = new_n5024 ^ new_n5022;
  assign new_n5026 = new_n4835 ^ new_n4834;
  assign new_n5027 = new_n5026 ^ new_n5025;
  assign new_n5028 = n18 & n60;
  assign new_n5029 = new_n5028 ^ new_n5025;
  assign new_n5030 = ~new_n5027 & new_n5029;
  assign new_n5031 = new_n5030 ^ new_n5028;
  assign new_n5032 = new_n4840 ^ new_n4839;
  assign new_n5033 = new_n5032 ^ new_n5031;
  assign new_n5034 = n17 & n60;
  assign new_n5035 = new_n5034 ^ new_n5032;
  assign new_n5036 = ~new_n5033 & new_n5035;
  assign new_n5037 = new_n5036 ^ new_n5034;
  assign new_n5038 = new_n4846 ^ new_n4845;
  assign new_n5039 = new_n5038 ^ new_n5037;
  assign new_n5040 = n16 & n60;
  assign new_n5041 = new_n5040 ^ new_n5037;
  assign new_n5042 = ~new_n5039 & new_n5041;
  assign new_n5043 = new_n5042 ^ new_n5040;
  assign new_n5044 = new_n4851 ^ new_n4850;
  assign new_n5045 = new_n5044 ^ new_n5043;
  assign new_n5046 = n15 & n60;
  assign new_n5047 = new_n5046 ^ new_n5044;
  assign new_n5048 = ~new_n5045 & new_n5047;
  assign new_n5049 = new_n5048 ^ new_n5046;
  assign new_n5050 = new_n4857 ^ new_n4856;
  assign new_n5051 = new_n5050 ^ new_n5049;
  assign new_n5052 = n14 & n60;
  assign new_n5053 = new_n5052 ^ new_n5049;
  assign new_n5054 = ~new_n5051 & new_n5053;
  assign new_n5055 = new_n5054 ^ new_n5052;
  assign new_n5056 = new_n4862 ^ new_n4861;
  assign new_n5057 = new_n5056 ^ new_n5055;
  assign new_n5058 = n13 & n60;
  assign new_n5059 = new_n5058 ^ new_n5056;
  assign new_n5060 = ~new_n5057 & new_n5059;
  assign new_n5061 = new_n5060 ^ new_n5058;
  assign new_n5062 = new_n4868 ^ new_n4867;
  assign new_n5063 = new_n5062 ^ new_n5061;
  assign new_n5064 = n12 & n60;
  assign new_n5065 = new_n5064 ^ new_n5061;
  assign new_n5066 = ~new_n5063 & new_n5065;
  assign new_n5067 = new_n5066 ^ new_n5064;
  assign new_n5068 = new_n4873 ^ new_n4872;
  assign new_n5069 = new_n5068 ^ new_n5067;
  assign new_n5070 = n11 & n60;
  assign new_n5071 = new_n5070 ^ new_n5068;
  assign new_n5072 = ~new_n5069 & new_n5071;
  assign new_n5073 = new_n5072 ^ new_n5070;
  assign new_n5074 = new_n4879 ^ new_n4878;
  assign new_n5075 = new_n5074 ^ new_n5073;
  assign new_n5076 = n10 & n60;
  assign new_n5077 = new_n5076 ^ new_n5073;
  assign new_n5078 = ~new_n5075 & new_n5077;
  assign new_n5079 = new_n5078 ^ new_n5076;
  assign new_n5080 = new_n4884 ^ new_n4883;
  assign new_n5081 = new_n5080 ^ new_n5079;
  assign new_n5082 = n9 & n60;
  assign new_n5083 = new_n5082 ^ new_n5080;
  assign new_n5084 = ~new_n5081 & new_n5083;
  assign new_n5085 = new_n5084 ^ new_n5082;
  assign new_n5086 = new_n4890 ^ new_n4889;
  assign new_n5087 = new_n5086 ^ new_n5085;
  assign new_n5088 = n8 & n60;
  assign new_n5089 = new_n5088 ^ new_n5085;
  assign new_n5090 = ~new_n5087 & new_n5089;
  assign new_n5091 = new_n5090 ^ new_n5088;
  assign new_n5092 = new_n4895 ^ new_n4894;
  assign new_n5093 = new_n5092 ^ new_n5091;
  assign new_n5094 = n7 & n60;
  assign new_n5095 = new_n5094 ^ new_n5092;
  assign new_n5096 = ~new_n5093 & new_n5095;
  assign new_n5097 = new_n5096 ^ new_n5094;
  assign new_n5098 = new_n4901 ^ new_n4900;
  assign new_n5099 = new_n5098 ^ new_n5097;
  assign new_n5100 = n6 & n60;
  assign new_n5101 = new_n5100 ^ new_n5097;
  assign new_n5102 = ~new_n5099 & new_n5101;
  assign new_n5103 = new_n5102 ^ new_n5100;
  assign new_n5104 = new_n4906 ^ new_n4905;
  assign new_n5105 = new_n5104 ^ new_n5103;
  assign new_n5106 = n5 & n60;
  assign new_n5107 = new_n5106 ^ new_n5104;
  assign new_n5108 = ~new_n5105 & new_n5107;
  assign new_n5109 = new_n5108 ^ new_n5106;
  assign new_n5110 = new_n4912 ^ new_n4911;
  assign new_n5111 = new_n5110 ^ new_n5109;
  assign new_n5112 = n4 & n60;
  assign new_n5113 = new_n5112 ^ new_n5109;
  assign new_n5114 = ~new_n5111 & new_n5113;
  assign new_n5115 = new_n5114 ^ new_n5112;
  assign new_n5116 = new_n4917 ^ new_n4916;
  assign new_n5117 = new_n5116 ^ new_n5115;
  assign new_n5118 = n3 & n60;
  assign new_n5119 = new_n5118 ^ new_n5115;
  assign new_n5120 = ~new_n5117 & new_n5119;
  assign new_n5121 = new_n5120 ^ new_n5118;
  assign new_n5122 = new_n4923 ^ new_n4922;
  assign new_n5123 = new_n5122 ^ new_n5121;
  assign new_n5124 = n2 & n60;
  assign new_n5125 = new_n5124 ^ new_n5122;
  assign new_n5126 = ~new_n5123 & new_n5125;
  assign new_n5127 = new_n5126 ^ new_n5124;
  assign new_n5128 = new_n4928 ^ new_n4927;
  assign new_n5129 = new_n5128 ^ new_n5127;
  assign new_n5130 = n1 & n60;
  assign new_n5131 = new_n5130 ^ new_n5128;
  assign new_n5132 = ~new_n5129 & new_n5131;
  assign new_n5133 = new_n5132 ^ new_n5130;
  assign new_n5134 = new_n4950 & new_n5133;
  assign new_n5135 = new_n4937 ^ new_n4754;
  assign new_n5136 = new_n5134 & new_n5135;
  assign new_n5137 = new_n5135 ^ new_n5134;
  assign new_n5138 = new_n5137 ^ new_n5136;
  assign new_n5139 = new_n4953 ^ new_n4952;
  assign new_n5140 = n31 & n61;
  assign new_n5141 = n32 & n60;
  assign new_n5142 = new_n5140 & new_n5141;
  assign new_n5143 = new_n5142 ^ new_n5139;
  assign new_n5144 = n30 & n61;
  assign new_n5145 = new_n5144 ^ new_n5142;
  assign new_n5146 = ~new_n5143 & new_n5145;
  assign new_n5147 = new_n5146 ^ new_n5144;
  assign new_n5148 = new_n4956 ^ new_n4955;
  assign new_n5149 = new_n5148 ^ new_n5147;
  assign new_n5150 = n29 & n61;
  assign new_n5151 = new_n5150 ^ new_n5148;
  assign new_n5152 = ~new_n5149 & new_n5151;
  assign new_n5153 = new_n5152 ^ new_n5150;
  assign new_n5154 = new_n4962 ^ new_n4961;
  assign new_n5155 = new_n5154 ^ new_n5153;
  assign new_n5156 = n28 & n61;
  assign new_n5157 = new_n5156 ^ new_n5153;
  assign new_n5158 = ~new_n5155 & new_n5157;
  assign new_n5159 = new_n5158 ^ new_n5156;
  assign new_n5160 = new_n4968 ^ new_n4967;
  assign new_n5161 = new_n5160 ^ new_n5159;
  assign new_n5162 = n27 & n61;
  assign new_n5163 = new_n5162 ^ new_n5160;
  assign new_n5164 = ~new_n5161 & new_n5163;
  assign new_n5165 = new_n5164 ^ new_n5162;
  assign new_n5166 = new_n4974 ^ new_n4973;
  assign new_n5167 = new_n5166 ^ new_n5165;
  assign new_n5168 = n26 & n61;
  assign new_n5169 = new_n5168 ^ new_n5165;
  assign new_n5170 = ~new_n5167 & new_n5169;
  assign new_n5171 = new_n5170 ^ new_n5168;
  assign new_n5172 = new_n4980 ^ new_n4979;
  assign new_n5173 = new_n5172 ^ new_n5171;
  assign new_n5174 = n25 & n61;
  assign new_n5175 = new_n5174 ^ new_n5172;
  assign new_n5176 = ~new_n5173 & new_n5175;
  assign new_n5177 = new_n5176 ^ new_n5174;
  assign new_n5178 = new_n4986 ^ new_n4985;
  assign new_n5179 = new_n5178 ^ new_n5177;
  assign new_n5180 = n24 & n61;
  assign new_n5181 = new_n5180 ^ new_n5177;
  assign new_n5182 = ~new_n5179 & new_n5181;
  assign new_n5183 = new_n5182 ^ new_n5180;
  assign new_n5184 = new_n4992 ^ new_n4991;
  assign new_n5185 = new_n5184 ^ new_n5183;
  assign new_n5186 = n23 & n61;
  assign new_n5187 = new_n5186 ^ new_n5184;
  assign new_n5188 = ~new_n5185 & new_n5187;
  assign new_n5189 = new_n5188 ^ new_n5186;
  assign new_n5190 = new_n4998 ^ new_n4997;
  assign new_n5191 = new_n5190 ^ new_n5189;
  assign new_n5192 = n22 & n61;
  assign new_n5193 = new_n5192 ^ new_n5189;
  assign new_n5194 = ~new_n5191 & new_n5193;
  assign new_n5195 = new_n5194 ^ new_n5192;
  assign new_n5196 = new_n5004 ^ new_n5003;
  assign new_n5197 = new_n5196 ^ new_n5195;
  assign new_n5198 = n21 & n61;
  assign new_n5199 = new_n5198 ^ new_n5196;
  assign new_n5200 = ~new_n5197 & new_n5199;
  assign new_n5201 = new_n5200 ^ new_n5198;
  assign new_n5202 = new_n5010 ^ new_n5009;
  assign new_n5203 = new_n5202 ^ new_n5201;
  assign new_n5204 = n20 & n61;
  assign new_n5205 = new_n5204 ^ new_n5201;
  assign new_n5206 = ~new_n5203 & new_n5205;
  assign new_n5207 = new_n5206 ^ new_n5204;
  assign new_n5208 = new_n5016 ^ new_n5015;
  assign new_n5209 = new_n5208 ^ new_n5207;
  assign new_n5210 = n19 & n61;
  assign new_n5211 = new_n5210 ^ new_n5208;
  assign new_n5212 = ~new_n5209 & new_n5211;
  assign new_n5213 = new_n5212 ^ new_n5210;
  assign new_n5214 = new_n5022 ^ new_n5021;
  assign new_n5215 = new_n5214 ^ new_n5213;
  assign new_n5216 = n18 & n61;
  assign new_n5217 = new_n5216 ^ new_n5213;
  assign new_n5218 = ~new_n5215 & new_n5217;
  assign new_n5219 = new_n5218 ^ new_n5216;
  assign new_n5220 = new_n5028 ^ new_n5027;
  assign new_n5221 = new_n5220 ^ new_n5219;
  assign new_n5222 = n17 & n61;
  assign new_n5223 = new_n5222 ^ new_n5220;
  assign new_n5224 = ~new_n5221 & new_n5223;
  assign new_n5225 = new_n5224 ^ new_n5222;
  assign new_n5226 = new_n5034 ^ new_n5033;
  assign new_n5227 = new_n5226 ^ new_n5225;
  assign new_n5228 = n16 & n61;
  assign new_n5229 = new_n5228 ^ new_n5225;
  assign new_n5230 = ~new_n5227 & new_n5229;
  assign new_n5231 = new_n5230 ^ new_n5228;
  assign new_n5232 = new_n5040 ^ new_n5039;
  assign new_n5233 = new_n5232 ^ new_n5231;
  assign new_n5234 = n15 & n61;
  assign new_n5235 = new_n5234 ^ new_n5232;
  assign new_n5236 = ~new_n5233 & new_n5235;
  assign new_n5237 = new_n5236 ^ new_n5234;
  assign new_n5238 = new_n5046 ^ new_n5045;
  assign new_n5239 = new_n5238 ^ new_n5237;
  assign new_n5240 = n14 & n61;
  assign new_n5241 = new_n5240 ^ new_n5237;
  assign new_n5242 = ~new_n5239 & new_n5241;
  assign new_n5243 = new_n5242 ^ new_n5240;
  assign new_n5244 = new_n5052 ^ new_n5051;
  assign new_n5245 = new_n5244 ^ new_n5243;
  assign new_n5246 = n13 & n61;
  assign new_n5247 = new_n5246 ^ new_n5244;
  assign new_n5248 = ~new_n5245 & new_n5247;
  assign new_n5249 = new_n5248 ^ new_n5246;
  assign new_n5250 = new_n5058 ^ new_n5057;
  assign new_n5251 = new_n5250 ^ new_n5249;
  assign new_n5252 = n12 & n61;
  assign new_n5253 = new_n5252 ^ new_n5249;
  assign new_n5254 = ~new_n5251 & new_n5253;
  assign new_n5255 = new_n5254 ^ new_n5252;
  assign new_n5256 = new_n5064 ^ new_n5063;
  assign new_n5257 = new_n5256 ^ new_n5255;
  assign new_n5258 = n11 & n61;
  assign new_n5259 = new_n5258 ^ new_n5256;
  assign new_n5260 = ~new_n5257 & new_n5259;
  assign new_n5261 = new_n5260 ^ new_n5258;
  assign new_n5262 = new_n5070 ^ new_n5069;
  assign new_n5263 = new_n5262 ^ new_n5261;
  assign new_n5264 = n10 & n61;
  assign new_n5265 = new_n5264 ^ new_n5261;
  assign new_n5266 = ~new_n5263 & new_n5265;
  assign new_n5267 = new_n5266 ^ new_n5264;
  assign new_n5268 = new_n5076 ^ new_n5075;
  assign new_n5269 = new_n5268 ^ new_n5267;
  assign new_n5270 = n9 & n61;
  assign new_n5271 = new_n5270 ^ new_n5268;
  assign new_n5272 = ~new_n5269 & new_n5271;
  assign new_n5273 = new_n5272 ^ new_n5270;
  assign new_n5274 = new_n5082 ^ new_n5081;
  assign new_n5275 = new_n5274 ^ new_n5273;
  assign new_n5276 = n8 & n61;
  assign new_n5277 = new_n5276 ^ new_n5273;
  assign new_n5278 = ~new_n5275 & new_n5277;
  assign new_n5279 = new_n5278 ^ new_n5276;
  assign new_n5280 = new_n5088 ^ new_n5087;
  assign new_n5281 = new_n5280 ^ new_n5279;
  assign new_n5282 = n7 & n61;
  assign new_n5283 = new_n5282 ^ new_n5280;
  assign new_n5284 = ~new_n5281 & new_n5283;
  assign new_n5285 = new_n5284 ^ new_n5282;
  assign new_n5286 = new_n5094 ^ new_n5093;
  assign new_n5287 = new_n5286 ^ new_n5285;
  assign new_n5288 = n6 & n61;
  assign new_n5289 = new_n5288 ^ new_n5285;
  assign new_n5290 = ~new_n5287 & new_n5289;
  assign new_n5291 = new_n5290 ^ new_n5288;
  assign new_n5292 = new_n5100 ^ new_n5099;
  assign new_n5293 = new_n5292 ^ new_n5291;
  assign new_n5294 = n5 & n61;
  assign new_n5295 = new_n5294 ^ new_n5292;
  assign new_n5296 = ~new_n5293 & new_n5295;
  assign new_n5297 = new_n5296 ^ new_n5294;
  assign new_n5298 = new_n5106 ^ new_n5105;
  assign new_n5299 = new_n5298 ^ new_n5297;
  assign new_n5300 = n4 & n61;
  assign new_n5301 = new_n5300 ^ new_n5297;
  assign new_n5302 = ~new_n5299 & new_n5301;
  assign new_n5303 = new_n5302 ^ new_n5300;
  assign new_n5304 = new_n5112 ^ new_n5111;
  assign new_n5305 = new_n5304 ^ new_n5303;
  assign new_n5306 = n3 & n61;
  assign new_n5307 = new_n5306 ^ new_n5304;
  assign new_n5308 = ~new_n5305 & new_n5307;
  assign new_n5309 = new_n5308 ^ new_n5306;
  assign new_n5310 = new_n5118 ^ new_n5117;
  assign new_n5311 = new_n5310 ^ new_n5309;
  assign new_n5312 = n2 & n61;
  assign new_n5313 = new_n5312 ^ new_n5309;
  assign new_n5314 = ~new_n5311 & new_n5313;
  assign new_n5315 = new_n5314 ^ new_n5312;
  assign new_n5316 = new_n5124 ^ new_n5123;
  assign new_n5317 = new_n5316 ^ new_n5315;
  assign new_n5318 = n1 & n61;
  assign new_n5319 = new_n5318 ^ new_n5316;
  assign new_n5320 = ~new_n5317 & new_n5319;
  assign new_n5321 = new_n5320 ^ new_n5318;
  assign new_n5322 = new_n5130 ^ new_n5129;
  assign new_n5323 = new_n5321 & new_n5322;
  assign new_n5324 = new_n5133 ^ new_n4950;
  assign new_n5325 = new_n5323 & new_n5324;
  assign new_n5326 = new_n5324 ^ new_n5323;
  assign new_n5327 = new_n5326 ^ new_n5325;
  assign new_n5328 = new_n5318 ^ new_n5317;
  assign new_n5329 = new_n5312 ^ new_n5311;
  assign new_n5330 = n2 & n62;
  assign new_n5331 = n3 & n62;
  assign new_n5332 = n4 & n62;
  assign new_n5333 = n5 & n62;
  assign new_n5334 = n6 & n62;
  assign new_n5335 = n7 & n62;
  assign new_n5336 = n8 & n62;
  assign new_n5337 = n9 & n62;
  assign new_n5338 = n10 & n62;
  assign new_n5339 = n11 & n62;
  assign new_n5340 = n12 & n62;
  assign new_n5341 = n13 & n62;
  assign new_n5342 = n14 & n62;
  assign new_n5343 = n15 & n62;
  assign new_n5344 = n16 & n62;
  assign new_n5345 = n17 & n62;
  assign new_n5346 = n18 & n62;
  assign new_n5347 = n19 & n62;
  assign new_n5348 = n20 & n62;
  assign new_n5349 = n21 & n62;
  assign new_n5350 = n22 & n62;
  assign new_n5351 = n23 & n62;
  assign new_n5352 = n24 & n62;
  assign new_n5353 = n25 & n62;
  assign new_n5354 = n26 & n62;
  assign new_n5355 = n27 & n62;
  assign new_n5356 = n28 & n62;
  assign new_n5357 = n29 & n62;
  assign new_n5358 = new_n5141 ^ new_n5140;
  assign new_n5359 = n32 & n61;
  assign new_n5360 = n31 & n62;
  assign new_n5361 = new_n5359 & new_n5360;
  assign new_n5362 = new_n5361 ^ new_n5358;
  assign new_n5363 = n30 & n62;
  assign new_n5364 = new_n5363 ^ new_n5361;
  assign new_n5365 = ~new_n5362 & new_n5364;
  assign new_n5366 = new_n5365 ^ new_n5363;
  assign new_n5367 = new_n5366 ^ new_n5357;
  assign new_n5368 = new_n5144 ^ new_n5143;
  assign new_n5369 = new_n5368 ^ new_n5366;
  assign new_n5370 = ~new_n5369 & new_n5367;
  assign new_n5371 = new_n5370 ^ new_n5357;
  assign new_n5372 = new_n5371 ^ new_n5356;
  assign new_n5373 = ~new_n5372 & new_n5356;
  assign new_n5374 = new_n5150 ^ new_n5149;
  assign new_n5375 = new_n5372 & new_n5374;
  assign new_n5376 = new_n5375 ^ new_n5373;
  assign new_n5377 = new_n5376 ^ new_n5355;
  assign new_n5378 = new_n5156 ^ new_n5155;
  assign new_n5379 = new_n5378 ^ new_n5376;
  assign new_n5380 = ~new_n5379 & new_n5377;
  assign new_n5381 = new_n5380 ^ new_n5355;
  assign new_n5382 = new_n5381 ^ new_n5354;
  assign new_n5383 = ~new_n5382 & new_n5354;
  assign new_n5384 = new_n5162 ^ new_n5161;
  assign new_n5385 = new_n5382 & new_n5384;
  assign new_n5386 = new_n5385 ^ new_n5383;
  assign new_n5387 = new_n5386 ^ new_n5353;
  assign new_n5388 = new_n5168 ^ new_n5167;
  assign new_n5389 = new_n5388 ^ new_n5386;
  assign new_n5390 = ~new_n5389 & new_n5387;
  assign new_n5391 = new_n5390 ^ new_n5353;
  assign new_n5392 = new_n5391 ^ new_n5352;
  assign new_n5393 = ~new_n5392 & new_n5352;
  assign new_n5394 = new_n5174 ^ new_n5173;
  assign new_n5395 = new_n5392 & new_n5394;
  assign new_n5396 = new_n5395 ^ new_n5393;
  assign new_n5397 = new_n5396 ^ new_n5351;
  assign new_n5398 = new_n5180 ^ new_n5179;
  assign new_n5399 = new_n5398 ^ new_n5396;
  assign new_n5400 = ~new_n5399 & new_n5397;
  assign new_n5401 = new_n5400 ^ new_n5351;
  assign new_n5402 = new_n5401 ^ new_n5350;
  assign new_n5403 = ~new_n5402 & new_n5350;
  assign new_n5404 = new_n5186 ^ new_n5185;
  assign new_n5405 = new_n5402 & new_n5404;
  assign new_n5406 = new_n5405 ^ new_n5403;
  assign new_n5407 = new_n5406 ^ new_n5349;
  assign new_n5408 = new_n5192 ^ new_n5191;
  assign new_n5409 = new_n5408 ^ new_n5406;
  assign new_n5410 = ~new_n5409 & new_n5407;
  assign new_n5411 = new_n5410 ^ new_n5349;
  assign new_n5412 = new_n5411 ^ new_n5348;
  assign new_n5413 = ~new_n5412 & new_n5348;
  assign new_n5414 = new_n5198 ^ new_n5197;
  assign new_n5415 = new_n5412 & new_n5414;
  assign new_n5416 = new_n5415 ^ new_n5413;
  assign new_n5417 = new_n5416 ^ new_n5347;
  assign new_n5418 = new_n5204 ^ new_n5203;
  assign new_n5419 = new_n5418 ^ new_n5416;
  assign new_n5420 = ~new_n5419 & new_n5417;
  assign new_n5421 = new_n5420 ^ new_n5347;
  assign new_n5422 = new_n5421 ^ new_n5346;
  assign new_n5423 = ~new_n5422 & new_n5346;
  assign new_n5424 = new_n5210 ^ new_n5209;
  assign new_n5425 = new_n5422 & new_n5424;
  assign new_n5426 = new_n5425 ^ new_n5423;
  assign new_n5427 = new_n5426 ^ new_n5345;
  assign new_n5428 = new_n5216 ^ new_n5215;
  assign new_n5429 = new_n5428 ^ new_n5426;
  assign new_n5430 = ~new_n5429 & new_n5427;
  assign new_n5431 = new_n5430 ^ new_n5345;
  assign new_n5432 = new_n5431 ^ new_n5344;
  assign new_n5433 = ~new_n5432 & new_n5344;
  assign new_n5434 = new_n5222 ^ new_n5221;
  assign new_n5435 = new_n5432 & new_n5434;
  assign new_n5436 = new_n5435 ^ new_n5433;
  assign new_n5437 = new_n5436 ^ new_n5343;
  assign new_n5438 = new_n5228 ^ new_n5227;
  assign new_n5439 = new_n5438 ^ new_n5436;
  assign new_n5440 = ~new_n5439 & new_n5437;
  assign new_n5441 = new_n5440 ^ new_n5343;
  assign new_n5442 = new_n5441 ^ new_n5342;
  assign new_n5443 = ~new_n5442 & new_n5342;
  assign new_n5444 = new_n5234 ^ new_n5233;
  assign new_n5445 = new_n5442 & new_n5444;
  assign new_n5446 = new_n5445 ^ new_n5443;
  assign new_n5447 = new_n5446 ^ new_n5341;
  assign new_n5448 = new_n5240 ^ new_n5239;
  assign new_n5449 = new_n5448 ^ new_n5446;
  assign new_n5450 = ~new_n5449 & new_n5447;
  assign new_n5451 = new_n5450 ^ new_n5341;
  assign new_n5452 = new_n5451 ^ new_n5340;
  assign new_n5453 = ~new_n5452 & new_n5340;
  assign new_n5454 = new_n5246 ^ new_n5245;
  assign new_n5455 = new_n5452 & new_n5454;
  assign new_n5456 = new_n5455 ^ new_n5453;
  assign new_n5457 = new_n5456 ^ new_n5339;
  assign new_n5458 = new_n5252 ^ new_n5251;
  assign new_n5459 = new_n5458 ^ new_n5456;
  assign new_n5460 = ~new_n5459 & new_n5457;
  assign new_n5461 = new_n5460 ^ new_n5339;
  assign new_n5462 = new_n5461 ^ new_n5338;
  assign new_n5463 = ~new_n5462 & new_n5338;
  assign new_n5464 = new_n5258 ^ new_n5257;
  assign new_n5465 = new_n5462 & new_n5464;
  assign new_n5466 = new_n5465 ^ new_n5463;
  assign new_n5467 = new_n5466 ^ new_n5337;
  assign new_n5468 = new_n5264 ^ new_n5263;
  assign new_n5469 = new_n5468 ^ new_n5466;
  assign new_n5470 = ~new_n5469 & new_n5467;
  assign new_n5471 = new_n5470 ^ new_n5337;
  assign new_n5472 = new_n5471 ^ new_n5336;
  assign new_n5473 = ~new_n5472 & new_n5336;
  assign new_n5474 = new_n5270 ^ new_n5269;
  assign new_n5475 = new_n5472 & new_n5474;
  assign new_n5476 = new_n5475 ^ new_n5473;
  assign new_n5477 = new_n5476 ^ new_n5335;
  assign new_n5478 = new_n5276 ^ new_n5275;
  assign new_n5479 = new_n5478 ^ new_n5476;
  assign new_n5480 = ~new_n5479 & new_n5477;
  assign new_n5481 = new_n5480 ^ new_n5335;
  assign new_n5482 = new_n5481 ^ new_n5334;
  assign new_n5483 = ~new_n5482 & new_n5334;
  assign new_n5484 = new_n5282 ^ new_n5281;
  assign new_n5485 = new_n5482 & new_n5484;
  assign new_n5486 = new_n5485 ^ new_n5483;
  assign new_n5487 = new_n5486 ^ new_n5333;
  assign new_n5488 = new_n5288 ^ new_n5287;
  assign new_n5489 = new_n5488 ^ new_n5486;
  assign new_n5490 = ~new_n5489 & new_n5487;
  assign new_n5491 = new_n5490 ^ new_n5333;
  assign new_n5492 = new_n5491 ^ new_n5332;
  assign new_n5493 = ~new_n5492 & new_n5332;
  assign new_n5494 = new_n5294 ^ new_n5293;
  assign new_n5495 = new_n5492 & new_n5494;
  assign new_n5496 = new_n5495 ^ new_n5493;
  assign new_n5497 = new_n5496 ^ new_n5331;
  assign new_n5498 = new_n5300 ^ new_n5299;
  assign new_n5499 = new_n5498 ^ new_n5496;
  assign new_n5500 = ~new_n5499 & new_n5497;
  assign new_n5501 = new_n5500 ^ new_n5331;
  assign new_n5502 = new_n5501 ^ new_n5330;
  assign new_n5503 = ~new_n5502 & new_n5330;
  assign new_n5504 = new_n5306 ^ new_n5305;
  assign new_n5505 = new_n5502 & new_n5504;
  assign new_n5506 = new_n5505 ^ new_n5503;
  assign new_n5507 = new_n5506 ^ new_n5329;
  assign new_n5508 = n1 & n62;
  assign new_n5509 = new_n5508 ^ new_n5506;
  assign new_n5510 = ~new_n5507 & new_n5509;
  assign new_n5511 = new_n5510 ^ new_n5508;
  assign new_n5512 = new_n5328 & new_n5511;
  assign new_n5513 = new_n5322 ^ new_n5321;
  assign new_n5514 = new_n5512 & new_n5513;
  assign new_n5515 = new_n5513 ^ new_n5512;
  assign new_n5516 = new_n5515 ^ new_n5514;
  assign new_n5517 = n1 & n63;
  assign new_n5518 = n2 & n63;
  assign new_n5519 = n3 & n63;
  assign new_n5520 = n4 & n63;
  assign new_n5521 = n5 & n63;
  assign new_n5522 = n6 & n63;
  assign new_n5523 = n7 & n63;
  assign new_n5524 = n8 & n63;
  assign new_n5525 = n9 & n63;
  assign new_n5526 = n10 & n63;
  assign new_n5527 = n11 & n63;
  assign new_n5528 = n12 & n63;
  assign new_n5529 = n13 & n63;
  assign new_n5530 = n14 & n63;
  assign new_n5531 = n15 & n63;
  assign new_n5532 = n16 & n63;
  assign new_n5533 = n17 & n63;
  assign new_n5534 = n18 & n63;
  assign new_n5535 = n19 & n63;
  assign new_n5536 = n20 & n63;
  assign new_n5537 = n21 & n63;
  assign new_n5538 = n22 & n63;
  assign new_n5539 = n23 & n63;
  assign new_n5540 = n24 & n63;
  assign new_n5541 = n25 & n63;
  assign new_n5542 = n26 & n63;
  assign new_n5543 = n27 & n63;
  assign new_n5544 = n28 & n63;
  assign new_n5545 = n29 & n63;
  assign new_n5546 = n31 & n63;
  assign new_n5547 = n32 & n62;
  assign new_n5548 = new_n5546 & new_n5547;
  assign new_n5549 = new_n5360 ^ new_n5359;
  assign new_n5550 = new_n5549 ^ new_n5548;
  assign new_n5551 = n30 & n63;
  assign new_n5552 = new_n5551 ^ new_n5548;
  assign new_n5553 = ~new_n5550 & new_n5552;
  assign new_n5554 = new_n5553 ^ new_n5551;
  assign new_n5555 = new_n5554 ^ new_n5545;
  assign new_n5556 = ~new_n5555 & new_n5545;
  assign new_n5557 = new_n5363 ^ new_n5362;
  assign new_n5558 = new_n5555 & new_n5557;
  assign new_n5559 = new_n5558 ^ new_n5556;
  assign new_n5560 = new_n5559 ^ new_n5544;
  assign new_n5561 = new_n5368 ^ new_n5367;
  assign new_n5562 = new_n5561 ^ new_n5544;
  assign new_n5563 = ~new_n5562 & new_n5560;
  assign new_n5564 = new_n5563 ^ new_n5559;
  assign new_n5565 = new_n5564 ^ new_n5543;
  assign new_n5566 = new_n5374 ^ new_n5372;
  assign new_n5567 = new_n5566 ^ new_n5564;
  assign new_n5568 = ~new_n5567 & new_n5565;
  assign new_n5569 = new_n5568 ^ new_n5543;
  assign new_n5570 = new_n5569 ^ new_n5542;
  assign new_n5571 = ~new_n5570 & new_n5542;
  assign new_n5572 = new_n5378 ^ new_n5377;
  assign new_n5573 = new_n5570 & new_n5572;
  assign new_n5574 = new_n5573 ^ new_n5571;
  assign new_n5575 = new_n5574 ^ new_n5541;
  assign new_n5576 = new_n5384 ^ new_n5382;
  assign new_n5577 = new_n5576 ^ new_n5541;
  assign new_n5578 = ~new_n5577 & new_n5575;
  assign new_n5579 = new_n5578 ^ new_n5574;
  assign new_n5580 = new_n5579 ^ new_n5540;
  assign new_n5581 = new_n5388 ^ new_n5387;
  assign new_n5582 = new_n5581 ^ new_n5579;
  assign new_n5583 = ~new_n5582 & new_n5580;
  assign new_n5584 = new_n5583 ^ new_n5540;
  assign new_n5585 = new_n5584 ^ new_n5539;
  assign new_n5586 = ~new_n5585 & new_n5539;
  assign new_n5587 = new_n5394 ^ new_n5392;
  assign new_n5588 = new_n5585 & new_n5587;
  assign new_n5589 = new_n5588 ^ new_n5586;
  assign new_n5590 = new_n5589 ^ new_n5538;
  assign new_n5591 = new_n5398 ^ new_n5397;
  assign new_n5592 = new_n5591 ^ new_n5538;
  assign new_n5593 = ~new_n5592 & new_n5590;
  assign new_n5594 = new_n5593 ^ new_n5589;
  assign new_n5595 = new_n5594 ^ new_n5537;
  assign new_n5596 = new_n5404 ^ new_n5402;
  assign new_n5597 = new_n5596 ^ new_n5594;
  assign new_n5598 = ~new_n5597 & new_n5595;
  assign new_n5599 = new_n5598 ^ new_n5537;
  assign new_n5600 = new_n5599 ^ new_n5536;
  assign new_n5601 = ~new_n5600 & new_n5536;
  assign new_n5602 = new_n5408 ^ new_n5407;
  assign new_n5603 = new_n5600 & new_n5602;
  assign new_n5604 = new_n5603 ^ new_n5601;
  assign new_n5605 = new_n5604 ^ new_n5535;
  assign new_n5606 = new_n5414 ^ new_n5412;
  assign new_n5607 = new_n5606 ^ new_n5535;
  assign new_n5608 = ~new_n5607 & new_n5605;
  assign new_n5609 = new_n5608 ^ new_n5604;
  assign new_n5610 = new_n5609 ^ new_n5534;
  assign new_n5611 = new_n5418 ^ new_n5417;
  assign new_n5612 = new_n5611 ^ new_n5609;
  assign new_n5613 = ~new_n5612 & new_n5610;
  assign new_n5614 = new_n5613 ^ new_n5534;
  assign new_n5615 = new_n5614 ^ new_n5533;
  assign new_n5616 = ~new_n5615 & new_n5533;
  assign new_n5617 = new_n5424 ^ new_n5422;
  assign new_n5618 = new_n5615 & new_n5617;
  assign new_n5619 = new_n5618 ^ new_n5616;
  assign new_n5620 = new_n5619 ^ new_n5532;
  assign new_n5621 = new_n5428 ^ new_n5427;
  assign new_n5622 = new_n5621 ^ new_n5532;
  assign new_n5623 = ~new_n5622 & new_n5620;
  assign new_n5624 = new_n5623 ^ new_n5619;
  assign new_n5625 = new_n5624 ^ new_n5531;
  assign new_n5626 = new_n5434 ^ new_n5432;
  assign new_n5627 = new_n5626 ^ new_n5624;
  assign new_n5628 = ~new_n5627 & new_n5625;
  assign new_n5629 = new_n5628 ^ new_n5531;
  assign new_n5630 = new_n5629 ^ new_n5530;
  assign new_n5631 = ~new_n5630 & new_n5530;
  assign new_n5632 = new_n5438 ^ new_n5437;
  assign new_n5633 = new_n5630 & new_n5632;
  assign new_n5634 = new_n5633 ^ new_n5631;
  assign new_n5635 = new_n5634 ^ new_n5529;
  assign new_n5636 = new_n5444 ^ new_n5442;
  assign new_n5637 = new_n5636 ^ new_n5529;
  assign new_n5638 = ~new_n5637 & new_n5635;
  assign new_n5639 = new_n5638 ^ new_n5634;
  assign new_n5640 = new_n5639 ^ new_n5528;
  assign new_n5641 = new_n5448 ^ new_n5447;
  assign new_n5642 = new_n5641 ^ new_n5639;
  assign new_n5643 = ~new_n5642 & new_n5640;
  assign new_n5644 = new_n5643 ^ new_n5528;
  assign new_n5645 = new_n5644 ^ new_n5527;
  assign new_n5646 = ~new_n5645 & new_n5527;
  assign new_n5647 = new_n5454 ^ new_n5452;
  assign new_n5648 = new_n5645 & new_n5647;
  assign new_n5649 = new_n5648 ^ new_n5646;
  assign new_n5650 = new_n5649 ^ new_n5526;
  assign new_n5651 = new_n5458 ^ new_n5457;
  assign new_n5652 = new_n5651 ^ new_n5526;
  assign new_n5653 = ~new_n5652 & new_n5650;
  assign new_n5654 = new_n5653 ^ new_n5649;
  assign new_n5655 = new_n5654 ^ new_n5525;
  assign new_n5656 = new_n5464 ^ new_n5462;
  assign new_n5657 = new_n5656 ^ new_n5654;
  assign new_n5658 = ~new_n5657 & new_n5655;
  assign new_n5659 = new_n5658 ^ new_n5525;
  assign new_n5660 = new_n5659 ^ new_n5524;
  assign new_n5661 = ~new_n5660 & new_n5524;
  assign new_n5662 = new_n5468 ^ new_n5467;
  assign new_n5663 = new_n5660 & new_n5662;
  assign new_n5664 = new_n5663 ^ new_n5661;
  assign new_n5665 = new_n5664 ^ new_n5523;
  assign new_n5666 = new_n5474 ^ new_n5472;
  assign new_n5667 = new_n5666 ^ new_n5523;
  assign new_n5668 = ~new_n5667 & new_n5665;
  assign new_n5669 = new_n5668 ^ new_n5664;
  assign new_n5670 = new_n5669 ^ new_n5522;
  assign new_n5671 = new_n5478 ^ new_n5477;
  assign new_n5672 = new_n5671 ^ new_n5669;
  assign new_n5673 = ~new_n5672 & new_n5670;
  assign new_n5674 = new_n5673 ^ new_n5522;
  assign new_n5675 = new_n5674 ^ new_n5521;
  assign new_n5676 = ~new_n5675 & new_n5521;
  assign new_n5677 = new_n5484 ^ new_n5482;
  assign new_n5678 = new_n5675 & new_n5677;
  assign new_n5679 = new_n5678 ^ new_n5676;
  assign new_n5680 = new_n5679 ^ new_n5520;
  assign new_n5681 = new_n5488 ^ new_n5487;
  assign new_n5682 = new_n5681 ^ new_n5520;
  assign new_n5683 = ~new_n5682 & new_n5680;
  assign new_n5684 = new_n5683 ^ new_n5679;
  assign new_n5685 = new_n5684 ^ new_n5519;
  assign new_n5686 = new_n5494 ^ new_n5492;
  assign new_n5687 = new_n5686 ^ new_n5684;
  assign new_n5688 = ~new_n5687 & new_n5685;
  assign new_n5689 = new_n5688 ^ new_n5519;
  assign new_n5690 = new_n5689 ^ new_n5518;
  assign new_n5691 = ~new_n5690 & new_n5518;
  assign new_n5692 = new_n5498 ^ new_n5497;
  assign new_n5693 = new_n5690 & new_n5692;
  assign new_n5694 = new_n5693 ^ new_n5691;
  assign new_n5695 = new_n5694 ^ new_n5517;
  assign new_n5696 = new_n5504 ^ new_n5502;
  assign new_n5697 = new_n5696 ^ new_n5517;
  assign new_n5698 = ~new_n5697 & new_n5695;
  assign new_n5699 = new_n5698 ^ new_n5694;
  assign new_n5700 = new_n5508 ^ new_n5507;
  assign new_n5701 = new_n5699 & new_n5700;
  assign new_n5702 = new_n5511 ^ new_n5328;
  assign new_n5703 = new_n5702 ^ new_n5701;
  assign new_n5704 = ~new_n5701 & ~new_n5702;
  assign new_n5705 = new_n5704 ^ new_n5703;
  assign new_n5706 = ~new_n5705 & new_n5516;
  assign new_n5707 = new_n5706 ^ new_n5514;
  assign new_n5708 = new_n5327 & new_n5707;
  assign new_n5709 = new_n5708 ^ new_n5325;
  assign new_n5710 = new_n5138 & new_n5709;
  assign new_n5711 = new_n5710 ^ new_n5136;
  assign new_n5712 = new_n5696 ^ new_n5695;
  assign new_n5713 = n1 & n64;
  assign new_n5714 = n2 & n64;
  assign new_n5715 = n3 & n64;
  assign new_n5716 = n4 & n64;
  assign new_n5717 = n5 & n64;
  assign new_n5718 = n6 & n64;
  assign new_n5719 = n7 & n64;
  assign new_n5720 = n8 & n64;
  assign new_n5721 = n9 & n64;
  assign new_n5722 = n10 & n64;
  assign new_n5723 = n11 & n64;
  assign new_n5724 = n12 & n64;
  assign new_n5725 = n13 & n64;
  assign new_n5726 = n14 & n64;
  assign new_n5727 = n15 & n64;
  assign new_n5728 = n16 & n64;
  assign new_n5729 = n17 & n64;
  assign new_n5730 = n18 & n64;
  assign new_n5731 = n19 & n64;
  assign new_n5732 = n20 & n64;
  assign new_n5733 = n21 & n64;
  assign new_n5734 = n22 & n64;
  assign new_n5735 = n23 & n64;
  assign new_n5736 = n24 & n64;
  assign new_n5737 = n25 & n64;
  assign new_n5738 = n26 & n64;
  assign new_n5739 = n27 & n64;
  assign new_n5740 = n28 & n64;
  assign new_n5741 = n29 & n64;
  assign new_n5742 = n31 & n64;
  assign new_n5743 = n32 & n63;
  assign new_n5744 = new_n5742 & new_n5743;
  assign new_n5745 = new_n5547 ^ new_n5546;
  assign new_n5746 = new_n5745 ^ new_n5744;
  assign new_n5747 = n30 & n64;
  assign new_n5748 = new_n5747 ^ new_n5744;
  assign new_n5749 = ~new_n5746 & new_n5748;
  assign new_n5750 = new_n5749 ^ new_n5747;
  assign new_n5751 = new_n5750 ^ new_n5741;
  assign new_n5752 = ~new_n5751 & new_n5741;
  assign new_n5753 = new_n5551 ^ new_n5550;
  assign new_n5754 = new_n5751 & new_n5753;
  assign new_n5755 = new_n5754 ^ new_n5752;
  assign new_n5756 = new_n5755 ^ new_n5740;
  assign new_n5757 = new_n5557 ^ new_n5555;
  assign new_n5758 = new_n5757 ^ new_n5740;
  assign new_n5759 = ~new_n5758 & new_n5756;
  assign new_n5760 = new_n5759 ^ new_n5755;
  assign new_n5761 = new_n5760 ^ new_n5739;
  assign new_n5762 = new_n5561 ^ new_n5560;
  assign new_n5763 = new_n5762 ^ new_n5760;
  assign new_n5764 = ~new_n5763 & new_n5761;
  assign new_n5765 = new_n5764 ^ new_n5739;
  assign new_n5766 = new_n5765 ^ new_n5738;
  assign new_n5767 = ~new_n5766 & new_n5738;
  assign new_n5768 = new_n5566 ^ new_n5565;
  assign new_n5769 = new_n5766 & new_n5768;
  assign new_n5770 = new_n5769 ^ new_n5767;
  assign new_n5771 = new_n5770 ^ new_n5737;
  assign new_n5772 = new_n5572 ^ new_n5570;
  assign new_n5773 = new_n5772 ^ new_n5737;
  assign new_n5774 = ~new_n5773 & new_n5771;
  assign new_n5775 = new_n5774 ^ new_n5770;
  assign new_n5776 = new_n5775 ^ new_n5736;
  assign new_n5777 = new_n5576 ^ new_n5575;
  assign new_n5778 = new_n5777 ^ new_n5775;
  assign new_n5779 = ~new_n5778 & new_n5776;
  assign new_n5780 = new_n5779 ^ new_n5736;
  assign new_n5781 = new_n5780 ^ new_n5735;
  assign new_n5782 = ~new_n5781 & new_n5735;
  assign new_n5783 = new_n5581 ^ new_n5580;
  assign new_n5784 = new_n5781 & new_n5783;
  assign new_n5785 = new_n5784 ^ new_n5782;
  assign new_n5786 = new_n5785 ^ new_n5734;
  assign new_n5787 = new_n5587 ^ new_n5585;
  assign new_n5788 = new_n5787 ^ new_n5734;
  assign new_n5789 = ~new_n5788 & new_n5786;
  assign new_n5790 = new_n5789 ^ new_n5785;
  assign new_n5791 = new_n5790 ^ new_n5733;
  assign new_n5792 = new_n5591 ^ new_n5590;
  assign new_n5793 = new_n5792 ^ new_n5790;
  assign new_n5794 = ~new_n5793 & new_n5791;
  assign new_n5795 = new_n5794 ^ new_n5733;
  assign new_n5796 = new_n5795 ^ new_n5732;
  assign new_n5797 = ~new_n5796 & new_n5732;
  assign new_n5798 = new_n5596 ^ new_n5595;
  assign new_n5799 = new_n5796 & new_n5798;
  assign new_n5800 = new_n5799 ^ new_n5797;
  assign new_n5801 = new_n5800 ^ new_n5731;
  assign new_n5802 = new_n5602 ^ new_n5600;
  assign new_n5803 = new_n5802 ^ new_n5731;
  assign new_n5804 = ~new_n5803 & new_n5801;
  assign new_n5805 = new_n5804 ^ new_n5800;
  assign new_n5806 = new_n5805 ^ new_n5730;
  assign new_n5807 = new_n5606 ^ new_n5605;
  assign new_n5808 = new_n5807 ^ new_n5805;
  assign new_n5809 = ~new_n5808 & new_n5806;
  assign new_n5810 = new_n5809 ^ new_n5730;
  assign new_n5811 = new_n5810 ^ new_n5729;
  assign new_n5812 = ~new_n5811 & new_n5729;
  assign new_n5813 = new_n5611 ^ new_n5610;
  assign new_n5814 = new_n5811 & new_n5813;
  assign new_n5815 = new_n5814 ^ new_n5812;
  assign new_n5816 = new_n5815 ^ new_n5728;
  assign new_n5817 = new_n5617 ^ new_n5615;
  assign new_n5818 = new_n5817 ^ new_n5728;
  assign new_n5819 = ~new_n5818 & new_n5816;
  assign new_n5820 = new_n5819 ^ new_n5815;
  assign new_n5821 = new_n5820 ^ new_n5727;
  assign new_n5822 = new_n5621 ^ new_n5620;
  assign new_n5823 = new_n5822 ^ new_n5820;
  assign new_n5824 = ~new_n5823 & new_n5821;
  assign new_n5825 = new_n5824 ^ new_n5727;
  assign new_n5826 = new_n5825 ^ new_n5726;
  assign new_n5827 = ~new_n5826 & new_n5726;
  assign new_n5828 = new_n5626 ^ new_n5625;
  assign new_n5829 = new_n5826 & new_n5828;
  assign new_n5830 = new_n5829 ^ new_n5827;
  assign new_n5831 = new_n5830 ^ new_n5725;
  assign new_n5832 = new_n5632 ^ new_n5630;
  assign new_n5833 = new_n5832 ^ new_n5725;
  assign new_n5834 = ~new_n5833 & new_n5831;
  assign new_n5835 = new_n5834 ^ new_n5830;
  assign new_n5836 = new_n5835 ^ new_n5724;
  assign new_n5837 = new_n5636 ^ new_n5635;
  assign new_n5838 = new_n5837 ^ new_n5835;
  assign new_n5839 = ~new_n5838 & new_n5836;
  assign new_n5840 = new_n5839 ^ new_n5724;
  assign new_n5841 = new_n5840 ^ new_n5723;
  assign new_n5842 = ~new_n5841 & new_n5723;
  assign new_n5843 = new_n5641 ^ new_n5640;
  assign new_n5844 = new_n5841 & new_n5843;
  assign new_n5845 = new_n5844 ^ new_n5842;
  assign new_n5846 = new_n5845 ^ new_n5722;
  assign new_n5847 = new_n5647 ^ new_n5645;
  assign new_n5848 = new_n5847 ^ new_n5722;
  assign new_n5849 = ~new_n5848 & new_n5846;
  assign new_n5850 = new_n5849 ^ new_n5845;
  assign new_n5851 = new_n5850 ^ new_n5721;
  assign new_n5852 = new_n5651 ^ new_n5650;
  assign new_n5853 = new_n5852 ^ new_n5850;
  assign new_n5854 = ~new_n5853 & new_n5851;
  assign new_n5855 = new_n5854 ^ new_n5721;
  assign new_n5856 = new_n5855 ^ new_n5720;
  assign new_n5857 = ~new_n5856 & new_n5720;
  assign new_n5858 = new_n5656 ^ new_n5655;
  assign new_n5859 = new_n5856 & new_n5858;
  assign new_n5860 = new_n5859 ^ new_n5857;
  assign new_n5861 = new_n5860 ^ new_n5719;
  assign new_n5862 = new_n5662 ^ new_n5660;
  assign new_n5863 = new_n5862 ^ new_n5719;
  assign new_n5864 = ~new_n5863 & new_n5861;
  assign new_n5865 = new_n5864 ^ new_n5860;
  assign new_n5866 = new_n5865 ^ new_n5718;
  assign new_n5867 = new_n5666 ^ new_n5665;
  assign new_n5868 = new_n5867 ^ new_n5865;
  assign new_n5869 = ~new_n5868 & new_n5866;
  assign new_n5870 = new_n5869 ^ new_n5718;
  assign new_n5871 = new_n5870 ^ new_n5717;
  assign new_n5872 = ~new_n5871 & new_n5717;
  assign new_n5873 = new_n5671 ^ new_n5670;
  assign new_n5874 = new_n5871 & new_n5873;
  assign new_n5875 = new_n5874 ^ new_n5872;
  assign new_n5876 = new_n5875 ^ new_n5716;
  assign new_n5877 = new_n5677 ^ new_n5675;
  assign new_n5878 = new_n5877 ^ new_n5716;
  assign new_n5879 = ~new_n5878 & new_n5876;
  assign new_n5880 = new_n5879 ^ new_n5875;
  assign new_n5881 = new_n5880 ^ new_n5715;
  assign new_n5882 = new_n5681 ^ new_n5680;
  assign new_n5883 = new_n5882 ^ new_n5880;
  assign new_n5884 = ~new_n5883 & new_n5881;
  assign new_n5885 = new_n5884 ^ new_n5715;
  assign new_n5886 = new_n5885 ^ new_n5714;
  assign new_n5887 = ~new_n5886 & new_n5714;
  assign new_n5888 = new_n5686 ^ new_n5685;
  assign new_n5889 = new_n5886 & new_n5888;
  assign new_n5890 = new_n5889 ^ new_n5887;
  assign new_n5891 = new_n5890 ^ new_n5713;
  assign new_n5892 = new_n5692 ^ new_n5690;
  assign new_n5893 = new_n5892 ^ new_n5713;
  assign new_n5894 = ~new_n5893 & new_n5891;
  assign new_n5895 = new_n5894 ^ new_n5890;
  assign new_n5896 = new_n5712 & new_n5895;
  assign new_n5897 = new_n5700 ^ new_n5699;
  assign new_n5898 = new_n5896 & new_n5897;
  assign new_n5899 = new_n5516 & new_n5898;
  assign new_n5900 = ~new_n5704 & new_n5327;
  assign new_n5901 = new_n5138 & new_n5900;
  assign new_n5902 = new_n5899 & new_n5901;
  assign new_n5903 = new_n5902 ^ new_n5711;
  assign new_n5904 = ~new_n4941 & new_n5903;
  assign new_n5905 = new_n4376 & new_n4753;
  assign new_n5906 = new_n5904 & new_n5905;
  assign new_n5907 = new_n5906 ^ new_n4949;
  assign new_n5908 = ~new_n4179 & new_n5907;
  assign new_n5909 = new_n3614 & new_n3991;
  assign new_n5910 = new_n5908 & new_n5909;
  assign new_n5911 = new_n5910 ^ new_n4187;
  assign new_n5912 = new_n5911 ^ new_n3239;
  assign new_n5913 = ~new_n5912 & new_n3425;
  assign new_n5914 = new_n5913 ^ new_n3424;
  assign new_n5915 = new_n5914 ^ new_n3052;
  assign new_n5916 = ~new_n5915 & new_n3238;
  assign new_n5917 = new_n5916 ^ new_n3237;
  assign new_n5918 = new_n5917 ^ new_n2865;
  assign new_n5919 = ~new_n5918 & new_n3051;
  assign new_n5920 = new_n5919 ^ new_n3050;
  assign new_n5921 = new_n5920 ^ new_n2678;
  assign new_n5922 = ~new_n5921 & new_n2864;
  assign new_n5923 = new_n5922 ^ new_n2863;
  assign new_n5924 = new_n5923 ^ new_n2491;
  assign new_n5925 = ~new_n5924 & new_n2677;
  assign new_n5926 = new_n5925 ^ new_n2676;
  assign new_n5927 = new_n5926 ^ new_n2304;
  assign new_n5928 = ~new_n5927 & new_n2490;
  assign new_n5929 = new_n5928 ^ new_n2489;
  assign new_n5930 = new_n5929 ^ new_n2117;
  assign new_n5931 = ~new_n5930 & new_n2303;
  assign new_n5932 = new_n5931 ^ new_n2302;
  assign new_n5933 = new_n5932 ^ new_n1930;
  assign new_n5934 = ~new_n5933 & new_n2116;
  assign new_n5935 = new_n5934 ^ new_n2115;
  assign new_n5936 = new_n5935 ^ new_n1743;
  assign new_n5937 = ~new_n5936 & new_n1929;
  assign new_n5938 = new_n5937 ^ new_n1928;
  assign new_n5939 = new_n5938 ^ new_n1556;
  assign new_n5940 = ~new_n5939 & new_n1742;
  assign new_n5941 = new_n5940 ^ new_n1741;
  assign new_n5942 = new_n5941 ^ new_n1369;
  assign new_n5943 = ~new_n5942 & new_n1555;
  assign new_n5944 = new_n5943 ^ new_n1554;
  assign new_n5945 = new_n5944 ^ new_n1182;
  assign new_n5946 = ~new_n5945 & new_n1368;
  assign new_n5947 = new_n5946 ^ new_n1367;
  assign new_n5948 = new_n5947 ^ new_n995;
  assign new_n5949 = ~new_n5948 & new_n1181;
  assign new_n5950 = new_n5949 ^ new_n1180;
  assign new_n5951 = new_n5950 ^ new_n808;
  assign new_n5952 = ~new_n5951 & new_n994;
  assign new_n5953 = new_n5952 ^ new_n993;
  assign new_n5954 = new_n5953 ^ new_n621;
  assign new_n5955 = ~new_n5954 & new_n807;
  assign new_n5956 = new_n5955 ^ new_n806;
  assign new_n5957 = new_n5956 ^ new_n434;
  assign new_n5958 = ~new_n5957 & new_n620;
  assign new_n5959 = new_n5958 ^ new_n619;
  assign new_n5960 = new_n433 & new_n5959;
  assign new_n5961 = new_n427 & new_n432;
  assign new_n5962 = new_n5961 ^ new_n5960;
  assign new_n5963 = new_n428 & new_n431;
  assign new_n5964 = new_n5963 ^ new_n5962;
  assign new_n5965 = new_n5959 ^ new_n433;
  assign new_n5966 = new_n5956 ^ new_n620;
  assign new_n5967 = new_n5953 ^ new_n807;
  assign new_n5968 = new_n5950 ^ new_n994;
  assign new_n5969 = new_n5947 ^ new_n1181;
  assign new_n5970 = new_n5944 ^ new_n1368;
  assign new_n5971 = new_n5941 ^ new_n1555;
  assign new_n5972 = new_n5938 ^ new_n1742;
  assign new_n5973 = new_n5935 ^ new_n1929;
  assign new_n5974 = new_n5932 ^ new_n2116;
  assign new_n5975 = new_n5929 ^ new_n2303;
  assign new_n5976 = new_n5926 ^ new_n2490;
  assign new_n5977 = new_n5923 ^ new_n2677;
  assign new_n5978 = new_n5920 ^ new_n2864;
  assign new_n5979 = new_n5917 ^ new_n3051;
  assign new_n5980 = new_n5914 ^ new_n3238;
  assign new_n5981 = new_n5911 ^ new_n3425;
  assign new_n5982 = new_n5908 ^ new_n4180;
  assign new_n5983 = ~new_n5982 & new_n3990;
  assign new_n5984 = new_n5983 ^ new_n3988;
  assign new_n5985 = ~new_n3801 & new_n5984;
  assign new_n5986 = new_n5985 ^ new_n4184;
  assign new_n5987 = new_n5986 ^ new_n3613;
  assign new_n5988 = new_n5984 ^ new_n4183;
  assign new_n5989 = new_n5982 ^ new_n3989;
  assign new_n5990 = new_n5907 ^ new_n4178;
  assign new_n5991 = new_n5904 ^ new_n4942;
  assign new_n5992 = ~new_n5991 & new_n4752;
  assign new_n5993 = new_n5992 ^ new_n4750;
  assign new_n5994 = ~new_n4563 & new_n5993;
  assign new_n5995 = new_n5994 ^ new_n4946;
  assign new_n5996 = new_n5995 ^ new_n4375;
  assign new_n5997 = new_n5993 ^ new_n4945;
  assign new_n5998 = new_n5991 ^ new_n4751;
  assign new_n5999 = new_n5903 ^ new_n4940;
  assign new_n6000 = new_n5898 ^ new_n5701;
  assign new_n6001 = new_n5702 & new_n6000;
  assign new_n6002 = new_n5516 & new_n6001;
  assign new_n6003 = new_n6002 ^ new_n5514;
  assign new_n6004 = new_n5327 & new_n6003;
  assign new_n6005 = new_n6004 ^ new_n5325;
  assign new_n6006 = new_n6005 ^ new_n5137;
  assign new_n6007 = new_n6003 ^ new_n5326;
  assign new_n6008 = new_n6001 ^ new_n5515;
  assign new_n6009 = new_n5898 ^ new_n5703;
  assign new_n6010 = new_n5897 ^ new_n5896;
  assign new_n6011 = new_n5895 ^ new_n5712;
  assign new_n6012 = new_n5892 ^ new_n5891;
  assign new_n6013 = new_n5888 ^ new_n5886;
  assign new_n6014 = new_n5882 ^ new_n5881;
  assign new_n6015 = new_n5877 ^ new_n5876;
  assign new_n6016 = new_n5873 ^ new_n5871;
  assign new_n6017 = new_n5867 ^ new_n5866;
  assign new_n6018 = new_n5862 ^ new_n5861;
  assign new_n6019 = new_n5858 ^ new_n5856;
  assign new_n6020 = new_n5852 ^ new_n5851;
  assign new_n6021 = new_n5847 ^ new_n5846;
  assign new_n6022 = new_n5843 ^ new_n5841;
  assign new_n6023 = new_n5837 ^ new_n5836;
  assign new_n6024 = new_n5832 ^ new_n5831;
  assign new_n6025 = new_n5828 ^ new_n5826;
  assign new_n6026 = new_n5822 ^ new_n5821;
  assign new_n6027 = new_n5817 ^ new_n5816;
  assign new_n6028 = new_n5813 ^ new_n5811;
  assign new_n6029 = new_n5807 ^ new_n5806;
  assign new_n6030 = new_n5802 ^ new_n5801;
  assign new_n6031 = new_n5798 ^ new_n5796;
  assign new_n6032 = new_n5792 ^ new_n5791;
  assign new_n6033 = new_n5787 ^ new_n5786;
  assign new_n6034 = new_n5783 ^ new_n5781;
  assign new_n6035 = new_n5777 ^ new_n5776;
  assign new_n6036 = new_n5772 ^ new_n5771;
  assign new_n6037 = new_n5768 ^ new_n5766;
  assign new_n6038 = new_n5762 ^ new_n5761;
  assign new_n6039 = new_n5757 ^ new_n5756;
  assign new_n6040 = new_n5753 ^ new_n5751;
  assign new_n6041 = new_n5747 ^ new_n5746;
  assign new_n6042 = new_n5743 ^ new_n5742;
  assign new_n6043 = n32 & n64;
  assign po0 = new_n5964;
  assign po1 = new_n5965;
  assign po2 = new_n5966;
  assign po3 = new_n5967;
  assign po4 = new_n5968;
  assign po5 = new_n5969;
  assign po6 = new_n5970;
  assign po7 = new_n5971;
  assign po8 = new_n5972;
  assign po9 = new_n5973;
  assign po10 = new_n5974;
  assign po11 = new_n5975;
  assign po12 = new_n5976;
  assign po13 = new_n5977;
  assign po14 = new_n5978;
  assign po15 = new_n5979;
  assign po16 = new_n5980;
  assign po17 = new_n5981;
  assign po18 = ~new_n5987;
  assign po19 = new_n5988;
  assign po20 = ~new_n5989;
  assign po21 = new_n5990;
  assign po22 = ~new_n5996;
  assign po23 = new_n5997;
  assign po24 = ~new_n5998;
  assign po25 = new_n5999;
  assign po26 = new_n6006;
  assign po27 = new_n6007;
  assign po28 = new_n6008;
  assign po29 = new_n6009;
  assign po30 = new_n6010;
  assign po31 = new_n6011;
  assign po32 = new_n6012;
  assign po33 = new_n6013;
  assign po34 = new_n6014;
  assign po35 = new_n6015;
  assign po36 = new_n6016;
  assign po37 = new_n6017;
  assign po38 = new_n6018;
  assign po39 = new_n6019;
  assign po40 = new_n6020;
  assign po41 = new_n6021;
  assign po42 = new_n6022;
  assign po43 = new_n6023;
  assign po44 = new_n6024;
  assign po45 = new_n6025;
  assign po46 = new_n6026;
  assign po47 = new_n6027;
  assign po48 = new_n6028;
  assign po49 = new_n6029;
  assign po50 = new_n6030;
  assign po51 = new_n6031;
  assign po52 = new_n6032;
  assign po53 = new_n6033;
  assign po54 = new_n6034;
  assign po55 = new_n6035;
  assign po56 = new_n6036;
  assign po57 = new_n6037;
  assign po58 = new_n6038;
  assign po59 = new_n6039;
  assign po60 = new_n6040;
  assign po61 = new_n6041;
  assign po62 = new_n6042;
  assign po63 = new_n6043;
endmodule


