module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 ;
  assign n17 = ~x2 & x3 ;
  assign n18 = ~x14 & x15 ;
  assign n19 = ~x12 & x13 ;
  assign n20 = ~x10 & x11 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = n19 & n20 ;
  assign n23 = ~n21 & ~n22 ;
  assign n24 = n18 & ~n23 ;
  assign n25 = ~n18 & n23 ;
  assign n26 = ~n24 & ~n25 ;
  assign n27 = n17 & ~n26 ;
  assign n28 = ~n17 & n26 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = ~x8 & x9 ;
  assign n31 = ~x6 & x7 ;
  assign n32 = ~x4 & x5 ;
  assign n33 = n31 & n32 ;
  assign n34 = ~n31 & ~n32 ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = n30 & ~n35 ;
  assign n37 = ~n30 & n35 ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = n29 & ~n38 ;
  assign n40 = ~n27 & ~n39 ;
  assign n41 = ~n18 & ~n22 ;
  assign n42 = ~n21 & ~n41 ;
  assign n43 = ~n40 & n42 ;
  assign n44 = ~x0 & x1 ;
  assign n45 = ~n29 & n38 ;
  assign n46 = ~n39 & ~n45 ;
  assign n47 = n44 & n46 ;
  assign n48 = n40 & ~n42 ;
  assign n49 = ~n43 & ~n48 ;
  assign n50 = ~n30 & ~n33 ;
  assign n51 = ~n34 & ~n50 ;
  assign n52 = n49 & n51 ;
  assign n53 = ~n49 & ~n51 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n47 & n54 ;
  assign n56 = n43 & n55 ;
  assign n57 = x2 & x3 ;
  assign n58 = x14 & x15 ;
  assign n59 = x12 & x13 ;
  assign n60 = x10 & x11 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = n59 & n60 ;
  assign n63 = ~n61 & ~n62 ;
  assign n64 = n58 & ~n63 ;
  assign n65 = ~n58 & n63 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = n57 & ~n66 ;
  assign n68 = ~n57 & n66 ;
  assign n69 = x8 & x9 ;
  assign n70 = x6 & x7 ;
  assign n71 = x4 & x5 ;
  assign n72 = n70 & n71 ;
  assign n73 = ~n70 & ~n71 ;
  assign n74 = ~n72 & ~n73 ;
  assign n75 = n69 & ~n74 ;
  assign n76 = ~n69 & n74 ;
  assign n77 = ~n75 & ~n76 ;
  assign n78 = ~n68 & ~n77 ;
  assign n79 = ~n67 & ~n78 ;
  assign n80 = ~n58 & ~n62 ;
  assign n81 = ~n61 & ~n80 ;
  assign n82 = ~n79 & n81 ;
  assign n83 = x0 & x1 ;
  assign n84 = ~n67 & ~n68 ;
  assign n85 = n77 & n84 ;
  assign n86 = ~n77 & ~n84 ;
  assign n87 = ~n85 & ~n86 ;
  assign n88 = n83 & ~n87 ;
  assign n89 = n79 & ~n81 ;
  assign n90 = ~n82 & ~n89 ;
  assign n91 = ~n69 & ~n72 ;
  assign n92 = ~n73 & ~n91 ;
  assign n93 = n90 & n92 ;
  assign n94 = ~n90 & ~n92 ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = n88 & n95 ;
  assign n97 = n82 & n96 ;
  assign n98 = ~n56 & n97 ;
  assign n99 = ~n82 & ~n93 ;
  assign n100 = ~n96 & n99 ;
  assign n101 = ~n97 & ~n100 ;
  assign n102 = ~n43 & ~n52 ;
  assign n103 = ~n55 & n102 ;
  assign n104 = ~n56 & ~n103 ;
  assign n105 = n101 & ~n104 ;
  assign n106 = ~n88 & ~n95 ;
  assign n107 = ~n96 & ~n106 ;
  assign n108 = ~n54 & n107 ;
  assign n109 = ~n83 & n87 ;
  assign n110 = ~n88 & ~n109 ;
  assign n111 = ~n44 & ~n46 ;
  assign n112 = ~n47 & ~n111 ;
  assign n113 = ~n110 & n112 ;
  assign n114 = ~n108 & n113 ;
  assign n115 = ~n47 & ~n54 ;
  assign n116 = ~n55 & ~n115 ;
  assign n117 = ~n107 & n116 ;
  assign n118 = ~n114 & ~n117 ;
  assign n119 = ~n105 & ~n118 ;
  assign n120 = n56 & ~n97 ;
  assign n121 = ~n101 & n104 ;
  assign n122 = ~n120 & ~n121 ;
  assign n123 = ~n119 & n122 ;
  assign n124 = ~n98 & ~n123 ;
  assign n125 = ~x0 & ~x1 ;
  assign n126 = ~x8 & ~x9 ;
  assign n127 = ~x6 & ~x7 ;
  assign n128 = ~x4 & ~x5 ;
  assign n129 = ~n127 & ~n128 ;
  assign n130 = n127 & n128 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = ~n126 & n131 ;
  assign n133 = n126 & ~n131 ;
  assign n134 = ~n132 & ~n133 ;
  assign n135 = ~x14 & ~x15 ;
  assign n136 = ~x12 & ~x13 ;
  assign n137 = ~x10 & ~x11 ;
  assign n138 = ~n136 & ~n137 ;
  assign n139 = n136 & n137 ;
  assign n140 = ~n138 & ~n139 ;
  assign n141 = ~n135 & n140 ;
  assign n142 = n135 & ~n140 ;
  assign n143 = ~n141 & ~n142 ;
  assign n144 = ~x2 & ~x3 ;
  assign n145 = n143 & ~n144 ;
  assign n146 = ~n143 & n144 ;
  assign n147 = ~n145 & ~n146 ;
  assign n148 = n134 & n147 ;
  assign n149 = ~n134 & ~n147 ;
  assign n150 = ~n148 & ~n149 ;
  assign n151 = n125 & ~n150 ;
  assign n152 = ~n129 & ~n132 ;
  assign n153 = ~n138 & ~n141 ;
  assign n154 = ~n145 & ~n148 ;
  assign n155 = ~n153 & ~n154 ;
  assign n156 = n153 & n154 ;
  assign n157 = ~n155 & ~n156 ;
  assign n158 = n152 & ~n157 ;
  assign n159 = ~n152 & n157 ;
  assign n160 = ~n158 & ~n159 ;
  assign n161 = n151 & ~n160 ;
  assign n162 = ~n155 & ~n159 ;
  assign n163 = n161 & n162 ;
  assign n164 = x2 & ~x3 ;
  assign n165 = x14 & ~x15 ;
  assign n166 = x12 & ~x13 ;
  assign n167 = x10 & ~x11 ;
  assign n168 = ~n166 & ~n167 ;
  assign n169 = n166 & n167 ;
  assign n170 = ~n168 & ~n169 ;
  assign n171 = n165 & ~n170 ;
  assign n172 = ~n165 & n170 ;
  assign n173 = ~n171 & ~n172 ;
  assign n174 = n164 & ~n173 ;
  assign n175 = ~n164 & n173 ;
  assign n176 = ~n174 & ~n175 ;
  assign n177 = x8 & ~x9 ;
  assign n178 = x6 & ~x7 ;
  assign n179 = x4 & ~x5 ;
  assign n180 = n178 & n179 ;
  assign n181 = ~n178 & ~n179 ;
  assign n182 = ~n180 & ~n181 ;
  assign n183 = n177 & ~n182 ;
  assign n184 = ~n177 & n182 ;
  assign n185 = ~n183 & ~n184 ;
  assign n186 = n176 & ~n185 ;
  assign n187 = ~n174 & ~n186 ;
  assign n188 = ~n165 & ~n169 ;
  assign n189 = ~n168 & ~n188 ;
  assign n190 = ~n187 & n189 ;
  assign n191 = x0 & ~x1 ;
  assign n192 = ~n176 & n185 ;
  assign n193 = ~n186 & ~n192 ;
  assign n194 = n191 & n193 ;
  assign n195 = n187 & ~n189 ;
  assign n196 = ~n190 & ~n195 ;
  assign n197 = ~n177 & ~n180 ;
  assign n198 = ~n181 & ~n197 ;
  assign n199 = n196 & n198 ;
  assign n200 = ~n196 & ~n198 ;
  assign n201 = ~n199 & ~n200 ;
  assign n202 = n194 & n201 ;
  assign n203 = n190 & n202 ;
  assign n204 = ~n163 & ~n203 ;
  assign n205 = ~n56 & ~n97 ;
  assign n206 = n204 & ~n205 ;
  assign n207 = ~n204 & n205 ;
  assign n208 = ~n190 & ~n199 ;
  assign n209 = ~n202 & n208 ;
  assign n210 = ~n161 & ~n162 ;
  assign n211 = n209 & n210 ;
  assign n212 = n204 & ~n211 ;
  assign n213 = n100 & n103 ;
  assign n214 = n205 & ~n213 ;
  assign n215 = ~n212 & n214 ;
  assign n216 = n107 & ~n124 ;
  assign n217 = n116 & n124 ;
  assign n218 = ~n216 & ~n217 ;
  assign n219 = ~n112 & n124 ;
  assign n220 = ~n110 & ~n124 ;
  assign n221 = ~n219 & ~n220 ;
  assign n222 = ~n125 & n150 ;
  assign n223 = ~n151 & ~n222 ;
  assign n224 = ~n163 & n203 ;
  assign n225 = ~n203 & ~n209 ;
  assign n226 = ~n163 & ~n210 ;
  assign n227 = n225 & ~n226 ;
  assign n228 = ~n151 & n160 ;
  assign n229 = ~n161 & ~n228 ;
  assign n230 = ~n191 & ~n193 ;
  assign n231 = ~n194 & ~n230 ;
  assign n232 = n223 & ~n231 ;
  assign n233 = ~n229 & ~n232 ;
  assign n234 = ~n194 & ~n201 ;
  assign n235 = ~n202 & ~n234 ;
  assign n236 = ~n160 & n232 ;
  assign n237 = n235 & ~n236 ;
  assign n238 = ~n233 & ~n237 ;
  assign n239 = ~n227 & n238 ;
  assign n240 = n163 & ~n203 ;
  assign n241 = ~n225 & n226 ;
  assign n242 = ~n240 & ~n241 ;
  assign n243 = ~n239 & n242 ;
  assign n244 = ~n224 & ~n243 ;
  assign n245 = ~n223 & n244 ;
  assign n246 = ~n231 & ~n244 ;
  assign n247 = ~n245 & ~n246 ;
  assign n248 = ~n221 & n247 ;
  assign n249 = ~n218 & ~n248 ;
  assign n250 = ~n229 & n244 ;
  assign n251 = ~n235 & ~n244 ;
  assign n252 = ~n250 & ~n251 ;
  assign n253 = ~n249 & n252 ;
  assign n254 = n212 & ~n214 ;
  assign n255 = n218 & n248 ;
  assign n256 = ~n254 & ~n255 ;
  assign n257 = ~n253 & n256 ;
  assign n258 = ~n215 & ~n257 ;
  assign n259 = ~n207 & ~n258 ;
  assign n260 = ~n206 & ~n259 ;
  assign n261 = ~n124 & ~n260 ;
  assign n262 = ~n244 & n260 ;
  assign n263 = ~n261 & ~n262 ;
  assign y0 = ~n263 ;
  assign y1 = ~n260 ;
endmodule
