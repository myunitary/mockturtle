module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 ;
  assign n25 = x5 & x13 ;
  assign n26 = x6 & x14 ;
  assign n27 = ~n25 & ~n26 ;
  assign n28 = ~x5 & ~x13 ;
  assign n29 = ~x4 & ~x12 ;
  assign n30 = ~n28 & ~n29 ;
  assign n31 = ~n27 & n30 ;
  assign n32 = x3 & x11 ;
  assign n33 = x4 & x12 ;
  assign n34 = ~n32 & ~n33 ;
  assign n22 = x10 ^ x2 ;
  assign n23 = ~x3 & ~x11 ;
  assign n35 = ~n22 & ~n23 ;
  assign n36 = n34 & n35 ;
  assign n37 = ~n31 & n36 ;
  assign n24 = ~n22 & n23 ;
  assign n38 = n37 ^ n24 ;
  assign n40 = x14 ^ x6 ;
  assign n41 = x7 & x15 ;
  assign n42 = n40 & n41 ;
  assign n43 = x13 ^ x5 ;
  assign n44 = n42 & n43 ;
  assign n20 = x1 & x9 ;
  assign n21 = ~x8 & n20 ;
  assign n45 = x12 ^ x4 ;
  assign n46 = x11 ^ x3 ;
  assign n47 = n45 & n46 ;
  assign n48 = ~n21 & n47 ;
  assign n49 = n44 & n48 ;
  assign n50 = ~n38 & n49 ;
  assign n39 = n21 & ~n38 ;
  assign n51 = n50 ^ n39 ;
  assign n53 = n44 & n47 ;
  assign n17 = x9 ^ x1 ;
  assign n18 = x2 & x10 ;
  assign n19 = ~n17 & ~n18 ;
  assign n54 = x0 & x8 ;
  assign n55 = ~n20 & n54 ;
  assign n56 = ~n21 & ~n55 ;
  assign n57 = ~n19 & ~n56 ;
  assign n58 = n53 & n57 ;
  assign n59 = n51 & n58 ;
  assign n52 = ~n19 & n51 ;
  assign n60 = n59 ^ n52 ;
  assign n61 = ~x2 & ~x10 ;
  assign n62 = ~n23 & ~n61 ;
  assign n63 = n34 & n62 ;
  assign n64 = ~n31 & n63 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = ~x0 & ~x8 ;
  assign n67 = ~n18 & ~n20 ;
  assign n68 = ~n66 & n67 ;
  assign n69 = ~n65 & n68 ;
  assign n70 = x2 & ~n23 ;
  assign n71 = n34 & n70 ;
  assign n72 = ~n31 & n71 ;
  assign n73 = n72 ^ n70 ;
  assign n74 = ~x0 & x10 ;
  assign n75 = n21 & n74 ;
  assign n76 = ~x1 & ~x9 ;
  assign n77 = ~n54 & ~n76 ;
  assign n78 = ~n66 & ~n77 ;
  assign n79 = n75 & ~n78 ;
  assign n80 = n73 & n79 ;
  assign n81 = n80 ^ n78 ;
  assign n82 = ~n69 & ~n81 ;
  assign n83 = ~n60 & ~n82 ;
  assign n84 = n73 ^ n17 ;
  assign n85 = ~n23 & n34 ;
  assign n86 = ~n31 & n85 ;
  assign n87 = n86 ^ n23 ;
  assign n88 = n87 ^ n22 ;
  assign n89 = n84 & ~n88 ;
  assign n90 = x8 ^ x0 ;
  assign n91 = n90 ^ n20 ;
  assign n92 = n91 ^ n53 ;
  assign n93 = n89 & ~n92 ;
  assign n94 = n17 & n61 ;
  assign n95 = ~n76 & ~n94 ;
  assign n96 = n95 ^ n90 ;
  assign n97 = ~n89 & ~n96 ;
  assign n98 = ~n93 & ~n97 ;
  assign n102 = n61 ^ n17 ;
  assign n103 = n88 & ~n102 ;
  assign n100 = ~n53 & ~n88 ;
  assign n99 = ~n84 & ~n88 ;
  assign n101 = n100 ^ n99 ;
  assign n104 = n103 ^ n101 ;
  assign n105 = n88 ^ n53 ;
  assign n106 = n27 & ~n42 ;
  assign n107 = ~n28 & ~n106 ;
  assign n108 = ~n33 & ~n107 ;
  assign n109 = ~n29 & ~n108 ;
  assign n110 = n109 ^ n46 ;
  assign n111 = ~n26 & ~n44 ;
  assign n112 = n43 & ~n111 ;
  assign n113 = ~n25 & ~n112 ;
  assign n114 = n113 ^ n45 ;
  assign n115 = ~n26 & ~n42 ;
  assign n116 = n115 ^ n43 ;
  assign n117 = n41 ^ n40 ;
  assign y0 = n83 ;
  assign y1 = n98 ;
  assign y2 = n104 ;
  assign y3 = ~n105 ;
  assign y4 = n110 ;
  assign y5 = ~n114 ;
  assign y6 = ~n116 ;
  assign y7 = n117 ;
endmodule
