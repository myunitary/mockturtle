module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ;
  assign n9 = x0 & x1 ;
  assign n10 = n9 ^ x0 ;
  assign n11 = x2 & n10 ;
  assign n12 = x2 ^ x0 ;
  assign n13 = x1 & n12 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = x3 & n16 ;
  assign n18 = x4 ^ x2 ;
  assign n19 = x3 & n18 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n16 & n22 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n16 ;
  assign n26 = x4 & n25 ;
  assign n27 = x5 & n25 ;
  assign n28 = x6 & ~n16 ;
  assign n29 = x4 & x5 ;
  assign n30 = n29 ^ x4 ;
  assign n31 = ~n22 & ~n30 ;
  assign n32 = n28 & n31 ;
  assign n33 = n32 ^ x6 ;
  assign n34 = n25 ^ x7 ;
  assign n35 = x6 ^ x4 ;
  assign n36 = x5 & n35 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = n37 ^ x5 ;
  assign n39 = n38 ^ x6 ;
  assign n40 = n39 ^ x7 ;
  assign n41 = n39 & ~n40 ;
  assign n42 = n41 ^ x7 ;
  assign n43 = ~n34 & ~n42 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = n44 ^ n25 ;
  assign n46 = n45 ^ x7 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = n11 ;
  assign y3 = n17 ;
  assign y4 = n26 ;
  assign y5 = n27 ;
  assign y6 = n33 ;
  assign y7 = ~n46 ;
endmodule
