module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 ;
  assign n526 = x38 & x128 ;
  assign n527 = n526 ^ x38 ;
  assign n528 = x129 & n527 ;
  assign n523 = x39 & x128 ;
  assign n524 = x129 & n523 ;
  assign n525 = n524 ^ n523 ;
  assign n529 = n528 ^ n525 ;
  assign n535 = x37 & x128 ;
  assign n536 = x129 & n535 ;
  assign n537 = n536 ^ x129 ;
  assign n530 = x40 & x128 ;
  assign n531 = n530 ^ x40 ;
  assign n532 = x129 & n531 ;
  assign n533 = n532 ^ x129 ;
  assign n534 = n533 ^ n531 ;
  assign n538 = n537 ^ n534 ;
  assign n539 = n529 & n538 ;
  assign n540 = n539 ^ n538 ;
  assign n541 = n540 ^ n529 ;
  assign n139 = x130 & x131 ;
  assign n155 = n139 ^ x131 ;
  assign n500 = x45 & x128 ;
  assign n498 = x46 & x128 ;
  assign n499 = n498 ^ x46 ;
  assign n501 = n500 ^ n499 ;
  assign n502 = x129 & n501 ;
  assign n494 = x47 & x128 ;
  assign n492 = x48 & x128 ;
  assign n493 = n492 ^ x48 ;
  assign n495 = n494 ^ n493 ;
  assign n496 = x129 & n495 ;
  assign n497 = n496 ^ n495 ;
  assign n503 = n502 ^ n497 ;
  assign n136 = x132 & x133 ;
  assign n137 = n136 ^ x132 ;
  assign n170 = n139 ^ x130 ;
  assign n171 = n170 ^ x131 ;
  assign n504 = n137 & n171 ;
  assign n505 = n504 ^ n137 ;
  assign n506 = n503 & n505 ;
  assign n507 = n506 ^ n137 ;
  assign n486 = x41 & x128 ;
  assign n484 = x42 & x128 ;
  assign n485 = n484 ^ x42 ;
  assign n487 = n486 ^ n485 ;
  assign n488 = x129 & n487 ;
  assign n480 = x43 & x128 ;
  assign n478 = x44 & x128 ;
  assign n479 = n478 ^ x44 ;
  assign n481 = n480 ^ n479 ;
  assign n482 = x129 & n481 ;
  assign n483 = n482 ^ n481 ;
  assign n489 = n488 ^ n483 ;
  assign n490 = n137 & n170 ;
  assign n491 = n489 & n490 ;
  assign n508 = n507 ^ n491 ;
  assign n542 = n155 & n508 ;
  assign n543 = n541 & n542 ;
  assign n544 = n543 ^ n542 ;
  assign n545 = n544 ^ n542 ;
  assign n546 = n545 ^ n508 ;
  assign n517 = x33 & x128 ;
  assign n515 = x34 & x128 ;
  assign n516 = n515 ^ x34 ;
  assign n518 = n517 ^ n516 ;
  assign n519 = x129 & n518 ;
  assign n511 = x35 & x128 ;
  assign n509 = x36 & x128 ;
  assign n510 = n509 ^ x36 ;
  assign n512 = n511 ^ n510 ;
  assign n513 = x129 & n512 ;
  assign n514 = n513 ^ n512 ;
  assign n520 = n519 ^ n514 ;
  assign n521 = n139 & n520 ;
  assign n522 = n508 & n521 ;
  assign n547 = n546 ^ n522 ;
  assign n548 = n547 ^ x133 ;
  assign n138 = n137 ^ x133 ;
  assign n439 = x57 & x128 ;
  assign n437 = x58 & x128 ;
  assign n438 = n437 ^ x58 ;
  assign n440 = n439 ^ n438 ;
  assign n441 = x129 & n440 ;
  assign n433 = x59 & x128 ;
  assign n431 = x60 & x128 ;
  assign n432 = n431 ^ x60 ;
  assign n434 = n433 ^ n432 ;
  assign n435 = x129 & n434 ;
  assign n436 = n435 ^ n434 ;
  assign n442 = n441 ^ n436 ;
  assign n443 = n170 & n442 ;
  assign n425 = x61 & x128 ;
  assign n423 = x62 & x128 ;
  assign n424 = n423 ^ x62 ;
  assign n426 = n425 ^ n424 ;
  assign n427 = x129 & n426 ;
  assign n419 = x63 & x128 ;
  assign n417 = x64 & x128 ;
  assign n418 = n417 ^ x64 ;
  assign n420 = n419 ^ n418 ;
  assign n421 = x129 & n420 ;
  assign n422 = n421 ^ n420 ;
  assign n428 = n427 ^ n422 ;
  assign n429 = n171 & n428 ;
  assign n430 = n429 ^ n428 ;
  assign n444 = n443 ^ n430 ;
  assign n466 = x53 & x128 ;
  assign n464 = x54 & x128 ;
  assign n465 = n464 ^ x54 ;
  assign n467 = n466 ^ n465 ;
  assign n468 = x129 & n467 ;
  assign n460 = x55 & x128 ;
  assign n458 = x56 & x128 ;
  assign n459 = n458 ^ x56 ;
  assign n461 = n460 ^ n459 ;
  assign n462 = x129 & n461 ;
  assign n463 = n462 ^ n461 ;
  assign n469 = n468 ^ n463 ;
  assign n470 = n155 & n469 ;
  assign n453 = x49 & x128 ;
  assign n451 = x50 & x128 ;
  assign n452 = n451 ^ x50 ;
  assign n454 = n453 ^ n452 ;
  assign n455 = x129 & n454 ;
  assign n447 = x51 & x128 ;
  assign n445 = x52 & x128 ;
  assign n446 = n445 ^ x52 ;
  assign n448 = n447 ^ n446 ;
  assign n449 = x129 & n448 ;
  assign n450 = n449 ^ n448 ;
  assign n456 = n455 ^ n450 ;
  assign n457 = n139 & n456 ;
  assign n471 = n470 ^ n457 ;
  assign n472 = n444 & n471 ;
  assign n473 = n472 ^ n444 ;
  assign n474 = n473 ^ n471 ;
  assign n475 = n138 & n474 ;
  assign n476 = n475 ^ n474 ;
  assign n477 = n476 ^ n138 ;
  assign n549 = n548 ^ n477 ;
  assign n635 = x9 & x128 ;
  assign n633 = x10 & x128 ;
  assign n634 = n633 ^ x10 ;
  assign n636 = n635 ^ n634 ;
  assign n637 = x129 & n636 ;
  assign n629 = x11 & x128 ;
  assign n627 = x12 & x128 ;
  assign n628 = n627 ^ x12 ;
  assign n630 = n629 ^ n628 ;
  assign n631 = x129 & n630 ;
  assign n632 = n631 ^ n630 ;
  assign n638 = n637 ^ n632 ;
  assign n639 = n170 & n638 ;
  assign n640 = n639 ^ n170 ;
  assign n641 = n640 ^ n170 ;
  assign n621 = x13 & x128 ;
  assign n619 = x14 & x128 ;
  assign n620 = n619 ^ x14 ;
  assign n622 = n621 ^ n620 ;
  assign n623 = x129 & n622 ;
  assign n615 = x15 & x128 ;
  assign n613 = x16 & x128 ;
  assign n614 = n613 ^ x16 ;
  assign n616 = n615 ^ n614 ;
  assign n617 = x129 & n616 ;
  assign n618 = n617 ^ n616 ;
  assign n624 = n623 ^ n618 ;
  assign n625 = n171 & n624 ;
  assign n626 = n625 ^ n624 ;
  assign n642 = n641 ^ n626 ;
  assign n664 = x5 & x128 ;
  assign n662 = x6 & x128 ;
  assign n663 = n662 ^ x6 ;
  assign n665 = n664 ^ n663 ;
  assign n666 = x129 & n665 ;
  assign n658 = x7 & x128 ;
  assign n656 = x8 & x128 ;
  assign n657 = n656 ^ x8 ;
  assign n659 = n658 ^ n657 ;
  assign n660 = x129 & n659 ;
  assign n661 = n660 ^ n659 ;
  assign n667 = n666 ^ n661 ;
  assign n668 = n155 & n667 ;
  assign n651 = x1 & x128 ;
  assign n649 = x2 & x128 ;
  assign n650 = n649 ^ x2 ;
  assign n652 = n651 ^ n650 ;
  assign n653 = x129 & n652 ;
  assign n645 = x3 & x128 ;
  assign n643 = x4 & x128 ;
  assign n644 = n643 ^ x4 ;
  assign n646 = n645 ^ n644 ;
  assign n647 = x129 & n646 ;
  assign n648 = n647 ^ n646 ;
  assign n654 = n653 ^ n648 ;
  assign n655 = n139 & n654 ;
  assign n669 = n668 ^ n655 ;
  assign n670 = n642 & n669 ;
  assign n671 = n670 ^ n669 ;
  assign n672 = n671 ^ n642 ;
  assign n673 = n136 & n672 ;
  assign n674 = n549 & n673 ;
  assign n675 = n674 ^ n673 ;
  assign n676 = n675 ^ n549 ;
  assign n402 = n136 ^ x133 ;
  assign n572 = x25 & x128 ;
  assign n570 = x26 & x128 ;
  assign n571 = n570 ^ x26 ;
  assign n573 = n572 ^ n571 ;
  assign n574 = x129 & n573 ;
  assign n566 = x27 & x128 ;
  assign n564 = x28 & x128 ;
  assign n565 = n564 ^ x28 ;
  assign n567 = n566 ^ n565 ;
  assign n568 = x129 & n567 ;
  assign n569 = n568 ^ n567 ;
  assign n575 = n574 ^ n569 ;
  assign n576 = n170 & n575 ;
  assign n558 = x29 & x128 ;
  assign n556 = x30 & x128 ;
  assign n557 = n556 ^ x30 ;
  assign n559 = n558 ^ n557 ;
  assign n560 = x129 & n559 ;
  assign n552 = x31 & x128 ;
  assign n550 = x32 & x128 ;
  assign n551 = n550 ^ x32 ;
  assign n553 = n552 ^ n551 ;
  assign n554 = x129 & n553 ;
  assign n555 = n554 ^ n553 ;
  assign n561 = n560 ^ n555 ;
  assign n562 = n171 & n561 ;
  assign n563 = n562 ^ n561 ;
  assign n577 = n576 ^ n563 ;
  assign n599 = x21 & x128 ;
  assign n597 = x22 & x128 ;
  assign n598 = n597 ^ x22 ;
  assign n600 = n599 ^ n598 ;
  assign n601 = x129 & n600 ;
  assign n593 = x23 & x128 ;
  assign n591 = x24 & x128 ;
  assign n592 = n591 ^ x24 ;
  assign n594 = n593 ^ n592 ;
  assign n595 = x129 & n594 ;
  assign n596 = n595 ^ n594 ;
  assign n602 = n601 ^ n596 ;
  assign n603 = n155 & n602 ;
  assign n586 = x17 & x128 ;
  assign n584 = x18 & x128 ;
  assign n585 = n584 ^ x18 ;
  assign n587 = n586 ^ n585 ;
  assign n588 = x129 & n587 ;
  assign n580 = x19 & x128 ;
  assign n578 = x20 & x128 ;
  assign n579 = n578 ^ x20 ;
  assign n581 = n580 ^ n579 ;
  assign n582 = x129 & n581 ;
  assign n583 = n582 ^ n581 ;
  assign n589 = n588 ^ n583 ;
  assign n590 = n139 & n589 ;
  assign n604 = n603 ^ n590 ;
  assign n605 = n577 & n604 ;
  assign n606 = n605 ^ n577 ;
  assign n607 = n606 ^ n604 ;
  assign n608 = n402 & n607 ;
  assign n609 = n608 ^ n402 ;
  assign n610 = n609 ^ n402 ;
  assign n611 = n549 & n610 ;
  assign n612 = n611 ^ n610 ;
  assign n677 = n676 ^ n612 ;
  assign n678 = x134 & n677 ;
  assign n679 = n678 ^ x134 ;
  assign n366 = x89 & x128 ;
  assign n364 = x90 & x128 ;
  assign n365 = n364 ^ x90 ;
  assign n367 = n366 ^ n365 ;
  assign n368 = x129 & n367 ;
  assign n360 = x91 & x128 ;
  assign n358 = x92 & x128 ;
  assign n359 = n358 ^ x92 ;
  assign n361 = n360 ^ n359 ;
  assign n362 = x129 & n361 ;
  assign n363 = n362 ^ n361 ;
  assign n369 = n368 ^ n363 ;
  assign n370 = n170 & n369 ;
  assign n353 = x93 & x128 ;
  assign n351 = x94 & x128 ;
  assign n352 = n351 ^ x94 ;
  assign n354 = n353 ^ n352 ;
  assign n355 = x129 & n354 ;
  assign n347 = x95 & x128 ;
  assign n345 = x96 & x128 ;
  assign n346 = n345 ^ x96 ;
  assign n348 = n347 ^ n346 ;
  assign n349 = x129 & n348 ;
  assign n350 = n349 ^ n348 ;
  assign n356 = n355 ^ n350 ;
  assign n357 = ~n171 & n356 ;
  assign n371 = n370 ^ n357 ;
  assign n393 = x85 & x128 ;
  assign n391 = x86 & x128 ;
  assign n392 = n391 ^ x86 ;
  assign n394 = n393 ^ n392 ;
  assign n395 = x129 & n394 ;
  assign n387 = x87 & x128 ;
  assign n385 = x88 & x128 ;
  assign n386 = n385 ^ x88 ;
  assign n388 = n387 ^ n386 ;
  assign n389 = x129 & n388 ;
  assign n390 = n389 ^ n388 ;
  assign n396 = n395 ^ n390 ;
  assign n397 = n155 & n396 ;
  assign n380 = x81 & x128 ;
  assign n378 = x82 & x128 ;
  assign n379 = n378 ^ x82 ;
  assign n381 = n380 ^ n379 ;
  assign n382 = x129 & n381 ;
  assign n374 = x83 & x128 ;
  assign n372 = x84 & x128 ;
  assign n373 = n372 ^ x84 ;
  assign n375 = n374 ^ n373 ;
  assign n376 = x129 & n375 ;
  assign n377 = n376 ^ n375 ;
  assign n383 = n382 ^ n377 ;
  assign n384 = n139 & n383 ;
  assign n398 = n397 ^ n384 ;
  assign n399 = ~n371 & ~n398 ;
  assign n680 = n679 ^ n399 ;
  assign n681 = n680 ^ x134 ;
  assign n231 = x105 & x128 ;
  assign n229 = x106 & x128 ;
  assign n230 = n229 ^ x106 ;
  assign n232 = n231 ^ n230 ;
  assign n233 = x129 & n232 ;
  assign n225 = x107 & x128 ;
  assign n223 = x108 & x128 ;
  assign n224 = n223 ^ x108 ;
  assign n226 = n225 ^ n224 ;
  assign n227 = x129 & n226 ;
  assign n228 = n227 ^ n226 ;
  assign n234 = n233 ^ n228 ;
  assign n235 = n170 & n234 ;
  assign n236 = n235 ^ n170 ;
  assign n237 = n236 ^ n170 ;
  assign n215 = x109 & x128 ;
  assign n213 = x110 & x128 ;
  assign n214 = n213 ^ x110 ;
  assign n216 = n215 ^ n214 ;
  assign n217 = x129 & n216 ;
  assign n209 = x111 & x128 ;
  assign n207 = x112 & x128 ;
  assign n208 = n207 ^ x112 ;
  assign n210 = n209 ^ n208 ;
  assign n211 = x129 & n210 ;
  assign n212 = n211 ^ n210 ;
  assign n218 = n217 ^ n212 ;
  assign n219 = n171 & n218 ;
  assign n220 = n219 ^ n218 ;
  assign n221 = n220 ^ n171 ;
  assign n222 = n221 ^ n171 ;
  assign n238 = n237 ^ n222 ;
  assign n262 = x101 & x128 ;
  assign n260 = x102 & x128 ;
  assign n261 = n260 ^ x102 ;
  assign n263 = n262 ^ n261 ;
  assign n264 = x129 & n263 ;
  assign n256 = x103 & x128 ;
  assign n254 = x104 & x128 ;
  assign n255 = n254 ^ x104 ;
  assign n257 = n256 ^ n255 ;
  assign n258 = x129 & n257 ;
  assign n259 = n258 ^ n257 ;
  assign n265 = n264 ^ n259 ;
  assign n266 = n155 & n265 ;
  assign n267 = n266 ^ n155 ;
  assign n268 = n267 ^ n155 ;
  assign n247 = x97 & x128 ;
  assign n245 = x98 & x128 ;
  assign n246 = n245 ^ x98 ;
  assign n248 = n247 ^ n246 ;
  assign n249 = x129 & n248 ;
  assign n241 = x99 & x128 ;
  assign n239 = x100 & x128 ;
  assign n240 = n239 ^ x100 ;
  assign n242 = n241 ^ n240 ;
  assign n243 = x129 & n242 ;
  assign n244 = n243 ^ n242 ;
  assign n250 = n249 ^ n244 ;
  assign n251 = n139 & n250 ;
  assign n252 = n251 ^ n139 ;
  assign n253 = n252 ^ n139 ;
  assign n269 = n268 ^ n253 ;
  assign n270 = n238 & n269 ;
  assign n271 = n270 ^ n238 ;
  assign n272 = n271 ^ n269 ;
  assign n273 = n137 & n272 ;
  assign n274 = n273 ^ n137 ;
  assign n275 = n274 ^ n137 ;
  assign n164 = x117 & x128 ;
  assign n162 = x118 & x128 ;
  assign n163 = n162 ^ x118 ;
  assign n165 = n164 ^ n163 ;
  assign n166 = x129 & n165 ;
  assign n158 = x119 & x128 ;
  assign n156 = x120 & x128 ;
  assign n157 = n156 ^ x120 ;
  assign n159 = n158 ^ n157 ;
  assign n160 = x129 & n159 ;
  assign n161 = n160 ^ n159 ;
  assign n167 = n166 ^ n161 ;
  assign n168 = n155 & n167 ;
  assign n148 = x113 & x128 ;
  assign n146 = x114 & x128 ;
  assign n147 = n146 ^ x114 ;
  assign n149 = n148 ^ n147 ;
  assign n150 = x129 & n149 ;
  assign n142 = x115 & x128 ;
  assign n140 = x116 & x128 ;
  assign n141 = n140 ^ x116 ;
  assign n143 = n142 ^ n141 ;
  assign n144 = x129 & n143 ;
  assign n145 = n144 ^ n143 ;
  assign n151 = n150 ^ n145 ;
  assign n152 = n139 & n151 ;
  assign n153 = n152 ^ n139 ;
  assign n154 = n153 ^ n139 ;
  assign n169 = n168 ^ n154 ;
  assign n194 = x121 & x128 ;
  assign n192 = x122 & x128 ;
  assign n193 = n192 ^ x122 ;
  assign n195 = n194 ^ n193 ;
  assign n196 = x129 & n195 ;
  assign n188 = x123 & x128 ;
  assign n186 = x124 & x128 ;
  assign n187 = n186 ^ x124 ;
  assign n189 = n188 ^ n187 ;
  assign n190 = x129 & n189 ;
  assign n191 = n190 ^ n189 ;
  assign n197 = n196 ^ n191 ;
  assign n198 = n170 & n197 ;
  assign n180 = x125 & x128 ;
  assign n178 = x126 & x128 ;
  assign n179 = n178 ^ x126 ;
  assign n181 = n180 ^ n179 ;
  assign n182 = x129 & n181 ;
  assign n173 = x0 & x128 ;
  assign n174 = n173 ^ x0 ;
  assign n172 = x127 & x128 ;
  assign n175 = n174 ^ n172 ;
  assign n176 = x129 & n175 ;
  assign n177 = n176 ^ n175 ;
  assign n183 = n182 ^ n177 ;
  assign n184 = n171 & n183 ;
  assign n185 = n184 ^ n183 ;
  assign n199 = n198 ^ n185 ;
  assign n200 = n169 & n199 ;
  assign n201 = n200 ^ n199 ;
  assign n202 = n201 ^ n169 ;
  assign n203 = n138 & n202 ;
  assign n204 = n203 ^ n202 ;
  assign n205 = n204 ^ n138 ;
  assign n206 = n205 ^ n138 ;
  assign n276 = n275 ^ n206 ;
  assign n400 = n399 ^ n276 ;
  assign n401 = n400 ^ x134 ;
  assign n403 = n402 ^ n276 ;
  assign n404 = n403 ^ x134 ;
  assign n405 = x134 & ~n402 ;
  assign n406 = n405 ^ n402 ;
  assign n407 = n406 ^ x134 ;
  assign n408 = n404 & n407 ;
  assign n409 = n408 ^ n404 ;
  assign n410 = n409 ^ n407 ;
  assign n411 = n410 ^ n405 ;
  assign n412 = n411 ^ n276 ;
  assign n413 = n401 & n412 ;
  assign n414 = n413 ^ n401 ;
  assign n415 = n414 ^ n410 ;
  assign n416 = n415 ^ n405 ;
  assign n682 = n681 ^ n416 ;
  assign n277 = x134 & n276 ;
  assign n278 = n277 ^ x134 ;
  assign n279 = n278 ^ n276 ;
  assign n301 = x69 & x128 ;
  assign n299 = x70 & x128 ;
  assign n300 = n299 ^ x70 ;
  assign n302 = n301 ^ n300 ;
  assign n303 = x129 & n302 ;
  assign n295 = x71 & x128 ;
  assign n293 = x72 & x128 ;
  assign n294 = n293 ^ x72 ;
  assign n296 = n295 ^ n294 ;
  assign n297 = x129 & n296 ;
  assign n298 = n297 ^ n296 ;
  assign n304 = n303 ^ n298 ;
  assign n305 = n155 & n304 ;
  assign n306 = n305 ^ n155 ;
  assign n307 = n306 ^ n155 ;
  assign n288 = x65 & x128 ;
  assign n286 = x66 & x128 ;
  assign n287 = n286 ^ x66 ;
  assign n289 = n288 ^ n287 ;
  assign n290 = x129 & n289 ;
  assign n282 = x67 & x128 ;
  assign n280 = x68 & x128 ;
  assign n281 = n280 ^ x68 ;
  assign n283 = n282 ^ n281 ;
  assign n284 = x129 & n283 ;
  assign n285 = n284 ^ n283 ;
  assign n291 = n290 ^ n285 ;
  assign n292 = n139 & n291 ;
  assign n308 = n307 ^ n292 ;
  assign n331 = x73 & x128 ;
  assign n329 = x74 & x128 ;
  assign n330 = n329 ^ x74 ;
  assign n332 = n331 ^ n330 ;
  assign n333 = x129 & n332 ;
  assign n325 = x75 & x128 ;
  assign n323 = x76 & x128 ;
  assign n324 = n323 ^ x76 ;
  assign n326 = n325 ^ n324 ;
  assign n327 = x129 & n326 ;
  assign n328 = n327 ^ n326 ;
  assign n334 = n333 ^ n328 ;
  assign n335 = n170 & n334 ;
  assign n317 = x77 & x128 ;
  assign n315 = x78 & x128 ;
  assign n316 = n315 ^ x78 ;
  assign n318 = n317 ^ n316 ;
  assign n319 = x129 & n318 ;
  assign n311 = x79 & x128 ;
  assign n309 = x80 & x128 ;
  assign n310 = n309 ^ x80 ;
  assign n312 = n311 ^ n310 ;
  assign n313 = x129 & n312 ;
  assign n314 = n313 ^ n312 ;
  assign n320 = n319 ^ n314 ;
  assign n321 = n171 & n320 ;
  assign n322 = n321 ^ n320 ;
  assign n336 = n335 ^ n322 ;
  assign n337 = n308 & n336 ;
  assign n338 = n337 ^ n336 ;
  assign n339 = n338 ^ n308 ;
  assign n340 = n136 & ~n339 ;
  assign n341 = n340 ^ n136 ;
  assign n342 = n279 & n341 ;
  assign n343 = n342 ^ n341 ;
  assign n344 = n343 ^ n279 ;
  assign n683 = n682 ^ n344 ;
  assign n789 = n225 ^ x107 ;
  assign n790 = x129 & n789 ;
  assign n787 = x129 & n223 ;
  assign n788 = n787 ^ n223 ;
  assign n791 = n790 ^ n788 ;
  assign n796 = x129 & n229 ;
  assign n797 = n796 ^ x129 ;
  assign n792 = n215 ^ x109 ;
  assign n793 = x129 & n792 ;
  assign n794 = n793 ^ x129 ;
  assign n795 = n794 ^ n792 ;
  assign n798 = n797 ^ n795 ;
  assign n799 = n791 & n798 ;
  assign n800 = n799 ^ n791 ;
  assign n801 = n800 ^ n798 ;
  assign n802 = n170 & n801 ;
  assign n803 = n802 ^ n170 ;
  assign n804 = n803 ^ n170 ;
  assign n770 = n209 ^ x111 ;
  assign n771 = x129 & n770 ;
  assign n768 = x129 & n207 ;
  assign n769 = n768 ^ n207 ;
  assign n772 = n771 ^ n769 ;
  assign n777 = x129 & n213 ;
  assign n778 = n777 ^ x129 ;
  assign n773 = n148 ^ x113 ;
  assign n774 = x129 & n773 ;
  assign n775 = n774 ^ x129 ;
  assign n776 = n775 ^ n773 ;
  assign n779 = n778 ^ n776 ;
  assign n780 = n772 & n779 ;
  assign n781 = n780 ^ n772 ;
  assign n782 = n781 ^ n779 ;
  assign n783 = n171 & n782 ;
  assign n784 = n783 ^ n171 ;
  assign n785 = n784 ^ n782 ;
  assign n786 = n785 ^ n171 ;
  assign n805 = n804 ^ n786 ;
  assign n824 = n256 ^ x103 ;
  assign n825 = x129 & n824 ;
  assign n822 = x129 & n254 ;
  assign n823 = n822 ^ n254 ;
  assign n826 = n825 ^ n823 ;
  assign n831 = x129 & n260 ;
  assign n832 = n831 ^ x129 ;
  assign n827 = n231 ^ x105 ;
  assign n828 = x129 & n827 ;
  assign n829 = n828 ^ x129 ;
  assign n830 = n829 ^ n827 ;
  assign n833 = n832 ^ n830 ;
  assign n834 = n826 & n833 ;
  assign n835 = n834 ^ n826 ;
  assign n836 = n835 ^ n833 ;
  assign n837 = n155 & n836 ;
  assign n838 = n837 ^ n155 ;
  assign n839 = n838 ^ n155 ;
  assign n808 = n241 ^ x99 ;
  assign n809 = x129 & n808 ;
  assign n806 = x129 & n239 ;
  assign n807 = n806 ^ n239 ;
  assign n810 = n809 ^ n807 ;
  assign n815 = x129 & n245 ;
  assign n816 = n815 ^ x129 ;
  assign n811 = n262 ^ x101 ;
  assign n812 = x129 & n811 ;
  assign n813 = n812 ^ x129 ;
  assign n814 = n813 ^ n811 ;
  assign n817 = n816 ^ n814 ;
  assign n818 = n810 & n817 ;
  assign n819 = n818 ^ n810 ;
  assign n820 = n819 ^ n817 ;
  assign n821 = n139 & n820 ;
  assign n840 = n839 ^ n821 ;
  assign n841 = n805 & n840 ;
  assign n842 = n841 ^ n840 ;
  assign n843 = n842 ^ n840 ;
  assign n844 = n843 ^ n805 ;
  assign n845 = n844 ^ n840 ;
  assign n846 = n137 & n845 ;
  assign n847 = n846 ^ n137 ;
  assign n848 = n847 ^ n137 ;
  assign n705 = n188 ^ x123 ;
  assign n706 = x129 & n705 ;
  assign n703 = x129 & n186 ;
  assign n704 = n703 ^ n186 ;
  assign n707 = n706 ^ n704 ;
  assign n712 = x129 & n192 ;
  assign n713 = n712 ^ x129 ;
  assign n708 = n180 ^ x125 ;
  assign n709 = x129 & n708 ;
  assign n710 = n709 ^ x129 ;
  assign n711 = n710 ^ n708 ;
  assign n714 = n713 ^ n711 ;
  assign n715 = n707 & n714 ;
  assign n716 = n715 ^ n707 ;
  assign n717 = n716 ^ n714 ;
  assign n718 = n170 & n717 ;
  assign n719 = n718 ^ n170 ;
  assign n720 = n719 ^ n170 ;
  assign n686 = n172 ^ x127 ;
  assign n687 = x129 & n686 ;
  assign n684 = x129 & n173 ;
  assign n685 = n684 ^ n173 ;
  assign n688 = n687 ^ n685 ;
  assign n693 = x129 & n178 ;
  assign n694 = n693 ^ x129 ;
  assign n689 = n651 ^ x1 ;
  assign n690 = x129 & n689 ;
  assign n691 = n690 ^ x129 ;
  assign n692 = n691 ^ n689 ;
  assign n695 = n694 ^ n692 ;
  assign n696 = n688 & n695 ;
  assign n697 = n696 ^ n688 ;
  assign n698 = n697 ^ n695 ;
  assign n699 = n171 & n698 ;
  assign n700 = n699 ^ n171 ;
  assign n701 = n700 ^ n698 ;
  assign n702 = n701 ^ n171 ;
  assign n721 = n720 ^ n702 ;
  assign n742 = n158 ^ x119 ;
  assign n743 = x129 & n742 ;
  assign n740 = x129 & n156 ;
  assign n741 = n740 ^ n156 ;
  assign n744 = n743 ^ n741 ;
  assign n749 = x129 & n162 ;
  assign n750 = n749 ^ x129 ;
  assign n745 = n194 ^ x121 ;
  assign n746 = x129 & n745 ;
  assign n747 = n746 ^ x129 ;
  assign n748 = n747 ^ n745 ;
  assign n751 = n750 ^ n748 ;
  assign n752 = n744 & n751 ;
  assign n753 = n752 ^ n744 ;
  assign n754 = n753 ^ n751 ;
  assign n755 = n155 & n754 ;
  assign n756 = n755 ^ n155 ;
  assign n757 = n756 ^ n155 ;
  assign n724 = n142 ^ x115 ;
  assign n725 = x129 & n724 ;
  assign n722 = x129 & n140 ;
  assign n723 = n722 ^ n140 ;
  assign n726 = n725 ^ n723 ;
  assign n731 = x129 & n146 ;
  assign n732 = n731 ^ x129 ;
  assign n727 = n164 ^ x117 ;
  assign n728 = x129 & n727 ;
  assign n729 = n728 ^ x129 ;
  assign n730 = n729 ^ n727 ;
  assign n733 = n732 ^ n730 ;
  assign n734 = n726 & n733 ;
  assign n735 = n734 ^ n726 ;
  assign n736 = n735 ^ n733 ;
  assign n737 = n139 & n736 ;
  assign n738 = n737 ^ n139 ;
  assign n739 = n738 ^ n139 ;
  assign n758 = n757 ^ n739 ;
  assign n759 = n721 & n758 ;
  assign n760 = n759 ^ n758 ;
  assign n761 = n760 ^ n758 ;
  assign n762 = n761 ^ n721 ;
  assign n763 = n762 ^ n758 ;
  assign n764 = n138 & n763 ;
  assign n765 = n764 ^ n138 ;
  assign n766 = n765 ^ n763 ;
  assign n767 = n766 ^ n138 ;
  assign n849 = n848 ^ n767 ;
  assign n1259 = ~x134 & n402 ;
  assign n1279 = n360 ^ x91 ;
  assign n1280 = x129 & n1279 ;
  assign n1277 = x129 & n358 ;
  assign n1278 = n1277 ^ n358 ;
  assign n1281 = n1280 ^ n1278 ;
  assign n1286 = x129 & n364 ;
  assign n1287 = n1286 ^ x129 ;
  assign n1282 = n353 ^ x93 ;
  assign n1283 = x129 & n1282 ;
  assign n1284 = n1283 ^ x129 ;
  assign n1285 = n1284 ^ n1282 ;
  assign n1288 = n1287 ^ n1285 ;
  assign n1289 = n1281 & n1288 ;
  assign n1290 = n1289 ^ n1281 ;
  assign n1291 = n1290 ^ n1288 ;
  assign n1292 = n170 & n1291 ;
  assign n1262 = n347 ^ x95 ;
  assign n1263 = x129 & n1262 ;
  assign n1260 = x129 & n345 ;
  assign n1261 = n1260 ^ n345 ;
  assign n1264 = n1263 ^ n1261 ;
  assign n1269 = x129 & n351 ;
  assign n1270 = n1269 ^ x129 ;
  assign n1265 = n247 ^ x97 ;
  assign n1266 = x129 & n1265 ;
  assign n1267 = n1266 ^ x129 ;
  assign n1268 = n1267 ^ n1265 ;
  assign n1271 = n1270 ^ n1268 ;
  assign n1272 = n1264 & n1271 ;
  assign n1273 = n1272 ^ n1264 ;
  assign n1274 = n1273 ^ n1271 ;
  assign n1275 = n171 & n1274 ;
  assign n1276 = n1275 ^ n1274 ;
  assign n1293 = n1292 ^ n1276 ;
  assign n1314 = n387 ^ x87 ;
  assign n1315 = x129 & n1314 ;
  assign n1312 = x129 & n385 ;
  assign n1313 = n1312 ^ n385 ;
  assign n1316 = n1315 ^ n1313 ;
  assign n1321 = x129 & n391 ;
  assign n1322 = n1321 ^ x129 ;
  assign n1317 = n366 ^ x89 ;
  assign n1318 = x129 & n1317 ;
  assign n1319 = n1318 ^ x129 ;
  assign n1320 = n1319 ^ n1317 ;
  assign n1323 = n1322 ^ n1320 ;
  assign n1324 = n1316 & n1323 ;
  assign n1325 = n1324 ^ n1316 ;
  assign n1326 = n1325 ^ n1323 ;
  assign n1327 = n155 & n1326 ;
  assign n1296 = n374 ^ x83 ;
  assign n1297 = x129 & n1296 ;
  assign n1294 = x129 & n372 ;
  assign n1295 = n1294 ^ n372 ;
  assign n1298 = n1297 ^ n1295 ;
  assign n1303 = x129 & n378 ;
  assign n1304 = n1303 ^ x129 ;
  assign n1299 = n393 ^ x85 ;
  assign n1300 = x129 & n1299 ;
  assign n1301 = n1300 ^ x129 ;
  assign n1302 = n1301 ^ n1299 ;
  assign n1305 = n1304 ^ n1302 ;
  assign n1306 = n1298 & n1305 ;
  assign n1307 = n1306 ^ n1298 ;
  assign n1308 = n1307 ^ n1305 ;
  assign n1309 = n139 & n1308 ;
  assign n1310 = n1309 ^ n139 ;
  assign n1311 = n1310 ^ n139 ;
  assign n1328 = n1327 ^ n1311 ;
  assign n1329 = n1293 & n1328 ;
  assign n1330 = n1329 ^ n1293 ;
  assign n1331 = n1330 ^ n1328 ;
  assign n1332 = n1259 & n1331 ;
  assign n1333 = ~n849 & n1332 ;
  assign n1334 = n1333 ^ n1332 ;
  assign n1335 = n1334 ^ n1332 ;
  assign n973 = n593 ^ x23 ;
  assign n974 = x129 & n973 ;
  assign n971 = x129 & n591 ;
  assign n972 = n971 ^ n591 ;
  assign n975 = n974 ^ n972 ;
  assign n980 = x129 & n597 ;
  assign n981 = n980 ^ x129 ;
  assign n976 = n572 ^ x25 ;
  assign n977 = x129 & n976 ;
  assign n978 = n977 ^ x129 ;
  assign n979 = n978 ^ n976 ;
  assign n982 = n981 ^ n979 ;
  assign n983 = n975 & n982 ;
  assign n984 = n983 ^ n975 ;
  assign n985 = n984 ^ n982 ;
  assign n986 = n155 & n985 ;
  assign n957 = n580 ^ x19 ;
  assign n958 = x129 & n957 ;
  assign n955 = x129 & n578 ;
  assign n956 = n955 ^ n578 ;
  assign n959 = n958 ^ n956 ;
  assign n964 = x129 & n584 ;
  assign n965 = n964 ^ x129 ;
  assign n960 = n599 ^ x21 ;
  assign n961 = x129 & n960 ;
  assign n962 = n961 ^ x129 ;
  assign n963 = n962 ^ n960 ;
  assign n966 = n965 ^ n963 ;
  assign n967 = n959 & n966 ;
  assign n968 = n967 ^ n959 ;
  assign n969 = n968 ^ n966 ;
  assign n970 = n139 & n969 ;
  assign n987 = n986 ^ n970 ;
  assign n1081 = n552 ^ x31 ;
  assign n1082 = x129 & n1081 ;
  assign n1079 = x129 & n550 ;
  assign n1080 = n1079 ^ n550 ;
  assign n1083 = n1082 ^ n1080 ;
  assign n1088 = x129 & n556 ;
  assign n1089 = n1088 ^ x129 ;
  assign n1084 = n517 ^ x33 ;
  assign n1085 = x129 & n1084 ;
  assign n1086 = n1085 ^ x129 ;
  assign n1087 = n1086 ^ n1084 ;
  assign n1090 = n1089 ^ n1087 ;
  assign n1091 = n1083 & n1090 ;
  assign n1092 = n1091 ^ n1083 ;
  assign n1093 = n1092 ^ n1090 ;
  assign n1094 = ~n171 & n402 ;
  assign n1095 = n1093 & n1094 ;
  assign n1096 = n987 & n1095 ;
  assign n1097 = n1096 ^ n1095 ;
  assign n1038 = ~x129 & n139 ;
  assign n1039 = n509 & n1038 ;
  assign n1032 = n526 ^ x128 ;
  assign n1030 = n523 ^ x39 ;
  assign n1031 = n1030 ^ x128 ;
  assign n1033 = n1032 ^ n1031 ;
  assign n1034 = x129 & n1033 ;
  assign n1035 = n1034 ^ x129 ;
  assign n1025 = n530 ^ x128 ;
  assign n1023 = n486 ^ x41 ;
  assign n1024 = n1023 ^ x128 ;
  assign n1026 = n1025 ^ n1024 ;
  assign n1027 = x129 & n1026 ;
  assign n1028 = n1027 ^ x129 ;
  assign n1029 = n1028 ^ n1026 ;
  assign n1036 = n1035 ^ n1029 ;
  assign n1037 = n155 & n1036 ;
  assign n1040 = n1039 ^ n1037 ;
  assign n1013 = x129 & n515 ;
  assign n1014 = n1013 ^ x129 ;
  assign n1009 = n535 ^ x37 ;
  assign n1010 = x129 & n1009 ;
  assign n1011 = n1010 ^ x129 ;
  assign n1012 = n1011 ^ n1009 ;
  assign n1015 = n1014 ^ n1012 ;
  assign n1016 = n511 ^ x35 ;
  assign n1017 = x129 & n1016 ;
  assign n1018 = n139 & n1017 ;
  assign n1019 = n1018 ^ n139 ;
  assign n1020 = n1015 & n1019 ;
  assign n1021 = n1020 ^ n1019 ;
  assign n1022 = n1021 ^ n139 ;
  assign n1041 = n1040 ^ n1022 ;
  assign n1042 = x129 & n171 ;
  assign n1043 = n1042 ^ x129 ;
  assign n1044 = n1043 ^ n171 ;
  assign n1072 = n492 & n1044 ;
  assign n1073 = n1072 ^ n492 ;
  assign n1066 = n484 ^ x128 ;
  assign n1064 = n480 ^ x43 ;
  assign n1065 = n1064 ^ x128 ;
  assign n1067 = n1066 ^ n1065 ;
  assign n1068 = x129 & n1067 ;
  assign n1069 = n1068 ^ x129 ;
  assign n1059 = n500 ^ x45 ;
  assign n1060 = n1059 ^ n478 ;
  assign n1061 = x129 & n1060 ;
  assign n1062 = n1061 ^ x129 ;
  assign n1063 = n1062 ^ n1060 ;
  assign n1070 = n1069 ^ n1063 ;
  assign n1071 = n170 & n1070 ;
  assign n1074 = n1073 ^ n1071 ;
  assign n1049 = x129 & n498 ;
  assign n1050 = n1049 ^ x129 ;
  assign n1051 = n494 ^ x47 ;
  assign n1052 = n171 & n1051 ;
  assign n1053 = n1052 ^ n171 ;
  assign n1054 = n1053 ^ n1051 ;
  assign n1055 = n1050 & n1054 ;
  assign n1056 = n1055 ^ n1050 ;
  assign n1045 = n453 ^ x49 ;
  assign n1046 = n1044 & n1045 ;
  assign n1047 = n1046 ^ n1045 ;
  assign n1048 = n1047 ^ n1044 ;
  assign n1057 = n1056 ^ n1048 ;
  assign n1058 = n1057 ^ n171 ;
  assign n1075 = n1074 ^ n1058 ;
  assign n1076 = n137 & ~n1075 ;
  assign n1077 = ~n1041 & n1076 ;
  assign n1078 = n1077 ^ n137 ;
  assign n1098 = n1097 ^ n1078 ;
  assign n990 = n566 ^ x27 ;
  assign n991 = x129 & n990 ;
  assign n988 = x129 & n564 ;
  assign n989 = n988 ^ n564 ;
  assign n992 = n991 ^ n989 ;
  assign n997 = x129 & n570 ;
  assign n998 = n997 ^ x129 ;
  assign n993 = n558 ^ x29 ;
  assign n994 = x129 & n993 ;
  assign n995 = n994 ^ x129 ;
  assign n996 = n995 ^ n993 ;
  assign n999 = n998 ^ n996 ;
  assign n1000 = n992 & n999 ;
  assign n1001 = n1000 ^ n992 ;
  assign n1002 = n1001 ^ n999 ;
  assign n1003 = n170 & n402 ;
  assign n1004 = n1002 & n1003 ;
  assign n1005 = n1004 ^ n402 ;
  assign n1006 = n987 & n1005 ;
  assign n1007 = n1006 ^ n1005 ;
  assign n1008 = n1007 ^ n402 ;
  assign n1099 = n1098 ^ n1008 ;
  assign n1180 = x134 & n136 ;
  assign n1200 = n629 ^ x11 ;
  assign n1201 = x129 & n1200 ;
  assign n1198 = x129 & n627 ;
  assign n1199 = n1198 ^ n627 ;
  assign n1202 = n1201 ^ n1199 ;
  assign n1207 = x129 & n633 ;
  assign n1208 = n1207 ^ x129 ;
  assign n1203 = n621 ^ x13 ;
  assign n1204 = x129 & n1203 ;
  assign n1205 = n1204 ^ x129 ;
  assign n1206 = n1205 ^ n1203 ;
  assign n1209 = n1208 ^ n1206 ;
  assign n1210 = n1202 & n1209 ;
  assign n1211 = n1210 ^ n1202 ;
  assign n1212 = n1211 ^ n1209 ;
  assign n1213 = n170 & n1212 ;
  assign n1183 = n615 ^ x15 ;
  assign n1184 = x129 & n1183 ;
  assign n1181 = x129 & n613 ;
  assign n1182 = n1181 ^ n613 ;
  assign n1185 = n1184 ^ n1182 ;
  assign n1190 = x129 & n619 ;
  assign n1191 = n1190 ^ x129 ;
  assign n1186 = n586 ^ x17 ;
  assign n1187 = x129 & n1186 ;
  assign n1188 = n1187 ^ x129 ;
  assign n1189 = n1188 ^ n1186 ;
  assign n1192 = n1191 ^ n1189 ;
  assign n1193 = n1185 & n1192 ;
  assign n1194 = n1193 ^ n1185 ;
  assign n1195 = n1194 ^ n1192 ;
  assign n1196 = n171 & n1195 ;
  assign n1197 = n1196 ^ n1195 ;
  assign n1214 = n1213 ^ n1197 ;
  assign n1235 = n658 ^ x7 ;
  assign n1236 = x129 & n1235 ;
  assign n1233 = x129 & n656 ;
  assign n1234 = n1233 ^ n656 ;
  assign n1237 = n1236 ^ n1234 ;
  assign n1242 = x129 & n662 ;
  assign n1243 = n1242 ^ x129 ;
  assign n1238 = n635 ^ x9 ;
  assign n1239 = x129 & n1238 ;
  assign n1240 = n1239 ^ x129 ;
  assign n1241 = n1240 ^ n1238 ;
  assign n1244 = n1243 ^ n1241 ;
  assign n1245 = n1237 & n1244 ;
  assign n1246 = n1245 ^ n1237 ;
  assign n1247 = n1246 ^ n1244 ;
  assign n1248 = n155 & n1247 ;
  assign n1249 = n1248 ^ n155 ;
  assign n1250 = n1249 ^ n155 ;
  assign n1217 = n645 ^ x3 ;
  assign n1218 = x129 & n1217 ;
  assign n1215 = x129 & n643 ;
  assign n1216 = n1215 ^ n643 ;
  assign n1219 = n1218 ^ n1216 ;
  assign n1224 = x129 & n649 ;
  assign n1225 = n1224 ^ x129 ;
  assign n1220 = n664 ^ x5 ;
  assign n1221 = x129 & n1220 ;
  assign n1222 = n1221 ^ x129 ;
  assign n1223 = n1222 ^ n1220 ;
  assign n1226 = n1225 ^ n1223 ;
  assign n1227 = n1219 & n1226 ;
  assign n1228 = n1227 ^ n1219 ;
  assign n1229 = n1228 ^ n1226 ;
  assign n1230 = n139 & n1229 ;
  assign n1231 = n1230 ^ n139 ;
  assign n1232 = n1231 ^ n139 ;
  assign n1251 = n1250 ^ n1232 ;
  assign n1252 = n1214 & n1251 ;
  assign n1253 = n1252 ^ n1214 ;
  assign n1254 = n1253 ^ n1251 ;
  assign n1255 = n1180 & n1254 ;
  assign n1256 = n1099 & n1255 ;
  assign n1257 = n1256 ^ n1255 ;
  assign n1157 = x130 & ~x131 ;
  assign n1160 = n433 ^ x59 ;
  assign n1161 = x129 & n1160 ;
  assign n1158 = x129 & n431 ;
  assign n1159 = n1158 ^ n431 ;
  assign n1162 = n1161 ^ n1159 ;
  assign n1167 = x129 & n437 ;
  assign n1168 = n1167 ^ x129 ;
  assign n1163 = n425 ^ x61 ;
  assign n1164 = x129 & n1163 ;
  assign n1165 = n1164 ^ x129 ;
  assign n1166 = n1165 ^ n1163 ;
  assign n1169 = n1168 ^ n1166 ;
  assign n1170 = n1162 & n1169 ;
  assign n1171 = n1170 ^ n1162 ;
  assign n1172 = n1171 ^ n1169 ;
  assign n1173 = n1157 & n1172 ;
  assign n1120 = n460 ^ x55 ;
  assign n1121 = x129 & n1120 ;
  assign n1118 = x129 & n458 ;
  assign n1119 = n1118 ^ n458 ;
  assign n1122 = n1121 ^ n1119 ;
  assign n1127 = x129 & n464 ;
  assign n1128 = n1127 ^ x129 ;
  assign n1123 = n439 ^ x57 ;
  assign n1124 = x129 & n1123 ;
  assign n1125 = n1124 ^ x129 ;
  assign n1126 = n1125 ^ n1123 ;
  assign n1129 = n1128 ^ n1126 ;
  assign n1130 = n1122 & n1129 ;
  assign n1131 = n1130 ^ n1122 ;
  assign n1132 = n1131 ^ n1129 ;
  assign n1133 = n155 & n1132 ;
  assign n1134 = n1133 ^ n155 ;
  assign n1135 = n1134 ^ n155 ;
  assign n1102 = n447 ^ x51 ;
  assign n1103 = x129 & n1102 ;
  assign n1100 = x129 & n445 ;
  assign n1101 = n1100 ^ n445 ;
  assign n1104 = n1103 ^ n1101 ;
  assign n1109 = x129 & n451 ;
  assign n1110 = n1109 ^ x129 ;
  assign n1105 = n466 ^ x53 ;
  assign n1106 = x129 & n1105 ;
  assign n1107 = n1106 ^ x129 ;
  assign n1108 = n1107 ^ n1105 ;
  assign n1111 = n1110 ^ n1108 ;
  assign n1112 = n1104 & n1111 ;
  assign n1113 = n1112 ^ n1104 ;
  assign n1114 = n1113 ^ n1111 ;
  assign n1115 = n139 & n1114 ;
  assign n1116 = n1115 ^ n139 ;
  assign n1117 = n1116 ^ n139 ;
  assign n1136 = n1135 ^ n1117 ;
  assign n1139 = n419 ^ x63 ;
  assign n1140 = x129 & n1139 ;
  assign n1137 = x129 & n417 ;
  assign n1138 = n1137 ^ n417 ;
  assign n1141 = n1140 ^ n1138 ;
  assign n1146 = x129 & n423 ;
  assign n1147 = n1146 ^ x129 ;
  assign n1142 = n288 ^ x65 ;
  assign n1143 = x129 & n1142 ;
  assign n1144 = n1143 ^ x129 ;
  assign n1145 = n1144 ^ n1142 ;
  assign n1148 = n1147 ^ n1145 ;
  assign n1149 = n1141 & n1148 ;
  assign n1150 = n1149 ^ n1141 ;
  assign n1151 = n1150 ^ n1148 ;
  assign n1152 = n171 & n1151 ;
  assign n1153 = n1152 ^ n1151 ;
  assign n1154 = n1136 & n1153 ;
  assign n1155 = n1154 ^ n1136 ;
  assign n1156 = n1155 ^ n1153 ;
  assign n1174 = n1173 ^ n1156 ;
  assign n1175 = x134 & ~n138 ;
  assign n1176 = n1174 & n1175 ;
  assign n1177 = n1176 ^ x134 ;
  assign n1178 = n1099 & n1177 ;
  assign n1179 = n1178 ^ n1177 ;
  assign n1258 = n1257 ^ n1179 ;
  assign n1336 = n1335 ^ n1258 ;
  assign n942 = n849 ^ x134 ;
  assign n872 = n325 ^ x75 ;
  assign n873 = x129 & n872 ;
  assign n870 = x129 & n323 ;
  assign n871 = n870 ^ n323 ;
  assign n874 = n873 ^ n871 ;
  assign n879 = x129 & n329 ;
  assign n880 = n879 ^ x129 ;
  assign n875 = n317 ^ x77 ;
  assign n876 = x129 & n875 ;
  assign n877 = n876 ^ x129 ;
  assign n878 = n877 ^ n875 ;
  assign n881 = n880 ^ n878 ;
  assign n882 = n874 & n881 ;
  assign n883 = n882 ^ n874 ;
  assign n884 = n883 ^ n881 ;
  assign n885 = n170 & n884 ;
  assign n886 = n885 ^ n170 ;
  assign n887 = n886 ^ n170 ;
  assign n853 = n311 ^ x79 ;
  assign n854 = x129 & n853 ;
  assign n851 = x129 & n309 ;
  assign n852 = n851 ^ n309 ;
  assign n855 = n854 ^ n852 ;
  assign n860 = x129 & n315 ;
  assign n861 = n860 ^ x129 ;
  assign n856 = n380 ^ x81 ;
  assign n857 = x129 & n856 ;
  assign n858 = n857 ^ x129 ;
  assign n859 = n858 ^ n856 ;
  assign n862 = n861 ^ n859 ;
  assign n863 = n855 & n862 ;
  assign n864 = n863 ^ n855 ;
  assign n865 = n864 ^ n862 ;
  assign n866 = n171 & n865 ;
  assign n867 = n866 ^ n171 ;
  assign n868 = n867 ^ n865 ;
  assign n869 = n868 ^ n171 ;
  assign n888 = n887 ^ n869 ;
  assign n909 = n295 ^ x71 ;
  assign n910 = x129 & n909 ;
  assign n907 = x129 & n293 ;
  assign n908 = n907 ^ n293 ;
  assign n911 = n910 ^ n908 ;
  assign n916 = x129 & n299 ;
  assign n917 = n916 ^ x129 ;
  assign n912 = n331 ^ x73 ;
  assign n913 = x129 & n912 ;
  assign n914 = n913 ^ x129 ;
  assign n915 = n914 ^ n912 ;
  assign n918 = n917 ^ n915 ;
  assign n919 = n911 & n918 ;
  assign n920 = n919 ^ n911 ;
  assign n921 = n920 ^ n918 ;
  assign n922 = n155 & n921 ;
  assign n923 = n922 ^ n155 ;
  assign n924 = n923 ^ n155 ;
  assign n891 = n282 ^ x67 ;
  assign n892 = x129 & n891 ;
  assign n889 = x129 & n280 ;
  assign n890 = n889 ^ n280 ;
  assign n893 = n892 ^ n890 ;
  assign n898 = x129 & n286 ;
  assign n899 = n898 ^ x129 ;
  assign n894 = n301 ^ x69 ;
  assign n895 = x129 & n894 ;
  assign n896 = n895 ^ x129 ;
  assign n897 = n896 ^ n894 ;
  assign n900 = n899 ^ n897 ;
  assign n901 = n893 & n900 ;
  assign n902 = n901 ^ n893 ;
  assign n903 = n902 ^ n900 ;
  assign n904 = n139 & n903 ;
  assign n905 = n904 ^ n139 ;
  assign n906 = n905 ^ n139 ;
  assign n925 = n924 ^ n906 ;
  assign n926 = n888 & n925 ;
  assign n927 = n926 ^ n925 ;
  assign n928 = n927 ^ n925 ;
  assign n929 = n928 ^ n888 ;
  assign n930 = n929 ^ n925 ;
  assign n943 = n930 ^ x134 ;
  assign n944 = n930 & n943 ;
  assign n945 = n944 ^ n930 ;
  assign n946 = n945 ^ n943 ;
  assign n947 = n946 ^ n930 ;
  assign n948 = n947 ^ n943 ;
  assign n949 = n948 ^ x134 ;
  assign n950 = ~n942 & ~n949 ;
  assign n951 = n950 ^ n942 ;
  assign n952 = n951 ^ n949 ;
  assign n953 = n952 ^ n948 ;
  assign n954 = n953 ^ n849 ;
  assign n1337 = n1336 ^ n954 ;
  assign n850 = ~x134 & ~n136 ;
  assign n931 = n930 ^ n850 ;
  assign n932 = n850 & n931 ;
  assign n933 = n932 ^ n850 ;
  assign n934 = n933 ^ n850 ;
  assign n935 = n934 ^ n931 ;
  assign n936 = n935 ^ n930 ;
  assign n937 = n936 ^ n849 ;
  assign n938 = ~n849 & ~n937 ;
  assign n939 = n938 ^ n937 ;
  assign n940 = n939 ^ n935 ;
  assign n941 = n940 ^ n930 ;
  assign n1338 = n1337 ^ n941 ;
  assign n1441 = n441 ^ n440 ;
  assign n1442 = n1441 ^ n462 ;
  assign n1443 = n155 & n1442 ;
  assign n1444 = n1443 ^ n155 ;
  assign n1445 = n1444 ^ n155 ;
  assign n1436 = n468 ^ n467 ;
  assign n1437 = n1436 ^ n449 ;
  assign n1438 = n139 & n1437 ;
  assign n1439 = n1438 ^ n139 ;
  assign n1440 = n1439 ^ n139 ;
  assign n1446 = n1445 ^ n1440 ;
  assign n1488 = n138 & n1446 ;
  assign n1489 = n1488 ^ n1446 ;
  assign n1490 = n1489 ^ n138 ;
  assign n1491 = n427 ^ n426 ;
  assign n1492 = n1491 ^ n435 ;
  assign n1493 = n170 & ~n1492 ;
  assign n1494 = n1493 ^ n170 ;
  assign n1495 = n1490 & n1494 ;
  assign n1496 = n1495 ^ n1494 ;
  assign n1497 = n1496 ^ n1490 ;
  assign n1467 = n171 & n617 ;
  assign n1468 = n1467 ^ n171 ;
  assign n1469 = n1468 ^ n617 ;
  assign n1463 = n588 ^ n587 ;
  assign n1464 = n171 & n1463 ;
  assign n1465 = n1464 ^ n171 ;
  assign n1466 = n1465 ^ n1463 ;
  assign n1470 = n1469 ^ n1466 ;
  assign n1460 = n623 ^ n622 ;
  assign n1461 = n1460 ^ n631 ;
  assign n1462 = n170 & n1461 ;
  assign n1471 = n1470 ^ n1462 ;
  assign n1478 = n139 & n647 ;
  assign n1479 = n1478 ^ n139 ;
  assign n1475 = n666 ^ n665 ;
  assign n1476 = n139 & n1475 ;
  assign n1477 = n1476 ^ n139 ;
  assign n1480 = n1479 ^ n1477 ;
  assign n1472 = n637 ^ n636 ;
  assign n1473 = n1472 ^ n660 ;
  assign n1474 = n155 & n1473 ;
  assign n1481 = n1480 ^ n1474 ;
  assign n1482 = n1471 & n1481 ;
  assign n1483 = n1482 ^ n1471 ;
  assign n1484 = n1483 ^ n1481 ;
  assign n1485 = n136 & n1484 ;
  assign n1486 = n1485 ^ n136 ;
  assign n1487 = n1486 ^ n136 ;
  assign n1498 = n1497 ^ n1487 ;
  assign n1447 = n290 ^ n289 ;
  assign n1448 = n1447 ^ n421 ;
  assign n1449 = n138 & n171 ;
  assign n1450 = n1449 ^ n171 ;
  assign n1451 = n1450 ^ n138 ;
  assign n1452 = n1451 ^ n1448 ;
  assign n1453 = ~n1448 & ~n1452 ;
  assign n1454 = n1453 ^ n1451 ;
  assign n1455 = n1454 ^ n1446 ;
  assign n1456 = n1446 & n1455 ;
  assign n1457 = n1456 ^ n1453 ;
  assign n1458 = n1457 ^ n1451 ;
  assign n1459 = n1458 ^ n138 ;
  assign n1499 = n1498 ^ n1459 ;
  assign n1552 = n171 & n402 ;
  assign n1553 = n1552 ^ n402 ;
  assign n1509 = n574 ^ n573 ;
  assign n1510 = n1509 ^ n595 ;
  assign n1511 = n155 & n1510 ;
  assign n1512 = n1511 ^ n155 ;
  assign n1513 = n1512 ^ n155 ;
  assign n1504 = n601 ^ n600 ;
  assign n1505 = n1504 ^ n582 ;
  assign n1506 = n139 & n1505 ;
  assign n1507 = n1506 ^ n139 ;
  assign n1508 = n1507 ^ n139 ;
  assign n1514 = n1513 ^ n1508 ;
  assign n1554 = n1553 ^ n1514 ;
  assign n1555 = n519 ^ n518 ;
  assign n1556 = n1555 ^ n554 ;
  assign n1557 = n1556 ^ n1553 ;
  assign n1558 = ~n1556 & n1557 ;
  assign n1559 = n1558 ^ n1553 ;
  assign n1560 = ~n1554 & ~n1559 ;
  assign n1561 = n1560 ^ n1558 ;
  assign n1562 = n1561 ^ n1514 ;
  assign n1532 = n531 ^ x128 ;
  assign n1531 = n523 ^ x128 ;
  assign n1533 = n1532 ^ n1531 ;
  assign n1534 = x129 & n1533 ;
  assign n1535 = n1534 ^ x129 ;
  assign n1529 = n488 ^ x129 ;
  assign n1530 = n1529 ^ n487 ;
  assign n1536 = n1535 ^ n1530 ;
  assign n1537 = n155 & n1536 ;
  assign n1526 = n513 ^ x129 ;
  assign n1521 = n535 ^ x128 ;
  assign n1520 = n527 ^ x128 ;
  assign n1522 = n1521 ^ n1520 ;
  assign n1523 = x129 & n1522 ;
  assign n1524 = n1523 ^ x129 ;
  assign n1525 = n1524 ^ n1522 ;
  assign n1527 = n1526 ^ n1525 ;
  assign n1528 = n139 & n1527 ;
  assign n1538 = n1537 ^ n1528 ;
  assign n1539 = n137 & n1538 ;
  assign n1540 = n1539 ^ n137 ;
  assign n1546 = n502 ^ n501 ;
  assign n1547 = n1546 ^ n482 ;
  assign n1548 = n170 & n1547 ;
  assign n1549 = n1540 & n1548 ;
  assign n1550 = n1549 ^ n137 ;
  assign n1541 = n455 ^ n454 ;
  assign n1542 = n1541 ^ n496 ;
  assign n1543 = ~n171 & n1542 ;
  assign n1544 = n1540 & n1543 ;
  assign n1545 = n1544 ^ n1540 ;
  assign n1551 = n1550 ^ n1545 ;
  assign n1563 = n1562 ^ n1551 ;
  assign n1500 = n560 ^ n559 ;
  assign n1501 = n1500 ^ n568 ;
  assign n1502 = n170 & ~n1501 ;
  assign n1503 = n1502 ^ n170 ;
  assign n1515 = n402 & n1514 ;
  assign n1516 = n1515 ^ n402 ;
  assign n1517 = n1503 & n1516 ;
  assign n1518 = n1517 ^ n1516 ;
  assign n1519 = n1518 ^ n402 ;
  assign n1564 = n1563 ^ n1519 ;
  assign n1565 = n1499 & n1564 ;
  assign n1566 = n1565 ^ n1499 ;
  assign n1567 = n1566 ^ n1564 ;
  assign n1568 = n1567 ^ n1499 ;
  assign n1569 = n1568 ^ n1564 ;
  assign n1570 = x134 & ~n1569 ;
  assign n1571 = n1570 ^ x134 ;
  assign n1370 = n395 ^ n394 ;
  assign n1371 = n1370 ^ n376 ;
  assign n1372 = n139 & ~n1371 ;
  assign n1373 = n1372 ^ n139 ;
  assign n1366 = n355 ^ n354 ;
  assign n1367 = n1366 ^ n362 ;
  assign n1368 = n170 & n1367 ;
  assign n1363 = n249 ^ n248 ;
  assign n1364 = n1363 ^ n349 ;
  assign n1365 = ~n171 & n1364 ;
  assign n1369 = n1368 ^ n1365 ;
  assign n1374 = n1373 ^ n1369 ;
  assign n1359 = n368 ^ n367 ;
  assign n1360 = n1359 ^ n389 ;
  assign n1361 = n155 & ~n1360 ;
  assign n1362 = n1361 ^ n155 ;
  assign n1375 = n1374 ^ n1362 ;
  assign n1376 = n402 & n1375 ;
  assign n1342 = n333 ^ n332 ;
  assign n1343 = n1342 ^ n297 ;
  assign n1344 = n155 & n1343 ;
  assign n1339 = n303 ^ n302 ;
  assign n1340 = n1339 ^ n284 ;
  assign n1341 = n139 & n1340 ;
  assign n1345 = n1344 ^ n1341 ;
  assign n1346 = n136 & n1345 ;
  assign n1347 = n1346 ^ n136 ;
  assign n1353 = n319 ^ n318 ;
  assign n1354 = n1353 ^ n327 ;
  assign n1355 = n170 & n1354 ;
  assign n1356 = n1347 & n1355 ;
  assign n1357 = n1356 ^ n136 ;
  assign n1348 = n382 ^ n381 ;
  assign n1349 = n1348 ^ n313 ;
  assign n1350 = ~n171 & n1349 ;
  assign n1351 = n1347 & n1350 ;
  assign n1352 = n1351 ^ n1347 ;
  assign n1358 = n1357 ^ n1352 ;
  assign n1377 = n1376 ^ n1358 ;
  assign n1410 = n217 ^ n216 ;
  assign n1411 = n1410 ^ n227 ;
  assign n1412 = n170 & n1411 ;
  assign n1406 = n150 ^ n149 ;
  assign n1407 = n1406 ^ n211 ;
  assign n1408 = n171 & n1407 ;
  assign n1409 = n1408 ^ n1407 ;
  assign n1413 = n1412 ^ n1409 ;
  assign n1417 = n233 ^ n232 ;
  assign n1418 = n1417 ^ n258 ;
  assign n1419 = n155 & n1418 ;
  assign n1414 = n264 ^ n263 ;
  assign n1415 = n1414 ^ n243 ;
  assign n1416 = n139 & n1415 ;
  assign n1420 = n1419 ^ n1416 ;
  assign n1421 = n1413 & n1420 ;
  assign n1422 = n1421 ^ n1413 ;
  assign n1423 = n1422 ^ n1420 ;
  assign n1424 = n137 & n1423 ;
  assign n1425 = n1424 ^ n137 ;
  assign n1426 = n1425 ^ n137 ;
  assign n1384 = n155 & n160 ;
  assign n1385 = n1384 ^ n155 ;
  assign n1381 = n196 ^ n195 ;
  assign n1382 = n155 & n1381 ;
  assign n1383 = n1382 ^ n155 ;
  assign n1386 = n1385 ^ n1383 ;
  assign n1378 = n166 ^ n165 ;
  assign n1379 = n1378 ^ n144 ;
  assign n1380 = n139 & n1379 ;
  assign n1387 = n1386 ^ n1380 ;
  assign n1388 = n138 & n1387 ;
  assign n1389 = n1388 ^ n1387 ;
  assign n1390 = n1389 ^ n138 ;
  assign n1399 = n182 ^ n181 ;
  assign n1400 = n1399 ^ n190 ;
  assign n1401 = n170 & n1400 ;
  assign n1402 = n1390 & n1401 ;
  assign n1403 = n1402 ^ n1401 ;
  assign n1404 = n1403 ^ n138 ;
  assign n1391 = n653 ^ n652 ;
  assign n1392 = n1391 ^ n176 ;
  assign n1393 = ~n171 & ~n1392 ;
  assign n1394 = n1393 ^ n171 ;
  assign n1395 = n1390 & n1394 ;
  assign n1396 = n1395 ^ n1394 ;
  assign n1397 = n1396 ^ n1390 ;
  assign n1398 = n1397 ^ n1390 ;
  assign n1405 = n1404 ^ n1398 ;
  assign n1427 = n1426 ^ n1405 ;
  assign n1428 = n1377 & n1427 ;
  assign n1429 = n1428 ^ n1377 ;
  assign n1430 = n1429 ^ n1377 ;
  assign n1431 = n1430 ^ n1427 ;
  assign n1432 = x134 & n1431 ;
  assign n1433 = n1432 ^ x134 ;
  assign n1434 = n1433 ^ x134 ;
  assign n1435 = n1434 ^ n1431 ;
  assign n1572 = n1571 ^ n1435 ;
  assign n1634 = n854 ^ n853 ;
  assign n1635 = n1634 ^ n870 ;
  assign n1636 = n861 ^ n315 ;
  assign n1637 = n1636 ^ n877 ;
  assign n1638 = n1635 & n1637 ;
  assign n1639 = n1638 ^ n1635 ;
  assign n1640 = n1639 ^ n1637 ;
  assign n1641 = n170 & n1640 ;
  assign n1625 = n1297 ^ n1296 ;
  assign n1626 = n1625 ^ n851 ;
  assign n1627 = n1304 ^ n378 ;
  assign n1628 = n1627 ^ n858 ;
  assign n1629 = n1626 & n1628 ;
  assign n1630 = n1629 ^ n1626 ;
  assign n1631 = n1630 ^ n1628 ;
  assign n1632 = n171 & n1631 ;
  assign n1633 = n1632 ^ n1631 ;
  assign n1642 = n1641 ^ n1633 ;
  assign n1653 = n873 ^ n872 ;
  assign n1654 = n1653 ^ n907 ;
  assign n1655 = n880 ^ n329 ;
  assign n1656 = n1655 ^ n914 ;
  assign n1657 = n1654 & n1656 ;
  assign n1658 = n1657 ^ n1654 ;
  assign n1659 = n1658 ^ n1656 ;
  assign n1660 = n155 & n1659 ;
  assign n1643 = n910 ^ n909 ;
  assign n1644 = n1643 ^ n889 ;
  assign n1645 = n917 ^ n299 ;
  assign n1646 = n1645 ^ n896 ;
  assign n1647 = n1644 & n1646 ;
  assign n1648 = n1647 ^ n1644 ;
  assign n1649 = n1648 ^ n1646 ;
  assign n1650 = n139 & n1649 ;
  assign n1651 = n1650 ^ n139 ;
  assign n1652 = n1651 ^ n139 ;
  assign n1661 = n1660 ^ n1652 ;
  assign n1662 = n1642 & n1661 ;
  assign n1663 = n1662 ^ n1642 ;
  assign n1664 = n1663 ^ n1661 ;
  assign n1665 = n136 & n1664 ;
  assign n1666 = n1665 ^ n136 ;
  assign n1667 = n1666 ^ n136 ;
  assign n1584 = n687 ^ n686 ;
  assign n1585 = n1584 ^ n703 ;
  assign n1586 = n694 ^ n178 ;
  assign n1587 = n1586 ^ n710 ;
  assign n1588 = n1585 & n1587 ;
  assign n1589 = n1588 ^ n1585 ;
  assign n1590 = n1589 ^ n1587 ;
  assign n1591 = n170 & n1590 ;
  assign n1592 = n1591 ^ n170 ;
  assign n1593 = n1592 ^ n170 ;
  assign n1573 = n1218 ^ n1217 ;
  assign n1574 = n1573 ^ n684 ;
  assign n1575 = n1225 ^ n649 ;
  assign n1576 = n1575 ^ n691 ;
  assign n1577 = n1574 & n1576 ;
  assign n1578 = n1577 ^ n1574 ;
  assign n1579 = n1578 ^ n1576 ;
  assign n1580 = n171 & n1579 ;
  assign n1581 = n1580 ^ n171 ;
  assign n1582 = n1581 ^ n1579 ;
  assign n1583 = n1582 ^ n171 ;
  assign n1594 = n1593 ^ n1583 ;
  assign n1605 = n706 ^ n705 ;
  assign n1606 = n1605 ^ n740 ;
  assign n1607 = n713 ^ n192 ;
  assign n1608 = n1607 ^ n747 ;
  assign n1609 = n1606 & n1608 ;
  assign n1610 = n1609 ^ n1606 ;
  assign n1611 = n1610 ^ n1608 ;
  assign n1612 = n155 & n1611 ;
  assign n1613 = n1612 ^ n155 ;
  assign n1614 = n1613 ^ n155 ;
  assign n1595 = n743 ^ n742 ;
  assign n1596 = n1595 ^ n722 ;
  assign n1597 = n750 ^ n162 ;
  assign n1598 = n1597 ^ n729 ;
  assign n1599 = n1596 & n1598 ;
  assign n1600 = n1599 ^ n1596 ;
  assign n1601 = n1600 ^ n1598 ;
  assign n1602 = n139 & n1601 ;
  assign n1603 = n1602 ^ n139 ;
  assign n1604 = n1603 ^ n139 ;
  assign n1615 = n1614 ^ n1604 ;
  assign n1616 = n1594 & n1615 ;
  assign n1617 = n1616 ^ n1615 ;
  assign n1618 = n1617 ^ n1615 ;
  assign n1619 = n1618 ^ n1594 ;
  assign n1620 = n1619 ^ n1615 ;
  assign n1621 = n138 & n1620 ;
  assign n1622 = n1621 ^ n138 ;
  assign n1623 = n1622 ^ n1620 ;
  assign n1624 = n1623 ^ n138 ;
  assign n1668 = n1667 ^ n1624 ;
  assign n1967 = n1263 ^ n1262 ;
  assign n1968 = n1967 ^ n1277 ;
  assign n1969 = n1270 ^ n351 ;
  assign n1970 = n1969 ^ n1284 ;
  assign n1971 = n1968 & n1970 ;
  assign n1972 = n1971 ^ n1968 ;
  assign n1973 = n1972 ^ n1970 ;
  assign n1974 = n170 & n1973 ;
  assign n1975 = n1974 ^ n170 ;
  assign n1976 = n1975 ^ n170 ;
  assign n1956 = n809 ^ n808 ;
  assign n1957 = n1956 ^ n1260 ;
  assign n1958 = n816 ^ n245 ;
  assign n1959 = n1958 ^ n1267 ;
  assign n1960 = n1957 & n1959 ;
  assign n1961 = n1960 ^ n1957 ;
  assign n1962 = n1961 ^ n1959 ;
  assign n1963 = n171 & n1962 ;
  assign n1964 = n1963 ^ n171 ;
  assign n1965 = n1964 ^ n1962 ;
  assign n1966 = n1965 ^ n171 ;
  assign n1977 = n1976 ^ n1966 ;
  assign n1986 = n1280 ^ n1279 ;
  assign n1987 = n1986 ^ n1312 ;
  assign n1988 = n1287 ^ n364 ;
  assign n1989 = n1988 ^ n1319 ;
  assign n1990 = n1987 & n1989 ;
  assign n1991 = n1990 ^ n1987 ;
  assign n1992 = n1991 ^ n1989 ;
  assign n1993 = n155 & n1992 ;
  assign n1978 = n1315 ^ n1314 ;
  assign n1979 = n1978 ^ n1294 ;
  assign n1980 = n1322 ^ n391 ;
  assign n1981 = n1980 ^ n1301 ;
  assign n1982 = n1979 & n1981 ;
  assign n1983 = n1982 ^ n1979 ;
  assign n1984 = n1983 ^ n1981 ;
  assign n1985 = n139 & n1984 ;
  assign n1994 = n1993 ^ n1985 ;
  assign n1995 = n1977 & n1994 ;
  assign n1996 = n1995 ^ n1994 ;
  assign n1997 = n1996 ^ n1994 ;
  assign n1998 = n1997 ^ n1977 ;
  assign n1999 = n1998 ^ n1994 ;
  assign n2000 = n1259 & n1999 ;
  assign n2001 = n2000 ^ n1259 ;
  assign n2002 = n2001 ^ n1259 ;
  assign n2003 = ~n1668 & n2002 ;
  assign n2004 = n2003 ^ n2002 ;
  assign n2005 = n2004 ^ n2002 ;
  assign n1917 = n1082 ^ n1081 ;
  assign n1918 = n1917 ^ n988 ;
  assign n1919 = n1089 ^ n556 ;
  assign n1920 = n1919 ^ n995 ;
  assign n1921 = n1918 & n1920 ;
  assign n1922 = n1921 ^ n1918 ;
  assign n1923 = n1922 ^ n1920 ;
  assign n1924 = n170 & n1923 ;
  assign n1908 = n1017 ^ n1016 ;
  assign n1909 = n1908 ^ n1079 ;
  assign n1910 = n1014 ^ n515 ;
  assign n1911 = n1910 ^ n1086 ;
  assign n1912 = n1909 & n1911 ;
  assign n1913 = n1912 ^ n1909 ;
  assign n1914 = n1913 ^ n1911 ;
  assign n1915 = n171 & n1914 ;
  assign n1916 = n1915 ^ n1914 ;
  assign n1925 = n1924 ^ n1916 ;
  assign n1936 = n991 ^ n990 ;
  assign n1937 = n1936 ^ n971 ;
  assign n1938 = n998 ^ n570 ;
  assign n1939 = n1938 ^ n978 ;
  assign n1940 = n1937 & n1939 ;
  assign n1941 = n1940 ^ n1937 ;
  assign n1942 = n1941 ^ n1939 ;
  assign n1943 = n155 & n1942 ;
  assign n1944 = n1943 ^ n155 ;
  assign n1945 = n1944 ^ n155 ;
  assign n1926 = n974 ^ n973 ;
  assign n1927 = n1926 ^ n955 ;
  assign n1928 = n981 ^ n597 ;
  assign n1929 = n1928 ^ n962 ;
  assign n1930 = n1927 & n1929 ;
  assign n1931 = n1930 ^ n1927 ;
  assign n1932 = n1931 ^ n1929 ;
  assign n1933 = n139 & n1932 ;
  assign n1934 = n1933 ^ n139 ;
  assign n1935 = n1934 ^ n139 ;
  assign n1946 = n1945 ^ n1935 ;
  assign n1947 = ~n1925 & n1946 ;
  assign n1948 = n1947 ^ n1925 ;
  assign n1796 = n1044 & n1102 ;
  assign n1797 = n1796 ^ n1102 ;
  assign n1787 = n498 ^ x128 ;
  assign n1786 = n1051 ^ x128 ;
  assign n1788 = n1787 ^ n1786 ;
  assign n1789 = x129 & n1788 ;
  assign n1790 = n1789 ^ x129 ;
  assign n1791 = n1790 ^ n1788 ;
  assign n1792 = n1791 ^ n1062 ;
  assign n1793 = n170 & n1792 ;
  assign n1794 = n1793 ^ n170 ;
  assign n1795 = n1794 ^ n170 ;
  assign n1798 = n1797 ^ n1795 ;
  assign n1777 = x129 & n492 ;
  assign n1778 = n1777 ^ x129 ;
  assign n1779 = n171 & n1045 ;
  assign n1780 = n1779 ^ n171 ;
  assign n1781 = n1780 ^ n1045 ;
  assign n1782 = n1778 & n1781 ;
  assign n1783 = n1782 ^ n1778 ;
  assign n1774 = n451 & n1044 ;
  assign n1775 = n1774 ^ n451 ;
  assign n1776 = n1775 ^ n1044 ;
  assign n1784 = n1783 ^ n1776 ;
  assign n1785 = n1784 ^ n171 ;
  assign n1799 = n1798 ^ n1785 ;
  assign n1839 = x129 & n1030 ;
  assign n1840 = n1839 ^ n1030 ;
  assign n1838 = x129 & n509 ;
  assign n1841 = n1840 ^ n1838 ;
  assign n1842 = x129 & n526 ;
  assign n1843 = n1842 ^ x129 ;
  assign n1844 = n1843 ^ n526 ;
  assign n1845 = n1844 ^ n1011 ;
  assign n1846 = n1841 & n1845 ;
  assign n1847 = n1846 ^ n1841 ;
  assign n1848 = n1847 ^ n1845 ;
  assign n1849 = n137 & n139 ;
  assign n1850 = n1848 & n1849 ;
  assign n1851 = n1850 ^ n137 ;
  assign n1852 = n1799 & n1851 ;
  assign n1853 = n1852 ^ n1851 ;
  assign n1854 = n1853 ^ n1851 ;
  assign n1855 = n1854 ^ n1851 ;
  assign n1751 = n1161 ^ n1160 ;
  assign n1752 = n1751 ^ n1118 ;
  assign n1753 = n1168 ^ n437 ;
  assign n1754 = n1753 ^ n1125 ;
  assign n1755 = n1752 & n1754 ;
  assign n1756 = n1755 ^ n1752 ;
  assign n1757 = n1756 ^ n1754 ;
  assign n1758 = n155 & n1757 ;
  assign n1759 = n1758 ^ n155 ;
  assign n1760 = n1759 ^ n155 ;
  assign n1741 = n1121 ^ n1120 ;
  assign n1742 = n1741 ^ n1100 ;
  assign n1743 = n1128 ^ n464 ;
  assign n1744 = n1743 ^ n1107 ;
  assign n1745 = n1742 & n1744 ;
  assign n1746 = n1745 ^ n1742 ;
  assign n1747 = n1746 ^ n1744 ;
  assign n1748 = n139 & n1747 ;
  assign n1749 = n1748 ^ n139 ;
  assign n1750 = n1749 ^ n139 ;
  assign n1761 = n1760 ^ n1750 ;
  assign n1820 = n1140 ^ n1139 ;
  assign n1821 = n1820 ^ n1158 ;
  assign n1822 = n1147 ^ n423 ;
  assign n1823 = n1822 ^ n1165 ;
  assign n1824 = n1821 & n1823 ;
  assign n1825 = n1824 ^ n1821 ;
  assign n1826 = n1825 ^ n1823 ;
  assign n1831 = n138 & n1826 ;
  assign n1832 = n1831 ^ n1826 ;
  assign n1833 = n1832 ^ n138 ;
  assign n1834 = n1761 & n1833 ;
  assign n1835 = n1834 ^ n1761 ;
  assign n1836 = n1835 ^ n1833 ;
  assign n1827 = ~n138 & ~n170 ;
  assign n1828 = n1826 & n1827 ;
  assign n1829 = n1761 & n1828 ;
  assign n1830 = n1829 ^ n1828 ;
  assign n1837 = n1836 ^ n1830 ;
  assign n1856 = n1855 ^ n1837 ;
  assign n1802 = x129 & n530 ;
  assign n1800 = x129 & n1064 ;
  assign n1801 = n1800 ^ n1064 ;
  assign n1803 = n1802 ^ n1801 ;
  assign n1807 = x129 & n1023 ;
  assign n1808 = n1807 ^ x129 ;
  assign n1804 = x129 & n484 ;
  assign n1805 = n1804 ^ x129 ;
  assign n1806 = n1805 ^ n484 ;
  assign n1809 = n1808 ^ n1806 ;
  assign n1810 = n1803 & n1809 ;
  assign n1811 = n1810 ^ n1803 ;
  assign n1812 = n1811 ^ n1809 ;
  assign n1813 = n137 & n155 ;
  assign n1814 = n1812 & n1813 ;
  assign n1815 = n1799 & n1814 ;
  assign n1816 = n1815 ^ n1814 ;
  assign n1817 = n1816 ^ n1814 ;
  assign n1818 = n1817 ^ n1814 ;
  assign n1819 = n1818 ^ n137 ;
  assign n1857 = n1856 ^ n1819 ;
  assign n1762 = n892 ^ n891 ;
  assign n1763 = n1762 ^ n1137 ;
  assign n1764 = n899 ^ n286 ;
  assign n1765 = n1764 ^ n1144 ;
  assign n1766 = n1763 & n1765 ;
  assign n1767 = n1766 ^ n1763 ;
  assign n1768 = n1767 ^ n1765 ;
  assign n1769 = n1451 & n1768 ;
  assign n1770 = n1769 ^ n1768 ;
  assign n1771 = n1761 & n1770 ;
  assign n1772 = n1771 ^ n1770 ;
  assign n1773 = n1772 ^ n138 ;
  assign n1858 = n1857 ^ n1773 ;
  assign n1949 = x134 & n402 ;
  assign n1950 = n1858 & n1949 ;
  assign n1951 = n1950 ^ n1949 ;
  assign n1952 = n1948 & n1951 ;
  assign n1953 = n1952 ^ n1951 ;
  assign n1954 = n1953 ^ n1951 ;
  assign n1868 = n1184 ^ n1183 ;
  assign n1869 = n1868 ^ n1198 ;
  assign n1870 = n1191 ^ n619 ;
  assign n1871 = n1870 ^ n1205 ;
  assign n1872 = n1869 & n1871 ;
  assign n1873 = n1872 ^ n1869 ;
  assign n1874 = n1873 ^ n1871 ;
  assign n1875 = n170 & n1874 ;
  assign n1859 = n958 ^ n957 ;
  assign n1860 = n1859 ^ n1181 ;
  assign n1861 = n965 ^ n584 ;
  assign n1862 = n1861 ^ n1188 ;
  assign n1863 = n1860 & n1862 ;
  assign n1864 = n1863 ^ n1860 ;
  assign n1865 = n1864 ^ n1862 ;
  assign n1866 = n171 & n1865 ;
  assign n1867 = n1866 ^ n1865 ;
  assign n1876 = n1875 ^ n1867 ;
  assign n1887 = n1201 ^ n1200 ;
  assign n1888 = n1887 ^ n1233 ;
  assign n1889 = n1208 ^ n633 ;
  assign n1890 = n1889 ^ n1240 ;
  assign n1891 = n1888 & n1890 ;
  assign n1892 = n1891 ^ n1888 ;
  assign n1893 = n1892 ^ n1890 ;
  assign n1894 = n155 & n1893 ;
  assign n1877 = n1236 ^ n1235 ;
  assign n1878 = n1877 ^ n1215 ;
  assign n1879 = n1243 ^ n662 ;
  assign n1880 = n1879 ^ n1222 ;
  assign n1881 = n1878 & n1880 ;
  assign n1882 = n1881 ^ n1878 ;
  assign n1883 = n1882 ^ n1880 ;
  assign n1884 = n139 & n1883 ;
  assign n1885 = n1884 ^ n139 ;
  assign n1886 = n1885 ^ n139 ;
  assign n1895 = n1894 ^ n1886 ;
  assign n1896 = n1876 & n1895 ;
  assign n1897 = n1896 ^ n1876 ;
  assign n1898 = n1897 ^ n1895 ;
  assign n1903 = x134 & n1898 ;
  assign n1904 = n1903 ^ x134 ;
  assign n1905 = n1858 & n1904 ;
  assign n1906 = n1905 ^ n1904 ;
  assign n1899 = x134 & ~n136 ;
  assign n1900 = n1898 & n1899 ;
  assign n1901 = n1858 & n1900 ;
  assign n1902 = n1901 ^ n1900 ;
  assign n1907 = n1906 ^ n1902 ;
  assign n1955 = n1954 ^ n1907 ;
  assign n2006 = n2005 ^ n1955 ;
  assign n1727 = n1668 ^ x134 ;
  assign n1681 = n771 ^ n770 ;
  assign n1682 = n1681 ^ n787 ;
  assign n1683 = n778 ^ n213 ;
  assign n1684 = n1683 ^ n794 ;
  assign n1685 = n1682 & n1684 ;
  assign n1686 = n1685 ^ n1682 ;
  assign n1687 = n1686 ^ n1684 ;
  assign n1688 = n170 & n1687 ;
  assign n1689 = n1688 ^ n170 ;
  assign n1690 = n1689 ^ n170 ;
  assign n1670 = n725 ^ n724 ;
  assign n1671 = n1670 ^ n768 ;
  assign n1672 = n732 ^ n146 ;
  assign n1673 = n1672 ^ n775 ;
  assign n1674 = n1671 & n1673 ;
  assign n1675 = n1674 ^ n1671 ;
  assign n1676 = n1675 ^ n1673 ;
  assign n1677 = n171 & n1676 ;
  assign n1678 = n1677 ^ n171 ;
  assign n1679 = n1678 ^ n1676 ;
  assign n1680 = n1679 ^ n171 ;
  assign n1691 = n1690 ^ n1680 ;
  assign n1702 = n790 ^ n789 ;
  assign n1703 = n1702 ^ n822 ;
  assign n1704 = n797 ^ n229 ;
  assign n1705 = n1704 ^ n829 ;
  assign n1706 = n1703 & n1705 ;
  assign n1707 = n1706 ^ n1703 ;
  assign n1708 = n1707 ^ n1705 ;
  assign n1709 = n155 & n1708 ;
  assign n1710 = n1709 ^ n155 ;
  assign n1711 = n1710 ^ n155 ;
  assign n1692 = n825 ^ n824 ;
  assign n1693 = n1692 ^ n806 ;
  assign n1694 = n832 ^ n260 ;
  assign n1695 = n1694 ^ n813 ;
  assign n1696 = n1693 & n1695 ;
  assign n1697 = n1696 ^ n1693 ;
  assign n1698 = n1697 ^ n1695 ;
  assign n1699 = n139 & n1698 ;
  assign n1700 = n1699 ^ n139 ;
  assign n1701 = n1700 ^ n139 ;
  assign n1712 = n1711 ^ n1701 ;
  assign n1713 = n1691 & n1712 ;
  assign n1714 = n1713 ^ n1712 ;
  assign n1715 = n1714 ^ n1691 ;
  assign n1728 = n1715 ^ x134 ;
  assign n1729 = n1715 & n1728 ;
  assign n1730 = n1729 ^ n1715 ;
  assign n1731 = n1730 ^ n1728 ;
  assign n1732 = n1731 ^ n1715 ;
  assign n1733 = n1732 ^ n1728 ;
  assign n1734 = n1733 ^ x134 ;
  assign n1735 = ~n1727 & ~n1734 ;
  assign n1736 = n1735 ^ n1727 ;
  assign n1737 = n1736 ^ n1734 ;
  assign n1738 = n1737 ^ n1733 ;
  assign n1739 = n1738 ^ n1668 ;
  assign n1669 = ~x134 & ~n137 ;
  assign n1716 = n1715 ^ n1669 ;
  assign n1717 = n1669 & n1716 ;
  assign n1718 = n1717 ^ n1669 ;
  assign n1719 = n1718 ^ n1669 ;
  assign n1720 = n1719 ^ n1716 ;
  assign n1721 = n1720 ^ n1715 ;
  assign n1722 = n1721 ^ n1668 ;
  assign n1723 = ~n1668 & ~n1722 ;
  assign n1724 = n1723 ^ n1722 ;
  assign n1725 = n1724 ^ n1720 ;
  assign n1726 = n1725 ^ n1715 ;
  assign n1740 = n1739 ^ n1726 ;
  assign n2007 = n2006 ^ n1740 ;
  assign n2026 = n170 & n218 ;
  assign n2027 = n2026 ^ n170 ;
  assign n2028 = n2027 ^ n170 ;
  assign n2022 = n151 & n171 ;
  assign n2023 = n2022 ^ n151 ;
  assign n2024 = n2023 ^ n171 ;
  assign n2025 = n2024 ^ n171 ;
  assign n2029 = n2028 ^ n2025 ;
  assign n2033 = n155 & n234 ;
  assign n2034 = n2033 ^ n155 ;
  assign n2035 = n2034 ^ n155 ;
  assign n2030 = n139 & n265 ;
  assign n2031 = n2030 ^ n139 ;
  assign n2032 = n2031 ^ n139 ;
  assign n2036 = n2035 ^ n2032 ;
  assign n2037 = n2029 & n2036 ;
  assign n2038 = n2037 ^ n2029 ;
  assign n2039 = n2038 ^ n2036 ;
  assign n2040 = n137 & n2039 ;
  assign n2041 = n2040 ^ n137 ;
  assign n2042 = n2041 ^ n137 ;
  assign n2010 = n170 & n183 ;
  assign n2008 = n171 & n654 ;
  assign n2009 = n2008 ^ n654 ;
  assign n2011 = n2010 ^ n2009 ;
  assign n2013 = n155 & n197 ;
  assign n2012 = n139 & n167 ;
  assign n2014 = n2013 ^ n2012 ;
  assign n2015 = n2011 & n2014 ;
  assign n2016 = n2015 ^ n2011 ;
  assign n2017 = n2016 ^ n2014 ;
  assign n2018 = n138 & n2017 ;
  assign n2019 = n2018 ^ n138 ;
  assign n2020 = n2019 ^ n2017 ;
  assign n2021 = n2020 ^ n138 ;
  assign n2043 = n2042 ^ n2021 ;
  assign n2141 = n2043 ^ n402 ;
  assign n2142 = n407 & ~n2141 ;
  assign n2143 = n2142 ^ n407 ;
  assign n2144 = n2143 ^ n407 ;
  assign n2145 = n2144 ^ n2141 ;
  assign n2146 = n2145 ^ n405 ;
  assign n2140 = n2043 ^ x134 ;
  assign n2147 = n2146 ^ n2140 ;
  assign n2065 = n170 & n356 ;
  assign n2064 = ~n171 & n250 ;
  assign n2066 = n2065 ^ n2064 ;
  assign n2068 = n155 & n369 ;
  assign n2067 = n139 & n396 ;
  assign n2069 = n2068 ^ n2067 ;
  assign n2070 = ~n2066 & ~n2069 ;
  assign n2148 = n2145 ^ n2070 ;
  assign n2149 = n2148 ^ x134 ;
  assign n2150 = n2147 & ~n2149 ;
  assign n2151 = n2150 ^ n2149 ;
  assign n2152 = n2151 ^ n405 ;
  assign n2085 = n171 & n291 ;
  assign n2086 = n2085 ^ n291 ;
  assign n2084 = n170 & n428 ;
  assign n2087 = n2086 ^ n2084 ;
  assign n2089 = n155 & n442 ;
  assign n2088 = n139 & n469 ;
  assign n2090 = n2089 ^ n2088 ;
  assign n2091 = n2087 & n2090 ;
  assign n2092 = n2091 ^ n2087 ;
  assign n2093 = n2092 ^ n2090 ;
  assign n2094 = n138 & n2093 ;
  assign n2095 = n2094 ^ n2093 ;
  assign n2096 = n2095 ^ n138 ;
  assign n2073 = n456 & n505 ;
  assign n2074 = n2073 ^ n137 ;
  assign n2072 = n490 & n503 ;
  assign n2075 = n2074 ^ n2072 ;
  assign n2080 = n155 & n489 ;
  assign n2081 = n2075 & n2080 ;
  assign n2082 = n2081 ^ n2075 ;
  assign n2076 = n139 & n2075 ;
  assign n2077 = n541 & n2076 ;
  assign n2078 = n2077 ^ n2076 ;
  assign n2079 = n2078 ^ n2076 ;
  assign n2083 = n2082 ^ n2079 ;
  assign n2097 = n2096 ^ n2083 ;
  assign n2098 = n2097 ^ x133 ;
  assign n2123 = n155 & n638 ;
  assign n2124 = n2123 ^ n155 ;
  assign n2125 = n2124 ^ n155 ;
  assign n2122 = n139 & n667 ;
  assign n2126 = n2125 ^ n2122 ;
  assign n2129 = n170 & n624 ;
  assign n2127 = n171 & n589 ;
  assign n2128 = n2127 ^ n589 ;
  assign n2130 = n2129 ^ n2128 ;
  assign n2131 = n2126 & n2130 ;
  assign n2132 = n2131 ^ n2130 ;
  assign n2133 = n2132 ^ n2126 ;
  assign n2134 = n136 & n2133 ;
  assign n2135 = n2098 & n2134 ;
  assign n2136 = n2135 ^ n2134 ;
  assign n2137 = n2136 ^ n2098 ;
  assign n2099 = n2098 ^ n402 ;
  assign n2102 = n170 & n561 ;
  assign n2100 = n171 & n520 ;
  assign n2101 = n2100 ^ n520 ;
  assign n2103 = n2102 ^ n2101 ;
  assign n2105 = n155 & n575 ;
  assign n2104 = n139 & n602 ;
  assign n2106 = n2105 ^ n2104 ;
  assign n2107 = n2103 & n2106 ;
  assign n2108 = n2107 ^ n2103 ;
  assign n2109 = n2108 ^ n2106 ;
  assign n2110 = n2109 ^ n402 ;
  assign n2111 = n2109 & n2110 ;
  assign n2112 = n2111 ^ n2109 ;
  assign n2113 = n2112 ^ n2110 ;
  assign n2114 = n2113 ^ n2109 ;
  assign n2115 = n2114 ^ n402 ;
  assign n2116 = n2099 & ~n2115 ;
  assign n2117 = n2116 ^ n2099 ;
  assign n2118 = n2117 ^ n2115 ;
  assign n2119 = n2118 ^ n2099 ;
  assign n2120 = n2119 ^ n2114 ;
  assign n2121 = n2120 ^ n2098 ;
  assign n2138 = n2137 ^ n2121 ;
  assign n2139 = x134 & ~n2138 ;
  assign n2153 = n2152 ^ n2139 ;
  assign n2071 = n2070 ^ n2043 ;
  assign n2154 = n2153 ^ n2071 ;
  assign n2044 = x134 & ~n2043 ;
  assign n2045 = n2044 ^ x134 ;
  assign n2046 = n2045 ^ x134 ;
  assign n2047 = n2046 ^ n2043 ;
  assign n2051 = n155 & n334 ;
  assign n2048 = n139 & n304 ;
  assign n2049 = n2048 ^ n139 ;
  assign n2050 = n2049 ^ n139 ;
  assign n2052 = n2051 ^ n2050 ;
  assign n2055 = n170 & n320 ;
  assign n2053 = n171 & n383 ;
  assign n2054 = n2053 ^ n383 ;
  assign n2056 = n2055 ^ n2054 ;
  assign n2057 = n2052 & n2056 ;
  assign n2058 = n2057 ^ n2056 ;
  assign n2059 = n2058 ^ n2052 ;
  assign n2060 = n136 & ~n2059 ;
  assign n2061 = n2060 ^ n136 ;
  assign n2062 = ~n2047 & n2061 ;
  assign n2063 = n2062 ^ n2047 ;
  assign n2155 = n2154 ^ n2063 ;
  assign n2347 = ~x132 & x133 ;
  assign n2348 = ~x134 & n2347 ;
  assign n2353 = n170 & n1274 ;
  assign n2354 = n2353 ^ n170 ;
  assign n2355 = n2354 ^ n170 ;
  assign n2349 = n171 & n820 ;
  assign n2350 = n2349 ^ n171 ;
  assign n2351 = n2350 ^ n820 ;
  assign n2352 = n2351 ^ n171 ;
  assign n2356 = n2355 ^ n2352 ;
  assign n2360 = n155 & n1291 ;
  assign n2361 = n2360 ^ n155 ;
  assign n2362 = n2361 ^ n155 ;
  assign n2357 = n139 & n1326 ;
  assign n2358 = n2357 ^ n139 ;
  assign n2359 = n2358 ^ n139 ;
  assign n2363 = n2362 ^ n2359 ;
  assign n2364 = n2356 & n2363 ;
  assign n2365 = n2364 ^ n2363 ;
  assign n2366 = n2365 ^ n2356 ;
  assign n2367 = n2348 & ~n2366 ;
  assign n2368 = n2367 ^ n2348 ;
  assign n2253 = n155 & n1172 ;
  assign n2250 = n139 & n1132 ;
  assign n2251 = n2250 ^ n139 ;
  assign n2252 = n2251 ^ n139 ;
  assign n2254 = n2253 ^ n2252 ;
  assign n2288 = n903 & n1451 ;
  assign n2289 = n2288 ^ n903 ;
  assign n2290 = n2254 & n2289 ;
  assign n2291 = n2290 ^ n2289 ;
  assign n2264 = n155 & n1070 ;
  assign n2263 = n139 & n1036 ;
  assign n2265 = n2264 ^ n2263 ;
  assign n2266 = n137 & n2265 ;
  assign n2267 = n2266 ^ n137 ;
  assign n2272 = x129 & n1045 ;
  assign n2273 = n2272 ^ x129 ;
  assign n2274 = n2273 ^ n1045 ;
  assign n2275 = n2274 ^ n1050 ;
  assign n2277 = n1777 ^ n492 ;
  assign n2276 = x129 & n1051 ;
  assign n2278 = n2277 ^ n2276 ;
  assign n2279 = n2275 & n2278 ;
  assign n2280 = n2279 ^ n2278 ;
  assign n2281 = n2280 ^ n2275 ;
  assign n2282 = n170 & n2281 ;
  assign n2283 = n2282 ^ n170 ;
  assign n2284 = n2283 ^ n170 ;
  assign n2285 = n2267 & n2284 ;
  assign n2286 = n2285 ^ n137 ;
  assign n2268 = n171 & n1114 ;
  assign n2269 = n2268 ^ n1114 ;
  assign n2270 = n2267 & n2269 ;
  assign n2271 = n2270 ^ n2267 ;
  assign n2287 = n2286 ^ n2271 ;
  assign n2292 = n2291 ^ n2287 ;
  assign n2255 = n138 & n170 ;
  assign n2256 = n2255 ^ n170 ;
  assign n2257 = n1151 & n2256 ;
  assign n2258 = n2257 ^ n138 ;
  assign n2259 = n2254 & n2258 ;
  assign n2260 = n2259 ^ n2254 ;
  assign n2261 = n2260 ^ n2258 ;
  assign n2262 = n2261 ^ n138 ;
  assign n2293 = n2292 ^ n2262 ;
  assign n2294 = x134 & n2293 ;
  assign n2295 = n2294 ^ x134 ;
  assign n2330 = n170 & n1195 ;
  assign n2326 = n171 & n969 ;
  assign n2327 = n2326 ^ n171 ;
  assign n2328 = n2327 ^ n969 ;
  assign n2329 = n2328 ^ n171 ;
  assign n2331 = n2330 ^ n2329 ;
  assign n2335 = n155 & n1212 ;
  assign n2332 = n139 & n1247 ;
  assign n2333 = n2332 ^ n139 ;
  assign n2334 = n2333 ^ n139 ;
  assign n2336 = n2335 ^ n2334 ;
  assign n2337 = n2331 & n2336 ;
  assign n2338 = n2337 ^ n2336 ;
  assign n2339 = n2338 ^ n2336 ;
  assign n2340 = n2339 ^ n2331 ;
  assign n2341 = n2340 ^ n2336 ;
  assign n2342 = n136 & n2341 ;
  assign n2343 = n2342 ^ n136 ;
  assign n2344 = n2343 ^ n136 ;
  assign n2345 = n2295 & n2344 ;
  assign n2305 = n170 & n1093 ;
  assign n2306 = n2305 ^ n170 ;
  assign n2307 = n2306 ^ n170 ;
  assign n2296 = n1838 ^ n509 ;
  assign n2297 = n2296 ^ n1017 ;
  assign n2298 = n1015 & n2297 ;
  assign n2299 = n2298 ^ n2297 ;
  assign n2300 = n2299 ^ n1015 ;
  assign n2301 = n171 & n2300 ;
  assign n2302 = n2301 ^ n171 ;
  assign n2303 = n2302 ^ n2300 ;
  assign n2304 = n2303 ^ n171 ;
  assign n2308 = n2307 ^ n2304 ;
  assign n2312 = n155 & n1002 ;
  assign n2313 = n2312 ^ n155 ;
  assign n2314 = n2313 ^ n155 ;
  assign n2309 = n139 & n985 ;
  assign n2310 = n2309 ^ n139 ;
  assign n2311 = n2310 ^ n139 ;
  assign n2315 = n2314 ^ n2311 ;
  assign n2316 = n2308 & n2315 ;
  assign n2317 = n2316 ^ n2315 ;
  assign n2318 = n2317 ^ n2315 ;
  assign n2319 = n2318 ^ n2308 ;
  assign n2320 = n2319 ^ n2315 ;
  assign n2321 = n402 & n2320 ;
  assign n2322 = n2321 ^ n402 ;
  assign n2323 = n2322 ^ n402 ;
  assign n2324 = n2295 & n2323 ;
  assign n2325 = n2324 ^ n2295 ;
  assign n2346 = n2345 ^ n2325 ;
  assign n2369 = n2368 ^ n2346 ;
  assign n2184 = n170 & n782 ;
  assign n2185 = n2184 ^ n170 ;
  assign n2186 = n2185 ^ n170 ;
  assign n2180 = n171 & n736 ;
  assign n2181 = n2180 ^ n171 ;
  assign n2182 = n2181 ^ n736 ;
  assign n2183 = n2182 ^ n171 ;
  assign n2187 = n2186 ^ n2183 ;
  assign n2191 = n155 & n801 ;
  assign n2192 = n2191 ^ n155 ;
  assign n2193 = n2192 ^ n155 ;
  assign n2188 = n139 & n836 ;
  assign n2189 = n2188 ^ n139 ;
  assign n2190 = n2189 ^ n139 ;
  assign n2194 = n2193 ^ n2190 ;
  assign n2195 = n2187 & n2194 ;
  assign n2196 = n2195 ^ n2194 ;
  assign n2197 = n2196 ^ n2194 ;
  assign n2198 = n2197 ^ n2187 ;
  assign n2199 = n2198 ^ n2194 ;
  assign n2200 = n137 & n2199 ;
  assign n2201 = n2200 ^ n137 ;
  assign n2202 = n2201 ^ n137 ;
  assign n2160 = n170 & n698 ;
  assign n2161 = n2160 ^ n170 ;
  assign n2162 = n2161 ^ n170 ;
  assign n2156 = n171 & n1229 ;
  assign n2157 = n2156 ^ n171 ;
  assign n2158 = n2157 ^ n1229 ;
  assign n2159 = n2158 ^ n171 ;
  assign n2163 = n2162 ^ n2159 ;
  assign n2167 = n155 & n717 ;
  assign n2168 = n2167 ^ n155 ;
  assign n2169 = n2168 ^ n155 ;
  assign n2164 = n139 & n754 ;
  assign n2165 = n2164 ^ n139 ;
  assign n2166 = n2165 ^ n139 ;
  assign n2170 = n2169 ^ n2166 ;
  assign n2171 = n2163 & n2170 ;
  assign n2172 = n2171 ^ n2170 ;
  assign n2173 = n2172 ^ n2170 ;
  assign n2174 = n2173 ^ n2163 ;
  assign n2175 = n2174 ^ n2170 ;
  assign n2176 = n138 & n2175 ;
  assign n2177 = n2176 ^ n138 ;
  assign n2178 = n2177 ^ n2175 ;
  assign n2179 = n2178 ^ n138 ;
  assign n2203 = n2202 ^ n2179 ;
  assign n2236 = n2203 ^ x134 ;
  assign n2221 = n865 & n1157 ;
  assign n2208 = n155 & n884 ;
  assign n2209 = n2208 ^ n155 ;
  assign n2210 = n2209 ^ n155 ;
  assign n2205 = n139 & n921 ;
  assign n2206 = n2205 ^ n139 ;
  assign n2207 = n2206 ^ n139 ;
  assign n2211 = n2210 ^ n2207 ;
  assign n2212 = n171 & n1308 ;
  assign n2213 = n2212 ^ n171 ;
  assign n2214 = n2213 ^ n1308 ;
  assign n2215 = n2214 ^ n171 ;
  assign n2216 = n2211 & n2215 ;
  assign n2217 = n2216 ^ n2211 ;
  assign n2218 = n2217 ^ n2211 ;
  assign n2219 = n2218 ^ n2211 ;
  assign n2220 = n2219 ^ n2215 ;
  assign n2222 = n2221 ^ n2220 ;
  assign n2237 = n2222 ^ x134 ;
  assign n2238 = n2222 & n2237 ;
  assign n2239 = n2238 ^ n2222 ;
  assign n2240 = n2239 ^ n2237 ;
  assign n2241 = n2240 ^ n2222 ;
  assign n2242 = n2241 ^ n2237 ;
  assign n2243 = n2242 ^ x134 ;
  assign n2244 = ~n2236 & ~n2243 ;
  assign n2245 = n2244 ^ n2236 ;
  assign n2246 = n2245 ^ n2243 ;
  assign n2247 = n2246 ^ n2242 ;
  assign n2248 = n2247 ^ n2203 ;
  assign n2204 = n2203 ^ n850 ;
  assign n2223 = n2222 ^ n850 ;
  assign n2224 = n2222 & n2223 ;
  assign n2225 = n2224 ^ n2222 ;
  assign n2226 = n2225 ^ n2223 ;
  assign n2227 = n2226 ^ n2222 ;
  assign n2228 = n2227 ^ n850 ;
  assign n2229 = ~n2204 & ~n2228 ;
  assign n2230 = n2229 ^ n2204 ;
  assign n2231 = n2230 ^ n2228 ;
  assign n2232 = n2231 ^ n2204 ;
  assign n2233 = n2232 ^ n2228 ;
  assign n2234 = n2233 ^ n2227 ;
  assign n2235 = n2234 ^ n2203 ;
  assign n2249 = n2248 ^ n2235 ;
  assign n2370 = n2369 ^ n2249 ;
  assign n2464 = n155 & ~n1492 ;
  assign n2465 = n2464 ^ n155 ;
  assign n2460 = n170 & n421 ;
  assign n2461 = n2460 ^ n170 ;
  assign n2458 = n170 & n1447 ;
  assign n2459 = n2458 ^ n170 ;
  assign n2462 = n2461 ^ n2459 ;
  assign n2457 = ~n171 & n1340 ;
  assign n2463 = n2462 ^ n2457 ;
  assign n2466 = n2465 ^ n2463 ;
  assign n2456 = n139 & n1442 ;
  assign n2467 = n2466 ^ n2456 ;
  assign n2468 = ~n138 & n2467 ;
  assign n2443 = n155 & n482 ;
  assign n2444 = n2443 ^ n155 ;
  assign n2441 = n155 & n1546 ;
  assign n2442 = n2441 ^ n155 ;
  assign n2445 = n2444 ^ n2442 ;
  assign n2440 = n139 & n1536 ;
  assign n2446 = n2445 ^ n2440 ;
  assign n2447 = n137 & n2446 ;
  assign n2448 = n2447 ^ n137 ;
  assign n2452 = n170 & n1542 ;
  assign n2453 = n2448 & n2452 ;
  assign n2454 = n2453 ^ n137 ;
  assign n2449 = ~n171 & n1437 ;
  assign n2450 = n2448 & n2449 ;
  assign n2451 = n2450 ^ n2448 ;
  assign n2455 = n2454 ^ n2451 ;
  assign n2469 = n2468 ^ n2455 ;
  assign n2485 = n155 & n1461 ;
  assign n2484 = n139 & n1473 ;
  assign n2486 = n2485 ^ n2484 ;
  assign n2487 = n136 & n2486 ;
  assign n2488 = n2487 ^ n136 ;
  assign n2492 = n1463 ^ n617 ;
  assign n2493 = n170 & n2492 ;
  assign n2494 = n2488 & n2493 ;
  assign n2495 = n2494 ^ n136 ;
  assign n2489 = ~n171 & n1505 ;
  assign n2490 = n2488 & n2489 ;
  assign n2491 = n2490 ^ n2488 ;
  assign n2496 = n2495 ^ n2491 ;
  assign n2479 = n155 & ~n1501 ;
  assign n2480 = n2479 ^ n155 ;
  assign n2475 = n170 & n554 ;
  assign n2476 = n2475 ^ n170 ;
  assign n2473 = n170 & n1555 ;
  assign n2474 = n2473 ^ n170 ;
  assign n2477 = n2476 ^ n2474 ;
  assign n2471 = ~n171 & ~n1527 ;
  assign n2472 = n2471 ^ n171 ;
  assign n2478 = n2477 ^ n2472 ;
  assign n2481 = n2480 ^ n2478 ;
  assign n2470 = n139 & n1510 ;
  assign n2482 = n2481 ^ n2470 ;
  assign n2483 = n402 & ~n2482 ;
  assign n2497 = n2496 ^ n2483 ;
  assign n2498 = n2469 & n2497 ;
  assign n2499 = n2498 ^ n2469 ;
  assign n2500 = n2499 ^ n2497 ;
  assign n2501 = x134 & n2500 ;
  assign n2502 = n2501 ^ x134 ;
  assign n2374 = n155 & ~n1400 ;
  assign n2375 = n2374 ^ n155 ;
  assign n2371 = n1381 ^ n160 ;
  assign n2372 = n139 & ~n2371 ;
  assign n2373 = n2372 ^ n139 ;
  assign n2376 = n2375 ^ n2373 ;
  assign n2392 = ~n138 & ~n2376 ;
  assign n2393 = n170 & n1392 ;
  assign n2394 = n2392 & ~n2393 ;
  assign n2383 = n170 & n1407 ;
  assign n2381 = n171 & n1379 ;
  assign n2382 = n2381 ^ n1379 ;
  assign n2384 = n2383 ^ n2382 ;
  assign n2386 = n155 & n1411 ;
  assign n2385 = n139 & n1418 ;
  assign n2387 = n2386 ^ n2385 ;
  assign n2388 = n2384 & n2387 ;
  assign n2389 = n2388 ^ n2384 ;
  assign n2390 = n2389 ^ n2387 ;
  assign n2391 = n137 & n2390 ;
  assign n2395 = n2394 ^ n2391 ;
  assign n2377 = n1475 ^ n647 ;
  assign n2378 = ~n2376 & n2377 ;
  assign n2379 = ~n1451 & n2378 ;
  assign n2380 = n2379 ^ n138 ;
  assign n2396 = n2395 ^ n2380 ;
  assign n2417 = n170 & n1364 ;
  assign n2415 = n171 & n1415 ;
  assign n2416 = n2415 ^ n1415 ;
  assign n2418 = n2417 ^ n2416 ;
  assign n2422 = n139 & n389 ;
  assign n2423 = n2422 ^ n139 ;
  assign n2420 = n139 & n1359 ;
  assign n2421 = n2420 ^ n139 ;
  assign n2424 = n2423 ^ n2421 ;
  assign n2419 = n155 & n1367 ;
  assign n2425 = n2424 ^ n2419 ;
  assign n2426 = n2418 & n2425 ;
  assign n2427 = n2426 ^ n2418 ;
  assign n2428 = n2427 ^ n2425 ;
  assign n2429 = n402 & n2428 ;
  assign n2430 = n2429 ^ n402 ;
  assign n2431 = n2430 ^ n402 ;
  assign n2400 = n155 & n327 ;
  assign n2401 = n2400 ^ n155 ;
  assign n2398 = n155 & n1353 ;
  assign n2399 = n2398 ^ n155 ;
  assign n2402 = n2401 ^ n2399 ;
  assign n2397 = n139 & n1343 ;
  assign n2403 = n2402 ^ n2397 ;
  assign n2404 = n136 & n2403 ;
  assign n2405 = n2404 ^ n136 ;
  assign n2411 = n170 & n1349 ;
  assign n2412 = n2405 & n2411 ;
  assign n2413 = n2412 ^ n136 ;
  assign n2406 = ~n171 & ~n1371 ;
  assign n2407 = n2406 ^ n171 ;
  assign n2408 = n2405 & n2407 ;
  assign n2409 = n2408 ^ n2405 ;
  assign n2410 = n2409 ^ n2405 ;
  assign n2414 = n2413 ^ n2410 ;
  assign n2432 = n2431 ^ n2414 ;
  assign n2433 = x134 & n2432 ;
  assign n2434 = n2433 ^ x134 ;
  assign n2435 = n2434 ^ n2432 ;
  assign n2436 = n2396 & n2435 ;
  assign n2437 = n2436 ^ n2435 ;
  assign n2438 = n2437 ^ n2396 ;
  assign n2439 = n2438 ^ n2435 ;
  assign n2503 = n2502 ^ n2439 ;
  assign n2532 = n170 & n1676 ;
  assign n2533 = n2532 ^ n170 ;
  assign n2534 = n2533 ^ n170 ;
  assign n2528 = n171 & n1601 ;
  assign n2529 = n2528 ^ n171 ;
  assign n2530 = n2529 ^ n1601 ;
  assign n2531 = n2530 ^ n171 ;
  assign n2535 = n2534 ^ n2531 ;
  assign n2539 = n155 & n1687 ;
  assign n2540 = n2539 ^ n155 ;
  assign n2541 = n2540 ^ n155 ;
  assign n2536 = n139 & n1708 ;
  assign n2537 = n2536 ^ n139 ;
  assign n2538 = n2537 ^ n139 ;
  assign n2542 = n2541 ^ n2538 ;
  assign n2543 = n2535 & n2542 ;
  assign n2544 = n2543 ^ n2542 ;
  assign n2545 = n2544 ^ n2542 ;
  assign n2546 = n2545 ^ n2535 ;
  assign n2547 = n2546 ^ n2542 ;
  assign n2548 = n137 & n2547 ;
  assign n2549 = n2548 ^ n137 ;
  assign n2550 = n2549 ^ n137 ;
  assign n2508 = n170 & n1579 ;
  assign n2509 = n2508 ^ n170 ;
  assign n2510 = n2509 ^ n170 ;
  assign n2504 = n171 & n1883 ;
  assign n2505 = n2504 ^ n171 ;
  assign n2506 = n2505 ^ n1883 ;
  assign n2507 = n2506 ^ n171 ;
  assign n2511 = n2510 ^ n2507 ;
  assign n2515 = n155 & n1590 ;
  assign n2516 = n2515 ^ n155 ;
  assign n2517 = n2516 ^ n155 ;
  assign n2512 = n139 & n1611 ;
  assign n2513 = n2512 ^ n139 ;
  assign n2514 = n2513 ^ n139 ;
  assign n2518 = n2517 ^ n2514 ;
  assign n2519 = n2511 & n2518 ;
  assign n2520 = n2519 ^ n2518 ;
  assign n2521 = n2520 ^ n2518 ;
  assign n2522 = n2521 ^ n2511 ;
  assign n2523 = n2522 ^ n2518 ;
  assign n2524 = n138 & n2523 ;
  assign n2525 = n2524 ^ n138 ;
  assign n2526 = n2525 ^ n2523 ;
  assign n2527 = n2526 ^ n138 ;
  assign n2551 = n2550 ^ n2527 ;
  assign n2695 = n170 & n1962 ;
  assign n2696 = n2695 ^ n170 ;
  assign n2697 = n2696 ^ n170 ;
  assign n2691 = n171 & n1698 ;
  assign n2692 = n2691 ^ n171 ;
  assign n2693 = n2692 ^ n1698 ;
  assign n2694 = n2693 ^ n171 ;
  assign n2698 = n2697 ^ n2694 ;
  assign n2700 = n155 & n1973 ;
  assign n2701 = n2700 ^ n155 ;
  assign n2702 = n2701 ^ n155 ;
  assign n2699 = n139 & n1992 ;
  assign n2703 = n2702 ^ n2699 ;
  assign n2704 = n2698 & n2703 ;
  assign n2705 = n2704 ^ n2703 ;
  assign n2706 = n2705 ^ n2703 ;
  assign n2707 = n2706 ^ n2698 ;
  assign n2708 = n2707 ^ n2703 ;
  assign n2709 = n1259 & n2708 ;
  assign n2710 = n2709 ^ n1259 ;
  assign n2711 = n2710 ^ n1259 ;
  assign n2712 = ~n2551 & n2711 ;
  assign n2713 = n2712 ^ n2711 ;
  assign n2714 = n2713 ^ n2711 ;
  assign n2599 = n155 & n1826 ;
  assign n2598 = n139 & n1757 ;
  assign n2600 = n2599 ^ n2598 ;
  assign n2637 = n1451 & n1649 ;
  assign n2638 = n2637 ^ n1649 ;
  assign n2639 = n2600 & n2638 ;
  assign n2640 = n2639 ^ n2638 ;
  assign n2612 = x129 & n170 ;
  assign n2613 = n2612 ^ n170 ;
  assign n2624 = n1102 & n2613 ;
  assign n2621 = n155 & n1792 ;
  assign n2622 = n2621 ^ n155 ;
  assign n2623 = n2622 ^ n155 ;
  assign n2625 = n2624 ^ n2623 ;
  assign n2616 = n170 & n1045 ;
  assign n2617 = n2616 ^ n170 ;
  assign n2618 = n1778 & n2617 ;
  assign n2614 = n451 & n2613 ;
  assign n2615 = n2614 ^ n2613 ;
  assign n2619 = n2618 ^ n2615 ;
  assign n2620 = n2619 ^ n170 ;
  assign n2626 = n2625 ^ n2620 ;
  assign n2627 = n137 & n2626 ;
  assign n2628 = n2627 ^ n137 ;
  assign n2632 = n171 & n1747 ;
  assign n2633 = n2632 ^ n1747 ;
  assign n2634 = n2628 & n2633 ;
  assign n2629 = n139 & n1812 ;
  assign n2630 = n2628 & n2629 ;
  assign n2631 = n2630 ^ n2628 ;
  assign n2635 = n2634 ^ n2631 ;
  assign n2636 = n2635 ^ n137 ;
  assign n2641 = n2640 ^ n2636 ;
  assign n2604 = n138 & n1768 ;
  assign n2605 = n2604 ^ n1768 ;
  assign n2606 = n2605 ^ n138 ;
  assign n2607 = n2600 & n2606 ;
  assign n2608 = n2607 ^ n2600 ;
  assign n2609 = n2608 ^ n2606 ;
  assign n2601 = n1768 & n1827 ;
  assign n2602 = n2600 & n2601 ;
  assign n2603 = n2602 ^ n2601 ;
  assign n2610 = n2609 ^ n2603 ;
  assign n2611 = n2610 ^ n138 ;
  assign n2642 = n2641 ^ n2611 ;
  assign n2643 = x134 & n2642 ;
  assign n2644 = n2643 ^ x134 ;
  assign n2672 = n170 & n1865 ;
  assign n2673 = n2672 ^ n170 ;
  assign n2674 = n2673 ^ n170 ;
  assign n2668 = n171 & n1932 ;
  assign n2669 = n2668 ^ n1932 ;
  assign n2670 = n2669 ^ n171 ;
  assign n2671 = n2670 ^ n171 ;
  assign n2675 = n2674 ^ n2671 ;
  assign n2679 = n155 & n1874 ;
  assign n2680 = n2679 ^ n155 ;
  assign n2681 = n2680 ^ n155 ;
  assign n2676 = n139 & n1893 ;
  assign n2677 = n2676 ^ n139 ;
  assign n2678 = n2677 ^ n139 ;
  assign n2682 = n2681 ^ n2678 ;
  assign n2683 = n2675 & n2682 ;
  assign n2684 = n2683 ^ n2675 ;
  assign n2685 = n2684 ^ n2682 ;
  assign n2686 = n136 & n2685 ;
  assign n2687 = n2686 ^ n136 ;
  assign n2688 = n2687 ^ n136 ;
  assign n2689 = n2644 & n2688 ;
  assign n2649 = n170 & n1914 ;
  assign n2650 = n2649 ^ n170 ;
  assign n2651 = n2650 ^ n170 ;
  assign n2645 = n171 & n1848 ;
  assign n2646 = n2645 ^ n171 ;
  assign n2647 = n2646 ^ n1848 ;
  assign n2648 = n2647 ^ n171 ;
  assign n2652 = n2651 ^ n2648 ;
  assign n2656 = n155 & n1923 ;
  assign n2657 = n2656 ^ n155 ;
  assign n2658 = n2657 ^ n155 ;
  assign n2653 = n139 & n1942 ;
  assign n2654 = n2653 ^ n139 ;
  assign n2655 = n2654 ^ n139 ;
  assign n2659 = n2658 ^ n2655 ;
  assign n2660 = n2652 & n2659 ;
  assign n2661 = n2660 ^ n2659 ;
  assign n2662 = n2661 ^ n2652 ;
  assign n2663 = n402 & n2662 ;
  assign n2664 = n2663 ^ n402 ;
  assign n2665 = n2664 ^ n402 ;
  assign n2666 = n2644 & n2665 ;
  assign n2667 = n2666 ^ n2644 ;
  assign n2690 = n2689 ^ n2667 ;
  assign n2715 = n2714 ^ n2690 ;
  assign n2584 = n2551 ^ x134 ;
  assign n2557 = n170 & n1631 ;
  assign n2558 = n2557 ^ n170 ;
  assign n2559 = n2558 ^ n170 ;
  assign n2553 = n171 & n1984 ;
  assign n2554 = n2553 ^ n171 ;
  assign n2555 = n2554 ^ n1984 ;
  assign n2556 = n2555 ^ n171 ;
  assign n2560 = n2559 ^ n2556 ;
  assign n2564 = n155 & n1640 ;
  assign n2565 = n2564 ^ n155 ;
  assign n2566 = n2565 ^ n155 ;
  assign n2561 = n139 & n1659 ;
  assign n2562 = n2561 ^ n139 ;
  assign n2563 = n2562 ^ n139 ;
  assign n2567 = n2566 ^ n2563 ;
  assign n2568 = n2560 & n2567 ;
  assign n2569 = n2568 ^ n2567 ;
  assign n2570 = n2569 ^ n2560 ;
  assign n2585 = n2570 ^ x134 ;
  assign n2586 = n2570 & n2585 ;
  assign n2587 = n2586 ^ n2570 ;
  assign n2588 = n2587 ^ n2585 ;
  assign n2589 = n2588 ^ n2570 ;
  assign n2590 = n2589 ^ n2585 ;
  assign n2591 = n2590 ^ x134 ;
  assign n2592 = ~n2584 & ~n2591 ;
  assign n2593 = n2592 ^ n2584 ;
  assign n2594 = n2593 ^ n2591 ;
  assign n2595 = n2594 ^ n2590 ;
  assign n2596 = n2595 ^ n2551 ;
  assign n2552 = n2551 ^ n850 ;
  assign n2571 = n2570 ^ n850 ;
  assign n2572 = n2570 & n2571 ;
  assign n2573 = n2572 ^ n2570 ;
  assign n2574 = n2573 ^ n2571 ;
  assign n2575 = n2574 ^ n2570 ;
  assign n2576 = n2575 ^ n850 ;
  assign n2577 = ~n2552 & ~n2576 ;
  assign n2578 = n2577 ^ n2552 ;
  assign n2579 = n2578 ^ n2576 ;
  assign n2580 = n2579 ^ n2552 ;
  assign n2581 = n2580 ^ n2576 ;
  assign n2582 = n2581 ^ n2575 ;
  assign n2583 = n2582 ^ n2551 ;
  assign n2597 = n2596 ^ n2583 ;
  assign n2716 = n2715 ^ n2597 ;
  assign n2730 = n151 & n170 ;
  assign n2731 = n2730 ^ n170 ;
  assign n2732 = n2731 ^ n170 ;
  assign n2728 = n167 & n171 ;
  assign n2729 = n2728 ^ n167 ;
  assign n2733 = n2732 ^ n2729 ;
  assign n2737 = n155 & n218 ;
  assign n2738 = n2737 ^ n155 ;
  assign n2739 = n2738 ^ n155 ;
  assign n2734 = n139 & n234 ;
  assign n2735 = n2734 ^ n139 ;
  assign n2736 = n2735 ^ n139 ;
  assign n2740 = n2739 ^ n2736 ;
  assign n2741 = n2733 & n2740 ;
  assign n2742 = n2741 ^ n2733 ;
  assign n2743 = n2742 ^ n2740 ;
  assign n2744 = n137 & n2743 ;
  assign n2745 = n2744 ^ n137 ;
  assign n2746 = n2745 ^ n137 ;
  assign n2719 = n170 & n654 ;
  assign n2717 = n171 & n667 ;
  assign n2718 = n2717 ^ n667 ;
  assign n2720 = n2719 ^ n2718 ;
  assign n2722 = n155 & n183 ;
  assign n2721 = n139 & n197 ;
  assign n2723 = n2722 ^ n2721 ;
  assign n2724 = n2720 & n2723 ;
  assign n2725 = n2724 ^ n2720 ;
  assign n2726 = n2725 ^ n2723 ;
  assign n2727 = ~n138 & n2726 ;
  assign n2747 = n2746 ^ n2727 ;
  assign n2828 = n2747 ^ n1259 ;
  assign n2833 = n170 & n250 ;
  assign n2834 = n2833 ^ n170 ;
  assign n2835 = n2834 ^ n170 ;
  assign n2829 = n171 & n265 ;
  assign n2830 = n2829 ^ n171 ;
  assign n2831 = n2830 ^ n265 ;
  assign n2832 = n2831 ^ n171 ;
  assign n2836 = n2835 ^ n2832 ;
  assign n2838 = n155 & n356 ;
  assign n2839 = n2838 ^ n155 ;
  assign n2840 = n2839 ^ n155 ;
  assign n2837 = n139 & n369 ;
  assign n2841 = n2840 ^ n2837 ;
  assign n2842 = n2836 & n2841 ;
  assign n2843 = n2842 ^ n2841 ;
  assign n2844 = n2843 ^ n2836 ;
  assign n2845 = n2844 ^ n1259 ;
  assign n2846 = ~n2844 & n2845 ;
  assign n2847 = n2846 ^ n1259 ;
  assign n2848 = ~n2828 & ~n2847 ;
  assign n2849 = n2848 ^ n2846 ;
  assign n2850 = n2849 ^ n2747 ;
  assign n2764 = n155 & n624 ;
  assign n2763 = n139 & n638 ;
  assign n2765 = n2764 ^ n2763 ;
  assign n2785 = n136 & n170 ;
  assign n2786 = n589 & n2785 ;
  assign n2787 = n2765 & n2786 ;
  assign n2788 = n2787 ^ n2786 ;
  assign n2773 = n139 & n402 ;
  assign n2774 = n575 & n2773 ;
  assign n2775 = n2774 ^ n402 ;
  assign n2771 = n155 & n402 ;
  assign n2772 = n561 & n2771 ;
  assign n2776 = n2775 ^ n2772 ;
  assign n2780 = n170 & n520 ;
  assign n2781 = n2776 & n2780 ;
  assign n2782 = n2781 ^ n2776 ;
  assign n2777 = n171 & n2776 ;
  assign n2778 = n2777 ^ n2776 ;
  assign n2779 = n541 & n2778 ;
  assign n2783 = n2782 ^ n2779 ;
  assign n2784 = n2783 ^ x133 ;
  assign n2789 = n2788 ^ n2784 ;
  assign n2766 = n136 & ~n171 ;
  assign n2767 = n602 & n2766 ;
  assign n2768 = n2767 ^ n136 ;
  assign n2769 = n2765 & n2768 ;
  assign n2770 = n2769 ^ n2768 ;
  assign n2790 = n2789 ^ n2770 ;
  assign n2807 = n2790 ^ x134 ;
  assign n2809 = n171 & n304 ;
  assign n2810 = n2809 ^ n171 ;
  assign n2811 = n2810 ^ n304 ;
  assign n2812 = n2811 ^ n171 ;
  assign n2808 = n170 & n291 ;
  assign n2813 = n2812 ^ n2808 ;
  assign n2815 = n155 & n428 ;
  assign n2814 = n139 & n442 ;
  assign n2816 = n2815 ^ n2814 ;
  assign n2817 = ~n2813 & n2816 ;
  assign n2818 = n2817 ^ n2813 ;
  assign n2819 = n1175 & n2818 ;
  assign n2820 = n2819 ^ x134 ;
  assign n2821 = n2820 ^ x134 ;
  assign n2822 = n2807 & n2821 ;
  assign n2823 = n2822 ^ n2807 ;
  assign n2824 = n2823 ^ n2821 ;
  assign n2825 = n2824 ^ n2820 ;
  assign n2826 = n2825 ^ n2790 ;
  assign n2791 = x134 & n2790 ;
  assign n2792 = n2791 ^ x134 ;
  assign n2795 = n170 & n456 ;
  assign n2793 = n171 & n469 ;
  assign n2794 = n2793 ^ n469 ;
  assign n2796 = n2795 ^ n2794 ;
  assign n2798 = n155 & n503 ;
  assign n2797 = n139 & n489 ;
  assign n2799 = n2798 ^ n2797 ;
  assign n2800 = n2796 & n2799 ;
  assign n2801 = n2800 ^ n2796 ;
  assign n2802 = n2801 ^ n2799 ;
  assign n2803 = n137 & ~n2802 ;
  assign n2804 = n2803 ^ n137 ;
  assign n2805 = n2792 & n2804 ;
  assign n2806 = n2805 ^ n2792 ;
  assign n2827 = n2826 ^ n2806 ;
  assign n2851 = n2850 ^ n2827 ;
  assign n2748 = ~x134 & n136 ;
  assign n2751 = n170 & n383 ;
  assign n2749 = n171 & n396 ;
  assign n2750 = n2749 ^ n396 ;
  assign n2752 = n2751 ^ n2750 ;
  assign n2754 = n155 & n320 ;
  assign n2753 = n139 & n334 ;
  assign n2755 = n2754 ^ n2753 ;
  assign n2756 = n2752 & n2755 ;
  assign n2757 = n2756 ^ n2752 ;
  assign n2758 = n2757 ^ n2755 ;
  assign n2759 = n2748 & n2758 ;
  assign n2760 = n2759 ^ x134 ;
  assign n2761 = n2747 & ~n2760 ;
  assign n2762 = n2761 ^ n2760 ;
  assign n2852 = n2851 ^ n2762 ;
  assign n2881 = n170 & n736 ;
  assign n2882 = n2881 ^ n170 ;
  assign n2883 = n2882 ^ n170 ;
  assign n2877 = n171 & n754 ;
  assign n2878 = n2877 ^ n171 ;
  assign n2879 = n2878 ^ n754 ;
  assign n2880 = n2879 ^ n171 ;
  assign n2884 = n2883 ^ n2880 ;
  assign n2888 = n155 & n782 ;
  assign n2889 = n2888 ^ n155 ;
  assign n2890 = n2889 ^ n155 ;
  assign n2885 = n139 & n801 ;
  assign n2886 = n2885 ^ n139 ;
  assign n2887 = n2886 ^ n139 ;
  assign n2891 = n2890 ^ n2887 ;
  assign n2892 = n2884 & n2891 ;
  assign n2893 = n2892 ^ n2891 ;
  assign n2894 = n2893 ^ n2891 ;
  assign n2895 = n2894 ^ n2884 ;
  assign n2896 = n2895 ^ n2891 ;
  assign n2897 = n137 & n2896 ;
  assign n2898 = n2897 ^ n137 ;
  assign n2899 = n2898 ^ n137 ;
  assign n2857 = n170 & n1229 ;
  assign n2858 = n2857 ^ n170 ;
  assign n2859 = n2858 ^ n170 ;
  assign n2853 = n171 & n1247 ;
  assign n2854 = n2853 ^ n171 ;
  assign n2855 = n2854 ^ n1247 ;
  assign n2856 = n2855 ^ n171 ;
  assign n2860 = n2859 ^ n2856 ;
  assign n2864 = n155 & n698 ;
  assign n2865 = n2864 ^ n155 ;
  assign n2866 = n2865 ^ n155 ;
  assign n2861 = n139 & n717 ;
  assign n2862 = n2861 ^ n139 ;
  assign n2863 = n2862 ^ n139 ;
  assign n2867 = n2866 ^ n2863 ;
  assign n2868 = n2860 & n2867 ;
  assign n2869 = n2868 ^ n2867 ;
  assign n2870 = n2869 ^ n2867 ;
  assign n2871 = n2870 ^ n2860 ;
  assign n2872 = n2871 ^ n2867 ;
  assign n2873 = n138 & n2872 ;
  assign n2874 = n2873 ^ n138 ;
  assign n2875 = n2874 ^ n2872 ;
  assign n2876 = n2875 ^ n138 ;
  assign n2900 = n2899 ^ n2876 ;
  assign n3029 = n170 & n820 ;
  assign n3025 = n171 & n836 ;
  assign n3026 = n3025 ^ n171 ;
  assign n3027 = n3026 ^ n836 ;
  assign n3028 = n3027 ^ n171 ;
  assign n3030 = n3029 ^ n3028 ;
  assign n3032 = n155 & n1274 ;
  assign n3031 = n139 & n1291 ;
  assign n3033 = n3032 ^ n3031 ;
  assign n3034 = n3030 & n3033 ;
  assign n3035 = n3034 ^ n3033 ;
  assign n3036 = n3035 ^ n3033 ;
  assign n3037 = n3036 ^ n3030 ;
  assign n3038 = n3037 ^ n3033 ;
  assign n3039 = n1259 & n3038 ;
  assign n3040 = n3039 ^ n1259 ;
  assign n3041 = n3040 ^ n1259 ;
  assign n3042 = ~n2900 & n3041 ;
  assign n3043 = n3042 ^ n3041 ;
  assign n3044 = n3043 ^ n3041 ;
  assign n2938 = n155 & n1151 ;
  assign n2939 = n2938 ^ n155 ;
  assign n2940 = n2939 ^ n155 ;
  assign n2935 = n139 & n1172 ;
  assign n2936 = n2935 ^ n139 ;
  assign n2937 = n2936 ^ n139 ;
  assign n2941 = n2940 ^ n2937 ;
  assign n2973 = n921 & n1451 ;
  assign n2974 = n2973 ^ n921 ;
  assign n2975 = n2941 & n2974 ;
  assign n2976 = n2975 ^ n2974 ;
  assign n2948 = x129 & n155 ;
  assign n2949 = n2948 ^ n155 ;
  assign n2960 = n492 & n2949 ;
  assign n2959 = n139 & n1070 ;
  assign n2961 = n2960 ^ n2959 ;
  assign n2952 = x47 ^ x46 ;
  assign n2953 = x128 & n2952 ;
  assign n2954 = n2953 ^ x47 ;
  assign n2955 = n2948 & n2954 ;
  assign n2956 = n2955 ^ n2948 ;
  assign n2950 = n1045 & n2949 ;
  assign n2951 = n2950 ^ n2949 ;
  assign n2957 = n2956 ^ n2951 ;
  assign n2958 = n2957 ^ n155 ;
  assign n2962 = n2961 ^ n2958 ;
  assign n2963 = n137 & n2962 ;
  assign n2964 = n2963 ^ n137 ;
  assign n2969 = n170 & n1114 ;
  assign n2970 = n2964 & n2969 ;
  assign n2971 = n2970 ^ n137 ;
  assign n2965 = n171 & n1132 ;
  assign n2966 = n2965 ^ n1132 ;
  assign n2967 = n2964 & n2966 ;
  assign n2968 = n2967 ^ n2964 ;
  assign n2972 = n2971 ^ n2968 ;
  assign n2977 = n2976 ^ n2972 ;
  assign n2942 = n903 & n2256 ;
  assign n2943 = n2942 ^ n138 ;
  assign n2944 = n2941 & n2943 ;
  assign n2945 = n2944 ^ n2941 ;
  assign n2946 = n2945 ^ n2943 ;
  assign n2947 = n2946 ^ n138 ;
  assign n2978 = n2977 ^ n2947 ;
  assign n2982 = n155 & n1195 ;
  assign n2983 = n2982 ^ n155 ;
  assign n2984 = n2983 ^ n155 ;
  assign n2979 = n139 & n1212 ;
  assign n2980 = n2979 ^ n139 ;
  assign n2981 = n2980 ^ n139 ;
  assign n2985 = n2984 ^ n2981 ;
  assign n3013 = n136 & n171 ;
  assign n3014 = n3013 ^ n136 ;
  assign n3015 = n985 & n3014 ;
  assign n3016 = n2985 & n3015 ;
  assign n3017 = n3016 ^ n3015 ;
  assign n3002 = ~n170 & n402 ;
  assign n2998 = n509 & n2613 ;
  assign n2996 = n171 & n1036 ;
  assign n2997 = n2996 ^ n1036 ;
  assign n2999 = n2998 ^ n2997 ;
  assign n3000 = n402 & n2999 ;
  assign n3001 = n3000 ^ n402 ;
  assign n3003 = n3002 ^ n3001 ;
  assign n2991 = n170 & n1017 ;
  assign n2992 = n2991 ^ n170 ;
  assign n2993 = n402 & n1015 ;
  assign n2994 = n2993 ^ n402 ;
  assign n2995 = n2992 & n2994 ;
  assign n3004 = n3003 ^ n2995 ;
  assign n3005 = n3004 ^ n402 ;
  assign n3009 = n155 & n1093 ;
  assign n3010 = n3005 & n3009 ;
  assign n3006 = n139 & n1002 ;
  assign n3007 = n3005 & n3006 ;
  assign n3008 = n3007 ^ n3005 ;
  assign n3011 = n3010 ^ n3008 ;
  assign n3012 = n3011 ^ n402 ;
  assign n3018 = n3017 ^ n3012 ;
  assign n2986 = n969 & n2785 ;
  assign n2987 = n2986 ^ n136 ;
  assign n2988 = n2985 & n2987 ;
  assign n2989 = n2988 ^ n2987 ;
  assign n2990 = n2989 ^ n136 ;
  assign n3019 = n3018 ^ n2990 ;
  assign n3020 = n2978 & n3019 ;
  assign n3021 = n3020 ^ n2978 ;
  assign n3022 = n3021 ^ n3019 ;
  assign n3023 = x134 & n3022 ;
  assign n3024 = n3023 ^ x134 ;
  assign n3045 = n3044 ^ n3024 ;
  assign n2926 = n2900 ^ x134 ;
  assign n2914 = n1157 & n1308 ;
  assign n2905 = n155 & n865 ;
  assign n2906 = n2905 ^ n155 ;
  assign n2907 = n2906 ^ n155 ;
  assign n2902 = n139 & n884 ;
  assign n2903 = n2902 ^ n139 ;
  assign n2904 = n2903 ^ n139 ;
  assign n2908 = n2907 ^ n2904 ;
  assign n2909 = n171 & n1326 ;
  assign n2910 = n2909 ^ n1326 ;
  assign n2911 = n2908 & n2910 ;
  assign n2912 = n2911 ^ n2908 ;
  assign n2913 = n2912 ^ n2910 ;
  assign n2915 = n2914 ^ n2913 ;
  assign n2927 = n2915 ^ x134 ;
  assign n2928 = n2915 & n2927 ;
  assign n2929 = n2928 ^ x134 ;
  assign n2930 = ~n2926 & n2929 ;
  assign n2931 = n2930 ^ n2929 ;
  assign n2932 = n2931 ^ n2928 ;
  assign n2933 = n2932 ^ n2900 ;
  assign n2901 = n2900 ^ n850 ;
  assign n2916 = n2915 ^ n850 ;
  assign n2917 = n2915 & n2916 ;
  assign n2918 = n2917 ^ n2916 ;
  assign n2919 = n2918 ^ n850 ;
  assign n2920 = ~n2901 & n2919 ;
  assign n2921 = n2920 ^ n2919 ;
  assign n2922 = n2921 ^ n2901 ;
  assign n2923 = n2922 ^ n2919 ;
  assign n2924 = n2923 ^ n2918 ;
  assign n2925 = n2924 ^ n2900 ;
  assign n2934 = n2933 ^ n2925 ;
  assign n3046 = n3045 ^ n2934 ;
  assign n3116 = n155 & n1542 ;
  assign n3117 = n3116 ^ n155 ;
  assign n3118 = n3117 ^ n155 ;
  assign n3113 = n139 & n1547 ;
  assign n3114 = n3113 ^ n139 ;
  assign n3115 = n3114 ^ n139 ;
  assign n3119 = n3118 ^ n3115 ;
  assign n3134 = n170 & n1437 ;
  assign n3135 = n137 & ~n3134 ;
  assign n3136 = ~n3119 & n3135 ;
  assign n3129 = n155 & ~n1448 ;
  assign n3130 = n3129 ^ n155 ;
  assign n3127 = n170 & n1340 ;
  assign n3126 = ~n171 & n1343 ;
  assign n3128 = n3127 ^ n3126 ;
  assign n3131 = n3130 ^ n3128 ;
  assign n3124 = n139 & ~n1492 ;
  assign n3125 = n3124 ^ n139 ;
  assign n3132 = n3131 ^ n3125 ;
  assign n3133 = ~n138 & n3132 ;
  assign n3137 = n3136 ^ n3133 ;
  assign n3120 = ~n171 & n1442 ;
  assign n3121 = n137 & n3120 ;
  assign n3122 = ~n3119 & n3121 ;
  assign n3123 = n3122 ^ n137 ;
  assign n3138 = n3137 ^ n3123 ;
  assign n3154 = n155 & n617 ;
  assign n3155 = n3154 ^ n155 ;
  assign n3152 = n155 & n1463 ;
  assign n3153 = n3152 ^ n155 ;
  assign n3156 = n3155 ^ n3153 ;
  assign n3151 = n139 & n1461 ;
  assign n3157 = n3156 ^ n3151 ;
  assign n3158 = n136 & n3157 ;
  assign n3159 = n3158 ^ n136 ;
  assign n3163 = n170 & n1505 ;
  assign n3164 = n3159 & n3163 ;
  assign n3165 = n3164 ^ n136 ;
  assign n3160 = ~n171 & n1510 ;
  assign n3161 = n3159 & n3160 ;
  assign n3162 = n3161 ^ n3159 ;
  assign n3166 = n3165 ^ n3162 ;
  assign n3146 = n155 & ~n1556 ;
  assign n3147 = n3146 ^ n155 ;
  assign n3143 = n170 & ~n1527 ;
  assign n3144 = n3143 ^ n170 ;
  assign n3141 = ~n171 & ~n1536 ;
  assign n3142 = n3141 ^ n171 ;
  assign n3145 = n3144 ^ n3142 ;
  assign n3148 = n3147 ^ n3145 ;
  assign n3139 = n139 & ~n1501 ;
  assign n3140 = n3139 ^ n139 ;
  assign n3149 = n3148 ^ n3140 ;
  assign n3150 = n402 & ~n3149 ;
  assign n3167 = n3166 ^ n3150 ;
  assign n3168 = x134 & n3167 ;
  assign n3169 = n3168 ^ x134 ;
  assign n3170 = n3138 & n3169 ;
  assign n3171 = n3170 ^ n3169 ;
  assign n3050 = n155 & n1349 ;
  assign n3051 = n3050 ^ n155 ;
  assign n3052 = n3051 ^ n155 ;
  assign n3047 = n139 & n1354 ;
  assign n3048 = n3047 ^ n139 ;
  assign n3049 = n3048 ^ n139 ;
  assign n3053 = n3052 ^ n3049 ;
  assign n3069 = n1371 & n2785 ;
  assign n3070 = n3069 ^ n136 ;
  assign n3071 = n3053 & n3070 ;
  assign n3072 = n3071 ^ n3070 ;
  assign n3060 = n170 & n1415 ;
  assign n3058 = n171 & n1418 ;
  assign n3059 = n3058 ^ n1418 ;
  assign n3061 = n3060 ^ n3059 ;
  assign n3063 = n155 & n1364 ;
  assign n3062 = n139 & n1367 ;
  assign n3064 = n3063 ^ n3062 ;
  assign n3065 = n3061 & n3064 ;
  assign n3066 = n3065 ^ n3061 ;
  assign n3067 = n3066 ^ n3064 ;
  assign n3068 = n402 & n3067 ;
  assign n3073 = n3072 ^ n3068 ;
  assign n3054 = n1360 & n3014 ;
  assign n3055 = n3053 & n3054 ;
  assign n3056 = n3055 ^ n3054 ;
  assign n3057 = n3056 ^ n136 ;
  assign n3074 = n3073 ^ n3057 ;
  assign n3092 = n160 & n171 ;
  assign n3093 = n3092 ^ n171 ;
  assign n3094 = n3093 ^ n160 ;
  assign n3089 = n171 & n1381 ;
  assign n3090 = n3089 ^ n171 ;
  assign n3091 = n3090 ^ n1381 ;
  assign n3095 = n3094 ^ n3091 ;
  assign n3088 = n170 & n1379 ;
  assign n3096 = n3095 ^ n3088 ;
  assign n3098 = n155 & n1407 ;
  assign n3097 = n139 & n1411 ;
  assign n3099 = n3098 ^ n3097 ;
  assign n3100 = n3096 & n3099 ;
  assign n3101 = n3100 ^ n3096 ;
  assign n3102 = n3101 ^ n3099 ;
  assign n3103 = n137 & n3102 ;
  assign n3104 = n3103 ^ n137 ;
  assign n3105 = n3104 ^ n137 ;
  assign n3083 = n155 & ~n1392 ;
  assign n3084 = n3083 ^ n155 ;
  assign n3079 = n170 & n647 ;
  assign n3080 = n3079 ^ n170 ;
  assign n3077 = n170 & n1475 ;
  assign n3078 = n3077 ^ n170 ;
  assign n3081 = n3080 ^ n3078 ;
  assign n3076 = ~n171 & n1473 ;
  assign n3082 = n3081 ^ n3076 ;
  assign n3085 = n3084 ^ n3082 ;
  assign n3075 = n139 & n1400 ;
  assign n3086 = n3085 ^ n3075 ;
  assign n3087 = ~n138 & n3086 ;
  assign n3106 = n3105 ^ n3087 ;
  assign n3107 = x134 & n3106 ;
  assign n3108 = n3107 ^ x134 ;
  assign n3109 = n3108 ^ n3106 ;
  assign n3110 = n3074 & n3109 ;
  assign n3111 = n3110 ^ n3074 ;
  assign n3112 = n3111 ^ n3109 ;
  assign n3172 = n3171 ^ n3112 ;
  assign n3197 = n170 & n1601 ;
  assign n3198 = n3197 ^ n170 ;
  assign n3199 = n3198 ^ n170 ;
  assign n3193 = n171 & n1611 ;
  assign n3194 = n3193 ^ n171 ;
  assign n3195 = n3194 ^ n1611 ;
  assign n3196 = n3195 ^ n171 ;
  assign n3200 = n3199 ^ n3196 ;
  assign n3204 = n155 & n1676 ;
  assign n3205 = n3204 ^ n155 ;
  assign n3206 = n3205 ^ n155 ;
  assign n3201 = n139 & n1687 ;
  assign n3202 = n3201 ^ n139 ;
  assign n3203 = n3202 ^ n139 ;
  assign n3207 = n3206 ^ n3203 ;
  assign n3208 = n3200 & n3207 ;
  assign n3209 = n3208 ^ n3207 ;
  assign n3210 = n3209 ^ n3207 ;
  assign n3211 = n3210 ^ n3200 ;
  assign n3212 = n3211 ^ n3207 ;
  assign n3213 = n137 & n3212 ;
  assign n3214 = n3213 ^ n137 ;
  assign n3215 = n3214 ^ n137 ;
  assign n3175 = n170 & n1883 ;
  assign n3176 = n3175 ^ n170 ;
  assign n3177 = n3176 ^ n170 ;
  assign n3173 = n171 & n1893 ;
  assign n3174 = n3173 ^ n1893 ;
  assign n3178 = n3177 ^ n3174 ;
  assign n3182 = n155 & n1579 ;
  assign n3183 = n3182 ^ n155 ;
  assign n3184 = n3183 ^ n155 ;
  assign n3179 = n139 & n1590 ;
  assign n3180 = n3179 ^ n139 ;
  assign n3181 = n3180 ^ n139 ;
  assign n3185 = n3184 ^ n3181 ;
  assign n3186 = n3178 & n3185 ;
  assign n3187 = n3186 ^ n3178 ;
  assign n3188 = n3187 ^ n3185 ;
  assign n3189 = n138 & n3188 ;
  assign n3190 = n3189 ^ n3188 ;
  assign n3191 = n3190 ^ n138 ;
  assign n3192 = n3191 ^ n138 ;
  assign n3216 = n3215 ^ n3192 ;
  assign n3344 = n170 & n1698 ;
  assign n3345 = n3344 ^ n170 ;
  assign n3346 = n3345 ^ n170 ;
  assign n3340 = n171 & n1708 ;
  assign n3341 = n3340 ^ n171 ;
  assign n3342 = n3341 ^ n1708 ;
  assign n3343 = n3342 ^ n171 ;
  assign n3347 = n3346 ^ n3343 ;
  assign n3351 = n155 & n1962 ;
  assign n3352 = n3351 ^ n155 ;
  assign n3353 = n3352 ^ n155 ;
  assign n3348 = n139 & n1973 ;
  assign n3349 = n3348 ^ n139 ;
  assign n3350 = n3349 ^ n139 ;
  assign n3354 = n3353 ^ n3350 ;
  assign n3355 = n3347 & n3354 ;
  assign n3356 = n3355 ^ n3354 ;
  assign n3357 = n3356 ^ n3354 ;
  assign n3358 = n3357 ^ n3347 ;
  assign n3359 = n3358 ^ n3354 ;
  assign n3360 = n1259 & n3359 ;
  assign n3361 = n3360 ^ n1259 ;
  assign n3362 = n3361 ^ n1259 ;
  assign n3363 = n3216 & n3362 ;
  assign n3364 = n3363 ^ n3362 ;
  assign n3262 = n155 & n1768 ;
  assign n3261 = n139 & n1826 ;
  assign n3263 = n3262 ^ n3261 ;
  assign n3300 = ~n1451 & n1659 ;
  assign n3301 = ~n3263 & n3300 ;
  assign n3278 = n1120 & n2613 ;
  assign n3275 = n139 & n1792 ;
  assign n3276 = n3275 ^ n139 ;
  assign n3277 = n3276 ^ n139 ;
  assign n3279 = n3278 ^ n3277 ;
  assign n3270 = n170 & n1100 ;
  assign n3271 = n3270 ^ n170 ;
  assign n3272 = n1744 & n3271 ;
  assign n3273 = n3272 ^ n3271 ;
  assign n3274 = n3273 ^ n170 ;
  assign n3280 = n3279 ^ n3274 ;
  assign n3281 = n137 & n3280 ;
  assign n3282 = n3281 ^ n137 ;
  assign n3287 = n1110 ^ n451 ;
  assign n3288 = n3287 ^ n2273 ;
  assign n3289 = n1103 ^ n1102 ;
  assign n3290 = n3289 ^ n1777 ;
  assign n3291 = n3288 & n3290 ;
  assign n3292 = n3291 ^ n3290 ;
  assign n3293 = n3292 ^ n3288 ;
  assign n3294 = n155 & n3293 ;
  assign n3295 = n3294 ^ n155 ;
  assign n3296 = n3295 ^ n155 ;
  assign n3297 = n3282 & n3296 ;
  assign n3298 = n3297 ^ n137 ;
  assign n3283 = n171 & n1757 ;
  assign n3284 = n3283 ^ n1757 ;
  assign n3285 = n3282 & n3284 ;
  assign n3286 = n3285 ^ n3282 ;
  assign n3299 = n3298 ^ n3286 ;
  assign n3302 = n3301 ^ n3299 ;
  assign n3266 = ~n138 & ~n1649 ;
  assign n3267 = ~n3263 & n3266 ;
  assign n3264 = n1649 & n1827 ;
  assign n3265 = ~n3263 & n3264 ;
  assign n3268 = n3267 ^ n3265 ;
  assign n3269 = n3268 ^ n138 ;
  assign n3303 = n3302 ^ n3269 ;
  assign n3327 = n170 & n1932 ;
  assign n3325 = n171 & n1942 ;
  assign n3326 = n3325 ^ n1942 ;
  assign n3328 = n3327 ^ n3326 ;
  assign n3330 = n155 & n1865 ;
  assign n3329 = n139 & n1874 ;
  assign n3331 = n3330 ^ n3329 ;
  assign n3332 = n3328 & n3331 ;
  assign n3333 = n3332 ^ n3328 ;
  assign n3334 = n3333 ^ n3331 ;
  assign n3335 = n1180 & n3334 ;
  assign n3336 = n3303 & n3335 ;
  assign n3337 = n3336 ^ n3335 ;
  assign n3338 = n3337 ^ n3335 ;
  assign n3308 = n170 & n1848 ;
  assign n3304 = n171 & n1812 ;
  assign n3305 = n3304 ^ n171 ;
  assign n3306 = n3305 ^ n1812 ;
  assign n3307 = n3306 ^ n171 ;
  assign n3309 = n3308 ^ n3307 ;
  assign n3311 = n155 & n1914 ;
  assign n3310 = n139 & n1923 ;
  assign n3312 = n3311 ^ n3310 ;
  assign n3313 = n3309 & n3312 ;
  assign n3314 = n3313 ^ n3312 ;
  assign n3315 = n3314 ^ n3312 ;
  assign n3316 = n3315 ^ n3309 ;
  assign n3317 = n3316 ^ n3312 ;
  assign n3318 = n1949 & n3317 ;
  assign n3319 = n3318 ^ n1949 ;
  assign n3320 = n3319 ^ n1949 ;
  assign n3321 = n3320 ^ x134 ;
  assign n3322 = n3303 & n3321 ;
  assign n3323 = n3322 ^ n3321 ;
  assign n3324 = n3323 ^ n3321 ;
  assign n3339 = n3338 ^ n3324 ;
  assign n3365 = n3364 ^ n3339 ;
  assign n3248 = n3216 ^ x134 ;
  assign n3222 = n170 & n1984 ;
  assign n3223 = n3222 ^ n170 ;
  assign n3224 = n3223 ^ n170 ;
  assign n3218 = n171 & n1992 ;
  assign n3219 = n3218 ^ n171 ;
  assign n3220 = n3219 ^ n1992 ;
  assign n3221 = n3220 ^ n171 ;
  assign n3225 = n3224 ^ n3221 ;
  assign n3229 = n155 & n1631 ;
  assign n3230 = n3229 ^ n155 ;
  assign n3231 = n3230 ^ n155 ;
  assign n3226 = n139 & n1640 ;
  assign n3227 = n3226 ^ n139 ;
  assign n3228 = n3227 ^ n139 ;
  assign n3232 = n3231 ^ n3228 ;
  assign n3233 = n3225 & n3232 ;
  assign n3234 = n3233 ^ n3232 ;
  assign n3235 = n3234 ^ n3225 ;
  assign n3249 = n3235 ^ x134 ;
  assign n3250 = n3235 & n3249 ;
  assign n3251 = n3250 ^ n3235 ;
  assign n3252 = n3251 ^ n3249 ;
  assign n3253 = n3252 ^ n3235 ;
  assign n3254 = n3253 ^ n3249 ;
  assign n3255 = n3254 ^ x134 ;
  assign n3256 = n3248 & ~n3255 ;
  assign n3257 = n3256 ^ n3248 ;
  assign n3258 = n3257 ^ n3254 ;
  assign n3259 = n3258 ^ n3216 ;
  assign n3217 = n3216 ^ n850 ;
  assign n3236 = n3235 ^ n850 ;
  assign n3237 = n3235 & n3236 ;
  assign n3238 = n3237 ^ n3235 ;
  assign n3239 = n3238 ^ n3236 ;
  assign n3240 = n3239 ^ n3235 ;
  assign n3241 = n3240 ^ n850 ;
  assign n3242 = n3217 & ~n3241 ;
  assign n3243 = n3242 ^ n3217 ;
  assign n3244 = n3243 ^ n3217 ;
  assign n3245 = n3244 ^ n3241 ;
  assign n3246 = n3245 ^ n3240 ;
  assign n3247 = n3246 ^ n3216 ;
  assign n3260 = n3259 ^ n3247 ;
  assign n3366 = n3365 ^ n3260 ;
  assign n3384 = n151 & n155 ;
  assign n3385 = n3384 ^ n155 ;
  assign n3386 = n3385 ^ n155 ;
  assign n3381 = n139 & n218 ;
  assign n3382 = n3381 ^ n139 ;
  assign n3383 = n3382 ^ n139 ;
  assign n3387 = n3386 ^ n3383 ;
  assign n3390 = n167 & n170 ;
  assign n3388 = n171 & n197 ;
  assign n3389 = n3388 ^ n197 ;
  assign n3391 = n3390 ^ n3389 ;
  assign n3392 = n3387 & n3391 ;
  assign n3393 = n3392 ^ n3391 ;
  assign n3394 = n3393 ^ n3387 ;
  assign n3395 = n137 & n3394 ;
  assign n3396 = n3395 ^ n137 ;
  assign n3397 = n3396 ^ n137 ;
  assign n3371 = n170 & n667 ;
  assign n3367 = n171 & n638 ;
  assign n3368 = n3367 ^ n171 ;
  assign n3369 = n3368 ^ n638 ;
  assign n3370 = n3369 ^ n171 ;
  assign n3372 = n3371 ^ n3370 ;
  assign n3374 = n155 & n654 ;
  assign n3373 = n139 & n183 ;
  assign n3375 = n3374 ^ n3373 ;
  assign n3376 = n3372 & n3375 ;
  assign n3377 = n3376 ^ n3375 ;
  assign n3378 = n3377 ^ n3372 ;
  assign n3379 = ~n138 & ~n3378 ;
  assign n3380 = n3379 ^ n138 ;
  assign n3398 = n3397 ^ n3380 ;
  assign n3490 = n3398 ^ n1259 ;
  assign n3495 = n170 & n265 ;
  assign n3496 = n3495 ^ n170 ;
  assign n3497 = n3496 ^ n170 ;
  assign n3491 = n171 & n234 ;
  assign n3492 = n3491 ^ n171 ;
  assign n3493 = n3492 ^ n234 ;
  assign n3494 = n3493 ^ n171 ;
  assign n3498 = n3497 ^ n3494 ;
  assign n3502 = n155 & n250 ;
  assign n3503 = n3502 ^ n155 ;
  assign n3504 = n3503 ^ n155 ;
  assign n3499 = n139 & n356 ;
  assign n3500 = n3499 ^ n139 ;
  assign n3501 = n3500 ^ n139 ;
  assign n3505 = n3504 ^ n3501 ;
  assign n3506 = n3498 & n3505 ;
  assign n3507 = n3506 ^ n3505 ;
  assign n3508 = n3507 ^ n3498 ;
  assign n3509 = n3508 ^ n1259 ;
  assign n3510 = ~n3508 & n3509 ;
  assign n3511 = n3510 ^ n1259 ;
  assign n3512 = n3490 & ~n3511 ;
  assign n3513 = n3512 ^ n3510 ;
  assign n3514 = n3513 ^ n3398 ;
  assign n3426 = n561 & n2773 ;
  assign n3427 = n3426 ^ n402 ;
  assign n3425 = n520 & n2771 ;
  assign n3428 = n3427 ^ n3425 ;
  assign n3431 = n170 & n3428 ;
  assign n3432 = n541 & n3431 ;
  assign n3433 = n3432 ^ n3431 ;
  assign n3434 = n3433 ^ n3431 ;
  assign n3435 = n3434 ^ n3428 ;
  assign n3429 = ~n171 & n489 ;
  assign n3430 = n3428 & n3429 ;
  assign n3436 = n3435 ^ n3430 ;
  assign n3437 = n3436 ^ x133 ;
  assign n3415 = n170 & n602 ;
  assign n3413 = n171 & n575 ;
  assign n3414 = n3413 ^ n575 ;
  assign n3416 = n3415 ^ n3414 ;
  assign n3418 = n155 & n589 ;
  assign n3417 = n139 & n624 ;
  assign n3419 = n3418 ^ n3417 ;
  assign n3420 = n3416 & n3419 ;
  assign n3421 = n3420 ^ n3416 ;
  assign n3422 = n3421 ^ n3419 ;
  assign n3423 = n136 & n3422 ;
  assign n3424 = n3423 ^ n136 ;
  assign n3438 = n3437 ^ n3424 ;
  assign n3472 = n170 & n469 ;
  assign n3470 = n171 & n442 ;
  assign n3471 = n3470 ^ n442 ;
  assign n3473 = n3472 ^ n3471 ;
  assign n3475 = n155 & n456 ;
  assign n3474 = n139 & n503 ;
  assign n3476 = n3475 ^ n3474 ;
  assign n3477 = n3473 & n3476 ;
  assign n3478 = n3477 ^ n3473 ;
  assign n3479 = n3478 ^ n3476 ;
  assign n3480 = n137 & n3479 ;
  assign n3481 = n3480 ^ n137 ;
  assign n3482 = n3438 & n3481 ;
  assign n3483 = n3482 ^ n3481 ;
  assign n3468 = n137 & n3438 ;
  assign n3469 = n3468 ^ n137 ;
  assign n3484 = n3483 ^ n3469 ;
  assign n3442 = n3438 ^ n138 ;
  assign n3445 = n170 & n304 ;
  assign n3446 = n3445 ^ n170 ;
  assign n3447 = n3446 ^ n170 ;
  assign n3443 = n171 & n334 ;
  assign n3444 = n3443 ^ n334 ;
  assign n3448 = n3447 ^ n3444 ;
  assign n3450 = n155 & n291 ;
  assign n3449 = n139 & n428 ;
  assign n3451 = n3450 ^ n3449 ;
  assign n3452 = n3448 & n3451 ;
  assign n3453 = n3452 ^ n3451 ;
  assign n3454 = n3453 ^ n3448 ;
  assign n3455 = n3454 ^ n138 ;
  assign n3456 = n3454 & n3455 ;
  assign n3457 = n3456 ^ n3454 ;
  assign n3458 = n3457 ^ n3454 ;
  assign n3459 = n3458 ^ n138 ;
  assign n3460 = n3442 & n3459 ;
  assign n3461 = n3460 ^ n3442 ;
  assign n3462 = n3461 ^ n3459 ;
  assign n3463 = n3462 ^ n3442 ;
  assign n3464 = n3463 ^ n3459 ;
  assign n3465 = n3464 ^ n3458 ;
  assign n3466 = n3465 ^ n3438 ;
  assign n3439 = n138 & n3438 ;
  assign n3440 = n3439 ^ n3438 ;
  assign n3441 = n3440 ^ n138 ;
  assign n3467 = n3466 ^ n3441 ;
  assign n3485 = n3484 ^ n3467 ;
  assign n3486 = n3485 ^ n3438 ;
  assign n3487 = x134 & ~n3486 ;
  assign n3488 = n3487 ^ x134 ;
  assign n3489 = n3488 ^ x134 ;
  assign n3515 = n3514 ^ n3489 ;
  assign n3401 = n170 & n396 ;
  assign n3399 = n171 & n369 ;
  assign n3400 = n3399 ^ n369 ;
  assign n3402 = n3401 ^ n3400 ;
  assign n3404 = n155 & n383 ;
  assign n3403 = n139 & n320 ;
  assign n3405 = n3404 ^ n3403 ;
  assign n3406 = n3402 & n3405 ;
  assign n3407 = n3406 ^ n3402 ;
  assign n3408 = n3407 ^ n3405 ;
  assign n3409 = n2748 & n3408 ;
  assign n3410 = n3409 ^ x134 ;
  assign n3411 = ~n3398 & ~n3410 ;
  assign n3412 = n3411 ^ n3410 ;
  assign n3516 = n3515 ^ n3412 ;
  assign n3533 = n170 & n754 ;
  assign n3531 = n171 & n717 ;
  assign n3532 = n3531 ^ n717 ;
  assign n3534 = n3533 ^ n3532 ;
  assign n3536 = n155 & n736 ;
  assign n3535 = n139 & n782 ;
  assign n3537 = n3536 ^ n3535 ;
  assign n3538 = n3534 & n3537 ;
  assign n3539 = n3538 ^ n3534 ;
  assign n3540 = n3539 ^ n3537 ;
  assign n3541 = n137 & n3540 ;
  assign n3542 = n3541 ^ n137 ;
  assign n3543 = n3542 ^ n137 ;
  assign n3519 = n170 & n1247 ;
  assign n3517 = n171 & n1212 ;
  assign n3518 = n3517 ^ n1212 ;
  assign n3520 = n3519 ^ n3518 ;
  assign n3522 = n155 & n1229 ;
  assign n3521 = n139 & n698 ;
  assign n3523 = n3522 ^ n3521 ;
  assign n3524 = n3520 & n3523 ;
  assign n3525 = n3524 ^ n3520 ;
  assign n3526 = n3525 ^ n3523 ;
  assign n3527 = n138 & n3526 ;
  assign n3528 = n3527 ^ n138 ;
  assign n3529 = n3528 ^ n3526 ;
  assign n3530 = n3529 ^ n138 ;
  assign n3544 = n3543 ^ n3530 ;
  assign n3644 = n170 & n836 ;
  assign n3645 = n3644 ^ n170 ;
  assign n3646 = n3645 ^ n170 ;
  assign n3640 = n171 & n801 ;
  assign n3641 = n3640 ^ n171 ;
  assign n3642 = n3641 ^ n801 ;
  assign n3643 = n3642 ^ n171 ;
  assign n3647 = n3646 ^ n3643 ;
  assign n3649 = n155 & n820 ;
  assign n3648 = n139 & n1274 ;
  assign n3650 = n3649 ^ n3648 ;
  assign n3651 = n3647 & n3650 ;
  assign n3652 = n3651 ^ n3650 ;
  assign n3653 = n3652 ^ n3650 ;
  assign n3654 = n3653 ^ n3647 ;
  assign n3655 = n3654 ^ n3650 ;
  assign n3656 = n1259 & n3655 ;
  assign n3657 = n3656 ^ n1259 ;
  assign n3658 = n3657 ^ n1259 ;
  assign n3659 = ~n3544 & n3658 ;
  assign n3660 = n3659 ^ n3658 ;
  assign n3661 = n3660 ^ n3658 ;
  assign n3572 = n155 & n969 ;
  assign n3571 = n139 & n1195 ;
  assign n3573 = n3572 ^ n3571 ;
  assign n3593 = n1002 & n2766 ;
  assign n3594 = n3573 & n3593 ;
  assign n3595 = n3594 ^ n3593 ;
  assign n3587 = n155 & n2300 ;
  assign n3588 = n3587 ^ n155 ;
  assign n3589 = n3588 ^ n155 ;
  assign n3584 = n170 & ~n1036 ;
  assign n3585 = n3584 ^ n170 ;
  assign n3582 = ~n171 & ~n1070 ;
  assign n3583 = n3582 ^ n171 ;
  assign n3586 = n3585 ^ n3583 ;
  assign n3590 = n3589 ^ n3586 ;
  assign n3579 = n139 & n1093 ;
  assign n3580 = n3579 ^ n139 ;
  assign n3581 = n3580 ^ n139 ;
  assign n3591 = n3590 ^ n3581 ;
  assign n3592 = n402 & ~n3591 ;
  assign n3596 = n3595 ^ n3592 ;
  assign n3574 = n985 & n2785 ;
  assign n3575 = n3574 ^ n136 ;
  assign n3576 = n3573 & n3575 ;
  assign n3577 = n3576 ^ n3575 ;
  assign n3578 = n3577 ^ n136 ;
  assign n3597 = n3596 ^ n3578 ;
  assign n3631 = ~x130 & x131 ;
  assign n3632 = n903 & n3631 ;
  assign n3625 = n170 & n921 ;
  assign n3623 = n171 & n884 ;
  assign n3624 = n3623 ^ n884 ;
  assign n3626 = n3625 ^ n3624 ;
  assign n3627 = n139 & n1151 ;
  assign n3628 = n3626 & n3627 ;
  assign n3629 = n3628 ^ n3626 ;
  assign n3630 = n3629 ^ n3627 ;
  assign n3633 = n3632 ^ n3630 ;
  assign n3634 = n1175 & n3633 ;
  assign n3635 = n3634 ^ n1175 ;
  assign n3636 = n3635 ^ n1175 ;
  assign n3637 = n3597 & n3636 ;
  assign n3638 = n3637 ^ n3636 ;
  assign n3601 = n155 & n1114 ;
  assign n3598 = n139 & n2281 ;
  assign n3599 = n3598 ^ n139 ;
  assign n3600 = n3599 ^ n139 ;
  assign n3602 = n3601 ^ n3600 ;
  assign n3608 = n170 & n1132 ;
  assign n3609 = n3602 & n3608 ;
  assign n3610 = n3609 ^ n3608 ;
  assign n3603 = n171 & n1172 ;
  assign n3604 = n3603 ^ n1172 ;
  assign n3605 = n3602 & n3604 ;
  assign n3606 = n3605 ^ n3602 ;
  assign n3607 = n3606 ^ n3604 ;
  assign n3611 = n3610 ^ n3607 ;
  assign n3618 = x134 & n3611 ;
  assign n3619 = n3618 ^ x134 ;
  assign n3620 = n3597 & n3619 ;
  assign n3621 = n3620 ^ n3619 ;
  assign n3612 = x134 & ~n137 ;
  assign n3613 = n3611 & n3612 ;
  assign n3614 = n3613 ^ n3612 ;
  assign n3615 = n3614 ^ n3612 ;
  assign n3616 = n3597 & n3615 ;
  assign n3617 = n3616 ^ n3615 ;
  assign n3622 = n3621 ^ n3617 ;
  assign n3639 = n3638 ^ n3622 ;
  assign n3662 = n3661 ^ n3639 ;
  assign n3547 = n170 & n1326 ;
  assign n3545 = n171 & n1291 ;
  assign n3546 = n3545 ^ n1291 ;
  assign n3548 = n3547 ^ n3546 ;
  assign n3552 = n155 & n1308 ;
  assign n3553 = n3552 ^ n155 ;
  assign n3554 = n3553 ^ n155 ;
  assign n3549 = n139 & n865 ;
  assign n3550 = n3549 ^ n139 ;
  assign n3551 = n3550 ^ n139 ;
  assign n3555 = n3554 ^ n3551 ;
  assign n3556 = n3548 & n3555 ;
  assign n3557 = n3556 ^ n3548 ;
  assign n3558 = n3557 ^ n3555 ;
  assign n3563 = x134 & n3558 ;
  assign n3564 = n3563 ^ x134 ;
  assign n3565 = n3564 ^ n3558 ;
  assign n3566 = ~n3544 & n3565 ;
  assign n3567 = n3566 ^ n3544 ;
  assign n3568 = n3567 ^ n3565 ;
  assign n3569 = n3568 ^ n3565 ;
  assign n3559 = n850 & n3558 ;
  assign n3560 = ~n3544 & n3559 ;
  assign n3561 = n3560 ^ n3559 ;
  assign n3562 = n3561 ^ n3559 ;
  assign n3570 = n3569 ^ n3562 ;
  assign n3663 = n3662 ^ n3570 ;
  assign n3717 = n155 & n1437 ;
  assign n3718 = n3717 ^ n155 ;
  assign n3719 = n3718 ^ n155 ;
  assign n3714 = n139 & n1542 ;
  assign n3715 = n3714 ^ n139 ;
  assign n3716 = n3715 ^ n139 ;
  assign n3720 = n3719 ^ n3716 ;
  assign n3756 = n3720 ^ x133 ;
  assign n3757 = n3756 ^ x132 ;
  assign n3758 = n3756 & n3757 ;
  assign n3747 = n170 ^ x133 ;
  assign n3748 = n3747 ^ x132 ;
  assign n3749 = n1442 ^ n170 ;
  assign n3750 = n3749 ^ x132 ;
  assign n3751 = n3748 & n3750 ;
  assign n3752 = n3751 ^ n3750 ;
  assign n3753 = n3720 & n3752 ;
  assign n3754 = n3753 ^ n3752 ;
  assign n3759 = n3758 ^ n3754 ;
  assign n3760 = n3759 ^ n3752 ;
  assign n3761 = n3760 ^ n3757 ;
  assign n3763 = n3758 ^ n3752 ;
  assign n3762 = x133 ^ x132 ;
  assign n3764 = n3763 ^ n3762 ;
  assign n3765 = n3761 & n3764 ;
  assign n3766 = n3765 ^ n3761 ;
  assign n3767 = n3766 ^ n3758 ;
  assign n3755 = n3754 ^ n3752 ;
  assign n3768 = n3767 ^ n3755 ;
  assign n3769 = n3768 ^ n3757 ;
  assign n3728 = n171 & n327 ;
  assign n3729 = n3728 ^ n171 ;
  assign n3730 = n3729 ^ n327 ;
  assign n3725 = n171 & n1353 ;
  assign n3726 = n3725 ^ n171 ;
  assign n3727 = n3726 ^ n1353 ;
  assign n3731 = n3730 ^ n3727 ;
  assign n3724 = n170 & n1343 ;
  assign n3732 = n3731 ^ n3724 ;
  assign n3736 = n139 & n421 ;
  assign n3737 = n3736 ^ n139 ;
  assign n3734 = n139 & n1447 ;
  assign n3735 = n3734 ^ n139 ;
  assign n3738 = n3737 ^ n3735 ;
  assign n3733 = n155 & n1340 ;
  assign n3739 = n3738 ^ n3733 ;
  assign n3740 = n3732 & n3739 ;
  assign n3741 = n3740 ^ n3732 ;
  assign n3742 = n3741 ^ n3739 ;
  assign n3743 = n138 & n3742 ;
  assign n3744 = n3743 ^ n138 ;
  assign n3745 = n3744 ^ n3742 ;
  assign n3746 = n3745 ^ n138 ;
  assign n3770 = n3769 ^ n3746 ;
  assign n3721 = n505 & n1492 ;
  assign n3722 = ~n3720 & n3721 ;
  assign n3723 = n3722 ^ n137 ;
  assign n3771 = n3770 ^ n3723 ;
  assign n3775 = n155 & n1505 ;
  assign n3776 = n3775 ^ n155 ;
  assign n3777 = n3776 ^ n155 ;
  assign n3772 = n139 & n2492 ;
  assign n3773 = n3772 ^ n139 ;
  assign n3774 = n3773 ^ n139 ;
  assign n3778 = n3777 ^ n3774 ;
  assign n3825 = n1501 & n3014 ;
  assign n3826 = ~n3778 & n3825 ;
  assign n3807 = n171 & n482 ;
  assign n3808 = n3807 ^ n171 ;
  assign n3809 = n3808 ^ n482 ;
  assign n3804 = n171 & n1546 ;
  assign n3805 = n3804 ^ n171 ;
  assign n3806 = n3805 ^ n1546 ;
  assign n3810 = n3809 ^ n3806 ;
  assign n3803 = n170 & n1536 ;
  assign n3811 = n3810 ^ n3803 ;
  assign n3815 = n139 & n554 ;
  assign n3816 = n3815 ^ n139 ;
  assign n3813 = n139 & n1555 ;
  assign n3814 = n3813 ^ n139 ;
  assign n3817 = n3816 ^ n3814 ;
  assign n3812 = n155 & n1527 ;
  assign n3818 = n3817 ^ n3812 ;
  assign n3819 = n3811 & n3818 ;
  assign n3820 = n3819 ^ n3811 ;
  assign n3821 = n3820 ^ n3818 ;
  assign n3822 = n402 & n3821 ;
  assign n3823 = n3822 ^ n402 ;
  assign n3824 = n3823 ^ n402 ;
  assign n3827 = n3826 ^ n3824 ;
  assign n3785 = n3778 ^ x133 ;
  assign n3786 = n3785 ^ x132 ;
  assign n3787 = n3785 & n3786 ;
  assign n3788 = n3787 ^ n3785 ;
  assign n3789 = n3788 ^ n3786 ;
  assign n3779 = n1510 ^ n170 ;
  assign n3780 = n3779 ^ x132 ;
  assign n3781 = n3748 & n3780 ;
  assign n3782 = n3778 & n3781 ;
  assign n3783 = n3782 ^ n3781 ;
  assign n3790 = n3789 ^ n3783 ;
  assign n3791 = n3790 ^ n3781 ;
  assign n3792 = n3791 ^ n3786 ;
  assign n3793 = n3789 ^ n3781 ;
  assign n3794 = n3793 ^ n3762 ;
  assign n3795 = n3792 & n3794 ;
  assign n3796 = n3795 ^ n3792 ;
  assign n3797 = n3796 ^ n3794 ;
  assign n3798 = n3797 ^ n3794 ;
  assign n3799 = n3798 ^ n3789 ;
  assign n3784 = n3783 ^ n3781 ;
  assign n3800 = n3799 ^ n3784 ;
  assign n3801 = n3800 ^ n3786 ;
  assign n3802 = n3801 ^ n136 ;
  assign n3828 = n3827 ^ n3802 ;
  assign n3829 = ~n3771 & ~n3828 ;
  assign n3830 = n3829 ^ n3828 ;
  assign n3831 = n3830 ^ n3771 ;
  assign n3832 = n3831 ^ n3771 ;
  assign n3833 = n3832 ^ n3828 ;
  assign n3834 = x134 & n3833 ;
  assign n3675 = n155 & n1379 ;
  assign n3674 = n139 & n1407 ;
  assign n3676 = n3675 ^ n3674 ;
  assign n3677 = n137 & ~n3676 ;
  assign n3680 = n170 & n2371 ;
  assign n3681 = n3677 & n3680 ;
  assign n3682 = n3681 ^ n137 ;
  assign n3678 = ~n171 & n1400 ;
  assign n3679 = n3677 & ~n3678 ;
  assign n3683 = n3682 ^ n3679 ;
  assign n3669 = n155 & ~n2377 ;
  assign n3670 = n3669 ^ n155 ;
  assign n3667 = n170 & n1473 ;
  assign n3666 = ~n171 & n1461 ;
  assign n3668 = n3667 ^ n3666 ;
  assign n3671 = n3670 ^ n3668 ;
  assign n3664 = n139 & ~n1392 ;
  assign n3665 = n3664 ^ n139 ;
  assign n3672 = n3671 ^ n3665 ;
  assign n3673 = ~n138 & n3672 ;
  assign n3684 = n3683 ^ n3673 ;
  assign n3707 = n155 & ~n1371 ;
  assign n3708 = n3707 ^ n155 ;
  assign n3703 = n170 & n389 ;
  assign n3704 = n3703 ^ n170 ;
  assign n3701 = n170 & n1359 ;
  assign n3702 = n3701 ^ n170 ;
  assign n3705 = n3704 ^ n3702 ;
  assign n3700 = ~n171 & n1367 ;
  assign n3706 = n3705 ^ n3700 ;
  assign n3709 = n3708 ^ n3706 ;
  assign n3699 = n139 & n1349 ;
  assign n3710 = n3709 ^ n3699 ;
  assign n3711 = n2748 & n3710 ;
  assign n3712 = ~n3684 & n3711 ;
  assign n3687 = n170 & n1418 ;
  assign n3685 = n171 & n1411 ;
  assign n3686 = n3685 ^ n1411 ;
  assign n3688 = n3687 ^ n3686 ;
  assign n3690 = n155 & n1415 ;
  assign n3689 = n139 & n1364 ;
  assign n3691 = n3690 ^ n3689 ;
  assign n3692 = n3688 & n3691 ;
  assign n3693 = n3692 ^ n3688 ;
  assign n3694 = n3693 ^ n3691 ;
  assign n3695 = n1259 & n3694 ;
  assign n3696 = n3695 ^ x134 ;
  assign n3697 = n3684 & ~n3696 ;
  assign n3698 = n3697 ^ n3696 ;
  assign n3713 = n3712 ^ n3698 ;
  assign n3835 = n3834 ^ n3713 ;
  assign n3852 = n170 & n1611 ;
  assign n3850 = n171 & n1590 ;
  assign n3851 = n3850 ^ n1590 ;
  assign n3853 = n3852 ^ n3851 ;
  assign n3855 = n155 & n1601 ;
  assign n3854 = n139 & n1676 ;
  assign n3856 = n3855 ^ n3854 ;
  assign n3857 = n3853 & n3856 ;
  assign n3858 = n3857 ^ n3853 ;
  assign n3859 = n3858 ^ n3856 ;
  assign n3860 = n137 & n3859 ;
  assign n3861 = n3860 ^ n137 ;
  assign n3862 = n3861 ^ n137 ;
  assign n3838 = n170 & n1893 ;
  assign n3836 = n171 & n1874 ;
  assign n3837 = n3836 ^ n1874 ;
  assign n3839 = n3838 ^ n3837 ;
  assign n3841 = n155 & n1883 ;
  assign n3840 = n139 & n1579 ;
  assign n3842 = n3841 ^ n3840 ;
  assign n3843 = n3839 & n3842 ;
  assign n3844 = n3843 ^ n3839 ;
  assign n3845 = n3844 ^ n3842 ;
  assign n3846 = n138 & n3845 ;
  assign n3847 = n3846 ^ n138 ;
  assign n3848 = n3847 ^ n3845 ;
  assign n3849 = n3848 ^ n138 ;
  assign n3863 = n3862 ^ n3849 ;
  assign n3968 = n170 & n1708 ;
  assign n3969 = n3968 ^ n170 ;
  assign n3970 = n3969 ^ n170 ;
  assign n3964 = n171 & n1687 ;
  assign n3965 = n3964 ^ n171 ;
  assign n3966 = n3965 ^ n1687 ;
  assign n3967 = n3966 ^ n171 ;
  assign n3971 = n3970 ^ n3967 ;
  assign n3975 = n155 & n1698 ;
  assign n3976 = n3975 ^ n155 ;
  assign n3977 = n3976 ^ n155 ;
  assign n3972 = n139 & n1962 ;
  assign n3973 = n3972 ^ n139 ;
  assign n3974 = n3973 ^ n139 ;
  assign n3978 = n3977 ^ n3974 ;
  assign n3979 = n3971 & n3978 ;
  assign n3980 = n3979 ^ n3978 ;
  assign n3981 = n3980 ^ n3978 ;
  assign n3982 = n3981 ^ n3971 ;
  assign n3983 = n3982 ^ n3978 ;
  assign n3984 = n1259 & n3983 ;
  assign n3985 = n3984 ^ n1259 ;
  assign n3986 = n3985 ^ n1259 ;
  assign n3987 = ~n3863 & n3986 ;
  assign n3988 = n3987 ^ n3986 ;
  assign n3989 = n3988 ^ n3986 ;
  assign n3893 = n155 & n1932 ;
  assign n3892 = n139 & n1865 ;
  assign n3894 = n3893 ^ n3892 ;
  assign n3921 = n1923 & n2766 ;
  assign n3922 = n3894 & n3921 ;
  assign n3923 = n3922 ^ n3921 ;
  assign n3909 = n1064 & n2613 ;
  assign n3905 = n171 & n1792 ;
  assign n3906 = n3905 ^ n171 ;
  assign n3907 = n3906 ^ n171 ;
  assign n3908 = n3907 ^ n1792 ;
  assign n3910 = n3909 ^ n3908 ;
  assign n3900 = n170 & n1802 ;
  assign n3901 = n3900 ^ n170 ;
  assign n3902 = n1809 & n3901 ;
  assign n3903 = n3902 ^ n3901 ;
  assign n3904 = n3903 ^ n170 ;
  assign n3911 = n3910 ^ n3904 ;
  assign n3912 = n402 & n3911 ;
  assign n3913 = n3912 ^ n402 ;
  assign n3917 = n155 & n1848 ;
  assign n3918 = n3913 & n3917 ;
  assign n3914 = n139 & n1914 ;
  assign n3915 = n3913 & n3914 ;
  assign n3916 = n3915 ^ n3913 ;
  assign n3919 = n3918 ^ n3916 ;
  assign n3920 = n3919 ^ n402 ;
  assign n3924 = n3923 ^ n3920 ;
  assign n3895 = n1942 & n2785 ;
  assign n3896 = n3895 ^ n136 ;
  assign n3897 = n3894 & n3896 ;
  assign n3898 = n3897 ^ n3896 ;
  assign n3899 = n3898 ^ n136 ;
  assign n3925 = n3924 ^ n3899 ;
  assign n3956 = n1157 & n1659 ;
  assign n3949 = n155 & n1649 ;
  assign n3948 = n139 & n1768 ;
  assign n3950 = n3949 ^ n3948 ;
  assign n3951 = n171 & n1640 ;
  assign n3952 = n3951 ^ n1640 ;
  assign n3953 = n3950 & n3952 ;
  assign n3954 = n3953 ^ n3950 ;
  assign n3955 = n3954 ^ n3952 ;
  assign n3957 = n3956 ^ n3955 ;
  assign n3958 = n1175 & n3957 ;
  assign n3959 = n3958 ^ n1175 ;
  assign n3960 = n3959 ^ n1175 ;
  assign n3961 = n3925 & n3960 ;
  assign n3962 = n3961 ^ n3960 ;
  assign n3928 = n170 & n1757 ;
  assign n3926 = n171 & n1826 ;
  assign n3927 = n3926 ^ n1826 ;
  assign n3929 = n3928 ^ n3927 ;
  assign n3933 = n155 & n1747 ;
  assign n3930 = n139 & n3293 ;
  assign n3931 = n3930 ^ n139 ;
  assign n3932 = n3931 ^ n139 ;
  assign n3934 = n3933 ^ n3932 ;
  assign n3935 = n3929 & n3934 ;
  assign n3936 = n3935 ^ n3929 ;
  assign n3937 = n3936 ^ n3934 ;
  assign n3943 = x134 & n3937 ;
  assign n3944 = n3943 ^ x134 ;
  assign n3945 = n3925 & n3944 ;
  assign n3946 = n3945 ^ n3944 ;
  assign n3938 = n3612 & n3937 ;
  assign n3939 = n3938 ^ n3612 ;
  assign n3940 = n3939 ^ n3612 ;
  assign n3941 = n3925 & n3940 ;
  assign n3942 = n3941 ^ n3940 ;
  assign n3947 = n3946 ^ n3942 ;
  assign n3963 = n3962 ^ n3947 ;
  assign n3990 = n3989 ^ n3963 ;
  assign n3868 = n170 & n1992 ;
  assign n3864 = n171 & n1973 ;
  assign n3865 = n3864 ^ n171 ;
  assign n3866 = n3865 ^ n1973 ;
  assign n3867 = n3866 ^ n171 ;
  assign n3869 = n3868 ^ n3867 ;
  assign n3871 = n155 & n1984 ;
  assign n3870 = n139 & n1631 ;
  assign n3872 = n3871 ^ n3870 ;
  assign n3873 = n3869 & n3872 ;
  assign n3874 = n3873 ^ n3872 ;
  assign n3875 = n3874 ^ n3872 ;
  assign n3876 = n3875 ^ n3869 ;
  assign n3877 = n3876 ^ n3872 ;
  assign n3884 = x134 & n3877 ;
  assign n3885 = n3884 ^ x134 ;
  assign n3886 = n3885 ^ n3877 ;
  assign n3887 = ~n3863 & n3886 ;
  assign n3888 = n3887 ^ n3863 ;
  assign n3889 = n3888 ^ n3886 ;
  assign n3890 = n3889 ^ n3886 ;
  assign n3878 = n850 & n3877 ;
  assign n3879 = n3878 ^ n850 ;
  assign n3880 = n3879 ^ n850 ;
  assign n3881 = ~n3863 & n3880 ;
  assign n3882 = n3881 ^ n3880 ;
  assign n3883 = n3882 ^ n3880 ;
  assign n3891 = n3890 ^ n3883 ;
  assign n3991 = n3990 ^ n3891 ;
  assign n4038 = n399 ^ n136 ;
  assign n4039 = n1180 ^ n399 ;
  assign n4040 = ~n4038 & ~n4039 ;
  assign n4034 = n137 & n202 ;
  assign n4035 = n4034 ^ n137 ;
  assign n4036 = n4035 ^ n137 ;
  assign n4031 = ~n138 & n672 ;
  assign n4032 = n4031 ^ n138 ;
  assign n4033 = n4032 ^ n138 ;
  assign n4037 = n4036 ^ n4033 ;
  assign n4041 = n4040 ^ n4037 ;
  assign n4042 = n4041 ^ n4038 ;
  assign n4044 = n4037 ^ n136 ;
  assign n4043 = n1180 ^ x134 ;
  assign n4045 = n4044 ^ n4043 ;
  assign n4046 = ~n4042 & n4045 ;
  assign n4047 = n4046 ^ n1180 ;
  assign n4028 = ~x134 & n272 ;
  assign n4029 = n402 & n4028 ;
  assign n4014 = n136 & ~n607 ;
  assign n4015 = n4014 ^ n136 ;
  assign n4026 = n4015 ^ x134 ;
  assign n3996 = n503 & n1553 ;
  assign n3997 = n3996 ^ n402 ;
  assign n3995 = n489 & n1003 ;
  assign n3998 = n3997 ^ n3995 ;
  assign n4000 = n155 & n3998 ;
  assign n4001 = n541 & n4000 ;
  assign n4002 = n4001 ^ n3998 ;
  assign n3999 = n521 & n3998 ;
  assign n4003 = n4002 ^ n3999 ;
  assign n4004 = n4003 ^ x132 ;
  assign n3993 = n137 & ~n474 ;
  assign n3994 = n3993 ^ x133 ;
  assign n4005 = n4004 ^ n3994 ;
  assign n4016 = n4015 ^ n4005 ;
  assign n4017 = n607 & n2748 ;
  assign n4018 = n4017 ^ x134 ;
  assign n4019 = n4018 ^ n4005 ;
  assign n4020 = n4019 ^ x134 ;
  assign n4021 = n4016 & ~n4020 ;
  assign n4022 = n4021 ^ n4016 ;
  assign n4023 = n4022 ^ n4020 ;
  assign n4024 = n4023 ^ n4018 ;
  assign n4006 = n4005 ^ x134 ;
  assign n4007 = n339 & n1175 ;
  assign n4008 = n4007 ^ x134 ;
  assign n4009 = n4006 & n4008 ;
  assign n4010 = n4009 ^ n4006 ;
  assign n4011 = n4010 ^ n4008 ;
  assign n4012 = n4011 ^ n4007 ;
  assign n4013 = n4012 ^ n4005 ;
  assign n4025 = n4024 ^ n4013 ;
  assign n4027 = n4026 ^ n4025 ;
  assign n4030 = n4029 ^ n4027 ;
  assign n4048 = n4047 ^ n4030 ;
  assign n3992 = n136 ^ x134 ;
  assign n4049 = n4048 ^ n3992 ;
  assign n4052 = n137 & n763 ;
  assign n4053 = n4052 ^ n137 ;
  assign n4054 = n4053 ^ n137 ;
  assign n4050 = n138 & n1254 ;
  assign n4051 = n4050 ^ n1254 ;
  assign n4055 = n4054 ^ n4051 ;
  assign n4087 = n845 & n1259 ;
  assign n4088 = n4087 ^ n1259 ;
  assign n4089 = n4088 ^ n1259 ;
  assign n4090 = n4055 & n4089 ;
  assign n4091 = n4090 ^ n4089 ;
  assign n4070 = n1002 & n2785 ;
  assign n4071 = n4070 ^ n136 ;
  assign n4072 = n987 & n4071 ;
  assign n4073 = n4072 ^ n4071 ;
  assign n4067 = n402 & ~n1075 ;
  assign n4068 = ~n1041 & n4067 ;
  assign n4069 = n4068 ^ n402 ;
  assign n4074 = n4073 ^ n4069 ;
  assign n4063 = n1093 & n2766 ;
  assign n4064 = n987 & n4063 ;
  assign n4065 = n4064 ^ n4063 ;
  assign n4066 = n4065 ^ n136 ;
  assign n4075 = n4074 ^ n4066 ;
  assign n4081 = n930 & n1175 ;
  assign n4082 = n4081 ^ n1175 ;
  assign n4083 = n4082 ^ n1175 ;
  assign n4084 = n4075 & n4083 ;
  assign n4085 = n4084 ^ n4083 ;
  assign n4076 = x134 & n137 ;
  assign n4077 = n1174 & n4076 ;
  assign n4078 = n4077 ^ x134 ;
  assign n4079 = n4075 & n4078 ;
  assign n4080 = n4079 ^ n4078 ;
  assign n4086 = n4085 ^ n4080 ;
  assign n4092 = n4091 ^ n4086 ;
  assign n4059 = n1331 & n2748 ;
  assign n4060 = n4055 & n4059 ;
  assign n4061 = n4060 ^ n4059 ;
  assign n4056 = x134 & n4055 ;
  assign n4057 = n4056 ^ x134 ;
  assign n4058 = n4057 ^ n4055 ;
  assign n4062 = n4061 ^ n4058 ;
  assign n4093 = n4092 ^ n4062 ;
  assign n4126 = n137 & n1446 ;
  assign n4127 = n4126 ^ n137 ;
  assign n4128 = n1494 & n4127 ;
  assign n4129 = n4128 ^ n4127 ;
  assign n4116 = n138 & n1345 ;
  assign n4117 = n4116 ^ n1345 ;
  assign n4118 = n4117 ^ n138 ;
  assign n4122 = n1355 & n4118 ;
  assign n4123 = n4122 ^ n1355 ;
  assign n4124 = n4123 ^ n138 ;
  assign n4119 = n1350 & n4118 ;
  assign n4120 = n4119 ^ n1350 ;
  assign n4121 = n4120 ^ n4118 ;
  assign n4125 = n4124 ^ n4121 ;
  assign n4130 = n4129 ^ n4125 ;
  assign n4108 = n1446 ^ n505 ;
  assign n4109 = n1448 ^ n505 ;
  assign n4110 = ~n1448 & n4109 ;
  assign n4111 = n4110 ^ n505 ;
  assign n4112 = ~n4108 & ~n4111 ;
  assign n4113 = n4112 ^ n4110 ;
  assign n4114 = n4113 ^ n1446 ;
  assign n4115 = n4114 ^ n137 ;
  assign n4131 = n4130 ^ n4115 ;
  assign n4147 = n136 & n1514 ;
  assign n4148 = n4147 ^ n136 ;
  assign n4149 = n1503 & n4148 ;
  assign n4150 = n4149 ^ n4148 ;
  assign n4140 = n402 & n1538 ;
  assign n4141 = n4140 ^ n402 ;
  assign n4144 = n1548 & n4141 ;
  assign n4145 = n4144 ^ n402 ;
  assign n4142 = n1543 & n4141 ;
  assign n4143 = n4142 ^ n4141 ;
  assign n4146 = n4145 ^ n4143 ;
  assign n4151 = n4150 ^ n4146 ;
  assign n4132 = n3014 ^ n1556 ;
  assign n4133 = ~n3014 & n4132 ;
  assign n4134 = n4133 ^ n1556 ;
  assign n4135 = n4134 ^ n1514 ;
  assign n4136 = n1514 & ~n4135 ;
  assign n4137 = n4136 ^ n4133 ;
  assign n4138 = n4137 ^ n1556 ;
  assign n4139 = n4138 ^ n136 ;
  assign n4152 = n4151 ^ n4139 ;
  assign n4153 = n4131 & n4152 ;
  assign n4154 = n4153 ^ n4152 ;
  assign n4155 = n4154 ^ n4131 ;
  assign n4156 = n4155 ^ n4152 ;
  assign n4157 = x134 & n4156 ;
  assign n4158 = n4157 ^ x134 ;
  assign n4159 = n4158 ^ x134 ;
  assign n4095 = n137 & ~n1387 ;
  assign n4097 = n1401 & n4095 ;
  assign n4098 = n4097 ^ n137 ;
  assign n4096 = n1394 & n4095 ;
  assign n4099 = n4098 ^ n4096 ;
  assign n4094 = ~n138 & n1484 ;
  assign n4100 = n4099 ^ n4094 ;
  assign n4105 = n1375 & n2748 ;
  assign n4106 = ~n4100 & n4105 ;
  assign n4101 = n1259 & n1423 ;
  assign n4102 = n4101 ^ x134 ;
  assign n4103 = n4100 & ~n4102 ;
  assign n4104 = n4103 ^ n4102 ;
  assign n4107 = n4106 ^ n4104 ;
  assign n4160 = n4159 ^ n4107 ;
  assign n4164 = n138 & n1898 ;
  assign n4165 = n4164 ^ n1898 ;
  assign n4166 = n4165 ^ n138 ;
  assign n4167 = n4166 ^ n138 ;
  assign n4161 = n137 & n1620 ;
  assign n4162 = n4161 ^ n137 ;
  assign n4163 = n4162 ^ n137 ;
  assign n4168 = n4167 ^ n4163 ;
  assign n4217 = n1999 & n2748 ;
  assign n4218 = n4217 ^ n2748 ;
  assign n4219 = n4218 ^ n2748 ;
  assign n4220 = n4168 & n4219 ;
  assign n4221 = n4220 ^ n4219 ;
  assign n4188 = n1923 & n2785 ;
  assign n4189 = n4188 ^ n136 ;
  assign n4190 = n1946 & n4189 ;
  assign n4191 = n4190 ^ n4189 ;
  assign n4179 = n402 & ~n1799 ;
  assign n4182 = n155 & n1812 ;
  assign n4183 = n4182 ^ n155 ;
  assign n4184 = n4183 ^ n155 ;
  assign n4185 = n4179 & n4184 ;
  assign n4180 = n139 & n1848 ;
  assign n4181 = n4179 & ~n4180 ;
  assign n4186 = n4185 ^ n4181 ;
  assign n4187 = n4186 ^ n402 ;
  assign n4192 = n4191 ^ n4187 ;
  assign n4175 = n1914 & n2766 ;
  assign n4176 = n1946 & n4175 ;
  assign n4177 = n4176 ^ n4175 ;
  assign n4178 = n4177 ^ n136 ;
  assign n4193 = n4192 ^ n4178 ;
  assign n4213 = n1175 & n1664 ;
  assign n4214 = n4193 & n4213 ;
  assign n4215 = n4214 ^ n4213 ;
  assign n4198 = n170 & n1826 ;
  assign n4199 = n4198 ^ n170 ;
  assign n4200 = n4199 ^ n170 ;
  assign n4194 = n171 & n1768 ;
  assign n4195 = n4194 ^ n171 ;
  assign n4196 = n4195 ^ n1768 ;
  assign n4197 = n4196 ^ n171 ;
  assign n4201 = n4200 ^ n4197 ;
  assign n4202 = n1761 & n4201 ;
  assign n4203 = n4202 ^ n1761 ;
  assign n4204 = n4203 ^ n1761 ;
  assign n4205 = n4204 ^ n1761 ;
  assign n4206 = n4205 ^ n4201 ;
  assign n4207 = n4076 & n4206 ;
  assign n4208 = n4207 ^ n4076 ;
  assign n4209 = n4208 ^ n4076 ;
  assign n4210 = n4209 ^ x134 ;
  assign n4211 = n4193 & n4210 ;
  assign n4212 = n4211 ^ n4210 ;
  assign n4216 = n4215 ^ n4212 ;
  assign n4222 = n4221 ^ n4216 ;
  assign n4172 = ~n1715 & n2348 ;
  assign n4173 = n4172 ^ n2348 ;
  assign n4169 = x134 & n4168 ;
  assign n4170 = n4169 ^ x134 ;
  assign n4171 = n4170 ^ n4168 ;
  assign n4174 = n4173 ^ n4171 ;
  assign n4223 = n4222 ^ n4174 ;
  assign n4230 = n137 & n2017 ;
  assign n4231 = n4230 ^ n137 ;
  assign n4232 = n4231 ^ n137 ;
  assign n4226 = n138 & n2133 ;
  assign n4227 = n4226 ^ n2133 ;
  assign n4228 = n4227 ^ n138 ;
  assign n4229 = n4228 ^ n138 ;
  assign n4233 = n4232 ^ n4229 ;
  assign n4274 = n1259 & n2039 ;
  assign n4275 = ~n4233 & n4274 ;
  assign n4255 = n320 & n2256 ;
  assign n4256 = n2052 & n4255 ;
  assign n4257 = n4256 ^ n4255 ;
  assign n4246 = n456 & n1553 ;
  assign n4247 = n4246 ^ n402 ;
  assign n4245 = n503 & n1003 ;
  assign n4248 = n4247 ^ n4245 ;
  assign n4251 = n2080 & n4248 ;
  assign n4252 = n4251 ^ n4248 ;
  assign n4249 = n139 & n4248 ;
  assign n4250 = n541 & n4249 ;
  assign n4253 = n4252 ^ n4250 ;
  assign n4254 = n4253 ^ x132 ;
  assign n4258 = n4257 ^ n4254 ;
  assign n4240 = ~n138 & ~n171 ;
  assign n4241 = n383 & n4240 ;
  assign n4242 = n4241 ^ n138 ;
  assign n4243 = n2052 & ~n4242 ;
  assign n4244 = n4243 ^ n4242 ;
  assign n4259 = n4258 ^ n4244 ;
  assign n4265 = n4259 ^ x134 ;
  assign n4266 = n2093 & n4076 ;
  assign n4267 = n4266 ^ x134 ;
  assign n4268 = n4267 ^ x134 ;
  assign n4269 = ~n4265 & n4268 ;
  assign n4270 = n4269 ^ n4265 ;
  assign n4271 = n4270 ^ n4267 ;
  assign n4272 = n4271 ^ n4259 ;
  assign n4260 = x134 & n4259 ;
  assign n4261 = n4260 ^ x134 ;
  assign n4262 = n136 & n2109 ;
  assign n4263 = n4261 & n4262 ;
  assign n4264 = n4263 ^ n4261 ;
  assign n4273 = n4272 ^ n4264 ;
  assign n4276 = n4275 ^ n4273 ;
  assign n4224 = n136 & n2070 ;
  assign n4225 = n4224 ^ n136 ;
  assign n4234 = x134 & n4233 ;
  assign n4235 = n4234 ^ x134 ;
  assign n4236 = n4235 ^ n4233 ;
  assign n4237 = n4225 & n4236 ;
  assign n4238 = n4237 ^ n4225 ;
  assign n4239 = n4238 ^ n4236 ;
  assign n4277 = n4276 ^ n4239 ;
  assign n4282 = n137 & n2175 ;
  assign n4283 = n4282 ^ n137 ;
  assign n4284 = n4283 ^ n137 ;
  assign n4278 = n138 & n2341 ;
  assign n4279 = n4278 ^ n138 ;
  assign n4280 = n4279 ^ n2341 ;
  assign n4281 = n4280 ^ n138 ;
  assign n4285 = n4284 ^ n4281 ;
  assign n4333 = n1259 & n2199 ;
  assign n4334 = n4333 ^ n1259 ;
  assign n4335 = n4334 ^ n1259 ;
  assign n4336 = ~n4285 & n4335 ;
  assign n4337 = n4336 ^ n4335 ;
  assign n4338 = n4337 ^ n4335 ;
  assign n4303 = ~n138 & ~n865 ;
  assign n4304 = ~n2211 & n4303 ;
  assign n4301 = n865 & n1827 ;
  assign n4302 = ~n2211 & n4301 ;
  assign n4305 = n4304 ^ n4302 ;
  assign n4296 = n402 & ~n2265 ;
  assign n4298 = n2284 & n4296 ;
  assign n4299 = n4298 ^ n402 ;
  assign n4297 = ~n2269 & n4296 ;
  assign n4300 = n4299 ^ n4297 ;
  assign n4306 = n4305 ^ n4300 ;
  assign n4293 = n1308 & ~n1451 ;
  assign n4294 = ~n2211 & n4293 ;
  assign n4295 = n4294 ^ n138 ;
  assign n4307 = n4306 ^ n4295 ;
  assign n4316 = n171 & n903 ;
  assign n4317 = n4316 ^ n171 ;
  assign n4318 = n4317 ^ n903 ;
  assign n4319 = n4318 ^ n171 ;
  assign n4315 = n170 & n1151 ;
  assign n4320 = n4319 ^ n4315 ;
  assign n4321 = n2254 & n4320 ;
  assign n4322 = n4321 ^ n2254 ;
  assign n4323 = n4322 ^ n2254 ;
  assign n4324 = n4323 ^ n2254 ;
  assign n4325 = n4324 ^ n4320 ;
  assign n4326 = n4076 & n4325 ;
  assign n4327 = n4326 ^ n4076 ;
  assign n4328 = n4327 ^ n4076 ;
  assign n4329 = n4307 & n4328 ;
  assign n4330 = n4329 ^ n4328 ;
  assign n4331 = n4330 ^ n4328 ;
  assign n4308 = n1180 & n2320 ;
  assign n4309 = n4308 ^ n1180 ;
  assign n4310 = n4309 ^ n1180 ;
  assign n4311 = n4310 ^ x134 ;
  assign n4312 = n4307 & n4311 ;
  assign n4313 = n4312 ^ n4311 ;
  assign n4314 = n4313 ^ n4311 ;
  assign n4332 = n4331 ^ n4314 ;
  assign n4339 = n4338 ^ n4332 ;
  assign n4290 = ~n2366 & n2748 ;
  assign n4291 = n4290 ^ n2748 ;
  assign n4286 = x134 & ~n4285 ;
  assign n4287 = n4286 ^ x134 ;
  assign n4288 = n4287 ^ x134 ;
  assign n4289 = n4288 ^ n4285 ;
  assign n4292 = n4291 ^ n4289 ;
  assign n4340 = n4339 ^ n4292 ;
  assign n4372 = n402 & ~n2446 ;
  assign n4374 = n2452 & n4372 ;
  assign n4375 = n4374 ^ n402 ;
  assign n4373 = ~n2449 & n4372 ;
  assign n4376 = n4375 ^ n4373 ;
  assign n4366 = ~n138 & ~n2403 ;
  assign n4369 = n2411 & n4366 ;
  assign n4370 = n4369 ^ n138 ;
  assign n4367 = ~n2407 & n4366 ;
  assign n4368 = n4367 ^ n4366 ;
  assign n4371 = n4370 ^ n4368 ;
  assign n4377 = n4376 ^ n4371 ;
  assign n4378 = n4377 ^ x134 ;
  assign n4380 = n137 & n2467 ;
  assign n4379 = n136 & ~n2482 ;
  assign n4381 = n4380 ^ n4379 ;
  assign n4382 = n4381 ^ x134 ;
  assign n4383 = n4381 & ~n4382 ;
  assign n4384 = n4383 ^ x134 ;
  assign n4385 = n4378 & ~n4384 ;
  assign n4386 = n4385 ^ n4383 ;
  assign n4387 = n4386 ^ n4377 ;
  assign n4348 = n137 & ~n2376 ;
  assign n4349 = ~n2393 & n4348 ;
  assign n4343 = ~n138 & ~n2486 ;
  assign n4345 = n2493 & n4343 ;
  assign n4346 = n4345 ^ n138 ;
  assign n4344 = ~n2489 & n4343 ;
  assign n4347 = n4346 ^ n4344 ;
  assign n4350 = n4349 ^ n4347 ;
  assign n4341 = n505 & n2378 ;
  assign n4342 = n4341 ^ n137 ;
  assign n4351 = n4350 ^ n4342 ;
  assign n4355 = n402 & n2390 ;
  assign n4356 = n4355 ^ n402 ;
  assign n4357 = n4356 ^ n402 ;
  assign n4352 = n136 & n2428 ;
  assign n4353 = n4352 ^ n136 ;
  assign n4354 = n4353 ^ n136 ;
  assign n4358 = n4357 ^ n4354 ;
  assign n4359 = x134 & n4358 ;
  assign n4360 = n4359 ^ x134 ;
  assign n4361 = n4360 ^ n4358 ;
  assign n4362 = n4351 & n4361 ;
  assign n4363 = n4362 ^ n4351 ;
  assign n4364 = n4363 ^ n4361 ;
  assign n4365 = n4364 ^ n4361 ;
  assign n4388 = n4387 ^ n4365 ;
  assign n4441 = ~x134 & ~n138 ;
  assign n4442 = ~n2685 & n4441 ;
  assign n4443 = n4442 ^ n4441 ;
  assign n4420 = n137 & n1768 ;
  assign n4421 = n4420 ^ n137 ;
  assign n4422 = n2600 & n4421 ;
  assign n4423 = n4422 ^ n4421 ;
  assign n4416 = n137 & ~n170 ;
  assign n4417 = n1768 & n4416 ;
  assign n4418 = n2600 & n4417 ;
  assign n4419 = n4418 ^ n4417 ;
  assign n4424 = n4423 ^ n4419 ;
  assign n4409 = n402 & n2626 ;
  assign n4410 = n4409 ^ n402 ;
  assign n4413 = n2633 & n4410 ;
  assign n4411 = n2629 & n4410 ;
  assign n4412 = n4411 ^ n4410 ;
  assign n4414 = n4413 ^ n4412 ;
  assign n4415 = n4414 ^ n402 ;
  assign n4425 = n4424 ^ n4415 ;
  assign n4405 = n505 & n1649 ;
  assign n4406 = n2600 & n4405 ;
  assign n4407 = n4406 ^ n4405 ;
  assign n4408 = n4407 ^ n137 ;
  assign n4426 = n4425 ^ n4408 ;
  assign n4427 = x134 & n4426 ;
  assign n4428 = n4427 ^ x134 ;
  assign n4434 = n138 & n2570 ;
  assign n4435 = n4434 ^ n138 ;
  assign n4436 = n4435 ^ n2570 ;
  assign n4437 = n4436 ^ n138 ;
  assign n4438 = n4428 & ~n4437 ;
  assign n4439 = n4438 ^ n4428 ;
  assign n4429 = n136 & n2662 ;
  assign n4430 = n4429 ^ n136 ;
  assign n4431 = n4430 ^ n136 ;
  assign n4432 = n4428 & n4431 ;
  assign n4433 = n4432 ^ n4428 ;
  assign n4440 = n4439 ^ n4433 ;
  assign n4444 = n4443 ^ n4440 ;
  assign n4392 = n402 & n2547 ;
  assign n4393 = n4392 ^ n402 ;
  assign n4394 = n4393 ^ n402 ;
  assign n4389 = n137 & n2523 ;
  assign n4390 = n4389 ^ n137 ;
  assign n4391 = n4390 ^ n137 ;
  assign n4395 = n4394 ^ n4391 ;
  assign n4399 = n2708 & n2748 ;
  assign n4400 = n4399 ^ n2748 ;
  assign n4401 = n4400 ^ n2748 ;
  assign n4402 = n4395 & n4401 ;
  assign n4403 = n4402 ^ n4401 ;
  assign n4396 = x134 & n4395 ;
  assign n4397 = n4396 ^ x134 ;
  assign n4398 = n4397 ^ n4395 ;
  assign n4404 = n4403 ^ n4398 ;
  assign n4445 = n4444 ^ n4404 ;
  assign n4493 = n136 & n139 ;
  assign n4494 = n575 & n4493 ;
  assign n4495 = n4494 ^ n136 ;
  assign n4491 = n136 & n155 ;
  assign n4492 = n561 & n4491 ;
  assign n4496 = n4495 ^ n4492 ;
  assign n4502 = n2780 & n4496 ;
  assign n4503 = n4502 ^ n4496 ;
  assign n4497 = n171 & n4496 ;
  assign n4498 = n4497 ^ n4496 ;
  assign n4499 = n541 & n4498 ;
  assign n4500 = n4499 ^ n4498 ;
  assign n4501 = n4500 ^ n4498 ;
  assign n4504 = n4503 ^ n4501 ;
  assign n4505 = n4504 ^ x132 ;
  assign n4487 = n138 & n2758 ;
  assign n4488 = n4487 ^ n138 ;
  assign n4489 = n4488 ^ n2758 ;
  assign n4490 = n4489 ^ x133 ;
  assign n4506 = n4505 ^ n4490 ;
  assign n4515 = x134 & ~n4506 ;
  assign n4516 = n402 & ~n2802 ;
  assign n4517 = n4516 ^ n402 ;
  assign n4518 = n4515 & n4517 ;
  assign n4519 = n4518 ^ n4515 ;
  assign n4520 = n4519 ^ n2818 ;
  assign n4511 = ~n2818 & n4076 ;
  assign n4512 = ~n4506 & n4511 ;
  assign n4507 = n4076 & ~n4506 ;
  assign n4508 = n4507 ^ n137 ;
  assign n4509 = n4508 ^ n2818 ;
  assign n4510 = n4509 ^ n137 ;
  assign n4513 = n4512 ^ n4510 ;
  assign n4480 = n170 & n589 ;
  assign n4478 = n171 & n602 ;
  assign n4479 = n4478 ^ n602 ;
  assign n4481 = n4480 ^ n4479 ;
  assign n4482 = n2765 & n4481 ;
  assign n4483 = n4482 ^ n2765 ;
  assign n4484 = n4483 ^ n4481 ;
  assign n4485 = n4441 & ~n4484 ;
  assign n4486 = n4485 ^ n4441 ;
  assign n4514 = n4513 ^ n4486 ;
  assign n4521 = n4520 ^ n4514 ;
  assign n4457 = n402 & n2743 ;
  assign n4458 = n4457 ^ n402 ;
  assign n4459 = n4458 ^ n402 ;
  assign n4454 = n137 & n2726 ;
  assign n4455 = n4454 ^ n137 ;
  assign n4456 = n4455 ^ n137 ;
  assign n4460 = n4459 ^ n4456 ;
  assign n4467 = n4460 ^ x134 ;
  assign n4468 = n4460 & n4467 ;
  assign n4469 = n4468 ^ n4467 ;
  assign n4446 = n2844 ^ x132 ;
  assign n4461 = n4460 ^ n2844 ;
  assign n4447 = n2844 ^ x134 ;
  assign n4448 = n2844 ^ x133 ;
  assign n4449 = n4448 ^ x134 ;
  assign n4450 = n4447 & n4449 ;
  assign n4451 = n4450 ^ n4447 ;
  assign n4452 = n4451 ^ n4449 ;
  assign n4453 = n4452 ^ x133 ;
  assign n4462 = n4461 ^ n4453 ;
  assign n4463 = n4446 & ~n4462 ;
  assign n4464 = n4463 ^ n4446 ;
  assign n4465 = n4464 ^ n4462 ;
  assign n4466 = n4465 ^ n4462 ;
  assign n4470 = n4469 ^ n4466 ;
  assign n4471 = n4470 ^ n4452 ;
  assign n4472 = n4471 ^ n4449 ;
  assign n4473 = n4469 ^ n4460 ;
  assign n4474 = n4472 & n4473 ;
  assign n4475 = n4474 ^ n4472 ;
  assign n4476 = n4475 ^ n4469 ;
  assign n4477 = n4476 ^ n4460 ;
  assign n4522 = n4521 ^ n4477 ;
  assign n4604 = ~n171 & ~n985 ;
  assign n4605 = n4604 ^ n171 ;
  assign n4602 = n170 & ~n969 ;
  assign n4603 = n4602 ^ n170 ;
  assign n4606 = n4605 ^ n4603 ;
  assign n4607 = n2985 & n4606 ;
  assign n4608 = n4607 ^ n4606 ;
  assign n4609 = n4441 & n4608 ;
  assign n4610 = n4609 ^ n4441 ;
  assign n4561 = n138 & n1308 ;
  assign n4562 = n4561 ^ n1308 ;
  assign n4563 = n4562 ^ n138 ;
  assign n4564 = n2908 & n4563 ;
  assign n4565 = n4564 ^ n2908 ;
  assign n4566 = n4565 ^ n4563 ;
  assign n4558 = n1308 & n1827 ;
  assign n4559 = n2908 & n4558 ;
  assign n4560 = n4559 ^ n4558 ;
  assign n4567 = n4566 ^ n4560 ;
  assign n4549 = n136 & ~n170 ;
  assign n4547 = n136 & n2999 ;
  assign n4548 = n4547 ^ n136 ;
  assign n4550 = n4549 ^ n4548 ;
  assign n4544 = n136 & n1015 ;
  assign n4545 = n4544 ^ n136 ;
  assign n4546 = n2992 & n4545 ;
  assign n4551 = n4550 ^ n4546 ;
  assign n4552 = n4551 ^ n136 ;
  assign n4555 = n3009 & n4552 ;
  assign n4553 = n3006 & n4552 ;
  assign n4554 = n4553 ^ n4552 ;
  assign n4556 = n4555 ^ n4554 ;
  assign n4557 = n4556 ^ n136 ;
  assign n4568 = n4567 ^ n4557 ;
  assign n4539 = n1326 & n1451 ;
  assign n4540 = n4539 ^ n1326 ;
  assign n4541 = n2908 & n4540 ;
  assign n4542 = n4541 ^ n4540 ;
  assign n4543 = n4542 ^ n138 ;
  assign n4569 = n4568 ^ n4543 ;
  assign n4591 = n490 & n903 ;
  assign n4592 = n4591 ^ n137 ;
  assign n4593 = n2941 & n4592 ;
  assign n4594 = n4593 ^ n4592 ;
  assign n4584 = n402 & n2962 ;
  assign n4585 = n4584 ^ n402 ;
  assign n4588 = n2969 & n4585 ;
  assign n4589 = n4588 ^ n402 ;
  assign n4586 = n2966 & n4585 ;
  assign n4587 = n4586 ^ n4585 ;
  assign n4590 = n4589 ^ n4587 ;
  assign n4595 = n4594 ^ n4590 ;
  assign n4596 = n4569 & n4595 ;
  assign n4597 = n4596 ^ n4595 ;
  assign n4581 = n137 & n4569 ;
  assign n4582 = n4581 ^ n137 ;
  assign n4583 = n4582 ^ n4569 ;
  assign n4598 = n4597 ^ n4583 ;
  assign n4570 = n4569 ^ n2941 ;
  assign n4571 = n505 & n921 ;
  assign n4572 = n4571 ^ n2941 ;
  assign n4573 = n4571 & n4572 ;
  assign n4574 = n4573 ^ n4571 ;
  assign n4575 = n4574 ^ n4572 ;
  assign n4576 = n4575 ^ n2941 ;
  assign n4577 = n4570 & n4576 ;
  assign n4578 = n4577 ^ n4570 ;
  assign n4579 = n4578 ^ n4575 ;
  assign n4580 = n4579 ^ n4569 ;
  assign n4599 = n4598 ^ n4580 ;
  assign n4600 = x134 & n4599 ;
  assign n4601 = n4600 ^ x134 ;
  assign n4611 = n4610 ^ n4601 ;
  assign n4526 = n402 & n2896 ;
  assign n4527 = n4526 ^ n402 ;
  assign n4528 = n4527 ^ n402 ;
  assign n4523 = n137 & n2872 ;
  assign n4524 = n4523 ^ n137 ;
  assign n4525 = n4524 ^ n137 ;
  assign n4529 = n4528 ^ n4525 ;
  assign n4533 = n2748 & n3038 ;
  assign n4534 = n4533 ^ n2748 ;
  assign n4535 = n4534 ^ n2748 ;
  assign n4536 = n4529 & n4535 ;
  assign n4537 = n4536 ^ n4535 ;
  assign n4530 = x134 & n4529 ;
  assign n4531 = n4530 ^ x134 ;
  assign n4532 = n4531 ^ n4529 ;
  assign n4538 = n4537 ^ n4532 ;
  assign n4612 = n4611 ^ n4538 ;
  assign n4642 = n1437 ^ n170 ;
  assign n4643 = n4642 ^ x132 ;
  assign n4644 = ~n3748 & ~n4643 ;
  assign n4645 = ~n3119 & n4644 ;
  assign n4653 = n4645 ^ n4644 ;
  assign n4639 = n3119 ^ x133 ;
  assign n4640 = n4639 ^ x132 ;
  assign n4641 = ~n4639 & n4640 ;
  assign n4646 = n4645 ^ n4641 ;
  assign n4647 = n4646 ^ n4644 ;
  assign n4648 = n4647 ^ n4640 ;
  assign n4649 = n4644 ^ n4641 ;
  assign n4650 = n4649 ^ n3762 ;
  assign n4651 = n4648 & ~n4650 ;
  assign n4652 = n4651 ^ n4641 ;
  assign n4654 = n4653 ^ n4652 ;
  assign n4655 = n4654 ^ n4640 ;
  assign n4638 = n137 & n3132 ;
  assign n4656 = n4655 ^ n4638 ;
  assign n4634 = n1442 & n3119 ;
  assign n4635 = n4634 ^ n1442 ;
  assign n4636 = n1553 & n4635 ;
  assign n4637 = n4636 ^ n402 ;
  assign n4657 = n4656 ^ n4637 ;
  assign n4658 = n4657 ^ x134 ;
  assign n4677 = n1451 ^ n1360 ;
  assign n4678 = n4677 ^ n3053 ;
  assign n4670 = ~n1360 & n1451 ;
  assign n4671 = n4670 ^ n1360 ;
  assign n4672 = n4671 ^ n1451 ;
  assign n4673 = n4670 ^ n3053 ;
  assign n4674 = ~n4672 & n4673 ;
  assign n4675 = n4674 ^ n138 ;
  assign n4666 = n136 & ~n3149 ;
  assign n4667 = n4666 ^ n138 ;
  assign n4668 = n4667 ^ n3053 ;
  assign n4659 = n1371 & n2256 ;
  assign n4660 = n4659 ^ n3053 ;
  assign n4661 = n4660 ^ n170 ;
  assign n4662 = n4659 ^ n138 ;
  assign n4663 = n4661 & n4662 ;
  assign n4664 = n4663 ^ n4659 ;
  assign n4665 = n4664 ^ n2255 ;
  assign n4669 = n4668 ^ n4665 ;
  assign n4676 = n4675 ^ n4669 ;
  assign n4679 = n4678 ^ n4676 ;
  assign n4680 = n4679 ^ x134 ;
  assign n4681 = n4679 & ~n4680 ;
  assign n4682 = n4681 ^ x134 ;
  assign n4683 = ~n4658 & ~n4682 ;
  assign n4684 = n4683 ^ n4681 ;
  assign n4685 = n4684 ^ n4657 ;
  assign n4618 = n137 & n3086 ;
  assign n4613 = ~n138 & ~n3157 ;
  assign n4615 = n3163 & n4613 ;
  assign n4616 = n4615 ^ n138 ;
  assign n4614 = ~n3160 & n4613 ;
  assign n4617 = n4616 ^ n4614 ;
  assign n4619 = n4618 ^ n4617 ;
  assign n4623 = n402 & n3102 ;
  assign n4624 = n4623 ^ n402 ;
  assign n4625 = n4624 ^ n402 ;
  assign n4620 = n136 & n3067 ;
  assign n4621 = n4620 ^ n136 ;
  assign n4622 = n4621 ^ n136 ;
  assign n4626 = n4625 ^ n4622 ;
  assign n4627 = x134 & n4626 ;
  assign n4628 = n4627 ^ x134 ;
  assign n4629 = n4628 ^ n4626 ;
  assign n4630 = n4619 & n4629 ;
  assign n4631 = n4630 ^ n4619 ;
  assign n4632 = n4631 ^ n4629 ;
  assign n4633 = n4632 ^ n4629 ;
  assign n4686 = n4685 ^ n4633 ;
  assign n4689 = n137 & n3188 ;
  assign n4687 = n138 & n3334 ;
  assign n4688 = n4687 ^ n3334 ;
  assign n4690 = n4689 ^ n4688 ;
  assign n4743 = n1259 & n3212 ;
  assign n4744 = n4743 ^ n1259 ;
  assign n4745 = n4744 ^ n1259 ;
  assign n4746 = n4690 & n4745 ;
  assign n4747 = n4746 ^ n4745 ;
  assign n4712 = n137 & ~n1649 ;
  assign n4713 = ~n3263 & n4712 ;
  assign n4710 = n1649 & n4416 ;
  assign n4711 = ~n3263 & n4710 ;
  assign n4714 = n4713 ^ n4711 ;
  assign n4703 = n402 & n3280 ;
  assign n4704 = n4703 ^ n402 ;
  assign n4707 = n3296 & n4704 ;
  assign n4708 = n4707 ^ n402 ;
  assign n4705 = n3284 & n4704 ;
  assign n4706 = n4705 ^ n4704 ;
  assign n4709 = n4708 ^ n4706 ;
  assign n4715 = n4714 ^ n4709 ;
  assign n4700 = n505 & n1659 ;
  assign n4701 = ~n3263 & n4700 ;
  assign n4702 = n4701 ^ n137 ;
  assign n4716 = n4715 ^ n4702 ;
  assign n4734 = n1180 & n3317 ;
  assign n4735 = n4734 ^ n1180 ;
  assign n4736 = n4735 ^ n1180 ;
  assign n4737 = n4736 ^ x134 ;
  assign n4738 = n4716 & n4737 ;
  assign n4739 = n4738 ^ n4737 ;
  assign n4740 = n4739 ^ n3235 ;
  assign n4741 = n4740 ^ n138 ;
  assign n4717 = n4716 ^ n138 ;
  assign n4718 = n4717 ^ x134 ;
  assign n4719 = ~x134 & n138 ;
  assign n4720 = n4719 ^ n138 ;
  assign n4721 = n4720 ^ x134 ;
  assign n4722 = n3249 & n4721 ;
  assign n4723 = n4722 ^ n3249 ;
  assign n4724 = n4723 ^ n4721 ;
  assign n4725 = n4724 ^ n4721 ;
  assign n4726 = n4725 ^ n4719 ;
  assign n4727 = n4726 ^ n4716 ;
  assign n4728 = n4727 ^ n3249 ;
  assign n4729 = n4718 & ~n4728 ;
  assign n4730 = n4729 ^ n4728 ;
  assign n4731 = n4730 ^ n4718 ;
  assign n4732 = n4731 ^ n4725 ;
  assign n4733 = n4732 ^ n4719 ;
  assign n4742 = n4741 ^ n4733 ;
  assign n4748 = n4747 ^ n4742 ;
  assign n4694 = n2748 & n3359 ;
  assign n4695 = n4694 ^ n2748 ;
  assign n4696 = n4695 ^ n2748 ;
  assign n4697 = n4690 & n4696 ;
  assign n4698 = n4697 ^ n4696 ;
  assign n4691 = x134 & n4690 ;
  assign n4692 = n4691 ^ x134 ;
  assign n4693 = n4692 ^ n4690 ;
  assign n4699 = n4698 ^ n4693 ;
  assign n4749 = n4748 ^ n4699 ;
  assign n4760 = n137 & n3378 ;
  assign n4761 = n4760 ^ n137 ;
  assign n4762 = n4761 ^ n137 ;
  assign n4758 = n138 & n3422 ;
  assign n4759 = n4758 ^ n3422 ;
  assign n4763 = n4762 ^ n4759 ;
  assign n4810 = n1259 & n3394 ;
  assign n4811 = ~n4763 & n4810 ;
  assign n4786 = n561 & n4493 ;
  assign n4787 = n4786 ^ n136 ;
  assign n4785 = n520 & n4491 ;
  assign n4788 = n4787 ^ n4785 ;
  assign n4790 = n170 & n4788 ;
  assign n4791 = n541 & n4790 ;
  assign n4792 = n4791 ^ n4788 ;
  assign n4789 = n3429 & n4788 ;
  assign n4793 = n4792 ^ n4789 ;
  assign n4794 = n4793 ^ x132 ;
  assign n4781 = n138 & n3408 ;
  assign n4782 = n4781 ^ n138 ;
  assign n4783 = n4782 ^ n3408 ;
  assign n4784 = n4783 ^ x133 ;
  assign n4795 = n4794 ^ n4784 ;
  assign n4801 = n4795 ^ x134 ;
  assign n4802 = n3454 & n4076 ;
  assign n4803 = n4802 ^ x134 ;
  assign n4804 = n4803 ^ x134 ;
  assign n4805 = ~n4801 & n4804 ;
  assign n4806 = n4805 ^ n4801 ;
  assign n4807 = n4806 ^ n4803 ;
  assign n4808 = n4807 ^ n4795 ;
  assign n4796 = x134 & ~n4795 ;
  assign n4797 = n402 & ~n3479 ;
  assign n4798 = n4797 ^ n402 ;
  assign n4799 = n4796 & n4798 ;
  assign n4800 = n4799 ^ n4796 ;
  assign n4809 = n4808 ^ n4800 ;
  assign n4812 = n4811 ^ n4809 ;
  assign n4770 = n4763 ^ x134 ;
  assign n4771 = n4763 & n4770 ;
  assign n4772 = n4771 ^ n4770 ;
  assign n4750 = n3508 ^ x132 ;
  assign n4764 = n4763 ^ n3508 ;
  assign n4751 = n3508 ^ x134 ;
  assign n4752 = n3508 ^ x133 ;
  assign n4753 = n4752 ^ x134 ;
  assign n4754 = n4751 & n4753 ;
  assign n4755 = n4754 ^ n4751 ;
  assign n4756 = n4755 ^ n4753 ;
  assign n4757 = n4756 ^ x133 ;
  assign n4765 = n4764 ^ n4757 ;
  assign n4766 = n4750 & ~n4765 ;
  assign n4767 = n4766 ^ n4750 ;
  assign n4768 = n4767 ^ n4765 ;
  assign n4769 = n4768 ^ n4765 ;
  assign n4773 = n4772 ^ n4769 ;
  assign n4774 = n4773 ^ n4756 ;
  assign n4775 = n4774 ^ n4753 ;
  assign n4776 = n4772 ^ n4763 ;
  assign n4777 = n4775 & n4776 ;
  assign n4778 = n4777 ^ n4775 ;
  assign n4779 = n4778 ^ n4772 ;
  assign n4780 = n4779 ^ n4763 ;
  assign n4813 = n4812 ^ n4780 ;
  assign n4829 = n137 & n3526 ;
  assign n4830 = n4829 ^ n137 ;
  assign n4831 = n4830 ^ n137 ;
  assign n4817 = n171 & n1002 ;
  assign n4818 = n4817 ^ n171 ;
  assign n4819 = n4818 ^ n1002 ;
  assign n4820 = n4819 ^ n171 ;
  assign n4814 = n170 & n985 ;
  assign n4815 = n4814 ^ n170 ;
  assign n4816 = n4815 ^ n170 ;
  assign n4821 = n4820 ^ n4816 ;
  assign n4822 = n3573 & n4821 ;
  assign n4823 = n4822 ^ n3573 ;
  assign n4824 = n4823 ^ n4821 ;
  assign n4825 = n138 & n4824 ;
  assign n4826 = n4825 ^ n138 ;
  assign n4827 = n4826 ^ n4824 ;
  assign n4828 = n4827 ^ n138 ;
  assign n4832 = n4831 ^ n4828 ;
  assign n4869 = n1259 & n3540 ;
  assign n4870 = n4869 ^ n1259 ;
  assign n4871 = n4870 ^ n1259 ;
  assign n4872 = ~n4832 & n4871 ;
  assign n4873 = n4872 ^ n4871 ;
  assign n4874 = n4873 ^ n4871 ;
  assign n4849 = n1326 & n2256 ;
  assign n4850 = n4849 ^ n138 ;
  assign n4851 = n3555 & ~n4850 ;
  assign n4852 = n4851 ^ n4850 ;
  assign n4848 = n136 & ~n3591 ;
  assign n4853 = n4852 ^ n4848 ;
  assign n4844 = n1291 & n4240 ;
  assign n4845 = n3555 & n4844 ;
  assign n4846 = n4845 ^ n4844 ;
  assign n4847 = n4846 ^ n138 ;
  assign n4854 = n4853 ^ n4847 ;
  assign n4863 = n3633 & n4076 ;
  assign n4864 = n4863 ^ n4076 ;
  assign n4865 = n4864 ^ n4076 ;
  assign n4866 = n4854 & n4865 ;
  assign n4867 = n4866 ^ n4865 ;
  assign n4857 = n1949 & n3611 ;
  assign n4858 = n4857 ^ n1949 ;
  assign n4859 = n4858 ^ n1949 ;
  assign n4860 = n4854 & n4859 ;
  assign n4861 = n4860 ^ n4859 ;
  assign n4855 = x134 & n4854 ;
  assign n4856 = n4855 ^ x134 ;
  assign n4862 = n4861 ^ n4856 ;
  assign n4868 = n4867 ^ n4862 ;
  assign n4875 = n4874 ^ n4868 ;
  assign n4837 = n2748 & n3655 ;
  assign n4838 = n4837 ^ n2748 ;
  assign n4839 = n4838 ^ n2748 ;
  assign n4840 = ~n4832 & n4839 ;
  assign n4841 = n4840 ^ n4839 ;
  assign n4842 = n4841 ^ n4839 ;
  assign n4833 = x134 & ~n4832 ;
  assign n4834 = n4833 ^ x134 ;
  assign n4835 = n4834 ^ x134 ;
  assign n4836 = n4835 ^ n4832 ;
  assign n4843 = n4842 ^ n4836 ;
  assign n4876 = n4875 ^ n4843 ;
  assign n4910 = n170 & n1442 ;
  assign n4911 = n402 & ~n4910 ;
  assign n4912 = ~n3720 & n4911 ;
  assign n4909 = n137 & n3742 ;
  assign n4913 = n4912 ^ n4909 ;
  assign n4905 = n1492 & n1553 ;
  assign n4906 = n3720 & n4905 ;
  assign n4907 = n4906 ^ n4905 ;
  assign n4908 = n4907 ^ n402 ;
  assign n4914 = n4913 ^ n4908 ;
  assign n4918 = ~n138 & n3710 ;
  assign n4915 = n136 & n3821 ;
  assign n4916 = n4915 ^ n136 ;
  assign n4917 = n4916 ^ n136 ;
  assign n4919 = n4918 ^ n4917 ;
  assign n4920 = x134 & n4919 ;
  assign n4921 = n4920 ^ x134 ;
  assign n4922 = n4914 & n4921 ;
  assign n4923 = n4922 ^ n4921 ;
  assign n4882 = n170 & n1510 ;
  assign n4883 = ~n138 & ~n4882 ;
  assign n4884 = ~n3778 & n4883 ;
  assign n4881 = n137 & n3672 ;
  assign n4885 = n4884 ^ n4881 ;
  assign n4877 = ~n1451 & n1501 ;
  assign n4878 = n3778 & n4877 ;
  assign n4879 = n4878 ^ n4877 ;
  assign n4880 = n4879 ^ n138 ;
  assign n4886 = n4885 ^ n4880 ;
  assign n4890 = n402 & n3676 ;
  assign n4891 = n4890 ^ n402 ;
  assign n4894 = n3680 & n4891 ;
  assign n4895 = n4894 ^ n402 ;
  assign n4892 = n3678 & n4891 ;
  assign n4893 = n4892 ^ n4891 ;
  assign n4896 = n4895 ^ n4893 ;
  assign n4887 = n136 & n3694 ;
  assign n4888 = n4887 ^ n136 ;
  assign n4889 = n4888 ^ n136 ;
  assign n4897 = n4896 ^ n4889 ;
  assign n4898 = x134 & n4897 ;
  assign n4899 = n4898 ^ x134 ;
  assign n4900 = n4899 ^ n4897 ;
  assign n4901 = n4886 & n4900 ;
  assign n4902 = n4901 ^ n4886 ;
  assign n4903 = n4902 ^ n4900 ;
  assign n4904 = n4903 ^ n4900 ;
  assign n4924 = n4923 ^ n4904 ;
  assign n4936 = n137 & n3845 ;
  assign n4937 = n4936 ^ n137 ;
  assign n4938 = n4937 ^ n137 ;
  assign n4926 = n171 & n1923 ;
  assign n4927 = n4926 ^ n1923 ;
  assign n4925 = n170 & n1942 ;
  assign n4928 = n4927 ^ n4925 ;
  assign n4929 = n3894 & n4928 ;
  assign n4930 = n4929 ^ n3894 ;
  assign n4931 = n4930 ^ n4928 ;
  assign n4932 = n138 & n4931 ;
  assign n4933 = n4932 ^ n138 ;
  assign n4934 = n4933 ^ n4931 ;
  assign n4935 = n4934 ^ n138 ;
  assign n4939 = n4938 ^ n4935 ;
  assign n4982 = n1259 & n3859 ;
  assign n4983 = n4982 ^ n1259 ;
  assign n4984 = n4983 ^ n1259 ;
  assign n4985 = ~n4939 & n4984 ;
  assign n4986 = n4985 ^ n4984 ;
  assign n4987 = n4986 ^ n4984 ;
  assign n4962 = n1992 & n2256 ;
  assign n4963 = n4962 ^ n138 ;
  assign n4964 = n3872 & ~n4963 ;
  assign n4965 = n4964 ^ n4963 ;
  assign n4955 = n136 & n3911 ;
  assign n4956 = n4955 ^ n136 ;
  assign n4959 = n3917 & n4956 ;
  assign n4957 = n3914 & n4956 ;
  assign n4958 = n4957 ^ n4956 ;
  assign n4960 = n4959 ^ n4958 ;
  assign n4961 = n4960 ^ n136 ;
  assign n4966 = n4965 ^ n4961 ;
  assign n4951 = n1973 & n4240 ;
  assign n4952 = n3872 & n4951 ;
  assign n4953 = n4952 ^ n4951 ;
  assign n4954 = n4953 ^ n138 ;
  assign n4967 = n4966 ^ n4954 ;
  assign n4976 = n3957 & n4076 ;
  assign n4977 = n4976 ^ n4076 ;
  assign n4978 = n4977 ^ n4076 ;
  assign n4979 = n4967 & n4978 ;
  assign n4980 = n4979 ^ n4978 ;
  assign n4970 = n1949 & n3937 ;
  assign n4971 = n4970 ^ n1949 ;
  assign n4972 = n4971 ^ n1949 ;
  assign n4973 = n4967 & n4972 ;
  assign n4974 = n4973 ^ n4972 ;
  assign n4968 = x134 & n4967 ;
  assign n4969 = n4968 ^ x134 ;
  assign n4975 = n4974 ^ n4969 ;
  assign n4981 = n4980 ^ n4975 ;
  assign n4988 = n4987 ^ n4981 ;
  assign n4944 = n2748 & n3983 ;
  assign n4945 = n4944 ^ n2748 ;
  assign n4946 = n4945 ^ n2748 ;
  assign n4947 = ~n4939 & n4946 ;
  assign n4948 = n4947 ^ n4946 ;
  assign n4949 = n4948 ^ n4946 ;
  assign n4940 = x134 & ~n4939 ;
  assign n4941 = n4940 ^ x134 ;
  assign n4942 = n4941 ^ x134 ;
  assign n4943 = n4942 ^ n4939 ;
  assign n4950 = n4949 ^ n4943 ;
  assign n4989 = n4988 ^ n4950 ;
  assign n5053 = ~x134 & n202 ;
  assign n5054 = n402 & n5053 ;
  assign n5041 = n402 & n474 ;
  assign n5042 = n5041 ^ n402 ;
  assign n5029 = n136 & n3631 ;
  assign n5030 = n541 & n5029 ;
  assign n5031 = n5030 ^ n5029 ;
  assign n5032 = n5031 ^ n5029 ;
  assign n5025 = n503 & n3014 ;
  assign n5026 = n5025 ^ n136 ;
  assign n5024 = n489 & n2785 ;
  assign n5027 = n5026 ^ n5024 ;
  assign n5033 = n5032 ^ n5027 ;
  assign n5028 = n521 & n5027 ;
  assign n5034 = n5033 ^ n5028 ;
  assign n5043 = n5042 ^ n5034 ;
  assign n5044 = n5043 ^ x133 ;
  assign n5045 = n137 & n339 ;
  assign n5046 = n5044 & n5045 ;
  assign n5047 = n5046 ^ n5045 ;
  assign n5035 = n138 & n5034 ;
  assign n5036 = n5035 ^ n5034 ;
  assign n5037 = n5036 ^ n138 ;
  assign n5038 = n399 & n5037 ;
  assign n5039 = n5038 ^ n399 ;
  assign n5040 = n5039 ^ n5037 ;
  assign n5048 = n5047 ^ n5040 ;
  assign n5049 = n5048 ^ n5044 ;
  assign n5050 = x134 & n5049 ;
  assign n5051 = n5050 ^ x134 ;
  assign n5052 = n5051 ^ x134 ;
  assign n5055 = n5054 ^ n5052 ;
  assign n4995 = n137 & n672 ;
  assign n4996 = n4995 ^ n137 ;
  assign n4997 = n4996 ^ n137 ;
  assign n4991 = n138 & n607 ;
  assign n4992 = n4991 ^ n138 ;
  assign n4993 = n4992 ^ n607 ;
  assign n4994 = n4993 ^ n138 ;
  assign n4998 = n4997 ^ n4994 ;
  assign n5010 = n4998 ^ x134 ;
  assign n5011 = ~n4998 & ~n5010 ;
  assign n5012 = n5011 ^ n4998 ;
  assign n5013 = n5012 ^ n5010 ;
  assign n5014 = n5013 ^ n5010 ;
  assign n4990 = n272 ^ x132 ;
  assign n5000 = n272 ^ x134 ;
  assign n5001 = n272 ^ x133 ;
  assign n5002 = n5001 ^ x134 ;
  assign n5003 = n5000 & n5002 ;
  assign n5004 = n5003 ^ n5002 ;
  assign n5005 = n5004 ^ n5000 ;
  assign n5006 = n5005 ^ x133 ;
  assign n4999 = n4998 ^ n272 ;
  assign n5007 = n5006 ^ n4999 ;
  assign n5008 = n4990 & ~n5007 ;
  assign n5009 = n5008 ^ n4990 ;
  assign n5015 = n5014 ^ n5009 ;
  assign n5016 = n5015 ^ n5005 ;
  assign n5017 = n5016 ^ n5002 ;
  assign n5018 = n5014 ^ n4998 ;
  assign n5019 = n5017 & ~n5018 ;
  assign n5020 = n5019 ^ n5017 ;
  assign n5021 = n5020 ^ n5018 ;
  assign n5022 = n5021 ^ n5014 ;
  assign n5023 = n5022 ^ n4998 ;
  assign n5056 = n5055 ^ n5023 ;
  assign n5072 = n137 & n1254 ;
  assign n5060 = n171 & n1093 ;
  assign n5061 = n5060 ^ n171 ;
  assign n5062 = n5061 ^ n1093 ;
  assign n5063 = n5062 ^ n171 ;
  assign n5057 = n170 & n1002 ;
  assign n5058 = n5057 ^ n170 ;
  assign n5059 = n5058 ^ n170 ;
  assign n5064 = n5063 ^ n5059 ;
  assign n5065 = n987 & n5064 ;
  assign n5066 = n5065 ^ n987 ;
  assign n5067 = n5066 ^ n5064 ;
  assign n5068 = n138 & n5067 ;
  assign n5069 = n5068 ^ n138 ;
  assign n5070 = n5069 ^ n5067 ;
  assign n5071 = n5070 ^ n138 ;
  assign n5073 = n5072 ^ n5071 ;
  assign n5108 = n763 & n1259 ;
  assign n5109 = n5108 ^ n1259 ;
  assign n5110 = n5109 ^ n1259 ;
  assign n5111 = ~n5073 & n5110 ;
  assign n5112 = n5111 ^ n5110 ;
  assign n5113 = n5112 ^ n5110 ;
  assign n5092 = n1291 & n2256 ;
  assign n5093 = n5092 ^ n138 ;
  assign n5094 = n1328 & ~n5093 ;
  assign n5095 = n5094 ^ n5093 ;
  assign n5089 = n136 & ~n1075 ;
  assign n5090 = ~n1041 & n5089 ;
  assign n5091 = n5090 ^ n136 ;
  assign n5096 = n5095 ^ n5091 ;
  assign n5085 = n1274 & n4240 ;
  assign n5086 = n1328 & n5085 ;
  assign n5087 = n5086 ^ n5085 ;
  assign n5088 = n5087 ^ n138 ;
  assign n5097 = n5096 ^ n5088 ;
  assign n5102 = n930 & n4076 ;
  assign n5103 = n5102 ^ n4076 ;
  assign n5104 = n5103 ^ n4076 ;
  assign n5105 = n5097 & n5104 ;
  assign n5106 = n5105 ^ n5104 ;
  assign n5098 = n1174 & n1949 ;
  assign n5099 = n5098 ^ x134 ;
  assign n5100 = n5097 & n5099 ;
  assign n5101 = n5100 ^ n5099 ;
  assign n5107 = n5106 ^ n5101 ;
  assign n5114 = n5113 ^ n5107 ;
  assign n5078 = n845 & n2748 ;
  assign n5079 = n5078 ^ n2748 ;
  assign n5080 = n5079 ^ n2748 ;
  assign n5081 = ~n5073 & n5080 ;
  assign n5082 = n5081 ^ n5080 ;
  assign n5083 = n5082 ^ n5080 ;
  assign n5074 = x134 & ~n5073 ;
  assign n5075 = n5074 ^ x134 ;
  assign n5076 = n5075 ^ x134 ;
  assign n5077 = n5076 ^ n5073 ;
  assign n5084 = n5083 ^ n5077 ;
  assign n5115 = n5114 ^ n5084 ;
  assign n5154 = n1003 & n1492 ;
  assign n5155 = n5154 ^ n402 ;
  assign n5156 = n1446 & n5155 ;
  assign n5157 = n5156 ^ n5155 ;
  assign n5149 = n137 & ~n1345 ;
  assign n5151 = n1355 & n5149 ;
  assign n5152 = n5151 ^ n137 ;
  assign n5150 = ~n1350 & n5149 ;
  assign n5153 = n5152 ^ n5150 ;
  assign n5158 = n5157 ^ n5153 ;
  assign n5145 = n1448 & n1553 ;
  assign n5146 = n1446 & n5145 ;
  assign n5147 = n5146 ^ n5145 ;
  assign n5148 = n5147 ^ n402 ;
  assign n5159 = n5158 ^ n5148 ;
  assign n5167 = ~n138 & n1375 ;
  assign n5160 = n136 & n1538 ;
  assign n5161 = n5160 ^ n136 ;
  assign n5164 = n1548 & n5161 ;
  assign n5165 = n5164 ^ n136 ;
  assign n5162 = n1543 & n5161 ;
  assign n5163 = n5162 ^ n5161 ;
  assign n5166 = n5165 ^ n5163 ;
  assign n5168 = n5167 ^ n5166 ;
  assign n5169 = x134 & n5168 ;
  assign n5170 = n5169 ^ x134 ;
  assign n5171 = n5159 & n5170 ;
  assign n5172 = n5171 ^ n5170 ;
  assign n5121 = n1501 & n2256 ;
  assign n5122 = n5121 ^ n138 ;
  assign n5123 = n1514 & ~n5122 ;
  assign n5124 = n5123 ^ n5122 ;
  assign n5120 = n137 & n1484 ;
  assign n5125 = n5124 ^ n5120 ;
  assign n5116 = ~n1451 & n1556 ;
  assign n5117 = n1514 & n5116 ;
  assign n5118 = n5117 ^ n5116 ;
  assign n5119 = n5118 ^ n138 ;
  assign n5126 = n5125 ^ n5119 ;
  assign n5130 = n402 & n1387 ;
  assign n5131 = n5130 ^ n402 ;
  assign n5135 = n1401 & n5131 ;
  assign n5136 = n5135 ^ n402 ;
  assign n5132 = n1394 & n5131 ;
  assign n5133 = n5132 ^ n5131 ;
  assign n5134 = n5133 ^ n5131 ;
  assign n5137 = n5136 ^ n5134 ;
  assign n5127 = n136 & n1423 ;
  assign n5128 = n5127 ^ n136 ;
  assign n5129 = n5128 ^ n136 ;
  assign n5138 = n5137 ^ n5129 ;
  assign n5139 = x134 & n5138 ;
  assign n5140 = n5139 ^ x134 ;
  assign n5141 = n5140 ^ n5138 ;
  assign n5142 = n5126 & n5141 ;
  assign n5143 = n5142 ^ n5126 ;
  assign n5144 = n5143 ^ n5141 ;
  assign n5173 = n5172 ^ n5144 ;
  assign n5215 = ~n1948 & n4441 ;
  assign n5216 = n5215 ^ n4441 ;
  assign n5197 = n490 & n1640 ;
  assign n5198 = n5197 ^ n137 ;
  assign n5199 = n1661 & n5198 ;
  assign n5200 = n5199 ^ n5198 ;
  assign n5192 = n136 & ~n1799 ;
  assign n5194 = n4184 & n5192 ;
  assign n5193 = ~n4180 & n5192 ;
  assign n5195 = n5194 ^ n5193 ;
  assign n5196 = n5195 ^ n136 ;
  assign n5201 = n5200 ^ n5196 ;
  assign n5187 = n137 & ~n171 ;
  assign n5188 = n1631 & n5187 ;
  assign n5189 = n1661 & n5188 ;
  assign n5190 = n5189 ^ n5188 ;
  assign n5191 = n5190 ^ n137 ;
  assign n5202 = n5201 ^ n5191 ;
  assign n5209 = n1175 & n1999 ;
  assign n5210 = n5209 ^ n1175 ;
  assign n5211 = n5210 ^ n1175 ;
  assign n5212 = n5202 & n5211 ;
  assign n5213 = n5212 ^ n5211 ;
  assign n5203 = n1949 & n4206 ;
  assign n5204 = n5203 ^ n1949 ;
  assign n5205 = n5204 ^ n1949 ;
  assign n5206 = n5205 ^ x134 ;
  assign n5207 = n5202 & n5206 ;
  assign n5208 = n5207 ^ n5206 ;
  assign n5214 = n5213 ^ n5208 ;
  assign n5217 = n5216 ^ n5214 ;
  assign n5184 = ~n1715 & n2748 ;
  assign n5185 = n5184 ^ n2748 ;
  assign n5177 = n137 & n1898 ;
  assign n5178 = n5177 ^ n137 ;
  assign n5179 = n5178 ^ n137 ;
  assign n5174 = n402 & n1620 ;
  assign n5175 = n5174 ^ n402 ;
  assign n5176 = n5175 ^ n402 ;
  assign n5180 = n5179 ^ n5176 ;
  assign n5181 = x134 & n5180 ;
  assign n5182 = n5181 ^ x134 ;
  assign n5183 = n5182 ^ n5180 ;
  assign n5186 = n5185 ^ n5183 ;
  assign n5218 = n5217 ^ n5186 ;
  assign n5230 = n138 & n2103 ;
  assign n5231 = n5230 ^ n2103 ;
  assign n5232 = n5231 ^ n138 ;
  assign n5233 = n2106 & n5232 ;
  assign n5234 = n5233 ^ n2106 ;
  assign n5235 = n5234 ^ n5232 ;
  assign n5236 = n5235 ^ n138 ;
  assign n5227 = n137 & n2133 ;
  assign n5228 = n5227 ^ n137 ;
  assign n5229 = n5228 ^ n137 ;
  assign n5237 = n5236 ^ n5229 ;
  assign n5284 = n1259 & n2017 ;
  assign n5285 = n5237 & n5284 ;
  assign n5286 = n5285 ^ n5284 ;
  assign n5260 = n456 & n3014 ;
  assign n5261 = n5260 ^ n136 ;
  assign n5259 = n503 & n2785 ;
  assign n5262 = n5261 ^ n5259 ;
  assign n5263 = n2080 & n5262 ;
  assign n5264 = n5263 ^ n5262 ;
  assign n5256 = n541 & n4493 ;
  assign n5257 = n5256 ^ n4493 ;
  assign n5258 = n5257 ^ n4493 ;
  assign n5265 = n5264 ^ n5258 ;
  assign n5274 = n5265 ^ x133 ;
  assign n5272 = n402 & n2093 ;
  assign n5273 = n5272 ^ n402 ;
  assign n5275 = n5274 ^ n5273 ;
  assign n5276 = n137 & n2059 ;
  assign n5277 = n5275 & n5276 ;
  assign n5278 = n5277 ^ n5276 ;
  assign n5266 = n138 & n5265 ;
  assign n5267 = n5266 ^ n5265 ;
  assign n5268 = n5267 ^ n138 ;
  assign n5269 = n2070 & n5268 ;
  assign n5270 = n5269 ^ n2070 ;
  assign n5271 = n5270 ^ n5268 ;
  assign n5279 = n5278 ^ n5271 ;
  assign n5280 = n5279 ^ n5275 ;
  assign n5281 = x134 & n5280 ;
  assign n5282 = n5281 ^ x134 ;
  assign n5283 = n5282 ^ x134 ;
  assign n5287 = n5286 ^ n5283 ;
  assign n5243 = n5237 ^ x134 ;
  assign n5244 = n5237 & n5243 ;
  assign n5245 = n5244 ^ n5243 ;
  assign n5219 = n2039 ^ x132 ;
  assign n5238 = n5237 ^ n2039 ;
  assign n5220 = n2039 ^ x134 ;
  assign n5221 = n2039 ^ x133 ;
  assign n5222 = n5221 ^ x134 ;
  assign n5223 = n5220 & n5222 ;
  assign n5224 = n5223 ^ n5220 ;
  assign n5225 = n5224 ^ n5222 ;
  assign n5226 = n5225 ^ x133 ;
  assign n5239 = n5238 ^ n5226 ;
  assign n5240 = n5219 & n5239 ;
  assign n5241 = n5240 ^ n5219 ;
  assign n5242 = n5241 ^ n5219 ;
  assign n5246 = n5245 ^ n5242 ;
  assign n5247 = n5246 ^ n5225 ;
  assign n5248 = n5247 ^ n5222 ;
  assign n5249 = n5245 ^ n5237 ;
  assign n5250 = n5248 & n5249 ;
  assign n5251 = n5250 ^ n5249 ;
  assign n5252 = n5251 ^ n5248 ;
  assign n5253 = n5252 ^ n5249 ;
  assign n5254 = n5253 ^ n5245 ;
  assign n5255 = n5254 ^ n5237 ;
  assign n5288 = n5287 ^ n5255 ;
  assign n5293 = n137 & n2341 ;
  assign n5294 = n5293 ^ n137 ;
  assign n5295 = n5294 ^ n137 ;
  assign n5289 = n138 & n2320 ;
  assign n5290 = n5289 ^ n138 ;
  assign n5291 = n5290 ^ n2320 ;
  assign n5292 = n5291 ^ n138 ;
  assign n5296 = n5295 ^ n5292 ;
  assign n5340 = n1259 & n2175 ;
  assign n5341 = n5340 ^ n1259 ;
  assign n5342 = n5341 ^ n1259 ;
  assign n5343 = ~n5296 & n5342 ;
  assign n5344 = n5343 ^ n5342 ;
  assign n5345 = n5344 ^ n5342 ;
  assign n5319 = n1003 & n1151 ;
  assign n5320 = n5319 ^ n402 ;
  assign n5321 = n2254 & n5320 ;
  assign n5322 = n5321 ^ n5320 ;
  assign n5312 = n136 & n2265 ;
  assign n5313 = n5312 ^ n136 ;
  assign n5316 = n2284 & n5313 ;
  assign n5317 = n5316 ^ n136 ;
  assign n5314 = n2269 & n5313 ;
  assign n5315 = n5314 ^ n5313 ;
  assign n5318 = n5317 ^ n5315 ;
  assign n5323 = n5322 ^ n5318 ;
  assign n5308 = n903 & n1553 ;
  assign n5309 = n2254 & n5308 ;
  assign n5310 = n5309 ^ n5308 ;
  assign n5311 = n5310 ^ n402 ;
  assign n5324 = n5323 ^ n5311 ;
  assign n5331 = x134 & n5324 ;
  assign n5332 = n5331 ^ x134 ;
  assign n5333 = n138 & n2366 ;
  assign n5334 = n5333 ^ n138 ;
  assign n5335 = n5334 ^ n2366 ;
  assign n5336 = n5335 ^ n138 ;
  assign n5337 = n5332 & ~n5336 ;
  assign n5338 = n5337 ^ n5332 ;
  assign n5325 = n2222 & n4076 ;
  assign n5326 = n5325 ^ n4076 ;
  assign n5327 = n5326 ^ n4076 ;
  assign n5328 = n5327 ^ x134 ;
  assign n5329 = n5324 & n5328 ;
  assign n5330 = n5329 ^ n5328 ;
  assign n5339 = n5338 ^ n5330 ;
  assign n5346 = n5345 ^ n5339 ;
  assign n5301 = n2199 & n2748 ;
  assign n5302 = n5301 ^ n2748 ;
  assign n5303 = n5302 ^ n2748 ;
  assign n5304 = ~n5296 & n5303 ;
  assign n5305 = n5304 ^ n5303 ;
  assign n5306 = n5305 ^ n5303 ;
  assign n5297 = x134 & ~n5296 ;
  assign n5298 = n5297 ^ x134 ;
  assign n5299 = n5298 ^ x134 ;
  assign n5300 = n5299 ^ n5296 ;
  assign n5307 = n5306 ^ n5300 ;
  assign n5347 = n5346 ^ n5307 ;
  assign n5378 = n138 & n2428 ;
  assign n5379 = n5378 ^ n138 ;
  assign n5380 = n5379 ^ n2428 ;
  assign n5381 = n5380 ^ n138 ;
  assign n5370 = n137 & n2403 ;
  assign n5371 = n5370 ^ n137 ;
  assign n5375 = n2411 & n5371 ;
  assign n5376 = n5375 ^ n137 ;
  assign n5372 = n2407 & n5371 ;
  assign n5373 = n5372 ^ n5371 ;
  assign n5374 = n5373 ^ n5371 ;
  assign n5377 = n5376 ^ n5374 ;
  assign n5382 = n5381 ^ n5377 ;
  assign n5384 = n136 & n2446 ;
  assign n5385 = n5384 ^ n136 ;
  assign n5388 = n2452 & n5385 ;
  assign n5389 = n5388 ^ n136 ;
  assign n5386 = n2449 & n5385 ;
  assign n5387 = n5386 ^ n5385 ;
  assign n5390 = n5389 ^ n5387 ;
  assign n5383 = n402 & n2467 ;
  assign n5391 = n5390 ^ n5383 ;
  assign n5392 = ~n5382 & n5391 ;
  assign n5393 = n5392 ^ n5391 ;
  assign n5394 = n5393 ^ n5382 ;
  assign n5395 = n5394 ^ n5391 ;
  assign n5396 = x134 & ~n5395 ;
  assign n5397 = n5396 ^ x134 ;
  assign n5398 = n5397 ^ x134 ;
  assign n5351 = n402 & ~n2376 ;
  assign n5352 = ~n2393 & n5351 ;
  assign n5350 = n136 & n2390 ;
  assign n5353 = n5352 ^ n5350 ;
  assign n5348 = n1553 & n2378 ;
  assign n5349 = n5348 ^ n402 ;
  assign n5354 = n5353 ^ n5349 ;
  assign n5356 = n137 & n2486 ;
  assign n5357 = n5356 ^ n137 ;
  assign n5360 = n2493 & n5357 ;
  assign n5361 = n5360 ^ n137 ;
  assign n5358 = n2489 & n5357 ;
  assign n5359 = n5358 ^ n5357 ;
  assign n5362 = n5361 ^ n5359 ;
  assign n5355 = ~n138 & ~n2482 ;
  assign n5363 = n5362 ^ n5355 ;
  assign n5364 = x134 & n5363 ;
  assign n5365 = n5364 ^ x134 ;
  assign n5366 = n5365 ^ n5363 ;
  assign n5367 = n5354 & n5366 ;
  assign n5368 = n5367 ^ n5354 ;
  assign n5369 = n5368 ^ n5366 ;
  assign n5399 = n5398 ^ n5369 ;
  assign n5456 = ~n2662 & n4441 ;
  assign n5457 = n5456 ^ n4441 ;
  assign n5427 = n402 & ~n1768 ;
  assign n5428 = ~n2600 & n5427 ;
  assign n5425 = n1768 & n3002 ;
  assign n5426 = ~n2600 & n5425 ;
  assign n5429 = n5428 ^ n5426 ;
  assign n5418 = n136 & n2626 ;
  assign n5419 = n5418 ^ n136 ;
  assign n5422 = n2633 & n5419 ;
  assign n5420 = n2629 & n5419 ;
  assign n5421 = n5420 ^ n5419 ;
  assign n5423 = n5422 ^ n5421 ;
  assign n5424 = n5423 ^ n136 ;
  assign n5430 = n5429 ^ n5424 ;
  assign n5415 = n1553 & n1649 ;
  assign n5416 = ~n2600 & n5415 ;
  assign n5417 = n5416 ^ n402 ;
  assign n5431 = n5430 ^ n5417 ;
  assign n5447 = n1175 & n2708 ;
  assign n5448 = n5447 ^ n1175 ;
  assign n5449 = n5448 ^ n1175 ;
  assign n5450 = n5449 ^ x134 ;
  assign n5451 = n5431 & n5450 ;
  assign n5452 = n5451 ^ n5450 ;
  assign n5453 = n5452 ^ n2570 ;
  assign n5454 = n5453 ^ n137 ;
  assign n5432 = n5431 ^ n137 ;
  assign n5433 = n5432 ^ x134 ;
  assign n5434 = n1669 ^ n137 ;
  assign n5435 = n5434 ^ x134 ;
  assign n5436 = n2585 & n5435 ;
  assign n5437 = n5436 ^ n5435 ;
  assign n5438 = n5437 ^ n5435 ;
  assign n5439 = n5438 ^ n1669 ;
  assign n5440 = n5439 ^ n5431 ;
  assign n5441 = n5440 ^ n2585 ;
  assign n5442 = n5433 & n5441 ;
  assign n5443 = n5442 ^ n5433 ;
  assign n5444 = n5443 ^ n5433 ;
  assign n5445 = n5444 ^ n5438 ;
  assign n5446 = n5445 ^ n1669 ;
  assign n5455 = n5454 ^ n5446 ;
  assign n5458 = n5457 ^ n5455 ;
  assign n5410 = x132 & ~x133 ;
  assign n5411 = ~x134 & n5410 ;
  assign n5412 = ~n2685 & n5411 ;
  assign n5413 = n5412 ^ n5411 ;
  assign n5403 = n136 & n2547 ;
  assign n5404 = n5403 ^ n136 ;
  assign n5405 = n5404 ^ n136 ;
  assign n5400 = n402 & n2523 ;
  assign n5401 = n5400 ^ n402 ;
  assign n5402 = n5401 ^ n402 ;
  assign n5406 = n5405 ^ n5402 ;
  assign n5407 = x134 & n5406 ;
  assign n5408 = n5407 ^ x134 ;
  assign n5409 = n5408 ^ n5406 ;
  assign n5414 = n5413 ^ n5409 ;
  assign n5459 = n5458 ^ n5414 ;
  assign n5464 = n137 & n2758 ;
  assign n5465 = n5464 ^ n137 ;
  assign n5466 = n5465 ^ n137 ;
  assign n5460 = n138 & n2844 ;
  assign n5461 = n5460 ^ n138 ;
  assign n5462 = n5461 ^ n2844 ;
  assign n5463 = n5462 ^ n138 ;
  assign n5467 = n5466 ^ n5463 ;
  assign n5468 = x134 & ~n5467 ;
  assign n5469 = n5468 ^ x134 ;
  assign n5470 = n5469 ^ x134 ;
  assign n5511 = n136 & ~n2802 ;
  assign n5512 = n5511 ^ n136 ;
  assign n5513 = n5470 & n5512 ;
  assign n5514 = n5513 ^ n5470 ;
  assign n5495 = n490 & n589 ;
  assign n5496 = n2765 & n5495 ;
  assign n5497 = n5496 ^ n5495 ;
  assign n5481 = n138 & n139 ;
  assign n5482 = n5481 ^ n139 ;
  assign n5483 = n575 & n5482 ;
  assign n5484 = n5483 ^ n138 ;
  assign n5478 = n138 & n155 ;
  assign n5479 = n5478 ^ n155 ;
  assign n5480 = n561 & n5479 ;
  assign n5485 = n5484 ^ n5480 ;
  assign n5491 = n2780 & ~n5485 ;
  assign n5492 = n5491 ^ n5485 ;
  assign n5486 = n171 & n5485 ;
  assign n5487 = n5486 ^ n171 ;
  assign n5488 = n5487 ^ n5485 ;
  assign n5489 = n541 & n5488 ;
  assign n5490 = n5489 ^ n541 ;
  assign n5493 = n5492 ^ n5490 ;
  assign n5494 = n5493 ^ x133 ;
  assign n5498 = n5497 ^ n5494 ;
  assign n5474 = n602 & n5187 ;
  assign n5475 = n5474 ^ n137 ;
  assign n5476 = n2765 & n5475 ;
  assign n5477 = n5476 ^ n5475 ;
  assign n5499 = n5498 ^ n5477 ;
  assign n5500 = x134 & n5499 ;
  assign n5501 = n5500 ^ x134 ;
  assign n5502 = n5501 ^ n5499 ;
  assign n5507 = n136 & n2743 ;
  assign n5508 = n5502 & n5507 ;
  assign n5509 = n5508 ^ n5507 ;
  assign n5503 = n402 & n2726 ;
  assign n5504 = n5502 & n5503 ;
  assign n5505 = n5504 ^ n5503 ;
  assign n5506 = n5505 ^ n5502 ;
  assign n5510 = n5509 ^ n5506 ;
  assign n5515 = n5514 ^ n5510 ;
  assign n5471 = n402 & ~n2818 ;
  assign n5472 = n5471 ^ n402 ;
  assign n5473 = n5470 & n5472 ;
  assign n5516 = n5515 ^ n5473 ;
  assign n5570 = n903 & n1003 ;
  assign n5571 = n5570 ^ n402 ;
  assign n5572 = n2941 & n5571 ;
  assign n5573 = n5572 ^ n5571 ;
  assign n5565 = n136 & ~n2962 ;
  assign n5567 = n2969 & n5565 ;
  assign n5568 = n5567 ^ n136 ;
  assign n5566 = ~n2966 & n5565 ;
  assign n5569 = n5568 ^ n5566 ;
  assign n5574 = n5573 ^ n5569 ;
  assign n5561 = n921 & n1094 ;
  assign n5562 = n2941 & n5561 ;
  assign n5563 = n5562 ^ n5561 ;
  assign n5564 = n5563 ^ n402 ;
  assign n5575 = n5574 ^ n5564 ;
  assign n5579 = n1175 & n3038 ;
  assign n5580 = n5579 ^ n1175 ;
  assign n5581 = n5580 ^ n1175 ;
  assign n5582 = n5581 ^ x134 ;
  assign n5583 = n5575 & n5582 ;
  assign n5584 = n5583 ^ n5582 ;
  assign n5576 = n2915 & n4076 ;
  assign n5577 = n5575 & n5576 ;
  assign n5578 = n5577 ^ n5576 ;
  assign n5585 = n5584 ^ n5578 ;
  assign n5537 = n490 & n969 ;
  assign n5538 = n5537 ^ n137 ;
  assign n5539 = n2985 & n5538 ;
  assign n5540 = n5539 ^ n5538 ;
  assign n5526 = n138 & n2999 ;
  assign n5527 = n5526 ^ n2999 ;
  assign n5528 = n5527 ^ n138 ;
  assign n5529 = n5528 ^ n1827 ;
  assign n5521 = n138 & n1015 ;
  assign n5522 = n5521 ^ n1015 ;
  assign n5523 = n5522 ^ n138 ;
  assign n5524 = n2992 & n5523 ;
  assign n5525 = n5524 ^ n2992 ;
  assign n5530 = n5529 ^ n5525 ;
  assign n5531 = n5530 ^ n138 ;
  assign n5534 = n3009 & n5531 ;
  assign n5532 = n3006 & n5531 ;
  assign n5533 = n5532 ^ n5531 ;
  assign n5535 = n5534 ^ n5533 ;
  assign n5536 = n5535 ^ n138 ;
  assign n5541 = n5540 ^ n5536 ;
  assign n5517 = n505 & n985 ;
  assign n5518 = n2985 & n5517 ;
  assign n5519 = n5518 ^ n5517 ;
  assign n5520 = n5519 ^ n137 ;
  assign n5542 = n5541 ^ n5520 ;
  assign n5543 = x134 & n5542 ;
  assign n5544 = n5543 ^ x134 ;
  assign n5545 = n5544 ^ x134 ;
  assign n5546 = n5545 ^ n5542 ;
  assign n5554 = n136 & n2896 ;
  assign n5555 = n5554 ^ n136 ;
  assign n5556 = n5555 ^ n136 ;
  assign n5557 = n5546 & n5556 ;
  assign n5558 = n5557 ^ n5556 ;
  assign n5559 = n5558 ^ n5556 ;
  assign n5547 = n402 & n2872 ;
  assign n5548 = n5547 ^ n402 ;
  assign n5549 = n5548 ^ n402 ;
  assign n5550 = n5546 & n5549 ;
  assign n5551 = n5550 ^ n5549 ;
  assign n5552 = n5551 ^ n5549 ;
  assign n5553 = n5552 ^ n5546 ;
  assign n5560 = n5559 ^ n5553 ;
  assign n5586 = n5585 ^ n5560 ;
  assign n5609 = n4639 & n4640 ;
  assign n5610 = n5609 ^ n4639 ;
  assign n5611 = n5610 ^ n4640 ;
  assign n5605 = n3748 & n4643 ;
  assign n5606 = n3119 & n5605 ;
  assign n5607 = n5606 ^ n5605 ;
  assign n5612 = n5611 ^ n5607 ;
  assign n5613 = n5612 ^ n5605 ;
  assign n5614 = n5613 ^ n4640 ;
  assign n5615 = n5611 ^ n5605 ;
  assign n5616 = n5615 ^ n3762 ;
  assign n5617 = n5614 & n5616 ;
  assign n5618 = n5617 ^ n5614 ;
  assign n5619 = n5618 ^ n5616 ;
  assign n5620 = n5619 ^ n5616 ;
  assign n5621 = n5620 ^ n5611 ;
  assign n5608 = n5607 ^ n5605 ;
  assign n5622 = n5621 ^ n5608 ;
  assign n5623 = n5622 ^ n4640 ;
  assign n5604 = n402 & n3132 ;
  assign n5624 = n5623 ^ n5604 ;
  assign n5601 = n1442 & n3014 ;
  assign n5602 = ~n3119 & n5601 ;
  assign n5603 = n5602 ^ n136 ;
  assign n5625 = n5624 ^ n5603 ;
  assign n5633 = n170 & ~n1371 ;
  assign n5634 = n5633 ^ n170 ;
  assign n5635 = n137 & n3053 ;
  assign n5636 = n5635 ^ n137 ;
  assign n5637 = n5634 & n5636 ;
  assign n5638 = n5637 ^ n5636 ;
  assign n5629 = n138 & n3067 ;
  assign n5630 = n5629 ^ n138 ;
  assign n5631 = n5630 ^ n3067 ;
  assign n5632 = n5631 ^ n138 ;
  assign n5639 = n5638 ^ n5632 ;
  assign n5626 = n505 & n1360 ;
  assign n5627 = ~n3053 & n5626 ;
  assign n5628 = n5627 ^ n137 ;
  assign n5640 = n5639 ^ n5628 ;
  assign n5641 = ~n5625 & ~n5640 ;
  assign n5642 = n5641 ^ n5625 ;
  assign n5643 = n5642 ^ n5640 ;
  assign n5644 = n5643 ^ n5625 ;
  assign n5645 = n5644 ^ n5640 ;
  assign n5646 = x134 & n5645 ;
  assign n5588 = n137 & ~n3157 ;
  assign n5590 = n3163 & n5588 ;
  assign n5591 = n5590 ^ n137 ;
  assign n5589 = ~n3160 & n5588 ;
  assign n5592 = n5591 ^ n5589 ;
  assign n5587 = ~n138 & ~n3149 ;
  assign n5593 = n5592 ^ n5587 ;
  assign n5598 = n1259 & n3086 ;
  assign n5599 = ~n5593 & n5598 ;
  assign n5594 = n2748 & n3102 ;
  assign n5595 = n5594 ^ x134 ;
  assign n5596 = n5593 & ~n5595 ;
  assign n5597 = n5596 ^ n5595 ;
  assign n5600 = n5599 ^ n5597 ;
  assign n5647 = n5646 ^ n5600 ;
  assign n5652 = n137 & n3334 ;
  assign n5648 = n138 & n3317 ;
  assign n5649 = n5648 ^ n138 ;
  assign n5650 = n5649 ^ n3317 ;
  assign n5651 = n5650 ^ n138 ;
  assign n5653 = n5652 ^ n5651 ;
  assign n5704 = n1259 & n3188 ;
  assign n5705 = ~n5653 & n5704 ;
  assign n5706 = n5705 ^ n5704 ;
  assign n5707 = n5706 ^ n5704 ;
  assign n5677 = n402 & ~n1649 ;
  assign n5678 = ~n3263 & n5677 ;
  assign n5675 = n1649 & n3002 ;
  assign n5676 = ~n3263 & n5675 ;
  assign n5679 = n5678 ^ n5676 ;
  assign n5668 = n136 & n3280 ;
  assign n5669 = n5668 ^ n136 ;
  assign n5672 = n3296 & n5669 ;
  assign n5673 = n5672 ^ n136 ;
  assign n5670 = n3284 & n5669 ;
  assign n5671 = n5670 ^ n5669 ;
  assign n5674 = n5673 ^ n5671 ;
  assign n5680 = n5679 ^ n5674 ;
  assign n5665 = n1553 & n1659 ;
  assign n5666 = ~n3263 & n5665 ;
  assign n5667 = n5666 ^ n402 ;
  assign n5681 = n5680 ^ n5667 ;
  assign n5695 = n1175 & n3359 ;
  assign n5696 = n5695 ^ n1175 ;
  assign n5697 = n5696 ^ n1175 ;
  assign n5698 = n5697 ^ x134 ;
  assign n5699 = n5681 & n5698 ;
  assign n5700 = n5699 ^ n5698 ;
  assign n5701 = n5700 ^ n3235 ;
  assign n5702 = n5701 ^ n137 ;
  assign n5682 = n5681 ^ n137 ;
  assign n5683 = n5682 ^ x134 ;
  assign n5684 = n3249 & n5435 ;
  assign n5685 = n5684 ^ n5435 ;
  assign n5686 = n5685 ^ n5435 ;
  assign n5687 = n5686 ^ n1669 ;
  assign n5688 = n5687 ^ n5681 ;
  assign n5689 = n5688 ^ n3249 ;
  assign n5690 = n5683 & n5689 ;
  assign n5691 = n5690 ^ n5683 ;
  assign n5692 = n5691 ^ n5683 ;
  assign n5693 = n5692 ^ n5686 ;
  assign n5694 = n5693 ^ n1669 ;
  assign n5703 = n5702 ^ n5694 ;
  assign n5708 = n5707 ^ n5703 ;
  assign n5658 = n2748 & n3212 ;
  assign n5659 = n5658 ^ n2748 ;
  assign n5660 = n5659 ^ n2748 ;
  assign n5661 = ~n5653 & n5660 ;
  assign n5662 = n5661 ^ n5660 ;
  assign n5663 = n5662 ^ n5660 ;
  assign n5654 = x134 & ~n5653 ;
  assign n5655 = n5654 ^ x134 ;
  assign n5656 = n5655 ^ x134 ;
  assign n5657 = n5656 ^ n5653 ;
  assign n5664 = n5663 ^ n5657 ;
  assign n5709 = n5708 ^ n5664 ;
  assign n5714 = n137 & n3408 ;
  assign n5715 = n5714 ^ n137 ;
  assign n5716 = n5715 ^ n137 ;
  assign n5710 = n138 & n3508 ;
  assign n5711 = n5710 ^ n138 ;
  assign n5712 = n5711 ^ n3508 ;
  assign n5713 = n5712 ^ n138 ;
  assign n5717 = n5716 ^ n5713 ;
  assign n5718 = x134 & ~n5717 ;
  assign n5719 = n5718 ^ x134 ;
  assign n5720 = n5719 ^ x134 ;
  assign n5753 = n136 & ~n3479 ;
  assign n5754 = n5753 ^ n136 ;
  assign n5755 = n5720 & n5754 ;
  assign n5756 = n5755 ^ n5720 ;
  assign n5727 = n561 & n5482 ;
  assign n5728 = n5727 ^ n138 ;
  assign n5726 = n520 & n5479 ;
  assign n5729 = n5728 ^ n5726 ;
  assign n5731 = n170 & n5729 ;
  assign n5732 = n5731 ^ n170 ;
  assign n5733 = n541 & n5732 ;
  assign n5734 = n5733 ^ n5732 ;
  assign n5735 = n5734 ^ n5732 ;
  assign n5736 = n5735 ^ n5729 ;
  assign n5730 = n3429 & ~n5729 ;
  assign n5737 = n5736 ^ n5730 ;
  assign n5738 = n5737 ^ x133 ;
  assign n5724 = n137 & n3422 ;
  assign n5725 = n5724 ^ n137 ;
  assign n5739 = n5738 ^ n5725 ;
  assign n5745 = n136 & n3394 ;
  assign n5746 = n5739 & n5745 ;
  assign n5747 = n5746 ^ n5745 ;
  assign n5748 = n5747 ^ n5739 ;
  assign n5740 = n402 & n3378 ;
  assign n5741 = n5740 ^ n402 ;
  assign n5742 = n5741 ^ n402 ;
  assign n5743 = n5739 & n5742 ;
  assign n5744 = n5743 ^ n5742 ;
  assign n5749 = n5748 ^ n5744 ;
  assign n5750 = x134 & n5749 ;
  assign n5751 = n5750 ^ x134 ;
  assign n5752 = n5751 ^ n5749 ;
  assign n5757 = n5756 ^ n5752 ;
  assign n5721 = n402 & ~n3454 ;
  assign n5722 = n5721 ^ n402 ;
  assign n5723 = n5720 & n5722 ;
  assign n5758 = n5757 ^ n5723 ;
  assign n5804 = n1180 & ~n3611 ;
  assign n5805 = n5804 ^ n1180 ;
  assign n5797 = n137 & n3558 ;
  assign n5798 = n5797 ^ n137 ;
  assign n5799 = n5798 ^ n137 ;
  assign n5793 = n138 & n3655 ;
  assign n5794 = n5793 ^ n138 ;
  assign n5795 = n5794 ^ n3655 ;
  assign n5796 = n5795 ^ n138 ;
  assign n5800 = n5799 ^ n5796 ;
  assign n5801 = x134 & ~n5800 ;
  assign n5802 = n5801 ^ x134 ;
  assign n5803 = n5802 ^ x134 ;
  assign n5806 = n5805 ^ n5803 ;
  assign n5769 = n490 & n985 ;
  assign n5770 = n5769 ^ n137 ;
  assign n5771 = n3573 & n5770 ;
  assign n5772 = n5771 ^ n5770 ;
  assign n5766 = n138 & n3591 ;
  assign n5767 = n5766 ^ n3591 ;
  assign n5768 = n5767 ^ n138 ;
  assign n5773 = n5772 ^ n5768 ;
  assign n5762 = n505 & n1002 ;
  assign n5763 = n3573 & n5762 ;
  assign n5764 = n5763 ^ n5762 ;
  assign n5765 = n5764 ^ n137 ;
  assign n5774 = n5773 ^ n5765 ;
  assign n5775 = x134 & n5774 ;
  assign n5776 = n5775 ^ x134 ;
  assign n5777 = n5776 ^ x134 ;
  assign n5778 = n5777 ^ n5774 ;
  assign n5786 = n402 & n3526 ;
  assign n5787 = n5786 ^ n402 ;
  assign n5788 = n5787 ^ n402 ;
  assign n5789 = n5778 & n5788 ;
  assign n5790 = n5789 ^ n5788 ;
  assign n5791 = n5790 ^ n5788 ;
  assign n5779 = n136 & n3540 ;
  assign n5780 = n5779 ^ n136 ;
  assign n5781 = n5780 ^ n136 ;
  assign n5782 = n5778 & n5781 ;
  assign n5783 = n5782 ^ n5781 ;
  assign n5784 = n5783 ^ n5781 ;
  assign n5785 = n5784 ^ n5778 ;
  assign n5792 = n5791 ^ n5785 ;
  assign n5807 = n5806 ^ n5792 ;
  assign n5759 = x134 & n2347 ;
  assign n5760 = ~n3633 & n5759 ;
  assign n5761 = n5760 ^ n5759 ;
  assign n5808 = n5807 ^ n5761 ;
  assign n5838 = n136 & ~n4910 ;
  assign n5839 = ~n3720 & n5838 ;
  assign n5837 = n402 & n3742 ;
  assign n5840 = n5839 ^ n5837 ;
  assign n5833 = n1492 & n3014 ;
  assign n5834 = n3720 & n5833 ;
  assign n5835 = n5834 ^ n5833 ;
  assign n5836 = n5835 ^ n136 ;
  assign n5841 = n5840 ^ n5836 ;
  assign n5846 = n137 & n3710 ;
  assign n5842 = n138 & n3694 ;
  assign n5843 = n5842 ^ n138 ;
  assign n5844 = n5843 ^ n3694 ;
  assign n5845 = n5844 ^ n138 ;
  assign n5847 = n5846 ^ n5845 ;
  assign n5848 = x134 & ~n5847 ;
  assign n5849 = n5848 ^ x134 ;
  assign n5850 = n5849 ^ x134 ;
  assign n5851 = n5841 & n5850 ;
  assign n5852 = n5851 ^ n5850 ;
  assign n5814 = n137 & ~n4882 ;
  assign n5815 = ~n3778 & n5814 ;
  assign n5813 = ~n138 & n3821 ;
  assign n5816 = n5815 ^ n5813 ;
  assign n5809 = n505 & n1501 ;
  assign n5810 = n3778 & n5809 ;
  assign n5811 = n5810 ^ n5809 ;
  assign n5812 = n5811 ^ n137 ;
  assign n5817 = n5816 ^ n5812 ;
  assign n5825 = n402 & n3672 ;
  assign n5818 = n136 & n3676 ;
  assign n5819 = n5818 ^ n136 ;
  assign n5822 = n3680 & n5819 ;
  assign n5823 = n5822 ^ n136 ;
  assign n5820 = n3678 & n5819 ;
  assign n5821 = n5820 ^ n5819 ;
  assign n5824 = n5823 ^ n5821 ;
  assign n5826 = n5825 ^ n5824 ;
  assign n5827 = x134 & n5826 ;
  assign n5828 = n5827 ^ x134 ;
  assign n5829 = n5828 ^ n5826 ;
  assign n5830 = n5817 & n5829 ;
  assign n5831 = n5830 ^ n5817 ;
  assign n5832 = n5831 ^ n5829 ;
  assign n5853 = n5852 ^ n5832 ;
  assign n5911 = n1180 & ~n3937 ;
  assign n5912 = n5911 ^ n1180 ;
  assign n5904 = n137 & n3877 ;
  assign n5905 = n5904 ^ n137 ;
  assign n5906 = n5905 ^ n137 ;
  assign n5900 = n138 & n3983 ;
  assign n5901 = n5900 ^ n138 ;
  assign n5902 = n5901 ^ n3983 ;
  assign n5903 = n5902 ^ n138 ;
  assign n5907 = n5906 ^ n5903 ;
  assign n5908 = x134 & ~n5907 ;
  assign n5909 = n5908 ^ x134 ;
  assign n5910 = n5909 ^ x134 ;
  assign n5913 = n5912 ^ n5910 ;
  assign n5876 = n490 & n1942 ;
  assign n5877 = n5876 ^ n137 ;
  assign n5878 = n3894 & n5877 ;
  assign n5879 = n5878 ^ n5877 ;
  assign n5865 = n138 & n3910 ;
  assign n5866 = n5865 ^ n3910 ;
  assign n5867 = n5866 ^ n138 ;
  assign n5868 = n5867 ^ n1827 ;
  assign n5860 = n138 & n1809 ;
  assign n5861 = n5860 ^ n1809 ;
  assign n5862 = n5861 ^ n138 ;
  assign n5863 = n3901 & n5862 ;
  assign n5864 = n5863 ^ n3901 ;
  assign n5869 = n5868 ^ n5864 ;
  assign n5870 = n5869 ^ n138 ;
  assign n5873 = n3917 & n5870 ;
  assign n5871 = n3914 & n5870 ;
  assign n5872 = n5871 ^ n5870 ;
  assign n5874 = n5873 ^ n5872 ;
  assign n5875 = n5874 ^ n138 ;
  assign n5880 = n5879 ^ n5875 ;
  assign n5856 = n505 & n1923 ;
  assign n5857 = n3894 & n5856 ;
  assign n5858 = n5857 ^ n5856 ;
  assign n5859 = n5858 ^ n137 ;
  assign n5881 = n5880 ^ n5859 ;
  assign n5882 = x134 & n5881 ;
  assign n5883 = n5882 ^ x134 ;
  assign n5884 = n5883 ^ x134 ;
  assign n5885 = n5884 ^ n5881 ;
  assign n5893 = n402 & n3845 ;
  assign n5894 = n5893 ^ n402 ;
  assign n5895 = n5894 ^ n402 ;
  assign n5896 = n5885 & n5895 ;
  assign n5897 = n5896 ^ n5895 ;
  assign n5898 = n5897 ^ n5895 ;
  assign n5886 = n136 & n3859 ;
  assign n5887 = n5886 ^ n136 ;
  assign n5888 = n5887 ^ n136 ;
  assign n5889 = n5885 & n5888 ;
  assign n5890 = n5889 ^ n5888 ;
  assign n5891 = n5890 ^ n5888 ;
  assign n5892 = n5891 ^ n5885 ;
  assign n5899 = n5898 ^ n5892 ;
  assign n5914 = n5913 ^ n5899 ;
  assign n5854 = ~n3957 & n5759 ;
  assign n5855 = n5854 ^ n5759 ;
  assign n5915 = n5914 ^ n5855 ;
  assign n6003 = ~n308 & n1949 ;
  assign n6004 = ~n336 & n6003 ;
  assign n5921 = n138 & n272 ;
  assign n5922 = n5921 ^ n272 ;
  assign n5923 = n5922 ^ n138 ;
  assign n5924 = n5923 ^ n138 ;
  assign n5918 = n136 & n474 ;
  assign n5919 = n5918 ^ n136 ;
  assign n5920 = n5919 ^ n136 ;
  assign n5925 = n5924 ^ n5920 ;
  assign n5990 = x134 & n308 ;
  assign n5999 = n5990 ^ x134 ;
  assign n6000 = n336 & n5999 ;
  assign n6001 = n6000 ^ n5999 ;
  assign n6002 = n5925 & n6001 ;
  assign n6005 = n6004 ^ n6002 ;
  assign n5997 = n308 & n1949 ;
  assign n5998 = n5925 & n5997 ;
  assign n6006 = n6005 ^ n5998 ;
  assign n5991 = n5990 ^ n308 ;
  assign n5992 = n336 & n5991 ;
  assign n5993 = n5925 & n5992 ;
  assign n5994 = n5993 ^ n5992 ;
  assign n5984 = ~x134 & ~n402 ;
  assign n5988 = n308 & n5984 ;
  assign n5989 = n336 & n5988 ;
  assign n5995 = n5994 ^ n5989 ;
  assign n5985 = ~n308 & n5984 ;
  assign n5986 = n5925 & n5985 ;
  assign n5987 = n5986 ^ n5985 ;
  assign n5996 = n5995 ^ n5987 ;
  assign n6007 = n6006 ^ n5996 ;
  assign n5960 = n5925 ^ n402 ;
  assign n5962 = n5925 ^ n336 ;
  assign n5963 = n5960 & n5962 ;
  assign n5964 = n5963 ^ n5960 ;
  assign n5965 = n5964 ^ n5960 ;
  assign n5966 = n5965 ^ n5962 ;
  assign n5967 = n5966 ^ n336 ;
  assign n5968 = n5967 ^ n308 ;
  assign n6008 = n6007 ^ n5968 ;
  assign n5982 = n5967 ^ n402 ;
  assign n5958 = n5925 ^ x134 ;
  assign n5983 = n5982 ^ n5958 ;
  assign n6009 = n6008 ^ n5983 ;
  assign n6021 = n6009 ^ n5966 ;
  assign n5977 = n336 & n405 ;
  assign n5978 = n5925 & n5977 ;
  assign n5974 = ~n336 & n1259 ;
  assign n5975 = n5925 & n5974 ;
  assign n5976 = n5975 ^ n5974 ;
  assign n5979 = n5978 ^ n5976 ;
  assign n5972 = ~x134 & ~n308 ;
  assign n5970 = n308 & n5925 ;
  assign n5971 = n5970 ^ n5925 ;
  assign n5973 = n5972 ^ n5971 ;
  assign n5980 = n5979 ^ n5973 ;
  assign n5961 = n5960 ^ x134 ;
  assign n5969 = n5968 ^ n5961 ;
  assign n5981 = n5980 ^ n5969 ;
  assign n6010 = n6009 ^ n5981 ;
  assign n6011 = n6010 ^ n5967 ;
  assign n6012 = n6011 ^ n5961 ;
  assign n6013 = n6009 ^ n308 ;
  assign n6014 = n6013 ^ x134 ;
  assign n6015 = n6012 & n6014 ;
  assign n6016 = n6015 ^ n6012 ;
  assign n6017 = n6016 ^ n6014 ;
  assign n6018 = n6017 ^ n6012 ;
  assign n6019 = n6018 ^ n6014 ;
  assign n6020 = n6019 ^ n5981 ;
  assign n6022 = n6021 ^ n6020 ;
  assign n5957 = n402 ^ n336 ;
  assign n5959 = n5958 ^ n5957 ;
  assign n6023 = n6022 ^ n5959 ;
  assign n5942 = n137 & n607 ;
  assign n5943 = n5942 ^ n137 ;
  assign n5930 = n503 & n1451 ;
  assign n5931 = n5930 ^ n503 ;
  assign n5932 = n5931 ^ n138 ;
  assign n5929 = n489 & n2256 ;
  assign n5933 = n5932 ^ n5929 ;
  assign n5935 = n155 & n5933 ;
  assign n5936 = n5935 ^ n155 ;
  assign n5937 = n541 & n5936 ;
  assign n5938 = n5937 ^ n5936 ;
  assign n5939 = n5938 ^ n5936 ;
  assign n5940 = n5939 ^ n5933 ;
  assign n5934 = n521 & ~n5933 ;
  assign n5941 = n5940 ^ n5934 ;
  assign n5944 = n5943 ^ n5941 ;
  assign n5945 = n5944 ^ x133 ;
  assign n5949 = n136 & n202 ;
  assign n5950 = n5945 & n5949 ;
  assign n5951 = n5950 ^ n5949 ;
  assign n5952 = n5951 ^ n5945 ;
  assign n5946 = n402 & n672 ;
  assign n5947 = n5945 & n5946 ;
  assign n5948 = n5947 ^ n5946 ;
  assign n5953 = n5952 ^ n5948 ;
  assign n5954 = x134 & n5953 ;
  assign n5955 = n5954 ^ x134 ;
  assign n5956 = n5955 ^ n5953 ;
  assign n6024 = n6023 ^ n5956 ;
  assign n5916 = n137 & n399 ;
  assign n5917 = n5916 ^ n137 ;
  assign n5926 = x134 & n5925 ;
  assign n5927 = n5926 ^ x134 ;
  assign n5928 = n5917 & n5927 ;
  assign n6025 = n6024 ^ n5928 ;
  assign n6071 = ~n1174 & n1180 ;
  assign n6072 = n6071 ^ n1180 ;
  assign n6064 = n137 & n1331 ;
  assign n6065 = n6064 ^ n137 ;
  assign n6066 = n6065 ^ n137 ;
  assign n6060 = n138 & n845 ;
  assign n6061 = n6060 ^ n138 ;
  assign n6062 = n6061 ^ n845 ;
  assign n6063 = n6062 ^ n138 ;
  assign n6067 = n6066 ^ n6063 ;
  assign n6068 = x134 & ~n6067 ;
  assign n6069 = n6068 ^ x134 ;
  assign n6070 = n6069 ^ x134 ;
  assign n6073 = n6072 ^ n6070 ;
  assign n6038 = n490 & n1002 ;
  assign n6039 = n6038 ^ n137 ;
  assign n6040 = n987 & n6039 ;
  assign n6041 = n6040 ^ n6039 ;
  assign n6032 = n138 & n1075 ;
  assign n6033 = n6032 ^ n138 ;
  assign n6034 = n6033 ^ n1075 ;
  assign n6035 = n1041 & ~n6034 ;
  assign n6036 = n6035 ^ n6034 ;
  assign n6037 = n6036 ^ n138 ;
  assign n6042 = n6041 ^ n6037 ;
  assign n6028 = n505 & n1093 ;
  assign n6029 = n987 & n6028 ;
  assign n6030 = n6029 ^ n6028 ;
  assign n6031 = n6030 ^ n137 ;
  assign n6043 = n6042 ^ n6031 ;
  assign n6044 = x134 & ~n6043 ;
  assign n6045 = n6044 ^ x134 ;
  assign n6046 = n6045 ^ x134 ;
  assign n6047 = n6046 ^ n6043 ;
  assign n6055 = n402 & n1254 ;
  assign n6056 = ~n6047 & n6055 ;
  assign n6057 = n6056 ^ n6055 ;
  assign n6058 = n6057 ^ n6055 ;
  assign n6048 = n136 & n763 ;
  assign n6049 = n6048 ^ n136 ;
  assign n6050 = n6049 ^ n136 ;
  assign n6051 = ~n6047 & n6050 ;
  assign n6052 = n6051 ^ n6050 ;
  assign n6053 = n6052 ^ n6050 ;
  assign n6054 = n6053 ^ n6047 ;
  assign n6059 = n6058 ^ n6054 ;
  assign n6074 = n6073 ^ n6059 ;
  assign n6026 = ~n930 & n5759 ;
  assign n6027 = n6026 ^ n5759 ;
  assign n6075 = n6074 ^ n6027 ;
  assign n6119 = n1492 & n2785 ;
  assign n6120 = n6119 ^ n136 ;
  assign n6121 = n1446 & n6120 ;
  assign n6122 = n6121 ^ n6120 ;
  assign n6114 = n402 & ~n1345 ;
  assign n6116 = n1355 & n6114 ;
  assign n6117 = n6116 ^ n402 ;
  assign n6115 = ~n1350 & n6114 ;
  assign n6118 = n6117 ^ n6115 ;
  assign n6123 = n6122 ^ n6118 ;
  assign n6110 = n1448 & n3014 ;
  assign n6111 = n1446 & n6110 ;
  assign n6112 = n6111 ^ n6110 ;
  assign n6113 = n6112 ^ n136 ;
  assign n6124 = n6123 ^ n6113 ;
  assign n6129 = n137 & n1375 ;
  assign n6125 = n138 & n1423 ;
  assign n6126 = n6125 ^ n138 ;
  assign n6127 = n6126 ^ n1423 ;
  assign n6128 = n6127 ^ n138 ;
  assign n6130 = n6129 ^ n6128 ;
  assign n6131 = x134 & ~n6130 ;
  assign n6132 = n6131 ^ x134 ;
  assign n6133 = n6132 ^ x134 ;
  assign n6134 = n6124 & n6133 ;
  assign n6135 = n6134 ^ n6133 ;
  assign n6085 = n490 & n1501 ;
  assign n6086 = n6085 ^ n137 ;
  assign n6087 = n1514 & n6086 ;
  assign n6088 = n6087 ^ n6086 ;
  assign n6080 = ~n138 & ~n1538 ;
  assign n6082 = n1548 & n6080 ;
  assign n6083 = n6082 ^ n138 ;
  assign n6081 = ~n1543 & n6080 ;
  assign n6084 = n6083 ^ n6081 ;
  assign n6089 = n6088 ^ n6084 ;
  assign n6076 = n505 & n1556 ;
  assign n6077 = n1514 & n6076 ;
  assign n6078 = n6077 ^ n6076 ;
  assign n6079 = n6078 ^ n137 ;
  assign n6090 = n6089 ^ n6079 ;
  assign n6099 = n402 & n1484 ;
  assign n6100 = n6099 ^ n402 ;
  assign n6101 = n6100 ^ n402 ;
  assign n6091 = n136 & n1387 ;
  assign n6092 = n6091 ^ n136 ;
  assign n6096 = n1401 & n6092 ;
  assign n6097 = n6096 ^ n136 ;
  assign n6093 = n1394 & n6092 ;
  assign n6094 = n6093 ^ n6092 ;
  assign n6095 = n6094 ^ n6092 ;
  assign n6098 = n6097 ^ n6095 ;
  assign n6102 = n6101 ^ n6098 ;
  assign n6103 = x134 & n6102 ;
  assign n6104 = n6103 ^ x134 ;
  assign n6105 = n6104 ^ n6102 ;
  assign n6106 = n6090 & n6105 ;
  assign n6107 = n6106 ^ n6105 ;
  assign n6108 = n6107 ^ n6090 ;
  assign n6109 = n6108 ^ n6105 ;
  assign n6136 = n6135 ^ n6109 ;
  assign n6184 = n1180 & ~n4206 ;
  assign n6185 = n6184 ^ n1180 ;
  assign n6178 = n137 & n1999 ;
  assign n6179 = n6178 ^ n137 ;
  assign n6180 = n6179 ^ n137 ;
  assign n6175 = n402 & n1664 ;
  assign n6176 = n6175 ^ n402 ;
  assign n6177 = n6176 ^ n402 ;
  assign n6181 = n6180 ^ n6177 ;
  assign n6182 = x134 & n6181 ;
  assign n6183 = n6182 ^ x134 ;
  assign n6186 = n6185 ^ n6183 ;
  assign n6153 = n490 & n1923 ;
  assign n6154 = n6153 ^ n137 ;
  assign n6155 = n1946 & n6154 ;
  assign n6156 = n6155 ^ n6154 ;
  assign n6143 = n138 & n1799 ;
  assign n6144 = n6143 ^ n138 ;
  assign n6145 = n6144 ^ n1799 ;
  assign n6146 = n6145 ^ n138 ;
  assign n6147 = n6146 ^ n138 ;
  assign n6150 = n4184 & ~n6147 ;
  assign n6148 = n4180 & ~n6147 ;
  assign n6149 = n6148 ^ n6147 ;
  assign n6151 = n6150 ^ n6149 ;
  assign n6152 = n6151 ^ n138 ;
  assign n6157 = n6156 ^ n6152 ;
  assign n6139 = n505 & n1914 ;
  assign n6140 = n1946 & n6139 ;
  assign n6141 = n6140 ^ n6139 ;
  assign n6142 = n6141 ^ n137 ;
  assign n6158 = n6157 ^ n6142 ;
  assign n6159 = x134 & ~n6158 ;
  assign n6160 = n6159 ^ x134 ;
  assign n6161 = n6160 ^ x134 ;
  assign n6162 = n6161 ^ n6158 ;
  assign n6170 = n402 & n1898 ;
  assign n6171 = ~n6162 & n6170 ;
  assign n6172 = n6171 ^ n6170 ;
  assign n6173 = n6172 ^ n6170 ;
  assign n6163 = n136 & n1620 ;
  assign n6164 = n6163 ^ n136 ;
  assign n6165 = n6164 ^ n136 ;
  assign n6166 = ~n6162 & n6165 ;
  assign n6167 = n6166 ^ n6165 ;
  assign n6168 = n6167 ^ n6165 ;
  assign n6169 = n6168 ^ n6162 ;
  assign n6174 = n6173 ^ n6169 ;
  assign n6187 = n6186 ^ n6174 ;
  assign n6137 = n1175 & ~n1715 ;
  assign n6138 = n6137 ^ n1175 ;
  assign n6188 = n6187 ^ n6138 ;
  assign n6206 = n456 & n1451 ;
  assign n6207 = n6206 ^ n456 ;
  assign n6208 = n6207 ^ n138 ;
  assign n6205 = n503 & n2256 ;
  assign n6209 = n6208 ^ n6205 ;
  assign n6213 = n2080 & ~n6209 ;
  assign n6214 = n6213 ^ n6209 ;
  assign n6210 = n139 & n6209 ;
  assign n6211 = n6210 ^ n139 ;
  assign n6212 = n541 & n6211 ;
  assign n6215 = n6214 ^ n6212 ;
  assign n6216 = n6215 ^ x132 ;
  assign n6202 = n136 & n2017 ;
  assign n6203 = n6202 ^ n136 ;
  assign n6204 = n6203 ^ x133 ;
  assign n6217 = n6216 ^ n6204 ;
  assign n6285 = n6217 ^ x134 ;
  assign n6290 = n2133 ^ n402 ;
  assign n6291 = n2133 & n6290 ;
  assign n6286 = n137 & n2109 ;
  assign n6287 = n6286 ^ n137 ;
  assign n6288 = n6287 ^ n137 ;
  assign n6289 = n6288 ^ n2133 ;
  assign n6292 = n6291 ^ n6289 ;
  assign n6293 = n6292 ^ x134 ;
  assign n6294 = n6292 & n6293 ;
  assign n6295 = n6294 ^ n6292 ;
  assign n6296 = n6295 ^ n6293 ;
  assign n6297 = n6296 ^ x134 ;
  assign n6298 = n6285 & n6297 ;
  assign n6299 = n6298 ^ n6285 ;
  assign n6300 = n6299 ^ n6297 ;
  assign n6301 = n6300 ^ n6297 ;
  assign n6302 = n6301 ^ n6296 ;
  assign n6303 = n6302 ^ n6217 ;
  assign n6264 = n1949 & ~n2052 ;
  assign n6265 = ~n2056 & n6264 ;
  assign n6195 = n136 & n2093 ;
  assign n6196 = n6195 ^ n136 ;
  assign n6197 = n6196 ^ n136 ;
  assign n6191 = n138 & n2039 ;
  assign n6192 = n6191 ^ n2039 ;
  assign n6193 = n6192 ^ n138 ;
  assign n6194 = n6193 ^ n138 ;
  assign n6198 = n6197 ^ n6194 ;
  assign n6251 = x134 & n2052 ;
  assign n6260 = n6251 ^ x134 ;
  assign n6261 = n2056 & n6260 ;
  assign n6262 = n6261 ^ n6260 ;
  assign n6263 = n6198 & n6262 ;
  assign n6266 = n6265 ^ n6263 ;
  assign n6258 = n1949 & n2052 ;
  assign n6259 = n6198 & n6258 ;
  assign n6267 = n6266 ^ n6259 ;
  assign n6252 = n6251 ^ n2052 ;
  assign n6253 = n2056 & n6252 ;
  assign n6254 = n6198 & n6253 ;
  assign n6255 = n6254 ^ n6253 ;
  assign n6249 = n2052 & n5984 ;
  assign n6250 = n2056 & n6249 ;
  assign n6256 = n6255 ^ n6250 ;
  assign n6246 = ~n2052 & n5984 ;
  assign n6247 = n6198 & n6246 ;
  assign n6248 = n6247 ^ n6246 ;
  assign n6257 = n6256 ^ n6248 ;
  assign n6268 = n6267 ^ n6257 ;
  assign n6222 = n6198 ^ n402 ;
  assign n6224 = n6198 ^ n2056 ;
  assign n6225 = n6222 & n6224 ;
  assign n6226 = n6225 ^ n6222 ;
  assign n6227 = n6226 ^ n6222 ;
  assign n6228 = n6227 ^ n6224 ;
  assign n6229 = n6228 ^ n2056 ;
  assign n6230 = n6229 ^ n2052 ;
  assign n6269 = n6268 ^ n6230 ;
  assign n6244 = n6229 ^ n402 ;
  assign n6220 = n6198 ^ x134 ;
  assign n6245 = n6244 ^ n6220 ;
  assign n6270 = n6269 ^ n6245 ;
  assign n6282 = n6270 ^ n6228 ;
  assign n6239 = n405 & n2056 ;
  assign n6240 = n6198 & n6239 ;
  assign n6236 = n1259 & ~n2056 ;
  assign n6237 = n6198 & n6236 ;
  assign n6238 = n6237 ^ n6236 ;
  assign n6241 = n6240 ^ n6238 ;
  assign n6234 = ~x134 & ~n2052 ;
  assign n6232 = n2052 & n6198 ;
  assign n6233 = n6232 ^ n6198 ;
  assign n6235 = n6234 ^ n6233 ;
  assign n6242 = n6241 ^ n6235 ;
  assign n6223 = n6222 ^ x134 ;
  assign n6231 = n6230 ^ n6223 ;
  assign n6243 = n6242 ^ n6231 ;
  assign n6271 = n6270 ^ n6243 ;
  assign n6272 = n6271 ^ n6229 ;
  assign n6273 = n6272 ^ n6223 ;
  assign n6274 = n6270 ^ n2052 ;
  assign n6275 = n6274 ^ x134 ;
  assign n6276 = n6273 & n6275 ;
  assign n6277 = n6276 ^ n6273 ;
  assign n6278 = n6277 ^ n6275 ;
  assign n6279 = n6278 ^ n6273 ;
  assign n6280 = n6279 ^ n6275 ;
  assign n6281 = n6280 ^ n6243 ;
  assign n6283 = n6282 ^ n6281 ;
  assign n6219 = n2056 ^ n402 ;
  assign n6221 = n6220 ^ n6219 ;
  assign n6284 = n6283 ^ n6221 ;
  assign n6304 = n6303 ^ n6284 ;
  assign n6218 = ~x134 & ~n6217 ;
  assign n6305 = n6304 ^ n6218 ;
  assign n6189 = n137 & n2070 ;
  assign n6190 = n6189 ^ n137 ;
  assign n6199 = x134 & n6198 ;
  assign n6200 = n6199 ^ x134 ;
  assign n6201 = n6190 & n6200 ;
  assign n6306 = n6305 ^ n6201 ;
  assign n6356 = ~n2222 & n5759 ;
  assign n6357 = n6356 ^ n5759 ;
  assign n6349 = n136 & n4325 ;
  assign n6350 = n6349 ^ n136 ;
  assign n6351 = n6350 ^ n136 ;
  assign n6345 = n138 & n2199 ;
  assign n6346 = n6345 ^ n138 ;
  assign n6347 = n6346 ^ n2199 ;
  assign n6348 = n6347 ^ n138 ;
  assign n6352 = n6351 ^ n6348 ;
  assign n6353 = x134 & ~n6352 ;
  assign n6354 = n6353 ^ x134 ;
  assign n6355 = n6354 ^ x134 ;
  assign n6358 = n6357 ^ n6355 ;
  assign n6324 = n698 & n2785 ;
  assign n6325 = n6324 ^ n136 ;
  assign n6326 = n2170 & n6325 ;
  assign n6327 = n6326 ^ n6325 ;
  assign n6314 = n138 & n2265 ;
  assign n6315 = n6314 ^ n2265 ;
  assign n6316 = n6315 ^ n138 ;
  assign n6320 = n2284 & n6316 ;
  assign n6321 = n6320 ^ n2284 ;
  assign n6322 = n6321 ^ n138 ;
  assign n6317 = n2269 & n6316 ;
  assign n6318 = n6317 ^ n2269 ;
  assign n6319 = n6318 ^ n6316 ;
  assign n6323 = n6322 ^ n6319 ;
  assign n6328 = n6327 ^ n6323 ;
  assign n6310 = n1229 & n3014 ;
  assign n6311 = n2170 & n6310 ;
  assign n6312 = n6311 ^ n6310 ;
  assign n6313 = n6312 ^ n136 ;
  assign n6329 = n6328 ^ n6313 ;
  assign n6330 = x134 & n6329 ;
  assign n6331 = n6330 ^ x134 ;
  assign n6332 = n6331 ^ n6329 ;
  assign n6339 = n402 & n2341 ;
  assign n6340 = n6339 ^ n402 ;
  assign n6341 = n6340 ^ n402 ;
  assign n6342 = n6332 & n6341 ;
  assign n6343 = n6342 ^ n6341 ;
  assign n6333 = n137 & n2320 ;
  assign n6334 = n6333 ^ n137 ;
  assign n6335 = n6334 ^ n137 ;
  assign n6336 = n6332 & n6335 ;
  assign n6337 = n6336 ^ n6335 ;
  assign n6338 = n6337 ^ n6332 ;
  assign n6344 = n6343 ^ n6338 ;
  assign n6359 = n6358 ^ n6344 ;
  assign n6307 = x134 & n5410 ;
  assign n6308 = ~n2366 & n6307 ;
  assign n6309 = n6308 ^ n6307 ;
  assign n6360 = n6359 ^ n6309 ;
  assign n6393 = n137 & n2428 ;
  assign n6388 = n402 & ~n2403 ;
  assign n6390 = n2411 & n6388 ;
  assign n6391 = n6390 ^ n402 ;
  assign n6389 = n2407 & n6388 ;
  assign n6392 = n6391 ^ n6389 ;
  assign n6394 = n6393 ^ n6392 ;
  assign n6399 = n1180 & n2467 ;
  assign n6400 = ~n6394 & n6399 ;
  assign n6395 = n1175 & n2390 ;
  assign n6396 = n6395 ^ x134 ;
  assign n6397 = n6394 & n6396 ;
  assign n6398 = n6397 ^ n6396 ;
  assign n6401 = n6400 ^ n6398 ;
  assign n6368 = n136 & ~n2376 ;
  assign n6369 = ~n2393 & n6368 ;
  assign n6363 = ~n138 & ~n2446 ;
  assign n6365 = n2452 & n6363 ;
  assign n6366 = n6365 ^ n138 ;
  assign n6364 = ~n2449 & n6363 ;
  assign n6367 = n6366 ^ n6364 ;
  assign n6370 = n6369 ^ n6367 ;
  assign n6361 = n2378 & n3014 ;
  assign n6362 = n6361 ^ n136 ;
  assign n6371 = n6370 ^ n6362 ;
  assign n6373 = n402 & n2486 ;
  assign n6374 = n6373 ^ n402 ;
  assign n6377 = n2493 & n6374 ;
  assign n6378 = n6377 ^ n402 ;
  assign n6375 = n2489 & n6374 ;
  assign n6376 = n6375 ^ n6374 ;
  assign n6379 = n6378 ^ n6376 ;
  assign n6372 = n137 & ~n2482 ;
  assign n6380 = n6379 ^ n6372 ;
  assign n6381 = x134 & n6380 ;
  assign n6382 = n6381 ^ x134 ;
  assign n6383 = n6382 ^ n6380 ;
  assign n6384 = n6371 & n6383 ;
  assign n6385 = n6384 ^ n6383 ;
  assign n6386 = n6385 ^ n6371 ;
  assign n6387 = n6386 ^ n6383 ;
  assign n6402 = n6401 ^ n6387 ;
  assign n6444 = n137 & n2708 ;
  assign n6445 = n6444 ^ n137 ;
  assign n6446 = n6445 ^ n137 ;
  assign n6440 = n138 & n2547 ;
  assign n6441 = n6440 ^ n138 ;
  assign n6442 = n6441 ^ n2547 ;
  assign n6443 = n6442 ^ n138 ;
  assign n6447 = n6446 ^ n6443 ;
  assign n6451 = n171 & n1649 ;
  assign n6452 = n6451 ^ n171 ;
  assign n6453 = n6452 ^ n1649 ;
  assign n6454 = n6453 ^ n171 ;
  assign n6448 = n170 & n1768 ;
  assign n6449 = n6448 ^ n170 ;
  assign n6450 = n6449 ^ n170 ;
  assign n6455 = n6454 ^ n6450 ;
  assign n6456 = n2600 & n6455 ;
  assign n6457 = n6456 ^ n2600 ;
  assign n6458 = n6457 ^ n6455 ;
  assign n6465 = x134 & n6458 ;
  assign n6466 = n6465 ^ x134 ;
  assign n6467 = ~n6447 & n6466 ;
  assign n6468 = n6467 ^ n6466 ;
  assign n6469 = n6468 ^ n6466 ;
  assign n6459 = n1899 & n6458 ;
  assign n6460 = n6459 ^ n1899 ;
  assign n6461 = n6460 ^ n1899 ;
  assign n6462 = ~n6447 & n6461 ;
  assign n6463 = n6462 ^ n6461 ;
  assign n6464 = n6463 ^ n6461 ;
  assign n6470 = n6469 ^ n6464 ;
  assign n6419 = n1003 & n1865 ;
  assign n6420 = n6419 ^ n402 ;
  assign n6421 = n2682 & n6420 ;
  assign n6422 = n6421 ^ n6420 ;
  assign n6409 = n138 & n2626 ;
  assign n6410 = n6409 ^ n2626 ;
  assign n6411 = n6410 ^ n138 ;
  assign n6415 = n2633 & n6411 ;
  assign n6416 = n6415 ^ n2633 ;
  assign n6412 = n2629 & n6411 ;
  assign n6413 = n6412 ^ n2629 ;
  assign n6414 = n6413 ^ n6411 ;
  assign n6417 = n6416 ^ n6414 ;
  assign n6418 = n6417 ^ n138 ;
  assign n6423 = n6422 ^ n6418 ;
  assign n6405 = n1553 & n1932 ;
  assign n6406 = n2682 & n6405 ;
  assign n6407 = n6406 ^ n6405 ;
  assign n6408 = n6407 ^ n402 ;
  assign n6424 = n6423 ^ n6408 ;
  assign n6425 = x134 & n6424 ;
  assign n6426 = n6425 ^ x134 ;
  assign n6427 = n6426 ^ n6424 ;
  assign n6434 = n137 & n2662 ;
  assign n6435 = n6434 ^ n137 ;
  assign n6436 = n6435 ^ n137 ;
  assign n6437 = n6427 & n6436 ;
  assign n6438 = n6437 ^ n6436 ;
  assign n6428 = n136 & n2523 ;
  assign n6429 = n6428 ^ n136 ;
  assign n6430 = n6429 ^ n136 ;
  assign n6431 = n6427 & n6430 ;
  assign n6432 = n6431 ^ n6430 ;
  assign n6433 = n6432 ^ n6427 ;
  assign n6439 = n6438 ^ n6433 ;
  assign n6471 = n6470 ^ n6439 ;
  assign n6403 = ~n2570 & n5759 ;
  assign n6404 = n6403 ^ n5759 ;
  assign n6472 = n6471 ^ n6404 ;
  assign n6477 = n137 & n2844 ;
  assign n6478 = n6477 ^ n137 ;
  assign n6479 = n6478 ^ n137 ;
  assign n6473 = n138 & n2743 ;
  assign n6474 = n6473 ^ n2743 ;
  assign n6475 = n6474 ^ n138 ;
  assign n6476 = n6475 ^ n138 ;
  assign n6480 = n6479 ^ n6476 ;
  assign n6522 = x134 & n6480 ;
  assign n6523 = n6522 ^ x134 ;
  assign n6524 = n136 & ~n2818 ;
  assign n6525 = n6524 ^ n136 ;
  assign n6526 = n6523 & n6525 ;
  assign n6527 = n6526 ^ n6523 ;
  assign n6496 = n136 & n2726 ;
  assign n6497 = n6496 ^ n136 ;
  assign n6485 = n575 & n1849 ;
  assign n6486 = n6485 ^ n137 ;
  assign n6484 = n561 & n1813 ;
  assign n6487 = n6486 ^ n6484 ;
  assign n6493 = n2780 & n6487 ;
  assign n6494 = n6493 ^ n6487 ;
  assign n6488 = n171 & n6487 ;
  assign n6489 = n6488 ^ n6487 ;
  assign n6490 = n541 & n6489 ;
  assign n6491 = n6490 ^ n6489 ;
  assign n6492 = n6491 ^ n6489 ;
  assign n6495 = n6494 ^ n6492 ;
  assign n6498 = n6497 ^ n6495 ;
  assign n6499 = n6498 ^ x132 ;
  assign n6510 = n138 & n2802 ;
  assign n6511 = n6510 ^ n138 ;
  assign n6512 = n6511 ^ n2802 ;
  assign n6513 = n6499 & ~n6512 ;
  assign n6514 = n6513 ^ n6512 ;
  assign n6507 = n138 & n6499 ;
  assign n6508 = n6507 ^ n6499 ;
  assign n6509 = n6508 ^ n138 ;
  assign n6515 = n6514 ^ n6509 ;
  assign n6516 = n6515 ^ n6499 ;
  assign n6502 = n402 & n4484 ;
  assign n6503 = n6502 ^ n402 ;
  assign n6504 = n6499 & n6503 ;
  assign n6505 = n6504 ^ n6503 ;
  assign n6500 = n402 & n6499 ;
  assign n6501 = n6500 ^ n402 ;
  assign n6506 = n6505 ^ n6501 ;
  assign n6517 = n6516 ^ n6506 ;
  assign n6518 = x134 & ~n6517 ;
  assign n6519 = n6518 ^ x134 ;
  assign n6520 = n6519 ^ x134 ;
  assign n6521 = n6520 ^ n6517 ;
  assign n6528 = n6527 ^ n6521 ;
  assign n6481 = n1949 & n2758 ;
  assign n6482 = n6480 & n6481 ;
  assign n6483 = n6482 ^ n6481 ;
  assign n6529 = n6528 ^ n6483 ;
  assign n6585 = n137 & n3038 ;
  assign n6586 = n6585 ^ n137 ;
  assign n6587 = n6586 ^ n137 ;
  assign n6581 = n138 & n2896 ;
  assign n6582 = n6581 ^ n138 ;
  assign n6583 = n6582 ^ n2896 ;
  assign n6584 = n6583 ^ n138 ;
  assign n6588 = n6587 ^ n6584 ;
  assign n6593 = n170 & n903 ;
  assign n6594 = n6593 ^ n170 ;
  assign n6595 = n6594 ^ n170 ;
  assign n6589 = n171 & n921 ;
  assign n6590 = n6589 ^ n171 ;
  assign n6591 = n6590 ^ n921 ;
  assign n6592 = n6591 ^ n171 ;
  assign n6596 = n6595 ^ n6592 ;
  assign n6597 = n2941 & n6596 ;
  assign n6598 = n6597 ^ n2941 ;
  assign n6599 = n6598 ^ n6596 ;
  assign n6606 = x134 & n6599 ;
  assign n6607 = n6606 ^ x134 ;
  assign n6608 = ~n6588 & n6607 ;
  assign n6609 = n6608 ^ n6607 ;
  assign n6610 = n6609 ^ n6607 ;
  assign n6600 = n1899 & n6599 ;
  assign n6601 = n6600 ^ n1899 ;
  assign n6602 = n6601 ^ n1899 ;
  assign n6603 = ~n6588 & n6602 ;
  assign n6604 = n6603 ^ n6602 ;
  assign n6605 = n6604 ^ n6602 ;
  assign n6611 = n6610 ^ n6605 ;
  assign n6546 = n969 & n1003 ;
  assign n6547 = n6546 ^ n402 ;
  assign n6548 = n2985 & n6547 ;
  assign n6549 = n6548 ^ n6547 ;
  assign n6536 = n138 & n2962 ;
  assign n6537 = n6536 ^ n2962 ;
  assign n6538 = n6537 ^ n138 ;
  assign n6542 = n2969 & n6538 ;
  assign n6543 = n6542 ^ n2969 ;
  assign n6544 = n6543 ^ n138 ;
  assign n6539 = n2966 & n6538 ;
  assign n6540 = n6539 ^ n2966 ;
  assign n6541 = n6540 ^ n6538 ;
  assign n6545 = n6544 ^ n6541 ;
  assign n6550 = n6549 ^ n6545 ;
  assign n6532 = n985 & n1553 ;
  assign n6533 = n2985 & n6532 ;
  assign n6534 = n6533 ^ n6532 ;
  assign n6535 = n6534 ^ n402 ;
  assign n6551 = n6550 ^ n6535 ;
  assign n6569 = n1229 & n2785 ;
  assign n6570 = n6569 ^ n136 ;
  assign n6571 = n2867 & n6570 ;
  assign n6572 = n6571 ^ n6570 ;
  assign n6559 = n137 & n2999 ;
  assign n6560 = n6559 ^ n137 ;
  assign n6561 = n6560 ^ n4416 ;
  assign n6556 = n137 & n1015 ;
  assign n6557 = n6556 ^ n137 ;
  assign n6558 = n2992 & n6557 ;
  assign n6562 = n6561 ^ n6558 ;
  assign n6563 = n6562 ^ n137 ;
  assign n6566 = n3009 & n6563 ;
  assign n6564 = n3006 & n6563 ;
  assign n6565 = n6564 ^ n6563 ;
  assign n6567 = n6566 ^ n6565 ;
  assign n6568 = n6567 ^ n137 ;
  assign n6573 = n6572 ^ n6568 ;
  assign n6552 = n1247 & n3014 ;
  assign n6553 = n2867 & n6552 ;
  assign n6554 = n6553 ^ n6552 ;
  assign n6555 = n6554 ^ n136 ;
  assign n6574 = n6573 ^ n6555 ;
  assign n6575 = n6551 & n6574 ;
  assign n6576 = n6575 ^ n6551 ;
  assign n6577 = n6576 ^ n6574 ;
  assign n6578 = x134 & n6577 ;
  assign n6579 = n6578 ^ x134 ;
  assign n6580 = n6579 ^ n6577 ;
  assign n6612 = n6611 ^ n6580 ;
  assign n6530 = ~n2915 & n5759 ;
  assign n6531 = n6530 ^ n5759 ;
  assign n6613 = n6612 ^ n6531 ;
  assign n6639 = n137 & n3067 ;
  assign n6638 = ~n138 & n3102 ;
  assign n6640 = n6639 ^ n6638 ;
  assign n6646 = n1003 & n1371 ;
  assign n6647 = n6646 ^ n402 ;
  assign n6648 = n3053 & n6647 ;
  assign n6649 = n6648 ^ n6647 ;
  assign n6645 = n136 & n3132 ;
  assign n6650 = n6649 ^ n6645 ;
  assign n6641 = n1360 & n1553 ;
  assign n6642 = n3053 & n6641 ;
  assign n6643 = n6642 ^ n6641 ;
  assign n6644 = n6643 ^ n402 ;
  assign n6651 = n6650 ^ n6644 ;
  assign n6652 = x134 & ~n6651 ;
  assign n6653 = ~n6640 & n6652 ;
  assign n6618 = ~n138 & ~n3134 ;
  assign n6619 = ~n3119 & n6618 ;
  assign n6617 = n136 & n3086 ;
  assign n6620 = n6619 ^ n6617 ;
  assign n6614 = ~n138 & n3120 ;
  assign n6615 = ~n3119 & n6614 ;
  assign n6616 = n6615 ^ n138 ;
  assign n6621 = n6620 ^ n6616 ;
  assign n6623 = n402 & n3157 ;
  assign n6624 = n6623 ^ n402 ;
  assign n6627 = n3163 & n6624 ;
  assign n6628 = n6627 ^ n402 ;
  assign n6625 = n3160 & n6624 ;
  assign n6626 = n6625 ^ n6624 ;
  assign n6629 = n6628 ^ n6626 ;
  assign n6622 = n137 & ~n3149 ;
  assign n6630 = n6629 ^ n6622 ;
  assign n6631 = x134 & n6630 ;
  assign n6632 = n6631 ^ x134 ;
  assign n6633 = n6632 ^ n6630 ;
  assign n6634 = n6621 & n6633 ;
  assign n6635 = n6634 ^ n6633 ;
  assign n6636 = n6635 ^ n6621 ;
  assign n6637 = n6636 ^ n6633 ;
  assign n6654 = n6653 ^ n6637 ;
  assign n6703 = n137 & n3359 ;
  assign n6704 = n6703 ^ n137 ;
  assign n6705 = n6704 ^ n137 ;
  assign n6699 = n138 & n3212 ;
  assign n6700 = n6699 ^ n138 ;
  assign n6701 = n6700 ^ n3212 ;
  assign n6702 = n6701 ^ n138 ;
  assign n6706 = n6705 ^ n6702 ;
  assign n6710 = n171 & n1659 ;
  assign n6711 = n6710 ^ n1659 ;
  assign n6707 = n170 & n1649 ;
  assign n6708 = n6707 ^ n170 ;
  assign n6709 = n6708 ^ n170 ;
  assign n6712 = n6711 ^ n6709 ;
  assign n6713 = n3263 & n6712 ;
  assign n6714 = n6713 ^ n3263 ;
  assign n6715 = n6714 ^ n6712 ;
  assign n6720 = x134 & n6715 ;
  assign n6721 = n6720 ^ x134 ;
  assign n6722 = ~n6706 & n6721 ;
  assign n6723 = n6722 ^ n6721 ;
  assign n6724 = n6723 ^ n6721 ;
  assign n6716 = n1899 & n6715 ;
  assign n6717 = ~n6706 & n6716 ;
  assign n6718 = n6717 ^ n6716 ;
  assign n6719 = n6718 ^ n6716 ;
  assign n6725 = n6724 ^ n6719 ;
  assign n6677 = n1883 & n2785 ;
  assign n6678 = n6677 ^ n136 ;
  assign n6679 = n3185 & n6678 ;
  assign n6680 = n6679 ^ n6678 ;
  assign n6666 = n138 & n3279 ;
  assign n6667 = n6666 ^ n3279 ;
  assign n6668 = n6667 ^ n138 ;
  assign n6669 = n6668 ^ n1827 ;
  assign n6661 = n138 & n1744 ;
  assign n6662 = n6661 ^ n1744 ;
  assign n6663 = n6662 ^ n138 ;
  assign n6664 = n3271 & n6663 ;
  assign n6665 = n6664 ^ n3271 ;
  assign n6670 = n6669 ^ n6665 ;
  assign n6671 = n6670 ^ n138 ;
  assign n6674 = n3296 & n6671 ;
  assign n6675 = n6674 ^ n138 ;
  assign n6672 = n3284 & n6671 ;
  assign n6673 = n6672 ^ n6671 ;
  assign n6676 = n6675 ^ n6673 ;
  assign n6681 = n6680 ^ n6676 ;
  assign n6657 = n1893 & n3014 ;
  assign n6658 = n3185 & n6657 ;
  assign n6659 = n6658 ^ n6657 ;
  assign n6660 = n6659 ^ n136 ;
  assign n6682 = n6681 ^ n6660 ;
  assign n6683 = x134 & n6682 ;
  assign n6684 = n6683 ^ x134 ;
  assign n6685 = n6684 ^ x134 ;
  assign n6686 = n6685 ^ n6682 ;
  assign n6694 = n402 & n3334 ;
  assign n6695 = n6686 & n6694 ;
  assign n6696 = n6695 ^ n6694 ;
  assign n6697 = n6696 ^ n6694 ;
  assign n6687 = n137 & n3317 ;
  assign n6688 = n6687 ^ n137 ;
  assign n6689 = n6688 ^ n137 ;
  assign n6690 = n6686 & n6689 ;
  assign n6691 = n6690 ^ n6689 ;
  assign n6692 = n6691 ^ n6689 ;
  assign n6693 = n6692 ^ n6686 ;
  assign n6698 = n6697 ^ n6693 ;
  assign n6726 = n6725 ^ n6698 ;
  assign n6655 = ~n3235 & n5759 ;
  assign n6656 = n6655 ^ n5759 ;
  assign n6727 = n6726 ^ n6656 ;
  assign n6732 = n137 & n3508 ;
  assign n6733 = n6732 ^ n137 ;
  assign n6734 = n6733 ^ n137 ;
  assign n6728 = n138 & n3394 ;
  assign n6729 = n6728 ^ n3394 ;
  assign n6730 = n6729 ^ n138 ;
  assign n6731 = n6730 ^ n138 ;
  assign n6735 = n6734 ^ n6731 ;
  assign n6766 = x134 & n6735 ;
  assign n6767 = n6766 ^ x134 ;
  assign n6768 = n136 & ~n3454 ;
  assign n6769 = n6768 ^ n136 ;
  assign n6770 = n6767 & n6769 ;
  assign n6771 = n6770 ^ n6767 ;
  assign n6743 = n561 & n1849 ;
  assign n6744 = n6743 ^ n137 ;
  assign n6742 = n520 & n1813 ;
  assign n6745 = n6744 ^ n6742 ;
  assign n6747 = n170 & n6745 ;
  assign n6748 = n541 & n6747 ;
  assign n6749 = n6748 ^ n6745 ;
  assign n6746 = n3429 & n6745 ;
  assign n6750 = n6749 ^ n6746 ;
  assign n6751 = n6750 ^ x132 ;
  assign n6739 = n402 & n3422 ;
  assign n6740 = n6739 ^ n402 ;
  assign n6741 = n6740 ^ x133 ;
  assign n6752 = n6751 ^ n6741 ;
  assign n6753 = x134 & n6752 ;
  assign n6754 = n6753 ^ x134 ;
  assign n6755 = n6754 ^ n6752 ;
  assign n6762 = n136 & n3378 ;
  assign n6763 = n6755 & n6762 ;
  assign n6764 = n6763 ^ n6762 ;
  assign n6756 = ~n138 & ~n3479 ;
  assign n6757 = n6756 ^ n138 ;
  assign n6758 = n6755 & n6757 ;
  assign n6759 = n6758 ^ n6755 ;
  assign n6760 = n6759 ^ n6757 ;
  assign n6761 = n6760 ^ n6755 ;
  assign n6765 = n6764 ^ n6761 ;
  assign n6772 = n6771 ^ n6765 ;
  assign n6736 = n1949 & n3408 ;
  assign n6737 = n6735 & n6736 ;
  assign n6738 = n6737 ^ n6736 ;
  assign n6773 = n6772 ^ n6738 ;
  assign n6778 = n137 & n3655 ;
  assign n6779 = n6778 ^ n137 ;
  assign n6780 = n6779 ^ n137 ;
  assign n6774 = n138 & n3540 ;
  assign n6775 = n6774 ^ n138 ;
  assign n6776 = n6775 ^ n3540 ;
  assign n6777 = n6776 ^ n138 ;
  assign n6781 = n6780 ^ n6777 ;
  assign n6815 = n1180 & n3633 ;
  assign n6816 = n6815 ^ n1180 ;
  assign n6817 = n6816 ^ n1180 ;
  assign n6818 = ~n6781 & n6817 ;
  assign n6819 = n6818 ^ n6817 ;
  assign n6820 = n6819 ^ n6817 ;
  assign n6794 = n985 & n1003 ;
  assign n6795 = n6794 ^ n402 ;
  assign n6796 = n3573 & n6795 ;
  assign n6797 = n6796 ^ n6795 ;
  assign n6793 = n137 & ~n3591 ;
  assign n6798 = n6797 ^ n6793 ;
  assign n6789 = n1002 & n1094 ;
  assign n6790 = n3573 & n6789 ;
  assign n6791 = n6790 ^ n6789 ;
  assign n6792 = n6791 ^ n402 ;
  assign n6799 = n6798 ^ n6792 ;
  assign n6809 = n2748 & n3526 ;
  assign n6810 = n6809 ^ n2748 ;
  assign n6811 = n6810 ^ n2748 ;
  assign n6812 = n6799 & n6811 ;
  assign n6813 = n6812 ^ n6811 ;
  assign n6803 = n3611 & n4441 ;
  assign n6804 = n6803 ^ n4441 ;
  assign n6805 = n6804 ^ n4441 ;
  assign n6806 = n6799 & n6805 ;
  assign n6807 = n6806 ^ n6805 ;
  assign n6800 = x134 & n6799 ;
  assign n6801 = n6800 ^ x134 ;
  assign n6802 = n6801 ^ n6799 ;
  assign n6808 = n6807 ^ n6802 ;
  assign n6814 = n6813 ^ n6808 ;
  assign n6821 = n6820 ^ n6814 ;
  assign n6786 = x134 & ~n6781 ;
  assign n6787 = n6786 ^ x134 ;
  assign n6788 = n6787 ^ x134 ;
  assign n6822 = n6821 ^ n6788 ;
  assign n6782 = n1949 & n3558 ;
  assign n6783 = ~n6781 & n6782 ;
  assign n6784 = n6783 ^ n6782 ;
  assign n6785 = n6784 ^ n6782 ;
  assign n6823 = n6822 ^ n6785 ;
  assign n6884 = n137 & n3694 ;
  assign n6879 = ~n138 & ~n3676 ;
  assign n6881 = n3680 & n6879 ;
  assign n6882 = n6881 ^ n138 ;
  assign n6880 = ~n3678 & n6879 ;
  assign n6883 = n6882 ^ n6880 ;
  assign n6885 = n6884 ^ n6883 ;
  assign n6890 = n1949 & n3710 ;
  assign n6891 = n6885 & n6890 ;
  assign n6886 = n1180 & n3742 ;
  assign n6887 = n6886 ^ x134 ;
  assign n6888 = ~n6885 & n6887 ;
  assign n6889 = n6888 ^ n6887 ;
  assign n6892 = n6891 ^ n6889 ;
  assign n6830 = n3748 & ~n3750 ;
  assign n6831 = ~n3720 & n6830 ;
  assign n6839 = n6831 ^ n6830 ;
  assign n6829 = n3756 & ~n3757 ;
  assign n6832 = n6831 ^ n6829 ;
  assign n6833 = n6832 ^ n6830 ;
  assign n6834 = n6833 ^ n3757 ;
  assign n6835 = n6830 ^ n6829 ;
  assign n6836 = n6835 ^ n3762 ;
  assign n6837 = ~n6834 & n6836 ;
  assign n6838 = n6837 ^ n6829 ;
  assign n6840 = n6839 ^ n6838 ;
  assign n6841 = n6840 ^ n3757 ;
  assign n6828 = n136 & n3672 ;
  assign n6842 = n6841 ^ n6828 ;
  assign n6824 = n1492 & n3720 ;
  assign n6825 = n6824 ^ n1492 ;
  assign n6826 = ~n1451 & n6825 ;
  assign n6827 = n6826 ^ n138 ;
  assign n6843 = n6842 ^ n6827 ;
  assign n6844 = n6843 ^ x134 ;
  assign n6857 = n3787 ^ n3786 ;
  assign n6851 = n3781 ^ n3748 ;
  assign n6852 = n6851 ^ n3780 ;
  assign n6853 = n3778 & n6852 ;
  assign n6854 = n6853 ^ n3778 ;
  assign n6855 = n6854 ^ n6852 ;
  assign n6858 = n6857 ^ n6855 ;
  assign n6859 = n6858 ^ n6852 ;
  assign n6860 = n6859 ^ n3786 ;
  assign n6861 = n6857 ^ n6852 ;
  assign n6862 = n6861 ^ n3762 ;
  assign n6863 = n6860 & n6862 ;
  assign n6864 = n6863 ^ n6860 ;
  assign n6865 = n6864 ^ n6860 ;
  assign n6866 = n6865 ^ n6857 ;
  assign n6856 = n6855 ^ n6852 ;
  assign n6867 = n6866 ^ n6856 ;
  assign n6868 = n6867 ^ n3786 ;
  assign n6848 = n137 & n3821 ;
  assign n6849 = n6848 ^ n137 ;
  assign n6850 = n6849 ^ n137 ;
  assign n6869 = n6868 ^ n6850 ;
  assign n6845 = n1501 & n1553 ;
  assign n6846 = ~n3778 & n6845 ;
  assign n6847 = n6846 ^ n402 ;
  assign n6870 = n6869 ^ n6847 ;
  assign n6871 = n6870 ^ x134 ;
  assign n6872 = n6870 & n6871 ;
  assign n6873 = n6872 ^ x134 ;
  assign n6874 = n6844 & n6873 ;
  assign n6875 = n6874 ^ n6873 ;
  assign n6876 = n6875 ^ n6873 ;
  assign n6877 = n6876 ^ n6872 ;
  assign n6878 = n6877 ^ n6843 ;
  assign n6893 = n6892 ^ n6878 ;
  assign n6898 = n137 & n3983 ;
  assign n6899 = n6898 ^ n137 ;
  assign n6900 = n6899 ^ n137 ;
  assign n6894 = n138 & n3859 ;
  assign n6895 = n6894 ^ n138 ;
  assign n6896 = n6895 ^ n3859 ;
  assign n6897 = n6896 ^ n138 ;
  assign n6901 = n6900 ^ n6897 ;
  assign n6943 = n1180 & n3957 ;
  assign n6944 = n6943 ^ n1180 ;
  assign n6945 = n6944 ^ n1180 ;
  assign n6946 = ~n6901 & n6945 ;
  assign n6947 = n6946 ^ n6945 ;
  assign n6948 = n6947 ^ n6945 ;
  assign n6922 = n1003 & n1942 ;
  assign n6923 = n6922 ^ n402 ;
  assign n6924 = n3894 & n6923 ;
  assign n6925 = n6924 ^ n6923 ;
  assign n6915 = n137 & n3911 ;
  assign n6916 = n6915 ^ n137 ;
  assign n6919 = n3917 & n6916 ;
  assign n6917 = n3914 & n6916 ;
  assign n6918 = n6917 ^ n6916 ;
  assign n6920 = n6919 ^ n6918 ;
  assign n6921 = n6920 ^ n137 ;
  assign n6926 = n6925 ^ n6921 ;
  assign n6911 = n1094 & n1923 ;
  assign n6912 = n3894 & n6911 ;
  assign n6913 = n6912 ^ n6911 ;
  assign n6914 = n6913 ^ n402 ;
  assign n6927 = n6926 ^ n6914 ;
  assign n6937 = n2748 & n3845 ;
  assign n6938 = n6937 ^ n2748 ;
  assign n6939 = n6938 ^ n2748 ;
  assign n6940 = n6927 & n6939 ;
  assign n6941 = n6940 ^ n6939 ;
  assign n6931 = n3937 & n4441 ;
  assign n6932 = n6931 ^ n4441 ;
  assign n6933 = n6932 ^ n4441 ;
  assign n6934 = n6927 & n6933 ;
  assign n6935 = n6934 ^ n6933 ;
  assign n6928 = x134 & n6927 ;
  assign n6929 = n6928 ^ x134 ;
  assign n6930 = n6929 ^ n6927 ;
  assign n6936 = n6935 ^ n6930 ;
  assign n6942 = n6941 ^ n6936 ;
  assign n6949 = n6948 ^ n6942 ;
  assign n6908 = x134 & ~n6901 ;
  assign n6909 = n6908 ^ x134 ;
  assign n6910 = n6909 ^ x134 ;
  assign n6950 = n6949 ^ n6910 ;
  assign n6902 = n1949 & n3877 ;
  assign n6903 = n6902 ^ n1949 ;
  assign n6904 = n6903 ^ n1949 ;
  assign n6905 = ~n6901 & n6904 ;
  assign n6906 = n6905 ^ n6904 ;
  assign n6907 = n6906 ^ n6904 ;
  assign n6951 = n6950 ^ n6907 ;
  assign n6963 = n679 ^ n677 ;
  assign n6964 = n6963 ^ n399 ;
  assign n6965 = n6964 ^ x134 ;
  assign n6954 = n5984 ^ n402 ;
  assign n6955 = n6954 ^ x134 ;
  assign n6956 = n404 & n6955 ;
  assign n6957 = n6956 ^ n5984 ;
  assign n6958 = n6957 ^ n276 ;
  assign n6959 = n401 & n6958 ;
  assign n6960 = n6959 ^ n6958 ;
  assign n6961 = n6960 ^ n6956 ;
  assign n6962 = n6961 ^ n5984 ;
  assign n6966 = n6965 ^ n6962 ;
  assign n6952 = n278 & n341 ;
  assign n6953 = n6952 ^ n278 ;
  assign n6967 = n6966 ^ n6953 ;
  assign n6998 = n1331 & n1949 ;
  assign n6999 = ~n849 & n6998 ;
  assign n7000 = n6999 ^ n6998 ;
  assign n7001 = n7000 ^ n6998 ;
  assign n6994 = n1254 & n2748 ;
  assign n6995 = n1099 & n6994 ;
  assign n6996 = n6995 ^ n6994 ;
  assign n6989 = n1174 & n4441 ;
  assign n6990 = n6989 ^ x134 ;
  assign n6991 = n1099 & n6990 ;
  assign n6992 = n6991 ^ n1099 ;
  assign n6993 = n6992 ^ n6990 ;
  assign n6997 = n6996 ^ n6993 ;
  assign n7002 = n7001 ^ n6997 ;
  assign n6979 = n946 ^ n943 ;
  assign n6980 = n6979 ^ x134 ;
  assign n6981 = ~n942 & ~n6980 ;
  assign n6982 = n6981 ^ n942 ;
  assign n6983 = n6982 ^ n6980 ;
  assign n6984 = n6983 ^ n942 ;
  assign n6985 = n6984 ^ n6980 ;
  assign n6986 = n6985 ^ n6979 ;
  assign n6987 = n6986 ^ n849 ;
  assign n6968 = n1899 ^ n930 ;
  assign n6969 = n1899 & n6968 ;
  assign n6970 = n6969 ^ n1899 ;
  assign n6971 = n6970 ^ n1899 ;
  assign n6972 = n6971 ^ n6968 ;
  assign n6973 = n6972 ^ n930 ;
  assign n6974 = n6973 ^ n849 ;
  assign n6975 = ~n849 & ~n6974 ;
  assign n6976 = n6975 ^ n6974 ;
  assign n6977 = n6976 ^ n6972 ;
  assign n6978 = n6977 ^ n930 ;
  assign n6988 = n6987 ^ n6978 ;
  assign n7003 = n7002 ^ n6988 ;
  assign n7004 = n1571 ^ n1569 ;
  assign n7005 = n7004 ^ n1434 ;
  assign n7041 = n1949 & n1999 ;
  assign n7042 = n7041 ^ n1949 ;
  assign n7043 = n7042 ^ n1949 ;
  assign n7044 = ~n1668 & n7043 ;
  assign n7045 = n7044 ^ n7043 ;
  assign n7046 = n7045 ^ n7043 ;
  assign n7035 = n1259 & n1858 ;
  assign n7036 = n7035 ^ n1259 ;
  assign n7037 = n1948 & n7036 ;
  assign n7038 = n7037 ^ n7036 ;
  assign n7039 = n7038 ^ n7036 ;
  assign n7030 = n1904 ^ n1898 ;
  assign n7031 = n1858 & n7030 ;
  assign n7032 = n7031 ^ n1858 ;
  assign n7033 = n7032 ^ n7030 ;
  assign n7027 = n850 & n1898 ;
  assign n7028 = n1858 & n7027 ;
  assign n7029 = n7028 ^ n7027 ;
  assign n7034 = n7033 ^ n7029 ;
  assign n7040 = n7039 ^ n7034 ;
  assign n7047 = n7046 ^ n7040 ;
  assign n7017 = n1731 ^ n1728 ;
  assign n7018 = n7017 ^ x134 ;
  assign n7019 = ~n1727 & ~n7018 ;
  assign n7020 = n7019 ^ n1727 ;
  assign n7021 = n7020 ^ n7018 ;
  assign n7022 = n7021 ^ n1727 ;
  assign n7023 = n7022 ^ n7018 ;
  assign n7024 = n7023 ^ n7017 ;
  assign n7025 = n7024 ^ n1668 ;
  assign n7006 = n3612 ^ n1715 ;
  assign n7007 = n3612 & n7006 ;
  assign n7008 = n7007 ^ n3612 ;
  assign n7009 = n7008 ^ n3612 ;
  assign n7010 = n7009 ^ n7006 ;
  assign n7011 = n7010 ^ n1715 ;
  assign n7012 = n7011 ^ n1668 ;
  assign n7013 = ~n1668 & ~n7012 ;
  assign n7014 = n7013 ^ n7012 ;
  assign n7015 = n7014 ^ n7010 ;
  assign n7016 = n7015 ^ n1715 ;
  assign n7026 = n7025 ^ n7016 ;
  assign n7048 = n7047 ^ n7026 ;
  assign n7052 = ~n2141 & n6955 ;
  assign n7053 = n7052 ^ n6955 ;
  assign n7054 = n7053 ^ n6955 ;
  assign n7055 = n7054 ^ n5984 ;
  assign n7056 = n7055 ^ n2140 ;
  assign n7057 = n7054 ^ n2070 ;
  assign n7058 = n7057 ^ x134 ;
  assign n7059 = ~n7056 & n7058 ;
  assign n7060 = n7059 ^ n7058 ;
  assign n7061 = n7060 ^ n7056 ;
  assign n7062 = n7061 ^ n7058 ;
  assign n7063 = n7062 ^ n5984 ;
  assign n7051 = n2139 ^ n2138 ;
  assign n7064 = n7063 ^ n7051 ;
  assign n7065 = n7064 ^ n2071 ;
  assign n7049 = n2046 & n2061 ;
  assign n7050 = n7049 ^ n2046 ;
  assign n7066 = n7065 ^ n7050 ;
  assign n7098 = ~n2366 & n5759 ;
  assign n7099 = n7098 ^ n5759 ;
  assign n7091 = n2295 ^ n2293 ;
  assign n7095 = n2344 & n7091 ;
  assign n7096 = n7095 ^ n2344 ;
  assign n7092 = n2323 & n7091 ;
  assign n7093 = n7092 ^ n2323 ;
  assign n7094 = n7093 ^ n7091 ;
  assign n7097 = n7096 ^ n7094 ;
  assign n7100 = n7099 ^ n7097 ;
  assign n7081 = n2240 ^ n2237 ;
  assign n7082 = n7081 ^ x134 ;
  assign n7083 = ~n2236 & ~n7082 ;
  assign n7084 = n7083 ^ n2236 ;
  assign n7085 = n7084 ^ n7082 ;
  assign n7086 = n7085 ^ n2236 ;
  assign n7087 = n7086 ^ n7082 ;
  assign n7088 = n7087 ^ n7081 ;
  assign n7089 = n7088 ^ n2203 ;
  assign n7067 = n2203 ^ n1899 ;
  assign n7068 = n2222 ^ n1899 ;
  assign n7069 = n2222 & n7068 ;
  assign n7070 = n7069 ^ n2222 ;
  assign n7071 = n7070 ^ n7068 ;
  assign n7072 = n7071 ^ n2222 ;
  assign n7073 = n7072 ^ n1899 ;
  assign n7074 = ~n7067 & ~n7073 ;
  assign n7075 = n7074 ^ n7067 ;
  assign n7076 = n7075 ^ n7073 ;
  assign n7077 = n7076 ^ n7067 ;
  assign n7078 = n7077 ^ n7073 ;
  assign n7079 = n7078 ^ n7072 ;
  assign n7080 = n7079 ^ n2203 ;
  assign n7090 = n7089 ^ n7080 ;
  assign n7101 = n7100 ^ n7090 ;
  assign n7103 = n2396 & n2434 ;
  assign n7104 = n7103 ^ n2434 ;
  assign n7105 = n7104 ^ n2434 ;
  assign n7102 = n2502 ^ n2500 ;
  assign n7106 = n7105 ^ n7102 ;
  assign n7138 = n1949 & n2708 ;
  assign n7139 = n7138 ^ n1949 ;
  assign n7140 = n7139 ^ n1949 ;
  assign n7141 = ~n2551 & n7140 ;
  assign n7142 = n7141 ^ n7140 ;
  assign n7143 = n7142 ^ n7140 ;
  assign n7131 = n2644 ^ n2642 ;
  assign n7135 = n2688 & n7131 ;
  assign n7136 = n7135 ^ n2688 ;
  assign n7132 = n2665 & n7131 ;
  assign n7133 = n7132 ^ n2665 ;
  assign n7134 = n7133 ^ n7131 ;
  assign n7137 = n7136 ^ n7134 ;
  assign n7144 = n7143 ^ n7137 ;
  assign n7121 = n2588 ^ n2585 ;
  assign n7122 = n7121 ^ x134 ;
  assign n7123 = ~n2584 & ~n7122 ;
  assign n7124 = n7123 ^ n2584 ;
  assign n7125 = n7124 ^ n7122 ;
  assign n7126 = n7125 ^ n2584 ;
  assign n7127 = n7126 ^ n7122 ;
  assign n7128 = n7127 ^ n7121 ;
  assign n7129 = n7128 ^ n2551 ;
  assign n7107 = n2551 ^ n1899 ;
  assign n7108 = n2570 ^ n1899 ;
  assign n7109 = n2570 & n7108 ;
  assign n7110 = n7109 ^ n2570 ;
  assign n7111 = n7110 ^ n7108 ;
  assign n7112 = n7111 ^ n2570 ;
  assign n7113 = n7112 ^ n1899 ;
  assign n7114 = ~n7107 & ~n7113 ;
  assign n7115 = n7114 ^ n7107 ;
  assign n7116 = n7115 ^ n7113 ;
  assign n7117 = n7116 ^ n7107 ;
  assign n7118 = n7117 ^ n7113 ;
  assign n7119 = n7118 ^ n7112 ;
  assign n7120 = n7119 ^ n2551 ;
  assign n7130 = n7129 ^ n7120 ;
  assign n7145 = n7144 ^ n7130 ;
  assign n7161 = n2747 ^ n1949 ;
  assign n7162 = n2844 ^ n1949 ;
  assign n7163 = ~n2844 & n7162 ;
  assign n7164 = n7163 ^ n1949 ;
  assign n7165 = ~n7161 & ~n7164 ;
  assign n7166 = n7165 ^ n7163 ;
  assign n7167 = n7166 ^ n2747 ;
  assign n7154 = n2818 & n4441 ;
  assign n7155 = n7154 ^ x134 ;
  assign n7156 = n7155 ^ x134 ;
  assign n7157 = n2807 & ~n7156 ;
  assign n7158 = n7157 ^ n7155 ;
  assign n7159 = n7158 ^ n2790 ;
  assign n7150 = n2792 ^ n2790 ;
  assign n7151 = n2804 & n7150 ;
  assign n7152 = n7151 ^ n2804 ;
  assign n7153 = n7152 ^ n7150 ;
  assign n7160 = n7159 ^ n7153 ;
  assign n7168 = n7167 ^ n7160 ;
  assign n7146 = n1180 & n2758 ;
  assign n7147 = n7146 ^ x134 ;
  assign n7148 = n2747 & n7147 ;
  assign n7149 = n7148 ^ n7147 ;
  assign n7169 = n7168 ^ n7149 ;
  assign n7191 = n1949 & n3038 ;
  assign n7192 = n7191 ^ n1949 ;
  assign n7193 = n7192 ^ n1949 ;
  assign n7194 = ~n2900 & n7193 ;
  assign n7195 = n7194 ^ n7193 ;
  assign n7196 = n7195 ^ n7193 ;
  assign n7190 = n3024 ^ n3022 ;
  assign n7197 = n7196 ^ n7190 ;
  assign n7181 = n2928 ^ n2915 ;
  assign n7182 = n7181 ^ x134 ;
  assign n7183 = ~n2926 & n7182 ;
  assign n7184 = n7183 ^ n7182 ;
  assign n7185 = n7184 ^ n2926 ;
  assign n7186 = n7185 ^ n7182 ;
  assign n7187 = n7186 ^ n7181 ;
  assign n7188 = n7187 ^ n2900 ;
  assign n7170 = n2900 ^ n1899 ;
  assign n7171 = n2915 ^ n1899 ;
  assign n7172 = n2915 & n7171 ;
  assign n7173 = n7172 ^ n7171 ;
  assign n7174 = n7173 ^ n1899 ;
  assign n7175 = ~n7170 & n7174 ;
  assign n7176 = n7175 ^ n7174 ;
  assign n7177 = n7176 ^ n7170 ;
  assign n7178 = n7177 ^ n7174 ;
  assign n7179 = n7178 ^ n7173 ;
  assign n7180 = n7179 ^ n2900 ;
  assign n7189 = n7188 ^ n7180 ;
  assign n7198 = n7197 ^ n7189 ;
  assign n7203 = n3074 & n3108 ;
  assign n7204 = n7203 ^ n3108 ;
  assign n7199 = n3169 ^ n3167 ;
  assign n7200 = n3138 & n7199 ;
  assign n7201 = n7200 ^ n3138 ;
  assign n7202 = n7201 ^ n7199 ;
  assign n7205 = n7204 ^ n7202 ;
  assign n7241 = n1949 & n3359 ;
  assign n7242 = n7241 ^ n1949 ;
  assign n7243 = n7242 ^ n1949 ;
  assign n7244 = n3216 & n7243 ;
  assign n7245 = n7244 ^ n7243 ;
  assign n7236 = n2748 & n3334 ;
  assign n7237 = n3303 & n7236 ;
  assign n7238 = n7237 ^ n7236 ;
  assign n7239 = n7238 ^ n7236 ;
  assign n7228 = n1259 & n3317 ;
  assign n7229 = n7228 ^ n1259 ;
  assign n7230 = n7229 ^ n1259 ;
  assign n7231 = n7230 ^ x134 ;
  assign n7232 = n3303 & n7231 ;
  assign n7233 = n7232 ^ n7231 ;
  assign n7234 = n7233 ^ n3303 ;
  assign n7235 = n7234 ^ n7231 ;
  assign n7240 = n7239 ^ n7235 ;
  assign n7246 = n7245 ^ n7240 ;
  assign n7219 = n3252 ^ n3249 ;
  assign n7220 = n7219 ^ x134 ;
  assign n7221 = n3248 & ~n7220 ;
  assign n7222 = n7221 ^ n3248 ;
  assign n7223 = n7222 ^ n3248 ;
  assign n7224 = n7223 ^ n7220 ;
  assign n7225 = n7224 ^ n7219 ;
  assign n7226 = n7225 ^ n3216 ;
  assign n7206 = n3216 ^ n1899 ;
  assign n7207 = n3235 ^ n1899 ;
  assign n7208 = n3235 & n7207 ;
  assign n7209 = n7208 ^ n3235 ;
  assign n7210 = n7209 ^ n7207 ;
  assign n7211 = n7210 ^ n3235 ;
  assign n7212 = n7211 ^ n1899 ;
  assign n7213 = n7206 & ~n7212 ;
  assign n7214 = n7213 ^ n7206 ;
  assign n7215 = n7214 ^ n7206 ;
  assign n7216 = n7215 ^ n7212 ;
  assign n7217 = n7216 ^ n7211 ;
  assign n7218 = n7217 ^ n3216 ;
  assign n7227 = n7226 ^ n7218 ;
  assign n7247 = n7246 ^ n7227 ;
  assign n7253 = n3398 ^ n1949 ;
  assign n7254 = n3508 ^ n1949 ;
  assign n7255 = ~n3508 & n7254 ;
  assign n7256 = n7255 ^ n1949 ;
  assign n7257 = n7253 & ~n7256 ;
  assign n7258 = n7257 ^ n7255 ;
  assign n7259 = n7258 ^ n3398 ;
  assign n7252 = n3489 ^ n3486 ;
  assign n7260 = n7259 ^ n7252 ;
  assign n7248 = n1180 & n3408 ;
  assign n7249 = n7248 ^ x134 ;
  assign n7250 = ~n3398 & n7249 ;
  assign n7251 = n7250 ^ n7249 ;
  assign n7261 = n7260 ^ n7251 ;
  assign n7286 = n1949 & n3655 ;
  assign n7287 = n7286 ^ n1949 ;
  assign n7288 = n7287 ^ n1949 ;
  assign n7289 = ~n3544 & n7288 ;
  assign n7290 = n7289 ^ n7288 ;
  assign n7291 = n7290 ^ n7288 ;
  assign n7280 = n3633 & n4441 ;
  assign n7281 = n7280 ^ n4441 ;
  assign n7282 = n7281 ^ n4441 ;
  assign n7283 = n3597 & n7282 ;
  assign n7284 = n7283 ^ n7282 ;
  assign n7275 = n3619 ^ n3611 ;
  assign n7276 = n3597 & n7275 ;
  assign n7277 = n7276 ^ n3597 ;
  assign n7278 = n7277 ^ n7275 ;
  assign n7270 = n1669 & n3611 ;
  assign n7271 = n7270 ^ n1669 ;
  assign n7272 = n7271 ^ n1669 ;
  assign n7273 = n3597 & n7272 ;
  assign n7274 = n7273 ^ n7272 ;
  assign n7279 = n7278 ^ n7274 ;
  assign n7285 = n7284 ^ n7279 ;
  assign n7292 = n7291 ^ n7285 ;
  assign n7266 = ~n3544 & n3564 ;
  assign n7267 = n7266 ^ n3564 ;
  assign n7268 = n7267 ^ n3564 ;
  assign n7262 = n1899 & n3558 ;
  assign n7263 = ~n3544 & n7262 ;
  assign n7264 = n7263 ^ n7262 ;
  assign n7265 = n7264 ^ n7262 ;
  assign n7269 = n7268 ^ n7265 ;
  assign n7293 = n7292 ^ n7269 ;
  assign n7299 = n1180 & n3710 ;
  assign n7300 = ~n3684 & n7299 ;
  assign n7295 = n1949 & n3694 ;
  assign n7296 = n7295 ^ x134 ;
  assign n7297 = n3684 & n7296 ;
  assign n7298 = n7297 ^ n7296 ;
  assign n7301 = n7300 ^ n7298 ;
  assign n7294 = n3834 ^ n3833 ;
  assign n7302 = n7301 ^ n7294 ;
  assign n7329 = n1949 & n3983 ;
  assign n7330 = n7329 ^ n1949 ;
  assign n7331 = n7330 ^ n1949 ;
  assign n7332 = ~n3863 & n7331 ;
  assign n7333 = n7332 ^ n7331 ;
  assign n7334 = n7333 ^ n7331 ;
  assign n7323 = n3957 & n4441 ;
  assign n7324 = n7323 ^ n4441 ;
  assign n7325 = n7324 ^ n4441 ;
  assign n7326 = n3925 & n7325 ;
  assign n7327 = n7326 ^ n7325 ;
  assign n7318 = n3944 ^ n3937 ;
  assign n7319 = n3925 & n7318 ;
  assign n7320 = n7319 ^ n3925 ;
  assign n7321 = n7320 ^ n7318 ;
  assign n7313 = n1669 & n3937 ;
  assign n7314 = n7313 ^ n1669 ;
  assign n7315 = n7314 ^ n1669 ;
  assign n7316 = n3925 & n7315 ;
  assign n7317 = n7316 ^ n7315 ;
  assign n7322 = n7321 ^ n7317 ;
  assign n7328 = n7327 ^ n7322 ;
  assign n7335 = n7334 ^ n7328 ;
  assign n7309 = ~n3863 & n3885 ;
  assign n7310 = n7309 ^ n3885 ;
  assign n7311 = n7310 ^ n3885 ;
  assign n7303 = n1899 & n3877 ;
  assign n7304 = n7303 ^ n1899 ;
  assign n7305 = n7304 ^ n1899 ;
  assign n7306 = ~n3863 & n7305 ;
  assign n7307 = n7306 ^ n7305 ;
  assign n7308 = n7307 ^ n7305 ;
  assign n7312 = n7311 ^ n7308 ;
  assign n7336 = n7335 ^ n7312 ;
  assign n7354 = n2748 ^ n399 ;
  assign n7355 = ~n4038 & ~n7354 ;
  assign n7356 = n7355 ^ n4037 ;
  assign n7357 = n7356 ^ n4038 ;
  assign n7358 = n2748 ^ x134 ;
  assign n7359 = n7358 ^ n4044 ;
  assign n7360 = ~n7357 & ~n7359 ;
  assign n7361 = n7360 ^ n2748 ;
  assign n7351 = x134 & n272 ;
  assign n7352 = n402 & n7351 ;
  assign n7342 = n607 & n1180 ;
  assign n7343 = n7342 ^ x134 ;
  assign n7344 = n7343 ^ n4005 ;
  assign n7345 = n7344 ^ x134 ;
  assign n7346 = n4016 & n7345 ;
  assign n7347 = n7346 ^ n7345 ;
  assign n7348 = n7347 ^ n7343 ;
  assign n7337 = n339 & n4441 ;
  assign n7338 = n7337 ^ x134 ;
  assign n7339 = n4006 & n7338 ;
  assign n7340 = n7339 ^ n7337 ;
  assign n7341 = n7340 ^ n4005 ;
  assign n7349 = n7348 ^ n7341 ;
  assign n7350 = n7349 ^ n4026 ;
  assign n7353 = n7352 ^ n7350 ;
  assign n7362 = n7361 ^ n7353 ;
  assign n7363 = n7362 ^ n3992 ;
  assign n7380 = n845 & n1949 ;
  assign n7381 = n7380 ^ n1949 ;
  assign n7382 = n7381 ^ n1949 ;
  assign n7383 = n4055 & n7382 ;
  assign n7384 = n7383 ^ n7382 ;
  assign n7374 = n930 & n4441 ;
  assign n7375 = n7374 ^ n4441 ;
  assign n7376 = n7375 ^ n4441 ;
  assign n7377 = n4075 & n7376 ;
  assign n7378 = n7377 ^ n7376 ;
  assign n7368 = ~x134 & n137 ;
  assign n7369 = n1174 & n7368 ;
  assign n7370 = n7369 ^ x134 ;
  assign n7371 = n4075 & n7370 ;
  assign n7372 = n7371 ^ n4075 ;
  assign n7373 = n7372 ^ n7370 ;
  assign n7379 = n7378 ^ n7373 ;
  assign n7385 = n7384 ^ n7379 ;
  assign n7364 = n1180 & n1331 ;
  assign n7365 = n4055 & n7364 ;
  assign n7366 = n7365 ^ n7364 ;
  assign n7367 = n7366 ^ n4057 ;
  assign n7386 = n7385 ^ n7367 ;
  assign n7392 = n1180 & n1375 ;
  assign n7393 = ~n4100 & n7392 ;
  assign n7388 = n1423 & n1949 ;
  assign n7389 = n7388 ^ x134 ;
  assign n7390 = n4100 & n7389 ;
  assign n7391 = n7390 ^ n7389 ;
  assign n7394 = n7393 ^ n7391 ;
  assign n7387 = n4159 ^ n4156 ;
  assign n7395 = n7394 ^ n7387 ;
  assign n7410 = n1180 & n1999 ;
  assign n7411 = n7410 ^ n1180 ;
  assign n7412 = n7411 ^ n1180 ;
  assign n7413 = n4168 & n7412 ;
  assign n7414 = n7413 ^ n7412 ;
  assign n7406 = n1664 & n4441 ;
  assign n7407 = n4193 & n7406 ;
  assign n7408 = n7407 ^ n7406 ;
  assign n7399 = n4206 & n7368 ;
  assign n7400 = n7399 ^ n7368 ;
  assign n7401 = n7400 ^ n7368 ;
  assign n7402 = n7401 ^ x134 ;
  assign n7403 = n4193 & n7402 ;
  assign n7404 = n7403 ^ n4193 ;
  assign n7405 = n7404 ^ n7402 ;
  assign n7409 = n7408 ^ n7405 ;
  assign n7415 = n7414 ^ n7409 ;
  assign n7396 = ~n1715 & n5759 ;
  assign n7397 = n7396 ^ n5759 ;
  assign n7398 = n7397 ^ n4170 ;
  assign n7416 = n7415 ^ n7398 ;
  assign n7431 = n1949 & n2039 ;
  assign n7432 = ~n4233 & n7431 ;
  assign n7423 = n2093 & n7368 ;
  assign n7424 = n7423 ^ x134 ;
  assign n7425 = n7424 ^ x134 ;
  assign n7426 = ~n4265 & ~n7425 ;
  assign n7427 = n7426 ^ n7425 ;
  assign n7428 = n7427 ^ n7424 ;
  assign n7429 = n7428 ^ n4259 ;
  assign n7419 = n4261 ^ n4259 ;
  assign n7420 = n4262 & n7419 ;
  assign n7421 = n7420 ^ n4262 ;
  assign n7422 = n7421 ^ n7419 ;
  assign n7430 = n7429 ^ n7422 ;
  assign n7433 = n7432 ^ n7430 ;
  assign n7417 = n4225 & n4235 ;
  assign n7418 = n7417 ^ n4235 ;
  assign n7434 = n7433 ^ n7418 ;
  assign n7453 = n1949 & n2199 ;
  assign n7454 = n7453 ^ n1949 ;
  assign n7455 = n7454 ^ n1949 ;
  assign n7456 = ~n4285 & n7455 ;
  assign n7457 = n7456 ^ n7455 ;
  assign n7458 = n7457 ^ n7455 ;
  assign n7446 = n4325 & n7368 ;
  assign n7447 = n7446 ^ n7368 ;
  assign n7448 = n7447 ^ n7368 ;
  assign n7449 = n4307 & n7448 ;
  assign n7450 = n7449 ^ n7448 ;
  assign n7451 = n7450 ^ n7448 ;
  assign n7438 = n2320 & n2748 ;
  assign n7439 = n7438 ^ n2748 ;
  assign n7440 = n7439 ^ n2748 ;
  assign n7441 = n7440 ^ x134 ;
  assign n7442 = n4307 & n7441 ;
  assign n7443 = n7442 ^ n7441 ;
  assign n7444 = n7443 ^ n4307 ;
  assign n7445 = n7444 ^ n7441 ;
  assign n7452 = n7451 ^ n7445 ;
  assign n7459 = n7458 ^ n7452 ;
  assign n7435 = n1180 & ~n2366 ;
  assign n7436 = n7435 ^ n1180 ;
  assign n7437 = n7436 ^ n4288 ;
  assign n7460 = n7459 ^ n7437 ;
  assign n7466 = n4351 & n4360 ;
  assign n7467 = n7466 ^ n4360 ;
  assign n7468 = n7467 ^ n4360 ;
  assign n7461 = n4381 & n4382 ;
  assign n7462 = n7461 ^ x134 ;
  assign n7463 = ~n4378 & n7462 ;
  assign n7464 = n7463 ^ n7461 ;
  assign n7465 = n7464 ^ n4377 ;
  assign n7469 = n7468 ^ n7465 ;
  assign n7484 = n1175 & ~n2685 ;
  assign n7485 = n7484 ^ n1175 ;
  assign n7476 = n4428 ^ n4426 ;
  assign n7480 = ~n4437 & n7476 ;
  assign n7481 = n7480 ^ n7476 ;
  assign n7482 = n7481 ^ n4437 ;
  assign n7477 = n4431 & n7476 ;
  assign n7478 = n7477 ^ n4431 ;
  assign n7479 = n7478 ^ n7476 ;
  assign n7483 = n7482 ^ n7479 ;
  assign n7486 = n7485 ^ n7483 ;
  assign n7470 = n1180 & n2708 ;
  assign n7471 = n7470 ^ n1180 ;
  assign n7472 = n7471 ^ n1180 ;
  assign n7473 = n4395 & n7472 ;
  assign n7474 = n7473 ^ n7472 ;
  assign n7475 = n7474 ^ n4397 ;
  assign n7487 = n7486 ^ n7475 ;
  assign n7520 = n4515 ^ n4506 ;
  assign n7521 = n4517 & ~n7520 ;
  assign n7522 = n7521 ^ n7520 ;
  assign n7523 = n7522 ^ n2818 ;
  assign n7510 = ~n4506 & n7368 ;
  assign n7511 = n7510 ^ n137 ;
  assign n7512 = n7511 ^ n137 ;
  assign n7513 = n7511 ^ n2818 ;
  assign n7514 = n7513 ^ n137 ;
  assign n7515 = n7512 & n7514 ;
  assign n7516 = n7515 ^ n7512 ;
  assign n7517 = n7516 ^ n7512 ;
  assign n7518 = n7517 ^ n7514 ;
  assign n7508 = n1175 & ~n4484 ;
  assign n7509 = n7508 ^ n1175 ;
  assign n7519 = n7518 ^ n7509 ;
  assign n7524 = n7523 ^ n7519 ;
  assign n7490 = n4452 ^ n4447 ;
  assign n7491 = n7490 ^ n4449 ;
  assign n7492 = n7491 ^ x133 ;
  assign n7493 = n7492 ^ n4461 ;
  assign n7494 = n4446 & ~n7493 ;
  assign n7495 = n7494 ^ n7493 ;
  assign n7496 = n7495 ^ n7493 ;
  assign n7488 = n4468 ^ n4460 ;
  assign n7489 = n7488 ^ n4467 ;
  assign n7497 = n7496 ^ n7489 ;
  assign n7498 = n7497 ^ n7491 ;
  assign n7499 = n7498 ^ n4449 ;
  assign n7500 = n7489 ^ n4460 ;
  assign n7501 = ~n7499 & n7500 ;
  assign n7502 = n7501 ^ n7499 ;
  assign n7503 = n7502 ^ n7500 ;
  assign n7504 = n7503 ^ n7499 ;
  assign n7505 = n7504 ^ n7500 ;
  assign n7506 = n7505 ^ n7489 ;
  assign n7507 = n7506 ^ n4460 ;
  assign n7525 = n7524 ^ n7507 ;
  assign n7533 = n1175 & n4608 ;
  assign n7534 = n7533 ^ n1175 ;
  assign n7532 = n4601 ^ n4599 ;
  assign n7535 = n7534 ^ n7532 ;
  assign n7526 = n1180 & n3038 ;
  assign n7527 = n7526 ^ n1180 ;
  assign n7528 = n7527 ^ n1180 ;
  assign n7529 = n4529 & n7528 ;
  assign n7530 = n7529 ^ n7528 ;
  assign n7531 = n7530 ^ n4531 ;
  assign n7536 = n7535 ^ n7531 ;
  assign n7541 = n4619 & n4628 ;
  assign n7542 = n7541 ^ n4628 ;
  assign n7543 = n7542 ^ n4628 ;
  assign n7537 = n4657 & n4679 ;
  assign n7538 = n7537 ^ n4657 ;
  assign n7539 = n7538 ^ n4679 ;
  assign n7540 = n7539 ^ n4685 ;
  assign n7544 = n7543 ^ n7540 ;
  assign n7576 = n1949 & n3212 ;
  assign n7577 = n7576 ^ n1949 ;
  assign n7578 = n7577 ^ n1949 ;
  assign n7579 = n4690 & n7578 ;
  assign n7580 = n7579 ^ n7578 ;
  assign n7566 = n2748 & n3317 ;
  assign n7567 = n7566 ^ n2748 ;
  assign n7568 = n7567 ^ n2748 ;
  assign n7569 = n7568 ^ x134 ;
  assign n7570 = n4716 & n7569 ;
  assign n7571 = n7570 ^ n4716 ;
  assign n7572 = n7571 ^ n7569 ;
  assign n7573 = n7572 ^ n3235 ;
  assign n7574 = n7573 ^ n138 ;
  assign n7551 = x134 & n138 ;
  assign n7552 = n7551 ^ n138 ;
  assign n7553 = n7552 ^ x134 ;
  assign n7554 = n3249 & n7553 ;
  assign n7555 = n7554 ^ n3249 ;
  assign n7556 = n7555 ^ n7553 ;
  assign n7557 = n7556 ^ n3249 ;
  assign n7558 = n7557 ^ n7551 ;
  assign n7559 = n7558 ^ n4716 ;
  assign n7560 = n7559 ^ n3249 ;
  assign n7561 = n4718 & ~n7560 ;
  assign n7562 = n7561 ^ n7560 ;
  assign n7563 = n7562 ^ n7560 ;
  assign n7564 = n7563 ^ n7557 ;
  assign n7565 = n7564 ^ n7551 ;
  assign n7575 = n7574 ^ n7565 ;
  assign n7581 = n7580 ^ n7575 ;
  assign n7545 = n1180 & n3359 ;
  assign n7546 = n7545 ^ n1180 ;
  assign n7547 = n7546 ^ n1180 ;
  assign n7548 = n4690 & n7547 ;
  assign n7549 = n7548 ^ n7547 ;
  assign n7550 = n7549 ^ n4692 ;
  assign n7582 = n7581 ^ n7550 ;
  assign n7614 = n1949 & n3394 ;
  assign n7615 = ~n4763 & n7614 ;
  assign n7606 = n3454 & n7368 ;
  assign n7607 = n7606 ^ x134 ;
  assign n7608 = n7607 ^ x134 ;
  assign n7609 = ~n4801 & ~n7608 ;
  assign n7610 = n7609 ^ n7608 ;
  assign n7611 = n7610 ^ n7607 ;
  assign n7612 = n7611 ^ n4795 ;
  assign n7603 = n4796 ^ n4795 ;
  assign n7604 = n4798 & ~n7603 ;
  assign n7605 = n7604 ^ n7603 ;
  assign n7613 = n7612 ^ n7605 ;
  assign n7616 = n7615 ^ n7613 ;
  assign n7585 = n4756 ^ n4751 ;
  assign n7586 = n7585 ^ n4753 ;
  assign n7587 = n7586 ^ x133 ;
  assign n7588 = n7587 ^ n4764 ;
  assign n7589 = n4750 & ~n7588 ;
  assign n7590 = n7589 ^ n7588 ;
  assign n7591 = n7590 ^ n7588 ;
  assign n7583 = n4771 ^ n4763 ;
  assign n7584 = n7583 ^ n4770 ;
  assign n7592 = n7591 ^ n7584 ;
  assign n7593 = n7592 ^ n7586 ;
  assign n7594 = n7593 ^ n4753 ;
  assign n7595 = n7584 ^ n4763 ;
  assign n7596 = ~n7594 & n7595 ;
  assign n7597 = n7596 ^ n7594 ;
  assign n7598 = n7597 ^ n7595 ;
  assign n7599 = n7598 ^ n7594 ;
  assign n7600 = n7599 ^ n7595 ;
  assign n7601 = n7600 ^ n7584 ;
  assign n7602 = n7601 ^ n4763 ;
  assign n7617 = n7616 ^ n7602 ;
  assign n7638 = n1949 & n3540 ;
  assign n7639 = n7638 ^ n1949 ;
  assign n7640 = n7639 ^ n1949 ;
  assign n7641 = ~n4832 & n7640 ;
  assign n7642 = n7641 ^ n7640 ;
  assign n7643 = n7642 ^ n7640 ;
  assign n7632 = n3633 & n7368 ;
  assign n7633 = n7632 ^ n7368 ;
  assign n7634 = n7633 ^ n7368 ;
  assign n7635 = n4854 & n7634 ;
  assign n7636 = n7635 ^ n7634 ;
  assign n7626 = n1259 & n3611 ;
  assign n7627 = n7626 ^ n1259 ;
  assign n7628 = n7627 ^ n1259 ;
  assign n7629 = n4854 & n7628 ;
  assign n7630 = n7629 ^ n7628 ;
  assign n7625 = n4856 ^ n4854 ;
  assign n7631 = n7630 ^ n7625 ;
  assign n7637 = n7636 ^ n7631 ;
  assign n7644 = n7643 ^ n7637 ;
  assign n7618 = n1180 & n3655 ;
  assign n7619 = n7618 ^ n1180 ;
  assign n7620 = n7619 ^ n1180 ;
  assign n7621 = ~n4832 & n7620 ;
  assign n7622 = n7621 ^ n7620 ;
  assign n7623 = n7622 ^ n7620 ;
  assign n7624 = n7623 ^ n4835 ;
  assign n7645 = n7644 ^ n7624 ;
  assign n7650 = n4886 & n4899 ;
  assign n7651 = n7650 ^ n4899 ;
  assign n7652 = n7651 ^ n4899 ;
  assign n7646 = n4921 ^ n4919 ;
  assign n7647 = n4914 & n7646 ;
  assign n7648 = n7647 ^ n4914 ;
  assign n7649 = n7648 ^ n7646 ;
  assign n7653 = n7652 ^ n7649 ;
  assign n7674 = n1949 & n3859 ;
  assign n7675 = n7674 ^ n1949 ;
  assign n7676 = n7675 ^ n1949 ;
  assign n7677 = ~n4939 & n7676 ;
  assign n7678 = n7677 ^ n7676 ;
  assign n7679 = n7678 ^ n7676 ;
  assign n7668 = n3957 & n7368 ;
  assign n7669 = n7668 ^ n7368 ;
  assign n7670 = n7669 ^ n7368 ;
  assign n7671 = n4967 & n7670 ;
  assign n7672 = n7671 ^ n7670 ;
  assign n7662 = n1259 & n3937 ;
  assign n7663 = n7662 ^ n1259 ;
  assign n7664 = n7663 ^ n1259 ;
  assign n7665 = n4967 & n7664 ;
  assign n7666 = n7665 ^ n7664 ;
  assign n7661 = n4969 ^ n4967 ;
  assign n7667 = n7666 ^ n7661 ;
  assign n7673 = n7672 ^ n7667 ;
  assign n7680 = n7679 ^ n7673 ;
  assign n7654 = n1180 & n3983 ;
  assign n7655 = n7654 ^ n1180 ;
  assign n7656 = n7655 ^ n1180 ;
  assign n7657 = ~n4939 & n7656 ;
  assign n7658 = n7657 ^ n7656 ;
  assign n7659 = n7658 ^ n7656 ;
  assign n7660 = n7659 ^ n4942 ;
  assign n7681 = n7680 ^ n7660 ;
  assign n7699 = x134 & n202 ;
  assign n7700 = n402 & n7699 ;
  assign n7698 = n5052 ^ n5049 ;
  assign n7701 = n7700 ^ n7698 ;
  assign n7684 = n5003 ^ x133 ;
  assign n7685 = n7684 ^ n4999 ;
  assign n7686 = n4990 & ~n7685 ;
  assign n7687 = n7686 ^ n4990 ;
  assign n7688 = n7687 ^ n4990 ;
  assign n7682 = n5013 ^ n4998 ;
  assign n7683 = n7682 ^ n5010 ;
  assign n7689 = n7688 ^ n7683 ;
  assign n7690 = n7689 ^ n5003 ;
  assign n7691 = n7690 ^ n5002 ;
  assign n7692 = n7683 ^ n4998 ;
  assign n7693 = ~n7691 & n7692 ;
  assign n7694 = n7693 ^ n7692 ;
  assign n7695 = n7694 ^ n7691 ;
  assign n7696 = n7695 ^ n7683 ;
  assign n7697 = n7696 ^ n4998 ;
  assign n7702 = n7701 ^ n7697 ;
  assign n7721 = n763 & n1949 ;
  assign n7722 = n7721 ^ n1949 ;
  assign n7723 = n7722 ^ n1949 ;
  assign n7724 = ~n5073 & n7723 ;
  assign n7725 = n7724 ^ n7723 ;
  assign n7726 = n7725 ^ n7723 ;
  assign n7715 = n930 & n7368 ;
  assign n7716 = n7715 ^ n7368 ;
  assign n7717 = n7716 ^ n7368 ;
  assign n7718 = n5097 & n7717 ;
  assign n7719 = n7718 ^ n7717 ;
  assign n7710 = n1174 & n1259 ;
  assign n7711 = n7710 ^ x134 ;
  assign n7712 = n5097 & n7711 ;
  assign n7713 = n7712 ^ n5097 ;
  assign n7714 = n7713 ^ n7711 ;
  assign n7720 = n7719 ^ n7714 ;
  assign n7727 = n7726 ^ n7720 ;
  assign n7703 = n845 & n1180 ;
  assign n7704 = n7703 ^ n1180 ;
  assign n7705 = n7704 ^ n1180 ;
  assign n7706 = ~n5073 & n7705 ;
  assign n7707 = n7706 ^ n7705 ;
  assign n7708 = n7707 ^ n7705 ;
  assign n7709 = n7708 ^ n5076 ;
  assign n7728 = n7727 ^ n7709 ;
  assign n7733 = n5126 & n5140 ;
  assign n7734 = n7733 ^ n5140 ;
  assign n7729 = n5170 ^ n5168 ;
  assign n7730 = n5159 & n7729 ;
  assign n7731 = n7730 ^ n5159 ;
  assign n7732 = n7731 ^ n7729 ;
  assign n7735 = n7734 ^ n7732 ;
  assign n7752 = n1175 & ~n1948 ;
  assign n7753 = n7752 ^ n1175 ;
  assign n7746 = n1999 & n4441 ;
  assign n7747 = n7746 ^ n4441 ;
  assign n7748 = n7747 ^ n4441 ;
  assign n7749 = n5202 & n7748 ;
  assign n7750 = n7749 ^ n7748 ;
  assign n7739 = n1259 & n4206 ;
  assign n7740 = n7739 ^ n1259 ;
  assign n7741 = n7740 ^ n1259 ;
  assign n7742 = n7741 ^ x134 ;
  assign n7743 = n5202 & n7742 ;
  assign n7744 = n7743 ^ n5202 ;
  assign n7745 = n7744 ^ n7742 ;
  assign n7751 = n7750 ^ n7745 ;
  assign n7754 = n7753 ^ n7751 ;
  assign n7736 = n1180 & ~n1715 ;
  assign n7737 = n7736 ^ n1180 ;
  assign n7738 = n7737 ^ n5182 ;
  assign n7755 = n7754 ^ n7738 ;
  assign n7773 = n1949 & n2017 ;
  assign n7774 = n5237 & n7773 ;
  assign n7775 = n7774 ^ n7773 ;
  assign n7772 = n5283 ^ n5280 ;
  assign n7776 = n7775 ^ n7772 ;
  assign n7758 = n5223 ^ x133 ;
  assign n7759 = n7758 ^ n5238 ;
  assign n7760 = n5219 & n7759 ;
  assign n7761 = n7760 ^ n5219 ;
  assign n7756 = n5244 ^ n5237 ;
  assign n7757 = n7756 ^ n5243 ;
  assign n7762 = n7761 ^ n7757 ;
  assign n7763 = n7762 ^ n5223 ;
  assign n7764 = n7763 ^ n5222 ;
  assign n7765 = n7757 ^ n5237 ;
  assign n7766 = n7764 & n7765 ;
  assign n7767 = n7766 ^ n7764 ;
  assign n7768 = n7767 ^ n7765 ;
  assign n7769 = n7768 ^ n7764 ;
  assign n7770 = n7769 ^ n7757 ;
  assign n7771 = n7770 ^ n5237 ;
  assign n7777 = n7776 ^ n7771 ;
  assign n7797 = n1949 & n2175 ;
  assign n7798 = n7797 ^ n1949 ;
  assign n7799 = n7798 ^ n1949 ;
  assign n7800 = ~n5296 & n7799 ;
  assign n7801 = n7800 ^ n7799 ;
  assign n7802 = n7801 ^ n7799 ;
  assign n7792 = n5332 ^ n5324 ;
  assign n7793 = ~n5336 & n7792 ;
  assign n7794 = n7793 ^ n7792 ;
  assign n7795 = n7794 ^ n5336 ;
  assign n7785 = n2222 & n7368 ;
  assign n7786 = n7785 ^ n7368 ;
  assign n7787 = n7786 ^ n7368 ;
  assign n7788 = n7787 ^ x134 ;
  assign n7789 = n5324 & n7788 ;
  assign n7790 = n7789 ^ n5324 ;
  assign n7791 = n7790 ^ n7788 ;
  assign n7796 = n7795 ^ n7791 ;
  assign n7803 = n7802 ^ n7796 ;
  assign n7778 = n1180 & n2199 ;
  assign n7779 = n7778 ^ n1180 ;
  assign n7780 = n7779 ^ n1180 ;
  assign n7781 = ~n5296 & n7780 ;
  assign n7782 = n7781 ^ n7780 ;
  assign n7783 = n7782 ^ n7780 ;
  assign n7784 = n7783 ^ n5299 ;
  assign n7804 = n7803 ^ n7784 ;
  assign n7806 = n5354 & n5365 ;
  assign n7807 = n7806 ^ n5365 ;
  assign n7805 = n5398 ^ n5395 ;
  assign n7808 = n7807 ^ n7805 ;
  assign n7834 = n1175 & ~n2662 ;
  assign n7835 = n7834 ^ n1175 ;
  assign n7824 = n2708 & n4441 ;
  assign n7825 = n7824 ^ n4441 ;
  assign n7826 = n7825 ^ n4441 ;
  assign n7827 = n7826 ^ x134 ;
  assign n7828 = n5431 & n7827 ;
  assign n7829 = n7828 ^ n5431 ;
  assign n7830 = n7829 ^ n7827 ;
  assign n7831 = n7830 ^ n2570 ;
  assign n7832 = n7831 ^ n137 ;
  assign n7812 = n3612 ^ n137 ;
  assign n7813 = n7812 ^ x134 ;
  assign n7814 = n2585 & n7813 ;
  assign n7815 = n7814 ^ n7813 ;
  assign n7816 = n7815 ^ n2585 ;
  assign n7817 = n7816 ^ n3612 ;
  assign n7818 = n7817 ^ n5431 ;
  assign n7819 = n7818 ^ n2585 ;
  assign n7820 = n5433 & n7819 ;
  assign n7821 = n7820 ^ n7819 ;
  assign n7822 = n7821 ^ n7816 ;
  assign n7823 = n7822 ^ n3612 ;
  assign n7833 = n7832 ^ n7823 ;
  assign n7836 = n7835 ^ n7833 ;
  assign n7809 = ~n2685 & n6307 ;
  assign n7810 = n7809 ^ n6307 ;
  assign n7811 = n7810 ^ n5408 ;
  assign n7837 = n7836 ^ n7811 ;
  assign n7838 = n5470 ^ n5467 ;
  assign n7855 = n5472 & ~n7838 ;
  assign n7856 = n7855 ^ n5499 ;
  assign n7843 = n5499 ^ x134 ;
  assign n7844 = n5507 ^ n5503 ;
  assign n7845 = x134 & n7844 ;
  assign n7846 = n7845 ^ x134 ;
  assign n7847 = n7846 ^ n7844 ;
  assign n7848 = n7847 ^ n5499 ;
  assign n7849 = n7848 ^ x134 ;
  assign n7850 = n7849 ^ n7844 ;
  assign n7851 = n7843 & n7850 ;
  assign n7852 = n7851 ^ n7850 ;
  assign n7853 = n7852 ^ n7843 ;
  assign n7854 = n7853 ^ n7847 ;
  assign n7857 = n7856 ^ n7854 ;
  assign n7841 = n5503 ^ x134 ;
  assign n7842 = n7841 ^ n5507 ;
  assign n7858 = n7857 ^ n7842 ;
  assign n7839 = n5512 & ~n7838 ;
  assign n7840 = n7839 ^ n7838 ;
  assign n7859 = n7858 ^ n7840 ;
  assign n7872 = n5545 & n5549 ;
  assign n7873 = n7872 ^ n5545 ;
  assign n7871 = n5545 & n5556 ;
  assign n7874 = n7873 ^ n7871 ;
  assign n7863 = n3038 & n4441 ;
  assign n7864 = n7863 ^ n4441 ;
  assign n7865 = n7864 ^ n4441 ;
  assign n7866 = n7865 ^ x134 ;
  assign n7867 = n5575 & n7866 ;
  assign n7868 = n7867 ^ n5575 ;
  assign n7869 = n7868 ^ n7866 ;
  assign n7860 = n2915 & n7368 ;
  assign n7861 = n5575 & n7860 ;
  assign n7862 = n7861 ^ n7860 ;
  assign n7870 = n7869 ^ n7862 ;
  assign n7875 = n7874 ^ n7870 ;
  assign n7881 = n1949 & n3086 ;
  assign n7882 = ~n5593 & n7881 ;
  assign n7877 = n1180 & n3102 ;
  assign n7878 = n7877 ^ x134 ;
  assign n7879 = n5593 & n7878 ;
  assign n7880 = n7879 ^ n7878 ;
  assign n7883 = n7882 ^ n7880 ;
  assign n7876 = n5646 ^ n5645 ;
  assign n7884 = n7883 ^ n7876 ;
  assign n7912 = n1949 & n3188 ;
  assign n7913 = ~n5653 & n7912 ;
  assign n7914 = n7913 ^ n7912 ;
  assign n7915 = n7914 ^ n7912 ;
  assign n7902 = n3359 & n4441 ;
  assign n7903 = n7902 ^ n4441 ;
  assign n7904 = n7903 ^ n4441 ;
  assign n7905 = n7904 ^ x134 ;
  assign n7906 = n5681 & n7905 ;
  assign n7907 = n7906 ^ n5681 ;
  assign n7908 = n7907 ^ n7905 ;
  assign n7909 = n7908 ^ n3235 ;
  assign n7910 = n7909 ^ n137 ;
  assign n7892 = n3249 & n7813 ;
  assign n7893 = n7892 ^ n7813 ;
  assign n7894 = n7893 ^ n3249 ;
  assign n7895 = n7894 ^ n3612 ;
  assign n7896 = n7895 ^ n5681 ;
  assign n7897 = n7896 ^ n3249 ;
  assign n7898 = n5683 & n7897 ;
  assign n7899 = n7898 ^ n7897 ;
  assign n7900 = n7899 ^ n7894 ;
  assign n7901 = n7900 ^ n3612 ;
  assign n7911 = n7910 ^ n7901 ;
  assign n7916 = n7915 ^ n7911 ;
  assign n7885 = n1180 & n3212 ;
  assign n7886 = n7885 ^ n1180 ;
  assign n7887 = n7886 ^ n1180 ;
  assign n7888 = ~n5653 & n7887 ;
  assign n7889 = n7888 ^ n7887 ;
  assign n7890 = n7889 ^ n7887 ;
  assign n7891 = n7890 ^ n5656 ;
  assign n7917 = n7916 ^ n7891 ;
  assign n7918 = n5720 ^ n5717 ;
  assign n7921 = n5722 & ~n7918 ;
  assign n7922 = n7921 ^ n5751 ;
  assign n7919 = n5754 & ~n7918 ;
  assign n7920 = n7919 ^ n7918 ;
  assign n7923 = n7922 ^ n7920 ;
  assign n7932 = n2348 & ~n3633 ;
  assign n7933 = n7932 ^ n2348 ;
  assign n7930 = n5777 & n5788 ;
  assign n7928 = n5777 & n5781 ;
  assign n7929 = n7928 ^ n5777 ;
  assign n7931 = n7930 ^ n7929 ;
  assign n7934 = n7933 ^ n7931 ;
  assign n7925 = n2748 & ~n3611 ;
  assign n7926 = n7925 ^ n2748 ;
  assign n7924 = n5803 ^ n5800 ;
  assign n7927 = n7926 ^ n7924 ;
  assign n7935 = n7934 ^ n7927 ;
  assign n7941 = n5817 & n5828 ;
  assign n7942 = n7941 ^ n5828 ;
  assign n7936 = n5850 ^ n5847 ;
  assign n7937 = n5841 & ~n7936 ;
  assign n7938 = n7937 ^ n5841 ;
  assign n7939 = n7938 ^ n5841 ;
  assign n7940 = n7939 ^ n7936 ;
  assign n7943 = n7942 ^ n7940 ;
  assign n7952 = n2348 & ~n3957 ;
  assign n7953 = n7952 ^ n2348 ;
  assign n7949 = n5884 & n5888 ;
  assign n7950 = n7949 ^ n5884 ;
  assign n7948 = n5884 & n5895 ;
  assign n7951 = n7950 ^ n7948 ;
  assign n7954 = n7953 ^ n7951 ;
  assign n7945 = n2748 & ~n3937 ;
  assign n7946 = n7945 ^ n2748 ;
  assign n7944 = n5910 ^ n5907 ;
  assign n7947 = n7946 ^ n7944 ;
  assign n7955 = n7954 ^ n7947 ;
  assign n7984 = n5955 ^ n399 ;
  assign n7985 = n7984 ^ x134 ;
  assign n7972 = n5925 ^ n399 ;
  assign n7973 = n7972 ^ x134 ;
  assign n7976 = n7813 ^ n5411 ;
  assign n7974 = n5925 ^ n137 ;
  assign n7975 = n7974 ^ x134 ;
  assign n7977 = n7976 ^ n7975 ;
  assign n7978 = n7977 ^ n3612 ;
  assign n7979 = n7978 ^ n5925 ;
  assign n7980 = n7973 & n7979 ;
  assign n7981 = n7980 ^ n7973 ;
  assign n7982 = n7981 ^ n7977 ;
  assign n7983 = n7982 ^ n3612 ;
  assign n7986 = n7985 ^ n7983 ;
  assign n7958 = n402 ^ n308 ;
  assign n7959 = n7958 ^ n5967 ;
  assign n7960 = n7959 ^ n5981 ;
  assign n7956 = n6007 ^ n5983 ;
  assign n7961 = n7960 ^ n7956 ;
  assign n7962 = n7961 ^ n5967 ;
  assign n7963 = n7962 ^ n5961 ;
  assign n7964 = n7956 ^ n308 ;
  assign n7965 = n7964 ^ x134 ;
  assign n7966 = n7963 & n7965 ;
  assign n7967 = n7966 ^ n7963 ;
  assign n7968 = n7967 ^ n7965 ;
  assign n7969 = n7968 ^ n7960 ;
  assign n7957 = n7956 ^ n5966 ;
  assign n7970 = n7969 ^ n7957 ;
  assign n7971 = n7970 ^ n5959 ;
  assign n7987 = n7986 ^ n7971 ;
  assign n7996 = ~n930 & n2348 ;
  assign n7997 = n7996 ^ n2348 ;
  assign n7993 = n6046 & n6050 ;
  assign n7994 = n7993 ^ n6046 ;
  assign n7992 = n6046 & n6055 ;
  assign n7995 = n7994 ^ n7992 ;
  assign n7998 = n7997 ^ n7995 ;
  assign n7989 = ~n1174 & n2748 ;
  assign n7990 = n7989 ^ n2748 ;
  assign n7988 = n6070 ^ n6067 ;
  assign n7991 = n7990 ^ n7988 ;
  assign n7999 = n7998 ^ n7991 ;
  assign n8005 = n6090 & n6104 ;
  assign n8006 = n8005 ^ n6104 ;
  assign n8007 = n8006 ^ n6104 ;
  assign n8000 = n6133 ^ n6130 ;
  assign n8001 = n6124 & ~n8000 ;
  assign n8002 = n8001 ^ n6124 ;
  assign n8003 = n8002 ^ n6124 ;
  assign n8004 = n8003 ^ n8000 ;
  assign n8008 = n8007 ^ n8004 ;
  assign n8017 = ~n1715 & n4441 ;
  assign n8018 = n8017 ^ n4441 ;
  assign n8014 = n6161 & n6165 ;
  assign n8015 = n8014 ^ n6161 ;
  assign n8013 = n6161 & n6170 ;
  assign n8016 = n8015 ^ n8013 ;
  assign n8019 = n8018 ^ n8016 ;
  assign n8010 = n2748 & ~n4206 ;
  assign n8011 = n8010 ^ n2748 ;
  assign n8009 = n6183 ^ n6181 ;
  assign n8012 = n8011 ^ n8009 ;
  assign n8020 = n8019 ^ n8012 ;
  assign n8044 = n6200 ^ n6198 ;
  assign n8045 = n6190 & n8044 ;
  assign n8046 = n8045 ^ n6190 ;
  assign n8037 = x134 & n6217 ;
  assign n8038 = n8037 ^ x134 ;
  assign n8041 = n402 & n2133 ;
  assign n8042 = n8038 & n8041 ;
  assign n8039 = n6288 & n8038 ;
  assign n8040 = n8039 ^ n8038 ;
  assign n8043 = n8042 ^ n8040 ;
  assign n8047 = n8046 ^ n8043 ;
  assign n8023 = n2052 ^ n402 ;
  assign n8024 = n8023 ^ n6229 ;
  assign n8025 = n8024 ^ n6243 ;
  assign n8021 = n6268 ^ n6245 ;
  assign n8026 = n8025 ^ n8021 ;
  assign n8027 = n8026 ^ n6229 ;
  assign n8028 = n8027 ^ n6223 ;
  assign n8029 = n8021 ^ n2052 ;
  assign n8030 = n8029 ^ x134 ;
  assign n8031 = n8028 & n8030 ;
  assign n8032 = n8031 ^ n8028 ;
  assign n8033 = n8032 ^ n8030 ;
  assign n8034 = n8033 ^ n8025 ;
  assign n8022 = n8021 ^ n6228 ;
  assign n8035 = n8034 ^ n8022 ;
  assign n8036 = n8035 ^ n6221 ;
  assign n8048 = n8047 ^ n8036 ;
  assign n8057 = ~n2366 & n5411 ;
  assign n8058 = n8057 ^ n5411 ;
  assign n8055 = n6331 & n6341 ;
  assign n8053 = n6331 & n6335 ;
  assign n8054 = n8053 ^ n6331 ;
  assign n8056 = n8055 ^ n8054 ;
  assign n8059 = n8058 ^ n8056 ;
  assign n8050 = ~n2222 & n2348 ;
  assign n8051 = n8050 ^ n2348 ;
  assign n8049 = n6355 ^ n6352 ;
  assign n8052 = n8051 ^ n8049 ;
  assign n8060 = n8059 ^ n8052 ;
  assign n8068 = n6371 & n6382 ;
  assign n8069 = n8068 ^ n6382 ;
  assign n8070 = n8069 ^ n6382 ;
  assign n8065 = n2467 & n2748 ;
  assign n8066 = ~n6394 & n8065 ;
  assign n8061 = n2390 & n4441 ;
  assign n8062 = n8061 ^ x134 ;
  assign n8063 = n6394 & ~n8062 ;
  assign n8064 = n8063 ^ n8062 ;
  assign n8067 = n8066 ^ n8064 ;
  assign n8071 = n8070 ^ n8067 ;
  assign n8088 = n2348 & ~n2570 ;
  assign n8089 = n8088 ^ n2348 ;
  assign n8085 = n6426 & n6430 ;
  assign n8086 = n8085 ^ n6426 ;
  assign n8084 = n6426 & n6436 ;
  assign n8087 = n8086 ^ n8084 ;
  assign n8090 = n8089 ^ n8087 ;
  assign n8078 = n6466 ^ n6458 ;
  assign n8079 = ~n6447 & n8078 ;
  assign n8080 = n8079 ^ n6447 ;
  assign n8081 = n8080 ^ n8078 ;
  assign n8082 = n8081 ^ n8078 ;
  assign n8072 = n850 & n6458 ;
  assign n8073 = n8072 ^ n850 ;
  assign n8074 = n8073 ^ n850 ;
  assign n8075 = ~n6447 & n8074 ;
  assign n8076 = n8075 ^ n8074 ;
  assign n8077 = n8076 ^ n8074 ;
  assign n8083 = n8082 ^ n8077 ;
  assign n8091 = n8090 ^ n8083 ;
  assign n8096 = n1259 & n2758 ;
  assign n8097 = n6480 & n8096 ;
  assign n8098 = n8097 ^ n8096 ;
  assign n8099 = n8098 ^ n6520 ;
  assign n8092 = n6523 ^ n6480 ;
  assign n8093 = n6525 & n8092 ;
  assign n8094 = n8093 ^ n6525 ;
  assign n8095 = n8094 ^ n8092 ;
  assign n8100 = n8099 ^ n8095 ;
  assign n8113 = n2348 & ~n2915 ;
  assign n8114 = n8113 ^ n2348 ;
  assign n8115 = n8114 ^ n6579 ;
  assign n8107 = n6607 ^ n6599 ;
  assign n8108 = ~n6588 & n8107 ;
  assign n8109 = n8108 ^ n6588 ;
  assign n8110 = n8109 ^ n8107 ;
  assign n8111 = n8110 ^ n8107 ;
  assign n8101 = n850 & n6599 ;
  assign n8102 = n8101 ^ n850 ;
  assign n8103 = n8102 ^ n850 ;
  assign n8104 = ~n6588 & n8103 ;
  assign n8105 = n8104 ^ n8103 ;
  assign n8106 = n8105 ^ n8103 ;
  assign n8112 = n8111 ^ n8106 ;
  assign n8116 = n8115 ^ n8112 ;
  assign n8119 = n6621 & n6632 ;
  assign n8120 = n8119 ^ n6632 ;
  assign n8121 = n8120 ^ n6632 ;
  assign n8117 = ~x134 & ~n6651 ;
  assign n8118 = ~n6640 & n8117 ;
  assign n8122 = n8121 ^ n8118 ;
  assign n8137 = n2348 & ~n3235 ;
  assign n8138 = n8137 ^ n2348 ;
  assign n8134 = n6685 & n6689 ;
  assign n8135 = n8134 ^ n6685 ;
  assign n8133 = n6685 & n6694 ;
  assign n8136 = n8135 ^ n8133 ;
  assign n8139 = n8138 ^ n8136 ;
  assign n8127 = n6721 ^ n6715 ;
  assign n8128 = ~n6706 & n8127 ;
  assign n8129 = n8128 ^ n6706 ;
  assign n8130 = n8129 ^ n8127 ;
  assign n8131 = n8130 ^ n8127 ;
  assign n8123 = n850 & n6715 ;
  assign n8124 = ~n6706 & n8123 ;
  assign n8125 = n8124 ^ n8123 ;
  assign n8126 = n8125 ^ n8123 ;
  assign n8132 = n8131 ^ n8126 ;
  assign n8140 = n8139 ^ n8132 ;
  assign n8164 = n3479 ^ n138 ;
  assign n8165 = n4441 ^ n3479 ;
  assign n8166 = ~n8164 & n8165 ;
  assign n8167 = n8166 ^ n6752 ;
  assign n8168 = n8167 ^ n8164 ;
  assign n8170 = n6752 ^ n138 ;
  assign n8169 = n4441 ^ x134 ;
  assign n8171 = n8170 ^ n8169 ;
  assign n8172 = ~n8168 & n8171 ;
  assign n8173 = n8172 ^ n4441 ;
  assign n8158 = n1259 & n3408 ;
  assign n8159 = n6735 & n8158 ;
  assign n8160 = n8159 ^ n8158 ;
  assign n8161 = n8160 ^ n3378 ;
  assign n8162 = n8161 ^ n136 ;
  assign n8146 = n6752 ^ n136 ;
  assign n8147 = n8146 ^ x134 ;
  assign n8148 = n850 ^ n136 ;
  assign n8149 = n8148 ^ x134 ;
  assign n8150 = n3378 ^ x134 ;
  assign n8151 = n8149 & n8150 ;
  assign n8152 = n8151 ^ n850 ;
  assign n8153 = n8152 ^ n6752 ;
  assign n8154 = n8153 ^ n8150 ;
  assign n8155 = n8147 & n8154 ;
  assign n8156 = n8155 ^ n8151 ;
  assign n8157 = n8156 ^ n850 ;
  assign n8163 = n8162 ^ n8157 ;
  assign n8174 = n8173 ^ n8163 ;
  assign n8145 = n138 ^ x134 ;
  assign n8175 = n8174 ^ n8145 ;
  assign n8141 = n6767 ^ n6735 ;
  assign n8142 = n6769 & n8141 ;
  assign n8143 = n8142 ^ n6769 ;
  assign n8144 = n8143 ^ n8141 ;
  assign n8176 = n8175 ^ n8144 ;
  assign n8195 = n2748 & n3633 ;
  assign n8196 = n8195 ^ n2748 ;
  assign n8197 = n8196 ^ n2748 ;
  assign n8198 = ~n6781 & n8197 ;
  assign n8199 = n8198 ^ n8197 ;
  assign n8200 = n8199 ^ n8197 ;
  assign n8194 = n6788 ^ n6781 ;
  assign n8201 = n8200 ^ n8194 ;
  assign n8189 = n1259 & n3558 ;
  assign n8190 = ~n6781 & n8189 ;
  assign n8191 = n8190 ^ n8189 ;
  assign n8192 = n8191 ^ n8189 ;
  assign n8183 = n1180 & n3526 ;
  assign n8184 = n8183 ^ n1180 ;
  assign n8185 = n8184 ^ n1180 ;
  assign n8186 = n6799 & n8185 ;
  assign n8187 = n8186 ^ n8185 ;
  assign n8177 = n1175 & n3611 ;
  assign n8178 = n8177 ^ n1175 ;
  assign n8179 = n8178 ^ n1175 ;
  assign n8180 = n6799 & n8179 ;
  assign n8181 = n8180 ^ n8179 ;
  assign n8182 = n8181 ^ n6801 ;
  assign n8188 = n8187 ^ n8182 ;
  assign n8193 = n8192 ^ n8188 ;
  assign n8202 = n8201 ^ n8193 ;
  assign n8210 = n6872 ^ n6870 ;
  assign n8211 = n8210 ^ x134 ;
  assign n8212 = n6844 & n8211 ;
  assign n8213 = n8212 ^ n8211 ;
  assign n8214 = n8213 ^ n6844 ;
  assign n8215 = n8214 ^ n8210 ;
  assign n8216 = n8215 ^ n6843 ;
  assign n8207 = n1259 & n3710 ;
  assign n8208 = n6885 & n8207 ;
  assign n8203 = n2748 & n3742 ;
  assign n8204 = n8203 ^ x134 ;
  assign n8205 = ~n6885 & ~n8204 ;
  assign n8206 = n8205 ^ n8204 ;
  assign n8209 = n8208 ^ n8206 ;
  assign n8217 = n8216 ^ n8209 ;
  assign n8238 = n2748 & n3957 ;
  assign n8239 = n8238 ^ n2748 ;
  assign n8240 = n8239 ^ n2748 ;
  assign n8241 = ~n6901 & n8240 ;
  assign n8242 = n8241 ^ n8240 ;
  assign n8243 = n8242 ^ n8240 ;
  assign n8231 = n1259 & n3877 ;
  assign n8232 = n8231 ^ n1259 ;
  assign n8233 = n8232 ^ n1259 ;
  assign n8234 = ~n6901 & n8233 ;
  assign n8235 = n8234 ^ n8233 ;
  assign n8236 = n8235 ^ n8233 ;
  assign n8225 = n1180 & n3845 ;
  assign n8226 = n8225 ^ n1180 ;
  assign n8227 = n8226 ^ n1180 ;
  assign n8228 = n6927 & n8227 ;
  assign n8229 = n8228 ^ n8227 ;
  assign n8219 = n1175 & n3937 ;
  assign n8220 = n8219 ^ n1175 ;
  assign n8221 = n8220 ^ n1175 ;
  assign n8222 = n6927 & n8221 ;
  assign n8223 = n8222 ^ n8221 ;
  assign n8224 = n8223 ^ n6929 ;
  assign n8230 = n8229 ^ n8224 ;
  assign n8237 = n8236 ^ n8230 ;
  assign n8244 = n8243 ^ n8237 ;
  assign n8218 = n6910 ^ n6901 ;
  assign n8245 = n8244 ^ n8218 ;
  assign y0 = n683 ;
  assign y1 = n1338 ;
  assign y2 = ~n1572 ;
  assign y3 = n2007 ;
  assign y4 = n2155 ;
  assign y5 = n2370 ;
  assign y6 = ~n2503 ;
  assign y7 = n2716 ;
  assign y8 = ~n2852 ;
  assign y9 = n3046 ;
  assign y10 = n3172 ;
  assign y11 = n3366 ;
  assign y12 = n3516 ;
  assign y13 = n3663 ;
  assign y14 = n3835 ;
  assign y15 = n3991 ;
  assign y16 = n4049 ;
  assign y17 = n4093 ;
  assign y18 = n4160 ;
  assign y19 = n4223 ;
  assign y20 = n4277 ;
  assign y21 = n4340 ;
  assign y22 = ~n4388 ;
  assign y23 = n4445 ;
  assign y24 = n4522 ;
  assign y25 = n4612 ;
  assign y26 = n4686 ;
  assign y27 = n4749 ;
  assign y28 = n4813 ;
  assign y29 = n4876 ;
  assign y30 = ~n4924 ;
  assign y31 = n4989 ;
  assign y32 = ~n5056 ;
  assign y33 = n5115 ;
  assign y34 = n5173 ;
  assign y35 = n5218 ;
  assign y36 = n5288 ;
  assign y37 = n5347 ;
  assign y38 = n5399 ;
  assign y39 = ~n5459 ;
  assign y40 = n5516 ;
  assign y41 = ~n5586 ;
  assign y42 = n5647 ;
  assign y43 = ~n5709 ;
  assign y44 = n5758 ;
  assign y45 = ~n5808 ;
  assign y46 = n5853 ;
  assign y47 = ~n5915 ;
  assign y48 = n6025 ;
  assign y49 = n6075 ;
  assign y50 = ~n6136 ;
  assign y51 = n6188 ;
  assign y52 = ~n6306 ;
  assign y53 = n6360 ;
  assign y54 = ~n6402 ;
  assign y55 = n6472 ;
  assign y56 = n6529 ;
  assign y57 = n6613 ;
  assign y58 = ~n6654 ;
  assign y59 = ~n6727 ;
  assign y60 = ~n6773 ;
  assign y61 = n6823 ;
  assign y62 = n6893 ;
  assign y63 = n6951 ;
  assign y64 = n6967 ;
  assign y65 = n7003 ;
  assign y66 = ~n7005 ;
  assign y67 = n7048 ;
  assign y68 = n7066 ;
  assign y69 = n7101 ;
  assign y70 = n7106 ;
  assign y71 = n7145 ;
  assign y72 = ~n7169 ;
  assign y73 = n7198 ;
  assign y74 = n7205 ;
  assign y75 = ~n7247 ;
  assign y76 = n7261 ;
  assign y77 = n7293 ;
  assign y78 = ~n7302 ;
  assign y79 = n7336 ;
  assign y80 = n7363 ;
  assign y81 = n7386 ;
  assign y82 = ~n7395 ;
  assign y83 = n7416 ;
  assign y84 = ~n7434 ;
  assign y85 = ~n7460 ;
  assign y86 = ~n7469 ;
  assign y87 = n7487 ;
  assign y88 = n7525 ;
  assign y89 = n7536 ;
  assign y90 = ~n7544 ;
  assign y91 = n7582 ;
  assign y92 = ~n7617 ;
  assign y93 = n7645 ;
  assign y94 = n7653 ;
  assign y95 = n7681 ;
  assign y96 = n7702 ;
  assign y97 = n7728 ;
  assign y98 = n7735 ;
  assign y99 = n7755 ;
  assign y100 = ~n7777 ;
  assign y101 = n7804 ;
  assign y102 = n7808 ;
  assign y103 = n7837 ;
  assign y104 = n7859 ;
  assign y105 = n7875 ;
  assign y106 = ~n7884 ;
  assign y107 = n7917 ;
  assign y108 = n7923 ;
  assign y109 = n7935 ;
  assign y110 = n7943 ;
  assign y111 = n7955 ;
  assign y112 = ~n7987 ;
  assign y113 = n7999 ;
  assign y114 = n8008 ;
  assign y115 = n8020 ;
  assign y116 = ~n8048 ;
  assign y117 = n8060 ;
  assign y118 = n8071 ;
  assign y119 = n8091 ;
  assign y120 = n8100 ;
  assign y121 = n8116 ;
  assign y122 = ~n8122 ;
  assign y123 = n8140 ;
  assign y124 = n8176 ;
  assign y125 = n8202 ;
  assign y126 = n8217 ;
  assign y127 = n8245 ;
endmodule
