module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 ;
  assign n462 = x40 ^ x16 ;
  assign n466 = x41 ^ x17 ;
  assign n467 = ~n462 & ~n466 ;
  assign n469 = x42 ^ x18 ;
  assign n475 = x43 ^ x19 ;
  assign n476 = ~n469 & ~n475 ;
  assign n477 = n467 & n476 ;
  assign n479 = x44 ^ x20 ;
  assign n483 = x45 ^ x21 ;
  assign n484 = ~n479 & ~n483 ;
  assign n486 = x46 ^ x22 ;
  assign n496 = x47 ^ x23 ;
  assign n497 = ~n486 & ~n496 ;
  assign n498 = n484 & n497 ;
  assign n499 = n477 & n498 ;
  assign n487 = x23 & x47 ;
  assign n488 = n487 ^ x23 ;
  assign n489 = n486 & n488 ;
  assign n490 = n489 ^ n488 ;
  assign n485 = x22 & ~x46 ;
  assign n491 = n490 ^ n485 ;
  assign n492 = n484 & n491 ;
  assign n480 = x21 & ~x45 ;
  assign n481 = ~n479 & n480 ;
  assign n478 = x20 & ~x44 ;
  assign n482 = n481 ^ n478 ;
  assign n493 = n492 ^ n482 ;
  assign n494 = n477 & n493 ;
  assign n470 = x19 & ~x43 ;
  assign n471 = ~n469 & n470 ;
  assign n468 = x18 & ~x42 ;
  assign n472 = n471 ^ n468 ;
  assign n473 = n467 & n472 ;
  assign n463 = x17 & ~x41 ;
  assign n464 = ~n462 & n463 ;
  assign n461 = x16 & ~x40 ;
  assign n465 = n464 ^ n461 ;
  assign n474 = n473 ^ n465 ;
  assign n495 = n494 ^ n474 ;
  assign n500 = n499 ^ n495 ;
  assign n275 = x40 ^ x8 ;
  assign n279 = x41 ^ x9 ;
  assign n280 = ~n275 & ~n279 ;
  assign n282 = x42 ^ x10 ;
  assign n288 = x43 ^ x11 ;
  assign n289 = ~n282 & ~n288 ;
  assign n290 = n280 & n289 ;
  assign n292 = x44 ^ x12 ;
  assign n296 = x45 ^ x13 ;
  assign n297 = ~n292 & ~n296 ;
  assign n299 = x46 ^ x14 ;
  assign n309 = x47 ^ x15 ;
  assign n310 = ~n299 & ~n309 ;
  assign n311 = n297 & n310 ;
  assign n312 = n290 & n311 ;
  assign n300 = x15 & x47 ;
  assign n301 = n300 ^ x15 ;
  assign n302 = n299 & n301 ;
  assign n303 = n302 ^ n301 ;
  assign n298 = x14 & ~x46 ;
  assign n304 = n303 ^ n298 ;
  assign n305 = n297 & n304 ;
  assign n293 = x13 & ~x45 ;
  assign n294 = ~n292 & n293 ;
  assign n291 = x12 & ~x44 ;
  assign n295 = n294 ^ n291 ;
  assign n306 = n305 ^ n295 ;
  assign n307 = n290 & n306 ;
  assign n283 = x11 & ~x43 ;
  assign n284 = ~n282 & n283 ;
  assign n281 = x10 & ~x42 ;
  assign n285 = n284 ^ n281 ;
  assign n286 = n280 & n285 ;
  assign n276 = x9 & ~x41 ;
  assign n277 = ~n275 & n276 ;
  assign n274 = x8 & ~x40 ;
  assign n278 = n277 ^ n274 ;
  assign n287 = n286 ^ n278 ;
  assign n308 = n307 ^ n287 ;
  assign n313 = n312 ^ n308 ;
  assign n793 = n500 ^ n313 ;
  assign n50 = x40 ^ x0 ;
  assign n54 = x41 ^ x1 ;
  assign n55 = ~n50 & ~n54 ;
  assign n57 = x42 ^ x2 ;
  assign n63 = x43 ^ x3 ;
  assign n64 = ~n57 & ~n63 ;
  assign n65 = n55 & n64 ;
  assign n67 = x44 ^ x4 ;
  assign n71 = x45 ^ x5 ;
  assign n72 = ~n67 & ~n71 ;
  assign n74 = x46 ^ x6 ;
  assign n84 = x47 ^ x7 ;
  assign n85 = ~n74 & ~n84 ;
  assign n86 = n72 & n85 ;
  assign n87 = n65 & n86 ;
  assign n75 = x7 & x47 ;
  assign n76 = n75 ^ x7 ;
  assign n77 = n74 & n76 ;
  assign n78 = n77 ^ n76 ;
  assign n73 = x6 & ~x46 ;
  assign n79 = n78 ^ n73 ;
  assign n80 = n72 & n79 ;
  assign n68 = x5 & ~x45 ;
  assign n69 = ~n67 & n68 ;
  assign n66 = x4 & ~x44 ;
  assign n70 = n69 ^ n66 ;
  assign n81 = n80 ^ n70 ;
  assign n82 = n65 & n81 ;
  assign n58 = x3 & ~x43 ;
  assign n59 = ~n57 & n58 ;
  assign n56 = x2 & ~x42 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n55 & n60 ;
  assign n51 = x1 & ~x41 ;
  assign n52 = ~n50 & n51 ;
  assign n49 = x0 & ~x40 ;
  assign n53 = n52 ^ n49 ;
  assign n62 = n61 ^ n53 ;
  assign n83 = n82 ^ n62 ;
  assign n88 = n87 ^ n83 ;
  assign n801 = n793 ^ n88 ;
  assign n731 = x40 ^ x32 ;
  assign n735 = x41 ^ x33 ;
  assign n736 = ~n731 & ~n735 ;
  assign n738 = x42 ^ x34 ;
  assign n744 = x43 ^ x35 ;
  assign n745 = ~n738 & ~n744 ;
  assign n746 = n736 & n745 ;
  assign n748 = x44 ^ x36 ;
  assign n752 = x45 ^ x37 ;
  assign n753 = ~n748 & ~n752 ;
  assign n755 = x46 ^ x38 ;
  assign n765 = x47 ^ x39 ;
  assign n766 = ~n755 & ~n765 ;
  assign n767 = n753 & n766 ;
  assign n768 = n746 & n767 ;
  assign n756 = x39 & x47 ;
  assign n757 = n756 ^ x39 ;
  assign n758 = n755 & n757 ;
  assign n759 = n758 ^ n757 ;
  assign n754 = x38 & ~x46 ;
  assign n760 = n759 ^ n754 ;
  assign n761 = n753 & n760 ;
  assign n749 = x37 & ~x45 ;
  assign n750 = ~n748 & n749 ;
  assign n747 = x36 & ~x44 ;
  assign n751 = n750 ^ n747 ;
  assign n762 = n761 ^ n751 ;
  assign n763 = n746 & n762 ;
  assign n739 = x35 & ~x43 ;
  assign n740 = ~n738 & n739 ;
  assign n737 = x34 & ~x42 ;
  assign n741 = n740 ^ n737 ;
  assign n742 = n736 & n741 ;
  assign n732 = x33 & ~x41 ;
  assign n733 = ~n731 & n732 ;
  assign n730 = x32 & ~x40 ;
  assign n734 = n733 ^ n730 ;
  assign n743 = n742 ^ n734 ;
  assign n764 = n763 ^ n743 ;
  assign n769 = n768 ^ n764 ;
  assign n661 = x40 ^ x24 ;
  assign n665 = x41 ^ x25 ;
  assign n666 = ~n661 & ~n665 ;
  assign n668 = x42 ^ x26 ;
  assign n674 = x43 ^ x27 ;
  assign n675 = ~n668 & ~n674 ;
  assign n676 = n666 & n675 ;
  assign n678 = x44 ^ x28 ;
  assign n682 = x45 ^ x29 ;
  assign n683 = ~n678 & ~n682 ;
  assign n685 = x46 ^ x30 ;
  assign n695 = x47 ^ x31 ;
  assign n696 = ~n685 & ~n695 ;
  assign n697 = n683 & n696 ;
  assign n698 = n676 & n697 ;
  assign n686 = x31 & x47 ;
  assign n687 = n686 ^ x31 ;
  assign n688 = n685 & n687 ;
  assign n689 = n688 ^ n687 ;
  assign n684 = x30 & ~x46 ;
  assign n690 = n689 ^ n684 ;
  assign n691 = n683 & n690 ;
  assign n679 = x29 & ~x45 ;
  assign n680 = ~n678 & n679 ;
  assign n677 = x28 & ~x44 ;
  assign n681 = n680 ^ n677 ;
  assign n692 = n691 ^ n681 ;
  assign n693 = n676 & n692 ;
  assign n669 = x27 & ~x43 ;
  assign n670 = ~n668 & n669 ;
  assign n667 = x26 & ~x42 ;
  assign n671 = n670 ^ n667 ;
  assign n672 = n666 & n671 ;
  assign n662 = x25 & ~x41 ;
  assign n663 = ~n661 & n662 ;
  assign n660 = x24 & ~x40 ;
  assign n664 = n663 ^ n660 ;
  assign n673 = n672 ^ n664 ;
  assign n694 = n693 ^ n673 ;
  assign n699 = n698 ^ n694 ;
  assign n802 = n769 ^ n699 ;
  assign n803 = n801 & n802 ;
  assign n804 = n803 ^ n802 ;
  assign n797 = n313 & n500 ;
  assign n798 = n797 ^ n500 ;
  assign n799 = n798 ^ n313 ;
  assign n794 = n88 & n793 ;
  assign n795 = n794 ^ n793 ;
  assign n800 = n799 ^ n795 ;
  assign n805 = n804 ^ n800 ;
  assign n806 = n699 & n769 ;
  assign n807 = n806 ^ n769 ;
  assign n808 = n807 ^ n699 ;
  assign n809 = n808 ^ n804 ;
  assign n810 = ~n805 & ~n809 ;
  assign n811 = n810 ^ n804 ;
  assign n791 = ~n88 & ~n313 ;
  assign n790 = ~n88 & ~n500 ;
  assign n792 = n791 ^ n790 ;
  assign n796 = n795 ^ n792 ;
  assign n812 = n811 ^ n796 ;
  assign n813 = n808 ^ n805 ;
  assign n814 = n802 ^ n801 ;
  assign n815 = x40 & n814 ;
  assign n816 = n813 & n815 ;
  assign n817 = n816 ^ n815 ;
  assign n818 = n812 & n817 ;
  assign n819 = n818 ^ n817 ;
  assign n543 = x32 ^ x16 ;
  assign n547 = x33 ^ x17 ;
  assign n548 = ~n543 & ~n547 ;
  assign n550 = x34 ^ x18 ;
  assign n556 = x35 ^ x19 ;
  assign n557 = ~n550 & ~n556 ;
  assign n558 = n548 & n557 ;
  assign n560 = x36 ^ x20 ;
  assign n564 = x37 ^ x21 ;
  assign n565 = ~n560 & ~n564 ;
  assign n567 = x38 ^ x22 ;
  assign n577 = x39 ^ x23 ;
  assign n578 = ~n567 & ~n577 ;
  assign n579 = n565 & n578 ;
  assign n580 = n558 & n579 ;
  assign n568 = x23 & x39 ;
  assign n569 = n568 ^ x23 ;
  assign n570 = n567 & n569 ;
  assign n571 = n570 ^ n569 ;
  assign n566 = x22 & ~x38 ;
  assign n572 = n571 ^ n566 ;
  assign n573 = n565 & n572 ;
  assign n561 = x21 & ~x37 ;
  assign n562 = ~n560 & n561 ;
  assign n559 = x20 & ~x36 ;
  assign n563 = n562 ^ n559 ;
  assign n574 = n573 ^ n563 ;
  assign n575 = n558 & n574 ;
  assign n551 = x19 & ~x35 ;
  assign n552 = ~n550 & n551 ;
  assign n549 = x18 & ~x34 ;
  assign n553 = n552 ^ n549 ;
  assign n554 = n548 & n553 ;
  assign n544 = x17 & ~x33 ;
  assign n545 = ~n543 & n544 ;
  assign n542 = x16 & ~x32 ;
  assign n546 = n545 ^ n542 ;
  assign n555 = n554 ^ n546 ;
  assign n576 = n575 ^ n555 ;
  assign n581 = n580 ^ n576 ;
  assign n356 = x32 ^ x8 ;
  assign n360 = x33 ^ x9 ;
  assign n361 = ~n356 & ~n360 ;
  assign n363 = x34 ^ x10 ;
  assign n369 = x35 ^ x11 ;
  assign n370 = ~n363 & ~n369 ;
  assign n371 = n361 & n370 ;
  assign n373 = x36 ^ x12 ;
  assign n377 = x37 ^ x13 ;
  assign n378 = ~n373 & ~n377 ;
  assign n380 = x38 ^ x14 ;
  assign n390 = x39 ^ x15 ;
  assign n391 = ~n380 & ~n390 ;
  assign n392 = n378 & n391 ;
  assign n393 = n371 & n392 ;
  assign n381 = x15 & x39 ;
  assign n382 = n381 ^ x15 ;
  assign n383 = n380 & n382 ;
  assign n384 = n383 ^ n382 ;
  assign n379 = x14 & ~x38 ;
  assign n385 = n384 ^ n379 ;
  assign n386 = n378 & n385 ;
  assign n374 = x13 & ~x37 ;
  assign n375 = ~n373 & n374 ;
  assign n372 = x12 & ~x36 ;
  assign n376 = n375 ^ n372 ;
  assign n387 = n386 ^ n376 ;
  assign n388 = n371 & n387 ;
  assign n364 = x11 & ~x35 ;
  assign n365 = ~n363 & n364 ;
  assign n362 = x10 & ~x34 ;
  assign n366 = n365 ^ n362 ;
  assign n367 = n361 & n366 ;
  assign n357 = x9 & ~x33 ;
  assign n358 = ~n356 & n357 ;
  assign n355 = x8 & ~x32 ;
  assign n359 = n358 ^ n355 ;
  assign n368 = n367 ^ n359 ;
  assign n389 = n388 ^ n368 ;
  assign n394 = n393 ^ n389 ;
  assign n721 = n581 ^ n394 ;
  assign n131 = x32 ^ x0 ;
  assign n135 = x33 ^ x1 ;
  assign n136 = ~n131 & ~n135 ;
  assign n138 = x34 ^ x2 ;
  assign n144 = x35 ^ x3 ;
  assign n145 = ~n138 & ~n144 ;
  assign n146 = n136 & n145 ;
  assign n148 = x36 ^ x4 ;
  assign n152 = x37 ^ x5 ;
  assign n153 = ~n148 & ~n152 ;
  assign n155 = x38 ^ x6 ;
  assign n165 = x39 ^ x7 ;
  assign n166 = ~n155 & ~n165 ;
  assign n167 = n153 & n166 ;
  assign n168 = n146 & n167 ;
  assign n156 = x7 & x39 ;
  assign n157 = n156 ^ x7 ;
  assign n158 = n155 & n157 ;
  assign n159 = n158 ^ n157 ;
  assign n154 = x6 & ~x38 ;
  assign n160 = n159 ^ n154 ;
  assign n161 = n153 & n160 ;
  assign n149 = x5 & ~x37 ;
  assign n150 = ~n148 & n149 ;
  assign n147 = x4 & ~x36 ;
  assign n151 = n150 ^ n147 ;
  assign n162 = n161 ^ n151 ;
  assign n163 = n146 & n162 ;
  assign n139 = x3 & ~x35 ;
  assign n140 = ~n138 & n139 ;
  assign n137 = x2 & ~x34 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n136 & n141 ;
  assign n132 = x1 & ~x33 ;
  assign n133 = ~n131 & n132 ;
  assign n130 = x0 & ~x32 ;
  assign n134 = n133 ^ n130 ;
  assign n143 = n142 ^ n134 ;
  assign n164 = n163 ^ n143 ;
  assign n169 = n168 ^ n164 ;
  assign n729 = n721 ^ n169 ;
  assign n621 = x32 ^ x24 ;
  assign n625 = x33 ^ x25 ;
  assign n626 = ~n621 & ~n625 ;
  assign n628 = x34 ^ x26 ;
  assign n634 = x35 ^ x27 ;
  assign n635 = ~n628 & ~n634 ;
  assign n636 = n626 & n635 ;
  assign n638 = x36 ^ x28 ;
  assign n642 = x37 ^ x29 ;
  assign n643 = ~n638 & ~n642 ;
  assign n645 = x38 ^ x30 ;
  assign n655 = x39 ^ x31 ;
  assign n656 = ~n645 & ~n655 ;
  assign n657 = n643 & n656 ;
  assign n658 = n636 & n657 ;
  assign n646 = x31 & x39 ;
  assign n647 = n646 ^ x31 ;
  assign n648 = n645 & n647 ;
  assign n649 = n648 ^ n647 ;
  assign n644 = x30 & ~x38 ;
  assign n650 = n649 ^ n644 ;
  assign n651 = n643 & n650 ;
  assign n639 = x29 & ~x37 ;
  assign n640 = ~n638 & n639 ;
  assign n637 = x28 & ~x36 ;
  assign n641 = n640 ^ n637 ;
  assign n652 = n651 ^ n641 ;
  assign n653 = n636 & n652 ;
  assign n629 = x27 & ~x35 ;
  assign n630 = ~n628 & n629 ;
  assign n627 = x26 & ~x34 ;
  assign n631 = n630 ^ n627 ;
  assign n632 = n626 & n631 ;
  assign n622 = x25 & ~x33 ;
  assign n623 = ~n621 & n622 ;
  assign n620 = x24 & ~x32 ;
  assign n624 = n623 ^ n620 ;
  assign n633 = n632 ^ n624 ;
  assign n654 = n653 ^ n633 ;
  assign n659 = n658 ^ n654 ;
  assign n770 = n769 ^ n659 ;
  assign n771 = n729 & n770 ;
  assign n772 = n771 ^ n729 ;
  assign n773 = n772 ^ n770 ;
  assign n725 = n394 & n581 ;
  assign n726 = n725 ^ n581 ;
  assign n727 = n726 ^ n394 ;
  assign n722 = n169 & n721 ;
  assign n723 = n722 ^ n721 ;
  assign n728 = n727 ^ n723 ;
  assign n774 = n773 ^ n728 ;
  assign n775 = n659 & n769 ;
  assign n776 = n775 ^ n769 ;
  assign n777 = n776 ^ n773 ;
  assign n778 = n774 & ~n777 ;
  assign n779 = n778 ^ n773 ;
  assign n719 = ~n169 & ~n394 ;
  assign n718 = ~n169 & ~n581 ;
  assign n720 = n719 ^ n718 ;
  assign n724 = n723 ^ n720 ;
  assign n780 = n779 ^ n724 ;
  assign n781 = n776 ^ n774 ;
  assign n782 = n770 ^ n729 ;
  assign n783 = x32 & n782 ;
  assign n784 = n783 ^ x32 ;
  assign n785 = n781 & n784 ;
  assign n786 = n785 ^ n784 ;
  assign n787 = ~n780 & n786 ;
  assign n788 = n787 ^ n786 ;
  assign n700 = n699 ^ n659 ;
  assign n502 = x24 ^ x16 ;
  assign n506 = x25 ^ x17 ;
  assign n507 = ~n502 & ~n506 ;
  assign n509 = x26 ^ x18 ;
  assign n515 = x27 ^ x19 ;
  assign n516 = ~n509 & ~n515 ;
  assign n517 = n507 & n516 ;
  assign n519 = x28 ^ x20 ;
  assign n523 = x29 ^ x21 ;
  assign n524 = ~n519 & ~n523 ;
  assign n526 = x30 ^ x22 ;
  assign n536 = x31 ^ x23 ;
  assign n537 = ~n526 & ~n536 ;
  assign n538 = n524 & n537 ;
  assign n539 = n517 & n538 ;
  assign n527 = x23 & x31 ;
  assign n528 = n527 ^ x23 ;
  assign n529 = n526 & n528 ;
  assign n530 = n529 ^ n528 ;
  assign n525 = x22 & ~x30 ;
  assign n531 = n530 ^ n525 ;
  assign n532 = n524 & n531 ;
  assign n520 = x21 & ~x29 ;
  assign n521 = ~n519 & n520 ;
  assign n518 = x20 & ~x28 ;
  assign n522 = n521 ^ n518 ;
  assign n533 = n532 ^ n522 ;
  assign n534 = n517 & n533 ;
  assign n510 = x19 & ~x27 ;
  assign n511 = ~n509 & n510 ;
  assign n508 = x18 & ~x26 ;
  assign n512 = n511 ^ n508 ;
  assign n513 = n507 & n512 ;
  assign n503 = x17 & ~x25 ;
  assign n504 = ~n502 & n503 ;
  assign n501 = x16 & ~x24 ;
  assign n505 = n504 ^ n501 ;
  assign n514 = n513 ^ n505 ;
  assign n535 = n534 ^ n514 ;
  assign n540 = n539 ^ n535 ;
  assign n315 = x24 ^ x8 ;
  assign n319 = x25 ^ x9 ;
  assign n320 = ~n315 & ~n319 ;
  assign n322 = x26 ^ x10 ;
  assign n328 = x27 ^ x11 ;
  assign n329 = ~n322 & ~n328 ;
  assign n330 = n320 & n329 ;
  assign n332 = x28 ^ x12 ;
  assign n336 = x29 ^ x13 ;
  assign n337 = ~n332 & ~n336 ;
  assign n339 = x30 ^ x14 ;
  assign n349 = x31 ^ x15 ;
  assign n350 = ~n339 & ~n349 ;
  assign n351 = n337 & n350 ;
  assign n352 = n330 & n351 ;
  assign n340 = x15 & x31 ;
  assign n341 = n340 ^ x15 ;
  assign n342 = n339 & n341 ;
  assign n343 = n342 ^ n341 ;
  assign n338 = x14 & ~x30 ;
  assign n344 = n343 ^ n338 ;
  assign n345 = n337 & n344 ;
  assign n333 = x13 & ~x29 ;
  assign n334 = ~n332 & n333 ;
  assign n331 = x12 & ~x28 ;
  assign n335 = n334 ^ n331 ;
  assign n346 = n345 ^ n335 ;
  assign n347 = n330 & n346 ;
  assign n323 = x11 & ~x27 ;
  assign n324 = ~n322 & n323 ;
  assign n321 = x10 & ~x26 ;
  assign n325 = n324 ^ n321 ;
  assign n326 = n320 & n325 ;
  assign n316 = x9 & ~x25 ;
  assign n317 = ~n315 & n316 ;
  assign n314 = x8 & ~x24 ;
  assign n318 = n317 ^ n314 ;
  assign n327 = n326 ^ n318 ;
  assign n348 = n347 ^ n327 ;
  assign n353 = n352 ^ n348 ;
  assign n612 = n540 ^ n353 ;
  assign n90 = x24 ^ x0 ;
  assign n94 = x25 ^ x1 ;
  assign n95 = ~n90 & ~n94 ;
  assign n97 = x26 ^ x2 ;
  assign n103 = x27 ^ x3 ;
  assign n104 = ~n97 & ~n103 ;
  assign n105 = n95 & n104 ;
  assign n107 = x28 ^ x4 ;
  assign n111 = x29 ^ x5 ;
  assign n112 = ~n107 & ~n111 ;
  assign n114 = x30 ^ x6 ;
  assign n124 = x31 ^ x7 ;
  assign n125 = ~n114 & ~n124 ;
  assign n126 = n112 & n125 ;
  assign n127 = n105 & n126 ;
  assign n115 = x7 & x31 ;
  assign n116 = n115 ^ x7 ;
  assign n117 = n114 & n116 ;
  assign n118 = n117 ^ n116 ;
  assign n113 = x6 & ~x30 ;
  assign n119 = n118 ^ n113 ;
  assign n120 = n112 & n119 ;
  assign n108 = x5 & ~x29 ;
  assign n109 = ~n107 & n108 ;
  assign n106 = x4 & ~x28 ;
  assign n110 = n109 ^ n106 ;
  assign n121 = n120 ^ n110 ;
  assign n122 = n105 & n121 ;
  assign n98 = x3 & ~x27 ;
  assign n99 = ~n97 & n98 ;
  assign n96 = x2 & ~x26 ;
  assign n100 = n99 ^ n96 ;
  assign n101 = n95 & n100 ;
  assign n91 = x1 & ~x25 ;
  assign n92 = ~n90 & n91 ;
  assign n89 = x0 & ~x24 ;
  assign n93 = n92 ^ n89 ;
  assign n102 = n101 ^ n93 ;
  assign n123 = n122 ^ n102 ;
  assign n128 = n127 ^ n123 ;
  assign n701 = n612 ^ n128 ;
  assign n702 = n700 & n701 ;
  assign n703 = n702 ^ n700 ;
  assign n616 = n353 & n540 ;
  assign n617 = n616 ^ n540 ;
  assign n618 = n617 ^ n353 ;
  assign n613 = n128 & n612 ;
  assign n614 = n613 ^ n612 ;
  assign n619 = n618 ^ n614 ;
  assign n704 = n703 ^ n619 ;
  assign n705 = n659 & n699 ;
  assign n706 = n705 ^ n703 ;
  assign n707 = ~n704 & n706 ;
  assign n708 = n707 ^ n703 ;
  assign n610 = ~n128 & ~n353 ;
  assign n609 = ~n128 & ~n540 ;
  assign n611 = n610 ^ n609 ;
  assign n615 = n614 ^ n611 ;
  assign n709 = n708 ^ n615 ;
  assign n710 = n705 ^ n704 ;
  assign n711 = n701 ^ n700 ;
  assign n712 = x24 & n711 ;
  assign n713 = ~n710 & n712 ;
  assign n714 = n713 ^ n712 ;
  assign n715 = n709 & n714 ;
  assign n716 = n715 ^ n714 ;
  assign n216 = x16 ^ x0 ;
  assign n220 = x17 ^ x1 ;
  assign n221 = ~n216 & ~n220 ;
  assign n223 = x18 ^ x2 ;
  assign n229 = x19 ^ x3 ;
  assign n230 = ~n223 & ~n229 ;
  assign n231 = n221 & n230 ;
  assign n233 = x20 ^ x4 ;
  assign n237 = x21 ^ x5 ;
  assign n238 = ~n233 & ~n237 ;
  assign n240 = x22 ^ x6 ;
  assign n250 = x23 ^ x7 ;
  assign n251 = ~n240 & ~n250 ;
  assign n252 = n238 & n251 ;
  assign n253 = n231 & n252 ;
  assign n241 = x7 & x23 ;
  assign n242 = n241 ^ x7 ;
  assign n243 = n240 & n242 ;
  assign n244 = n243 ^ n242 ;
  assign n239 = x6 & ~x22 ;
  assign n245 = n244 ^ n239 ;
  assign n246 = n238 & n245 ;
  assign n234 = x5 & ~x21 ;
  assign n235 = ~n233 & n234 ;
  assign n232 = x4 & ~x20 ;
  assign n236 = n235 ^ n232 ;
  assign n247 = n246 ^ n236 ;
  assign n248 = n231 & n247 ;
  assign n224 = x3 & ~x19 ;
  assign n225 = ~n223 & n224 ;
  assign n222 = x2 & ~x18 ;
  assign n226 = n225 ^ n222 ;
  assign n227 = n221 & n226 ;
  assign n217 = x1 & ~x17 ;
  assign n218 = ~n216 & n217 ;
  assign n215 = x0 & ~x16 ;
  assign n219 = n218 ^ n215 ;
  assign n228 = n227 ^ n219 ;
  assign n249 = n248 ^ n228 ;
  assign n254 = n253 ^ n249 ;
  assign n401 = x16 ^ x8 ;
  assign n405 = x17 ^ x9 ;
  assign n406 = ~n401 & ~n405 ;
  assign n408 = x18 ^ x10 ;
  assign n414 = x19 ^ x11 ;
  assign n415 = ~n408 & ~n414 ;
  assign n416 = n406 & n415 ;
  assign n418 = x20 ^ x12 ;
  assign n422 = x21 ^ x13 ;
  assign n423 = ~n418 & ~n422 ;
  assign n425 = x22 ^ x14 ;
  assign n435 = x23 ^ x15 ;
  assign n436 = ~n425 & ~n435 ;
  assign n437 = n423 & n436 ;
  assign n438 = n416 & n437 ;
  assign n426 = x15 & x23 ;
  assign n427 = n426 ^ x15 ;
  assign n428 = n425 & n427 ;
  assign n429 = n428 ^ n427 ;
  assign n424 = x14 & ~x22 ;
  assign n430 = n429 ^ n424 ;
  assign n431 = n423 & n430 ;
  assign n419 = x13 & ~x21 ;
  assign n420 = ~n418 & n419 ;
  assign n417 = x12 & ~x20 ;
  assign n421 = n420 ^ n417 ;
  assign n432 = n431 ^ n421 ;
  assign n433 = n416 & n432 ;
  assign n409 = x11 & ~x19 ;
  assign n410 = ~n408 & n409 ;
  assign n407 = x10 & ~x18 ;
  assign n411 = n410 ^ n407 ;
  assign n412 = n406 & n411 ;
  assign n402 = x9 & ~x17 ;
  assign n403 = ~n401 & n402 ;
  assign n400 = x8 & ~x16 ;
  assign n404 = n403 ^ n400 ;
  assign n413 = n412 ^ n404 ;
  assign n434 = n433 ^ n413 ;
  assign n439 = n438 ^ n434 ;
  assign n590 = n254 & n439 ;
  assign n591 = n590 ^ n254 ;
  assign n592 = n591 ^ n439 ;
  assign n587 = n439 ^ n254 ;
  assign n584 = n581 ^ n500 ;
  assign n588 = n584 ^ n540 ;
  assign n589 = n587 & n588 ;
  assign n593 = n592 ^ n589 ;
  assign n594 = n500 & n581 ;
  assign n585 = n540 & n584 ;
  assign n595 = n594 ^ n585 ;
  assign n596 = n595 ^ n589 ;
  assign n597 = ~n593 & n596 ;
  assign n598 = n597 ^ n589 ;
  assign n582 = n540 & ~n581 ;
  assign n541 = ~n500 & n540 ;
  assign n583 = n582 ^ n541 ;
  assign n586 = n585 ^ n583 ;
  assign n599 = n598 ^ n586 ;
  assign n600 = n595 ^ n593 ;
  assign n601 = n588 ^ n587 ;
  assign n602 = x16 & n601 ;
  assign n603 = n602 ^ x16 ;
  assign n604 = ~n600 & n603 ;
  assign n605 = n604 ^ n603 ;
  assign n606 = n599 & n605 ;
  assign n607 = n606 ^ n605 ;
  assign n176 = x8 ^ x0 ;
  assign n180 = x9 ^ x1 ;
  assign n181 = ~n176 & ~n180 ;
  assign n183 = x10 ^ x2 ;
  assign n189 = x11 ^ x3 ;
  assign n190 = ~n183 & ~n189 ;
  assign n191 = n181 & n190 ;
  assign n193 = x12 ^ x4 ;
  assign n197 = x13 ^ x5 ;
  assign n198 = ~n193 & ~n197 ;
  assign n200 = x14 ^ x6 ;
  assign n210 = x15 ^ x7 ;
  assign n211 = ~n200 & ~n210 ;
  assign n212 = n198 & n211 ;
  assign n213 = n191 & n212 ;
  assign n201 = x7 & x15 ;
  assign n202 = n201 ^ x7 ;
  assign n203 = n200 & n202 ;
  assign n204 = n203 ^ n202 ;
  assign n199 = x6 & ~x14 ;
  assign n205 = n204 ^ n199 ;
  assign n206 = n198 & n205 ;
  assign n194 = x5 & ~x13 ;
  assign n195 = ~n193 & n194 ;
  assign n192 = x4 & ~x12 ;
  assign n196 = n195 ^ n192 ;
  assign n207 = n206 ^ n196 ;
  assign n208 = n191 & n207 ;
  assign n184 = x3 & ~x11 ;
  assign n185 = ~n183 & n184 ;
  assign n182 = x2 & ~x10 ;
  assign n186 = n185 ^ n182 ;
  assign n187 = n181 & n186 ;
  assign n177 = x1 & ~x9 ;
  assign n178 = ~n176 & n177 ;
  assign n175 = x0 & ~x8 ;
  assign n179 = n178 ^ n175 ;
  assign n188 = n187 ^ n179 ;
  assign n209 = n208 ^ n188 ;
  assign n214 = n213 ^ n209 ;
  assign n444 = n214 & n439 ;
  assign n445 = n444 ^ n439 ;
  assign n440 = n439 ^ n214 ;
  assign n397 = n394 ^ n313 ;
  assign n441 = n397 ^ n353 ;
  assign n442 = n440 & n441 ;
  assign n443 = n442 ^ n441 ;
  assign n446 = n445 ^ n443 ;
  assign n447 = n313 & n394 ;
  assign n398 = n353 & n397 ;
  assign n448 = n447 ^ n398 ;
  assign n449 = n448 ^ n443 ;
  assign n450 = n446 & n449 ;
  assign n451 = n450 ^ n443 ;
  assign n395 = n353 & ~n394 ;
  assign n354 = ~n313 & n353 ;
  assign n396 = n395 ^ n354 ;
  assign n399 = n398 ^ n396 ;
  assign n452 = n451 ^ n399 ;
  assign n453 = n448 ^ n446 ;
  assign n454 = n441 ^ n440 ;
  assign n455 = x8 & n454 ;
  assign n456 = n453 & n455 ;
  assign n457 = n456 ^ n455 ;
  assign n458 = n452 & n457 ;
  assign n459 = n458 ^ n457 ;
  assign n258 = n214 & n254 ;
  assign n255 = n254 ^ n214 ;
  assign n172 = n169 ^ n88 ;
  assign n256 = n172 ^ n128 ;
  assign n257 = n255 & n256 ;
  assign n259 = n258 ^ n257 ;
  assign n260 = n88 & n169 ;
  assign n173 = n128 & n172 ;
  assign n261 = n260 ^ n173 ;
  assign n262 = n261 ^ n257 ;
  assign n263 = n259 & n262 ;
  assign n264 = n263 ^ n257 ;
  assign n170 = n128 & ~n169 ;
  assign n129 = ~n88 & n128 ;
  assign n171 = n170 ^ n129 ;
  assign n174 = n173 ^ n171 ;
  assign n265 = n264 ^ n174 ;
  assign n266 = n261 ^ n259 ;
  assign n267 = n256 ^ n255 ;
  assign n268 = x0 & n267 ;
  assign n269 = n268 ^ x0 ;
  assign n270 = n266 & n269 ;
  assign n271 = n270 ^ n269 ;
  assign n272 = n265 & n271 ;
  assign n273 = n272 ^ n271 ;
  assign n460 = n459 ^ n273 ;
  assign n608 = n607 ^ n460 ;
  assign n717 = n716 ^ n608 ;
  assign n789 = n788 ^ n717 ;
  assign n820 = n819 ^ n789 ;
  assign n853 = x41 & n814 ;
  assign n854 = n813 & n853 ;
  assign n855 = n854 ^ n853 ;
  assign n856 = n812 & n855 ;
  assign n857 = n856 ^ n855 ;
  assign n846 = x33 & n782 ;
  assign n847 = n846 ^ x33 ;
  assign n848 = n781 & n847 ;
  assign n849 = n848 ^ n847 ;
  assign n850 = ~n780 & n849 ;
  assign n851 = n850 ^ n849 ;
  assign n840 = x25 & n711 ;
  assign n841 = ~n710 & n840 ;
  assign n842 = n841 ^ n840 ;
  assign n843 = n709 & n842 ;
  assign n844 = n843 ^ n842 ;
  assign n833 = x17 & n601 ;
  assign n834 = n833 ^ x17 ;
  assign n835 = ~n600 & n834 ;
  assign n836 = n835 ^ n834 ;
  assign n837 = n599 & n836 ;
  assign n838 = n837 ^ n836 ;
  assign n827 = x9 & n454 ;
  assign n828 = n453 & n827 ;
  assign n829 = n828 ^ n827 ;
  assign n830 = n452 & n829 ;
  assign n831 = n830 ^ n829 ;
  assign n821 = x1 & n267 ;
  assign n822 = n821 ^ x1 ;
  assign n823 = n266 & n822 ;
  assign n824 = n823 ^ n822 ;
  assign n825 = n265 & n824 ;
  assign n826 = n825 ^ n824 ;
  assign n832 = n831 ^ n826 ;
  assign n839 = n838 ^ n832 ;
  assign n845 = n844 ^ n839 ;
  assign n852 = n851 ^ n845 ;
  assign n858 = n857 ^ n852 ;
  assign n891 = x42 & n814 ;
  assign n892 = n813 & n891 ;
  assign n893 = n892 ^ n891 ;
  assign n894 = n812 & n893 ;
  assign n895 = n894 ^ n893 ;
  assign n884 = x34 & n782 ;
  assign n885 = n884 ^ x34 ;
  assign n886 = n781 & n885 ;
  assign n887 = n886 ^ n885 ;
  assign n888 = ~n780 & n887 ;
  assign n889 = n888 ^ n887 ;
  assign n878 = x26 & n711 ;
  assign n879 = ~n710 & n878 ;
  assign n880 = n879 ^ n878 ;
  assign n881 = n709 & n880 ;
  assign n882 = n881 ^ n880 ;
  assign n871 = x18 & n601 ;
  assign n872 = n871 ^ x18 ;
  assign n873 = ~n600 & n872 ;
  assign n874 = n873 ^ n872 ;
  assign n875 = n599 & n874 ;
  assign n876 = n875 ^ n874 ;
  assign n865 = x10 & n454 ;
  assign n866 = n453 & n865 ;
  assign n867 = n866 ^ n865 ;
  assign n868 = n452 & n867 ;
  assign n869 = n868 ^ n867 ;
  assign n859 = x2 & n267 ;
  assign n860 = n859 ^ x2 ;
  assign n861 = n266 & n860 ;
  assign n862 = n861 ^ n860 ;
  assign n863 = n265 & n862 ;
  assign n864 = n863 ^ n862 ;
  assign n870 = n869 ^ n864 ;
  assign n877 = n876 ^ n870 ;
  assign n883 = n882 ^ n877 ;
  assign n890 = n889 ^ n883 ;
  assign n896 = n895 ^ n890 ;
  assign n929 = x43 & n814 ;
  assign n930 = n813 & n929 ;
  assign n931 = n930 ^ n929 ;
  assign n932 = n812 & n931 ;
  assign n933 = n932 ^ n931 ;
  assign n922 = x35 & n782 ;
  assign n923 = n922 ^ x35 ;
  assign n924 = n781 & n923 ;
  assign n925 = n924 ^ n923 ;
  assign n926 = ~n780 & n925 ;
  assign n927 = n926 ^ n925 ;
  assign n916 = x27 & n711 ;
  assign n917 = ~n710 & n916 ;
  assign n918 = n917 ^ n916 ;
  assign n919 = n709 & n918 ;
  assign n920 = n919 ^ n918 ;
  assign n909 = x19 & n601 ;
  assign n910 = n909 ^ x19 ;
  assign n911 = ~n600 & n910 ;
  assign n912 = n911 ^ n910 ;
  assign n913 = n599 & n912 ;
  assign n914 = n913 ^ n912 ;
  assign n903 = x11 & n454 ;
  assign n904 = n453 & n903 ;
  assign n905 = n904 ^ n903 ;
  assign n906 = n452 & n905 ;
  assign n907 = n906 ^ n905 ;
  assign n897 = x3 & n267 ;
  assign n898 = n897 ^ x3 ;
  assign n899 = n266 & n898 ;
  assign n900 = n899 ^ n898 ;
  assign n901 = n265 & n900 ;
  assign n902 = n901 ^ n900 ;
  assign n908 = n907 ^ n902 ;
  assign n915 = n914 ^ n908 ;
  assign n921 = n920 ^ n915 ;
  assign n928 = n927 ^ n921 ;
  assign n934 = n933 ^ n928 ;
  assign n967 = x44 & n814 ;
  assign n968 = n813 & n967 ;
  assign n969 = n968 ^ n967 ;
  assign n970 = n812 & n969 ;
  assign n971 = n970 ^ n969 ;
  assign n960 = x36 & n782 ;
  assign n961 = n960 ^ x36 ;
  assign n962 = n781 & n961 ;
  assign n963 = n962 ^ n961 ;
  assign n964 = ~n780 & n963 ;
  assign n965 = n964 ^ n963 ;
  assign n954 = x28 & n711 ;
  assign n955 = ~n710 & n954 ;
  assign n956 = n955 ^ n954 ;
  assign n957 = n709 & n956 ;
  assign n958 = n957 ^ n956 ;
  assign n947 = x20 & n601 ;
  assign n948 = n947 ^ x20 ;
  assign n949 = ~n600 & n948 ;
  assign n950 = n949 ^ n948 ;
  assign n951 = n599 & n950 ;
  assign n952 = n951 ^ n950 ;
  assign n941 = x12 & n454 ;
  assign n942 = n453 & n941 ;
  assign n943 = n942 ^ n941 ;
  assign n944 = n452 & n943 ;
  assign n945 = n944 ^ n943 ;
  assign n935 = x4 & n267 ;
  assign n936 = n935 ^ x4 ;
  assign n937 = n266 & n936 ;
  assign n938 = n937 ^ n936 ;
  assign n939 = n265 & n938 ;
  assign n940 = n939 ^ n938 ;
  assign n946 = n945 ^ n940 ;
  assign n953 = n952 ^ n946 ;
  assign n959 = n958 ^ n953 ;
  assign n966 = n965 ^ n959 ;
  assign n972 = n971 ^ n966 ;
  assign n1005 = x45 & n814 ;
  assign n1006 = n813 & n1005 ;
  assign n1007 = n1006 ^ n1005 ;
  assign n1008 = n812 & n1007 ;
  assign n1009 = n1008 ^ n1007 ;
  assign n998 = x37 & n782 ;
  assign n999 = n998 ^ x37 ;
  assign n1000 = n781 & n999 ;
  assign n1001 = n1000 ^ n999 ;
  assign n1002 = ~n780 & n1001 ;
  assign n1003 = n1002 ^ n1001 ;
  assign n992 = x29 & n711 ;
  assign n993 = ~n710 & n992 ;
  assign n994 = n993 ^ n992 ;
  assign n995 = n709 & n994 ;
  assign n996 = n995 ^ n994 ;
  assign n985 = x21 & n601 ;
  assign n986 = n985 ^ x21 ;
  assign n987 = ~n600 & n986 ;
  assign n988 = n987 ^ n986 ;
  assign n989 = n599 & n988 ;
  assign n990 = n989 ^ n988 ;
  assign n979 = x13 & n454 ;
  assign n980 = n453 & n979 ;
  assign n981 = n980 ^ n979 ;
  assign n982 = n452 & n981 ;
  assign n983 = n982 ^ n981 ;
  assign n973 = x5 & n267 ;
  assign n974 = n973 ^ x5 ;
  assign n975 = n266 & n974 ;
  assign n976 = n975 ^ n974 ;
  assign n977 = n265 & n976 ;
  assign n978 = n977 ^ n976 ;
  assign n984 = n983 ^ n978 ;
  assign n991 = n990 ^ n984 ;
  assign n997 = n996 ^ n991 ;
  assign n1004 = n1003 ^ n997 ;
  assign n1010 = n1009 ^ n1004 ;
  assign n1043 = x46 & n814 ;
  assign n1044 = n813 & n1043 ;
  assign n1045 = n1044 ^ n1043 ;
  assign n1046 = n812 & n1045 ;
  assign n1047 = n1046 ^ n1045 ;
  assign n1036 = x38 & n782 ;
  assign n1037 = n1036 ^ x38 ;
  assign n1038 = n781 & n1037 ;
  assign n1039 = n1038 ^ n1037 ;
  assign n1040 = ~n780 & n1039 ;
  assign n1041 = n1040 ^ n1039 ;
  assign n1030 = x30 & n711 ;
  assign n1031 = ~n710 & n1030 ;
  assign n1032 = n1031 ^ n1030 ;
  assign n1033 = n709 & n1032 ;
  assign n1034 = n1033 ^ n1032 ;
  assign n1023 = x22 & n601 ;
  assign n1024 = n1023 ^ x22 ;
  assign n1025 = ~n600 & n1024 ;
  assign n1026 = n1025 ^ n1024 ;
  assign n1027 = n599 & n1026 ;
  assign n1028 = n1027 ^ n1026 ;
  assign n1017 = x14 & n454 ;
  assign n1018 = n453 & n1017 ;
  assign n1019 = n1018 ^ n1017 ;
  assign n1020 = n452 & n1019 ;
  assign n1021 = n1020 ^ n1019 ;
  assign n1011 = x6 & n267 ;
  assign n1012 = n1011 ^ x6 ;
  assign n1013 = n266 & n1012 ;
  assign n1014 = n1013 ^ n1012 ;
  assign n1015 = n265 & n1014 ;
  assign n1016 = n1015 ^ n1014 ;
  assign n1022 = n1021 ^ n1016 ;
  assign n1029 = n1028 ^ n1022 ;
  assign n1035 = n1034 ^ n1029 ;
  assign n1042 = n1041 ^ n1035 ;
  assign n1048 = n1047 ^ n1042 ;
  assign n1081 = x47 & n814 ;
  assign n1082 = n813 & n1081 ;
  assign n1083 = n1082 ^ n1081 ;
  assign n1084 = n812 & n1083 ;
  assign n1085 = n1084 ^ n1083 ;
  assign n1074 = x39 & n782 ;
  assign n1075 = n1074 ^ x39 ;
  assign n1076 = n781 & n1075 ;
  assign n1077 = n1076 ^ n1075 ;
  assign n1078 = ~n780 & n1077 ;
  assign n1079 = n1078 ^ n1077 ;
  assign n1068 = x31 & n711 ;
  assign n1069 = ~n710 & n1068 ;
  assign n1070 = n1069 ^ n1068 ;
  assign n1071 = n709 & n1070 ;
  assign n1072 = n1071 ^ n1070 ;
  assign n1061 = x23 & n601 ;
  assign n1062 = n1061 ^ x23 ;
  assign n1063 = ~n600 & n1062 ;
  assign n1064 = n1063 ^ n1062 ;
  assign n1065 = n599 & n1064 ;
  assign n1066 = n1065 ^ n1064 ;
  assign n1055 = x15 & n454 ;
  assign n1056 = n453 & n1055 ;
  assign n1057 = n1056 ^ n1055 ;
  assign n1058 = n452 & n1057 ;
  assign n1059 = n1058 ^ n1057 ;
  assign n1049 = x7 & n267 ;
  assign n1050 = n1049 ^ x7 ;
  assign n1051 = n266 & n1050 ;
  assign n1052 = n1051 ^ n1050 ;
  assign n1053 = n265 & n1052 ;
  assign n1054 = n1053 ^ n1052 ;
  assign n1060 = n1059 ^ n1054 ;
  assign n1067 = n1066 ^ n1060 ;
  assign n1073 = n1072 ^ n1067 ;
  assign n1080 = n1079 ^ n1073 ;
  assign n1086 = n1085 ^ n1080 ;
  assign n1113 = n815 ^ x40 ;
  assign n1114 = n813 & n1113 ;
  assign n1115 = n1114 ^ n1113 ;
  assign n1116 = n812 & n1115 ;
  assign n1117 = n1116 ^ n1115 ;
  assign n1108 = n781 & n783 ;
  assign n1109 = n1108 ^ n783 ;
  assign n1110 = ~n780 & n1109 ;
  assign n1111 = n1110 ^ n1109 ;
  assign n1102 = n712 ^ x24 ;
  assign n1103 = ~n710 & n1102 ;
  assign n1104 = n1103 ^ n1102 ;
  assign n1105 = n709 & n1104 ;
  assign n1106 = n1105 ^ n1104 ;
  assign n1097 = ~n600 & n602 ;
  assign n1098 = n1097 ^ n602 ;
  assign n1099 = n599 & n1098 ;
  assign n1100 = n1099 ^ n1098 ;
  assign n1091 = n455 ^ x8 ;
  assign n1092 = n453 & n1091 ;
  assign n1093 = n1092 ^ n1091 ;
  assign n1094 = n452 & n1093 ;
  assign n1095 = n1094 ^ n1093 ;
  assign n1087 = n266 & n268 ;
  assign n1088 = n1087 ^ n268 ;
  assign n1089 = n265 & n1088 ;
  assign n1090 = n1089 ^ n1088 ;
  assign n1096 = n1095 ^ n1090 ;
  assign n1101 = n1100 ^ n1096 ;
  assign n1107 = n1106 ^ n1101 ;
  assign n1112 = n1111 ^ n1107 ;
  assign n1118 = n1117 ^ n1112 ;
  assign n1145 = n853 ^ x41 ;
  assign n1146 = n813 & n1145 ;
  assign n1147 = n1146 ^ n1145 ;
  assign n1148 = n812 & n1147 ;
  assign n1149 = n1148 ^ n1147 ;
  assign n1140 = n781 & n846 ;
  assign n1141 = n1140 ^ n846 ;
  assign n1142 = ~n780 & n1141 ;
  assign n1143 = n1142 ^ n1141 ;
  assign n1134 = n840 ^ x25 ;
  assign n1135 = ~n710 & n1134 ;
  assign n1136 = n1135 ^ n1134 ;
  assign n1137 = n709 & n1136 ;
  assign n1138 = n1137 ^ n1136 ;
  assign n1129 = ~n600 & n833 ;
  assign n1130 = n1129 ^ n833 ;
  assign n1131 = n599 & n1130 ;
  assign n1132 = n1131 ^ n1130 ;
  assign n1123 = n827 ^ x9 ;
  assign n1124 = n453 & n1123 ;
  assign n1125 = n1124 ^ n1123 ;
  assign n1126 = n452 & n1125 ;
  assign n1127 = n1126 ^ n1125 ;
  assign n1119 = n266 & n821 ;
  assign n1120 = n1119 ^ n821 ;
  assign n1121 = n265 & n1120 ;
  assign n1122 = n1121 ^ n1120 ;
  assign n1128 = n1127 ^ n1122 ;
  assign n1133 = n1132 ^ n1128 ;
  assign n1139 = n1138 ^ n1133 ;
  assign n1144 = n1143 ^ n1139 ;
  assign n1150 = n1149 ^ n1144 ;
  assign n1177 = n891 ^ x42 ;
  assign n1178 = n813 & n1177 ;
  assign n1179 = n1178 ^ n1177 ;
  assign n1180 = n812 & n1179 ;
  assign n1181 = n1180 ^ n1179 ;
  assign n1172 = n781 & n884 ;
  assign n1173 = n1172 ^ n884 ;
  assign n1174 = ~n780 & n1173 ;
  assign n1175 = n1174 ^ n1173 ;
  assign n1166 = n878 ^ x26 ;
  assign n1167 = ~n710 & n1166 ;
  assign n1168 = n1167 ^ n1166 ;
  assign n1169 = n709 & n1168 ;
  assign n1170 = n1169 ^ n1168 ;
  assign n1161 = ~n600 & n871 ;
  assign n1162 = n1161 ^ n871 ;
  assign n1163 = n599 & n1162 ;
  assign n1164 = n1163 ^ n1162 ;
  assign n1155 = n865 ^ x10 ;
  assign n1156 = n453 & n1155 ;
  assign n1157 = n1156 ^ n1155 ;
  assign n1158 = n452 & n1157 ;
  assign n1159 = n1158 ^ n1157 ;
  assign n1151 = n266 & n859 ;
  assign n1152 = n1151 ^ n859 ;
  assign n1153 = n265 & n1152 ;
  assign n1154 = n1153 ^ n1152 ;
  assign n1160 = n1159 ^ n1154 ;
  assign n1165 = n1164 ^ n1160 ;
  assign n1171 = n1170 ^ n1165 ;
  assign n1176 = n1175 ^ n1171 ;
  assign n1182 = n1181 ^ n1176 ;
  assign n1209 = n929 ^ x43 ;
  assign n1210 = n813 & n1209 ;
  assign n1211 = n1210 ^ n1209 ;
  assign n1212 = n812 & n1211 ;
  assign n1213 = n1212 ^ n1211 ;
  assign n1204 = n781 & n922 ;
  assign n1205 = n1204 ^ n922 ;
  assign n1206 = ~n780 & n1205 ;
  assign n1207 = n1206 ^ n1205 ;
  assign n1198 = n916 ^ x27 ;
  assign n1199 = ~n710 & n1198 ;
  assign n1200 = n1199 ^ n1198 ;
  assign n1201 = n709 & n1200 ;
  assign n1202 = n1201 ^ n1200 ;
  assign n1193 = ~n600 & n909 ;
  assign n1194 = n1193 ^ n909 ;
  assign n1195 = n599 & n1194 ;
  assign n1196 = n1195 ^ n1194 ;
  assign n1187 = n903 ^ x11 ;
  assign n1188 = n453 & n1187 ;
  assign n1189 = n1188 ^ n1187 ;
  assign n1190 = n452 & n1189 ;
  assign n1191 = n1190 ^ n1189 ;
  assign n1183 = n266 & n897 ;
  assign n1184 = n1183 ^ n897 ;
  assign n1185 = n265 & n1184 ;
  assign n1186 = n1185 ^ n1184 ;
  assign n1192 = n1191 ^ n1186 ;
  assign n1197 = n1196 ^ n1192 ;
  assign n1203 = n1202 ^ n1197 ;
  assign n1208 = n1207 ^ n1203 ;
  assign n1214 = n1213 ^ n1208 ;
  assign n1241 = n967 ^ x44 ;
  assign n1242 = n813 & n1241 ;
  assign n1243 = n1242 ^ n1241 ;
  assign n1244 = n812 & n1243 ;
  assign n1245 = n1244 ^ n1243 ;
  assign n1236 = n781 & n960 ;
  assign n1237 = n1236 ^ n960 ;
  assign n1238 = ~n780 & n1237 ;
  assign n1239 = n1238 ^ n1237 ;
  assign n1230 = n954 ^ x28 ;
  assign n1231 = ~n710 & n1230 ;
  assign n1232 = n1231 ^ n1230 ;
  assign n1233 = n709 & n1232 ;
  assign n1234 = n1233 ^ n1232 ;
  assign n1225 = ~n600 & n947 ;
  assign n1226 = n1225 ^ n947 ;
  assign n1227 = n599 & n1226 ;
  assign n1228 = n1227 ^ n1226 ;
  assign n1219 = n941 ^ x12 ;
  assign n1220 = n453 & n1219 ;
  assign n1221 = n1220 ^ n1219 ;
  assign n1222 = n452 & n1221 ;
  assign n1223 = n1222 ^ n1221 ;
  assign n1215 = n266 & n935 ;
  assign n1216 = n1215 ^ n935 ;
  assign n1217 = n265 & n1216 ;
  assign n1218 = n1217 ^ n1216 ;
  assign n1224 = n1223 ^ n1218 ;
  assign n1229 = n1228 ^ n1224 ;
  assign n1235 = n1234 ^ n1229 ;
  assign n1240 = n1239 ^ n1235 ;
  assign n1246 = n1245 ^ n1240 ;
  assign n1273 = n1005 ^ x45 ;
  assign n1274 = n813 & n1273 ;
  assign n1275 = n1274 ^ n1273 ;
  assign n1276 = n812 & n1275 ;
  assign n1277 = n1276 ^ n1275 ;
  assign n1268 = n781 & n998 ;
  assign n1269 = n1268 ^ n998 ;
  assign n1270 = ~n780 & n1269 ;
  assign n1271 = n1270 ^ n1269 ;
  assign n1262 = n992 ^ x29 ;
  assign n1263 = ~n710 & n1262 ;
  assign n1264 = n1263 ^ n1262 ;
  assign n1265 = n709 & n1264 ;
  assign n1266 = n1265 ^ n1264 ;
  assign n1257 = ~n600 & n985 ;
  assign n1258 = n1257 ^ n985 ;
  assign n1259 = n599 & n1258 ;
  assign n1260 = n1259 ^ n1258 ;
  assign n1251 = n979 ^ x13 ;
  assign n1252 = n453 & n1251 ;
  assign n1253 = n1252 ^ n1251 ;
  assign n1254 = n452 & n1253 ;
  assign n1255 = n1254 ^ n1253 ;
  assign n1247 = n266 & n973 ;
  assign n1248 = n1247 ^ n973 ;
  assign n1249 = n265 & n1248 ;
  assign n1250 = n1249 ^ n1248 ;
  assign n1256 = n1255 ^ n1250 ;
  assign n1261 = n1260 ^ n1256 ;
  assign n1267 = n1266 ^ n1261 ;
  assign n1272 = n1271 ^ n1267 ;
  assign n1278 = n1277 ^ n1272 ;
  assign n1305 = n1043 ^ x46 ;
  assign n1306 = n813 & n1305 ;
  assign n1307 = n1306 ^ n1305 ;
  assign n1308 = n812 & n1307 ;
  assign n1309 = n1308 ^ n1307 ;
  assign n1300 = n781 & n1036 ;
  assign n1301 = n1300 ^ n1036 ;
  assign n1302 = ~n780 & n1301 ;
  assign n1303 = n1302 ^ n1301 ;
  assign n1294 = n1030 ^ x30 ;
  assign n1295 = ~n710 & n1294 ;
  assign n1296 = n1295 ^ n1294 ;
  assign n1297 = n709 & n1296 ;
  assign n1298 = n1297 ^ n1296 ;
  assign n1289 = ~n600 & n1023 ;
  assign n1290 = n1289 ^ n1023 ;
  assign n1291 = n599 & n1290 ;
  assign n1292 = n1291 ^ n1290 ;
  assign n1283 = n1017 ^ x14 ;
  assign n1284 = n453 & n1283 ;
  assign n1285 = n1284 ^ n1283 ;
  assign n1286 = n452 & n1285 ;
  assign n1287 = n1286 ^ n1285 ;
  assign n1279 = n266 & n1011 ;
  assign n1280 = n1279 ^ n1011 ;
  assign n1281 = n265 & n1280 ;
  assign n1282 = n1281 ^ n1280 ;
  assign n1288 = n1287 ^ n1282 ;
  assign n1293 = n1292 ^ n1288 ;
  assign n1299 = n1298 ^ n1293 ;
  assign n1304 = n1303 ^ n1299 ;
  assign n1310 = n1309 ^ n1304 ;
  assign n1337 = n1081 ^ x47 ;
  assign n1338 = n813 & n1337 ;
  assign n1339 = n1338 ^ n1337 ;
  assign n1340 = n812 & n1339 ;
  assign n1341 = n1340 ^ n1339 ;
  assign n1332 = n781 & n1074 ;
  assign n1333 = n1332 ^ n1074 ;
  assign n1334 = ~n780 & n1333 ;
  assign n1335 = n1334 ^ n1333 ;
  assign n1326 = n1068 ^ x31 ;
  assign n1327 = ~n710 & n1326 ;
  assign n1328 = n1327 ^ n1326 ;
  assign n1329 = n709 & n1328 ;
  assign n1330 = n1329 ^ n1328 ;
  assign n1321 = ~n600 & n1061 ;
  assign n1322 = n1321 ^ n1061 ;
  assign n1323 = n599 & n1322 ;
  assign n1324 = n1323 ^ n1322 ;
  assign n1315 = n1055 ^ x15 ;
  assign n1316 = n453 & n1315 ;
  assign n1317 = n1316 ^ n1315 ;
  assign n1318 = n452 & n1317 ;
  assign n1319 = n1318 ^ n1317 ;
  assign n1311 = n266 & n1049 ;
  assign n1312 = n1311 ^ n1049 ;
  assign n1313 = n265 & n1312 ;
  assign n1314 = n1313 ^ n1312 ;
  assign n1320 = n1319 ^ n1314 ;
  assign n1325 = n1324 ^ n1320 ;
  assign n1331 = n1330 ^ n1325 ;
  assign n1336 = n1335 ^ n1331 ;
  assign n1342 = n1341 ^ n1336 ;
  assign n1357 = n812 & n816 ;
  assign n1358 = n1357 ^ n816 ;
  assign n1354 = ~n780 & n785 ;
  assign n1355 = n1354 ^ n785 ;
  assign n1351 = n709 & n713 ;
  assign n1352 = n1351 ^ n713 ;
  assign n1348 = n599 & n604 ;
  assign n1349 = n1348 ^ n604 ;
  assign n1345 = n452 & n456 ;
  assign n1346 = n1345 ^ n456 ;
  assign n1343 = n265 & n270 ;
  assign n1344 = n1343 ^ n270 ;
  assign n1347 = n1346 ^ n1344 ;
  assign n1350 = n1349 ^ n1347 ;
  assign n1353 = n1352 ^ n1350 ;
  assign n1356 = n1355 ^ n1353 ;
  assign n1359 = n1358 ^ n1356 ;
  assign n1374 = n812 & n854 ;
  assign n1375 = n1374 ^ n854 ;
  assign n1371 = ~n780 & n848 ;
  assign n1372 = n1371 ^ n848 ;
  assign n1368 = n709 & n841 ;
  assign n1369 = n1368 ^ n841 ;
  assign n1365 = n599 & n835 ;
  assign n1366 = n1365 ^ n835 ;
  assign n1362 = n452 & n828 ;
  assign n1363 = n1362 ^ n828 ;
  assign n1360 = n265 & n823 ;
  assign n1361 = n1360 ^ n823 ;
  assign n1364 = n1363 ^ n1361 ;
  assign n1367 = n1366 ^ n1364 ;
  assign n1370 = n1369 ^ n1367 ;
  assign n1373 = n1372 ^ n1370 ;
  assign n1376 = n1375 ^ n1373 ;
  assign n1391 = n812 & n892 ;
  assign n1392 = n1391 ^ n892 ;
  assign n1388 = ~n780 & n886 ;
  assign n1389 = n1388 ^ n886 ;
  assign n1385 = n709 & n879 ;
  assign n1386 = n1385 ^ n879 ;
  assign n1382 = n599 & n873 ;
  assign n1383 = n1382 ^ n873 ;
  assign n1379 = n452 & n866 ;
  assign n1380 = n1379 ^ n866 ;
  assign n1377 = n265 & n861 ;
  assign n1378 = n1377 ^ n861 ;
  assign n1381 = n1380 ^ n1378 ;
  assign n1384 = n1383 ^ n1381 ;
  assign n1387 = n1386 ^ n1384 ;
  assign n1390 = n1389 ^ n1387 ;
  assign n1393 = n1392 ^ n1390 ;
  assign n1408 = n812 & n930 ;
  assign n1409 = n1408 ^ n930 ;
  assign n1405 = ~n780 & n924 ;
  assign n1406 = n1405 ^ n924 ;
  assign n1402 = n709 & n917 ;
  assign n1403 = n1402 ^ n917 ;
  assign n1399 = n599 & n911 ;
  assign n1400 = n1399 ^ n911 ;
  assign n1396 = n452 & n904 ;
  assign n1397 = n1396 ^ n904 ;
  assign n1394 = n265 & n899 ;
  assign n1395 = n1394 ^ n899 ;
  assign n1398 = n1397 ^ n1395 ;
  assign n1401 = n1400 ^ n1398 ;
  assign n1404 = n1403 ^ n1401 ;
  assign n1407 = n1406 ^ n1404 ;
  assign n1410 = n1409 ^ n1407 ;
  assign n1425 = n812 & n968 ;
  assign n1426 = n1425 ^ n968 ;
  assign n1422 = ~n780 & n962 ;
  assign n1423 = n1422 ^ n962 ;
  assign n1419 = n709 & n955 ;
  assign n1420 = n1419 ^ n955 ;
  assign n1416 = n599 & n949 ;
  assign n1417 = n1416 ^ n949 ;
  assign n1413 = n452 & n942 ;
  assign n1414 = n1413 ^ n942 ;
  assign n1411 = n265 & n937 ;
  assign n1412 = n1411 ^ n937 ;
  assign n1415 = n1414 ^ n1412 ;
  assign n1418 = n1417 ^ n1415 ;
  assign n1421 = n1420 ^ n1418 ;
  assign n1424 = n1423 ^ n1421 ;
  assign n1427 = n1426 ^ n1424 ;
  assign n1442 = n812 & n1006 ;
  assign n1443 = n1442 ^ n1006 ;
  assign n1439 = ~n780 & n1000 ;
  assign n1440 = n1439 ^ n1000 ;
  assign n1436 = n709 & n993 ;
  assign n1437 = n1436 ^ n993 ;
  assign n1433 = n599 & n987 ;
  assign n1434 = n1433 ^ n987 ;
  assign n1430 = n452 & n980 ;
  assign n1431 = n1430 ^ n980 ;
  assign n1428 = n265 & n975 ;
  assign n1429 = n1428 ^ n975 ;
  assign n1432 = n1431 ^ n1429 ;
  assign n1435 = n1434 ^ n1432 ;
  assign n1438 = n1437 ^ n1435 ;
  assign n1441 = n1440 ^ n1438 ;
  assign n1444 = n1443 ^ n1441 ;
  assign n1459 = n812 & n1044 ;
  assign n1460 = n1459 ^ n1044 ;
  assign n1456 = ~n780 & n1038 ;
  assign n1457 = n1456 ^ n1038 ;
  assign n1453 = n709 & n1031 ;
  assign n1454 = n1453 ^ n1031 ;
  assign n1450 = n599 & n1025 ;
  assign n1451 = n1450 ^ n1025 ;
  assign n1447 = n452 & n1018 ;
  assign n1448 = n1447 ^ n1018 ;
  assign n1445 = n265 & n1013 ;
  assign n1446 = n1445 ^ n1013 ;
  assign n1449 = n1448 ^ n1446 ;
  assign n1452 = n1451 ^ n1449 ;
  assign n1455 = n1454 ^ n1452 ;
  assign n1458 = n1457 ^ n1455 ;
  assign n1461 = n1460 ^ n1458 ;
  assign n1476 = n812 & n1082 ;
  assign n1477 = n1476 ^ n1082 ;
  assign n1473 = ~n780 & n1076 ;
  assign n1474 = n1473 ^ n1076 ;
  assign n1470 = n709 & n1069 ;
  assign n1471 = n1470 ^ n1069 ;
  assign n1467 = n599 & n1063 ;
  assign n1468 = n1467 ^ n1063 ;
  assign n1464 = n452 & n1056 ;
  assign n1465 = n1464 ^ n1056 ;
  assign n1462 = n265 & n1051 ;
  assign n1463 = n1462 ^ n1051 ;
  assign n1466 = n1465 ^ n1463 ;
  assign n1469 = n1468 ^ n1466 ;
  assign n1472 = n1471 ^ n1469 ;
  assign n1475 = n1474 ^ n1472 ;
  assign n1478 = n1477 ^ n1475 ;
  assign n1493 = n812 & n1114 ;
  assign n1494 = n1493 ^ n1114 ;
  assign n1490 = ~n780 & n1108 ;
  assign n1491 = n1490 ^ n1108 ;
  assign n1487 = n709 & n1103 ;
  assign n1488 = n1487 ^ n1103 ;
  assign n1484 = n599 & n1097 ;
  assign n1485 = n1484 ^ n1097 ;
  assign n1481 = n452 & n1092 ;
  assign n1482 = n1481 ^ n1092 ;
  assign n1479 = n265 & n1087 ;
  assign n1480 = n1479 ^ n1087 ;
  assign n1483 = n1482 ^ n1480 ;
  assign n1486 = n1485 ^ n1483 ;
  assign n1489 = n1488 ^ n1486 ;
  assign n1492 = n1491 ^ n1489 ;
  assign n1495 = n1494 ^ n1492 ;
  assign n1510 = n812 & n1146 ;
  assign n1511 = n1510 ^ n1146 ;
  assign n1507 = ~n780 & n1140 ;
  assign n1508 = n1507 ^ n1140 ;
  assign n1504 = n709 & n1135 ;
  assign n1505 = n1504 ^ n1135 ;
  assign n1501 = n599 & n1129 ;
  assign n1502 = n1501 ^ n1129 ;
  assign n1498 = n452 & n1124 ;
  assign n1499 = n1498 ^ n1124 ;
  assign n1496 = n265 & n1119 ;
  assign n1497 = n1496 ^ n1119 ;
  assign n1500 = n1499 ^ n1497 ;
  assign n1503 = n1502 ^ n1500 ;
  assign n1506 = n1505 ^ n1503 ;
  assign n1509 = n1508 ^ n1506 ;
  assign n1512 = n1511 ^ n1509 ;
  assign n1527 = n812 & n1178 ;
  assign n1528 = n1527 ^ n1178 ;
  assign n1524 = ~n780 & n1172 ;
  assign n1525 = n1524 ^ n1172 ;
  assign n1521 = n709 & n1167 ;
  assign n1522 = n1521 ^ n1167 ;
  assign n1518 = n599 & n1161 ;
  assign n1519 = n1518 ^ n1161 ;
  assign n1515 = n452 & n1156 ;
  assign n1516 = n1515 ^ n1156 ;
  assign n1513 = n265 & n1151 ;
  assign n1514 = n1513 ^ n1151 ;
  assign n1517 = n1516 ^ n1514 ;
  assign n1520 = n1519 ^ n1517 ;
  assign n1523 = n1522 ^ n1520 ;
  assign n1526 = n1525 ^ n1523 ;
  assign n1529 = n1528 ^ n1526 ;
  assign n1544 = n812 & n1210 ;
  assign n1545 = n1544 ^ n1210 ;
  assign n1541 = ~n780 & n1204 ;
  assign n1542 = n1541 ^ n1204 ;
  assign n1538 = n709 & n1199 ;
  assign n1539 = n1538 ^ n1199 ;
  assign n1535 = n599 & n1193 ;
  assign n1536 = n1535 ^ n1193 ;
  assign n1532 = n452 & n1188 ;
  assign n1533 = n1532 ^ n1188 ;
  assign n1530 = n265 & n1183 ;
  assign n1531 = n1530 ^ n1183 ;
  assign n1534 = n1533 ^ n1531 ;
  assign n1537 = n1536 ^ n1534 ;
  assign n1540 = n1539 ^ n1537 ;
  assign n1543 = n1542 ^ n1540 ;
  assign n1546 = n1545 ^ n1543 ;
  assign n1561 = n812 & n1242 ;
  assign n1562 = n1561 ^ n1242 ;
  assign n1558 = ~n780 & n1236 ;
  assign n1559 = n1558 ^ n1236 ;
  assign n1555 = n709 & n1231 ;
  assign n1556 = n1555 ^ n1231 ;
  assign n1552 = n599 & n1225 ;
  assign n1553 = n1552 ^ n1225 ;
  assign n1549 = n452 & n1220 ;
  assign n1550 = n1549 ^ n1220 ;
  assign n1547 = n265 & n1215 ;
  assign n1548 = n1547 ^ n1215 ;
  assign n1551 = n1550 ^ n1548 ;
  assign n1554 = n1553 ^ n1551 ;
  assign n1557 = n1556 ^ n1554 ;
  assign n1560 = n1559 ^ n1557 ;
  assign n1563 = n1562 ^ n1560 ;
  assign n1578 = n812 & n1274 ;
  assign n1579 = n1578 ^ n1274 ;
  assign n1575 = ~n780 & n1268 ;
  assign n1576 = n1575 ^ n1268 ;
  assign n1572 = n709 & n1263 ;
  assign n1573 = n1572 ^ n1263 ;
  assign n1569 = n599 & n1257 ;
  assign n1570 = n1569 ^ n1257 ;
  assign n1566 = n452 & n1252 ;
  assign n1567 = n1566 ^ n1252 ;
  assign n1564 = n265 & n1247 ;
  assign n1565 = n1564 ^ n1247 ;
  assign n1568 = n1567 ^ n1565 ;
  assign n1571 = n1570 ^ n1568 ;
  assign n1574 = n1573 ^ n1571 ;
  assign n1577 = n1576 ^ n1574 ;
  assign n1580 = n1579 ^ n1577 ;
  assign n1595 = n812 & n1306 ;
  assign n1596 = n1595 ^ n1306 ;
  assign n1592 = ~n780 & n1300 ;
  assign n1593 = n1592 ^ n1300 ;
  assign n1589 = n709 & n1295 ;
  assign n1590 = n1589 ^ n1295 ;
  assign n1586 = n599 & n1289 ;
  assign n1587 = n1586 ^ n1289 ;
  assign n1583 = n452 & n1284 ;
  assign n1584 = n1583 ^ n1284 ;
  assign n1581 = n265 & n1279 ;
  assign n1582 = n1581 ^ n1279 ;
  assign n1585 = n1584 ^ n1582 ;
  assign n1588 = n1587 ^ n1585 ;
  assign n1591 = n1590 ^ n1588 ;
  assign n1594 = n1593 ^ n1591 ;
  assign n1597 = n1596 ^ n1594 ;
  assign n1612 = n812 & n1338 ;
  assign n1613 = n1612 ^ n1338 ;
  assign n1609 = ~n780 & n1332 ;
  assign n1610 = n1609 ^ n1332 ;
  assign n1606 = n709 & n1327 ;
  assign n1607 = n1606 ^ n1327 ;
  assign n1603 = n599 & n1321 ;
  assign n1604 = n1603 ^ n1321 ;
  assign n1600 = n452 & n1316 ;
  assign n1601 = n1600 ^ n1316 ;
  assign n1598 = n265 & n1311 ;
  assign n1599 = n1598 ^ n1311 ;
  assign n1602 = n1601 ^ n1599 ;
  assign n1605 = n1604 ^ n1602 ;
  assign n1608 = n1607 ^ n1605 ;
  assign n1611 = n1610 ^ n1608 ;
  assign n1614 = n1613 ^ n1611 ;
  assign n1615 = n458 ^ n272 ;
  assign n1616 = n1615 ^ n606 ;
  assign n1617 = n1616 ^ n715 ;
  assign n1618 = n1617 ^ n787 ;
  assign n1619 = n1618 ^ n818 ;
  assign n1620 = n830 ^ n825 ;
  assign n1621 = n1620 ^ n837 ;
  assign n1622 = n1621 ^ n843 ;
  assign n1623 = n1622 ^ n850 ;
  assign n1624 = n1623 ^ n856 ;
  assign n1625 = n868 ^ n863 ;
  assign n1626 = n1625 ^ n875 ;
  assign n1627 = n1626 ^ n881 ;
  assign n1628 = n1627 ^ n888 ;
  assign n1629 = n1628 ^ n894 ;
  assign n1630 = n906 ^ n901 ;
  assign n1631 = n1630 ^ n913 ;
  assign n1632 = n1631 ^ n919 ;
  assign n1633 = n1632 ^ n926 ;
  assign n1634 = n1633 ^ n932 ;
  assign n1635 = n944 ^ n939 ;
  assign n1636 = n1635 ^ n951 ;
  assign n1637 = n1636 ^ n957 ;
  assign n1638 = n1637 ^ n964 ;
  assign n1639 = n1638 ^ n970 ;
  assign n1640 = n982 ^ n977 ;
  assign n1641 = n1640 ^ n989 ;
  assign n1642 = n1641 ^ n995 ;
  assign n1643 = n1642 ^ n1002 ;
  assign n1644 = n1643 ^ n1008 ;
  assign n1645 = n1020 ^ n1015 ;
  assign n1646 = n1645 ^ n1027 ;
  assign n1647 = n1646 ^ n1033 ;
  assign n1648 = n1647 ^ n1040 ;
  assign n1649 = n1648 ^ n1046 ;
  assign n1650 = n1058 ^ n1053 ;
  assign n1651 = n1650 ^ n1065 ;
  assign n1652 = n1651 ^ n1071 ;
  assign n1653 = n1652 ^ n1078 ;
  assign n1654 = n1653 ^ n1084 ;
  assign n1655 = n1094 ^ n1089 ;
  assign n1656 = n1655 ^ n1099 ;
  assign n1657 = n1656 ^ n1105 ;
  assign n1658 = n1657 ^ n1110 ;
  assign n1659 = n1658 ^ n1116 ;
  assign n1660 = n1126 ^ n1121 ;
  assign n1661 = n1660 ^ n1131 ;
  assign n1662 = n1661 ^ n1137 ;
  assign n1663 = n1662 ^ n1142 ;
  assign n1664 = n1663 ^ n1148 ;
  assign n1665 = n1158 ^ n1153 ;
  assign n1666 = n1665 ^ n1163 ;
  assign n1667 = n1666 ^ n1169 ;
  assign n1668 = n1667 ^ n1174 ;
  assign n1669 = n1668 ^ n1180 ;
  assign n1670 = n1190 ^ n1185 ;
  assign n1671 = n1670 ^ n1195 ;
  assign n1672 = n1671 ^ n1201 ;
  assign n1673 = n1672 ^ n1206 ;
  assign n1674 = n1673 ^ n1212 ;
  assign n1675 = n1222 ^ n1217 ;
  assign n1676 = n1675 ^ n1227 ;
  assign n1677 = n1676 ^ n1233 ;
  assign n1678 = n1677 ^ n1238 ;
  assign n1679 = n1678 ^ n1244 ;
  assign n1680 = n1254 ^ n1249 ;
  assign n1681 = n1680 ^ n1259 ;
  assign n1682 = n1681 ^ n1265 ;
  assign n1683 = n1682 ^ n1270 ;
  assign n1684 = n1683 ^ n1276 ;
  assign n1685 = n1286 ^ n1281 ;
  assign n1686 = n1685 ^ n1291 ;
  assign n1687 = n1686 ^ n1297 ;
  assign n1688 = n1687 ^ n1302 ;
  assign n1689 = n1688 ^ n1308 ;
  assign n1690 = n1318 ^ n1313 ;
  assign n1691 = n1690 ^ n1323 ;
  assign n1692 = n1691 ^ n1329 ;
  assign n1693 = n1692 ^ n1334 ;
  assign n1694 = n1693 ^ n1340 ;
  assign y0 = n820 ;
  assign y1 = n858 ;
  assign y2 = n896 ;
  assign y3 = n934 ;
  assign y4 = n972 ;
  assign y5 = n1010 ;
  assign y6 = n1048 ;
  assign y7 = n1086 ;
  assign y8 = n1118 ;
  assign y9 = n1150 ;
  assign y10 = n1182 ;
  assign y11 = n1214 ;
  assign y12 = n1246 ;
  assign y13 = n1278 ;
  assign y14 = n1310 ;
  assign y15 = n1342 ;
  assign y16 = n1359 ;
  assign y17 = n1376 ;
  assign y18 = n1393 ;
  assign y19 = n1410 ;
  assign y20 = n1427 ;
  assign y21 = n1444 ;
  assign y22 = n1461 ;
  assign y23 = n1478 ;
  assign y24 = n1495 ;
  assign y25 = n1512 ;
  assign y26 = n1529 ;
  assign y27 = n1546 ;
  assign y28 = n1563 ;
  assign y29 = n1580 ;
  assign y30 = n1597 ;
  assign y31 = n1614 ;
  assign y32 = n1619 ;
  assign y33 = n1624 ;
  assign y34 = n1629 ;
  assign y35 = n1634 ;
  assign y36 = n1639 ;
  assign y37 = n1644 ;
  assign y38 = n1649 ;
  assign y39 = n1654 ;
  assign y40 = n1659 ;
  assign y41 = n1664 ;
  assign y42 = n1669 ;
  assign y43 = n1674 ;
  assign y44 = n1679 ;
  assign y45 = n1684 ;
  assign y46 = n1689 ;
  assign y47 = n1694 ;
endmodule
