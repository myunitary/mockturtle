module bitonic_sort_inc_1_8 (in_array_0, in_array_1, in_array_2, in_array_3, in_array_4, in_array_5, in_array_6, in_array_7, out_array_0, out_array_1, out_array_2, out_array_3, out_array_4, out_array_5, out_array_6, out_array_7);
input in_array_0, in_array_1, in_array_2, in_array_3, in_array_4, in_array_5, in_array_6, in_array_7;
output out_array_0, out_array_1, out_array_2, out_array_3, out_array_4, out_array_5, out_array_6, out_array_7;
wire _000_, _001_, _002_, _003_, _004_, _005_, _005__neg, _006_, _006__neg, _007_, _008_, _008__neg, _009_, _009__neg, _010_, _011_, _011__neg, _012_, _013_, _014_, _015_, _016_, _017_, _017__neg, _018_, _019_, _020_, _021_, _022_, _023_, _024_, _024__neg, _025_, _026_, _027_, _028_, _029_, _030_, _030__neg, _031_, _031__neg, _032_, _033_, _034_, _035_, _036_, _037_, _038_, _039_, _040_, _041_, _042_, _043_, _044_, _045_, _046_, _047_, _048_, _049_, _050_, _051_, _052_, _053_, _054_, _055_, _056_, _057_, _058_, _058__neg, _059_, _059__neg, _060_, _061_, _062_, _063_, _064_, _065_, _066_, _066__neg, _067_, _067__neg, _068_, _069_, _070_, _070__neg, _071_, _071__neg, _072_, _073_, _074_, _075_, _076_, _076__neg, _077_, _078_, _079_, _079__neg, _080_, _081_, _082_, _082__neg, _083_, _084_, _085_, _086_, _087_, out_array_1_neg, out_array_5_neg;
assign _009__neg = in_array_1 | in_array_0;
assign _009_ = ~_009__neg;
assign _010_ = in_array_3 & in_array_2;
assign _011__neg = _010_ | _009_;
assign _011_ = ~_011__neg;
assign _012_ = _011_ ^ _009_;
assign _013_ = ~_009_;
assign _014_ = _011_ ^ _013_;
assign _015_ = in_array_1 & in_array_0;
assign _016_ = ~_015_;
assign _017__neg = in_array_3 | in_array_2;
assign _017_ = ~_017__neg;
assign _018_ = _017_ & _015_;
assign _019_ = _018_ ^ _016_;
assign _020_ = _019_ & _014_;
assign _021_ = _020_ ^ _012_;
assign _022_ = _018_ ^ _015_;
assign _023_ = _022_ & _014_;
assign _024__neg = in_array_5 | in_array_4;
assign _024_ = ~_024__neg;
assign _025_ = in_array_7 & in_array_6;
assign _026_ = _025_ & _024_;
assign _027_ = _026_ ^ _024_;
assign _028_ = in_array_5 & in_array_4;
assign _029_ = ~_028_;
assign _030__neg = in_array_7 | in_array_6;
assign _030_ = ~_030__neg;
assign _031__neg = _030_ | _028_;
assign _031_ = ~_031__neg;
assign _032_ = _031_ ^ _029_;
assign _033_ = _032_ & _027_;
assign _034_ = _033_ & _023_;
assign _035_ = _034_ ^ _021_;
assign _036_ = ~_010_;
assign _037_ = _011_ ^ _036_;
assign _038_ = _011_ ^ _010_;
assign _039_ = _018_ ^ _017_;
assign _040_ = _039_ & _038_;
assign _041_ = _040_ ^ _037_;
assign _042_ = ~_017_;
assign _043_ = _018_ ^ _042_;
assign _044_ = _043_ & _038_;
assign _045_ = ~_025_;
assign _046_ = _026_ ^ _045_;
assign _047_ = _031_ ^ _030_;
assign _048_ = _047_ & _046_;
assign _049_ = _048_ & _044_;
assign _050_ = _049_ ^ _041_;
assign _051_ = _050_ & _035_;
assign _052_ = _020_ ^ _022_;
assign _053_ = _019_ & _012_;
assign _054_ = ~_024_;
assign _055_ = _026_ ^ _054_;
assign _056_ = _031_ ^ _028_;
assign _057_ = _056_ & _055_;
assign _058__neg = _057_ | _053_;
assign _058_ = ~_058__neg;
assign _059__neg = _058_ ^ _052_;
assign _059_ = ~_059__neg;
assign _060_ = _040_ ^ _043_;
assign _061_ = _039_ & _037_;
assign _062_ = _026_ ^ _025_;
assign _063_ = ~_030_;
assign _064_ = _031_ ^ _063_;
assign _065_ = _064_ & _062_;
assign _066__neg = _065_ | _061_;
assign _066_ = ~_066__neg;
assign _067__neg = _066_ ^ _060_;
assign _067_ = ~_067__neg;
assign _068_ = _067_ & _059_;
assign _069_ = _068_ & _051_;
assign out_array_4 = ~_069_;
assign _070__neg = _034_ ^ _021_;
assign _070_ = ~_070__neg;
assign _071__neg = _049_ ^ _041_;
assign _071_ = ~_071__neg;
assign _072_ = _071_ & _070_;
assign _073_ = _058_ ^ _052_;
assign _074_ = _066_ ^ _060_;
assign _075_ = _074_ & _073_;
assign _076__neg = _075_ | _072_;
assign _076_ = ~_076__neg;
assign out_array_6 = ~_076_;
assign out_array_5_neg = _068_ | _051_;
assign out_array_5 = ~out_array_5_neg;
assign out_array_7 = _075_ & _072_;
assign _077_ = _056_ & _027_;
assign _078_ = _077_ ^ _055_;
assign _079__neg = _034_ ^ _078_;
assign _079_ = ~_079__neg;
assign _080_ = _064_ & _046_;
assign _081_ = _080_ ^ _062_;
assign _082__neg = _049_ ^ _081_;
assign _082_ = ~_082__neg;
assign _083_ = _082_ & _079_;
assign _084_ = _077_ ^ _032_;
assign _085_ = _058_ ^ _084_;
assign _086_ = _080_ ^ _047_;
assign _087_ = _066_ ^ _086_;
assign _000_ = _087_ & _085_;
assign _001_ = _000_ & _083_;
assign out_array_0 = ~_001_;
assign _002_ = _034_ ^ _078_;
assign _003_ = _049_ ^ _081_;
assign _004_ = _003_ & _002_;
assign _005__neg = _058_ ^ _084_;
assign _005_ = ~_005__neg;
assign _006__neg = _066_ ^ _086_;
assign _006_ = ~_006__neg;
assign _007_ = _006_ & _005_;
assign _008__neg = _007_ | _004_;
assign _008_ = ~_008__neg;
assign out_array_2 = ~_008_;
assign out_array_1_neg = _000_ | _083_;
assign out_array_1 = ~out_array_1_neg;
assign out_array_3 = _007_ & _004_;
endmodule
