module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 ;
  assign n33 = x31 ^ x0 ;
  assign n34 = n33 ^ x31 ;
  assign n36 = x31 ^ x1 ;
  assign n35 = ~x0 & x31 ;
  assign n37 = n36 ^ n35 ;
  assign n39 = x31 ^ x2 ;
  assign n38 = n35 & n36 ;
  assign n40 = n39 ^ n38 ;
  assign n42 = x31 ^ x3 ;
  assign n41 = n38 & n39 ;
  assign n43 = n42 ^ n41 ;
  assign n46 = x31 ^ x4 ;
  assign n44 = n39 & n42 ;
  assign n45 = n38 & n44 ;
  assign n47 = n46 ^ n45 ;
  assign n49 = x31 ^ x5 ;
  assign n48 = n45 & n46 ;
  assign n50 = n49 ^ n48 ;
  assign n53 = x31 ^ x6 ;
  assign n51 = n46 & n49 ;
  assign n52 = n45 & n51 ;
  assign n54 = n53 ^ n52 ;
  assign n57 = x31 ^ x7 ;
  assign n55 = n51 & n53 ;
  assign n56 = n45 & n55 ;
  assign n58 = n57 ^ n56 ;
  assign n62 = x31 ^ x8 ;
  assign n59 = n53 & n57 ;
  assign n60 = n51 & n59 ;
  assign n61 = n45 & n60 ;
  assign n63 = n62 ^ n61 ;
  assign n65 = x31 ^ x9 ;
  assign n64 = n61 & n62 ;
  assign n66 = n65 ^ n64 ;
  assign n69 = x31 ^ x10 ;
  assign n67 = n62 & n65 ;
  assign n68 = n61 & n67 ;
  assign n70 = n69 ^ n68 ;
  assign n73 = x31 ^ x11 ;
  assign n71 = n67 & n69 ;
  assign n72 = n61 & n71 ;
  assign n74 = n73 ^ n72 ;
  assign n78 = x31 ^ x12 ;
  assign n75 = n69 & n73 ;
  assign n76 = n67 & n75 ;
  assign n77 = n61 & n76 ;
  assign n79 = n78 ^ n77 ;
  assign n82 = x31 ^ x13 ;
  assign n80 = n76 & n78 ;
  assign n81 = n61 & n80 ;
  assign n83 = n82 ^ n81 ;
  assign n87 = x31 ^ x14 ;
  assign n84 = n78 & n82 ;
  assign n85 = n76 & n84 ;
  assign n86 = n61 & n85 ;
  assign n88 = n87 ^ n86 ;
  assign n92 = x31 ^ x15 ;
  assign n89 = n84 & n87 ;
  assign n90 = n76 & n89 ;
  assign n91 = n61 & n90 ;
  assign n93 = n92 ^ n91 ;
  assign n98 = x31 ^ x16 ;
  assign n94 = n87 & n92 ;
  assign n95 = n84 & n94 ;
  assign n96 = n76 & n95 ;
  assign n97 = n61 & n96 ;
  assign n99 = n98 ^ n97 ;
  assign n101 = x31 ^ x17 ;
  assign n100 = n97 & n98 ;
  assign n102 = n101 ^ n100 ;
  assign n105 = x31 ^ x18 ;
  assign n103 = n98 & n101 ;
  assign n104 = n97 & n103 ;
  assign n106 = n105 ^ n104 ;
  assign n109 = x31 ^ x19 ;
  assign n107 = n103 & n105 ;
  assign n108 = n97 & n107 ;
  assign n110 = n109 ^ n108 ;
  assign n114 = x31 ^ x20 ;
  assign n111 = n105 & n109 ;
  assign n112 = n103 & n111 ;
  assign n113 = n97 & n112 ;
  assign n115 = n114 ^ n113 ;
  assign n118 = x31 ^ x21 ;
  assign n116 = n112 & n114 ;
  assign n117 = n97 & n116 ;
  assign n119 = n118 ^ n117 ;
  assign n123 = x31 ^ x22 ;
  assign n120 = n114 & n118 ;
  assign n121 = n112 & n120 ;
  assign n122 = n97 & n121 ;
  assign n124 = n123 ^ n122 ;
  assign n128 = x31 ^ x23 ;
  assign n125 = n120 & n123 ;
  assign n126 = n112 & n125 ;
  assign n127 = n97 & n126 ;
  assign n129 = n128 ^ n127 ;
  assign n134 = x31 ^ x24 ;
  assign n130 = n123 & n128 ;
  assign n131 = n120 & n130 ;
  assign n132 = n112 & n131 ;
  assign n133 = n97 & n132 ;
  assign n135 = n134 ^ n133 ;
  assign n138 = x31 ^ x25 ;
  assign n136 = n132 & n134 ;
  assign n137 = n97 & n136 ;
  assign n139 = n138 ^ n137 ;
  assign n143 = x31 ^ x26 ;
  assign n140 = n134 & n138 ;
  assign n141 = n132 & n140 ;
  assign n142 = n97 & n141 ;
  assign n144 = n143 ^ n142 ;
  assign n148 = x31 ^ x27 ;
  assign n145 = n140 & n143 ;
  assign n146 = n132 & n145 ;
  assign n147 = n97 & n146 ;
  assign n149 = n148 ^ n147 ;
  assign n154 = x31 ^ x28 ;
  assign n150 = n143 & n148 ;
  assign n151 = n140 & n150 ;
  assign n152 = n132 & n151 ;
  assign n153 = n97 & n152 ;
  assign n155 = n154 ^ n153 ;
  assign n159 = x31 ^ x29 ;
  assign n156 = n151 & n154 ;
  assign n157 = n132 & n156 ;
  assign n158 = n97 & n157 ;
  assign n160 = n159 ^ n158 ;
  assign n165 = x31 ^ x30 ;
  assign n161 = n154 & n159 ;
  assign n162 = n151 & n161 ;
  assign n163 = n132 & n162 ;
  assign n164 = n97 & n163 ;
  assign n166 = n165 ^ n164 ;
  assign n167 = n161 & n165 ;
  assign n168 = n151 & n167 ;
  assign n169 = n132 & n168 ;
  assign n170 = n97 & n169 ;
  assign y0 = n34 ;
  assign y1 = n37 ;
  assign y2 = n40 ;
  assign y3 = n43 ;
  assign y4 = n47 ;
  assign y5 = n50 ;
  assign y6 = n54 ;
  assign y7 = n58 ;
  assign y8 = n63 ;
  assign y9 = n66 ;
  assign y10 = n70 ;
  assign y11 = n74 ;
  assign y12 = n79 ;
  assign y13 = n83 ;
  assign y14 = n88 ;
  assign y15 = n93 ;
  assign y16 = n99 ;
  assign y17 = n102 ;
  assign y18 = n106 ;
  assign y19 = n110 ;
  assign y20 = n115 ;
  assign y21 = n119 ;
  assign y22 = n124 ;
  assign y23 = n129 ;
  assign y24 = n135 ;
  assign y25 = n139 ;
  assign y26 = n144 ;
  assign y27 = n149 ;
  assign y28 = n155 ;
  assign y29 = n160 ;
  assign y30 = n166 ;
  assign y31 = n170 ;
endmodule
