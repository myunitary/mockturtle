module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 ;
  assign n148 = ~x4 & ~x19 ;
  assign n149 = ~x18 & n148 ;
  assign n150 = ~x16 & n149 ;
  assign n151 = ~x9 & ~x11 ;
  assign n152 = ~x7 & ~x13 ;
  assign n153 = ~x14 & ~x22 ;
  assign n154 = n152 & n153 ;
  assign n155 = n151 & n154 ;
  assign n156 = ~x17 & ~x21 ;
  assign n157 = ~x8 & n156 ;
  assign n158 = ~x6 & ~x12 ;
  assign n159 = ~x5 & n158 ;
  assign n160 = n157 & n159 ;
  assign n161 = n155 & n160 ;
  assign n162 = n150 & n161 ;
  assign n163 = x54 & ~n162 ;
  assign n164 = ~x0 & ~n163 ;
  assign n165 = ~x5 & ~x22 ;
  assign n168 = ~x56 & ~n151 ;
  assign n169 = n165 & n168 ;
  assign n172 = n169 ^ n151 ;
  assign n212 = n172 ^ x54 ;
  assign n181 = x21 ^ x13 ;
  assign n179 = x21 ^ x8 ;
  assign n178 = x21 ^ x7 ;
  assign n180 = n179 ^ n178 ;
  assign n182 = n181 ^ n180 ;
  assign n183 = n179 ^ x21 ;
  assign n184 = n183 ^ x21 ;
  assign n185 = n181 ^ x21 ;
  assign n186 = n185 ^ n183 ;
  assign n187 = n184 & n186 ;
  assign n188 = n187 ^ n183 ;
  assign n189 = n182 & n188 ;
  assign n190 = n189 ^ n182 ;
  assign n192 = n190 ^ x14 ;
  assign n176 = x14 ^ x10 ;
  assign n177 = n176 ^ x14 ;
  assign n191 = n190 ^ n177 ;
  assign n193 = n192 ^ n191 ;
  assign n195 = x8 & x21 ;
  assign n196 = n195 ^ x8 ;
  assign n197 = n196 ^ x21 ;
  assign n198 = n152 & ~n197 ;
  assign n194 = n190 & n191 ;
  assign n199 = n198 ^ n194 ;
  assign n200 = n193 & n199 ;
  assign n201 = n200 ^ n194 ;
  assign n202 = ~x17 & n158 ;
  assign n203 = n165 & n202 ;
  assign n204 = n150 & n203 ;
  assign n205 = ~n201 & n204 ;
  assign n206 = n205 ^ n204 ;
  assign n166 = ~x56 & ~n165 ;
  assign n173 = n169 ^ n166 ;
  assign n174 = ~n172 & n173 ;
  assign n175 = n174 ^ n166 ;
  assign n207 = n206 ^ n175 ;
  assign n213 = n212 ^ n207 ;
  assign n214 = n206 ^ n151 ;
  assign n215 = n214 ^ n175 ;
  assign n216 = ~n213 & n215 ;
  assign n208 = n175 ^ n151 ;
  assign n170 = n169 ^ x54 ;
  assign n209 = n208 ^ n170 ;
  assign n210 = n207 & n209 ;
  assign n217 = n216 ^ n210 ;
  assign n218 = n217 ^ n175 ;
  assign n219 = n218 ^ n212 ;
  assign n220 = n210 ^ n206 ;
  assign n221 = n220 ^ x54 ;
  assign n222 = n219 & ~n221 ;
  assign n223 = n222 ^ n216 ;
  assign n211 = n210 ^ n174 ;
  assign n224 = n223 ^ n211 ;
  assign n167 = n166 ^ n151 ;
  assign n171 = n170 ^ n167 ;
  assign n225 = n224 ^ n171 ;
  assign n226 = n225 ^ x54 ;
  assign n227 = n164 & n226 ;
  assign n228 = n227 ^ n164 ;
  assign n229 = n228 ^ n226 ;
  assign n230 = ~x3 & ~x129 ;
  assign n231 = ~n229 & n230 ;
  assign n232 = n231 ^ n230 ;
  assign n233 = ~x17 & x54 ;
  assign n234 = ~x5 & ~x6 ;
  assign n235 = n152 & n234 ;
  assign n236 = n150 & n235 ;
  assign n237 = ~x14 & ~n197 ;
  assign n238 = ~x11 & ~x12 ;
  assign n239 = ~x10 & ~x22 ;
  assign n240 = n238 & n239 ;
  assign n241 = n237 & n240 ;
  assign n242 = n236 & n241 ;
  assign n243 = n233 & ~n242 ;
  assign n244 = ~x1 & ~n243 ;
  assign n245 = ~x7 & ~x12 ;
  assign n246 = ~n234 & ~n245 ;
  assign n247 = ~x13 & ~n246 ;
  assign n248 = ~x5 & ~x7 ;
  assign n249 = n248 ^ n158 ;
  assign n250 = n247 & n249 ;
  assign n251 = x13 & n158 ;
  assign n252 = n248 & n251 ;
  assign n253 = ~x9 & ~n252 ;
  assign n254 = ~n250 & n253 ;
  assign n255 = n152 & n159 ;
  assign n256 = x9 & ~n255 ;
  assign n257 = ~x10 & x54 ;
  assign n258 = n153 & n257 ;
  assign n259 = ~x8 & ~x11 ;
  assign n260 = n156 & n259 ;
  assign n261 = n258 & n260 ;
  assign n262 = n150 & n261 ;
  assign n263 = ~n256 & n262 ;
  assign n264 = ~n254 & n263 ;
  assign n265 = ~n244 & ~n264 ;
  assign n266 = n230 & ~n265 ;
  assign n269 = x42 & x44 ;
  assign n270 = n269 ^ x42 ;
  assign n271 = n270 ^ x44 ;
  assign n272 = x40 & ~n271 ;
  assign n273 = n272 ^ n271 ;
  assign n274 = x24 & x49 ;
  assign n275 = n274 ^ x24 ;
  assign n276 = n275 ^ x49 ;
  assign n277 = x15 & x20 ;
  assign n278 = n277 ^ x15 ;
  assign n279 = n278 ^ x20 ;
  assign n280 = x45 & n279 ;
  assign n281 = n280 ^ x45 ;
  assign n282 = n281 ^ n279 ;
  assign n283 = n276 & ~n282 ;
  assign n284 = n283 ^ n282 ;
  assign n285 = x43 & x47 ;
  assign n286 = n285 ^ x43 ;
  assign n287 = n286 ^ x47 ;
  assign n288 = ~x2 & ~x48 ;
  assign n289 = ~n287 & n288 ;
  assign n290 = x38 & x50 ;
  assign n291 = n290 ^ x38 ;
  assign n292 = n291 ^ x50 ;
  assign n293 = ~x41 & ~x46 ;
  assign n294 = ~n292 & n293 ;
  assign n295 = n294 ^ n289 ;
  assign n296 = ~n289 & n295 ;
  assign n297 = n296 ^ n294 ;
  assign n298 = n297 ^ n284 ;
  assign n299 = n284 & ~n298 ;
  assign n300 = n299 ^ n296 ;
  assign n301 = n300 ^ n294 ;
  assign n302 = ~n273 & n301 ;
  assign n303 = x82 & ~n302 ;
  assign n267 = x122 & x127 ;
  assign n268 = ~x65 & ~n267 ;
  assign n304 = n303 ^ n268 ;
  assign n305 = ~x40 & ~x46 ;
  assign n306 = ~n292 & n305 ;
  assign n307 = ~x41 & ~x43 ;
  assign n308 = ~n271 & n307 ;
  assign n309 = n306 & n308 ;
  assign n310 = ~x47 & ~x48 ;
  assign n311 = n309 & n310 ;
  assign n312 = x82 & ~n284 ;
  assign n313 = n311 & n312 ;
  assign n314 = ~x82 & ~n267 ;
  assign n315 = x2 & ~n314 ;
  assign n316 = n313 & n315 ;
  assign n317 = n316 ^ n315 ;
  assign n318 = n317 ^ n268 ;
  assign n319 = n317 & n318 ;
  assign n320 = n319 ^ n317 ;
  assign n321 = n320 ^ n303 ;
  assign n322 = ~n304 & ~n321 ;
  assign n323 = n322 ^ n319 ;
  assign n324 = n323 ^ n303 ;
  assign n325 = x129 & n324 ;
  assign n326 = n325 ^ x129 ;
  assign n327 = n326 ^ n324 ;
  assign n328 = x0 & ~x113 ;
  assign n329 = ~x123 & n328 ;
  assign n330 = ~x9 & ~x14 ;
  assign n331 = n239 & n330 ;
  assign n332 = ~x12 & n260 ;
  assign n333 = n331 & n332 ;
  assign n334 = n236 & n333 ;
  assign n335 = ~x61 & ~x118 ;
  assign n336 = ~n334 & n335 ;
  assign n337 = ~n329 & ~n336 ;
  assign n338 = ~x129 & ~n337 ;
  assign n339 = x4 & ~x54 ;
  assign n340 = n255 & n330 ;
  assign n341 = ~x16 & x54 ;
  assign n342 = n156 & n341 ;
  assign n343 = n149 & n342 ;
  assign n344 = n259 & n343 ;
  assign n345 = x10 & ~x22 ;
  assign n346 = n344 & n345 ;
  assign n347 = n340 & n346 ;
  assign n348 = ~n339 & ~n347 ;
  assign n349 = n230 & ~n348 ;
  assign n350 = x5 & ~x54 ;
  assign n351 = ~x13 & n331 ;
  assign n352 = ~x59 & n260 ;
  assign n353 = n351 & n352 ;
  assign n354 = n158 & n248 ;
  assign n355 = n341 & n354 ;
  assign n356 = ~x25 & x28 ;
  assign n357 = ~x29 & n356 ;
  assign n358 = n149 & n357 ;
  assign n359 = n355 & n358 ;
  assign n360 = n353 & n359 ;
  assign n361 = ~n350 & ~n360 ;
  assign n362 = n230 & ~n361 ;
  assign n363 = x6 & ~x54 ;
  assign n364 = ~x28 & ~x29 ;
  assign n365 = x25 & n364 ;
  assign n366 = n149 & n365 ;
  assign n367 = n355 & n366 ;
  assign n368 = n353 & n367 ;
  assign n369 = ~n363 & ~n368 ;
  assign n370 = n230 & ~n369 ;
  assign n371 = x7 & ~x54 ;
  assign n372 = x8 & n343 ;
  assign n373 = ~x11 & n354 ;
  assign n374 = n351 & n373 ;
  assign n375 = n372 & n374 ;
  assign n376 = ~n371 & ~n375 ;
  assign n377 = n230 & ~n376 ;
  assign n378 = x8 & ~x54 ;
  assign n379 = ~x12 & n331 ;
  assign n380 = n235 & n379 ;
  assign n381 = n148 & n341 ;
  assign n382 = ~x17 & ~x18 ;
  assign n383 = n259 & n382 ;
  assign n384 = x21 & n383 ;
  assign n385 = n381 & n384 ;
  assign n386 = n380 & n385 ;
  assign n387 = ~n378 & ~n386 ;
  assign n388 = n230 & ~n387 ;
  assign n389 = x9 & ~x54 ;
  assign n390 = ~x8 & n343 ;
  assign n391 = x11 & n354 ;
  assign n392 = n351 & n391 ;
  assign n393 = n390 & n392 ;
  assign n394 = ~n389 & ~n393 ;
  assign n395 = n230 & ~n394 ;
  assign n396 = x10 & ~x54 ;
  assign n397 = ~x9 & ~x18 ;
  assign n398 = n157 & n397 ;
  assign n399 = n239 & n398 ;
  assign n400 = ~x13 & x14 ;
  assign n401 = n381 & n400 ;
  assign n402 = n373 & n401 ;
  assign n403 = n399 & n402 ;
  assign n404 = ~n396 & ~n403 ;
  assign n405 = n230 & ~n404 ;
  assign n406 = x11 & ~x54 ;
  assign n407 = ~x10 & ~x11 ;
  assign n408 = x22 & n407 ;
  assign n409 = n340 & n408 ;
  assign n410 = n390 & n409 ;
  assign n411 = ~n406 & ~n410 ;
  assign n412 = n230 & ~n411 ;
  assign n413 = x12 & ~x54 ;
  assign n414 = x18 & n235 ;
  assign n415 = n331 & n381 ;
  assign n416 = n414 & n415 ;
  assign n417 = n332 & n416 ;
  assign n418 = ~n413 & ~n417 ;
  assign n419 = n230 & ~n418 ;
  assign n420 = x13 & ~x54 ;
  assign n421 = ~x25 & ~x28 ;
  assign n422 = x29 & n421 ;
  assign n423 = ~x59 & n239 ;
  assign n424 = n422 & n423 ;
  assign n425 = n344 & n424 ;
  assign n426 = n340 & n425 ;
  assign n427 = ~n420 & ~n426 ;
  assign n428 = n230 & ~n427 ;
  assign n429 = x14 & ~x54 ;
  assign n430 = x13 & ~x16 ;
  assign n431 = n148 & n430 ;
  assign n432 = n258 & n431 ;
  assign n433 = n373 & n432 ;
  assign n434 = n398 & n433 ;
  assign n435 = ~n429 & ~n434 ;
  assign n436 = n230 & ~n435 ;
  assign n437 = ~n273 & n294 ;
  assign n438 = x48 & ~n287 ;
  assign n439 = n438 ^ n287 ;
  assign n440 = x45 & ~n276 ;
  assign n441 = n440 ^ n276 ;
  assign n442 = ~n439 & ~n441 ;
  assign n443 = n437 & n442 ;
  assign n444 = x15 & ~n443 ;
  assign n445 = ~x15 & ~n276 ;
  assign n446 = ~x45 & n310 ;
  assign n447 = ~x2 & ~x20 ;
  assign n448 = n446 & ~n447 ;
  assign n449 = n445 & n448 ;
  assign n450 = n309 & n449 ;
  assign n451 = ~n444 & ~n450 ;
  assign n452 = x82 & ~n451 ;
  assign n453 = ~x82 & n267 ;
  assign n454 = x15 & n453 ;
  assign n455 = n271 & n306 ;
  assign n456 = n455 ^ n306 ;
  assign n457 = ~x15 & n307 ;
  assign n458 = n310 & n457 ;
  assign n459 = ~n441 & n458 ;
  assign n460 = n456 & n459 ;
  assign n461 = x82 & ~n460 ;
  assign n462 = ~x70 & ~n267 ;
  assign n463 = ~n461 & n462 ;
  assign n464 = ~n454 & ~n463 ;
  assign n465 = ~n452 & n464 ;
  assign n466 = ~x129 & ~n465 ;
  assign n467 = x16 & ~x54 ;
  assign n468 = x6 & ~x13 ;
  assign n469 = n248 & n468 ;
  assign n470 = n379 & n469 ;
  assign n471 = n344 & n470 ;
  assign n472 = ~n467 & ~n471 ;
  assign n473 = n230 & ~n472 ;
  assign n474 = x17 & ~x54 ;
  assign n475 = ~x25 & x59 ;
  assign n476 = ~n197 & n475 ;
  assign n477 = n233 & n364 ;
  assign n478 = n476 & n477 ;
  assign n479 = n150 & n478 ;
  assign n480 = n374 & n479 ;
  assign n481 = ~n474 & ~n480 ;
  assign n482 = n230 & ~n481 ;
  assign n483 = x18 & ~x54 ;
  assign n484 = n149 & n380 ;
  assign n485 = x16 & x54 ;
  assign n486 = n260 & n485 ;
  assign n487 = n484 & n486 ;
  assign n488 = ~n483 & ~n487 ;
  assign n489 = n230 & ~n488 ;
  assign n490 = x19 & ~x54 ;
  assign n491 = x17 & ~x21 ;
  assign n492 = n259 & n491 ;
  assign n493 = n341 & n492 ;
  assign n494 = n484 & n493 ;
  assign n495 = ~n490 & ~n494 ;
  assign n496 = n230 & ~n495 ;
  assign n506 = ~x46 & ~x50 ;
  assign n507 = ~x38 & ~x40 ;
  assign n508 = ~n271 & n507 ;
  assign n509 = n506 & n508 ;
  assign n510 = ~x45 & n307 ;
  assign n511 = ~n276 & n310 ;
  assign n512 = n510 & n511 ;
  assign n513 = n509 & n512 ;
  assign n534 = x2 & ~n279 ;
  assign n535 = n513 & n534 ;
  assign n536 = ~x15 & x20 ;
  assign n537 = n513 & n536 ;
  assign n538 = n537 ^ x20 ;
  assign n539 = n535 & n538 ;
  assign n540 = n539 ^ n535 ;
  assign n541 = n540 ^ n538 ;
  assign n542 = x82 & ~n541 ;
  assign n543 = n542 ^ x82 ;
  assign n499 = ~x71 & ~n267 ;
  assign n502 = n499 ^ x82 ;
  assign n498 = x20 & n453 ;
  assign n519 = n502 ^ n498 ;
  assign n503 = n499 ^ n279 ;
  assign n504 = n502 & ~n503 ;
  assign n505 = n504 ^ n279 ;
  assign n514 = n513 ^ n505 ;
  assign n520 = n519 ^ n514 ;
  assign n521 = n513 ^ x82 ;
  assign n522 = n521 ^ n505 ;
  assign n523 = n520 & ~n522 ;
  assign n515 = n505 ^ x82 ;
  assign n500 = n499 ^ n498 ;
  assign n516 = n515 ^ n500 ;
  assign n517 = ~n514 & n516 ;
  assign n524 = n523 ^ n517 ;
  assign n525 = n524 ^ n505 ;
  assign n526 = n525 ^ n519 ;
  assign n527 = n517 ^ n513 ;
  assign n528 = n527 ^ n498 ;
  assign n529 = n526 & ~n528 ;
  assign n530 = n529 ^ n523 ;
  assign n518 = n517 ^ n504 ;
  assign n531 = n530 ^ n518 ;
  assign n497 = n279 ^ x82 ;
  assign n501 = n500 ^ n497 ;
  assign n532 = n531 ^ n501 ;
  assign n533 = n532 ^ n498 ;
  assign n544 = n543 ^ n533 ;
  assign n545 = n533 ^ x129 ;
  assign n546 = x129 & ~n545 ;
  assign n547 = n546 ^ x129 ;
  assign n548 = n547 ^ n543 ;
  assign n549 = n544 & ~n548 ;
  assign n550 = n549 ^ n546 ;
  assign n551 = n550 ^ n543 ;
  assign n552 = x21 & ~x54 ;
  assign n553 = ~x4 & x19 ;
  assign n554 = ~x21 & n553 ;
  assign n555 = n341 & n554 ;
  assign n556 = n383 & n555 ;
  assign n557 = n380 & n556 ;
  assign n558 = ~n552 & ~n557 ;
  assign n559 = n230 & ~n558 ;
  assign n560 = x22 & ~x54 ;
  assign n561 = x5 & ~x6 ;
  assign n562 = ~x14 & n561 ;
  assign n563 = n152 & n238 ;
  assign n564 = n562 & n563 ;
  assign n565 = n381 & n564 ;
  assign n566 = n399 & n565 ;
  assign n567 = ~n560 & ~n566 ;
  assign n568 = n230 & ~n567 ;
  assign n569 = ~x23 & x55 ;
  assign n570 = x61 & ~x129 ;
  assign n571 = ~n569 & n570 ;
  assign n577 = n307 & n446 ;
  assign n578 = n509 & n577 ;
  assign n579 = x24 & x82 ;
  assign n580 = n578 & n579 ;
  assign n581 = ~x129 & ~n580 ;
  assign n597 = n581 ^ x24 ;
  assign n572 = n534 ^ n279 ;
  assign n582 = ~x45 & ~x49 ;
  assign n583 = ~n572 & n582 ;
  assign n584 = n583 ^ n311 ;
  assign n585 = n583 ^ x82 ;
  assign n586 = ~x82 & ~n585 ;
  assign n587 = n586 ^ x82 ;
  assign n588 = n587 ^ n311 ;
  assign n589 = n584 & ~n588 ;
  assign n590 = n589 ^ n586 ;
  assign n591 = n590 ^ n311 ;
  assign n592 = x63 & ~n267 ;
  assign n593 = ~n591 & n592 ;
  assign n594 = n593 ^ n592 ;
  assign n608 = n597 ^ n594 ;
  assign n601 = n456 & n577 ;
  assign n602 = x82 & ~n601 ;
  assign n573 = ~x49 & ~n572 ;
  assign n574 = x82 & ~n573 ;
  assign n575 = n267 & ~n574 ;
  assign n598 = n581 ^ n575 ;
  assign n599 = ~n597 & ~n598 ;
  assign n600 = n599 ^ n575 ;
  assign n603 = n602 ^ n600 ;
  assign n609 = n608 ^ n603 ;
  assign n610 = n602 ^ x24 ;
  assign n611 = n610 ^ n600 ;
  assign n612 = n609 & ~n611 ;
  assign n604 = n600 ^ x24 ;
  assign n595 = n594 ^ n581 ;
  assign n605 = n604 ^ n595 ;
  assign n606 = n603 & ~n605 ;
  assign n613 = n612 ^ n606 ;
  assign n614 = n613 ^ n600 ;
  assign n615 = n614 ^ n608 ;
  assign n616 = n606 ^ n602 ;
  assign n617 = n616 ^ n594 ;
  assign n618 = ~n615 & n617 ;
  assign n619 = n618 ^ n612 ;
  assign n607 = n606 ^ n599 ;
  assign n620 = n619 ^ n607 ;
  assign n576 = n575 ^ x24 ;
  assign n596 = n595 ^ n576 ;
  assign n621 = n620 ^ n596 ;
  assign n666 = x58 ^ x53 ;
  assign n669 = n666 ^ x53 ;
  assign n659 = ~x53 & ~x58 ;
  assign n660 = ~x27 & ~x85 ;
  assign n661 = x25 & ~x116 ;
  assign n662 = ~x26 & n661 ;
  assign n663 = n660 & n662 ;
  assign n664 = ~n659 & ~n663 ;
  assign n665 = n230 & ~n664 ;
  assign n697 = n669 ^ n665 ;
  assign n642 = x39 & x52 ;
  assign n643 = n642 ^ x39 ;
  assign n644 = n643 ^ x52 ;
  assign n645 = ~x51 & x116 ;
  assign n646 = ~n644 & n645 ;
  assign n673 = ~n646 & ~n661 ;
  assign n674 = x27 & ~n673 ;
  assign n675 = x51 & x52 ;
  assign n676 = n675 ^ x51 ;
  assign n677 = n676 ^ x52 ;
  assign n678 = x39 & ~n677 ;
  assign n679 = n678 ^ n677 ;
  assign n680 = x27 & n679 ;
  assign n681 = x95 & x100 ;
  assign n682 = n681 ^ x95 ;
  assign n683 = n682 ^ x100 ;
  assign n684 = ~x97 & ~x110 ;
  assign n685 = ~n683 & n684 ;
  assign n686 = n685 ^ x110 ;
  assign n687 = x25 & n686 ;
  assign n688 = ~n680 & n687 ;
  assign n689 = ~n674 & ~n688 ;
  assign n690 = ~x26 & ~x85 ;
  assign n691 = ~n689 & n690 ;
  assign n625 = x116 ^ x110 ;
  assign n624 = x116 ^ x96 ;
  assign n626 = n625 ^ n624 ;
  assign n627 = n624 ^ x116 ;
  assign n628 = n626 & ~n627 ;
  assign n629 = n628 ^ n624 ;
  assign n630 = ~x85 & ~n629 ;
  assign n631 = n630 ^ x116 ;
  assign n632 = x100 & ~n631 ;
  assign n633 = n632 ^ x100 ;
  assign n622 = x85 & ~x116 ;
  assign n623 = x25 & n622 ;
  assign n634 = n633 ^ n623 ;
  assign n635 = n623 ^ x26 ;
  assign n636 = x26 & ~n635 ;
  assign n637 = n636 ^ x26 ;
  assign n638 = n637 ^ n633 ;
  assign n639 = n634 & ~n638 ;
  assign n640 = n639 ^ n636 ;
  assign n641 = n640 ^ n633 ;
  assign n647 = x26 & ~x85 ;
  assign n648 = ~n646 & n647 ;
  assign n649 = ~x25 & ~x116 ;
  assign n650 = n648 & n649 ;
  assign n651 = n650 ^ n648 ;
  assign n652 = n641 & n651 ;
  assign n653 = n652 ^ n641 ;
  assign n654 = n653 ^ n651 ;
  assign n655 = x27 & ~n654 ;
  assign n656 = n655 ^ x27 ;
  assign n657 = n656 ^ n654 ;
  assign n670 = n666 ^ n657 ;
  assign n671 = n669 & n670 ;
  assign n672 = n671 ^ n657 ;
  assign n692 = n691 ^ n672 ;
  assign n698 = n697 ^ n692 ;
  assign n699 = n691 ^ x53 ;
  assign n700 = n699 ^ n672 ;
  assign n701 = n698 & ~n700 ;
  assign n693 = n672 ^ x53 ;
  assign n667 = n666 ^ n665 ;
  assign n694 = n693 ^ n667 ;
  assign n695 = n692 & ~n694 ;
  assign n702 = n701 ^ n695 ;
  assign n703 = n702 ^ n672 ;
  assign n704 = n703 ^ n697 ;
  assign n705 = n695 ^ n691 ;
  assign n706 = n705 ^ n665 ;
  assign n707 = ~n704 & ~n706 ;
  assign n708 = n707 ^ n701 ;
  assign n696 = n695 ^ n671 ;
  assign n709 = n708 ^ n696 ;
  assign n658 = n657 ^ x53 ;
  assign n668 = n667 ^ n658 ;
  assign n710 = n709 ^ n668 ;
  assign n711 = n710 ^ n665 ;
  assign n712 = x26 & x116 ;
  assign n713 = n633 & ~n712 ;
  assign n714 = ~n648 & ~n713 ;
  assign n715 = ~x27 & ~x53 ;
  assign n716 = ~x58 & n715 ;
  assign n717 = n230 & n716 ;
  assign n718 = ~n714 & n717 ;
  assign n719 = x85 & n646 ;
  assign n720 = n719 ^ x85 ;
  assign n721 = n720 ^ n646 ;
  assign n722 = x27 & ~n721 ;
  assign n723 = x85 & x116 ;
  assign n724 = x85 & x110 ;
  assign n725 = n724 ^ x85 ;
  assign n726 = n725 ^ x110 ;
  assign n727 = x95 & ~x96 ;
  assign n728 = ~n726 & n727 ;
  assign n729 = ~n723 & ~n728 ;
  assign n730 = ~x27 & ~x100 ;
  assign n731 = ~n729 & n730 ;
  assign n732 = ~n722 & ~n731 ;
  assign n733 = ~x26 & n230 ;
  assign n734 = n659 & n733 ;
  assign n735 = ~n732 & n734 ;
  assign n758 = ~x27 & x28 ;
  assign n759 = ~x116 & n758 ;
  assign n760 = x53 & n690 ;
  assign n761 = n759 & n760 ;
  assign n750 = x100 & x116 ;
  assign n751 = ~x26 & ~x27 ;
  assign n752 = ~x28 & ~x116 ;
  assign n753 = n751 & ~n752 ;
  assign n754 = ~n750 & n753 ;
  assign n755 = x85 & ~n754 ;
  assign n756 = ~x53 & ~n755 ;
  assign n764 = n761 ^ n756 ;
  assign n792 = n764 ^ x58 ;
  assign n768 = ~x26 & n680 ;
  assign n769 = x116 & n768 ;
  assign n770 = x51 & n644 ;
  assign n771 = n770 ^ x51 ;
  assign n772 = n771 ^ n644 ;
  assign n773 = n712 & ~n772 ;
  assign n774 = x26 & x100 ;
  assign n775 = n774 ^ x26 ;
  assign n776 = n775 ^ x100 ;
  assign n777 = x110 & ~n776 ;
  assign n778 = n777 ^ n776 ;
  assign n779 = n727 & ~n778 ;
  assign n780 = n773 & n779 ;
  assign n781 = n780 ^ n773 ;
  assign n782 = n781 ^ n779 ;
  assign n783 = n660 & n782 ;
  assign n784 = n783 ^ x85 ;
  assign n785 = n769 & ~n784 ;
  assign n786 = n785 ^ n784 ;
  assign n736 = ~x51 & ~x52 ;
  assign n737 = x27 ^ x26 ;
  assign n738 = ~x39 & n737 ;
  assign n739 = n736 & n738 ;
  assign n740 = n739 ^ n737 ;
  assign n741 = n740 ^ x27 ;
  assign n742 = n686 & n741 ;
  assign n743 = n742 ^ n686 ;
  assign n744 = ~x116 & n737 ;
  assign n745 = n743 & n744 ;
  assign n746 = n745 ^ n743 ;
  assign n747 = n746 ^ n744 ;
  assign n748 = x28 & ~n747 ;
  assign n749 = n748 ^ x28 ;
  assign n765 = n761 ^ n749 ;
  assign n766 = ~n764 & n765 ;
  assign n767 = n766 ^ n749 ;
  assign n787 = n786 ^ n767 ;
  assign n793 = n792 ^ n787 ;
  assign n794 = n786 ^ n756 ;
  assign n795 = n794 ^ n767 ;
  assign n796 = n793 & n795 ;
  assign n788 = n767 ^ n756 ;
  assign n762 = n761 ^ x58 ;
  assign n789 = n788 ^ n762 ;
  assign n790 = n787 & ~n789 ;
  assign n797 = n796 ^ n790 ;
  assign n798 = n797 ^ n767 ;
  assign n799 = n798 ^ n792 ;
  assign n800 = n790 ^ n786 ;
  assign n801 = n800 ^ x58 ;
  assign n802 = ~n799 & n801 ;
  assign n803 = n802 ^ n796 ;
  assign n791 = n790 ^ n766 ;
  assign n804 = n803 ^ n791 ;
  assign n757 = n756 ^ n749 ;
  assign n763 = n762 ^ n757 ;
  assign n805 = n804 ^ n763 ;
  assign n806 = n805 ^ x58 ;
  assign n807 = ~x26 & ~x53 ;
  assign n808 = ~x85 & n807 ;
  assign n809 = x58 & n759 ;
  assign n810 = n808 & n809 ;
  assign n811 = n806 & n810 ;
  assign n812 = n811 ^ n806 ;
  assign n813 = n812 ^ n810 ;
  assign n814 = n230 & ~n813 ;
  assign n815 = n814 ^ n230 ;
  assign n816 = x29 & ~x116 ;
  assign n817 = x26 & ~x27 ;
  assign n818 = ~x85 & n659 ;
  assign n819 = n817 & n818 ;
  assign n820 = n816 & n819 ;
  assign n824 = n820 ^ x129 ;
  assign n894 = n824 ^ x3 ;
  assign n831 = x85 & n816 ;
  assign n832 = n716 & n831 ;
  assign n828 = x27 & n659 ;
  assign n829 = n816 & n828 ;
  assign n835 = n832 ^ n829 ;
  assign n874 = n835 ^ x85 ;
  assign n848 = x96 & x110 ;
  assign n849 = n848 ^ x96 ;
  assign n850 = n849 ^ x110 ;
  assign n851 = x97 & ~n850 ;
  assign n852 = n851 ^ x97 ;
  assign n853 = ~x110 & ~n683 ;
  assign n854 = ~n852 & n853 ;
  assign n855 = n854 ^ x110 ;
  assign n856 = x29 & ~n855 ;
  assign n857 = n856 ^ x29 ;
  assign n858 = ~x58 & x97 ;
  assign n859 = ~n683 & ~n850 ;
  assign n860 = n858 & n859 ;
  assign n861 = n860 ^ x58 ;
  assign n862 = n857 & ~n861 ;
  assign n863 = n862 ^ n861 ;
  assign n839 = x53 & ~x58 ;
  assign n840 = n816 & n839 ;
  assign n841 = x97 & x116 ;
  assign n842 = x58 & ~n816 ;
  assign n843 = ~n841 & n842 ;
  assign n844 = ~x53 & ~n843 ;
  assign n845 = n844 ^ n840 ;
  assign n846 = n840 & n845 ;
  assign n847 = n846 ^ n840 ;
  assign n864 = n863 ^ n847 ;
  assign n865 = n863 ^ n844 ;
  assign n866 = n864 & n865 ;
  assign n867 = n866 ^ n846 ;
  assign n868 = n867 ^ n863 ;
  assign n836 = n832 ^ x27 ;
  assign n837 = n835 & n836 ;
  assign n838 = n837 ^ x27 ;
  assign n869 = n868 ^ n838 ;
  assign n875 = n874 ^ n869 ;
  assign n876 = n868 ^ n829 ;
  assign n877 = n876 ^ n838 ;
  assign n878 = n875 & n877 ;
  assign n870 = n838 ^ n829 ;
  assign n833 = n832 ^ x85 ;
  assign n871 = n870 ^ n833 ;
  assign n872 = ~n869 & n871 ;
  assign n879 = n878 ^ n872 ;
  assign n880 = n879 ^ n838 ;
  assign n881 = n880 ^ n874 ;
  assign n882 = n872 ^ n868 ;
  assign n883 = n882 ^ x85 ;
  assign n884 = n881 & ~n883 ;
  assign n885 = n884 ^ n878 ;
  assign n873 = n872 ^ n837 ;
  assign n886 = n885 ^ n873 ;
  assign n830 = n829 ^ x27 ;
  assign n834 = n833 ^ n830 ;
  assign n887 = n886 ^ n834 ;
  assign n888 = n887 ^ n832 ;
  assign n825 = x129 ^ x26 ;
  assign n826 = n824 & n825 ;
  assign n827 = n826 ^ x26 ;
  assign n889 = n888 ^ n827 ;
  assign n895 = n894 ^ n889 ;
  assign n896 = n888 ^ n820 ;
  assign n897 = n896 ^ n827 ;
  assign n898 = n895 & n897 ;
  assign n890 = n827 ^ n820 ;
  assign n822 = x129 ^ x3 ;
  assign n891 = n890 ^ n822 ;
  assign n892 = ~n889 & n891 ;
  assign n899 = n898 ^ n892 ;
  assign n900 = n899 ^ n827 ;
  assign n901 = n900 ^ n894 ;
  assign n902 = n892 ^ n888 ;
  assign n903 = n902 ^ x3 ;
  assign n904 = n901 & ~n903 ;
  assign n905 = n904 ^ n898 ;
  assign n893 = n892 ^ n826 ;
  assign n906 = n905 ^ n893 ;
  assign n821 = n820 ^ x26 ;
  assign n823 = n822 ^ n821 ;
  assign n907 = n906 ^ n823 ;
  assign n908 = ~x30 & ~x109 ;
  assign n909 = ~x60 & x109 ;
  assign n910 = ~n908 & ~n909 ;
  assign n911 = ~x106 & ~n910 ;
  assign n912 = ~x88 & x106 ;
  assign n913 = ~x129 & ~n912 ;
  assign n914 = ~n911 & n913 ;
  assign n915 = ~x31 & ~x109 ;
  assign n916 = ~x30 & x109 ;
  assign n917 = ~n915 & ~n916 ;
  assign n918 = ~x106 & ~n917 ;
  assign n919 = ~x89 & x106 ;
  assign n920 = ~x129 & ~n919 ;
  assign n921 = ~n918 & n920 ;
  assign n922 = ~x32 & ~x109 ;
  assign n923 = ~x31 & x109 ;
  assign n924 = ~n922 & ~n923 ;
  assign n925 = ~x106 & ~n924 ;
  assign n926 = ~x99 & x106 ;
  assign n927 = ~x129 & ~n926 ;
  assign n928 = ~n925 & n927 ;
  assign n929 = ~x33 & ~x109 ;
  assign n930 = ~x32 & x109 ;
  assign n931 = ~n929 & ~n930 ;
  assign n932 = ~x106 & ~n931 ;
  assign n933 = ~x90 & x106 ;
  assign n934 = ~x129 & ~n933 ;
  assign n935 = ~n932 & n934 ;
  assign n936 = ~x34 & ~x109 ;
  assign n937 = ~x33 & x109 ;
  assign n938 = ~n936 & ~n937 ;
  assign n939 = ~x106 & ~n938 ;
  assign n940 = ~x91 & x106 ;
  assign n941 = ~x129 & ~n940 ;
  assign n942 = ~n939 & n941 ;
  assign n943 = ~x35 & ~x109 ;
  assign n944 = ~x34 & x109 ;
  assign n945 = ~n943 & ~n944 ;
  assign n946 = ~x106 & ~n945 ;
  assign n947 = ~x92 & x106 ;
  assign n948 = ~x129 & ~n947 ;
  assign n949 = ~n946 & n948 ;
  assign n950 = ~x36 & ~x109 ;
  assign n951 = ~x35 & x109 ;
  assign n952 = ~n950 & ~n951 ;
  assign n953 = ~x106 & ~n952 ;
  assign n954 = ~x98 & x106 ;
  assign n955 = ~x129 & ~n954 ;
  assign n956 = ~n953 & n955 ;
  assign n957 = ~x37 & ~x109 ;
  assign n958 = ~x36 & x109 ;
  assign n959 = ~n957 & ~n958 ;
  assign n960 = ~x106 & ~n959 ;
  assign n961 = ~x93 & x106 ;
  assign n962 = ~x129 & ~n961 ;
  assign n963 = ~n960 & n962 ;
  assign n964 = x82 & n273 ;
  assign n965 = n293 & ~n439 ;
  assign n966 = ~n441 & ~n572 ;
  assign n967 = ~x50 & n966 ;
  assign n968 = n965 & n967 ;
  assign n969 = x82 & ~n968 ;
  assign n970 = n267 & ~n969 ;
  assign n971 = ~n964 & ~n970 ;
  assign n972 = ~x38 & ~n971 ;
  assign n973 = ~x48 & n966 ;
  assign n974 = ~n287 & n293 ;
  assign n975 = ~x50 & n974 ;
  assign n976 = n973 & n975 ;
  assign n977 = ~n273 & n976 ;
  assign n978 = x82 & ~n977 ;
  assign n979 = x74 & ~n267 ;
  assign n980 = ~n978 & n979 ;
  assign n981 = ~x44 & x82 ;
  assign n982 = ~x40 & ~x42 ;
  assign n983 = x38 & n982 ;
  assign n984 = n981 & n983 ;
  assign n985 = ~x129 & ~n984 ;
  assign n986 = ~n980 & n985 ;
  assign n987 = ~n972 & n986 ;
  assign n988 = x109 & ~n677 ;
  assign n989 = x39 & ~n988 ;
  assign n990 = ~x51 & x109 ;
  assign n991 = ~n644 & n990 ;
  assign n992 = ~x106 & ~n991 ;
  assign n993 = ~n989 & n992 ;
  assign n994 = ~x129 & ~n993 ;
  assign n995 = ~x46 & n307 ;
  assign n996 = ~n292 & n310 ;
  assign n997 = n995 & n996 ;
  assign n998 = n966 & n997 ;
  assign n999 = ~n271 & n998 ;
  assign n1000 = x82 & ~n999 ;
  assign n1001 = x73 & ~n267 ;
  assign n1002 = ~n1000 & n1001 ;
  assign n1003 = x82 & n267 ;
  assign n1004 = ~n301 & n1003 ;
  assign n1005 = n1004 ^ n267 ;
  assign n1006 = x82 & n271 ;
  assign n1007 = ~x40 & ~n1006 ;
  assign n1008 = ~n1005 & n1007 ;
  assign n1009 = n1008 ^ x40 ;
  assign n1010 = ~x42 & n981 ;
  assign n1011 = x40 & n1010 ;
  assign n1012 = ~x129 & ~n1011 ;
  assign n1013 = ~n1009 & n1012 ;
  assign n1014 = n1013 ^ n1012 ;
  assign n1015 = n1002 & n1014 ;
  assign n1016 = n1015 ^ n1014 ;
  assign n1017 = ~n284 & n289 ;
  assign n1018 = n509 & n1017 ;
  assign n1019 = x82 & ~n1018 ;
  assign n1020 = x76 & ~n267 ;
  assign n1021 = ~n1019 & n1020 ;
  assign n1022 = x82 & ~n456 ;
  assign n1023 = x82 & ~n1017 ;
  assign n1024 = n267 & ~n1023 ;
  assign n1025 = ~n1022 & ~n1024 ;
  assign n1026 = ~x41 & ~n1025 ;
  assign n1027 = x41 & n1010 ;
  assign n1028 = n306 & n1027 ;
  assign n1029 = ~x129 & ~n1028 ;
  assign n1030 = ~n1026 & n1029 ;
  assign n1031 = ~n1021 & n1030 ;
  assign n1043 = x42 & n981 ;
  assign n1044 = ~x129 & ~n1043 ;
  assign n1047 = n1044 ^ x72 ;
  assign n1033 = ~x40 & x82 ;
  assign n1034 = n998 & n1033 ;
  assign n1035 = n1034 ^ x82 ;
  assign n1036 = x44 & x82 ;
  assign n1037 = n267 & ~n1036 ;
  assign n1038 = ~n1035 & n1037 ;
  assign n1039 = n1038 ^ n1036 ;
  assign n1040 = x42 & ~n1039 ;
  assign n1041 = n1040 ^ x42 ;
  assign n1042 = n1041 ^ n1039 ;
  assign n1057 = n1047 ^ n1042 ;
  assign n1051 = n982 & n998 ;
  assign n1048 = n1044 ^ n314 ;
  assign n1049 = n1047 & ~n1048 ;
  assign n1050 = n1049 ^ n314 ;
  assign n1052 = n1051 ^ n1050 ;
  assign n1058 = n1057 ^ n1052 ;
  assign n1059 = n1051 ^ x72 ;
  assign n1060 = n1059 ^ n1050 ;
  assign n1061 = ~n1058 & n1060 ;
  assign n1053 = n1050 ^ x72 ;
  assign n1045 = n1044 ^ n1042 ;
  assign n1054 = n1053 ^ n1045 ;
  assign n1055 = n1052 & n1054 ;
  assign n1062 = n1061 ^ n1055 ;
  assign n1063 = n1062 ^ n1050 ;
  assign n1064 = n1063 ^ n1057 ;
  assign n1065 = n1055 ^ n1051 ;
  assign n1066 = n1065 ^ n1042 ;
  assign n1067 = n1064 & n1066 ;
  assign n1068 = n1067 ^ n1061 ;
  assign n1056 = n1055 ^ n1049 ;
  assign n1069 = n1068 ^ n1056 ;
  assign n1032 = n314 ^ x72 ;
  assign n1046 = n1045 ^ n1032 ;
  assign n1070 = n1069 ^ n1046 ;
  assign n1071 = x82 & ~n437 ;
  assign n1072 = n445 & n447 ;
  assign n1073 = n446 & n1072 ;
  assign n1074 = x82 & ~n1073 ;
  assign n1075 = n267 & ~n1074 ;
  assign n1076 = ~n1071 & ~n1075 ;
  assign n1077 = ~x43 & ~n1076 ;
  assign n1078 = n310 & n966 ;
  assign n1079 = n437 & n1078 ;
  assign n1080 = x82 & ~n1079 ;
  assign n1081 = x77 & ~n267 ;
  assign n1082 = ~n1080 & n1081 ;
  assign n1083 = n981 & n982 ;
  assign n1084 = n294 & n1083 ;
  assign n1085 = x43 & n1084 ;
  assign n1086 = ~x129 & ~n1085 ;
  assign n1087 = ~n1082 & n1086 ;
  assign n1088 = ~n1077 & n1087 ;
  assign n1089 = x82 & ~n1051 ;
  assign n1090 = ~x67 & ~n267 ;
  assign n1091 = x44 & n267 ;
  assign n1092 = ~n1090 & ~n1091 ;
  assign n1093 = ~n1089 & n1092 ;
  assign n1094 = ~x129 & ~n1036 ;
  assign n1095 = ~n1093 & n1094 ;
  assign n1104 = n1072 ^ n311 ;
  assign n1105 = n1072 ^ x82 ;
  assign n1106 = ~x82 & ~n1105 ;
  assign n1107 = n1106 ^ x82 ;
  assign n1108 = n1107 ^ n311 ;
  assign n1109 = n1104 & ~n1108 ;
  assign n1110 = n1109 ^ n1106 ;
  assign n1111 = n1110 ^ n311 ;
  assign n1112 = x68 & ~n267 ;
  assign n1113 = ~n1111 & n1112 ;
  assign n1114 = n1113 ^ n1112 ;
  assign n1096 = x82 & ~n1072 ;
  assign n1097 = n267 & ~n1096 ;
  assign n1098 = x50 & n508 ;
  assign n1099 = n1098 ^ n508 ;
  assign n1100 = n965 & n1099 ;
  assign n1101 = x82 & ~n1100 ;
  assign n1102 = ~n1097 & ~n1101 ;
  assign n1103 = ~x45 & ~n1102 ;
  assign n1115 = n1114 ^ n1103 ;
  assign n1116 = x45 & x82 ;
  assign n1117 = n1100 & n1116 ;
  assign n1118 = ~x129 & ~n1117 ;
  assign n1119 = n1118 ^ n1114 ;
  assign n1120 = ~n1118 & ~n1119 ;
  assign n1121 = n1120 ^ n1114 ;
  assign n1122 = n1115 & n1121 ;
  assign n1123 = n1122 ^ n1120 ;
  assign n1124 = n1123 ^ n1103 ;
  assign n1125 = ~x75 & ~n267 ;
  assign n1126 = n307 & n310 ;
  assign n1127 = n966 & n1126 ;
  assign n1128 = x82 & ~n1127 ;
  assign n1129 = ~n1125 & ~n1128 ;
  assign n1130 = n509 & ~n1129 ;
  assign n1131 = ~x75 & n314 ;
  assign n1132 = x82 & n1099 ;
  assign n1133 = x46 & ~n314 ;
  assign n1134 = ~n1132 & n1133 ;
  assign n1135 = ~n1131 & ~n1134 ;
  assign n1136 = ~n1130 & n1135 ;
  assign n1137 = ~x129 & ~n1136 ;
  assign n1138 = n309 & n973 ;
  assign n1139 = x82 & ~n1138 ;
  assign n1140 = x64 & ~n267 ;
  assign n1141 = ~n1139 & n1140 ;
  assign n1142 = x82 & ~n309 ;
  assign n1143 = x82 & ~n973 ;
  assign n1144 = n267 & ~n1143 ;
  assign n1145 = ~n1142 & ~n1144 ;
  assign n1146 = ~x47 & ~n1145 ;
  assign n1147 = ~x43 & x47 ;
  assign n1148 = n1084 & n1147 ;
  assign n1149 = ~x129 & ~n1148 ;
  assign n1150 = ~n1146 & n1149 ;
  assign n1151 = ~n1141 & n1150 ;
  assign n1152 = x47 & n309 ;
  assign n1153 = n1152 ^ n309 ;
  assign n1154 = n966 & n1153 ;
  assign n1155 = x82 & ~n1154 ;
  assign n1156 = x62 & ~n267 ;
  assign n1157 = ~n1155 & n1156 ;
  assign n1158 = x82 & ~n966 ;
  assign n1159 = n267 & ~n1158 ;
  assign n1160 = n974 & n1099 ;
  assign n1161 = x82 & ~n1160 ;
  assign n1162 = ~n1159 & ~n1161 ;
  assign n1163 = ~x48 & ~n1162 ;
  assign n1164 = n438 & n1084 ;
  assign n1165 = ~x129 & ~n1164 ;
  assign n1166 = ~n1163 & n1165 ;
  assign n1167 = ~n1157 & n1166 ;
  assign n1168 = x46 & ~n292 ;
  assign n1169 = n1168 ^ n292 ;
  assign n1170 = ~x24 & ~x40 ;
  assign n1171 = ~n271 & n1170 ;
  assign n1172 = ~n1169 & n1171 ;
  assign n1173 = n577 & n1172 ;
  assign n1174 = x49 & ~n1173 ;
  assign n1175 = n513 & n572 ;
  assign n1176 = ~n1174 & ~n1175 ;
  assign n1177 = x82 & ~n1176 ;
  assign n1178 = x49 & n453 ;
  assign n1179 = x82 & ~n513 ;
  assign n1180 = ~x69 & ~n267 ;
  assign n1181 = ~n1179 & n1180 ;
  assign n1182 = ~n1178 & ~n1181 ;
  assign n1183 = ~n1177 & n1182 ;
  assign n1184 = ~x129 & ~n1183 ;
  assign n1185 = x82 & ~n508 ;
  assign n1186 = n293 & n1017 ;
  assign n1187 = x82 & ~n1186 ;
  assign n1188 = n267 & ~n1187 ;
  assign n1189 = ~n1185 & ~n1188 ;
  assign n1190 = ~x50 & ~n1189 ;
  assign n1191 = x82 & ~n976 ;
  assign n1192 = x66 & ~n267 ;
  assign n1193 = ~n1191 & n1192 ;
  assign n1194 = x50 & x82 ;
  assign n1195 = n508 & n1194 ;
  assign n1196 = ~x129 & ~n1195 ;
  assign n1197 = ~n1193 & n1196 ;
  assign n1198 = ~n1190 & n1197 ;
  assign n1199 = x51 & ~x109 ;
  assign n1200 = ~x106 & ~n990 ;
  assign n1201 = ~n1199 & n1200 ;
  assign n1202 = ~x129 & ~n1201 ;
  assign n1203 = x52 & ~n990 ;
  assign n1204 = ~x106 & ~n988 ;
  assign n1205 = ~n1203 & n1204 ;
  assign n1206 = ~x129 & ~n1205 ;
  assign n1207 = ~x116 & n839 ;
  assign n1208 = x58 & x116 ;
  assign n1209 = ~x58 & ~n683 ;
  assign n1210 = ~n850 & n1209 ;
  assign n1211 = ~n1208 & ~n1210 ;
  assign n1212 = ~x53 & x97 ;
  assign n1213 = ~n1211 & n1212 ;
  assign n1214 = ~n1207 & ~n1213 ;
  assign n1215 = n660 & n733 ;
  assign n1216 = ~n1214 & n1215 ;
  assign n1217 = ~n267 & n1072 ;
  assign n1218 = n601 & n1217 ;
  assign n1219 = ~x129 & ~n314 ;
  assign n1220 = ~n1218 & n1219 ;
  assign n1221 = ~x123 & ~x129 ;
  assign n1222 = x114 & ~x122 ;
  assign n1223 = n1221 & n1222 ;
  assign n1224 = ~x26 & x37 ;
  assign n1227 = n818 & n1224 ;
  assign n1225 = n659 & n1224 ;
  assign n1230 = n1227 ^ n1225 ;
  assign n1266 = n1230 ^ x27 ;
  assign n1238 = x116 ^ x58 ;
  assign n1236 = x116 ^ x26 ;
  assign n1237 = n1236 ^ x37 ;
  assign n1239 = n1238 ^ n1237 ;
  assign n1240 = n1239 ^ x37 ;
  assign n1242 = n1240 ^ n1238 ;
  assign n1234 = x116 ^ x94 ;
  assign n1235 = n1234 ^ x116 ;
  assign n1243 = n1242 ^ n1235 ;
  assign n1241 = n1240 ^ n1235 ;
  assign n1244 = n1243 ^ n1241 ;
  assign n1247 = ~n1235 & ~n1243 ;
  assign n1245 = n1240 ^ x37 ;
  assign n1246 = ~x116 & n1245 ;
  assign n1248 = n1247 ^ n1246 ;
  assign n1249 = ~n1244 & n1248 ;
  assign n1250 = n1249 ^ n1247 ;
  assign n1251 = n1250 ^ n1240 ;
  assign n1252 = n1251 ^ x116 ;
  assign n1253 = n1252 ^ x116 ;
  assign n1254 = x53 & ~n1253 ;
  assign n1255 = n1254 ^ x53 ;
  assign n1256 = n1255 ^ n1253 ;
  assign n1257 = ~x58 & n1224 ;
  assign n1258 = n1256 & n1257 ;
  assign n1259 = n1258 ^ n1256 ;
  assign n1260 = n1259 ^ n1257 ;
  assign n1231 = n1227 ^ x85 ;
  assign n1232 = n1230 & n1231 ;
  assign n1233 = n1232 ^ x85 ;
  assign n1261 = n1260 ^ n1233 ;
  assign n1267 = n1266 ^ n1261 ;
  assign n1268 = n1260 ^ n1225 ;
  assign n1269 = n1268 ^ n1233 ;
  assign n1270 = n1267 & n1269 ;
  assign n1262 = n1233 ^ n1225 ;
  assign n1228 = n1227 ^ x27 ;
  assign n1263 = n1262 ^ n1228 ;
  assign n1264 = ~n1261 & n1263 ;
  assign n1271 = n1270 ^ n1264 ;
  assign n1272 = n1271 ^ n1233 ;
  assign n1273 = n1272 ^ n1266 ;
  assign n1274 = n1264 ^ n1260 ;
  assign n1275 = n1274 ^ x27 ;
  assign n1276 = n1273 & ~n1275 ;
  assign n1277 = n1276 ^ n1270 ;
  assign n1265 = n1264 ^ n1232 ;
  assign n1278 = n1277 ^ n1265 ;
  assign n1226 = n1225 ^ x85 ;
  assign n1229 = n1228 ^ n1226 ;
  assign n1279 = n1278 ^ n1229 ;
  assign n1280 = n1279 ^ n1227 ;
  assign n1281 = n230 & ~n1280 ;
  assign n1282 = n1281 ^ n230 ;
  assign n1283 = ~x116 & n808 ;
  assign n1284 = x85 & ~n807 ;
  assign n1285 = x26 & x53 ;
  assign n1286 = ~x58 & ~n1285 ;
  assign n1287 = ~n1284 & n1286 ;
  assign n1288 = ~n1283 & ~n1287 ;
  assign n1289 = x57 & ~n1288 ;
  assign n1290 = x60 & n1208 ;
  assign n1291 = n808 & n1290 ;
  assign n1292 = ~n1289 & ~n1291 ;
  assign n1293 = ~x27 & ~n1292 ;
  assign n1294 = x57 & ~x58 ;
  assign n1295 = n808 & n1294 ;
  assign n1296 = ~n1293 & ~n1295 ;
  assign n1297 = n230 & ~n1296 ;
  assign n1298 = x58 & ~x116 ;
  assign n1299 = n751 & n1298 ;
  assign n1300 = ~x58 & n737 ;
  assign n1301 = n646 & n1300 ;
  assign n1302 = ~n1299 & ~n1301 ;
  assign n1303 = ~x53 & ~x85 ;
  assign n1304 = n230 & n1303 ;
  assign n1305 = ~n1302 & n1304 ;
  assign n1309 = n686 ^ x96 ;
  assign n1307 = x96 ^ x59 ;
  assign n1308 = n1307 ^ x96 ;
  assign n1310 = n1309 ^ n1308 ;
  assign n1311 = n1309 ^ x96 ;
  assign n1312 = n1310 & n1311 ;
  assign n1313 = n1312 ^ n1309 ;
  assign n1314 = x59 & ~x116 ;
  assign n1315 = n666 & n1314 ;
  assign n1316 = n659 & ~n1315 ;
  assign n1317 = n1313 & n1316 ;
  assign n1318 = n1317 ^ n1315 ;
  assign n1319 = n1318 ^ x85 ;
  assign n1320 = x85 & n659 ;
  assign n1321 = n1314 & n1320 ;
  assign n1322 = n1321 ^ x85 ;
  assign n1323 = n1321 & ~n1322 ;
  assign n1324 = n1323 ^ n1321 ;
  assign n1325 = n1324 ^ n1318 ;
  assign n1326 = ~n1319 & n1325 ;
  assign n1327 = n1326 ^ n1323 ;
  assign n1328 = n1327 ^ n1318 ;
  assign n1330 = n1328 ^ x27 ;
  assign n1306 = n737 ^ x27 ;
  assign n1329 = n1328 ^ n1306 ;
  assign n1331 = n1330 ^ n1329 ;
  assign n1333 = n818 & n1314 ;
  assign n1332 = n1328 & n1329 ;
  assign n1334 = n1333 ^ n1332 ;
  assign n1335 = n1331 & n1334 ;
  assign n1336 = n1335 ^ n1332 ;
  assign n1337 = n230 & ~n1336 ;
  assign n1338 = n1337 ^ n230 ;
  assign n1339 = ~x117 & ~x122 ;
  assign n1340 = x60 & ~n1339 ;
  assign n1341 = x123 & n1339 ;
  assign n1342 = ~n1340 & ~n1341 ;
  assign n1343 = ~x114 & ~x122 ;
  assign n1344 = x123 & ~x129 ;
  assign n1345 = n1343 & n1344 ;
  assign n1346 = x136 & ~x137 ;
  assign n1347 = x131 & x132 ;
  assign n1348 = x133 & n1347 ;
  assign n1349 = ~x138 & n1348 ;
  assign n1350 = n1346 & n1349 ;
  assign n1351 = x140 & n1350 ;
  assign n1352 = ~x62 & ~n1350 ;
  assign n1353 = ~x129 & ~n1352 ;
  assign n1354 = ~n1351 & n1353 ;
  assign n1355 = x142 & n1350 ;
  assign n1356 = ~x63 & ~n1350 ;
  assign n1357 = ~x129 & ~n1356 ;
  assign n1358 = ~n1355 & n1357 ;
  assign n1359 = x139 & n1350 ;
  assign n1360 = ~x64 & ~n1350 ;
  assign n1361 = ~x129 & ~n1360 ;
  assign n1362 = ~n1359 & n1361 ;
  assign n1363 = x146 & n1350 ;
  assign n1364 = ~x65 & ~n1350 ;
  assign n1365 = ~x129 & ~n1364 ;
  assign n1366 = ~n1363 & n1365 ;
  assign n1367 = ~x136 & ~x137 ;
  assign n1368 = n1349 & n1367 ;
  assign n1369 = x143 & n1368 ;
  assign n1370 = ~x66 & ~n1368 ;
  assign n1371 = ~x129 & ~n1370 ;
  assign n1372 = ~n1369 & n1371 ;
  assign n1373 = x139 & n1368 ;
  assign n1374 = ~x67 & ~n1368 ;
  assign n1375 = ~x129 & ~n1374 ;
  assign n1376 = ~n1373 & n1375 ;
  assign n1377 = x141 & n1350 ;
  assign n1378 = ~x68 & ~n1350 ;
  assign n1379 = ~x129 & ~n1378 ;
  assign n1380 = ~n1377 & n1379 ;
  assign n1381 = x143 & n1350 ;
  assign n1382 = ~x69 & ~n1350 ;
  assign n1383 = ~x129 & ~n1382 ;
  assign n1384 = ~n1381 & n1383 ;
  assign n1385 = x144 & n1350 ;
  assign n1386 = ~x70 & ~n1350 ;
  assign n1387 = ~x129 & ~n1386 ;
  assign n1388 = ~n1385 & n1387 ;
  assign n1389 = x145 & n1350 ;
  assign n1390 = ~x71 & ~n1350 ;
  assign n1391 = ~x129 & ~n1390 ;
  assign n1392 = ~n1389 & n1391 ;
  assign n1393 = x140 & n1368 ;
  assign n1394 = ~x72 & ~n1368 ;
  assign n1395 = ~x129 & ~n1394 ;
  assign n1396 = ~n1393 & n1395 ;
  assign n1397 = x141 & n1368 ;
  assign n1398 = ~x73 & ~n1368 ;
  assign n1399 = ~x129 & ~n1398 ;
  assign n1400 = ~n1397 & n1399 ;
  assign n1401 = x142 & n1368 ;
  assign n1402 = ~x74 & ~n1368 ;
  assign n1403 = ~x129 & ~n1402 ;
  assign n1404 = ~n1401 & n1403 ;
  assign n1405 = x144 & n1368 ;
  assign n1406 = ~x75 & ~n1368 ;
  assign n1407 = ~x129 & ~n1406 ;
  assign n1408 = ~n1405 & n1407 ;
  assign n1409 = x145 & n1368 ;
  assign n1410 = ~x76 & ~n1368 ;
  assign n1411 = ~x129 & ~n1410 ;
  assign n1412 = ~n1409 & n1411 ;
  assign n1413 = x146 & n1368 ;
  assign n1414 = ~x77 & ~n1368 ;
  assign n1415 = ~x129 & ~n1414 ;
  assign n1416 = ~n1413 & n1415 ;
  assign n1417 = ~x136 & x137 ;
  assign n1418 = n1349 & n1417 ;
  assign n1419 = ~x142 & n1418 ;
  assign n1420 = ~x78 & ~n1418 ;
  assign n1421 = ~x129 & ~n1420 ;
  assign n1422 = ~n1419 & n1421 ;
  assign n1423 = ~x143 & n1418 ;
  assign n1424 = ~x79 & ~n1418 ;
  assign n1425 = ~x129 & ~n1424 ;
  assign n1426 = ~n1423 & n1425 ;
  assign n1427 = ~x144 & n1418 ;
  assign n1428 = ~x80 & ~n1418 ;
  assign n1429 = ~x129 & ~n1428 ;
  assign n1430 = ~n1427 & n1429 ;
  assign n1431 = ~x145 & n1418 ;
  assign n1432 = ~x81 & ~n1418 ;
  assign n1433 = ~x129 & ~n1432 ;
  assign n1434 = ~n1431 & n1433 ;
  assign n1435 = ~x146 & n1418 ;
  assign n1436 = ~x82 & ~n1418 ;
  assign n1437 = ~x129 & ~n1436 ;
  assign n1438 = ~n1435 & n1437 ;
  assign n1439 = x136 & ~x138 ;
  assign n1440 = x31 & n1439 ;
  assign n1441 = x115 & x138 ;
  assign n1442 = ~x87 & ~x138 ;
  assign n1443 = ~x136 & ~n1442 ;
  assign n1444 = ~n1441 & n1443 ;
  assign n1445 = ~n1440 & ~n1444 ;
  assign n1446 = x137 & ~n1445 ;
  assign n1447 = x62 & ~x138 ;
  assign n1448 = ~x89 & x138 ;
  assign n1449 = x136 & ~n1448 ;
  assign n1450 = ~n1447 & n1449 ;
  assign n1451 = x72 & ~x138 ;
  assign n1452 = ~x119 & x138 ;
  assign n1453 = ~x136 & ~n1452 ;
  assign n1454 = ~n1451 & n1453 ;
  assign n1455 = ~n1450 & ~n1454 ;
  assign n1456 = ~x137 & ~n1455 ;
  assign n1457 = ~n1446 & ~n1456 ;
  assign n1458 = ~x141 & n1418 ;
  assign n1459 = ~x84 & ~n1418 ;
  assign n1460 = ~x129 & ~n1459 ;
  assign n1461 = ~n1458 & n1460 ;
  assign n1462 = x97 & ~n683 ;
  assign n1463 = n1462 ^ n683 ;
  assign n1464 = ~n726 & n1463 ;
  assign n1465 = x96 & n1464 ;
  assign n1466 = ~n622 & ~n1465 ;
  assign n1467 = n716 & n733 ;
  assign n1468 = ~n1466 & n1467 ;
  assign n1469 = ~x139 & n1418 ;
  assign n1470 = ~x86 & ~n1418 ;
  assign n1471 = ~x129 & ~n1470 ;
  assign n1472 = ~n1469 & n1471 ;
  assign n1473 = ~x140 & n1418 ;
  assign n1474 = ~x87 & ~n1418 ;
  assign n1475 = ~x129 & ~n1474 ;
  assign n1476 = ~n1473 & n1475 ;
  assign n1477 = x137 & n1439 ;
  assign n1478 = n1348 & n1477 ;
  assign n1479 = ~x139 & n1478 ;
  assign n1480 = ~x88 & ~n1478 ;
  assign n1481 = ~x129 & ~n1480 ;
  assign n1482 = ~n1479 & n1481 ;
  assign n1483 = ~x140 & n1478 ;
  assign n1484 = ~x89 & ~n1478 ;
  assign n1485 = ~x129 & ~n1484 ;
  assign n1486 = ~n1483 & n1485 ;
  assign n1487 = ~x142 & n1478 ;
  assign n1488 = ~x90 & ~n1478 ;
  assign n1489 = ~x129 & ~n1488 ;
  assign n1490 = ~n1487 & n1489 ;
  assign n1491 = ~x143 & n1478 ;
  assign n1492 = ~x91 & ~n1478 ;
  assign n1493 = ~x129 & ~n1492 ;
  assign n1494 = ~n1491 & n1493 ;
  assign n1495 = ~x144 & n1478 ;
  assign n1496 = ~x92 & ~n1478 ;
  assign n1497 = ~x129 & ~n1496 ;
  assign n1498 = ~n1495 & n1497 ;
  assign n1499 = ~x146 & n1478 ;
  assign n1500 = ~x93 & ~n1478 ;
  assign n1501 = ~x129 & ~n1500 ;
  assign n1502 = ~n1499 & n1501 ;
  assign n1503 = x82 & x138 ;
  assign n1504 = n1367 & n1503 ;
  assign n1505 = n1348 & n1504 ;
  assign n1506 = ~x142 & n1505 ;
  assign n1507 = ~x94 & ~n1505 ;
  assign n1508 = ~x129 & ~n1507 ;
  assign n1509 = ~n1506 & n1508 ;
  assign n1510 = ~x3 & ~x110 ;
  assign n1511 = ~n1348 & ~n1510 ;
  assign n1512 = ~n1505 & ~n1511 ;
  assign n1513 = x95 & n1512 ;
  assign n1514 = x143 & n1505 ;
  assign n1515 = ~n1513 & ~n1514 ;
  assign n1516 = ~x129 & ~n1515 ;
  assign n1517 = x96 & n1512 ;
  assign n1518 = x146 & n1505 ;
  assign n1519 = ~n1517 & ~n1518 ;
  assign n1520 = ~x129 & ~n1519 ;
  assign n1521 = x97 & n1512 ;
  assign n1522 = x145 & n1505 ;
  assign n1523 = ~n1521 & ~n1522 ;
  assign n1524 = ~x129 & ~n1523 ;
  assign n1525 = ~x145 & n1478 ;
  assign n1526 = ~x98 & ~n1478 ;
  assign n1527 = ~x129 & ~n1526 ;
  assign n1528 = ~n1525 & n1527 ;
  assign n1529 = ~x141 & n1478 ;
  assign n1530 = ~x99 & ~n1478 ;
  assign n1531 = ~x129 & ~n1530 ;
  assign n1532 = ~n1529 & n1531 ;
  assign n1533 = x100 & n1512 ;
  assign n1534 = x144 & n1505 ;
  assign n1535 = ~n1533 & ~n1534 ;
  assign n1536 = ~x129 & ~n1535 ;
  assign n1537 = x37 & n1439 ;
  assign n1538 = ~x96 & x138 ;
  assign n1539 = ~x82 & ~x138 ;
  assign n1540 = ~x136 & ~n1539 ;
  assign n1541 = ~n1538 & n1540 ;
  assign n1542 = ~n1537 & ~n1541 ;
  assign n1543 = x137 & ~n1542 ;
  assign n1544 = x65 & ~x138 ;
  assign n1545 = ~x93 & x138 ;
  assign n1546 = x136 & ~n1545 ;
  assign n1547 = ~n1544 & n1546 ;
  assign n1548 = x77 & ~x138 ;
  assign n1549 = ~x124 & x138 ;
  assign n1550 = ~x136 & ~n1549 ;
  assign n1551 = ~n1548 & n1550 ;
  assign n1552 = ~n1547 & ~n1551 ;
  assign n1553 = ~x137 & ~n1552 ;
  assign n1554 = ~n1543 & ~n1553 ;
  assign n1555 = x91 & n1346 ;
  assign n1556 = x95 & n1417 ;
  assign n1557 = ~n1555 & ~n1556 ;
  assign n1558 = x138 & ~n1557 ;
  assign n1559 = ~x34 & x136 ;
  assign n1560 = ~x79 & ~x136 ;
  assign n1561 = x137 & ~n1560 ;
  assign n1562 = ~n1559 & n1561 ;
  assign n1563 = x69 & x136 ;
  assign n1564 = x66 & ~x136 ;
  assign n1565 = ~x137 & ~n1564 ;
  assign n1566 = ~n1563 & n1565 ;
  assign n1567 = ~n1562 & ~n1566 ;
  assign n1568 = ~x138 & ~n1567 ;
  assign n1569 = ~n1558 & ~n1568 ;
  assign n1570 = x90 & n1346 ;
  assign n1571 = x94 & n1417 ;
  assign n1572 = ~n1570 & ~n1571 ;
  assign n1573 = x138 & ~n1572 ;
  assign n1574 = ~x33 & x136 ;
  assign n1575 = ~x78 & ~x136 ;
  assign n1576 = x137 & ~n1575 ;
  assign n1577 = ~n1574 & n1576 ;
  assign n1578 = x63 & x136 ;
  assign n1579 = x74 & ~x136 ;
  assign n1580 = ~x137 & ~n1579 ;
  assign n1581 = ~n1578 & n1580 ;
  assign n1582 = ~n1577 & ~n1581 ;
  assign n1583 = ~x138 & ~n1582 ;
  assign n1584 = ~n1573 & ~n1583 ;
  assign n1585 = x99 & n1346 ;
  assign n1586 = ~x112 & n1417 ;
  assign n1587 = ~n1585 & ~n1586 ;
  assign n1588 = x138 & ~n1587 ;
  assign n1589 = ~x32 & x136 ;
  assign n1590 = ~x84 & ~x136 ;
  assign n1591 = x137 & ~n1590 ;
  assign n1592 = ~n1589 & n1591 ;
  assign n1593 = x68 & x136 ;
  assign n1594 = x73 & ~x136 ;
  assign n1595 = ~x137 & ~n1594 ;
  assign n1596 = ~n1593 & n1595 ;
  assign n1597 = ~n1592 & ~n1596 ;
  assign n1598 = ~x138 & ~n1597 ;
  assign n1599 = ~n1588 & ~n1598 ;
  assign n1600 = x35 & n1439 ;
  assign n1601 = ~x100 & x138 ;
  assign n1602 = ~x80 & ~x138 ;
  assign n1603 = ~x136 & ~n1602 ;
  assign n1604 = ~n1601 & n1603 ;
  assign n1605 = ~n1600 & ~n1604 ;
  assign n1606 = x137 & ~n1605 ;
  assign n1607 = x70 & ~x138 ;
  assign n1608 = ~x92 & x138 ;
  assign n1609 = x136 & ~n1608 ;
  assign n1610 = ~n1607 & n1609 ;
  assign n1611 = x75 & ~x138 ;
  assign n1612 = ~x125 & x138 ;
  assign n1613 = ~x136 & ~n1612 ;
  assign n1614 = ~n1611 & n1613 ;
  assign n1615 = ~n1610 & ~n1614 ;
  assign n1616 = ~x137 & ~n1615 ;
  assign n1617 = ~n1606 & ~n1616 ;
  assign n1618 = ~x26 & n716 ;
  assign n1619 = n1464 & n1618 ;
  assign n1620 = ~n723 & ~n1619 ;
  assign n1621 = n230 & ~n1620 ;
  assign n1622 = x36 & n1439 ;
  assign n1623 = ~x97 & x138 ;
  assign n1624 = ~x81 & ~x138 ;
  assign n1625 = ~x136 & ~n1624 ;
  assign n1626 = ~n1623 & n1625 ;
  assign n1627 = ~n1622 & ~n1626 ;
  assign n1628 = x137 & ~n1627 ;
  assign n1629 = x71 & ~x138 ;
  assign n1630 = ~x98 & x138 ;
  assign n1631 = x136 & ~n1630 ;
  assign n1632 = ~n1629 & n1631 ;
  assign n1633 = x76 & ~x138 ;
  assign n1634 = ~x23 & x138 ;
  assign n1635 = ~x136 & ~n1634 ;
  assign n1636 = ~n1633 & n1635 ;
  assign n1637 = ~n1632 & ~n1636 ;
  assign n1638 = ~x137 & ~n1637 ;
  assign n1639 = ~n1628 & ~n1638 ;
  assign n1640 = x30 & n1439 ;
  assign n1641 = ~x111 & x138 ;
  assign n1642 = ~x86 & ~x138 ;
  assign n1643 = ~x136 & ~n1642 ;
  assign n1644 = ~n1641 & n1643 ;
  assign n1645 = ~n1640 & ~n1644 ;
  assign n1646 = x137 & ~n1645 ;
  assign n1647 = x64 & ~x138 ;
  assign n1648 = ~x88 & x138 ;
  assign n1649 = x136 & ~n1648 ;
  assign n1650 = ~n1647 & n1649 ;
  assign n1651 = x67 & ~x138 ;
  assign n1652 = ~x120 & x138 ;
  assign n1653 = ~x136 & ~n1652 ;
  assign n1654 = ~n1651 & n1653 ;
  assign n1655 = ~n1650 & ~n1654 ;
  assign n1656 = ~x137 & ~n1655 ;
  assign n1657 = ~n1646 & ~n1656 ;
  assign n1658 = ~n768 & ~n817 ;
  assign n1659 = x116 & n230 ;
  assign n1660 = ~n1658 & n1659 ;
  assign n1661 = ~x53 & x58 ;
  assign n1662 = ~x97 & n1661 ;
  assign n1663 = ~n839 & ~n1662 ;
  assign n1664 = n1659 & ~n1663 ;
  assign n1665 = ~x139 & n1504 ;
  assign n1666 = ~x129 & n1348 ;
  assign n1667 = ~x111 & ~n1504 ;
  assign n1668 = n1666 & ~n1667 ;
  assign n1669 = ~n1665 & n1668 ;
  assign n1670 = x112 & ~n1504 ;
  assign n1671 = ~x141 & n1504 ;
  assign n1672 = n1666 & ~n1671 ;
  assign n1673 = ~n1670 & n1672 ;
  assign n1674 = ~x11 & ~x22 ;
  assign n1675 = x54 & n1674 ;
  assign n1676 = ~x54 & x113 ;
  assign n1677 = n230 & ~n1676 ;
  assign n1678 = ~n1675 & n1677 ;
  assign n1679 = x115 & ~n1504 ;
  assign n1680 = ~x140 & n1504 ;
  assign n1681 = n1666 & ~n1680 ;
  assign n1682 = ~n1679 & n1681 ;
  assign n1683 = ~x4 & ~x9 ;
  assign n1684 = n245 & n1683 ;
  assign n1685 = x54 & n230 ;
  assign n1686 = ~n1684 & n1685 ;
  assign n1687 = x122 & ~x129 ;
  assign n1688 = ~x54 & x118 ;
  assign n1689 = x54 & ~x59 ;
  assign n1690 = n422 & n1689 ;
  assign n1691 = ~n1688 & ~n1690 ;
  assign n1692 = ~x129 & ~n1691 ;
  assign n1693 = ~x129 & n683 ;
  assign n1694 = ~x120 & n1510 ;
  assign n1695 = ~x111 & ~x129 ;
  assign n1696 = ~n1694 & n1695 ;
  assign n1697 = x81 & x120 ;
  assign n1698 = ~x129 & n1697 ;
  assign n1699 = ~x129 & ~x134 ;
  assign n1700 = ~x129 & ~x135 ;
  assign n1701 = x57 & ~x129 ;
  assign n1702 = ~x96 & x125 ;
  assign n1703 = ~x3 & ~n1702 ;
  assign n1704 = ~x129 & ~n1703 ;
  assign n1705 = ~x126 & x132 ;
  assign n1706 = x133 & n1705 ;
  assign y0 = x108 ;
  assign y1 = x83 ;
  assign y2 = x104 ;
  assign y3 = x103 ;
  assign y4 = x102 ;
  assign y5 = x105 ;
  assign y6 = x107 ;
  assign y7 = x101 ;
  assign y8 = x126 ;
  assign y9 = x121 ;
  assign y10 = x1 ;
  assign y11 = x0 ;
  assign y12 = ~1'b0 ;
  assign y13 = x130 ;
  assign y14 = x128 ;
  assign y15 = ~n232 ;
  assign y16 = ~n266 ;
  assign y17 = ~n327 ;
  assign y18 = n338 ;
  assign y19 = n349 ;
  assign y20 = n362 ;
  assign y21 = n370 ;
  assign y22 = n377 ;
  assign y23 = n388 ;
  assign y24 = n395 ;
  assign y25 = n405 ;
  assign y26 = n412 ;
  assign y27 = n419 ;
  assign y28 = n428 ;
  assign y29 = n436 ;
  assign y30 = n466 ;
  assign y31 = n473 ;
  assign y32 = n482 ;
  assign y33 = n489 ;
  assign y34 = n496 ;
  assign y35 = n551 ;
  assign y36 = n559 ;
  assign y37 = n568 ;
  assign y38 = n571 ;
  assign y39 = ~n621 ;
  assign y40 = ~n711 ;
  assign y41 = n718 ;
  assign y42 = n735 ;
  assign y43 = n815 ;
  assign y44 = n907 ;
  assign y45 = n914 ;
  assign y46 = n921 ;
  assign y47 = n928 ;
  assign y48 = n935 ;
  assign y49 = n942 ;
  assign y50 = n949 ;
  assign y51 = n956 ;
  assign y52 = n963 ;
  assign y53 = n987 ;
  assign y54 = n994 ;
  assign y55 = n1016 ;
  assign y56 = n1031 ;
  assign y57 = n1070 ;
  assign y58 = n1088 ;
  assign y59 = n1095 ;
  assign y60 = ~n1124 ;
  assign y61 = n1137 ;
  assign y62 = n1151 ;
  assign y63 = n1167 ;
  assign y64 = n1184 ;
  assign y65 = n1198 ;
  assign y66 = n1202 ;
  assign y67 = n1206 ;
  assign y68 = n1216 ;
  assign y69 = ~n1220 ;
  assign y70 = n1223 ;
  assign y71 = n1282 ;
  assign y72 = n1297 ;
  assign y73 = n1305 ;
  assign y74 = n1338 ;
  assign y75 = ~n1342 ;
  assign y76 = n1345 ;
  assign y77 = ~n1354 ;
  assign y78 = ~n1358 ;
  assign y79 = ~n1362 ;
  assign y80 = ~n1366 ;
  assign y81 = ~n1372 ;
  assign y82 = ~n1376 ;
  assign y83 = ~n1380 ;
  assign y84 = ~n1384 ;
  assign y85 = ~n1388 ;
  assign y86 = ~n1392 ;
  assign y87 = ~n1396 ;
  assign y88 = ~n1400 ;
  assign y89 = ~n1404 ;
  assign y90 = ~n1408 ;
  assign y91 = ~n1412 ;
  assign y92 = ~n1416 ;
  assign y93 = n1422 ;
  assign y94 = n1426 ;
  assign y95 = n1430 ;
  assign y96 = n1434 ;
  assign y97 = n1438 ;
  assign y98 = ~n1457 ;
  assign y99 = n1461 ;
  assign y100 = n1468 ;
  assign y101 = n1472 ;
  assign y102 = n1476 ;
  assign y103 = n1482 ;
  assign y104 = n1486 ;
  assign y105 = n1490 ;
  assign y106 = n1494 ;
  assign y107 = n1498 ;
  assign y108 = n1502 ;
  assign y109 = n1509 ;
  assign y110 = n1516 ;
  assign y111 = n1520 ;
  assign y112 = n1524 ;
  assign y113 = n1528 ;
  assign y114 = n1532 ;
  assign y115 = n1536 ;
  assign y116 = ~n1554 ;
  assign y117 = ~n1569 ;
  assign y118 = ~n1584 ;
  assign y119 = ~n1599 ;
  assign y120 = ~n1617 ;
  assign y121 = n1621 ;
  assign y122 = ~n1639 ;
  assign y123 = ~n1657 ;
  assign y124 = n1660 ;
  assign y125 = n1664 ;
  assign y126 = n1669 ;
  assign y127 = n1673 ;
  assign y128 = n1678 ;
  assign y129 = ~n1221 ;
  assign y130 = n1682 ;
  assign y131 = n1686 ;
  assign y132 = ~n1687 ;
  assign y133 = n1692 ;
  assign y134 = n1693 ;
  assign y135 = n1696 ;
  assign y136 = n1698 ;
  assign y137 = ~n1699 ;
  assign y138 = ~n1700 ;
  assign y139 = n1701 ;
  assign y140 = n1704 ;
  assign y141 = n1706 ;
endmodule
