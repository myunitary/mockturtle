module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , y0 , y1 , y2 , y3 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 ;
  output y0 , y1 , y2 , y3 ;
  wire n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 ;
  assign n278 = x61 ^ x5 ;
  assign n311 = x62 ^ x6 ;
  assign n279 = x67 ^ x11 ;
  assign n280 = x66 ^ x10 ;
  assign n281 = n279 & n280 ;
  assign n282 = x65 ^ x9 ;
  assign n283 = x64 ^ x8 ;
  assign n284 = ~n282 & ~n283 ;
  assign n285 = n281 & n284 ;
  assign n286 = x69 ^ x13 ;
  assign n287 = x68 ^ x12 ;
  assign n303 = n286 & ~n287 ;
  assign n304 = n303 ^ n287 ;
  assign n300 = ~n286 & ~n287 ;
  assign n290 = x70 ^ x14 ;
  assign n291 = x71 ^ x15 ;
  assign n301 = n290 & n291 ;
  assign n302 = n300 & n301 ;
  assign n305 = n304 ^ n302 ;
  assign n306 = n285 & n305 ;
  assign n113 = x63 ^ x7 ;
  assign n296 = n282 & ~n283 ;
  assign n297 = n296 ^ n283 ;
  assign n307 = n113 & ~n297 ;
  assign n308 = ~n306 & n307 ;
  assign n309 = n308 ^ n113 ;
  assign n298 = ~n113 & n297 ;
  assign n288 = n286 & n287 ;
  assign n289 = n285 & n288 ;
  assign n292 = ~n290 & n291 ;
  assign n293 = n292 ^ n290 ;
  assign n294 = ~n113 & n293 ;
  assign n295 = n289 & n294 ;
  assign n299 = n298 ^ n295 ;
  assign n310 = n309 ^ n299 ;
  assign n312 = n311 ^ n310 ;
  assign n327 = n278 & n312 ;
  assign n330 = n298 & n309 ;
  assign n329 = n295 & n309 ;
  assign n331 = n330 ^ n329 ;
  assign n328 = n310 & n311 ;
  assign n332 = n331 ^ n328 ;
  assign n347 = n327 & n332 ;
  assign n348 = n328 & n331 ;
  assign n363 = n347 & n348 ;
  assign n277 = x60 ^ x4 ;
  assign n313 = n312 ^ n278 ;
  assign n326 = n277 & n313 ;
  assign n333 = n332 ^ n327 ;
  assign n346 = n326 & n333 ;
  assign n349 = n348 ^ n347 ;
  assign n362 = n346 & n349 ;
  assign n364 = n363 ^ n362 ;
  assign n276 = x59 ^ x3 ;
  assign n314 = n313 ^ n277 ;
  assign n325 = n276 & n314 ;
  assign n334 = n333 ^ n326 ;
  assign n345 = n325 & n334 ;
  assign n350 = n349 ^ n346 ;
  assign n361 = n345 & n350 ;
  assign n365 = n364 ^ n361 ;
  assign n248 = x73 ^ x17 ;
  assign n249 = x72 ^ x16 ;
  assign n271 = n248 & ~n249 ;
  assign n272 = n271 ^ n249 ;
  assign n250 = ~n248 & ~n249 ;
  assign n251 = x75 ^ x19 ;
  assign n252 = x74 ^ x18 ;
  assign n269 = n251 & n252 ;
  assign n270 = n250 & n269 ;
  assign n273 = n272 ^ n270 ;
  assign n253 = ~n251 & n252 ;
  assign n254 = n250 & n253 ;
  assign n255 = x77 ^ x21 ;
  assign n256 = x76 ^ x20 ;
  assign n266 = n255 & n256 ;
  assign n257 = ~n255 & n256 ;
  assign n258 = x79 ^ x23 ;
  assign n259 = x78 ^ x22 ;
  assign n263 = n258 & ~n259 ;
  assign n264 = n263 ^ n259 ;
  assign n265 = n257 & n264 ;
  assign n267 = n266 ^ n265 ;
  assign n268 = n254 & n267 ;
  assign n274 = n273 ^ n268 ;
  assign n260 = ~n258 & ~n259 ;
  assign n261 = n257 & n260 ;
  assign n262 = n254 & n261 ;
  assign n275 = n274 ^ n262 ;
  assign n315 = n314 ^ n276 ;
  assign n324 = ~n275 & n315 ;
  assign n335 = n334 ^ n325 ;
  assign n344 = n324 & n335 ;
  assign n351 = n350 ^ n345 ;
  assign n360 = n344 & n351 ;
  assign n366 = n365 ^ n360 ;
  assign n168 = x80 ^ x24 ;
  assign n187 = x88 ^ x32 ;
  assign n169 = x94 ^ x38 ;
  assign n170 = x93 ^ x37 ;
  assign n171 = ~n169 & n170 ;
  assign n172 = n171 ^ n169 ;
  assign n173 = x92 ^ x36 ;
  assign n178 = n172 & ~n173 ;
  assign n179 = n178 ^ n172 ;
  assign n174 = x91 ^ x35 ;
  assign n175 = n173 & n174 ;
  assign n176 = n172 & n175 ;
  assign n177 = n176 ^ n174 ;
  assign n180 = n179 ^ n177 ;
  assign n181 = x90 ^ x34 ;
  assign n184 = ~n180 & n181 ;
  assign n185 = n184 ^ n180 ;
  assign n167 = x89 ^ x33 ;
  assign n182 = n167 & ~n181 ;
  assign n183 = ~n180 & n182 ;
  assign n186 = n185 ^ n183 ;
  assign n188 = n187 ^ n186 ;
  assign n244 = ~n168 & ~n188 ;
  assign n189 = n188 ^ n168 ;
  assign n193 = x81 ^ x25 ;
  assign n194 = n189 & ~n193 ;
  assign n191 = ~n185 & n189 ;
  assign n190 = n167 & n189 ;
  assign n192 = n191 ^ n190 ;
  assign n195 = n194 ^ n192 ;
  assign n223 = x82 ^ x26 ;
  assign n237 = n181 ^ n180 ;
  assign n241 = ~n223 & ~n237 ;
  assign n238 = n237 ^ n223 ;
  assign n218 = x83 ^ x27 ;
  assign n219 = n179 ^ n174 ;
  assign n239 = ~n218 & ~n219 ;
  assign n240 = n238 & n239 ;
  assign n242 = n241 ^ n240 ;
  assign n243 = n195 & n242 ;
  assign n245 = n244 ^ n243 ;
  assign n231 = n185 ^ n167 ;
  assign n234 = ~n188 & ~n193 ;
  assign n235 = ~n231 & n234 ;
  assign n232 = ~n168 & ~n193 ;
  assign n233 = ~n231 & n232 ;
  assign n236 = n235 ^ n233 ;
  assign n246 = n245 ^ n236 ;
  assign n196 = x84 ^ x28 ;
  assign n197 = n173 ^ n172 ;
  assign n215 = ~n196 & n197 ;
  assign n198 = n197 ^ n196 ;
  assign n202 = x85 ^ x29 ;
  assign n203 = n170 ^ n169 ;
  assign n213 = ~n202 & ~n203 ;
  assign n214 = ~n198 & n213 ;
  assign n216 = n215 ^ n214 ;
  assign n204 = n203 ^ n202 ;
  assign n205 = x86 ^ x30 ;
  assign n209 = ~n169 & ~n205 ;
  assign n210 = n204 & n209 ;
  assign n199 = x87 ^ x31 ;
  assign n200 = x95 ^ x39 ;
  assign n201 = ~n199 & n200 ;
  assign n206 = n205 ^ n169 ;
  assign n207 = n204 & n206 ;
  assign n208 = n201 & n207 ;
  assign n211 = n210 ^ n208 ;
  assign n212 = ~n198 & n211 ;
  assign n217 = n216 ^ n212 ;
  assign n220 = n219 ^ n218 ;
  assign n227 = ~n180 & n220 ;
  assign n228 = n217 & n227 ;
  assign n224 = n220 & ~n223 ;
  assign n225 = n217 & n224 ;
  assign n221 = n181 & n220 ;
  assign n222 = n217 & n221 ;
  assign n226 = n225 ^ n222 ;
  assign n229 = n228 ^ n226 ;
  assign n230 = n195 & n229 ;
  assign n247 = n246 ^ n230 ;
  assign n316 = n315 ^ n275 ;
  assign n323 = n247 & ~n316 ;
  assign n336 = n335 ^ n324 ;
  assign n343 = n323 & n336 ;
  assign n352 = n351 ^ n344 ;
  assign n359 = n343 & n352 ;
  assign n367 = n366 ^ n359 ;
  assign n143 = x97 ^ x41 ;
  assign n144 = x96 ^ x40 ;
  assign n162 = n143 & ~n144 ;
  assign n163 = n162 ^ n144 ;
  assign n145 = ~n143 & ~n144 ;
  assign n146 = x98 ^ x42 ;
  assign n161 = n145 & n146 ;
  assign n164 = n163 ^ n161 ;
  assign n147 = x99 ^ x43 ;
  assign n148 = ~n146 & n147 ;
  assign n149 = n145 & n148 ;
  assign n150 = x101 ^ x45 ;
  assign n151 = x100 ^ x44 ;
  assign n152 = n150 & n151 ;
  assign n153 = x103 ^ x47 ;
  assign n154 = x102 ^ x46 ;
  assign n158 = n153 & n154 ;
  assign n159 = n152 & n158 ;
  assign n160 = n149 & n159 ;
  assign n165 = n164 ^ n160 ;
  assign n155 = ~n153 & n154 ;
  assign n156 = n152 & n155 ;
  assign n157 = n149 & n156 ;
  assign n166 = n165 ^ n157 ;
  assign n317 = n316 ^ n247 ;
  assign n322 = ~n166 & ~n317 ;
  assign n337 = n336 ^ n323 ;
  assign n342 = n322 & n337 ;
  assign n353 = n352 ^ n343 ;
  assign n358 = n342 & n353 ;
  assign n368 = n367 ^ n358 ;
  assign n114 = x105 ^ x49 ;
  assign n115 = x104 ^ x48 ;
  assign n116 = ~n114 & ~n115 ;
  assign n117 = x107 ^ x51 ;
  assign n118 = x106 ^ x50 ;
  assign n119 = ~n117 & ~n118 ;
  assign n120 = n116 & n119 ;
  assign n124 = x109 ^ x53 ;
  assign n125 = x108 ^ x52 ;
  assign n128 = n124 & ~n125 ;
  assign n129 = n128 ^ n125 ;
  assign n140 = n120 & n129 ;
  assign n135 = n114 & ~n115 ;
  assign n136 = n135 ^ n115 ;
  assign n132 = n117 & ~n118 ;
  assign n133 = n132 ^ n118 ;
  assign n134 = n116 & n133 ;
  assign n137 = n136 ^ n134 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n113 & n141 ;
  assign n318 = n317 ^ n166 ;
  assign n321 = n142 & n318 ;
  assign n338 = n337 ^ n322 ;
  assign n341 = n321 & n338 ;
  assign n354 = n353 ^ n342 ;
  assign n357 = n341 & n354 ;
  assign n369 = n368 ^ n357 ;
  assign n121 = x111 ^ x55 ;
  assign n122 = x110 ^ x54 ;
  assign n123 = n121 & n122 ;
  assign n126 = ~n124 & ~n125 ;
  assign n127 = n123 & n126 ;
  assign n130 = n129 ^ n127 ;
  assign n131 = n120 & n130 ;
  assign n138 = n137 ^ n131 ;
  assign n139 = ~n113 & n138 ;
  assign n319 = n318 ^ n142 ;
  assign n320 = n139 & n319 ;
  assign n339 = n338 ^ n321 ;
  assign n340 = n320 & n339 ;
  assign n355 = n354 ^ n341 ;
  assign n356 = n340 & n355 ;
  assign n370 = n369 ^ n356 ;
  assign n371 = n355 ^ n340 ;
  assign n372 = n339 ^ n320 ;
  assign n373 = n319 ^ n139 ;
  assign y0 = n370 ;
  assign y1 = n371 ;
  assign y2 = n372 ;
  assign y3 = n373 ;
endmodule
