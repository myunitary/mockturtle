module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 ;
  assign n33 = x29 & x30 ;
  assign n34 = x27 & x28 ;
  assign n35 = n33 & n34 ;
  assign n36 = x26 & x27 ;
  assign n37 = n35 & n36 ;
  assign n38 = x22 & x23 ;
  assign n39 = x23 & x24 ;
  assign n40 = n38 & n39 ;
  assign n41 = x25 & x26 ;
  assign n42 = x24 & x25 ;
  assign n43 = n41 & n42 ;
  assign n44 = n40 & n43 ;
  assign n45 = ~n37 & ~n44 ;
  assign n46 = n34 & n36 ;
  assign n47 = n43 & n46 ;
  assign n48 = ~n45 & n47 ;
  assign n49 = x28 & x29 ;
  assign n50 = x30 & x31 ;
  assign n51 = n49 & n50 ;
  assign n52 = n34 & n51 ;
  assign n53 = n36 & n41 ;
  assign n54 = n39 & n42 ;
  assign n55 = n53 & n54 ;
  assign n56 = n52 & n55 ;
  assign n57 = n56 ^ n52 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n34 & n49 ;
  assign n60 = n53 & n59 ;
  assign n61 = ~n58 & n60 ;
  assign n62 = n61 ^ n60 ;
  assign n63 = n48 & n62 ;
  assign n64 = x10 & x11 ;
  assign n65 = x17 & x18 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = x12 & x13 ;
  assign n68 = x13 & x14 ;
  assign n69 = n67 & n68 ;
  assign n70 = x14 & x15 ;
  assign n71 = x15 & x16 ;
  assign n72 = n70 & n71 ;
  assign n73 = n69 & n72 ;
  assign n74 = n66 & n73 ;
  assign n75 = n74 ^ n73 ;
  assign n76 = x16 & x17 ;
  assign n77 = n71 & n76 ;
  assign n78 = x19 & x20 ;
  assign n79 = n65 & n78 ;
  assign n80 = n77 & n79 ;
  assign n81 = n75 & n80 ;
  assign n82 = n81 ^ n75 ;
  assign n83 = n82 ^ n80 ;
  assign n84 = x18 & x19 ;
  assign n85 = x11 & x12 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = n68 & n70 ;
  assign n88 = n77 & n87 ;
  assign n89 = n86 & n88 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = ~n83 & n90 ;
  assign n92 = n91 ^ n90 ;
  assign n93 = x21 & x22 ;
  assign n94 = ~n70 & ~n93 ;
  assign n95 = n78 & n84 ;
  assign n96 = n65 & n76 ;
  assign n97 = n95 & n96 ;
  assign n98 = n94 & n97 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = n65 & n84 ;
  assign n101 = n77 & n100 ;
  assign n102 = x20 & x21 ;
  assign n103 = n84 & n102 ;
  assign n104 = n96 & n103 ;
  assign n105 = n101 & n104 ;
  assign n106 = n99 & n105 ;
  assign n107 = n92 & n106 ;
  assign n108 = n107 ^ n92 ;
  assign n109 = n108 ^ n106 ;
  assign n110 = n63 & ~n109 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = n78 & n93 ;
  assign n113 = n95 & n112 ;
  assign n114 = n38 & n102 ;
  assign n115 = n113 & n114 ;
  assign n116 = n65 & n103 ;
  assign n117 = n115 & n116 ;
  assign n118 = ~n39 & ~n76 ;
  assign n119 = n117 & ~n118 ;
  assign n120 = ~n41 & ~n84 ;
  assign n121 = n39 & n93 ;
  assign n122 = n102 & n121 ;
  assign n123 = ~n120 & n122 ;
  assign n124 = n34 & n41 ;
  assign n125 = n54 & n124 ;
  assign n126 = ~n123 & ~n125 ;
  assign n127 = ~n36 & ~n78 ;
  assign n128 = n38 & n93 ;
  assign n129 = n54 & n128 ;
  assign n130 = ~n127 & n129 ;
  assign n131 = ~n126 & n130 ;
  assign n132 = ~n119 & ~n131 ;
  assign n133 = ~n111 & n132 ;
  assign n135 = n67 & n85 ;
  assign n139 = x9 & x10 ;
  assign n148 = n64 & n139 ;
  assign n159 = n135 & n148 ;
  assign n142 = x7 & x8 ;
  assign n160 = ~n70 & ~n142 ;
  assign n161 = n159 & n160 ;
  assign n162 = n161 ^ n159 ;
  assign n134 = n68 & n71 ;
  assign n136 = n134 & n135 ;
  assign n163 = n162 ^ n136 ;
  assign n164 = ~n162 & n163 ;
  assign n165 = n164 ^ n162 ;
  assign n137 = x8 & x9 ;
  assign n138 = x7 & n137 ;
  assign n140 = n85 & n139 ;
  assign n141 = n138 & n140 ;
  assign n143 = n139 & n142 ;
  assign n144 = x6 & x7 ;
  assign n145 = n142 & n144 ;
  assign n146 = n143 & n145 ;
  assign n147 = n141 & n146 ;
  assign n149 = n68 & n85 ;
  assign n150 = n148 & n149 ;
  assign n151 = n137 & n139 ;
  assign n152 = n64 & n85 ;
  assign n153 = n151 & n152 ;
  assign n154 = n150 & n153 ;
  assign n155 = n147 & n154 ;
  assign n156 = n155 ^ n147 ;
  assign n157 = n156 ^ n154 ;
  assign n166 = n165 ^ n157 ;
  assign n158 = n157 ^ n136 ;
  assign n167 = n166 ^ n158 ;
  assign n168 = n167 ^ n164 ;
  assign n169 = n168 ^ n157 ;
  assign n170 = x4 & x5 ;
  assign n171 = x3 & x4 ;
  assign n172 = n170 & n171 ;
  assign n173 = x5 & x6 ;
  assign n174 = n142 & n173 ;
  assign n175 = n172 & n174 ;
  assign n176 = n170 & n173 ;
  assign n177 = x2 & x3 ;
  assign n178 = n171 & n177 ;
  assign n179 = n176 & n178 ;
  assign n180 = n175 & n179 ;
  assign n181 = n137 & n144 ;
  assign n182 = n173 & n181 ;
  assign n183 = n143 & n182 ;
  assign n184 = n170 & n177 ;
  assign n185 = x1 & x2 ;
  assign n186 = n171 & n185 ;
  assign n187 = x0 & x1 ;
  assign n188 = n186 & n187 ;
  assign n189 = n184 & n188 ;
  assign n190 = n183 & n189 ;
  assign n191 = n190 ^ n183 ;
  assign n192 = n191 ^ n189 ;
  assign n193 = n180 & ~n192 ;
  assign n194 = n193 ^ n192 ;
  assign n195 = n144 & n173 ;
  assign n196 = n172 & n195 ;
  assign n197 = n176 & n181 ;
  assign n198 = n196 & n197 ;
  assign n199 = n177 & n185 ;
  assign n200 = n172 & n199 ;
  assign n201 = n144 & n170 ;
  assign n202 = n178 & n201 ;
  assign n203 = n200 & n202 ;
  assign n204 = n198 & n203 ;
  assign n205 = n204 ^ n198 ;
  assign n206 = n205 ^ n203 ;
  assign n207 = ~n194 & ~n206 ;
  assign n208 = n207 ^ n194 ;
  assign n209 = n208 ^ n206 ;
  assign n210 = n145 & n176 ;
  assign n211 = n183 & n210 ;
  assign n212 = n147 & n211 ;
  assign n213 = n212 ^ n147 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = n64 & n137 ;
  assign n216 = n146 & n215 ;
  assign n217 = n182 & n216 ;
  assign n218 = ~n214 & n217 ;
  assign n219 = n218 ^ n217 ;
  assign n220 = ~n209 & n219 ;
  assign n221 = n220 ^ n209 ;
  assign n222 = n221 ^ n219 ;
  assign n223 = n169 & n222 ;
  assign n224 = n223 ^ n222 ;
  assign n225 = n133 & n224 ;
  assign n520 = ~n71 & ~n177 ;
  assign n521 = ~n33 & ~n49 ;
  assign n522 = n520 & n521 ;
  assign n523 = ~n64 & ~n85 ;
  assign n524 = ~n67 & ~n68 ;
  assign n525 = n523 & n524 ;
  assign n526 = n522 & n525 ;
  assign n527 = ~n50 & ~n93 ;
  assign n528 = ~n42 & n527 ;
  assign n529 = ~n34 & ~n36 ;
  assign n530 = n120 & n529 ;
  assign n531 = n528 & n530 ;
  assign n532 = n526 & n531 ;
  assign n533 = ~n144 & ~n173 ;
  assign n534 = n118 & n533 ;
  assign n461 = ~n38 & ~n102 ;
  assign n535 = ~n65 & ~n78 ;
  assign n536 = n461 & n535 ;
  assign n537 = n534 & n536 ;
  assign n538 = ~n137 & ~n139 ;
  assign n539 = ~n185 & ~n187 ;
  assign n540 = n538 & n539 ;
  assign n541 = ~n170 & ~n171 ;
  assign n542 = n160 & n541 ;
  assign n543 = n540 & n542 ;
  assign n544 = n537 & n543 ;
  assign n545 = n532 & n544 ;
  assign n491 = ~x18 & ~x19 ;
  assign n492 = ~x21 & ~x22 ;
  assign n493 = n491 & n492 ;
  assign n494 = ~x14 & ~x15 ;
  assign n495 = ~x16 & ~x17 ;
  assign n496 = n494 & n495 ;
  assign n497 = n493 & n496 ;
  assign n498 = ~x28 & ~x29 ;
  assign n499 = ~x30 & ~x31 ;
  assign n500 = n498 & n499 ;
  assign n501 = ~x23 & ~x24 ;
  assign n502 = ~x25 & ~x27 ;
  assign n503 = n501 & n502 ;
  assign n504 = n500 & n503 ;
  assign n505 = n497 & n504 ;
  assign n506 = ~x1 & ~x2 ;
  assign n507 = ~x4 & ~x5 ;
  assign n508 = n506 & n507 ;
  assign n271 = ~x20 & ~x26 ;
  assign n446 = ~x0 & ~x3 ;
  assign n509 = n271 & n446 ;
  assign n510 = n508 & n509 ;
  assign n511 = ~x10 & ~x11 ;
  assign n512 = ~x12 & ~x13 ;
  assign n513 = n511 & n512 ;
  assign n514 = ~x6 & ~x7 ;
  assign n515 = ~x8 & ~x9 ;
  assign n516 = n514 & n515 ;
  assign n517 = n513 & n516 ;
  assign n518 = n510 & n517 ;
  assign n519 = n505 & n518 ;
  assign n546 = n545 ^ n519 ;
  assign n430 = n44 ^ n40 ;
  assign n431 = n430 ^ n43 ;
  assign n432 = n33 & n50 ;
  assign n433 = n46 & n432 ;
  assign n434 = n433 ^ n46 ;
  assign n435 = n434 ^ n432 ;
  assign n436 = ~n431 & ~n435 ;
  assign n437 = n87 & n151 ;
  assign n438 = n437 ^ n87 ;
  assign n439 = n438 ^ n151 ;
  assign n440 = n33 & n49 ;
  assign n441 = n72 & n440 ;
  assign n442 = n441 ^ n72 ;
  assign n443 = n442 ^ n440 ;
  assign n444 = ~n439 & ~n443 ;
  assign n445 = n436 & n444 ;
  assign n447 = n185 & ~n446 ;
  assign n448 = ~x15 & x16 ;
  assign n449 = x17 & ~x18 ;
  assign n450 = n448 & n449 ;
  assign n451 = n450 ^ n76 ;
  assign n452 = ~n447 & ~n451 ;
  assign n453 = n55 ^ n53 ;
  assign n454 = n453 ^ n54 ;
  assign n281 = x19 & n102 ;
  assign n455 = n59 & n281 ;
  assign n456 = n455 ^ n59 ;
  assign n457 = n456 ^ n281 ;
  assign n458 = ~n454 & ~n457 ;
  assign n459 = n452 & n458 ;
  assign n460 = n445 & n459 ;
  assign n462 = n93 & ~n461 ;
  assign n463 = ~x17 & x18 ;
  assign n464 = x19 & ~x20 ;
  assign n465 = n463 & n464 ;
  assign n466 = n465 ^ n84 ;
  assign n467 = n196 ^ n195 ;
  assign n468 = n467 ^ n172 ;
  assign n469 = n466 & ~n468 ;
  assign n470 = n469 ^ n468 ;
  assign n471 = n462 & ~n470 ;
  assign n472 = n471 ^ n470 ;
  assign n473 = ~x9 & x10 ;
  assign n474 = x11 & ~x12 ;
  assign n475 = n473 & n474 ;
  assign n476 = n475 ^ n64 ;
  assign n477 = ~x11 & x12 ;
  assign n478 = x13 & ~x14 ;
  assign n479 = n477 & n478 ;
  assign n480 = n479 ^ n67 ;
  assign n481 = ~n476 & ~n480 ;
  assign n482 = n210 ^ n145 ;
  assign n483 = n482 ^ n176 ;
  assign n484 = n138 & n178 ;
  assign n485 = n484 ^ n138 ;
  assign n486 = n485 ^ n178 ;
  assign n487 = ~n483 & ~n486 ;
  assign n488 = n481 & n487 ;
  assign n489 = ~n472 & n488 ;
  assign n490 = n460 & n489 ;
  assign n547 = n546 ^ n490 ;
  assign n370 = n38 & n42 ;
  assign n371 = n177 & n187 ;
  assign n372 = n370 & n371 ;
  assign n373 = n372 ^ n370 ;
  assign n374 = n373 ^ n371 ;
  assign n375 = n65 & n71 ;
  assign n376 = n64 & n67 ;
  assign n377 = n375 & n376 ;
  assign n378 = n377 ^ n376 ;
  assign n379 = n378 ^ n375 ;
  assign n380 = ~n374 & ~n379 ;
  assign n233 = n171 & n173 ;
  assign n381 = n149 & n233 ;
  assign n382 = n381 ^ n233 ;
  assign n383 = n382 ^ n149 ;
  assign n384 = n124 & n174 ;
  assign n385 = n384 ^ n174 ;
  assign n386 = n385 ^ n124 ;
  assign n387 = ~n383 & ~n386 ;
  assign n388 = n380 & n387 ;
  assign n389 = n76 & n84 ;
  assign n390 = n201 & n389 ;
  assign n391 = n390 ^ n201 ;
  assign n392 = n391 ^ n389 ;
  assign n393 = n79 & ~n392 ;
  assign n394 = n393 ^ n392 ;
  assign n395 = n134 & n140 ;
  assign n396 = n395 ^ n134 ;
  assign n397 = n396 ^ n140 ;
  assign n257 = n67 & n70 ;
  assign n398 = n39 & n41 ;
  assign n399 = n257 & n398 ;
  assign n400 = n399 ^ n398 ;
  assign n401 = n400 ^ n257 ;
  assign n402 = ~n397 & ~n401 ;
  assign n403 = ~n394 & n402 ;
  assign n404 = n388 & n403 ;
  assign n255 = n36 & n42 ;
  assign n292 = n51 & n255 ;
  assign n293 = n292 ^ n51 ;
  assign n294 = n293 ^ n255 ;
  assign n405 = n143 & n181 ;
  assign n406 = n405 ^ n143 ;
  assign n407 = n406 ^ n181 ;
  assign n408 = n184 & n186 ;
  assign n409 = n408 ^ n186 ;
  assign n410 = n409 ^ n184 ;
  assign n411 = ~n407 & ~n410 ;
  assign n412 = ~n294 & n411 ;
  assign n413 = n103 & n121 ;
  assign n414 = n413 ^ n103 ;
  assign n415 = n414 ^ n121 ;
  assign n291 = n36 & n49 ;
  assign n297 = n70 & n76 ;
  assign n416 = n291 & n297 ;
  assign n417 = n416 ^ n291 ;
  assign n418 = n417 ^ n297 ;
  assign n419 = ~n415 & ~n418 ;
  assign n420 = n35 & n215 ;
  assign n421 = n420 ^ n35 ;
  assign n422 = n421 ^ n215 ;
  assign n423 = n112 & n114 ;
  assign n424 = n423 ^ n112 ;
  assign n425 = n424 ^ n114 ;
  assign n426 = ~n422 & ~n425 ;
  assign n427 = n419 & n426 ;
  assign n428 = n412 & n427 ;
  assign n429 = n404 & n428 ;
  assign n548 = n547 ^ n429 ;
  assign n322 = n179 & n196 ;
  assign n323 = n322 ^ n196 ;
  assign n324 = n323 ^ n179 ;
  assign n325 = n182 & ~n324 ;
  assign n326 = n325 ^ n324 ;
  assign n327 = ~n146 & ~n188 ;
  assign n328 = ~n326 & n327 ;
  assign n329 = n87 & n135 ;
  assign n330 = n153 & n329 ;
  assign n331 = n330 ^ n153 ;
  assign n332 = n331 ^ n329 ;
  assign n333 = n47 & n60 ;
  assign n334 = n333 ^ n47 ;
  assign n335 = n334 ^ n60 ;
  assign n336 = ~n332 & ~n335 ;
  assign n337 = n138 & n148 ;
  assign n338 = n200 & n337 ;
  assign n339 = n338 ^ n337 ;
  assign n340 = n339 ^ n200 ;
  assign n341 = n159 & n210 ;
  assign n342 = n341 ^ n159 ;
  assign n343 = n342 ^ n210 ;
  assign n344 = ~n340 & ~n343 ;
  assign n345 = n336 & n344 ;
  assign n346 = n328 & n345 ;
  assign n347 = n69 & n152 ;
  assign n348 = n129 & n347 ;
  assign n349 = n348 ^ n129 ;
  assign n350 = n349 ^ n347 ;
  assign n274 = n72 & n96 ;
  assign n351 = n128 & n281 ;
  assign n352 = n274 & n351 ;
  assign n353 = n352 ^ n274 ;
  assign n354 = n353 ^ n351 ;
  assign n355 = ~n350 & ~n354 ;
  assign n356 = n73 & n101 ;
  assign n357 = n356 ^ n73 ;
  assign n358 = n357 ^ n101 ;
  assign n359 = n88 & n97 ;
  assign n360 = n359 ^ n88 ;
  assign n361 = n360 ^ n97 ;
  assign n362 = ~n358 & ~n361 ;
  assign n363 = n355 & n362 ;
  assign n364 = n45 & ~n58 ;
  assign n365 = ~n113 & ~n116 ;
  assign n366 = ~n122 & n365 ;
  assign n367 = n364 & n366 ;
  assign n368 = n363 & n367 ;
  assign n369 = n346 & n368 ;
  assign n549 = n548 ^ n369 ;
  assign n234 = n199 & n233 ;
  assign n252 = n125 & n234 ;
  assign n253 = n252 ^ n125 ;
  assign n254 = n253 ^ n234 ;
  assign n256 = n40 & n255 ;
  assign n258 = n152 & n257 ;
  assign n259 = n256 & n258 ;
  assign n260 = n259 ^ n256 ;
  assign n261 = n260 ^ n258 ;
  assign n262 = ~n254 & ~n261 ;
  assign n263 = n136 & n150 ;
  assign n264 = n263 ^ n150 ;
  assign n265 = n264 ^ n136 ;
  assign n266 = n80 & n104 ;
  assign n267 = n266 ^ n80 ;
  assign n268 = n267 ^ n104 ;
  assign n269 = ~n265 & ~n268 ;
  assign n270 = n262 & n269 ;
  assign n272 = n129 & n271 ;
  assign n273 = n272 ^ n129 ;
  assign n275 = ~x13 & ~x19 ;
  assign n276 = n274 & n275 ;
  assign n277 = n276 ^ n274 ;
  assign n278 = n273 & n277 ;
  assign n279 = n278 ^ n273 ;
  assign n280 = n279 ^ n277 ;
  assign n282 = n121 & n281 ;
  assign n283 = n35 & n53 ;
  assign n284 = n282 & n283 ;
  assign n285 = n284 ^ n282 ;
  assign n286 = n285 ^ n283 ;
  assign n287 = ~n280 & ~n286 ;
  assign n288 = ~n192 & n287 ;
  assign n289 = n270 & n288 ;
  assign n290 = n112 & n116 ;
  assign n295 = n291 & ~n294 ;
  assign n296 = n295 ^ n291 ;
  assign n298 = n297 ^ n153 ;
  assign n299 = n297 ^ n67 ;
  assign n300 = ~n67 & n299 ;
  assign n301 = n300 ^ n67 ;
  assign n302 = n301 ^ n153 ;
  assign n303 = n298 & n302 ;
  assign n304 = n303 ^ n300 ;
  assign n305 = n304 ^ n153 ;
  assign n306 = n296 & n305 ;
  assign n307 = n306 ^ n296 ;
  assign n308 = n307 ^ n305 ;
  assign n309 = n290 & ~n308 ;
  assign n310 = n309 ^ n308 ;
  assign n311 = n175 & n197 ;
  assign n312 = n311 ^ n175 ;
  assign n313 = n312 ^ n197 ;
  assign n314 = n141 & n202 ;
  assign n315 = n314 ^ n141 ;
  assign n316 = n315 ^ n202 ;
  assign n317 = ~n313 & ~n316 ;
  assign n318 = ~n115 & ~n216 ;
  assign n319 = n317 & n318 ;
  assign n320 = ~n310 & n319 ;
  assign n321 = n289 & n320 ;
  assign n550 = n549 ^ n321 ;
  assign n226 = ~n48 & ~n62 ;
  assign n227 = ~n117 & n226 ;
  assign n228 = ~n206 & n211 ;
  assign n229 = n228 ^ n206 ;
  assign n230 = ~n157 & n217 ;
  assign n231 = n230 ^ n157 ;
  assign n232 = ~n229 & ~n231 ;
  assign n235 = n188 & n234 ;
  assign n236 = ~n105 & ~n123 ;
  assign n237 = ~n235 & n236 ;
  assign n238 = n90 & n99 ;
  assign n239 = n238 ^ n90 ;
  assign n240 = n239 ^ n99 ;
  assign n241 = n130 & ~n240 ;
  assign n242 = n241 ^ n240 ;
  assign n243 = n75 & n162 ;
  assign n244 = n243 ^ n75 ;
  assign n245 = n244 ^ n162 ;
  assign n246 = n180 & ~n245 ;
  assign n247 = n246 ^ n245 ;
  assign n248 = ~n242 & ~n247 ;
  assign n249 = n237 & n248 ;
  assign n250 = n232 & n249 ;
  assign n251 = n227 & n250 ;
  assign n551 = n550 ^ n251 ;
  assign n552 = n225 & n551 ;
  assign n553 = n552 ^ n225 ;
  assign n554 = n553 ^ n551 ;
  assign n567 = ~n429 & ~n519 ;
  assign n566 = n429 & ~n545 ;
  assign n568 = n567 ^ n566 ;
  assign n563 = ~n519 & n545 ;
  assign n564 = ~n490 & n563 ;
  assign n561 = ~n429 & ~n490 ;
  assign n559 = n519 & ~n545 ;
  assign n560 = n490 & n559 ;
  assign n562 = n561 ^ n560 ;
  assign n565 = n564 ^ n562 ;
  assign n569 = n568 ^ n565 ;
  assign n558 = n369 & ~n548 ;
  assign n570 = n569 ^ n558 ;
  assign n556 = n321 & n548 ;
  assign n555 = n321 & ~n369 ;
  assign n557 = n556 ^ n555 ;
  assign n571 = n570 ^ n557 ;
  assign n572 = ~n554 & n571 ;
  assign n573 = n572 ^ n554 ;
  assign n582 = n569 ^ n547 ;
  assign n574 = n346 & n366 ;
  assign n575 = n363 & n364 ;
  assign n578 = n429 & n575 ;
  assign n579 = n574 & n578 ;
  assign n576 = n547 & n575 ;
  assign n577 = n574 & n576 ;
  assign n580 = n579 ^ n577 ;
  assign n581 = n580 ^ n429 ;
  assign n583 = n582 ^ n581 ;
  assign n588 = n321 & n583 ;
  assign n589 = n588 ^ n583 ;
  assign n590 = n251 & n589 ;
  assign n591 = n590 ^ n589 ;
  assign n584 = n549 & n583 ;
  assign n585 = n584 ^ n583 ;
  assign n586 = n251 & n585 ;
  assign n587 = n586 ^ n585 ;
  assign n592 = n591 ^ n587 ;
  assign n599 = n369 & n548 ;
  assign n600 = n599 ^ n548 ;
  assign n594 = ~n490 & n519 ;
  assign n593 = n490 & n545 ;
  assign n595 = n594 ^ n593 ;
  assign n596 = n595 ^ n559 ;
  assign n601 = n569 & ~n596 ;
  assign n602 = n600 & n601 ;
  assign n603 = n602 ^ n601 ;
  assign n604 = n592 & n603 ;
  assign n605 = n604 ^ n603 ;
  assign n597 = n592 & n596 ;
  assign n598 = n597 ^ n596 ;
  assign n606 = n605 ^ n598 ;
  assign n607 = ~n573 & n606 ;
  assign n608 = n607 ^ n573 ;
  assign n609 = n569 ^ n549 ;
  assign n610 = ~n569 & ~n609 ;
  assign n611 = n610 ^ n549 ;
  assign n612 = n611 ^ n321 ;
  assign n613 = n321 & n612 ;
  assign n614 = n613 ^ n610 ;
  assign n615 = n614 ^ n549 ;
  assign n627 = n615 ^ n592 ;
  assign n628 = n603 ^ n596 ;
  assign n629 = ~n615 & n628 ;
  assign n630 = n629 ^ n592 ;
  assign n631 = n630 ^ n615 ;
  assign n632 = n631 ^ n628 ;
  assign n633 = ~n627 & ~n632 ;
  assign n634 = n633 ^ n629 ;
  assign n618 = n321 & n549 ;
  assign n619 = n618 ^ n321 ;
  assign n620 = n619 ^ n549 ;
  assign n621 = n583 ^ n569 ;
  assign n622 = ~n620 & n621 ;
  assign n623 = n622 ^ n583 ;
  assign n624 = n623 ^ n620 ;
  assign n625 = ~n554 & ~n624 ;
  assign n626 = n625 ^ n592 ;
  assign n635 = n634 ^ n626 ;
  assign n616 = n615 ^ n603 ;
  assign n617 = n616 ^ n596 ;
  assign n636 = n635 ^ n617 ;
  assign n637 = ~n251 & n550 ;
  assign n638 = n554 & ~n637 ;
  assign n639 = n638 ^ n571 ;
  assign n640 = n551 ^ n225 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = 1'b0 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = ~n608 ;
  assign y29 = n636 ;
  assign y30 = n639 ;
  assign y31 = n640 ;
endmodule
