module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 ;
  assign n185 = x132 & x133 ;
  assign n148 = ~x130 & ~x131 ;
  assign n386 = x80 & ~x128 ;
  assign n385 = x79 & x128 ;
  assign n387 = n386 ^ n385 ;
  assign n388 = ~x129 & n387 ;
  assign n382 = x78 & ~x128 ;
  assign n381 = x77 & x128 ;
  assign n383 = n382 ^ n381 ;
  assign n384 = x129 & n383 ;
  assign n389 = n388 ^ n384 ;
  assign n390 = n148 & n389 ;
  assign n137 = x130 & ~x131 ;
  assign n376 = x76 & ~x128 ;
  assign n375 = x75 & x128 ;
  assign n377 = n376 ^ n375 ;
  assign n378 = ~x129 & n377 ;
  assign n372 = x74 & ~x128 ;
  assign n371 = x73 & x128 ;
  assign n373 = n372 ^ n371 ;
  assign n374 = x129 & n373 ;
  assign n379 = n378 ^ n374 ;
  assign n380 = n137 & n379 ;
  assign n391 = n390 ^ n380 ;
  assign n171 = x130 & x131 ;
  assign n407 = x68 & ~x128 ;
  assign n406 = x67 & x128 ;
  assign n408 = n407 ^ n406 ;
  assign n409 = ~x129 & n408 ;
  assign n403 = x66 & ~x128 ;
  assign n402 = x65 & x128 ;
  assign n404 = n403 ^ n402 ;
  assign n405 = x129 & n404 ;
  assign n410 = n409 ^ n405 ;
  assign n411 = n171 & n410 ;
  assign n160 = ~x130 & x131 ;
  assign n397 = x72 & ~x128 ;
  assign n396 = x71 & x128 ;
  assign n398 = n397 ^ n396 ;
  assign n399 = ~x129 & n398 ;
  assign n393 = x70 & ~x128 ;
  assign n392 = x69 & x128 ;
  assign n394 = n393 ^ n392 ;
  assign n395 = x129 & n394 ;
  assign n400 = n399 ^ n395 ;
  assign n401 = n160 & n400 ;
  assign n412 = n411 ^ n401 ;
  assign n413 = ~n391 & ~n412 ;
  assign n414 = n185 & ~n413 ;
  assign n136 = ~x132 & x133 ;
  assign n342 = x96 & ~x128 ;
  assign n341 = x95 & x128 ;
  assign n343 = n342 ^ n341 ;
  assign n344 = ~x129 & n343 ;
  assign n338 = x94 & ~x128 ;
  assign n337 = x93 & x128 ;
  assign n339 = n338 ^ n337 ;
  assign n340 = x129 & n339 ;
  assign n345 = n344 ^ n340 ;
  assign n346 = n148 & n345 ;
  assign n332 = x92 & ~x128 ;
  assign n331 = x91 & x128 ;
  assign n333 = n332 ^ n331 ;
  assign n334 = ~x129 & n333 ;
  assign n328 = x90 & ~x128 ;
  assign n327 = x89 & x128 ;
  assign n329 = n328 ^ n327 ;
  assign n330 = x129 & n329 ;
  assign n335 = n334 ^ n330 ;
  assign n336 = n137 & n335 ;
  assign n347 = n346 ^ n336 ;
  assign n363 = x84 & ~x128 ;
  assign n362 = x83 & x128 ;
  assign n364 = n363 ^ n362 ;
  assign n365 = ~x129 & n364 ;
  assign n359 = x82 & ~x128 ;
  assign n358 = x81 & x128 ;
  assign n360 = n359 ^ n358 ;
  assign n361 = x129 & n360 ;
  assign n366 = n365 ^ n361 ;
  assign n367 = n171 & n366 ;
  assign n353 = x88 & ~x128 ;
  assign n352 = x87 & x128 ;
  assign n354 = n353 ^ n352 ;
  assign n355 = ~x129 & n354 ;
  assign n349 = x86 & ~x128 ;
  assign n348 = x85 & x128 ;
  assign n350 = n349 ^ n348 ;
  assign n351 = x129 & n350 ;
  assign n356 = n355 ^ n351 ;
  assign n357 = n160 & n356 ;
  assign n368 = n367 ^ n357 ;
  assign n369 = ~n347 & ~n368 ;
  assign n370 = n136 & ~n369 ;
  assign n415 = n414 ^ n370 ;
  assign n279 = ~x132 & ~x133 ;
  assign n475 = x127 & x128 ;
  assign n474 = x0 & ~x128 ;
  assign n476 = n475 ^ n474 ;
  assign n477 = ~x129 & n476 ;
  assign n471 = x126 & ~x128 ;
  assign n470 = x125 & x128 ;
  assign n472 = n471 ^ n470 ;
  assign n473 = x129 & n472 ;
  assign n478 = n477 ^ n473 ;
  assign n479 = n148 & n478 ;
  assign n465 = x124 & ~x128 ;
  assign n464 = x123 & x128 ;
  assign n466 = n465 ^ n464 ;
  assign n467 = ~x129 & n466 ;
  assign n461 = x122 & ~x128 ;
  assign n460 = x121 & x128 ;
  assign n462 = n461 ^ n460 ;
  assign n463 = x129 & n462 ;
  assign n468 = n467 ^ n463 ;
  assign n469 = n137 & n468 ;
  assign n480 = n479 ^ n469 ;
  assign n496 = x116 & ~x128 ;
  assign n495 = x115 & x128 ;
  assign n497 = n496 ^ n495 ;
  assign n498 = ~x129 & n497 ;
  assign n492 = x114 & ~x128 ;
  assign n491 = x113 & x128 ;
  assign n493 = n492 ^ n491 ;
  assign n494 = x129 & n493 ;
  assign n499 = n498 ^ n494 ;
  assign n500 = n171 & n499 ;
  assign n486 = x120 & ~x128 ;
  assign n485 = x119 & x128 ;
  assign n487 = n486 ^ n485 ;
  assign n488 = ~x129 & n487 ;
  assign n482 = x118 & ~x128 ;
  assign n481 = x117 & x128 ;
  assign n483 = n482 ^ n481 ;
  assign n484 = x129 & n483 ;
  assign n489 = n488 ^ n484 ;
  assign n490 = n160 & n489 ;
  assign n501 = n500 ^ n490 ;
  assign n502 = ~n480 & ~n501 ;
  assign n503 = n279 & ~n502 ;
  assign n254 = x132 & ~x133 ;
  assign n431 = x112 & ~x128 ;
  assign n430 = x111 & x128 ;
  assign n432 = n431 ^ n430 ;
  assign n433 = ~x129 & n432 ;
  assign n427 = x110 & ~x128 ;
  assign n426 = x109 & x128 ;
  assign n428 = n427 ^ n426 ;
  assign n429 = x129 & n428 ;
  assign n434 = n433 ^ n429 ;
  assign n435 = n148 & n434 ;
  assign n421 = x108 & ~x128 ;
  assign n420 = x107 & x128 ;
  assign n422 = n421 ^ n420 ;
  assign n423 = ~x129 & n422 ;
  assign n417 = x106 & ~x128 ;
  assign n416 = x105 & x128 ;
  assign n418 = n417 ^ n416 ;
  assign n419 = x129 & n418 ;
  assign n424 = n423 ^ n419 ;
  assign n425 = n137 & n424 ;
  assign n436 = n435 ^ n425 ;
  assign n452 = x100 & ~x128 ;
  assign n451 = x99 & x128 ;
  assign n453 = n452 ^ n451 ;
  assign n454 = ~x129 & n453 ;
  assign n448 = x98 & ~x128 ;
  assign n447 = x97 & x128 ;
  assign n449 = n448 ^ n447 ;
  assign n450 = x129 & n449 ;
  assign n455 = n454 ^ n450 ;
  assign n456 = n171 & n455 ;
  assign n442 = x104 & ~x128 ;
  assign n441 = x103 & x128 ;
  assign n443 = n442 ^ n441 ;
  assign n444 = ~x129 & n443 ;
  assign n438 = x102 & ~x128 ;
  assign n437 = x101 & x128 ;
  assign n439 = n438 ^ n437 ;
  assign n440 = x129 & n439 ;
  assign n445 = n444 ^ n440 ;
  assign n446 = n160 & n445 ;
  assign n457 = n456 ^ n446 ;
  assign n458 = ~n436 & ~n457 ;
  assign n459 = n254 & ~n458 ;
  assign n504 = n503 ^ n459 ;
  assign n505 = ~n415 & ~n504 ;
  assign n506 = ~x134 & n505 ;
  assign n201 = x16 & ~x128 ;
  assign n200 = x15 & x128 ;
  assign n202 = n201 ^ n200 ;
  assign n203 = ~x129 & n202 ;
  assign n197 = x14 & ~x128 ;
  assign n196 = x13 & x128 ;
  assign n198 = n197 ^ n196 ;
  assign n199 = x129 & n198 ;
  assign n204 = n203 ^ n199 ;
  assign n205 = n148 & n204 ;
  assign n191 = x12 & ~x128 ;
  assign n190 = x11 & x128 ;
  assign n192 = n191 ^ n190 ;
  assign n193 = ~x129 & n192 ;
  assign n187 = x10 & ~x128 ;
  assign n186 = x9 & x128 ;
  assign n188 = n187 ^ n186 ;
  assign n189 = x129 & n188 ;
  assign n194 = n193 ^ n189 ;
  assign n195 = n137 & n194 ;
  assign n206 = n205 ^ n195 ;
  assign n222 = x4 & ~x128 ;
  assign n221 = x3 & x128 ;
  assign n223 = n222 ^ n221 ;
  assign n224 = ~x129 & n223 ;
  assign n218 = x2 & ~x128 ;
  assign n217 = x1 & x128 ;
  assign n219 = n218 ^ n217 ;
  assign n220 = x129 & n219 ;
  assign n225 = n224 ^ n220 ;
  assign n226 = n171 & n225 ;
  assign n212 = x8 & ~x128 ;
  assign n211 = x7 & x128 ;
  assign n213 = n212 ^ n211 ;
  assign n214 = ~x129 & n213 ;
  assign n208 = x6 & ~x128 ;
  assign n207 = x5 & x128 ;
  assign n209 = n208 ^ n207 ;
  assign n210 = x129 & n209 ;
  assign n215 = n214 ^ n210 ;
  assign n216 = n160 & n215 ;
  assign n227 = n226 ^ n216 ;
  assign n228 = ~n206 & ~n227 ;
  assign n229 = n185 & ~n228 ;
  assign n154 = x32 & ~x128 ;
  assign n153 = x31 & x128 ;
  assign n155 = n154 ^ n153 ;
  assign n156 = ~x129 & n155 ;
  assign n150 = x30 & ~x128 ;
  assign n149 = x29 & x128 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = x129 & n151 ;
  assign n157 = n156 ^ n152 ;
  assign n158 = n148 & n157 ;
  assign n143 = x28 & ~x128 ;
  assign n142 = x27 & x128 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = ~x129 & n144 ;
  assign n139 = x26 & ~x128 ;
  assign n138 = x25 & x128 ;
  assign n140 = n139 ^ n138 ;
  assign n141 = x129 & n140 ;
  assign n146 = n145 ^ n141 ;
  assign n147 = n137 & n146 ;
  assign n159 = n158 ^ n147 ;
  assign n177 = x20 & ~x128 ;
  assign n176 = x19 & x128 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = ~x129 & n178 ;
  assign n173 = x18 & ~x128 ;
  assign n172 = x17 & x128 ;
  assign n174 = n173 ^ n172 ;
  assign n175 = x129 & n174 ;
  assign n180 = n179 ^ n175 ;
  assign n181 = n171 & n180 ;
  assign n166 = x24 & ~x128 ;
  assign n165 = x23 & x128 ;
  assign n167 = n166 ^ n165 ;
  assign n168 = ~x129 & n167 ;
  assign n162 = x22 & ~x128 ;
  assign n161 = x21 & x128 ;
  assign n163 = n162 ^ n161 ;
  assign n164 = x129 & n163 ;
  assign n169 = n168 ^ n164 ;
  assign n170 = n160 & n169 ;
  assign n182 = n181 ^ n170 ;
  assign n183 = ~n159 & ~n182 ;
  assign n184 = n136 & ~n183 ;
  assign n230 = n229 ^ n184 ;
  assign n295 = x64 & ~x128 ;
  assign n294 = x63 & x128 ;
  assign n296 = n295 ^ n294 ;
  assign n297 = ~x129 & n296 ;
  assign n291 = x62 & ~x128 ;
  assign n290 = x61 & x128 ;
  assign n292 = n291 ^ n290 ;
  assign n293 = x129 & n292 ;
  assign n298 = n297 ^ n293 ;
  assign n299 = n148 & n298 ;
  assign n285 = x60 & ~x128 ;
  assign n284 = x59 & x128 ;
  assign n286 = n285 ^ n284 ;
  assign n287 = ~x129 & n286 ;
  assign n281 = x58 & ~x128 ;
  assign n280 = x57 & x128 ;
  assign n282 = n281 ^ n280 ;
  assign n283 = x129 & n282 ;
  assign n288 = n287 ^ n283 ;
  assign n289 = n137 & n288 ;
  assign n300 = n299 ^ n289 ;
  assign n316 = x52 & ~x128 ;
  assign n315 = x51 & x128 ;
  assign n317 = n316 ^ n315 ;
  assign n318 = ~x129 & n317 ;
  assign n312 = x50 & ~x128 ;
  assign n311 = x49 & x128 ;
  assign n313 = n312 ^ n311 ;
  assign n314 = x129 & n313 ;
  assign n319 = n318 ^ n314 ;
  assign n320 = n171 & n319 ;
  assign n306 = x56 & ~x128 ;
  assign n305 = x55 & x128 ;
  assign n307 = n306 ^ n305 ;
  assign n308 = ~x129 & n307 ;
  assign n302 = x54 & ~x128 ;
  assign n301 = x53 & x128 ;
  assign n303 = n302 ^ n301 ;
  assign n304 = x129 & n303 ;
  assign n309 = n308 ^ n304 ;
  assign n310 = n160 & n309 ;
  assign n321 = n320 ^ n310 ;
  assign n322 = ~n300 & ~n321 ;
  assign n323 = n279 & n322 ;
  assign n248 = x36 & ~x128 ;
  assign n247 = x35 & x128 ;
  assign n249 = n248 ^ n247 ;
  assign n250 = ~x129 & n249 ;
  assign n244 = x34 & ~x128 ;
  assign n243 = x33 & x128 ;
  assign n245 = n244 ^ n243 ;
  assign n246 = x129 & n245 ;
  assign n251 = n250 ^ n246 ;
  assign n252 = n171 & n251 ;
  assign n233 = x39 & x128 ;
  assign n234 = ~x129 & n233 ;
  assign n231 = x38 & ~x128 ;
  assign n232 = x129 & n231 ;
  assign n235 = n234 ^ n232 ;
  assign n238 = x40 & ~x128 ;
  assign n239 = ~x129 & ~n238 ;
  assign n236 = x37 & x128 ;
  assign n237 = x129 & ~n236 ;
  assign n240 = n239 ^ n237 ;
  assign n241 = ~n235 & n240 ;
  assign n242 = n160 & ~n241 ;
  assign n253 = n252 ^ n242 ;
  assign n270 = x48 & ~x128 ;
  assign n269 = x47 & x128 ;
  assign n271 = n270 ^ n269 ;
  assign n272 = ~x129 & n271 ;
  assign n266 = x46 & ~x128 ;
  assign n265 = x45 & x128 ;
  assign n267 = n266 ^ n265 ;
  assign n268 = x129 & n267 ;
  assign n273 = n272 ^ n268 ;
  assign n274 = n148 & n273 ;
  assign n260 = x44 & ~x128 ;
  assign n259 = x43 & x128 ;
  assign n261 = n260 ^ n259 ;
  assign n262 = ~x129 & n261 ;
  assign n256 = x42 & ~x128 ;
  assign n255 = x41 & x128 ;
  assign n257 = n256 ^ n255 ;
  assign n258 = x129 & n257 ;
  assign n263 = n262 ^ n258 ;
  assign n264 = n137 & n263 ;
  assign n275 = n274 ^ n264 ;
  assign n276 = n254 & ~n275 ;
  assign n277 = ~n253 & n276 ;
  assign n278 = n277 ^ x133 ;
  assign n324 = n323 ^ n278 ;
  assign n325 = ~n230 & n324 ;
  assign n326 = x134 & n325 ;
  assign n507 = n506 ^ n326 ;
  assign n913 = x80 & x128 ;
  assign n914 = x129 & n913 ;
  assign n915 = n914 ^ n913 ;
  assign n911 = n385 ^ x79 ;
  assign n912 = x129 & n911 ;
  assign n916 = n915 ^ n912 ;
  assign n920 = n358 ^ x81 ;
  assign n921 = x129 & n920 ;
  assign n922 = n921 ^ x129 ;
  assign n923 = n922 ^ n920 ;
  assign n917 = x78 & x128 ;
  assign n918 = x129 & n917 ;
  assign n919 = n918 ^ x129 ;
  assign n924 = n923 ^ n919 ;
  assign n925 = n916 & ~n924 ;
  assign n926 = n925 ^ n924 ;
  assign n927 = n148 & ~n926 ;
  assign n928 = n927 ^ n148 ;
  assign n895 = x76 & x128 ;
  assign n896 = x129 & n895 ;
  assign n897 = n896 ^ n895 ;
  assign n893 = n375 ^ x75 ;
  assign n894 = x129 & n893 ;
  assign n898 = n897 ^ n894 ;
  assign n902 = n381 ^ x77 ;
  assign n903 = x129 & n902 ;
  assign n904 = n903 ^ x129 ;
  assign n905 = n904 ^ n902 ;
  assign n899 = x74 & x128 ;
  assign n900 = x129 & n899 ;
  assign n901 = n900 ^ x129 ;
  assign n906 = n905 ^ n901 ;
  assign n907 = n898 & ~n906 ;
  assign n908 = n907 ^ n906 ;
  assign n909 = n137 & ~n908 ;
  assign n910 = n909 ^ n137 ;
  assign n929 = n928 ^ n910 ;
  assign n950 = x68 & x128 ;
  assign n951 = x129 & n950 ;
  assign n952 = n951 ^ n950 ;
  assign n948 = n406 ^ x67 ;
  assign n949 = x129 & n948 ;
  assign n953 = n952 ^ n949 ;
  assign n957 = n392 ^ x69 ;
  assign n958 = x129 & n957 ;
  assign n959 = n958 ^ x129 ;
  assign n960 = n959 ^ n957 ;
  assign n954 = x66 & x128 ;
  assign n955 = x129 & n954 ;
  assign n956 = n955 ^ x129 ;
  assign n961 = n960 ^ n956 ;
  assign n962 = n953 & ~n961 ;
  assign n963 = n962 ^ n961 ;
  assign n964 = n171 & ~n963 ;
  assign n965 = n964 ^ n171 ;
  assign n932 = x72 & x128 ;
  assign n933 = x129 & n932 ;
  assign n934 = n933 ^ n932 ;
  assign n930 = n396 ^ x71 ;
  assign n931 = x129 & n930 ;
  assign n935 = n934 ^ n931 ;
  assign n939 = n371 ^ x73 ;
  assign n940 = x129 & n939 ;
  assign n941 = n940 ^ x129 ;
  assign n942 = n941 ^ n939 ;
  assign n936 = x70 & x128 ;
  assign n937 = x129 & n936 ;
  assign n938 = n937 ^ x129 ;
  assign n943 = n942 ^ n938 ;
  assign n944 = n935 & ~n943 ;
  assign n945 = n944 ^ n943 ;
  assign n946 = n160 & ~n945 ;
  assign n947 = n946 ^ n160 ;
  assign n966 = n965 ^ n947 ;
  assign n967 = n929 & n966 ;
  assign n968 = n967 ^ n929 ;
  assign n969 = n968 ^ n966 ;
  assign n970 = n185 & ~n969 ;
  assign n971 = n970 ^ n185 ;
  assign n834 = x96 & x128 ;
  assign n835 = x129 & n834 ;
  assign n836 = n835 ^ n834 ;
  assign n832 = n341 ^ x95 ;
  assign n833 = x129 & n832 ;
  assign n837 = n836 ^ n833 ;
  assign n841 = n447 ^ x97 ;
  assign n842 = x129 & n841 ;
  assign n843 = n842 ^ x129 ;
  assign n844 = n843 ^ n841 ;
  assign n838 = x94 & x128 ;
  assign n839 = x129 & n838 ;
  assign n840 = n839 ^ x129 ;
  assign n845 = n844 ^ n840 ;
  assign n846 = n837 & ~n845 ;
  assign n847 = n846 ^ n845 ;
  assign n848 = n148 & ~n847 ;
  assign n849 = n848 ^ n148 ;
  assign n816 = x92 & x128 ;
  assign n817 = x129 & n816 ;
  assign n818 = n817 ^ n816 ;
  assign n814 = n331 ^ x91 ;
  assign n815 = x129 & n814 ;
  assign n819 = n818 ^ n815 ;
  assign n823 = n337 ^ x93 ;
  assign n824 = x129 & n823 ;
  assign n825 = n824 ^ x129 ;
  assign n826 = n825 ^ n823 ;
  assign n820 = x90 & x128 ;
  assign n821 = x129 & n820 ;
  assign n822 = n821 ^ x129 ;
  assign n827 = n826 ^ n822 ;
  assign n828 = n819 & ~n827 ;
  assign n829 = n828 ^ n827 ;
  assign n830 = n137 & ~n829 ;
  assign n831 = n830 ^ n137 ;
  assign n850 = n849 ^ n831 ;
  assign n871 = x84 & x128 ;
  assign n872 = x129 & n871 ;
  assign n873 = n872 ^ n871 ;
  assign n869 = n362 ^ x83 ;
  assign n870 = x129 & n869 ;
  assign n874 = n873 ^ n870 ;
  assign n878 = n348 ^ x85 ;
  assign n879 = x129 & n878 ;
  assign n880 = n879 ^ x129 ;
  assign n881 = n880 ^ n878 ;
  assign n875 = x82 & x128 ;
  assign n876 = x129 & n875 ;
  assign n877 = n876 ^ x129 ;
  assign n882 = n881 ^ n877 ;
  assign n883 = n874 & ~n882 ;
  assign n884 = n883 ^ n882 ;
  assign n885 = n171 & ~n884 ;
  assign n886 = n885 ^ n171 ;
  assign n853 = x88 & x128 ;
  assign n854 = x129 & n853 ;
  assign n855 = n854 ^ n853 ;
  assign n851 = n352 ^ x87 ;
  assign n852 = x129 & n851 ;
  assign n856 = n855 ^ n852 ;
  assign n860 = n327 ^ x89 ;
  assign n861 = x129 & n860 ;
  assign n862 = n861 ^ x129 ;
  assign n863 = n862 ^ n860 ;
  assign n857 = x86 & x128 ;
  assign n858 = x129 & n857 ;
  assign n859 = n858 ^ x129 ;
  assign n864 = n863 ^ n859 ;
  assign n865 = n856 & ~n864 ;
  assign n866 = n865 ^ n864 ;
  assign n867 = n160 & ~n866 ;
  assign n868 = n867 ^ n160 ;
  assign n887 = n886 ^ n868 ;
  assign n888 = n850 & n887 ;
  assign n889 = n888 ^ n850 ;
  assign n890 = n889 ^ n887 ;
  assign n891 = n136 & ~n890 ;
  assign n892 = n891 ^ n136 ;
  assign n972 = n971 ^ n892 ;
  assign n1072 = x0 & x128 ;
  assign n1073 = x129 & n1072 ;
  assign n1074 = n1073 ^ n1072 ;
  assign n1070 = n475 ^ x127 ;
  assign n1071 = x129 & n1070 ;
  assign n1075 = n1074 ^ n1071 ;
  assign n1079 = n217 ^ x1 ;
  assign n1080 = x129 & n1079 ;
  assign n1081 = n1080 ^ x129 ;
  assign n1082 = n1081 ^ n1079 ;
  assign n1076 = x126 & x128 ;
  assign n1077 = x129 & n1076 ;
  assign n1078 = n1077 ^ x129 ;
  assign n1083 = n1082 ^ n1078 ;
  assign n1084 = n1075 & ~n1083 ;
  assign n1085 = n1084 ^ n1083 ;
  assign n1086 = n148 & ~n1085 ;
  assign n1087 = n1086 ^ n148 ;
  assign n1054 = x124 & x128 ;
  assign n1055 = x129 & n1054 ;
  assign n1056 = n1055 ^ n1054 ;
  assign n1052 = n464 ^ x123 ;
  assign n1053 = x129 & n1052 ;
  assign n1057 = n1056 ^ n1053 ;
  assign n1061 = n470 ^ x125 ;
  assign n1062 = x129 & n1061 ;
  assign n1063 = n1062 ^ x129 ;
  assign n1064 = n1063 ^ n1061 ;
  assign n1058 = x122 & x128 ;
  assign n1059 = x129 & n1058 ;
  assign n1060 = n1059 ^ x129 ;
  assign n1065 = n1064 ^ n1060 ;
  assign n1066 = n1057 & ~n1065 ;
  assign n1067 = n1066 ^ n1065 ;
  assign n1068 = n137 & ~n1067 ;
  assign n1069 = n1068 ^ n137 ;
  assign n1088 = n1087 ^ n1069 ;
  assign n1109 = x116 & x128 ;
  assign n1110 = x129 & n1109 ;
  assign n1111 = n1110 ^ n1109 ;
  assign n1107 = n495 ^ x115 ;
  assign n1108 = x129 & n1107 ;
  assign n1112 = n1111 ^ n1108 ;
  assign n1116 = n481 ^ x117 ;
  assign n1117 = x129 & n1116 ;
  assign n1118 = n1117 ^ x129 ;
  assign n1119 = n1118 ^ n1116 ;
  assign n1113 = x114 & x128 ;
  assign n1114 = x129 & n1113 ;
  assign n1115 = n1114 ^ x129 ;
  assign n1120 = n1119 ^ n1115 ;
  assign n1121 = n1112 & ~n1120 ;
  assign n1122 = n1121 ^ n1120 ;
  assign n1123 = n171 & ~n1122 ;
  assign n1124 = n1123 ^ n171 ;
  assign n1091 = x120 & x128 ;
  assign n1092 = x129 & n1091 ;
  assign n1093 = n1092 ^ n1091 ;
  assign n1089 = n485 ^ x119 ;
  assign n1090 = x129 & n1089 ;
  assign n1094 = n1093 ^ n1090 ;
  assign n1098 = n460 ^ x121 ;
  assign n1099 = x129 & n1098 ;
  assign n1100 = n1099 ^ x129 ;
  assign n1101 = n1100 ^ n1098 ;
  assign n1095 = x118 & x128 ;
  assign n1096 = x129 & n1095 ;
  assign n1097 = n1096 ^ x129 ;
  assign n1102 = n1101 ^ n1097 ;
  assign n1103 = n1094 & ~n1102 ;
  assign n1104 = n1103 ^ n1102 ;
  assign n1105 = n160 & ~n1104 ;
  assign n1106 = n1105 ^ n160 ;
  assign n1125 = n1124 ^ n1106 ;
  assign n1126 = n1088 & n1125 ;
  assign n1127 = n1126 ^ n1088 ;
  assign n1128 = n1127 ^ n1125 ;
  assign n1129 = n279 & ~n1128 ;
  assign n1130 = n1129 ^ n279 ;
  assign n993 = x112 & x128 ;
  assign n994 = x129 & n993 ;
  assign n995 = n994 ^ n993 ;
  assign n991 = n430 ^ x111 ;
  assign n992 = x129 & n991 ;
  assign n996 = n995 ^ n992 ;
  assign n1000 = n491 ^ x113 ;
  assign n1001 = x129 & n1000 ;
  assign n1002 = n1001 ^ x129 ;
  assign n1003 = n1002 ^ n1000 ;
  assign n997 = x110 & x128 ;
  assign n998 = x129 & n997 ;
  assign n999 = n998 ^ x129 ;
  assign n1004 = n1003 ^ n999 ;
  assign n1005 = n996 & ~n1004 ;
  assign n1006 = n1005 ^ n1004 ;
  assign n1007 = n148 & ~n1006 ;
  assign n1008 = n1007 ^ n148 ;
  assign n975 = x108 & x128 ;
  assign n976 = x129 & n975 ;
  assign n977 = n976 ^ n975 ;
  assign n973 = n420 ^ x107 ;
  assign n974 = x129 & n973 ;
  assign n978 = n977 ^ n974 ;
  assign n982 = n426 ^ x109 ;
  assign n983 = x129 & n982 ;
  assign n984 = n983 ^ x129 ;
  assign n985 = n984 ^ n982 ;
  assign n979 = x106 & x128 ;
  assign n980 = x129 & n979 ;
  assign n981 = n980 ^ x129 ;
  assign n986 = n985 ^ n981 ;
  assign n987 = n978 & ~n986 ;
  assign n988 = n987 ^ n986 ;
  assign n989 = n137 & ~n988 ;
  assign n990 = n989 ^ n137 ;
  assign n1009 = n1008 ^ n990 ;
  assign n1030 = x100 & x128 ;
  assign n1031 = x129 & n1030 ;
  assign n1032 = n1031 ^ n1030 ;
  assign n1028 = n451 ^ x99 ;
  assign n1029 = x129 & n1028 ;
  assign n1033 = n1032 ^ n1029 ;
  assign n1037 = n437 ^ x101 ;
  assign n1038 = x129 & n1037 ;
  assign n1039 = n1038 ^ x129 ;
  assign n1040 = n1039 ^ n1037 ;
  assign n1034 = x98 & x128 ;
  assign n1035 = x129 & n1034 ;
  assign n1036 = n1035 ^ x129 ;
  assign n1041 = n1040 ^ n1036 ;
  assign n1042 = n1033 & ~n1041 ;
  assign n1043 = n1042 ^ n1041 ;
  assign n1044 = n171 & ~n1043 ;
  assign n1045 = n1044 ^ n171 ;
  assign n1012 = x104 & x128 ;
  assign n1013 = x129 & n1012 ;
  assign n1014 = n1013 ^ n1012 ;
  assign n1010 = n441 ^ x103 ;
  assign n1011 = x129 & n1010 ;
  assign n1015 = n1014 ^ n1011 ;
  assign n1019 = n416 ^ x105 ;
  assign n1020 = x129 & n1019 ;
  assign n1021 = n1020 ^ x129 ;
  assign n1022 = n1021 ^ n1019 ;
  assign n1016 = x102 & x128 ;
  assign n1017 = x129 & n1016 ;
  assign n1018 = n1017 ^ x129 ;
  assign n1023 = n1022 ^ n1018 ;
  assign n1024 = n1015 & ~n1023 ;
  assign n1025 = n1024 ^ n1023 ;
  assign n1026 = n160 & ~n1025 ;
  assign n1027 = n1026 ^ n160 ;
  assign n1046 = n1045 ^ n1027 ;
  assign n1047 = n1009 & n1046 ;
  assign n1048 = n1047 ^ n1009 ;
  assign n1049 = n1048 ^ n1046 ;
  assign n1050 = n254 & ~n1049 ;
  assign n1051 = n1050 ^ n254 ;
  assign n1131 = n1130 ^ n1051 ;
  assign n1132 = n972 & n1131 ;
  assign n1133 = n1132 ^ n972 ;
  assign n1134 = n1133 ^ n1131 ;
  assign n1135 = x134 & ~n1134 ;
  assign n1136 = n1135 ^ n1134 ;
  assign n607 = x64 & x128 ;
  assign n608 = x129 & n607 ;
  assign n609 = n608 ^ n607 ;
  assign n605 = n294 ^ x63 ;
  assign n606 = x129 & n605 ;
  assign n610 = n609 ^ n606 ;
  assign n614 = n402 ^ x65 ;
  assign n615 = x129 & n614 ;
  assign n616 = n615 ^ x129 ;
  assign n617 = n616 ^ n614 ;
  assign n611 = x62 & x128 ;
  assign n612 = x129 & n611 ;
  assign n613 = n612 ^ x129 ;
  assign n618 = n617 ^ n613 ;
  assign n619 = n610 & ~n618 ;
  assign n620 = n619 ^ n618 ;
  assign n621 = n148 & ~n620 ;
  assign n622 = n621 ^ n148 ;
  assign n589 = x60 & x128 ;
  assign n590 = x129 & n589 ;
  assign n591 = n590 ^ n589 ;
  assign n587 = n284 ^ x59 ;
  assign n588 = x129 & n587 ;
  assign n592 = n591 ^ n588 ;
  assign n596 = n290 ^ x61 ;
  assign n597 = x129 & n596 ;
  assign n598 = n597 ^ x129 ;
  assign n599 = n598 ^ n596 ;
  assign n593 = x58 & x128 ;
  assign n594 = x129 & n593 ;
  assign n595 = n594 ^ x129 ;
  assign n600 = n599 ^ n595 ;
  assign n601 = n592 & ~n600 ;
  assign n602 = n601 ^ n600 ;
  assign n603 = n137 & ~n602 ;
  assign n604 = n603 ^ n137 ;
  assign n623 = n622 ^ n604 ;
  assign n644 = x52 & x128 ;
  assign n645 = x129 & n644 ;
  assign n646 = n645 ^ n644 ;
  assign n642 = n315 ^ x51 ;
  assign n643 = x129 & n642 ;
  assign n647 = n646 ^ n643 ;
  assign n651 = n301 ^ x53 ;
  assign n652 = x129 & n651 ;
  assign n653 = n652 ^ x129 ;
  assign n654 = n653 ^ n651 ;
  assign n648 = x50 & x128 ;
  assign n649 = x129 & n648 ;
  assign n650 = n649 ^ x129 ;
  assign n655 = n654 ^ n650 ;
  assign n656 = n647 & ~n655 ;
  assign n657 = n656 ^ n655 ;
  assign n658 = n171 & ~n657 ;
  assign n659 = n658 ^ n171 ;
  assign n626 = x56 & x128 ;
  assign n627 = x129 & n626 ;
  assign n628 = n627 ^ n626 ;
  assign n624 = n305 ^ x55 ;
  assign n625 = x129 & n624 ;
  assign n629 = n628 ^ n625 ;
  assign n633 = n280 ^ x57 ;
  assign n634 = x129 & n633 ;
  assign n635 = n634 ^ x129 ;
  assign n636 = n635 ^ n633 ;
  assign n630 = x54 & x128 ;
  assign n631 = x129 & n630 ;
  assign n632 = n631 ^ x129 ;
  assign n637 = n636 ^ n632 ;
  assign n638 = n629 & ~n637 ;
  assign n639 = n638 ^ n637 ;
  assign n640 = n160 & ~n639 ;
  assign n641 = n640 ^ n160 ;
  assign n660 = n659 ^ n641 ;
  assign n661 = n623 & n660 ;
  assign n662 = n661 ^ n623 ;
  assign n663 = n662 ^ n660 ;
  assign n664 = n279 & ~n663 ;
  assign n665 = n664 ^ n279 ;
  assign n528 = x16 & x128 ;
  assign n529 = x129 & n528 ;
  assign n530 = n529 ^ n528 ;
  assign n526 = n200 ^ x15 ;
  assign n527 = x129 & n526 ;
  assign n531 = n530 ^ n527 ;
  assign n535 = n172 ^ x17 ;
  assign n536 = x129 & n535 ;
  assign n537 = n536 ^ x129 ;
  assign n538 = n537 ^ n535 ;
  assign n532 = x14 & x128 ;
  assign n533 = x129 & n532 ;
  assign n534 = n533 ^ x129 ;
  assign n539 = n538 ^ n534 ;
  assign n540 = n531 & ~n539 ;
  assign n541 = n540 ^ n539 ;
  assign n542 = n148 & ~n541 ;
  assign n543 = n542 ^ n148 ;
  assign n510 = x12 & x128 ;
  assign n511 = x129 & n510 ;
  assign n512 = n511 ^ n510 ;
  assign n508 = n190 ^ x11 ;
  assign n509 = x129 & n508 ;
  assign n513 = n512 ^ n509 ;
  assign n517 = n196 ^ x13 ;
  assign n518 = x129 & n517 ;
  assign n519 = n518 ^ x129 ;
  assign n520 = n519 ^ n517 ;
  assign n514 = x10 & x128 ;
  assign n515 = x129 & n514 ;
  assign n516 = n515 ^ x129 ;
  assign n521 = n520 ^ n516 ;
  assign n522 = n513 & ~n521 ;
  assign n523 = n522 ^ n521 ;
  assign n524 = n137 & ~n523 ;
  assign n525 = n524 ^ n137 ;
  assign n544 = n543 ^ n525 ;
  assign n565 = x4 & x128 ;
  assign n566 = x129 & n565 ;
  assign n567 = n566 ^ n565 ;
  assign n563 = n221 ^ x3 ;
  assign n564 = x129 & n563 ;
  assign n568 = n567 ^ n564 ;
  assign n572 = n207 ^ x5 ;
  assign n573 = x129 & n572 ;
  assign n574 = n573 ^ x129 ;
  assign n575 = n574 ^ n572 ;
  assign n569 = x2 & x128 ;
  assign n570 = x129 & n569 ;
  assign n571 = n570 ^ x129 ;
  assign n576 = n575 ^ n571 ;
  assign n577 = n568 & ~n576 ;
  assign n578 = n577 ^ n576 ;
  assign n579 = n171 & ~n578 ;
  assign n580 = n579 ^ n171 ;
  assign n547 = x8 & x128 ;
  assign n548 = x129 & n547 ;
  assign n549 = n548 ^ n547 ;
  assign n545 = n211 ^ x7 ;
  assign n546 = x129 & n545 ;
  assign n550 = n549 ^ n546 ;
  assign n554 = n186 ^ x9 ;
  assign n555 = x129 & n554 ;
  assign n556 = n555 ^ x129 ;
  assign n557 = n556 ^ n554 ;
  assign n551 = x6 & x128 ;
  assign n552 = x129 & n551 ;
  assign n553 = n552 ^ x129 ;
  assign n558 = n557 ^ n553 ;
  assign n559 = n550 & ~n558 ;
  assign n560 = n559 ^ n558 ;
  assign n561 = n160 & ~n560 ;
  assign n562 = n561 ^ n160 ;
  assign n581 = n580 ^ n562 ;
  assign n582 = n544 & n581 ;
  assign n583 = n582 ^ n544 ;
  assign n584 = n583 ^ n581 ;
  assign n585 = n185 & ~n584 ;
  assign n586 = n585 ^ n185 ;
  assign n666 = n665 ^ n586 ;
  assign n758 = x48 & x128 ;
  assign n759 = x129 & n758 ;
  assign n760 = n759 ^ n758 ;
  assign n756 = n269 ^ x47 ;
  assign n757 = x129 & n756 ;
  assign n761 = n760 ^ n757 ;
  assign n765 = n311 ^ x49 ;
  assign n766 = x129 & n765 ;
  assign n767 = n766 ^ x129 ;
  assign n768 = n767 ^ n765 ;
  assign n762 = x46 & x128 ;
  assign n763 = x129 & n762 ;
  assign n764 = n763 ^ x129 ;
  assign n769 = n768 ^ n764 ;
  assign n770 = n761 & ~n769 ;
  assign n771 = n770 ^ n769 ;
  assign n772 = n148 & ~n771 ;
  assign n773 = n772 ^ n148 ;
  assign n751 = x45 & ~x128 ;
  assign n750 = x44 & x128 ;
  assign n752 = n751 ^ n750 ;
  assign n753 = ~x129 & ~n752 ;
  assign n747 = ~x43 & ~x128 ;
  assign n746 = ~x42 & x128 ;
  assign n748 = n747 ^ n746 ;
  assign n749 = x129 & n748 ;
  assign n754 = n753 ^ n749 ;
  assign n755 = n137 & ~n754 ;
  assign n774 = n773 ^ n755 ;
  assign n787 = x36 & x128 ;
  assign n788 = x129 & n787 ;
  assign n789 = n788 ^ n787 ;
  assign n785 = n247 ^ x35 ;
  assign n786 = x129 & n785 ;
  assign n790 = n789 ^ n786 ;
  assign n794 = n236 ^ x37 ;
  assign n795 = x129 & n794 ;
  assign n796 = n795 ^ x129 ;
  assign n797 = n796 ^ n794 ;
  assign n791 = x34 & x128 ;
  assign n792 = x129 & n791 ;
  assign n793 = n792 ^ x129 ;
  assign n798 = n797 ^ n793 ;
  assign n799 = n790 & ~n798 ;
  assign n800 = n799 ^ n798 ;
  assign n801 = n171 & ~n800 ;
  assign n802 = n801 ^ n171 ;
  assign n780 = ~x41 & ~x128 ;
  assign n779 = ~x40 & x128 ;
  assign n781 = n780 ^ n779 ;
  assign n782 = ~x129 & n781 ;
  assign n776 = ~x39 & ~x128 ;
  assign n775 = ~x38 & x128 ;
  assign n777 = n776 ^ n775 ;
  assign n778 = x129 & n777 ;
  assign n783 = n782 ^ n778 ;
  assign n784 = n160 & ~n783 ;
  assign n803 = n802 ^ n784 ;
  assign n804 = n774 & n803 ;
  assign n805 = n804 ^ n774 ;
  assign n806 = n805 ^ n803 ;
  assign n807 = n254 & ~n806 ;
  assign n808 = n807 ^ n254 ;
  assign n687 = x32 & x128 ;
  assign n688 = x129 & n687 ;
  assign n689 = n688 ^ n687 ;
  assign n685 = n153 ^ x31 ;
  assign n686 = x129 & n685 ;
  assign n690 = n689 ^ n686 ;
  assign n694 = n243 ^ x33 ;
  assign n695 = x129 & n694 ;
  assign n696 = n695 ^ x129 ;
  assign n697 = n696 ^ n694 ;
  assign n691 = x30 & x128 ;
  assign n692 = x129 & n691 ;
  assign n693 = n692 ^ x129 ;
  assign n698 = n697 ^ n693 ;
  assign n699 = n690 & ~n698 ;
  assign n700 = n699 ^ n698 ;
  assign n701 = n148 & ~n700 ;
  assign n702 = n701 ^ n148 ;
  assign n669 = x28 & x128 ;
  assign n670 = x129 & n669 ;
  assign n671 = n670 ^ n669 ;
  assign n667 = n142 ^ x27 ;
  assign n668 = x129 & n667 ;
  assign n672 = n671 ^ n668 ;
  assign n676 = n149 ^ x29 ;
  assign n677 = x129 & n676 ;
  assign n678 = n677 ^ x129 ;
  assign n679 = n678 ^ n676 ;
  assign n673 = x26 & x128 ;
  assign n674 = x129 & n673 ;
  assign n675 = n674 ^ x129 ;
  assign n680 = n679 ^ n675 ;
  assign n681 = n672 & ~n680 ;
  assign n682 = n681 ^ n680 ;
  assign n683 = n137 & ~n682 ;
  assign n684 = n683 ^ n137 ;
  assign n703 = n702 ^ n684 ;
  assign n724 = x20 & x128 ;
  assign n725 = x129 & n724 ;
  assign n726 = n725 ^ n724 ;
  assign n722 = n176 ^ x19 ;
  assign n723 = x129 & n722 ;
  assign n727 = n726 ^ n723 ;
  assign n731 = n161 ^ x21 ;
  assign n732 = x129 & n731 ;
  assign n733 = n732 ^ x129 ;
  assign n734 = n733 ^ n731 ;
  assign n728 = x18 & x128 ;
  assign n729 = x129 & n728 ;
  assign n730 = n729 ^ x129 ;
  assign n735 = n734 ^ n730 ;
  assign n736 = n727 & ~n735 ;
  assign n737 = n736 ^ n735 ;
  assign n738 = n171 & ~n737 ;
  assign n739 = n738 ^ n171 ;
  assign n706 = x24 & x128 ;
  assign n707 = x129 & n706 ;
  assign n708 = n707 ^ n706 ;
  assign n704 = n165 ^ x23 ;
  assign n705 = x129 & n704 ;
  assign n709 = n708 ^ n705 ;
  assign n713 = n138 ^ x25 ;
  assign n714 = x129 & n713 ;
  assign n715 = n714 ^ x129 ;
  assign n716 = n715 ^ n713 ;
  assign n710 = x22 & x128 ;
  assign n711 = x129 & n710 ;
  assign n712 = n711 ^ x129 ;
  assign n717 = n716 ^ n712 ;
  assign n718 = n709 & ~n717 ;
  assign n719 = n718 ^ n717 ;
  assign n720 = n160 & ~n719 ;
  assign n721 = n720 ^ n160 ;
  assign n740 = n739 ^ n721 ;
  assign n741 = n703 & n740 ;
  assign n742 = n741 ^ n703 ;
  assign n743 = n742 ^ n740 ;
  assign n744 = n136 & ~n743 ;
  assign n745 = n744 ^ n136 ;
  assign n809 = n808 ^ n745 ;
  assign n810 = n666 & n809 ;
  assign n811 = n810 ^ n666 ;
  assign n812 = n811 ^ n809 ;
  assign n813 = x134 & ~n812 ;
  assign n1137 = n1136 ^ n813 ;
  assign n1253 = ~x129 & n360 ;
  assign n1252 = x129 & n387 ;
  assign n1254 = n1253 ^ n1252 ;
  assign n1255 = n148 & n1254 ;
  assign n1249 = ~x129 & n383 ;
  assign n1248 = x129 & n377 ;
  assign n1250 = n1249 ^ n1248 ;
  assign n1251 = n137 & n1250 ;
  assign n1256 = n1255 ^ n1251 ;
  assign n1262 = ~x129 & n394 ;
  assign n1261 = x129 & n408 ;
  assign n1263 = n1262 ^ n1261 ;
  assign n1264 = n171 & n1263 ;
  assign n1258 = ~x129 & n373 ;
  assign n1257 = x129 & n398 ;
  assign n1259 = n1258 ^ n1257 ;
  assign n1260 = n160 & n1259 ;
  assign n1265 = n1264 ^ n1260 ;
  assign n1266 = ~n1256 & ~n1265 ;
  assign n1267 = n185 & ~n1266 ;
  assign n1233 = ~x129 & n449 ;
  assign n1232 = x129 & n343 ;
  assign n1234 = n1233 ^ n1232 ;
  assign n1235 = n148 & n1234 ;
  assign n1229 = ~x129 & n339 ;
  assign n1228 = x129 & n333 ;
  assign n1230 = n1229 ^ n1228 ;
  assign n1231 = n137 & n1230 ;
  assign n1236 = n1235 ^ n1231 ;
  assign n1242 = ~x129 & n350 ;
  assign n1241 = x129 & n364 ;
  assign n1243 = n1242 ^ n1241 ;
  assign n1244 = n171 & n1243 ;
  assign n1238 = ~x129 & n329 ;
  assign n1237 = x129 & n354 ;
  assign n1239 = n1238 ^ n1237 ;
  assign n1240 = n160 & n1239 ;
  assign n1245 = n1244 ^ n1240 ;
  assign n1246 = ~n1236 & ~n1245 ;
  assign n1247 = n136 & ~n1246 ;
  assign n1268 = n1267 ^ n1247 ;
  assign n1294 = ~x129 & n219 ;
  assign n1293 = x129 & n476 ;
  assign n1295 = n1294 ^ n1293 ;
  assign n1296 = n148 & n1295 ;
  assign n1290 = ~x129 & n472 ;
  assign n1289 = x129 & n466 ;
  assign n1291 = n1290 ^ n1289 ;
  assign n1292 = n137 & n1291 ;
  assign n1297 = n1296 ^ n1292 ;
  assign n1303 = ~x129 & n483 ;
  assign n1302 = x129 & n497 ;
  assign n1304 = n1303 ^ n1302 ;
  assign n1305 = n171 & n1304 ;
  assign n1299 = ~x129 & n462 ;
  assign n1298 = x129 & n487 ;
  assign n1300 = n1299 ^ n1298 ;
  assign n1301 = n160 & n1300 ;
  assign n1306 = n1305 ^ n1301 ;
  assign n1307 = ~n1297 & ~n1306 ;
  assign n1308 = n279 & ~n1307 ;
  assign n1274 = ~x129 & n493 ;
  assign n1273 = x129 & n432 ;
  assign n1275 = n1274 ^ n1273 ;
  assign n1276 = n148 & n1275 ;
  assign n1270 = ~x129 & n428 ;
  assign n1269 = x129 & n422 ;
  assign n1271 = n1270 ^ n1269 ;
  assign n1272 = n137 & n1271 ;
  assign n1277 = n1276 ^ n1272 ;
  assign n1283 = ~x129 & n439 ;
  assign n1282 = x129 & n453 ;
  assign n1284 = n1283 ^ n1282 ;
  assign n1285 = n171 & n1284 ;
  assign n1279 = ~x129 & n418 ;
  assign n1278 = x129 & n443 ;
  assign n1280 = n1279 ^ n1278 ;
  assign n1281 = n160 & n1280 ;
  assign n1286 = n1285 ^ n1281 ;
  assign n1287 = ~n1277 & ~n1286 ;
  assign n1288 = n254 & ~n1287 ;
  assign n1309 = n1308 ^ n1288 ;
  assign n1310 = ~n1268 & ~n1309 ;
  assign n1311 = ~x134 & n1310 ;
  assign n1163 = ~x129 & n404 ;
  assign n1162 = x129 & n296 ;
  assign n1164 = n1163 ^ n1162 ;
  assign n1165 = n148 & n1164 ;
  assign n1159 = ~x129 & n292 ;
  assign n1158 = x129 & n286 ;
  assign n1160 = n1159 ^ n1158 ;
  assign n1161 = n137 & n1160 ;
  assign n1166 = n1165 ^ n1161 ;
  assign n1172 = ~x129 & n303 ;
  assign n1171 = x129 & n317 ;
  assign n1173 = n1172 ^ n1171 ;
  assign n1174 = n171 & n1173 ;
  assign n1168 = ~x129 & n282 ;
  assign n1167 = x129 & n307 ;
  assign n1169 = n1168 ^ n1167 ;
  assign n1170 = n160 & n1169 ;
  assign n1175 = n1174 ^ n1170 ;
  assign n1176 = ~n1166 & ~n1175 ;
  assign n1177 = n279 & ~n1176 ;
  assign n1143 = ~x129 & n174 ;
  assign n1142 = x129 & n202 ;
  assign n1144 = n1143 ^ n1142 ;
  assign n1145 = n148 & n1144 ;
  assign n1139 = ~x129 & n198 ;
  assign n1138 = x129 & n192 ;
  assign n1140 = n1139 ^ n1138 ;
  assign n1141 = n137 & n1140 ;
  assign n1146 = n1145 ^ n1141 ;
  assign n1152 = ~x129 & n209 ;
  assign n1151 = x129 & n223 ;
  assign n1153 = n1152 ^ n1151 ;
  assign n1154 = n171 & n1153 ;
  assign n1148 = ~x129 & n188 ;
  assign n1147 = x129 & n213 ;
  assign n1149 = n1148 ^ n1147 ;
  assign n1150 = n160 & n1149 ;
  assign n1155 = n1154 ^ n1150 ;
  assign n1156 = ~n1146 & ~n1155 ;
  assign n1157 = n185 & ~n1156 ;
  assign n1178 = n1177 ^ n1157 ;
  assign n1204 = ~x129 & n313 ;
  assign n1203 = x129 & n271 ;
  assign n1205 = n1204 ^ n1203 ;
  assign n1206 = n148 & n1205 ;
  assign n1200 = ~x129 & n267 ;
  assign n1199 = x129 & n261 ;
  assign n1201 = n1200 ^ n1199 ;
  assign n1202 = n137 & n1201 ;
  assign n1207 = n1206 ^ n1202 ;
  assign n1217 = ~x38 & ~x128 ;
  assign n1216 = ~x37 & x128 ;
  assign n1218 = n1217 ^ n1216 ;
  assign n1219 = ~x129 & n1218 ;
  assign n1215 = x129 & ~n249 ;
  assign n1220 = n1219 ^ n1215 ;
  assign n1221 = n171 & ~n1220 ;
  assign n1212 = ~x129 & ~n257 ;
  assign n1209 = ~x40 & ~x128 ;
  assign n1208 = ~x39 & x128 ;
  assign n1210 = n1209 ^ n1208 ;
  assign n1211 = x129 & n1210 ;
  assign n1213 = n1212 ^ n1211 ;
  assign n1214 = n160 & ~n1213 ;
  assign n1222 = n1221 ^ n1214 ;
  assign n1223 = ~n1207 & ~n1222 ;
  assign n1224 = n254 & ~n1223 ;
  assign n1184 = ~x129 & n245 ;
  assign n1183 = x129 & n155 ;
  assign n1185 = n1184 ^ n1183 ;
  assign n1186 = n148 & n1185 ;
  assign n1180 = ~x129 & n151 ;
  assign n1179 = x129 & n144 ;
  assign n1181 = n1180 ^ n1179 ;
  assign n1182 = n137 & n1181 ;
  assign n1187 = n1186 ^ n1182 ;
  assign n1193 = ~x129 & n163 ;
  assign n1192 = x129 & n178 ;
  assign n1194 = n1193 ^ n1192 ;
  assign n1195 = n171 & n1194 ;
  assign n1189 = ~x129 & n140 ;
  assign n1188 = x129 & n167 ;
  assign n1190 = n1189 ^ n1188 ;
  assign n1191 = n160 & n1190 ;
  assign n1196 = n1195 ^ n1191 ;
  assign n1197 = ~n1187 & ~n1196 ;
  assign n1198 = n136 & ~n1197 ;
  assign n1225 = n1224 ^ n1198 ;
  assign n1226 = ~n1178 & ~n1225 ;
  assign n1227 = x134 & n1226 ;
  assign n1312 = n1311 ^ n1227 ;
  assign n1536 = n1108 ^ n1107 ;
  assign n1537 = n1536 ^ n994 ;
  assign n1538 = n1115 ^ n1113 ;
  assign n1539 = n1538 ^ n1002 ;
  assign n1540 = n1537 & ~n1539 ;
  assign n1541 = n1540 ^ n1539 ;
  assign n1542 = n148 & ~n1541 ;
  assign n1543 = n1542 ^ n148 ;
  assign n1528 = n992 ^ n991 ;
  assign n1529 = n1528 ^ n976 ;
  assign n1530 = n999 ^ n997 ;
  assign n1531 = n1530 ^ n984 ;
  assign n1532 = n1529 & ~n1531 ;
  assign n1533 = n1532 ^ n1531 ;
  assign n1534 = n137 & ~n1533 ;
  assign n1535 = n1534 ^ n137 ;
  assign n1544 = n1543 ^ n1535 ;
  assign n1553 = n1011 ^ n1010 ;
  assign n1554 = n1553 ^ n1031 ;
  assign n1555 = n1018 ^ n1016 ;
  assign n1556 = n1555 ^ n1039 ;
  assign n1557 = n1554 & ~n1556 ;
  assign n1558 = n1557 ^ n1556 ;
  assign n1559 = n171 & ~n1558 ;
  assign n1560 = n1559 ^ n171 ;
  assign n1545 = n974 ^ n973 ;
  assign n1546 = n1545 ^ n1013 ;
  assign n1547 = n981 ^ n979 ;
  assign n1548 = n1547 ^ n1021 ;
  assign n1549 = n1546 & ~n1548 ;
  assign n1550 = n1549 ^ n1548 ;
  assign n1551 = n160 & ~n1550 ;
  assign n1552 = n1551 ^ n160 ;
  assign n1561 = n1560 ^ n1552 ;
  assign n1562 = n1544 & n1561 ;
  assign n1563 = n1562 ^ n1544 ;
  assign n1564 = n1563 ^ n1561 ;
  assign n1565 = n254 & ~n1564 ;
  assign n1566 = n1565 ^ n254 ;
  assign n1497 = n1029 ^ n1028 ;
  assign n1498 = n1497 ^ n835 ;
  assign n1499 = n1036 ^ n1034 ;
  assign n1500 = n1499 ^ n843 ;
  assign n1501 = n1498 & ~n1500 ;
  assign n1502 = n1501 ^ n1500 ;
  assign n1503 = n148 & ~n1502 ;
  assign n1504 = n1503 ^ n148 ;
  assign n1489 = n833 ^ n832 ;
  assign n1490 = n1489 ^ n817 ;
  assign n1491 = n840 ^ n838 ;
  assign n1492 = n1491 ^ n825 ;
  assign n1493 = n1490 & ~n1492 ;
  assign n1494 = n1493 ^ n1492 ;
  assign n1495 = n137 & ~n1494 ;
  assign n1496 = n1495 ^ n137 ;
  assign n1505 = n1504 ^ n1496 ;
  assign n1514 = n852 ^ n851 ;
  assign n1515 = n1514 ^ n872 ;
  assign n1516 = n859 ^ n857 ;
  assign n1517 = n1516 ^ n880 ;
  assign n1518 = n1515 & ~n1517 ;
  assign n1519 = n1518 ^ n1517 ;
  assign n1520 = n171 & ~n1519 ;
  assign n1521 = n1520 ^ n171 ;
  assign n1506 = n815 ^ n814 ;
  assign n1507 = n1506 ^ n854 ;
  assign n1508 = n822 ^ n820 ;
  assign n1509 = n1508 ^ n862 ;
  assign n1510 = n1507 & ~n1509 ;
  assign n1511 = n1510 ^ n1509 ;
  assign n1512 = n160 & ~n1511 ;
  assign n1513 = n1512 ^ n160 ;
  assign n1522 = n1521 ^ n1513 ;
  assign n1523 = n1505 & n1522 ;
  assign n1524 = n1523 ^ n1505 ;
  assign n1525 = n1524 ^ n1522 ;
  assign n1526 = n136 & ~n1525 ;
  assign n1527 = n1526 ^ n136 ;
  assign n1567 = n1566 ^ n1527 ;
  assign n1615 = n564 ^ n563 ;
  assign n1616 = n1615 ^ n1073 ;
  assign n1617 = n571 ^ n569 ;
  assign n1618 = n1617 ^ n1081 ;
  assign n1619 = n1616 & ~n1618 ;
  assign n1620 = n1619 ^ n1618 ;
  assign n1621 = n148 & ~n1620 ;
  assign n1622 = n1621 ^ n148 ;
  assign n1607 = n1071 ^ n1070 ;
  assign n1608 = n1607 ^ n1055 ;
  assign n1609 = n1078 ^ n1076 ;
  assign n1610 = n1609 ^ n1063 ;
  assign n1611 = n1608 & ~n1610 ;
  assign n1612 = n1611 ^ n1610 ;
  assign n1613 = n137 & ~n1612 ;
  assign n1614 = n1613 ^ n137 ;
  assign n1623 = n1622 ^ n1614 ;
  assign n1632 = n1090 ^ n1089 ;
  assign n1633 = n1632 ^ n1110 ;
  assign n1634 = n1097 ^ n1095 ;
  assign n1635 = n1634 ^ n1118 ;
  assign n1636 = n1633 & ~n1635 ;
  assign n1637 = n1636 ^ n1635 ;
  assign n1638 = n171 & ~n1637 ;
  assign n1639 = n1638 ^ n171 ;
  assign n1624 = n1053 ^ n1052 ;
  assign n1625 = n1624 ^ n1092 ;
  assign n1626 = n1060 ^ n1058 ;
  assign n1627 = n1626 ^ n1100 ;
  assign n1628 = n1625 & ~n1627 ;
  assign n1629 = n1628 ^ n1627 ;
  assign n1630 = n160 & ~n1629 ;
  assign n1631 = n1630 ^ n160 ;
  assign n1640 = n1639 ^ n1631 ;
  assign n1641 = n1623 & n1640 ;
  assign n1642 = n1641 ^ n1623 ;
  assign n1643 = n1642 ^ n1640 ;
  assign n1644 = n279 & ~n1643 ;
  assign n1645 = n1644 ^ n279 ;
  assign n1576 = n870 ^ n869 ;
  assign n1577 = n1576 ^ n914 ;
  assign n1578 = n877 ^ n875 ;
  assign n1579 = n1578 ^ n922 ;
  assign n1580 = n1577 & ~n1579 ;
  assign n1581 = n1580 ^ n1579 ;
  assign n1582 = n148 & ~n1581 ;
  assign n1583 = n1582 ^ n148 ;
  assign n1568 = n912 ^ n911 ;
  assign n1569 = n1568 ^ n896 ;
  assign n1570 = n919 ^ n917 ;
  assign n1571 = n1570 ^ n904 ;
  assign n1572 = n1569 & ~n1571 ;
  assign n1573 = n1572 ^ n1571 ;
  assign n1574 = n137 & ~n1573 ;
  assign n1575 = n1574 ^ n137 ;
  assign n1584 = n1583 ^ n1575 ;
  assign n1593 = n931 ^ n930 ;
  assign n1594 = n1593 ^ n951 ;
  assign n1595 = n938 ^ n936 ;
  assign n1596 = n1595 ^ n959 ;
  assign n1597 = n1594 & ~n1596 ;
  assign n1598 = n1597 ^ n1596 ;
  assign n1599 = n171 & ~n1598 ;
  assign n1600 = n1599 ^ n171 ;
  assign n1585 = n894 ^ n893 ;
  assign n1586 = n1585 ^ n933 ;
  assign n1587 = n901 ^ n899 ;
  assign n1588 = n1587 ^ n941 ;
  assign n1589 = n1586 & ~n1588 ;
  assign n1590 = n1589 ^ n1588 ;
  assign n1591 = n160 & ~n1590 ;
  assign n1592 = n1591 ^ n160 ;
  assign n1601 = n1600 ^ n1592 ;
  assign n1602 = n1584 & n1601 ;
  assign n1603 = n1602 ^ n1584 ;
  assign n1604 = n1603 ^ n1601 ;
  assign n1605 = n185 & ~n1604 ;
  assign n1606 = n1605 ^ n185 ;
  assign n1646 = n1645 ^ n1606 ;
  assign n1647 = n1567 & n1646 ;
  assign n1648 = n1647 ^ n1567 ;
  assign n1649 = n1648 ^ n1646 ;
  assign n1650 = x134 & ~n1649 ;
  assign n1651 = n1650 ^ n1649 ;
  assign n1374 = n949 ^ n948 ;
  assign n1375 = n1374 ^ n608 ;
  assign n1376 = n956 ^ n954 ;
  assign n1377 = n1376 ^ n616 ;
  assign n1378 = n1375 & ~n1377 ;
  assign n1379 = n1378 ^ n1377 ;
  assign n1380 = n148 & ~n1379 ;
  assign n1381 = n1380 ^ n148 ;
  assign n1366 = n606 ^ n605 ;
  assign n1367 = n1366 ^ n590 ;
  assign n1368 = n613 ^ n611 ;
  assign n1369 = n1368 ^ n598 ;
  assign n1370 = n1367 & ~n1369 ;
  assign n1371 = n1370 ^ n1369 ;
  assign n1372 = n137 & ~n1371 ;
  assign n1373 = n1372 ^ n137 ;
  assign n1382 = n1381 ^ n1373 ;
  assign n1391 = n625 ^ n624 ;
  assign n1392 = n1391 ^ n645 ;
  assign n1393 = n632 ^ n630 ;
  assign n1394 = n1393 ^ n653 ;
  assign n1395 = n1392 & ~n1394 ;
  assign n1396 = n1395 ^ n1394 ;
  assign n1397 = n171 & ~n1396 ;
  assign n1398 = n1397 ^ n171 ;
  assign n1383 = n588 ^ n587 ;
  assign n1384 = n1383 ^ n627 ;
  assign n1385 = n595 ^ n593 ;
  assign n1386 = n1385 ^ n635 ;
  assign n1387 = n1384 & ~n1386 ;
  assign n1388 = n1387 ^ n1386 ;
  assign n1389 = n160 & ~n1388 ;
  assign n1390 = n1389 ^ n160 ;
  assign n1399 = n1398 ^ n1390 ;
  assign n1400 = n1382 & n1399 ;
  assign n1401 = n1400 ^ n1382 ;
  assign n1402 = n1401 ^ n1399 ;
  assign n1403 = n279 & ~n1402 ;
  assign n1404 = n1403 ^ n279 ;
  assign n1320 = n643 ^ n642 ;
  assign n1321 = n1320 ^ n759 ;
  assign n1322 = n650 ^ n648 ;
  assign n1323 = n1322 ^ n767 ;
  assign n1324 = n1321 & ~n1323 ;
  assign n1325 = n1324 ^ n1323 ;
  assign n1326 = n148 & ~n1325 ;
  assign n1327 = n1326 ^ n148 ;
  assign n1315 = ~x47 & ~x128 ;
  assign n1314 = ~x46 & x128 ;
  assign n1316 = n1315 ^ n1314 ;
  assign n1317 = ~x129 & n1316 ;
  assign n1313 = x129 & ~n752 ;
  assign n1318 = n1317 ^ n1313 ;
  assign n1319 = n137 & ~n1318 ;
  assign n1328 = n1327 ^ n1319 ;
  assign n1347 = n233 ^ x39 ;
  assign n1348 = x129 & n1347 ;
  assign n1349 = n1348 ^ n1347 ;
  assign n1350 = n1349 ^ n788 ;
  assign n1351 = x38 & x128 ;
  assign n1352 = x129 & n1351 ;
  assign n1353 = n1352 ^ x129 ;
  assign n1354 = n1353 ^ n1351 ;
  assign n1355 = n1354 ^ n796 ;
  assign n1356 = n1350 & ~n1355 ;
  assign n1357 = n1356 ^ n1355 ;
  assign n1358 = n171 & ~n1357 ;
  assign n1359 = n1358 ^ n171 ;
  assign n1331 = n259 ^ x43 ;
  assign n1332 = x129 & n1331 ;
  assign n1333 = n1332 ^ n1331 ;
  assign n1329 = x40 & x128 ;
  assign n1330 = x129 & n1329 ;
  assign n1334 = n1333 ^ n1330 ;
  assign n1338 = x42 & x128 ;
  assign n1339 = x129 & n1338 ;
  assign n1340 = n1339 ^ x129 ;
  assign n1341 = n1340 ^ n1338 ;
  assign n1335 = n255 ^ x41 ;
  assign n1336 = x129 & n1335 ;
  assign n1337 = n1336 ^ x129 ;
  assign n1342 = n1341 ^ n1337 ;
  assign n1343 = n1334 & ~n1342 ;
  assign n1344 = n1343 ^ n1342 ;
  assign n1345 = n160 & ~n1344 ;
  assign n1346 = n1345 ^ n160 ;
  assign n1360 = n1359 ^ n1346 ;
  assign n1361 = n1328 & n1360 ;
  assign n1362 = n1361 ^ n1328 ;
  assign n1363 = n1362 ^ n1360 ;
  assign n1364 = n254 & ~n1363 ;
  assign n1365 = n1364 ^ n254 ;
  assign n1405 = n1404 ^ n1365 ;
  assign n1453 = n723 ^ n722 ;
  assign n1454 = n1453 ^ n529 ;
  assign n1455 = n730 ^ n728 ;
  assign n1456 = n1455 ^ n537 ;
  assign n1457 = n1454 & ~n1456 ;
  assign n1458 = n1457 ^ n1456 ;
  assign n1459 = n148 & ~n1458 ;
  assign n1460 = n1459 ^ n148 ;
  assign n1445 = n527 ^ n526 ;
  assign n1446 = n1445 ^ n511 ;
  assign n1447 = n534 ^ n532 ;
  assign n1448 = n1447 ^ n519 ;
  assign n1449 = n1446 & ~n1448 ;
  assign n1450 = n1449 ^ n1448 ;
  assign n1451 = n137 & ~n1450 ;
  assign n1452 = n1451 ^ n137 ;
  assign n1461 = n1460 ^ n1452 ;
  assign n1470 = n546 ^ n545 ;
  assign n1471 = n1470 ^ n566 ;
  assign n1472 = n553 ^ n551 ;
  assign n1473 = n1472 ^ n574 ;
  assign n1474 = n1471 & ~n1473 ;
  assign n1475 = n1474 ^ n1473 ;
  assign n1476 = n171 & ~n1475 ;
  assign n1477 = n1476 ^ n171 ;
  assign n1462 = n509 ^ n508 ;
  assign n1463 = n1462 ^ n548 ;
  assign n1464 = n516 ^ n514 ;
  assign n1465 = n1464 ^ n556 ;
  assign n1466 = n1463 & ~n1465 ;
  assign n1467 = n1466 ^ n1465 ;
  assign n1468 = n160 & ~n1467 ;
  assign n1469 = n1468 ^ n160 ;
  assign n1478 = n1477 ^ n1469 ;
  assign n1479 = n1461 & n1478 ;
  assign n1480 = n1479 ^ n1461 ;
  assign n1481 = n1480 ^ n1478 ;
  assign n1482 = n185 & ~n1481 ;
  assign n1483 = n1482 ^ n185 ;
  assign n1414 = n786 ^ n785 ;
  assign n1415 = n1414 ^ n688 ;
  assign n1416 = n793 ^ n791 ;
  assign n1417 = n1416 ^ n696 ;
  assign n1418 = n1415 & ~n1417 ;
  assign n1419 = n1418 ^ n1417 ;
  assign n1420 = n148 & ~n1419 ;
  assign n1421 = n1420 ^ n148 ;
  assign n1406 = n686 ^ n685 ;
  assign n1407 = n1406 ^ n670 ;
  assign n1408 = n693 ^ n691 ;
  assign n1409 = n1408 ^ n678 ;
  assign n1410 = n1407 & ~n1409 ;
  assign n1411 = n1410 ^ n1409 ;
  assign n1412 = n137 & ~n1411 ;
  assign n1413 = n1412 ^ n137 ;
  assign n1422 = n1421 ^ n1413 ;
  assign n1431 = n705 ^ n704 ;
  assign n1432 = n1431 ^ n725 ;
  assign n1433 = n712 ^ n710 ;
  assign n1434 = n1433 ^ n733 ;
  assign n1435 = n1432 & ~n1434 ;
  assign n1436 = n1435 ^ n1434 ;
  assign n1437 = n171 & ~n1436 ;
  assign n1438 = n1437 ^ n171 ;
  assign n1423 = n668 ^ n667 ;
  assign n1424 = n1423 ^ n707 ;
  assign n1425 = n675 ^ n673 ;
  assign n1426 = n1425 ^ n715 ;
  assign n1427 = n1424 & ~n1426 ;
  assign n1428 = n1427 ^ n1426 ;
  assign n1429 = n160 & ~n1428 ;
  assign n1430 = n1429 ^ n160 ;
  assign n1439 = n1438 ^ n1430 ;
  assign n1440 = n1422 & n1439 ;
  assign n1441 = n1440 ^ n1422 ;
  assign n1442 = n1441 ^ n1439 ;
  assign n1443 = n136 & ~n1442 ;
  assign n1444 = n1443 ^ n136 ;
  assign n1484 = n1483 ^ n1444 ;
  assign n1485 = n1405 & n1484 ;
  assign n1486 = n1485 ^ n1405 ;
  assign n1487 = n1486 ^ n1484 ;
  assign n1488 = x134 & ~n1487 ;
  assign n1652 = n1651 ^ n1488 ;
  assign n1699 = n148 & n366 ;
  assign n1698 = n137 & n389 ;
  assign n1700 = n1699 ^ n1698 ;
  assign n1702 = n171 & n400 ;
  assign n1701 = n160 & n379 ;
  assign n1703 = n1702 ^ n1701 ;
  assign n1704 = ~n1700 & ~n1703 ;
  assign n1705 = n185 & ~n1704 ;
  assign n1691 = n148 & n455 ;
  assign n1690 = n137 & n345 ;
  assign n1692 = n1691 ^ n1690 ;
  assign n1694 = n171 & n356 ;
  assign n1693 = n160 & n335 ;
  assign n1695 = n1694 ^ n1693 ;
  assign n1696 = ~n1692 & ~n1695 ;
  assign n1697 = n136 & ~n1696 ;
  assign n1706 = n1705 ^ n1697 ;
  assign n1716 = n148 & n225 ;
  assign n1715 = n137 & n478 ;
  assign n1717 = n1716 ^ n1715 ;
  assign n1719 = n171 & n489 ;
  assign n1718 = n160 & n468 ;
  assign n1720 = n1719 ^ n1718 ;
  assign n1721 = ~n1717 & ~n1720 ;
  assign n1722 = n279 & ~n1721 ;
  assign n1708 = n148 & n499 ;
  assign n1707 = n137 & n434 ;
  assign n1709 = n1708 ^ n1707 ;
  assign n1711 = n171 & n445 ;
  assign n1710 = n160 & n424 ;
  assign n1712 = n1711 ^ n1710 ;
  assign n1713 = ~n1709 & ~n1712 ;
  assign n1714 = n254 & ~n1713 ;
  assign n1723 = n1722 ^ n1714 ;
  assign n1724 = ~n1706 & ~n1723 ;
  assign n1725 = ~x134 & n1724 ;
  assign n1662 = n171 & ~n241 ;
  assign n1661 = n160 & n263 ;
  assign n1663 = n1662 ^ n1661 ;
  assign n1665 = n148 & n319 ;
  assign n1664 = n137 & n273 ;
  assign n1666 = n1665 ^ n1664 ;
  assign n1667 = n254 & ~n1666 ;
  assign n1668 = ~n1663 & n1667 ;
  assign n1654 = n148 & n410 ;
  assign n1653 = n137 & n298 ;
  assign n1655 = n1654 ^ n1653 ;
  assign n1657 = n171 & n309 ;
  assign n1656 = n160 & n288 ;
  assign n1658 = n1657 ^ n1656 ;
  assign n1659 = ~n1655 & ~n1658 ;
  assign n1660 = n279 & n1659 ;
  assign n1669 = n1668 ^ n1660 ;
  assign n1670 = n1669 ^ x133 ;
  assign n1680 = n148 & n251 ;
  assign n1679 = n137 & n157 ;
  assign n1681 = n1680 ^ n1679 ;
  assign n1683 = n169 & n171 ;
  assign n1682 = n146 & n160 ;
  assign n1684 = n1683 ^ n1682 ;
  assign n1685 = ~n1681 & ~n1684 ;
  assign n1686 = n136 & ~n1685 ;
  assign n1672 = n148 & n180 ;
  assign n1671 = n137 & n204 ;
  assign n1673 = n1672 ^ n1671 ;
  assign n1675 = n171 & n215 ;
  assign n1674 = n160 & n194 ;
  assign n1676 = n1675 ^ n1674 ;
  assign n1677 = ~n1673 & ~n1676 ;
  assign n1678 = n185 & ~n1677 ;
  assign n1687 = n1686 ^ n1678 ;
  assign n1688 = n1670 & ~n1687 ;
  assign n1689 = x134 & n1688 ;
  assign n1726 = n1725 ^ n1689 ;
  assign n1811 = n148 & ~n884 ;
  assign n1812 = n1811 ^ n148 ;
  assign n1809 = n137 & ~n926 ;
  assign n1810 = n1809 ^ n137 ;
  assign n1813 = n1812 ^ n1810 ;
  assign n1816 = n171 & ~n945 ;
  assign n1817 = n1816 ^ n171 ;
  assign n1814 = n160 & ~n908 ;
  assign n1815 = n1814 ^ n160 ;
  assign n1818 = n1817 ^ n1815 ;
  assign n1819 = n1813 & n1818 ;
  assign n1820 = n1819 ^ n1813 ;
  assign n1821 = n1820 ^ n1818 ;
  assign n1822 = n185 & ~n1821 ;
  assign n1823 = n1822 ^ n185 ;
  assign n1796 = n148 & ~n1043 ;
  assign n1797 = n1796 ^ n148 ;
  assign n1794 = n137 & ~n847 ;
  assign n1795 = n1794 ^ n137 ;
  assign n1798 = n1797 ^ n1795 ;
  assign n1801 = n171 & ~n866 ;
  assign n1802 = n1801 ^ n171 ;
  assign n1799 = n160 & ~n829 ;
  assign n1800 = n1799 ^ n160 ;
  assign n1803 = n1802 ^ n1800 ;
  assign n1804 = n1798 & n1803 ;
  assign n1805 = n1804 ^ n1798 ;
  assign n1806 = n1805 ^ n1803 ;
  assign n1807 = n136 & ~n1806 ;
  assign n1808 = n1807 ^ n136 ;
  assign n1824 = n1823 ^ n1808 ;
  assign n1842 = n148 & ~n578 ;
  assign n1843 = n1842 ^ n148 ;
  assign n1840 = n137 & ~n1085 ;
  assign n1841 = n1840 ^ n137 ;
  assign n1844 = n1843 ^ n1841 ;
  assign n1847 = n171 & ~n1104 ;
  assign n1848 = n1847 ^ n171 ;
  assign n1845 = n160 & ~n1067 ;
  assign n1846 = n1845 ^ n160 ;
  assign n1849 = n1848 ^ n1846 ;
  assign n1850 = n1844 & n1849 ;
  assign n1851 = n1850 ^ n1844 ;
  assign n1852 = n1851 ^ n1849 ;
  assign n1853 = n279 & ~n1852 ;
  assign n1854 = n1853 ^ n279 ;
  assign n1827 = n148 & ~n1122 ;
  assign n1828 = n1827 ^ n148 ;
  assign n1825 = n137 & ~n1006 ;
  assign n1826 = n1825 ^ n137 ;
  assign n1829 = n1828 ^ n1826 ;
  assign n1832 = n171 & ~n1025 ;
  assign n1833 = n1832 ^ n171 ;
  assign n1830 = n160 & ~n988 ;
  assign n1831 = n1830 ^ n160 ;
  assign n1834 = n1833 ^ n1831 ;
  assign n1835 = n1829 & n1834 ;
  assign n1836 = n1835 ^ n1829 ;
  assign n1837 = n1836 ^ n1834 ;
  assign n1838 = n254 & ~n1837 ;
  assign n1839 = n1838 ^ n254 ;
  assign n1855 = n1854 ^ n1839 ;
  assign n1856 = n1824 & n1855 ;
  assign n1857 = n1856 ^ n1824 ;
  assign n1858 = n1857 ^ n1855 ;
  assign n1859 = x134 & ~n1858 ;
  assign n1860 = n1859 ^ n1858 ;
  assign n1747 = n148 & ~n657 ;
  assign n1748 = n1747 ^ n148 ;
  assign n1745 = n137 & ~n771 ;
  assign n1746 = n1745 ^ n137 ;
  assign n1749 = n1748 ^ n1746 ;
  assign n1743 = n171 & ~n783 ;
  assign n1742 = n160 & ~n754 ;
  assign n1744 = n1743 ^ n1742 ;
  assign n1750 = n1749 ^ n1744 ;
  assign n1751 = n1744 ^ n254 ;
  assign n1752 = ~n254 & n1751 ;
  assign n1753 = n1752 ^ n254 ;
  assign n1754 = n1753 ^ n1749 ;
  assign n1755 = n1750 & n1754 ;
  assign n1756 = n1755 ^ n1752 ;
  assign n1757 = n1756 ^ n1749 ;
  assign n1729 = n148 & ~n963 ;
  assign n1730 = n1729 ^ n148 ;
  assign n1727 = n137 & ~n620 ;
  assign n1728 = n1727 ^ n137 ;
  assign n1731 = n1730 ^ n1728 ;
  assign n1734 = n171 & ~n639 ;
  assign n1735 = n1734 ^ n171 ;
  assign n1732 = n160 & ~n602 ;
  assign n1733 = n1732 ^ n160 ;
  assign n1736 = n1735 ^ n1733 ;
  assign n1737 = n1731 & n1736 ;
  assign n1738 = n1737 ^ n1731 ;
  assign n1739 = n1738 ^ n1736 ;
  assign n1740 = n279 & ~n1739 ;
  assign n1741 = n1740 ^ n279 ;
  assign n1758 = n1757 ^ n1741 ;
  assign n1776 = n148 & ~n800 ;
  assign n1777 = n1776 ^ n148 ;
  assign n1774 = n137 & ~n700 ;
  assign n1775 = n1774 ^ n137 ;
  assign n1778 = n1777 ^ n1775 ;
  assign n1781 = n171 & ~n719 ;
  assign n1782 = n1781 ^ n171 ;
  assign n1779 = n160 & ~n682 ;
  assign n1780 = n1779 ^ n160 ;
  assign n1783 = n1782 ^ n1780 ;
  assign n1784 = n1778 & n1783 ;
  assign n1785 = n1784 ^ n1778 ;
  assign n1786 = n1785 ^ n1783 ;
  assign n1787 = n136 & ~n1786 ;
  assign n1788 = n1787 ^ n136 ;
  assign n1761 = n148 & ~n737 ;
  assign n1762 = n1761 ^ n148 ;
  assign n1759 = n137 & ~n541 ;
  assign n1760 = n1759 ^ n137 ;
  assign n1763 = n1762 ^ n1760 ;
  assign n1766 = n171 & ~n560 ;
  assign n1767 = n1766 ^ n171 ;
  assign n1764 = n160 & ~n523 ;
  assign n1765 = n1764 ^ n160 ;
  assign n1768 = n1767 ^ n1765 ;
  assign n1769 = n1763 & n1768 ;
  assign n1770 = n1769 ^ n1763 ;
  assign n1771 = n1770 ^ n1768 ;
  assign n1772 = n185 & ~n1771 ;
  assign n1773 = n1772 ^ n185 ;
  assign n1789 = n1788 ^ n1773 ;
  assign n1790 = n1758 & n1789 ;
  assign n1791 = n1790 ^ n1758 ;
  assign n1792 = n1791 ^ n1789 ;
  assign n1793 = x134 & ~n1792 ;
  assign n1861 = n1860 ^ n1793 ;
  assign n1907 = n148 & n1243 ;
  assign n1906 = n137 & n1254 ;
  assign n1908 = n1907 ^ n1906 ;
  assign n1910 = n171 & n1259 ;
  assign n1909 = n160 & n1250 ;
  assign n1911 = n1910 ^ n1909 ;
  assign n1912 = ~n1908 & ~n1911 ;
  assign n1913 = n185 & ~n1912 ;
  assign n1899 = n148 & n1284 ;
  assign n1898 = n137 & n1234 ;
  assign n1900 = n1899 ^ n1898 ;
  assign n1902 = n171 & n1239 ;
  assign n1901 = n160 & n1230 ;
  assign n1903 = n1902 ^ n1901 ;
  assign n1904 = ~n1900 & ~n1903 ;
  assign n1905 = n136 & ~n1904 ;
  assign n1914 = n1913 ^ n1905 ;
  assign n1924 = n148 & n1153 ;
  assign n1923 = n137 & n1295 ;
  assign n1925 = n1924 ^ n1923 ;
  assign n1927 = n171 & n1300 ;
  assign n1926 = n160 & n1291 ;
  assign n1928 = n1927 ^ n1926 ;
  assign n1929 = ~n1925 & ~n1928 ;
  assign n1930 = n279 & ~n1929 ;
  assign n1916 = n148 & n1304 ;
  assign n1915 = n137 & n1275 ;
  assign n1917 = n1916 ^ n1915 ;
  assign n1919 = n171 & n1280 ;
  assign n1918 = n160 & n1271 ;
  assign n1920 = n1919 ^ n1918 ;
  assign n1921 = ~n1917 & ~n1920 ;
  assign n1922 = n254 & ~n1921 ;
  assign n1931 = n1930 ^ n1922 ;
  assign n1932 = ~n1914 & ~n1931 ;
  assign n1933 = ~x134 & n1932 ;
  assign n1871 = n148 & n1173 ;
  assign n1870 = n137 & n1205 ;
  assign n1872 = n1871 ^ n1870 ;
  assign n1874 = n171 & ~n1213 ;
  assign n1873 = n160 & n1201 ;
  assign n1875 = n1874 ^ n1873 ;
  assign n1876 = ~n1872 & ~n1875 ;
  assign n1877 = n254 & ~n1876 ;
  assign n1863 = n148 & n1263 ;
  assign n1862 = n137 & n1164 ;
  assign n1864 = n1863 ^ n1862 ;
  assign n1866 = n171 & n1169 ;
  assign n1865 = n160 & n1160 ;
  assign n1867 = n1866 ^ n1865 ;
  assign n1868 = ~n1864 & ~n1867 ;
  assign n1869 = n279 & ~n1868 ;
  assign n1878 = n1877 ^ n1869 ;
  assign n1888 = n148 & ~n1220 ;
  assign n1887 = n137 & n1185 ;
  assign n1889 = n1888 ^ n1887 ;
  assign n1891 = n171 & n1190 ;
  assign n1890 = n160 & n1181 ;
  assign n1892 = n1891 ^ n1890 ;
  assign n1893 = ~n1889 & ~n1892 ;
  assign n1894 = n136 & ~n1893 ;
  assign n1880 = n148 & n1194 ;
  assign n1879 = n137 & n1144 ;
  assign n1881 = n1880 ^ n1879 ;
  assign n1883 = n171 & n1149 ;
  assign n1882 = n160 & n1140 ;
  assign n1884 = n1883 ^ n1882 ;
  assign n1885 = ~n1881 & ~n1884 ;
  assign n1886 = n185 & ~n1885 ;
  assign n1895 = n1894 ^ n1886 ;
  assign n1896 = ~n1878 & ~n1895 ;
  assign n1897 = x134 & n1896 ;
  assign n1934 = n1933 ^ n1897 ;
  assign n2017 = n148 & ~n1519 ;
  assign n2018 = n2017 ^ n148 ;
  assign n2015 = n137 & ~n1581 ;
  assign n2016 = n2015 ^ n137 ;
  assign n2019 = n2018 ^ n2016 ;
  assign n2022 = n171 & ~n1590 ;
  assign n2023 = n2022 ^ n171 ;
  assign n2020 = n160 & ~n1573 ;
  assign n2021 = n2020 ^ n160 ;
  assign n2024 = n2023 ^ n2021 ;
  assign n2025 = n2019 & n2024 ;
  assign n2026 = n2025 ^ n2019 ;
  assign n2027 = n2026 ^ n2024 ;
  assign n2028 = n185 & ~n2027 ;
  assign n2029 = n2028 ^ n185 ;
  assign n2002 = n148 & ~n1558 ;
  assign n2003 = n2002 ^ n148 ;
  assign n2000 = n137 & ~n1502 ;
  assign n2001 = n2000 ^ n137 ;
  assign n2004 = n2003 ^ n2001 ;
  assign n2007 = n171 & ~n1511 ;
  assign n2008 = n2007 ^ n171 ;
  assign n2005 = n160 & ~n1494 ;
  assign n2006 = n2005 ^ n160 ;
  assign n2009 = n2008 ^ n2006 ;
  assign n2010 = n2004 & n2009 ;
  assign n2011 = n2010 ^ n2004 ;
  assign n2012 = n2011 ^ n2009 ;
  assign n2013 = n136 & ~n2012 ;
  assign n2014 = n2013 ^ n136 ;
  assign n2030 = n2029 ^ n2014 ;
  assign n2048 = n148 & ~n1475 ;
  assign n2049 = n2048 ^ n148 ;
  assign n2046 = n137 & ~n1620 ;
  assign n2047 = n2046 ^ n137 ;
  assign n2050 = n2049 ^ n2047 ;
  assign n2053 = n171 & ~n1629 ;
  assign n2054 = n2053 ^ n171 ;
  assign n2051 = n160 & ~n1612 ;
  assign n2052 = n2051 ^ n160 ;
  assign n2055 = n2054 ^ n2052 ;
  assign n2056 = n2050 & n2055 ;
  assign n2057 = n2056 ^ n2050 ;
  assign n2058 = n2057 ^ n2055 ;
  assign n2059 = n279 & ~n2058 ;
  assign n2060 = n2059 ^ n279 ;
  assign n2033 = n148 & ~n1637 ;
  assign n2034 = n2033 ^ n148 ;
  assign n2031 = n137 & ~n1541 ;
  assign n2032 = n2031 ^ n137 ;
  assign n2035 = n2034 ^ n2032 ;
  assign n2038 = n171 & ~n1550 ;
  assign n2039 = n2038 ^ n171 ;
  assign n2036 = n160 & ~n1533 ;
  assign n2037 = n2036 ^ n160 ;
  assign n2040 = n2039 ^ n2037 ;
  assign n2041 = n2035 & n2040 ;
  assign n2042 = n2041 ^ n2035 ;
  assign n2043 = n2042 ^ n2040 ;
  assign n2044 = n254 & ~n2043 ;
  assign n2045 = n2044 ^ n254 ;
  assign n2061 = n2060 ^ n2045 ;
  assign n2062 = n2030 & n2061 ;
  assign n2063 = n2062 ^ n2030 ;
  assign n2064 = n2063 ^ n2061 ;
  assign n2065 = x134 & ~n2064 ;
  assign n2066 = n2065 ^ n2064 ;
  assign n1951 = n137 & ~n1325 ;
  assign n1952 = n1951 ^ n137 ;
  assign n1950 = n160 & ~n1318 ;
  assign n1953 = n1952 ^ n1950 ;
  assign n1956 = n171 & ~n1344 ;
  assign n1957 = n1956 ^ n171 ;
  assign n1954 = n148 & ~n1396 ;
  assign n1955 = n1954 ^ n148 ;
  assign n1958 = n1957 ^ n1955 ;
  assign n1959 = n1953 & n1958 ;
  assign n1960 = n1959 ^ n1953 ;
  assign n1961 = n1960 ^ n1958 ;
  assign n1962 = n254 & ~n1961 ;
  assign n1963 = n1962 ^ n254 ;
  assign n1937 = n148 & ~n1598 ;
  assign n1938 = n1937 ^ n148 ;
  assign n1935 = n137 & ~n1379 ;
  assign n1936 = n1935 ^ n137 ;
  assign n1939 = n1938 ^ n1936 ;
  assign n1942 = n171 & ~n1388 ;
  assign n1943 = n1942 ^ n171 ;
  assign n1940 = n160 & ~n1371 ;
  assign n1941 = n1940 ^ n160 ;
  assign n1944 = n1943 ^ n1941 ;
  assign n1945 = n1939 & n1944 ;
  assign n1946 = n1945 ^ n1939 ;
  assign n1947 = n1946 ^ n1944 ;
  assign n1948 = n279 & ~n1947 ;
  assign n1949 = n1948 ^ n279 ;
  assign n1964 = n1963 ^ n1949 ;
  assign n1982 = n148 & ~n1357 ;
  assign n1983 = n1982 ^ n148 ;
  assign n1980 = n137 & ~n1419 ;
  assign n1981 = n1980 ^ n137 ;
  assign n1984 = n1983 ^ n1981 ;
  assign n1987 = n171 & ~n1428 ;
  assign n1988 = n1987 ^ n171 ;
  assign n1985 = n160 & ~n1411 ;
  assign n1986 = n1985 ^ n160 ;
  assign n1989 = n1988 ^ n1986 ;
  assign n1990 = n1984 & n1989 ;
  assign n1991 = n1990 ^ n1984 ;
  assign n1992 = n1991 ^ n1989 ;
  assign n1993 = n136 & ~n1992 ;
  assign n1994 = n1993 ^ n136 ;
  assign n1967 = n148 & ~n1436 ;
  assign n1968 = n1967 ^ n148 ;
  assign n1965 = n137 & ~n1458 ;
  assign n1966 = n1965 ^ n137 ;
  assign n1969 = n1968 ^ n1966 ;
  assign n1972 = n171 & ~n1467 ;
  assign n1973 = n1972 ^ n171 ;
  assign n1970 = n160 & ~n1450 ;
  assign n1971 = n1970 ^ n160 ;
  assign n1974 = n1973 ^ n1971 ;
  assign n1975 = n1969 & n1974 ;
  assign n1976 = n1975 ^ n1969 ;
  assign n1977 = n1976 ^ n1974 ;
  assign n1978 = n185 & ~n1977 ;
  assign n1979 = n1978 ^ n185 ;
  assign n1995 = n1994 ^ n1979 ;
  assign n1996 = n1964 & n1995 ;
  assign n1997 = n1996 ^ n1964 ;
  assign n1998 = n1997 ^ n1995 ;
  assign n1999 = x134 & ~n1998 ;
  assign n2067 = n2066 ^ n1999 ;
  assign n2114 = n148 & n356 ;
  assign n2113 = n137 & n366 ;
  assign n2115 = n2114 ^ n2113 ;
  assign n2117 = n171 & n379 ;
  assign n2116 = n160 & n389 ;
  assign n2118 = n2117 ^ n2116 ;
  assign n2119 = ~n2115 & ~n2118 ;
  assign n2120 = n185 & ~n2119 ;
  assign n2106 = n148 & n445 ;
  assign n2105 = n137 & n455 ;
  assign n2107 = n2106 ^ n2105 ;
  assign n2109 = n171 & n335 ;
  assign n2108 = n160 & n345 ;
  assign n2110 = n2109 ^ n2108 ;
  assign n2111 = ~n2107 & ~n2110 ;
  assign n2112 = n136 & ~n2111 ;
  assign n2121 = n2120 ^ n2112 ;
  assign n2131 = n148 & n215 ;
  assign n2130 = n137 & n225 ;
  assign n2132 = n2131 ^ n2130 ;
  assign n2134 = n171 & n468 ;
  assign n2133 = n160 & n478 ;
  assign n2135 = n2134 ^ n2133 ;
  assign n2136 = ~n2132 & ~n2135 ;
  assign n2137 = n279 & ~n2136 ;
  assign n2123 = n148 & n489 ;
  assign n2122 = n137 & n499 ;
  assign n2124 = n2123 ^ n2122 ;
  assign n2126 = n171 & n424 ;
  assign n2125 = n160 & n434 ;
  assign n2127 = n2126 ^ n2125 ;
  assign n2128 = ~n2124 & ~n2127 ;
  assign n2129 = n254 & ~n2128 ;
  assign n2138 = n2137 ^ n2129 ;
  assign n2139 = ~n2121 & ~n2138 ;
  assign n2140 = ~x134 & n2139 ;
  assign n2077 = n148 & n309 ;
  assign n2076 = n137 & n319 ;
  assign n2078 = n2077 ^ n2076 ;
  assign n2080 = n171 & n263 ;
  assign n2079 = n160 & n273 ;
  assign n2081 = n2080 ^ n2079 ;
  assign n2082 = ~n2078 & ~n2081 ;
  assign n2083 = n254 & ~n2082 ;
  assign n2069 = n148 & n400 ;
  assign n2068 = n137 & n410 ;
  assign n2070 = n2069 ^ n2068 ;
  assign n2072 = n171 & n288 ;
  assign n2071 = n160 & n298 ;
  assign n2073 = n2072 ^ n2071 ;
  assign n2074 = ~n2070 & ~n2073 ;
  assign n2075 = n279 & ~n2074 ;
  assign n2084 = n2083 ^ n2075 ;
  assign n2095 = n148 & n169 ;
  assign n2094 = n137 & n180 ;
  assign n2096 = n2095 ^ n2094 ;
  assign n2098 = n171 & n194 ;
  assign n2097 = n160 & n204 ;
  assign n2099 = n2098 ^ n2097 ;
  assign n2100 = ~n2096 & ~n2099 ;
  assign n2101 = n185 & n2100 ;
  assign n2086 = n148 & ~n241 ;
  assign n2085 = n137 & n251 ;
  assign n2087 = n2086 ^ n2085 ;
  assign n2089 = n146 & n171 ;
  assign n2088 = n157 & n160 ;
  assign n2090 = n2089 ^ n2088 ;
  assign n2091 = n136 & ~n2090 ;
  assign n2092 = ~n2087 & n2091 ;
  assign n2093 = n2092 ^ x133 ;
  assign n2102 = n2101 ^ n2093 ;
  assign n2103 = ~n2084 & ~n2102 ;
  assign n2104 = x134 & n2103 ;
  assign n2141 = n2140 ^ n2104 ;
  assign n2223 = n148 & ~n866 ;
  assign n2224 = n2223 ^ n148 ;
  assign n2221 = n137 & ~n884 ;
  assign n2222 = n2221 ^ n137 ;
  assign n2225 = n2224 ^ n2222 ;
  assign n2228 = n171 & ~n908 ;
  assign n2229 = n2228 ^ n171 ;
  assign n2226 = n160 & ~n926 ;
  assign n2227 = n2226 ^ n160 ;
  assign n2230 = n2229 ^ n2227 ;
  assign n2231 = n2225 & n2230 ;
  assign n2232 = n2231 ^ n2225 ;
  assign n2233 = n2232 ^ n2230 ;
  assign n2234 = n185 & ~n2233 ;
  assign n2235 = n2234 ^ n185 ;
  assign n2208 = n148 & ~n1025 ;
  assign n2209 = n2208 ^ n148 ;
  assign n2206 = n137 & ~n1043 ;
  assign n2207 = n2206 ^ n137 ;
  assign n2210 = n2209 ^ n2207 ;
  assign n2213 = n171 & ~n829 ;
  assign n2214 = n2213 ^ n171 ;
  assign n2211 = n160 & ~n847 ;
  assign n2212 = n2211 ^ n160 ;
  assign n2215 = n2214 ^ n2212 ;
  assign n2216 = n2210 & n2215 ;
  assign n2217 = n2216 ^ n2210 ;
  assign n2218 = n2217 ^ n2215 ;
  assign n2219 = n136 & ~n2218 ;
  assign n2220 = n2219 ^ n136 ;
  assign n2236 = n2235 ^ n2220 ;
  assign n2254 = n148 & ~n560 ;
  assign n2255 = n2254 ^ n148 ;
  assign n2252 = n137 & ~n578 ;
  assign n2253 = n2252 ^ n137 ;
  assign n2256 = n2255 ^ n2253 ;
  assign n2259 = n171 & ~n1067 ;
  assign n2260 = n2259 ^ n171 ;
  assign n2257 = n160 & ~n1085 ;
  assign n2258 = n2257 ^ n160 ;
  assign n2261 = n2260 ^ n2258 ;
  assign n2262 = n2256 & n2261 ;
  assign n2263 = n2262 ^ n2256 ;
  assign n2264 = n2263 ^ n2261 ;
  assign n2265 = n279 & ~n2264 ;
  assign n2266 = n2265 ^ n279 ;
  assign n2239 = n148 & ~n1104 ;
  assign n2240 = n2239 ^ n148 ;
  assign n2237 = n137 & ~n1122 ;
  assign n2238 = n2237 ^ n137 ;
  assign n2241 = n2240 ^ n2238 ;
  assign n2244 = n171 & ~n988 ;
  assign n2245 = n2244 ^ n171 ;
  assign n2242 = n160 & ~n1006 ;
  assign n2243 = n2242 ^ n160 ;
  assign n2246 = n2245 ^ n2243 ;
  assign n2247 = n2241 & n2246 ;
  assign n2248 = n2247 ^ n2241 ;
  assign n2249 = n2248 ^ n2246 ;
  assign n2250 = n254 & ~n2249 ;
  assign n2251 = n2250 ^ n254 ;
  assign n2267 = n2266 ^ n2251 ;
  assign n2268 = n2236 & n2267 ;
  assign n2269 = n2268 ^ n2236 ;
  assign n2270 = n2269 ^ n2267 ;
  assign n2271 = x134 & ~n2270 ;
  assign n2272 = n2271 ^ n2270 ;
  assign n2159 = n148 & ~n639 ;
  assign n2160 = n2159 ^ n148 ;
  assign n2157 = n137 & ~n657 ;
  assign n2158 = n2157 ^ n137 ;
  assign n2161 = n2160 ^ n2158 ;
  assign n2164 = n171 & ~n754 ;
  assign n2162 = n160 & ~n771 ;
  assign n2163 = n2162 ^ n160 ;
  assign n2165 = n2164 ^ n2163 ;
  assign n2166 = n2161 & n2165 ;
  assign n2167 = n2166 ^ n2161 ;
  assign n2168 = n2167 ^ n2165 ;
  assign n2169 = n254 & ~n2168 ;
  assign n2170 = n2169 ^ n254 ;
  assign n2144 = n148 & ~n945 ;
  assign n2145 = n2144 ^ n148 ;
  assign n2142 = n137 & ~n963 ;
  assign n2143 = n2142 ^ n137 ;
  assign n2146 = n2145 ^ n2143 ;
  assign n2149 = n171 & ~n602 ;
  assign n2150 = n2149 ^ n171 ;
  assign n2147 = n160 & ~n620 ;
  assign n2148 = n2147 ^ n160 ;
  assign n2151 = n2150 ^ n2148 ;
  assign n2152 = n2146 & n2151 ;
  assign n2153 = n2152 ^ n2146 ;
  assign n2154 = n2153 ^ n2151 ;
  assign n2155 = n279 & ~n2154 ;
  assign n2156 = n2155 ^ n279 ;
  assign n2171 = n2170 ^ n2156 ;
  assign n2189 = n148 & ~n783 ;
  assign n2187 = n137 & ~n800 ;
  assign n2188 = n2187 ^ n137 ;
  assign n2190 = n2189 ^ n2188 ;
  assign n2193 = n171 & ~n682 ;
  assign n2194 = n2193 ^ n171 ;
  assign n2191 = n160 & ~n700 ;
  assign n2192 = n2191 ^ n160 ;
  assign n2195 = n2194 ^ n2192 ;
  assign n2196 = n2190 & n2195 ;
  assign n2197 = n2196 ^ n2190 ;
  assign n2198 = n2197 ^ n2195 ;
  assign n2199 = n136 & ~n2198 ;
  assign n2200 = n2199 ^ n136 ;
  assign n2174 = n148 & ~n719 ;
  assign n2175 = n2174 ^ n148 ;
  assign n2172 = n137 & ~n737 ;
  assign n2173 = n2172 ^ n137 ;
  assign n2176 = n2175 ^ n2173 ;
  assign n2179 = n171 & ~n523 ;
  assign n2180 = n2179 ^ n171 ;
  assign n2177 = n160 & ~n541 ;
  assign n2178 = n2177 ^ n160 ;
  assign n2181 = n2180 ^ n2178 ;
  assign n2182 = n2176 & n2181 ;
  assign n2183 = n2182 ^ n2176 ;
  assign n2184 = n2183 ^ n2181 ;
  assign n2185 = n185 & ~n2184 ;
  assign n2186 = n2185 ^ n185 ;
  assign n2201 = n2200 ^ n2186 ;
  assign n2202 = n2171 & n2201 ;
  assign n2203 = n2202 ^ n2171 ;
  assign n2204 = n2203 ^ n2201 ;
  assign n2205 = x134 & ~n2204 ;
  assign n2273 = n2272 ^ n2205 ;
  assign n2319 = n148 & n1239 ;
  assign n2318 = n137 & n1243 ;
  assign n2320 = n2319 ^ n2318 ;
  assign n2322 = n171 & n1250 ;
  assign n2321 = n160 & n1254 ;
  assign n2323 = n2322 ^ n2321 ;
  assign n2324 = ~n2320 & ~n2323 ;
  assign n2325 = n185 & ~n2324 ;
  assign n2311 = n148 & n1280 ;
  assign n2310 = n137 & n1284 ;
  assign n2312 = n2311 ^ n2310 ;
  assign n2314 = n171 & n1230 ;
  assign n2313 = n160 & n1234 ;
  assign n2315 = n2314 ^ n2313 ;
  assign n2316 = ~n2312 & ~n2315 ;
  assign n2317 = n136 & ~n2316 ;
  assign n2326 = n2325 ^ n2317 ;
  assign n2336 = n148 & n1149 ;
  assign n2335 = n137 & n1153 ;
  assign n2337 = n2336 ^ n2335 ;
  assign n2339 = n171 & n1291 ;
  assign n2338 = n160 & n1295 ;
  assign n2340 = n2339 ^ n2338 ;
  assign n2341 = ~n2337 & ~n2340 ;
  assign n2342 = n279 & ~n2341 ;
  assign n2328 = n148 & n1300 ;
  assign n2327 = n137 & n1304 ;
  assign n2329 = n2328 ^ n2327 ;
  assign n2331 = n171 & n1271 ;
  assign n2330 = n160 & n1275 ;
  assign n2332 = n2331 ^ n2330 ;
  assign n2333 = ~n2329 & ~n2332 ;
  assign n2334 = n254 & ~n2333 ;
  assign n2343 = n2342 ^ n2334 ;
  assign n2344 = ~n2326 & ~n2343 ;
  assign n2345 = ~x134 & n2344 ;
  assign n2283 = n148 & n1169 ;
  assign n2282 = n137 & n1173 ;
  assign n2284 = n2283 ^ n2282 ;
  assign n2286 = n171 & n1201 ;
  assign n2285 = n160 & n1205 ;
  assign n2287 = n2286 ^ n2285 ;
  assign n2288 = ~n2284 & ~n2287 ;
  assign n2289 = n254 & ~n2288 ;
  assign n2275 = n148 & n1259 ;
  assign n2274 = n137 & n1263 ;
  assign n2276 = n2275 ^ n2274 ;
  assign n2278 = n171 & n1160 ;
  assign n2277 = n160 & n1164 ;
  assign n2279 = n2278 ^ n2277 ;
  assign n2280 = ~n2276 & ~n2279 ;
  assign n2281 = n279 & ~n2280 ;
  assign n2290 = n2289 ^ n2281 ;
  assign n2300 = n148 & ~n1213 ;
  assign n2299 = n137 & ~n1220 ;
  assign n2301 = n2300 ^ n2299 ;
  assign n2303 = n171 & n1181 ;
  assign n2302 = n160 & n1185 ;
  assign n2304 = n2303 ^ n2302 ;
  assign n2305 = ~n2301 & ~n2304 ;
  assign n2306 = n136 & ~n2305 ;
  assign n2292 = n148 & n1190 ;
  assign n2291 = n137 & n1194 ;
  assign n2293 = n2292 ^ n2291 ;
  assign n2295 = n171 & n1140 ;
  assign n2294 = n160 & n1144 ;
  assign n2296 = n2295 ^ n2294 ;
  assign n2297 = ~n2293 & ~n2296 ;
  assign n2298 = n185 & ~n2297 ;
  assign n2307 = n2306 ^ n2298 ;
  assign n2308 = ~n2290 & ~n2307 ;
  assign n2309 = x134 & n2308 ;
  assign n2346 = n2345 ^ n2309 ;
  assign n2429 = n148 & ~n1511 ;
  assign n2430 = n2429 ^ n148 ;
  assign n2427 = n137 & ~n1519 ;
  assign n2428 = n2427 ^ n137 ;
  assign n2431 = n2430 ^ n2428 ;
  assign n2434 = n171 & ~n1573 ;
  assign n2435 = n2434 ^ n171 ;
  assign n2432 = n160 & ~n1581 ;
  assign n2433 = n2432 ^ n160 ;
  assign n2436 = n2435 ^ n2433 ;
  assign n2437 = n2431 & n2436 ;
  assign n2438 = n2437 ^ n2431 ;
  assign n2439 = n2438 ^ n2436 ;
  assign n2440 = n185 & ~n2439 ;
  assign n2441 = n2440 ^ n185 ;
  assign n2414 = n148 & ~n1550 ;
  assign n2415 = n2414 ^ n148 ;
  assign n2412 = n137 & ~n1558 ;
  assign n2413 = n2412 ^ n137 ;
  assign n2416 = n2415 ^ n2413 ;
  assign n2419 = n171 & ~n1494 ;
  assign n2420 = n2419 ^ n171 ;
  assign n2417 = n160 & ~n1502 ;
  assign n2418 = n2417 ^ n160 ;
  assign n2421 = n2420 ^ n2418 ;
  assign n2422 = n2416 & n2421 ;
  assign n2423 = n2422 ^ n2416 ;
  assign n2424 = n2423 ^ n2421 ;
  assign n2425 = n136 & ~n2424 ;
  assign n2426 = n2425 ^ n136 ;
  assign n2442 = n2441 ^ n2426 ;
  assign n2460 = n148 & ~n1467 ;
  assign n2461 = n2460 ^ n148 ;
  assign n2458 = n137 & ~n1475 ;
  assign n2459 = n2458 ^ n137 ;
  assign n2462 = n2461 ^ n2459 ;
  assign n2465 = n171 & ~n1612 ;
  assign n2466 = n2465 ^ n171 ;
  assign n2463 = n160 & ~n1620 ;
  assign n2464 = n2463 ^ n160 ;
  assign n2467 = n2466 ^ n2464 ;
  assign n2468 = n2462 & n2467 ;
  assign n2469 = n2468 ^ n2462 ;
  assign n2470 = n2469 ^ n2467 ;
  assign n2471 = n279 & ~n2470 ;
  assign n2472 = n2471 ^ n279 ;
  assign n2445 = n148 & ~n1629 ;
  assign n2446 = n2445 ^ n148 ;
  assign n2443 = n137 & ~n1637 ;
  assign n2444 = n2443 ^ n137 ;
  assign n2447 = n2446 ^ n2444 ;
  assign n2450 = n171 & ~n1533 ;
  assign n2451 = n2450 ^ n171 ;
  assign n2448 = n160 & ~n1541 ;
  assign n2449 = n2448 ^ n160 ;
  assign n2452 = n2451 ^ n2449 ;
  assign n2453 = n2447 & n2452 ;
  assign n2454 = n2453 ^ n2447 ;
  assign n2455 = n2454 ^ n2452 ;
  assign n2456 = n254 & ~n2455 ;
  assign n2457 = n2456 ^ n254 ;
  assign n2473 = n2472 ^ n2457 ;
  assign n2474 = n2442 & n2473 ;
  assign n2475 = n2474 ^ n2442 ;
  assign n2476 = n2475 ^ n2473 ;
  assign n2477 = x134 & ~n2476 ;
  assign n2478 = n2477 ^ n2476 ;
  assign n2364 = n148 & ~n1388 ;
  assign n2365 = n2364 ^ n148 ;
  assign n2362 = n160 & ~n1325 ;
  assign n2363 = n2362 ^ n160 ;
  assign n2366 = n2365 ^ n2363 ;
  assign n2369 = n171 & ~n1318 ;
  assign n2367 = n137 & ~n1396 ;
  assign n2368 = n2367 ^ n137 ;
  assign n2370 = n2369 ^ n2368 ;
  assign n2371 = n2366 & n2370 ;
  assign n2372 = n2371 ^ n2366 ;
  assign n2373 = n2372 ^ n2370 ;
  assign n2374 = n254 & ~n2373 ;
  assign n2375 = n2374 ^ n254 ;
  assign n2349 = n148 & ~n1590 ;
  assign n2350 = n2349 ^ n148 ;
  assign n2347 = n137 & ~n1598 ;
  assign n2348 = n2347 ^ n137 ;
  assign n2351 = n2350 ^ n2348 ;
  assign n2354 = n171 & ~n1371 ;
  assign n2355 = n2354 ^ n171 ;
  assign n2352 = n160 & ~n1379 ;
  assign n2353 = n2352 ^ n160 ;
  assign n2356 = n2355 ^ n2353 ;
  assign n2357 = n2351 & n2356 ;
  assign n2358 = n2357 ^ n2351 ;
  assign n2359 = n2358 ^ n2356 ;
  assign n2360 = n279 & ~n2359 ;
  assign n2361 = n2360 ^ n279 ;
  assign n2376 = n2375 ^ n2361 ;
  assign n2394 = n148 & ~n1344 ;
  assign n2395 = n2394 ^ n148 ;
  assign n2392 = n137 & ~n1357 ;
  assign n2393 = n2392 ^ n137 ;
  assign n2396 = n2395 ^ n2393 ;
  assign n2399 = n171 & ~n1411 ;
  assign n2400 = n2399 ^ n171 ;
  assign n2397 = n160 & ~n1419 ;
  assign n2398 = n2397 ^ n160 ;
  assign n2401 = n2400 ^ n2398 ;
  assign n2402 = n2396 & n2401 ;
  assign n2403 = n2402 ^ n2396 ;
  assign n2404 = n2403 ^ n2401 ;
  assign n2405 = n136 & ~n2404 ;
  assign n2406 = n2405 ^ n136 ;
  assign n2379 = n148 & ~n1428 ;
  assign n2380 = n2379 ^ n148 ;
  assign n2377 = n137 & ~n1436 ;
  assign n2378 = n2377 ^ n137 ;
  assign n2381 = n2380 ^ n2378 ;
  assign n2384 = n171 & ~n1450 ;
  assign n2385 = n2384 ^ n171 ;
  assign n2382 = n160 & ~n1458 ;
  assign n2383 = n2382 ^ n160 ;
  assign n2386 = n2385 ^ n2383 ;
  assign n2387 = n2381 & n2386 ;
  assign n2388 = n2387 ^ n2381 ;
  assign n2389 = n2388 ^ n2386 ;
  assign n2390 = n185 & ~n2389 ;
  assign n2391 = n2390 ^ n185 ;
  assign n2407 = n2406 ^ n2391 ;
  assign n2408 = n2376 & n2407 ;
  assign n2409 = n2408 ^ n2376 ;
  assign n2410 = n2409 ^ n2407 ;
  assign n2411 = x134 & ~n2410 ;
  assign n2479 = n2478 ^ n2411 ;
  assign n2526 = n148 & n335 ;
  assign n2525 = n137 & n356 ;
  assign n2527 = n2526 ^ n2525 ;
  assign n2529 = n171 & n389 ;
  assign n2528 = n160 & n366 ;
  assign n2530 = n2529 ^ n2528 ;
  assign n2531 = ~n2527 & ~n2530 ;
  assign n2532 = n185 & ~n2531 ;
  assign n2518 = n148 & n424 ;
  assign n2517 = n137 & n445 ;
  assign n2519 = n2518 ^ n2517 ;
  assign n2521 = n171 & n345 ;
  assign n2520 = n160 & n455 ;
  assign n2522 = n2521 ^ n2520 ;
  assign n2523 = ~n2519 & ~n2522 ;
  assign n2524 = n136 & ~n2523 ;
  assign n2533 = n2532 ^ n2524 ;
  assign n2543 = n148 & n194 ;
  assign n2542 = n137 & n215 ;
  assign n2544 = n2543 ^ n2542 ;
  assign n2546 = n171 & n478 ;
  assign n2545 = n160 & n225 ;
  assign n2547 = n2546 ^ n2545 ;
  assign n2548 = ~n2544 & ~n2547 ;
  assign n2549 = n279 & ~n2548 ;
  assign n2535 = n148 & n468 ;
  assign n2534 = n137 & n489 ;
  assign n2536 = n2535 ^ n2534 ;
  assign n2538 = n171 & n434 ;
  assign n2537 = n160 & n499 ;
  assign n2539 = n2538 ^ n2537 ;
  assign n2540 = ~n2536 & ~n2539 ;
  assign n2541 = n254 & ~n2540 ;
  assign n2550 = n2549 ^ n2541 ;
  assign n2551 = ~n2533 & ~n2550 ;
  assign n2552 = ~x134 & n2551 ;
  assign n2489 = n148 & n288 ;
  assign n2488 = n137 & n309 ;
  assign n2490 = n2489 ^ n2488 ;
  assign n2492 = n171 & n273 ;
  assign n2491 = n160 & n319 ;
  assign n2493 = n2492 ^ n2491 ;
  assign n2494 = ~n2490 & ~n2493 ;
  assign n2495 = n254 & ~n2494 ;
  assign n2481 = n148 & n379 ;
  assign n2480 = n137 & n400 ;
  assign n2482 = n2481 ^ n2480 ;
  assign n2484 = n171 & n298 ;
  assign n2483 = n160 & n410 ;
  assign n2485 = n2484 ^ n2483 ;
  assign n2486 = ~n2482 & ~n2485 ;
  assign n2487 = n279 & ~n2486 ;
  assign n2496 = n2495 ^ n2487 ;
  assign n2507 = n146 & n148 ;
  assign n2506 = n137 & n169 ;
  assign n2508 = n2507 ^ n2506 ;
  assign n2510 = n171 & n204 ;
  assign n2509 = n160 & n180 ;
  assign n2511 = n2510 ^ n2509 ;
  assign n2512 = ~n2508 & ~n2511 ;
  assign n2513 = n185 & n2512 ;
  assign n2498 = n148 & n263 ;
  assign n2497 = n137 & ~n241 ;
  assign n2499 = n2498 ^ n2497 ;
  assign n2501 = n157 & n171 ;
  assign n2500 = n160 & n251 ;
  assign n2502 = n2501 ^ n2500 ;
  assign n2503 = n136 & ~n2502 ;
  assign n2504 = ~n2499 & n2503 ;
  assign n2505 = n2504 ^ x133 ;
  assign n2514 = n2513 ^ n2505 ;
  assign n2515 = ~n2496 & ~n2514 ;
  assign n2516 = x134 & n2515 ;
  assign n2553 = n2552 ^ n2516 ;
  assign n2633 = n148 & ~n829 ;
  assign n2634 = n2633 ^ n148 ;
  assign n2631 = n137 & ~n866 ;
  assign n2632 = n2631 ^ n137 ;
  assign n2635 = n2634 ^ n2632 ;
  assign n2638 = n171 & ~n926 ;
  assign n2639 = n2638 ^ n171 ;
  assign n2636 = n160 & ~n884 ;
  assign n2637 = n2636 ^ n160 ;
  assign n2640 = n2639 ^ n2637 ;
  assign n2641 = n2635 & n2640 ;
  assign n2642 = n2641 ^ n2635 ;
  assign n2643 = n2642 ^ n2640 ;
  assign n2644 = n185 & ~n2643 ;
  assign n2645 = n2644 ^ n185 ;
  assign n2618 = n148 & ~n988 ;
  assign n2619 = n2618 ^ n148 ;
  assign n2616 = n137 & ~n1025 ;
  assign n2617 = n2616 ^ n137 ;
  assign n2620 = n2619 ^ n2617 ;
  assign n2623 = n171 & ~n847 ;
  assign n2624 = n2623 ^ n171 ;
  assign n2621 = n160 & ~n1043 ;
  assign n2622 = n2621 ^ n160 ;
  assign n2625 = n2624 ^ n2622 ;
  assign n2626 = n2620 & n2625 ;
  assign n2627 = n2626 ^ n2620 ;
  assign n2628 = n2627 ^ n2625 ;
  assign n2629 = n136 & ~n2628 ;
  assign n2630 = n2629 ^ n136 ;
  assign n2646 = n2645 ^ n2630 ;
  assign n2664 = n148 & ~n523 ;
  assign n2665 = n2664 ^ n148 ;
  assign n2662 = n137 & ~n560 ;
  assign n2663 = n2662 ^ n137 ;
  assign n2666 = n2665 ^ n2663 ;
  assign n2669 = n171 & ~n1085 ;
  assign n2670 = n2669 ^ n171 ;
  assign n2667 = n160 & ~n578 ;
  assign n2668 = n2667 ^ n160 ;
  assign n2671 = n2670 ^ n2668 ;
  assign n2672 = n2666 & n2671 ;
  assign n2673 = n2672 ^ n2666 ;
  assign n2674 = n2673 ^ n2671 ;
  assign n2675 = n279 & ~n2674 ;
  assign n2676 = n2675 ^ n279 ;
  assign n2649 = n148 & ~n1067 ;
  assign n2650 = n2649 ^ n148 ;
  assign n2647 = n137 & ~n1104 ;
  assign n2648 = n2647 ^ n137 ;
  assign n2651 = n2650 ^ n2648 ;
  assign n2654 = n171 & ~n1006 ;
  assign n2655 = n2654 ^ n171 ;
  assign n2652 = n160 & ~n1122 ;
  assign n2653 = n2652 ^ n160 ;
  assign n2656 = n2655 ^ n2653 ;
  assign n2657 = n2651 & n2656 ;
  assign n2658 = n2657 ^ n2651 ;
  assign n2659 = n2658 ^ n2656 ;
  assign n2660 = n254 & ~n2659 ;
  assign n2661 = n2660 ^ n254 ;
  assign n2677 = n2676 ^ n2661 ;
  assign n2678 = n2646 & n2677 ;
  assign n2679 = n2678 ^ n2646 ;
  assign n2680 = n2679 ^ n2677 ;
  assign n2681 = x134 & ~n2680 ;
  assign n2682 = n2681 ^ n2680 ;
  assign n2571 = n148 & ~n602 ;
  assign n2572 = n2571 ^ n148 ;
  assign n2569 = n137 & ~n639 ;
  assign n2570 = n2569 ^ n137 ;
  assign n2573 = n2572 ^ n2570 ;
  assign n2576 = n171 & ~n771 ;
  assign n2577 = n2576 ^ n171 ;
  assign n2574 = n160 & ~n657 ;
  assign n2575 = n2574 ^ n160 ;
  assign n2578 = n2577 ^ n2575 ;
  assign n2579 = n2573 & n2578 ;
  assign n2580 = n2579 ^ n2573 ;
  assign n2581 = n2580 ^ n2578 ;
  assign n2582 = n254 & ~n2581 ;
  assign n2583 = n2582 ^ n254 ;
  assign n2556 = n148 & ~n908 ;
  assign n2557 = n2556 ^ n148 ;
  assign n2554 = n137 & ~n945 ;
  assign n2555 = n2554 ^ n137 ;
  assign n2558 = n2557 ^ n2555 ;
  assign n2561 = n171 & ~n620 ;
  assign n2562 = n2561 ^ n171 ;
  assign n2559 = n160 & ~n963 ;
  assign n2560 = n2559 ^ n160 ;
  assign n2563 = n2562 ^ n2560 ;
  assign n2564 = n2558 & n2563 ;
  assign n2565 = n2564 ^ n2558 ;
  assign n2566 = n2565 ^ n2563 ;
  assign n2567 = n279 & ~n2566 ;
  assign n2568 = n2567 ^ n279 ;
  assign n2584 = n2583 ^ n2568 ;
  assign n2602 = n171 & ~n700 ;
  assign n2603 = n2602 ^ n171 ;
  assign n2600 = n160 & ~n800 ;
  assign n2601 = n2600 ^ n160 ;
  assign n2604 = n2603 ^ n2601 ;
  assign n2606 = n148 & ~n754 ;
  assign n2605 = n137 & ~n783 ;
  assign n2607 = n2606 ^ n2605 ;
  assign n2608 = n136 & ~n2607 ;
  assign n2609 = ~n2604 & n2608 ;
  assign n2610 = n2609 ^ n136 ;
  assign n2587 = n148 & ~n682 ;
  assign n2588 = n2587 ^ n148 ;
  assign n2585 = n137 & ~n719 ;
  assign n2586 = n2585 ^ n137 ;
  assign n2589 = n2588 ^ n2586 ;
  assign n2592 = n171 & ~n541 ;
  assign n2593 = n2592 ^ n171 ;
  assign n2590 = n160 & ~n737 ;
  assign n2591 = n2590 ^ n160 ;
  assign n2594 = n2593 ^ n2591 ;
  assign n2595 = n2589 & n2594 ;
  assign n2596 = n2595 ^ n2589 ;
  assign n2597 = n2596 ^ n2594 ;
  assign n2598 = n185 & ~n2597 ;
  assign n2599 = n2598 ^ n185 ;
  assign n2611 = n2610 ^ n2599 ;
  assign n2612 = n2584 & n2611 ;
  assign n2613 = n2612 ^ n2584 ;
  assign n2614 = n2613 ^ n2611 ;
  assign n2615 = x134 & ~n2614 ;
  assign n2683 = n2682 ^ n2615 ;
  assign n2729 = n148 & n1230 ;
  assign n2728 = n137 & n1239 ;
  assign n2730 = n2729 ^ n2728 ;
  assign n2732 = n171 & n1254 ;
  assign n2731 = n160 & n1243 ;
  assign n2733 = n2732 ^ n2731 ;
  assign n2734 = ~n2730 & ~n2733 ;
  assign n2735 = n185 & ~n2734 ;
  assign n2721 = n148 & n1271 ;
  assign n2720 = n137 & n1280 ;
  assign n2722 = n2721 ^ n2720 ;
  assign n2724 = n171 & n1234 ;
  assign n2723 = n160 & n1284 ;
  assign n2725 = n2724 ^ n2723 ;
  assign n2726 = ~n2722 & ~n2725 ;
  assign n2727 = n136 & ~n2726 ;
  assign n2736 = n2735 ^ n2727 ;
  assign n2746 = n148 & n1140 ;
  assign n2745 = n137 & n1149 ;
  assign n2747 = n2746 ^ n2745 ;
  assign n2749 = n171 & n1295 ;
  assign n2748 = n160 & n1153 ;
  assign n2750 = n2749 ^ n2748 ;
  assign n2751 = ~n2747 & ~n2750 ;
  assign n2752 = n279 & ~n2751 ;
  assign n2738 = n148 & n1291 ;
  assign n2737 = n137 & n1300 ;
  assign n2739 = n2738 ^ n2737 ;
  assign n2741 = n171 & n1275 ;
  assign n2740 = n160 & n1304 ;
  assign n2742 = n2741 ^ n2740 ;
  assign n2743 = ~n2739 & ~n2742 ;
  assign n2744 = n254 & ~n2743 ;
  assign n2753 = n2752 ^ n2744 ;
  assign n2754 = ~n2736 & ~n2753 ;
  assign n2755 = ~x134 & n2754 ;
  assign n2693 = n148 & n1160 ;
  assign n2692 = n137 & n1169 ;
  assign n2694 = n2693 ^ n2692 ;
  assign n2696 = n171 & n1205 ;
  assign n2695 = n160 & n1173 ;
  assign n2697 = n2696 ^ n2695 ;
  assign n2698 = ~n2694 & ~n2697 ;
  assign n2699 = n254 & ~n2698 ;
  assign n2685 = n148 & n1250 ;
  assign n2684 = n137 & n1259 ;
  assign n2686 = n2685 ^ n2684 ;
  assign n2688 = n171 & n1164 ;
  assign n2687 = n160 & n1263 ;
  assign n2689 = n2688 ^ n2687 ;
  assign n2690 = ~n2686 & ~n2689 ;
  assign n2691 = n279 & ~n2690 ;
  assign n2700 = n2699 ^ n2691 ;
  assign n2710 = n148 & n1201 ;
  assign n2709 = n137 & ~n1213 ;
  assign n2711 = n2710 ^ n2709 ;
  assign n2713 = n171 & n1185 ;
  assign n2712 = n160 & ~n1220 ;
  assign n2714 = n2713 ^ n2712 ;
  assign n2715 = ~n2711 & ~n2714 ;
  assign n2716 = n136 & ~n2715 ;
  assign n2702 = n148 & n1181 ;
  assign n2701 = n137 & n1190 ;
  assign n2703 = n2702 ^ n2701 ;
  assign n2705 = n171 & n1144 ;
  assign n2704 = n160 & n1194 ;
  assign n2706 = n2705 ^ n2704 ;
  assign n2707 = ~n2703 & ~n2706 ;
  assign n2708 = n185 & ~n2707 ;
  assign n2717 = n2716 ^ n2708 ;
  assign n2718 = ~n2700 & ~n2717 ;
  assign n2719 = x134 & n2718 ;
  assign n2756 = n2755 ^ n2719 ;
  assign n2839 = n148 & ~n1494 ;
  assign n2840 = n2839 ^ n148 ;
  assign n2837 = n137 & ~n1511 ;
  assign n2838 = n2837 ^ n137 ;
  assign n2841 = n2840 ^ n2838 ;
  assign n2844 = n171 & ~n1581 ;
  assign n2845 = n2844 ^ n171 ;
  assign n2842 = n160 & ~n1519 ;
  assign n2843 = n2842 ^ n160 ;
  assign n2846 = n2845 ^ n2843 ;
  assign n2847 = n2841 & n2846 ;
  assign n2848 = n2847 ^ n2841 ;
  assign n2849 = n2848 ^ n2846 ;
  assign n2850 = n185 & ~n2849 ;
  assign n2851 = n2850 ^ n185 ;
  assign n2824 = n148 & ~n1533 ;
  assign n2825 = n2824 ^ n148 ;
  assign n2822 = n137 & ~n1550 ;
  assign n2823 = n2822 ^ n137 ;
  assign n2826 = n2825 ^ n2823 ;
  assign n2829 = n171 & ~n1502 ;
  assign n2830 = n2829 ^ n171 ;
  assign n2827 = n160 & ~n1558 ;
  assign n2828 = n2827 ^ n160 ;
  assign n2831 = n2830 ^ n2828 ;
  assign n2832 = n2826 & n2831 ;
  assign n2833 = n2832 ^ n2826 ;
  assign n2834 = n2833 ^ n2831 ;
  assign n2835 = n136 & ~n2834 ;
  assign n2836 = n2835 ^ n136 ;
  assign n2852 = n2851 ^ n2836 ;
  assign n2870 = n148 & ~n1450 ;
  assign n2871 = n2870 ^ n148 ;
  assign n2868 = n137 & ~n1467 ;
  assign n2869 = n2868 ^ n137 ;
  assign n2872 = n2871 ^ n2869 ;
  assign n2875 = n171 & ~n1620 ;
  assign n2876 = n2875 ^ n171 ;
  assign n2873 = n160 & ~n1475 ;
  assign n2874 = n2873 ^ n160 ;
  assign n2877 = n2876 ^ n2874 ;
  assign n2878 = n2872 & n2877 ;
  assign n2879 = n2878 ^ n2872 ;
  assign n2880 = n2879 ^ n2877 ;
  assign n2881 = n279 & ~n2880 ;
  assign n2882 = n2881 ^ n279 ;
  assign n2855 = n148 & ~n1612 ;
  assign n2856 = n2855 ^ n148 ;
  assign n2853 = n137 & ~n1629 ;
  assign n2854 = n2853 ^ n137 ;
  assign n2857 = n2856 ^ n2854 ;
  assign n2860 = n171 & ~n1541 ;
  assign n2861 = n2860 ^ n171 ;
  assign n2858 = n160 & ~n1637 ;
  assign n2859 = n2858 ^ n160 ;
  assign n2862 = n2861 ^ n2859 ;
  assign n2863 = n2857 & n2862 ;
  assign n2864 = n2863 ^ n2857 ;
  assign n2865 = n2864 ^ n2862 ;
  assign n2866 = n254 & ~n2865 ;
  assign n2867 = n2866 ^ n254 ;
  assign n2883 = n2882 ^ n2867 ;
  assign n2884 = n2852 & n2883 ;
  assign n2885 = n2884 ^ n2852 ;
  assign n2886 = n2885 ^ n2883 ;
  assign n2887 = x134 & ~n2886 ;
  assign n2888 = n2887 ^ n2886 ;
  assign n2774 = n148 & ~n1371 ;
  assign n2775 = n2774 ^ n148 ;
  assign n2772 = n137 & ~n1388 ;
  assign n2773 = n2772 ^ n137 ;
  assign n2776 = n2775 ^ n2773 ;
  assign n2779 = n171 & ~n1325 ;
  assign n2780 = n2779 ^ n171 ;
  assign n2777 = n160 & ~n1396 ;
  assign n2778 = n2777 ^ n160 ;
  assign n2781 = n2780 ^ n2778 ;
  assign n2782 = n2776 & n2781 ;
  assign n2783 = n2782 ^ n2776 ;
  assign n2784 = n2783 ^ n2781 ;
  assign n2785 = n254 & ~n2784 ;
  assign n2786 = n2785 ^ n254 ;
  assign n2759 = n148 & ~n1573 ;
  assign n2760 = n2759 ^ n148 ;
  assign n2757 = n137 & ~n1590 ;
  assign n2758 = n2757 ^ n137 ;
  assign n2761 = n2760 ^ n2758 ;
  assign n2764 = n171 & ~n1379 ;
  assign n2765 = n2764 ^ n171 ;
  assign n2762 = n160 & ~n1598 ;
  assign n2763 = n2762 ^ n160 ;
  assign n2766 = n2765 ^ n2763 ;
  assign n2767 = n2761 & n2766 ;
  assign n2768 = n2767 ^ n2761 ;
  assign n2769 = n2768 ^ n2766 ;
  assign n2770 = n279 & ~n2769 ;
  assign n2771 = n2770 ^ n279 ;
  assign n2787 = n2786 ^ n2771 ;
  assign n2805 = n148 & ~n1318 ;
  assign n2803 = n137 & ~n1344 ;
  assign n2804 = n2803 ^ n137 ;
  assign n2806 = n2805 ^ n2804 ;
  assign n2809 = n171 & ~n1419 ;
  assign n2810 = n2809 ^ n171 ;
  assign n2807 = n160 & ~n1357 ;
  assign n2808 = n2807 ^ n160 ;
  assign n2811 = n2810 ^ n2808 ;
  assign n2812 = n2806 & n2811 ;
  assign n2813 = n2812 ^ n2806 ;
  assign n2814 = n2813 ^ n2811 ;
  assign n2815 = n136 & ~n2814 ;
  assign n2816 = n2815 ^ n136 ;
  assign n2790 = n148 & ~n1411 ;
  assign n2791 = n2790 ^ n148 ;
  assign n2788 = n137 & ~n1428 ;
  assign n2789 = n2788 ^ n137 ;
  assign n2792 = n2791 ^ n2789 ;
  assign n2795 = n171 & ~n1458 ;
  assign n2796 = n2795 ^ n171 ;
  assign n2793 = n160 & ~n1436 ;
  assign n2794 = n2793 ^ n160 ;
  assign n2797 = n2796 ^ n2794 ;
  assign n2798 = n2792 & n2797 ;
  assign n2799 = n2798 ^ n2792 ;
  assign n2800 = n2799 ^ n2797 ;
  assign n2801 = n185 & ~n2800 ;
  assign n2802 = n2801 ^ n185 ;
  assign n2817 = n2816 ^ n2802 ;
  assign n2818 = n2787 & n2817 ;
  assign n2819 = n2818 ^ n2787 ;
  assign n2820 = n2819 ^ n2817 ;
  assign n2821 = x134 & ~n2820 ;
  assign n2889 = n2888 ^ n2821 ;
  assign n2902 = n185 & ~n369 ;
  assign n2901 = n136 & ~n458 ;
  assign n2903 = n2902 ^ n2901 ;
  assign n2905 = ~n228 & n279 ;
  assign n2904 = n254 & ~n502 ;
  assign n2906 = n2905 ^ n2904 ;
  assign n2907 = ~n2903 & ~n2906 ;
  assign n2908 = ~x134 & n2907 ;
  assign n2891 = n279 & ~n413 ;
  assign n2890 = ~n183 & n185 ;
  assign n2892 = n2891 ^ n2890 ;
  assign n2896 = n254 & n322 ;
  assign n2897 = n2896 ^ x133 ;
  assign n2893 = n136 & ~n275 ;
  assign n2894 = ~n253 & n2893 ;
  assign n2895 = n2894 ^ x132 ;
  assign n2898 = n2897 ^ n2895 ;
  assign n2899 = ~n2892 & ~n2898 ;
  assign n2900 = x134 & n2899 ;
  assign n2909 = n2908 ^ n2900 ;
  assign n2926 = n185 & ~n890 ;
  assign n2927 = n2926 ^ n185 ;
  assign n2924 = n136 & ~n1049 ;
  assign n2925 = n2924 ^ n136 ;
  assign n2928 = n2927 ^ n2925 ;
  assign n2931 = n279 & ~n584 ;
  assign n2932 = n2931 ^ n279 ;
  assign n2929 = n254 & ~n1128 ;
  assign n2930 = n2929 ^ n254 ;
  assign n2933 = n2932 ^ n2930 ;
  assign n2934 = n2928 & n2933 ;
  assign n2935 = n2934 ^ n2928 ;
  assign n2936 = n2935 ^ n2933 ;
  assign n2937 = x134 & ~n2936 ;
  assign n2938 = n2937 ^ n2936 ;
  assign n2912 = n254 & ~n663 ;
  assign n2913 = n2912 ^ n254 ;
  assign n2910 = n279 & ~n969 ;
  assign n2911 = n2910 ^ n279 ;
  assign n2914 = n2913 ^ n2911 ;
  assign n2917 = n136 & ~n806 ;
  assign n2918 = n2917 ^ n136 ;
  assign n2915 = n185 & ~n743 ;
  assign n2916 = n2915 ^ n185 ;
  assign n2919 = n2918 ^ n2916 ;
  assign n2920 = n2914 & n2919 ;
  assign n2921 = n2920 ^ n2914 ;
  assign n2922 = n2921 ^ n2919 ;
  assign n2923 = x134 & ~n2922 ;
  assign n2939 = n2938 ^ n2923 ;
  assign n2949 = n185 & ~n1246 ;
  assign n2948 = n136 & ~n1287 ;
  assign n2950 = n2949 ^ n2948 ;
  assign n2952 = n279 & ~n1156 ;
  assign n2951 = n254 & ~n1307 ;
  assign n2953 = n2952 ^ n2951 ;
  assign n2954 = ~n2950 & ~n2953 ;
  assign n2955 = ~x134 & n2954 ;
  assign n2941 = n254 & ~n1176 ;
  assign n2940 = n279 & ~n1266 ;
  assign n2942 = n2941 ^ n2940 ;
  assign n2944 = n136 & ~n1223 ;
  assign n2943 = n185 & ~n1197 ;
  assign n2945 = n2944 ^ n2943 ;
  assign n2946 = ~n2942 & ~n2945 ;
  assign n2947 = x134 & n2946 ;
  assign n2956 = n2955 ^ n2947 ;
  assign n2973 = n136 & ~n1564 ;
  assign n2974 = n2973 ^ n136 ;
  assign n2971 = n185 & ~n1525 ;
  assign n2972 = n2971 ^ n185 ;
  assign n2975 = n2974 ^ n2972 ;
  assign n2978 = n254 & ~n1643 ;
  assign n2979 = n2978 ^ n254 ;
  assign n2976 = n279 & ~n1481 ;
  assign n2977 = n2976 ^ n279 ;
  assign n2980 = n2979 ^ n2977 ;
  assign n2981 = n2975 & n2980 ;
  assign n2982 = n2981 ^ n2975 ;
  assign n2983 = n2982 ^ n2980 ;
  assign n2984 = x134 & ~n2983 ;
  assign n2985 = n2984 ^ n2983 ;
  assign n2959 = n254 & ~n1402 ;
  assign n2960 = n2959 ^ n254 ;
  assign n2957 = n279 & ~n1604 ;
  assign n2958 = n2957 ^ n279 ;
  assign n2961 = n2960 ^ n2958 ;
  assign n2964 = n185 & ~n1442 ;
  assign n2965 = n2964 ^ n185 ;
  assign n2962 = n136 & ~n1363 ;
  assign n2963 = n2962 ^ n136 ;
  assign n2966 = n2965 ^ n2963 ;
  assign n2967 = n2961 & n2966 ;
  assign n2968 = n2967 ^ n2961 ;
  assign n2969 = n2968 ^ n2966 ;
  assign n2970 = x134 & ~n2969 ;
  assign n2986 = n2985 ^ n2970 ;
  assign n2998 = n185 & ~n1696 ;
  assign n2997 = n136 & ~n1713 ;
  assign n2999 = n2998 ^ n2997 ;
  assign n3001 = n279 & ~n1677 ;
  assign n3000 = n254 & ~n1721 ;
  assign n3002 = n3001 ^ n3000 ;
  assign n3003 = ~n2999 & ~n3002 ;
  assign n3004 = ~x134 & n3003 ;
  assign n2990 = n279 & n1704 ;
  assign n2987 = n136 & ~n1666 ;
  assign n2988 = ~n1663 & n2987 ;
  assign n2989 = n2988 ^ x132 ;
  assign n2991 = n2990 ^ n2989 ;
  assign n2993 = n185 & ~n1685 ;
  assign n2992 = n254 & ~n1659 ;
  assign n2994 = n2993 ^ n2992 ;
  assign n2995 = n2991 & ~n2994 ;
  assign n2996 = x134 & n2995 ;
  assign n3005 = n3004 ^ n2996 ;
  assign n3027 = n185 & ~n1806 ;
  assign n3028 = n3027 ^ n185 ;
  assign n3025 = n136 & ~n1837 ;
  assign n3026 = n3025 ^ n136 ;
  assign n3029 = n3028 ^ n3026 ;
  assign n3032 = n279 & ~n1771 ;
  assign n3033 = n3032 ^ n279 ;
  assign n3030 = n254 & ~n1852 ;
  assign n3031 = n3030 ^ n254 ;
  assign n3034 = n3033 ^ n3031 ;
  assign n3035 = n3029 & n3034 ;
  assign n3036 = n3035 ^ n3029 ;
  assign n3037 = n3036 ^ n3034 ;
  assign n3038 = x134 & ~n3037 ;
  assign n3039 = n3038 ^ n3037 ;
  assign n3013 = n279 & ~n1821 ;
  assign n3014 = n3013 ^ n279 ;
  assign n3006 = n1744 ^ n136 ;
  assign n3007 = ~n136 & n3006 ;
  assign n3008 = n3007 ^ n136 ;
  assign n3009 = n3008 ^ n1749 ;
  assign n3010 = n1750 & n3009 ;
  assign n3011 = n3010 ^ n3007 ;
  assign n3012 = n3011 ^ n1749 ;
  assign n3015 = n3014 ^ n3012 ;
  assign n3018 = n185 & ~n1786 ;
  assign n3019 = n3018 ^ n185 ;
  assign n3016 = n254 & ~n1739 ;
  assign n3017 = n3016 ^ n254 ;
  assign n3020 = n3019 ^ n3017 ;
  assign n3021 = n3015 & n3020 ;
  assign n3022 = n3021 ^ n3015 ;
  assign n3023 = n3022 ^ n3020 ;
  assign n3024 = x134 & ~n3023 ;
  assign n3040 = n3039 ^ n3024 ;
  assign n3050 = n185 & ~n1904 ;
  assign n3049 = n136 & ~n1921 ;
  assign n3051 = n3050 ^ n3049 ;
  assign n3053 = n279 & ~n1885 ;
  assign n3052 = n254 & ~n1929 ;
  assign n3054 = n3053 ^ n3052 ;
  assign n3055 = ~n3051 & ~n3054 ;
  assign n3056 = ~x134 & n3055 ;
  assign n3042 = n279 & ~n1912 ;
  assign n3041 = n136 & ~n1876 ;
  assign n3043 = n3042 ^ n3041 ;
  assign n3045 = n185 & ~n1893 ;
  assign n3044 = n254 & ~n1868 ;
  assign n3046 = n3045 ^ n3044 ;
  assign n3047 = ~n3043 & ~n3046 ;
  assign n3048 = x134 & n3047 ;
  assign n3057 = n3056 ^ n3048 ;
  assign n3074 = n185 & ~n2012 ;
  assign n3075 = n3074 ^ n185 ;
  assign n3072 = n279 & ~n1977 ;
  assign n3073 = n3072 ^ n279 ;
  assign n3076 = n3075 ^ n3073 ;
  assign n3079 = n254 & ~n2058 ;
  assign n3080 = n3079 ^ n254 ;
  assign n3077 = n136 & ~n2043 ;
  assign n3078 = n3077 ^ n136 ;
  assign n3081 = n3080 ^ n3078 ;
  assign n3082 = n3076 & n3081 ;
  assign n3083 = n3082 ^ n3076 ;
  assign n3084 = n3083 ^ n3081 ;
  assign n3085 = x134 & ~n3084 ;
  assign n3086 = n3085 ^ n3084 ;
  assign n3060 = n136 & ~n1961 ;
  assign n3061 = n3060 ^ n136 ;
  assign n3058 = n254 & ~n1947 ;
  assign n3059 = n3058 ^ n254 ;
  assign n3062 = n3061 ^ n3059 ;
  assign n3065 = n185 & ~n1992 ;
  assign n3066 = n3065 ^ n185 ;
  assign n3063 = n279 & ~n2027 ;
  assign n3064 = n3063 ^ n279 ;
  assign n3067 = n3066 ^ n3064 ;
  assign n3068 = n3062 & n3067 ;
  assign n3069 = n3068 ^ n3062 ;
  assign n3070 = n3069 ^ n3067 ;
  assign n3071 = x134 & ~n3070 ;
  assign n3087 = n3086 ^ n3071 ;
  assign n3100 = n185 & ~n2111 ;
  assign n3099 = n279 & ~n2100 ;
  assign n3101 = n3100 ^ n3099 ;
  assign n3103 = n254 & ~n2136 ;
  assign n3102 = n136 & ~n2128 ;
  assign n3104 = n3103 ^ n3102 ;
  assign n3105 = ~n3101 & ~n3104 ;
  assign n3106 = ~x134 & n3105 ;
  assign n3089 = n136 & ~n2082 ;
  assign n3088 = n254 & ~n2074 ;
  assign n3090 = n3089 ^ n3088 ;
  assign n3094 = n279 & n2119 ;
  assign n3095 = n3094 ^ x133 ;
  assign n3091 = n185 & ~n2090 ;
  assign n3092 = ~n2087 & n3091 ;
  assign n3093 = n3092 ^ x132 ;
  assign n3096 = n3095 ^ n3093 ;
  assign n3097 = ~n3090 & n3096 ;
  assign n3098 = x134 & n3097 ;
  assign n3107 = n3106 ^ n3098 ;
  assign n3124 = n185 & ~n2218 ;
  assign n3125 = n3124 ^ n185 ;
  assign n3122 = n279 & ~n2184 ;
  assign n3123 = n3122 ^ n279 ;
  assign n3126 = n3125 ^ n3123 ;
  assign n3129 = n254 & ~n2264 ;
  assign n3130 = n3129 ^ n254 ;
  assign n3127 = n136 & ~n2249 ;
  assign n3128 = n3127 ^ n136 ;
  assign n3131 = n3130 ^ n3128 ;
  assign n3132 = n3126 & n3131 ;
  assign n3133 = n3132 ^ n3126 ;
  assign n3134 = n3133 ^ n3131 ;
  assign n3135 = x134 & ~n3134 ;
  assign n3136 = n3135 ^ n3134 ;
  assign n3110 = n136 & ~n2168 ;
  assign n3111 = n3110 ^ n136 ;
  assign n3108 = n254 & ~n2154 ;
  assign n3109 = n3108 ^ n254 ;
  assign n3112 = n3111 ^ n3109 ;
  assign n3115 = n185 & ~n2198 ;
  assign n3116 = n3115 ^ n185 ;
  assign n3113 = n279 & ~n2233 ;
  assign n3114 = n3113 ^ n279 ;
  assign n3117 = n3116 ^ n3114 ;
  assign n3118 = n3112 & n3117 ;
  assign n3119 = n3118 ^ n3112 ;
  assign n3120 = n3119 ^ n3117 ;
  assign n3121 = x134 & ~n3120 ;
  assign n3137 = n3136 ^ n3121 ;
  assign n3147 = n185 & ~n2316 ;
  assign n3146 = n136 & ~n2333 ;
  assign n3148 = n3147 ^ n3146 ;
  assign n3150 = n279 & ~n2297 ;
  assign n3149 = n254 & ~n2341 ;
  assign n3151 = n3150 ^ n3149 ;
  assign n3152 = ~n3148 & ~n3151 ;
  assign n3153 = ~x134 & n3152 ;
  assign n3139 = n136 & ~n2288 ;
  assign n3138 = n254 & ~n2280 ;
  assign n3140 = n3139 ^ n3138 ;
  assign n3142 = n185 & ~n2305 ;
  assign n3141 = n279 & ~n2324 ;
  assign n3143 = n3142 ^ n3141 ;
  assign n3144 = ~n3140 & ~n3143 ;
  assign n3145 = x134 & n3144 ;
  assign n3154 = n3153 ^ n3145 ;
  assign n3171 = n185 & ~n2424 ;
  assign n3172 = n3171 ^ n185 ;
  assign n3169 = n136 & ~n2455 ;
  assign n3170 = n3169 ^ n136 ;
  assign n3173 = n3172 ^ n3170 ;
  assign n3176 = n279 & ~n2389 ;
  assign n3177 = n3176 ^ n279 ;
  assign n3174 = n254 & ~n2470 ;
  assign n3175 = n3174 ^ n254 ;
  assign n3178 = n3177 ^ n3175 ;
  assign n3179 = n3173 & n3178 ;
  assign n3180 = n3179 ^ n3173 ;
  assign n3181 = n3180 ^ n3178 ;
  assign n3182 = x134 & ~n3181 ;
  assign n3183 = n3182 ^ n3181 ;
  assign n3157 = n136 & ~n2373 ;
  assign n3158 = n3157 ^ n136 ;
  assign n3155 = n254 & ~n2359 ;
  assign n3156 = n3155 ^ n254 ;
  assign n3159 = n3158 ^ n3156 ;
  assign n3162 = n185 & ~n2404 ;
  assign n3163 = n3162 ^ n185 ;
  assign n3160 = n279 & ~n2439 ;
  assign n3161 = n3160 ^ n279 ;
  assign n3164 = n3163 ^ n3161 ;
  assign n3165 = n3159 & n3164 ;
  assign n3166 = n3165 ^ n3159 ;
  assign n3167 = n3166 ^ n3164 ;
  assign n3168 = x134 & ~n3167 ;
  assign n3184 = n3183 ^ n3168 ;
  assign n3197 = n185 & ~n2523 ;
  assign n3196 = n136 & ~n2540 ;
  assign n3198 = n3197 ^ n3196 ;
  assign n3200 = n279 & ~n2512 ;
  assign n3199 = n254 & ~n2548 ;
  assign n3201 = n3200 ^ n3199 ;
  assign n3202 = ~n3198 & ~n3201 ;
  assign n3203 = ~x134 & n3202 ;
  assign n3186 = n136 & ~n2494 ;
  assign n3185 = n254 & ~n2486 ;
  assign n3187 = n3186 ^ n3185 ;
  assign n3191 = n279 & n2531 ;
  assign n3192 = n3191 ^ x133 ;
  assign n3188 = n185 & ~n2502 ;
  assign n3189 = ~n2499 & n3188 ;
  assign n3190 = n3189 ^ x132 ;
  assign n3193 = n3192 ^ n3190 ;
  assign n3194 = ~n3187 & n3193 ;
  assign n3195 = x134 & n3194 ;
  assign n3204 = n3203 ^ n3195 ;
  assign n3222 = n185 & ~n2628 ;
  assign n3223 = n3222 ^ n185 ;
  assign n3220 = n136 & ~n2659 ;
  assign n3221 = n3220 ^ n136 ;
  assign n3224 = n3223 ^ n3221 ;
  assign n3227 = n279 & ~n2597 ;
  assign n3228 = n3227 ^ n279 ;
  assign n3225 = n254 & ~n2674 ;
  assign n3226 = n3225 ^ n254 ;
  assign n3229 = n3228 ^ n3226 ;
  assign n3230 = n3224 & n3229 ;
  assign n3231 = n3230 ^ n3224 ;
  assign n3232 = n3231 ^ n3229 ;
  assign n3233 = x134 & ~n3232 ;
  assign n3234 = n3233 ^ n3232 ;
  assign n3207 = n136 & ~n2581 ;
  assign n3208 = n3207 ^ n136 ;
  assign n3205 = n254 & ~n2566 ;
  assign n3206 = n3205 ^ n254 ;
  assign n3209 = n3208 ^ n3206 ;
  assign n3212 = n185 & ~n2607 ;
  assign n3213 = ~n2604 & n3212 ;
  assign n3214 = n3213 ^ n185 ;
  assign n3210 = n279 & ~n2643 ;
  assign n3211 = n3210 ^ n279 ;
  assign n3215 = n3214 ^ n3211 ;
  assign n3216 = n3209 & n3215 ;
  assign n3217 = n3216 ^ n3209 ;
  assign n3218 = n3217 ^ n3215 ;
  assign n3219 = x134 & ~n3218 ;
  assign n3235 = n3234 ^ n3219 ;
  assign n3245 = n185 & ~n2726 ;
  assign n3244 = n136 & ~n2743 ;
  assign n3246 = n3245 ^ n3244 ;
  assign n3248 = n279 & ~n2707 ;
  assign n3247 = n254 & ~n2751 ;
  assign n3249 = n3248 ^ n3247 ;
  assign n3250 = ~n3246 & ~n3249 ;
  assign n3251 = ~x134 & n3250 ;
  assign n3237 = n136 & ~n2698 ;
  assign n3236 = n254 & ~n2690 ;
  assign n3238 = n3237 ^ n3236 ;
  assign n3240 = n185 & ~n2715 ;
  assign n3239 = n279 & ~n2734 ;
  assign n3241 = n3240 ^ n3239 ;
  assign n3242 = ~n3238 & ~n3241 ;
  assign n3243 = x134 & n3242 ;
  assign n3252 = n3251 ^ n3243 ;
  assign n3269 = n185 & ~n2834 ;
  assign n3270 = n3269 ^ n185 ;
  assign n3267 = n136 & ~n2865 ;
  assign n3268 = n3267 ^ n136 ;
  assign n3271 = n3270 ^ n3268 ;
  assign n3274 = n279 & ~n2800 ;
  assign n3275 = n3274 ^ n279 ;
  assign n3272 = n254 & ~n2880 ;
  assign n3273 = n3272 ^ n254 ;
  assign n3276 = n3275 ^ n3273 ;
  assign n3277 = n3271 & n3276 ;
  assign n3278 = n3277 ^ n3271 ;
  assign n3279 = n3278 ^ n3276 ;
  assign n3280 = x134 & ~n3279 ;
  assign n3281 = n3280 ^ n3279 ;
  assign n3255 = n136 & ~n2784 ;
  assign n3256 = n3255 ^ n136 ;
  assign n3253 = n254 & ~n2769 ;
  assign n3254 = n3253 ^ n254 ;
  assign n3257 = n3256 ^ n3254 ;
  assign n3260 = n185 & ~n2814 ;
  assign n3261 = n3260 ^ n185 ;
  assign n3258 = n279 & ~n2849 ;
  assign n3259 = n3258 ^ n279 ;
  assign n3262 = n3261 ^ n3259 ;
  assign n3263 = n3257 & n3262 ;
  assign n3264 = n3263 ^ n3257 ;
  assign n3265 = n3264 ^ n3262 ;
  assign n3266 = x134 & ~n3265 ;
  assign n3282 = n3281 ^ n3266 ;
  assign n3294 = n185 & ~n458 ;
  assign n3293 = n136 & ~n502 ;
  assign n3295 = n3294 ^ n3293 ;
  assign n3297 = ~n183 & n279 ;
  assign n3296 = ~n228 & n254 ;
  assign n3298 = n3297 ^ n3296 ;
  assign n3299 = ~n3295 & ~n3298 ;
  assign n3300 = ~x134 & n3299 ;
  assign n3284 = n254 & ~n413 ;
  assign n3283 = n279 & ~n369 ;
  assign n3285 = n3284 ^ n3283 ;
  assign n3287 = n185 & ~n275 ;
  assign n3288 = ~n253 & n3287 ;
  assign n3286 = n136 & n322 ;
  assign n3289 = n3288 ^ n3286 ;
  assign n3290 = n3289 ^ x133 ;
  assign n3291 = ~n3285 & ~n3290 ;
  assign n3292 = x134 & n3291 ;
  assign n3301 = n3300 ^ n3292 ;
  assign n3318 = n185 & ~n1049 ;
  assign n3319 = n3318 ^ n185 ;
  assign n3316 = n136 & ~n1128 ;
  assign n3317 = n3316 ^ n136 ;
  assign n3320 = n3319 ^ n3317 ;
  assign n3323 = n279 & ~n743 ;
  assign n3324 = n3323 ^ n279 ;
  assign n3321 = n254 & ~n584 ;
  assign n3322 = n3321 ^ n254 ;
  assign n3325 = n3324 ^ n3322 ;
  assign n3326 = n3320 & n3325 ;
  assign n3327 = n3326 ^ n3320 ;
  assign n3328 = n3327 ^ n3325 ;
  assign n3329 = x134 & ~n3328 ;
  assign n3330 = n3329 ^ n3328 ;
  assign n3304 = n136 & ~n663 ;
  assign n3305 = n3304 ^ n136 ;
  assign n3302 = n254 & ~n969 ;
  assign n3303 = n3302 ^ n254 ;
  assign n3306 = n3305 ^ n3303 ;
  assign n3309 = n185 & ~n806 ;
  assign n3310 = n3309 ^ n185 ;
  assign n3307 = n279 & ~n890 ;
  assign n3308 = n3307 ^ n279 ;
  assign n3311 = n3310 ^ n3308 ;
  assign n3312 = n3306 & n3311 ;
  assign n3313 = n3312 ^ n3306 ;
  assign n3314 = n3313 ^ n3311 ;
  assign n3315 = x134 & ~n3314 ;
  assign n3331 = n3330 ^ n3315 ;
  assign n3341 = n185 & ~n1287 ;
  assign n3340 = n136 & ~n1307 ;
  assign n3342 = n3341 ^ n3340 ;
  assign n3344 = n279 & ~n1197 ;
  assign n3343 = n254 & ~n1156 ;
  assign n3345 = n3344 ^ n3343 ;
  assign n3346 = ~n3342 & ~n3345 ;
  assign n3347 = ~x134 & n3346 ;
  assign n3333 = n136 & ~n1176 ;
  assign n3332 = n254 & ~n1266 ;
  assign n3334 = n3333 ^ n3332 ;
  assign n3336 = n185 & ~n1223 ;
  assign n3335 = n279 & ~n1246 ;
  assign n3337 = n3336 ^ n3335 ;
  assign n3338 = ~n3334 & ~n3337 ;
  assign n3339 = x134 & n3338 ;
  assign n3348 = n3347 ^ n3339 ;
  assign n3365 = n185 & ~n1564 ;
  assign n3366 = n3365 ^ n185 ;
  assign n3363 = n279 & ~n1442 ;
  assign n3364 = n3363 ^ n279 ;
  assign n3367 = n3366 ^ n3364 ;
  assign n3370 = n136 & ~n1643 ;
  assign n3371 = n3370 ^ n136 ;
  assign n3368 = n254 & ~n1481 ;
  assign n3369 = n3368 ^ n254 ;
  assign n3372 = n3371 ^ n3369 ;
  assign n3373 = n3367 & n3372 ;
  assign n3374 = n3373 ^ n3367 ;
  assign n3375 = n3374 ^ n3372 ;
  assign n3376 = x134 & ~n3375 ;
  assign n3377 = n3376 ^ n3375 ;
  assign n3351 = n136 & ~n1402 ;
  assign n3352 = n3351 ^ n136 ;
  assign n3349 = n279 & ~n1525 ;
  assign n3350 = n3349 ^ n279 ;
  assign n3353 = n3352 ^ n3350 ;
  assign n3356 = n185 & ~n1363 ;
  assign n3357 = n3356 ^ n185 ;
  assign n3354 = n254 & ~n1604 ;
  assign n3355 = n3354 ^ n254 ;
  assign n3358 = n3357 ^ n3355 ;
  assign n3359 = n3353 & n3358 ;
  assign n3360 = n3359 ^ n3353 ;
  assign n3361 = n3360 ^ n3358 ;
  assign n3362 = x134 & ~n3361 ;
  assign n3378 = n3377 ^ n3362 ;
  assign n3390 = n185 & ~n1713 ;
  assign n3389 = n136 & ~n1721 ;
  assign n3391 = n3390 ^ n3389 ;
  assign n3393 = n279 & ~n1685 ;
  assign n3392 = n254 & ~n1677 ;
  assign n3394 = n3393 ^ n3392 ;
  assign n3395 = ~n3391 & ~n3394 ;
  assign n3396 = ~x134 & n3395 ;
  assign n3380 = n254 & ~n1704 ;
  assign n3379 = n279 & ~n1696 ;
  assign n3381 = n3380 ^ n3379 ;
  assign n3385 = n136 & n1659 ;
  assign n3382 = n185 & ~n1666 ;
  assign n3383 = ~n1663 & n3382 ;
  assign n3384 = n3383 ^ x133 ;
  assign n3386 = n3385 ^ n3384 ;
  assign n3387 = ~n3381 & ~n3386 ;
  assign n3388 = x134 & n3387 ;
  assign n3397 = n3396 ^ n3388 ;
  assign n3419 = n185 & ~n1837 ;
  assign n3420 = n3419 ^ n185 ;
  assign n3417 = n136 & ~n1852 ;
  assign n3418 = n3417 ^ n136 ;
  assign n3421 = n3420 ^ n3418 ;
  assign n3424 = n279 & ~n1786 ;
  assign n3425 = n3424 ^ n279 ;
  assign n3422 = n254 & ~n1771 ;
  assign n3423 = n3422 ^ n254 ;
  assign n3426 = n3425 ^ n3423 ;
  assign n3427 = n3421 & n3426 ;
  assign n3428 = n3427 ^ n3421 ;
  assign n3429 = n3428 ^ n3426 ;
  assign n3430 = x134 & ~n3429 ;
  assign n3431 = n3430 ^ n3429 ;
  assign n3400 = n254 & ~n1821 ;
  assign n3401 = n3400 ^ n254 ;
  assign n3398 = n279 & ~n1806 ;
  assign n3399 = n3398 ^ n279 ;
  assign n3402 = n3401 ^ n3399 ;
  assign n3410 = n136 & ~n1739 ;
  assign n3411 = n3410 ^ n136 ;
  assign n3403 = n1744 ^ n185 ;
  assign n3404 = ~n185 & n3403 ;
  assign n3405 = n3404 ^ n185 ;
  assign n3406 = n3405 ^ n1749 ;
  assign n3407 = n1750 & n3406 ;
  assign n3408 = n3407 ^ n3404 ;
  assign n3409 = n3408 ^ n1749 ;
  assign n3412 = n3411 ^ n3409 ;
  assign n3413 = n3402 & n3412 ;
  assign n3414 = n3413 ^ n3402 ;
  assign n3415 = n3414 ^ n3412 ;
  assign n3416 = x134 & ~n3415 ;
  assign n3432 = n3431 ^ n3416 ;
  assign n3442 = n185 & ~n1921 ;
  assign n3441 = n136 & ~n1929 ;
  assign n3443 = n3442 ^ n3441 ;
  assign n3445 = n279 & ~n1893 ;
  assign n3444 = n254 & ~n1885 ;
  assign n3446 = n3445 ^ n3444 ;
  assign n3447 = ~n3443 & ~n3446 ;
  assign n3448 = ~x134 & n3447 ;
  assign n3434 = n254 & ~n1912 ;
  assign n3433 = n279 & ~n1904 ;
  assign n3435 = n3434 ^ n3433 ;
  assign n3437 = n136 & ~n1868 ;
  assign n3436 = n185 & ~n1876 ;
  assign n3438 = n3437 ^ n3436 ;
  assign n3439 = ~n3435 & ~n3438 ;
  assign n3440 = x134 & n3439 ;
  assign n3449 = n3448 ^ n3440 ;
  assign n3466 = n254 & ~n1977 ;
  assign n3467 = n3466 ^ n254 ;
  assign n3464 = n279 & ~n1992 ;
  assign n3465 = n3464 ^ n279 ;
  assign n3468 = n3467 ^ n3465 ;
  assign n3471 = n136 & ~n2058 ;
  assign n3472 = n3471 ^ n136 ;
  assign n3469 = n185 & ~n2043 ;
  assign n3470 = n3469 ^ n185 ;
  assign n3473 = n3472 ^ n3470 ;
  assign n3474 = n3468 & n3473 ;
  assign n3475 = n3474 ^ n3468 ;
  assign n3476 = n3475 ^ n3473 ;
  assign n3477 = x134 & ~n3476 ;
  assign n3478 = n3477 ^ n3476 ;
  assign n3452 = n185 & ~n1961 ;
  assign n3453 = n3452 ^ n185 ;
  assign n3450 = n136 & ~n1947 ;
  assign n3451 = n3450 ^ n136 ;
  assign n3454 = n3453 ^ n3451 ;
  assign n3457 = n279 & ~n2012 ;
  assign n3458 = n3457 ^ n279 ;
  assign n3455 = n254 & ~n2027 ;
  assign n3456 = n3455 ^ n254 ;
  assign n3459 = n3458 ^ n3456 ;
  assign n3460 = n3454 & n3459 ;
  assign n3461 = n3460 ^ n3454 ;
  assign n3462 = n3461 ^ n3459 ;
  assign n3463 = x134 & ~n3462 ;
  assign n3479 = n3478 ^ n3463 ;
  assign n3491 = n254 & n2100 ;
  assign n3488 = n279 & ~n2090 ;
  assign n3489 = ~n2087 & n3488 ;
  assign n3490 = n3489 ^ x133 ;
  assign n3492 = n3491 ^ n3490 ;
  assign n3494 = n136 & ~n2136 ;
  assign n3493 = n185 & ~n2128 ;
  assign n3495 = n3494 ^ n3493 ;
  assign n3496 = n3492 & ~n3495 ;
  assign n3497 = ~x134 & n3496 ;
  assign n3481 = n185 & ~n2082 ;
  assign n3480 = n136 & ~n2074 ;
  assign n3482 = n3481 ^ n3480 ;
  assign n3484 = n279 & ~n2111 ;
  assign n3483 = n254 & ~n2119 ;
  assign n3485 = n3484 ^ n3483 ;
  assign n3486 = ~n3482 & ~n3485 ;
  assign n3487 = x134 & n3486 ;
  assign n3498 = n3497 ^ n3487 ;
  assign n3515 = n254 & ~n2184 ;
  assign n3516 = n3515 ^ n254 ;
  assign n3513 = n279 & ~n2198 ;
  assign n3514 = n3513 ^ n279 ;
  assign n3517 = n3516 ^ n3514 ;
  assign n3520 = n136 & ~n2264 ;
  assign n3521 = n3520 ^ n136 ;
  assign n3518 = n185 & ~n2249 ;
  assign n3519 = n3518 ^ n185 ;
  assign n3522 = n3521 ^ n3519 ;
  assign n3523 = n3517 & n3522 ;
  assign n3524 = n3523 ^ n3517 ;
  assign n3525 = n3524 ^ n3522 ;
  assign n3526 = x134 & ~n3525 ;
  assign n3527 = n3526 ^ n3525 ;
  assign n3501 = n185 & ~n2168 ;
  assign n3502 = n3501 ^ n185 ;
  assign n3499 = n136 & ~n2154 ;
  assign n3500 = n3499 ^ n136 ;
  assign n3503 = n3502 ^ n3500 ;
  assign n3506 = n279 & ~n2218 ;
  assign n3507 = n3506 ^ n279 ;
  assign n3504 = n254 & ~n2233 ;
  assign n3505 = n3504 ^ n254 ;
  assign n3508 = n3507 ^ n3505 ;
  assign n3509 = n3503 & n3508 ;
  assign n3510 = n3509 ^ n3503 ;
  assign n3511 = n3510 ^ n3508 ;
  assign n3512 = x134 & ~n3511 ;
  assign n3528 = n3527 ^ n3512 ;
  assign n3538 = n185 & ~n2333 ;
  assign n3537 = n136 & ~n2341 ;
  assign n3539 = n3538 ^ n3537 ;
  assign n3541 = n279 & ~n2305 ;
  assign n3540 = n254 & ~n2297 ;
  assign n3542 = n3541 ^ n3540 ;
  assign n3543 = ~n3539 & ~n3542 ;
  assign n3544 = ~x134 & n3543 ;
  assign n3530 = n185 & ~n2288 ;
  assign n3529 = n136 & ~n2280 ;
  assign n3531 = n3530 ^ n3529 ;
  assign n3533 = n279 & ~n2316 ;
  assign n3532 = n254 & ~n2324 ;
  assign n3534 = n3533 ^ n3532 ;
  assign n3535 = ~n3531 & ~n3534 ;
  assign n3536 = x134 & n3535 ;
  assign n3545 = n3544 ^ n3536 ;
  assign n3562 = n185 & ~n2455 ;
  assign n3563 = n3562 ^ n185 ;
  assign n3560 = n136 & ~n2470 ;
  assign n3561 = n3560 ^ n136 ;
  assign n3564 = n3563 ^ n3561 ;
  assign n3567 = n279 & ~n2404 ;
  assign n3568 = n3567 ^ n279 ;
  assign n3565 = n254 & ~n2389 ;
  assign n3566 = n3565 ^ n254 ;
  assign n3569 = n3568 ^ n3566 ;
  assign n3570 = n3564 & n3569 ;
  assign n3571 = n3570 ^ n3564 ;
  assign n3572 = n3571 ^ n3569 ;
  assign n3573 = x134 & ~n3572 ;
  assign n3574 = n3573 ^ n3572 ;
  assign n3548 = n185 & ~n2373 ;
  assign n3549 = n3548 ^ n185 ;
  assign n3546 = n136 & ~n2359 ;
  assign n3547 = n3546 ^ n136 ;
  assign n3550 = n3549 ^ n3547 ;
  assign n3553 = n279 & ~n2424 ;
  assign n3554 = n3553 ^ n279 ;
  assign n3551 = n254 & ~n2439 ;
  assign n3552 = n3551 ^ n254 ;
  assign n3555 = n3554 ^ n3552 ;
  assign n3556 = n3550 & n3555 ;
  assign n3557 = n3556 ^ n3550 ;
  assign n3558 = n3557 ^ n3555 ;
  assign n3559 = x134 & ~n3558 ;
  assign n3575 = n3574 ^ n3559 ;
  assign n3585 = n185 & ~n2540 ;
  assign n3584 = n136 & ~n2548 ;
  assign n3586 = n3585 ^ n3584 ;
  assign n3590 = n254 & n2512 ;
  assign n3587 = n279 & ~n2502 ;
  assign n3588 = ~n2499 & n3587 ;
  assign n3589 = n3588 ^ x133 ;
  assign n3591 = n3590 ^ n3589 ;
  assign n3592 = ~n3586 & n3591 ;
  assign n3593 = ~x134 & n3592 ;
  assign n3577 = n185 & ~n2494 ;
  assign n3576 = n136 & ~n2486 ;
  assign n3578 = n3577 ^ n3576 ;
  assign n3580 = n279 & ~n2523 ;
  assign n3579 = n254 & ~n2531 ;
  assign n3581 = n3580 ^ n3579 ;
  assign n3582 = ~n3578 & ~n3581 ;
  assign n3583 = x134 & n3582 ;
  assign n3594 = n3593 ^ n3583 ;
  assign n3611 = n185 & ~n2659 ;
  assign n3612 = n3611 ^ n185 ;
  assign n3609 = n136 & ~n2674 ;
  assign n3610 = n3609 ^ n136 ;
  assign n3613 = n3612 ^ n3610 ;
  assign n3616 = n279 & ~n2607 ;
  assign n3617 = ~n2604 & n3616 ;
  assign n3618 = n3617 ^ n279 ;
  assign n3614 = n254 & ~n2597 ;
  assign n3615 = n3614 ^ n254 ;
  assign n3619 = n3618 ^ n3615 ;
  assign n3620 = n3613 & n3619 ;
  assign n3621 = n3620 ^ n3613 ;
  assign n3622 = n3621 ^ n3619 ;
  assign n3623 = x134 & ~n3622 ;
  assign n3624 = n3623 ^ n3622 ;
  assign n3597 = n185 & ~n2581 ;
  assign n3598 = n3597 ^ n185 ;
  assign n3595 = n136 & ~n2566 ;
  assign n3596 = n3595 ^ n136 ;
  assign n3599 = n3598 ^ n3596 ;
  assign n3602 = n279 & ~n2628 ;
  assign n3603 = n3602 ^ n279 ;
  assign n3600 = n254 & ~n2643 ;
  assign n3601 = n3600 ^ n254 ;
  assign n3604 = n3603 ^ n3601 ;
  assign n3605 = n3599 & n3604 ;
  assign n3606 = n3605 ^ n3599 ;
  assign n3607 = n3606 ^ n3604 ;
  assign n3608 = x134 & ~n3607 ;
  assign n3625 = n3624 ^ n3608 ;
  assign n3635 = n185 & ~n2743 ;
  assign n3634 = n136 & ~n2751 ;
  assign n3636 = n3635 ^ n3634 ;
  assign n3638 = n279 & ~n2715 ;
  assign n3637 = n254 & ~n2707 ;
  assign n3639 = n3638 ^ n3637 ;
  assign n3640 = ~n3636 & ~n3639 ;
  assign n3641 = ~x134 & n3640 ;
  assign n3627 = n185 & ~n2698 ;
  assign n3626 = n136 & ~n2690 ;
  assign n3628 = n3627 ^ n3626 ;
  assign n3630 = n279 & ~n2726 ;
  assign n3629 = n254 & ~n2734 ;
  assign n3631 = n3630 ^ n3629 ;
  assign n3632 = ~n3628 & ~n3631 ;
  assign n3633 = x134 & n3632 ;
  assign n3642 = n3641 ^ n3633 ;
  assign n3659 = n185 & ~n2865 ;
  assign n3660 = n3659 ^ n185 ;
  assign n3657 = n136 & ~n2880 ;
  assign n3658 = n3657 ^ n136 ;
  assign n3661 = n3660 ^ n3658 ;
  assign n3664 = n279 & ~n2814 ;
  assign n3665 = n3664 ^ n279 ;
  assign n3662 = n254 & ~n2800 ;
  assign n3663 = n3662 ^ n254 ;
  assign n3666 = n3665 ^ n3663 ;
  assign n3667 = n3661 & n3666 ;
  assign n3668 = n3667 ^ n3661 ;
  assign n3669 = n3668 ^ n3666 ;
  assign n3670 = x134 & ~n3669 ;
  assign n3671 = n3670 ^ n3669 ;
  assign n3645 = n185 & ~n2784 ;
  assign n3646 = n3645 ^ n185 ;
  assign n3643 = n136 & ~n2769 ;
  assign n3644 = n3643 ^ n136 ;
  assign n3647 = n3646 ^ n3644 ;
  assign n3650 = n279 & ~n2834 ;
  assign n3651 = n3650 ^ n279 ;
  assign n3648 = n254 & ~n2849 ;
  assign n3649 = n3648 ^ n254 ;
  assign n3652 = n3651 ^ n3649 ;
  assign n3653 = n3647 & n3652 ;
  assign n3654 = n3653 ^ n3647 ;
  assign n3655 = n3654 ^ n3652 ;
  assign n3656 = x134 & ~n3655 ;
  assign n3672 = n3671 ^ n3656 ;
  assign n3682 = n185 & ~n502 ;
  assign n3681 = n136 & ~n228 ;
  assign n3683 = n3682 ^ n3681 ;
  assign n3685 = ~n275 & n279 ;
  assign n3686 = ~n253 & n3685 ;
  assign n3684 = n183 & n254 ;
  assign n3687 = n3686 ^ n3684 ;
  assign n3688 = n3687 ^ x133 ;
  assign n3689 = ~n3683 & n3688 ;
  assign n3690 = ~x134 & n3689 ;
  assign n3674 = n136 & ~n413 ;
  assign n3673 = n254 & ~n369 ;
  assign n3675 = n3674 ^ n3673 ;
  assign n3677 = n185 & ~n322 ;
  assign n3676 = n279 & ~n458 ;
  assign n3678 = n3677 ^ n3676 ;
  assign n3679 = ~n3675 & ~n3678 ;
  assign n3680 = x134 & n3679 ;
  assign n3691 = n3690 ^ n3680 ;
  assign n3708 = n185 & ~n1128 ;
  assign n3709 = n3708 ^ n185 ;
  assign n3706 = n136 & ~n584 ;
  assign n3707 = n3706 ^ n136 ;
  assign n3710 = n3709 ^ n3707 ;
  assign n3713 = n279 & ~n806 ;
  assign n3714 = n3713 ^ n279 ;
  assign n3711 = n254 & ~n743 ;
  assign n3712 = n3711 ^ n254 ;
  assign n3715 = n3714 ^ n3712 ;
  assign n3716 = n3710 & n3715 ;
  assign n3717 = n3716 ^ n3710 ;
  assign n3718 = n3717 ^ n3715 ;
  assign n3719 = x134 & ~n3718 ;
  assign n3720 = n3719 ^ n3718 ;
  assign n3694 = n185 & ~n663 ;
  assign n3695 = n3694 ^ n185 ;
  assign n3692 = n136 & ~n969 ;
  assign n3693 = n3692 ^ n136 ;
  assign n3696 = n3695 ^ n3693 ;
  assign n3699 = n279 & ~n1049 ;
  assign n3700 = n3699 ^ n279 ;
  assign n3697 = n254 & ~n890 ;
  assign n3698 = n3697 ^ n254 ;
  assign n3701 = n3700 ^ n3698 ;
  assign n3702 = n3696 & n3701 ;
  assign n3703 = n3702 ^ n3696 ;
  assign n3704 = n3703 ^ n3701 ;
  assign n3705 = x134 & ~n3704 ;
  assign n3721 = n3720 ^ n3705 ;
  assign n3731 = n185 & ~n1307 ;
  assign n3730 = n136 & ~n1156 ;
  assign n3732 = n3731 ^ n3730 ;
  assign n3734 = n279 & ~n1223 ;
  assign n3733 = n254 & ~n1197 ;
  assign n3735 = n3734 ^ n3733 ;
  assign n3736 = ~n3732 & ~n3735 ;
  assign n3737 = ~x134 & n3736 ;
  assign n3723 = n185 & ~n1176 ;
  assign n3722 = n136 & ~n1266 ;
  assign n3724 = n3723 ^ n3722 ;
  assign n3726 = n279 & ~n1287 ;
  assign n3725 = n254 & ~n1246 ;
  assign n3727 = n3726 ^ n3725 ;
  assign n3728 = ~n3724 & ~n3727 ;
  assign n3729 = x134 & n3728 ;
  assign n3738 = n3737 ^ n3729 ;
  assign n3755 = n279 & ~n1363 ;
  assign n3756 = n3755 ^ n279 ;
  assign n3753 = n254 & ~n1442 ;
  assign n3754 = n3753 ^ n254 ;
  assign n3757 = n3756 ^ n3754 ;
  assign n3760 = n185 & ~n1643 ;
  assign n3761 = n3760 ^ n185 ;
  assign n3758 = n136 & ~n1481 ;
  assign n3759 = n3758 ^ n136 ;
  assign n3762 = n3761 ^ n3759 ;
  assign n3763 = n3757 & n3762 ;
  assign n3764 = n3763 ^ n3757 ;
  assign n3765 = n3764 ^ n3762 ;
  assign n3766 = x134 & ~n3765 ;
  assign n3767 = n3766 ^ n3765 ;
  assign n3741 = n185 & ~n1402 ;
  assign n3742 = n3741 ^ n185 ;
  assign n3739 = n279 & ~n1564 ;
  assign n3740 = n3739 ^ n279 ;
  assign n3743 = n3742 ^ n3740 ;
  assign n3746 = n136 & ~n1604 ;
  assign n3747 = n3746 ^ n136 ;
  assign n3744 = n254 & ~n1525 ;
  assign n3745 = n3744 ^ n254 ;
  assign n3748 = n3747 ^ n3745 ;
  assign n3749 = n3743 & n3748 ;
  assign n3750 = n3749 ^ n3743 ;
  assign n3751 = n3750 ^ n3748 ;
  assign n3752 = x134 & ~n3751 ;
  assign n3768 = n3767 ^ n3752 ;
  assign n3780 = n185 & n1721 ;
  assign n3781 = n3780 ^ x133 ;
  assign n3777 = n279 & ~n1666 ;
  assign n3778 = ~n1663 & n3777 ;
  assign n3779 = n3778 ^ x132 ;
  assign n3782 = n3781 ^ n3779 ;
  assign n3784 = n254 & ~n1685 ;
  assign n3783 = n136 & ~n1677 ;
  assign n3785 = n3784 ^ n3783 ;
  assign n3786 = n3782 & ~n3785 ;
  assign n3787 = ~x134 & n3786 ;
  assign n3770 = n136 & ~n1704 ;
  assign n3769 = n254 & ~n1696 ;
  assign n3771 = n3770 ^ n3769 ;
  assign n3773 = n279 & ~n1713 ;
  assign n3772 = n185 & ~n1659 ;
  assign n3774 = n3773 ^ n3772 ;
  assign n3775 = ~n3771 & ~n3774 ;
  assign n3776 = x134 & n3775 ;
  assign n3788 = n3787 ^ n3776 ;
  assign n3805 = n1744 ^ n279 ;
  assign n3806 = ~n279 & n3805 ;
  assign n3807 = n3806 ^ n279 ;
  assign n3808 = n3807 ^ n1749 ;
  assign n3809 = n1750 & n3808 ;
  assign n3810 = n3809 ^ n3806 ;
  assign n3811 = n3810 ^ n1749 ;
  assign n3803 = n185 & ~n1852 ;
  assign n3804 = n3803 ^ n185 ;
  assign n3812 = n3811 ^ n3804 ;
  assign n3815 = n254 & ~n1786 ;
  assign n3816 = n3815 ^ n254 ;
  assign n3813 = n136 & ~n1771 ;
  assign n3814 = n3813 ^ n136 ;
  assign n3817 = n3816 ^ n3814 ;
  assign n3818 = n3812 & n3817 ;
  assign n3819 = n3818 ^ n3812 ;
  assign n3820 = n3819 ^ n3817 ;
  assign n3821 = x134 & ~n3820 ;
  assign n3822 = n3821 ^ n3820 ;
  assign n3791 = n136 & ~n1821 ;
  assign n3792 = n3791 ^ n136 ;
  assign n3789 = n254 & ~n1806 ;
  assign n3790 = n3789 ^ n254 ;
  assign n3793 = n3792 ^ n3790 ;
  assign n3796 = n279 & ~n1837 ;
  assign n3797 = n3796 ^ n279 ;
  assign n3794 = n185 & ~n1739 ;
  assign n3795 = n3794 ^ n185 ;
  assign n3798 = n3797 ^ n3795 ;
  assign n3799 = n3793 & n3798 ;
  assign n3800 = n3799 ^ n3793 ;
  assign n3801 = n3800 ^ n3798 ;
  assign n3802 = x134 & ~n3801 ;
  assign n3823 = n3822 ^ n3802 ;
  assign n3833 = n279 & ~n1876 ;
  assign n3832 = n185 & ~n1929 ;
  assign n3834 = n3833 ^ n3832 ;
  assign n3836 = n254 & ~n1893 ;
  assign n3835 = n136 & ~n1885 ;
  assign n3837 = n3836 ^ n3835 ;
  assign n3838 = ~n3834 & ~n3837 ;
  assign n3839 = ~x134 & n3838 ;
  assign n3825 = n136 & ~n1912 ;
  assign n3824 = n254 & ~n1904 ;
  assign n3826 = n3825 ^ n3824 ;
  assign n3828 = n279 & ~n1921 ;
  assign n3827 = n185 & ~n1868 ;
  assign n3829 = n3828 ^ n3827 ;
  assign n3830 = ~n3826 & ~n3829 ;
  assign n3831 = x134 & n3830 ;
  assign n3840 = n3839 ^ n3831 ;
  assign n3857 = n279 & ~n1961 ;
  assign n3858 = n3857 ^ n279 ;
  assign n3855 = n136 & ~n1977 ;
  assign n3856 = n3855 ^ n136 ;
  assign n3859 = n3858 ^ n3856 ;
  assign n3862 = n185 & ~n2058 ;
  assign n3863 = n3862 ^ n185 ;
  assign n3860 = n254 & ~n1992 ;
  assign n3861 = n3860 ^ n254 ;
  assign n3864 = n3863 ^ n3861 ;
  assign n3865 = n3859 & n3864 ;
  assign n3866 = n3865 ^ n3859 ;
  assign n3867 = n3866 ^ n3864 ;
  assign n3868 = x134 & ~n3867 ;
  assign n3869 = n3868 ^ n3867 ;
  assign n3843 = n185 & ~n1947 ;
  assign n3844 = n3843 ^ n185 ;
  assign n3841 = n136 & ~n2027 ;
  assign n3842 = n3841 ^ n136 ;
  assign n3845 = n3844 ^ n3842 ;
  assign n3848 = n279 & ~n2043 ;
  assign n3849 = n3848 ^ n279 ;
  assign n3846 = n254 & ~n2012 ;
  assign n3847 = n3846 ^ n254 ;
  assign n3850 = n3849 ^ n3847 ;
  assign n3851 = n3845 & n3850 ;
  assign n3852 = n3851 ^ n3845 ;
  assign n3853 = n3852 ^ n3850 ;
  assign n3854 = x134 & ~n3853 ;
  assign n3870 = n3869 ^ n3854 ;
  assign n3880 = n279 & ~n2082 ;
  assign n3879 = n136 & ~n2100 ;
  assign n3881 = n3880 ^ n3879 ;
  assign n3883 = n254 & ~n2090 ;
  assign n3884 = ~n2087 & n3883 ;
  assign n3882 = n185 & n2136 ;
  assign n3885 = n3884 ^ n3882 ;
  assign n3886 = n3885 ^ x132 ;
  assign n3887 = ~n3881 & ~n3886 ;
  assign n3888 = ~x134 & n3887 ;
  assign n3872 = n185 & ~n2074 ;
  assign n3871 = n136 & ~n2119 ;
  assign n3873 = n3872 ^ n3871 ;
  assign n3875 = n279 & ~n2128 ;
  assign n3874 = n254 & ~n2111 ;
  assign n3876 = n3875 ^ n3874 ;
  assign n3877 = ~n3873 & ~n3876 ;
  assign n3878 = x134 & n3877 ;
  assign n3889 = n3888 ^ n3878 ;
  assign n3906 = n279 & ~n2168 ;
  assign n3907 = n3906 ^ n279 ;
  assign n3904 = n136 & ~n2184 ;
  assign n3905 = n3904 ^ n136 ;
  assign n3908 = n3907 ^ n3905 ;
  assign n3911 = n185 & ~n2264 ;
  assign n3912 = n3911 ^ n185 ;
  assign n3909 = n254 & ~n2198 ;
  assign n3910 = n3909 ^ n254 ;
  assign n3913 = n3912 ^ n3910 ;
  assign n3914 = n3908 & n3913 ;
  assign n3915 = n3914 ^ n3908 ;
  assign n3916 = n3915 ^ n3913 ;
  assign n3917 = x134 & ~n3916 ;
  assign n3918 = n3917 ^ n3916 ;
  assign n3892 = n185 & ~n2154 ;
  assign n3893 = n3892 ^ n185 ;
  assign n3890 = n136 & ~n2233 ;
  assign n3891 = n3890 ^ n136 ;
  assign n3894 = n3893 ^ n3891 ;
  assign n3897 = n279 & ~n2249 ;
  assign n3898 = n3897 ^ n279 ;
  assign n3895 = n254 & ~n2218 ;
  assign n3896 = n3895 ^ n254 ;
  assign n3899 = n3898 ^ n3896 ;
  assign n3900 = n3894 & n3899 ;
  assign n3901 = n3900 ^ n3894 ;
  assign n3902 = n3901 ^ n3899 ;
  assign n3903 = x134 & ~n3902 ;
  assign n3919 = n3918 ^ n3903 ;
  assign n3929 = n279 & ~n2288 ;
  assign n3928 = n185 & ~n2341 ;
  assign n3930 = n3929 ^ n3928 ;
  assign n3932 = n254 & ~n2305 ;
  assign n3931 = n136 & ~n2297 ;
  assign n3933 = n3932 ^ n3931 ;
  assign n3934 = ~n3930 & ~n3933 ;
  assign n3935 = ~x134 & n3934 ;
  assign n3921 = n185 & ~n2280 ;
  assign n3920 = n136 & ~n2324 ;
  assign n3922 = n3921 ^ n3920 ;
  assign n3924 = n279 & ~n2333 ;
  assign n3923 = n254 & ~n2316 ;
  assign n3925 = n3924 ^ n3923 ;
  assign n3926 = ~n3922 & ~n3925 ;
  assign n3927 = x134 & n3926 ;
  assign n3936 = n3935 ^ n3927 ;
  assign n3953 = n279 & ~n2373 ;
  assign n3954 = n3953 ^ n279 ;
  assign n3951 = n185 & ~n2470 ;
  assign n3952 = n3951 ^ n185 ;
  assign n3955 = n3954 ^ n3952 ;
  assign n3958 = n254 & ~n2404 ;
  assign n3959 = n3958 ^ n254 ;
  assign n3956 = n136 & ~n2389 ;
  assign n3957 = n3956 ^ n136 ;
  assign n3960 = n3959 ^ n3957 ;
  assign n3961 = n3955 & n3960 ;
  assign n3962 = n3961 ^ n3955 ;
  assign n3963 = n3962 ^ n3960 ;
  assign n3964 = x134 & ~n3963 ;
  assign n3965 = n3964 ^ n3963 ;
  assign n3939 = n185 & ~n2359 ;
  assign n3940 = n3939 ^ n185 ;
  assign n3937 = n136 & ~n2439 ;
  assign n3938 = n3937 ^ n136 ;
  assign n3941 = n3940 ^ n3938 ;
  assign n3944 = n279 & ~n2455 ;
  assign n3945 = n3944 ^ n279 ;
  assign n3942 = n254 & ~n2424 ;
  assign n3943 = n3942 ^ n254 ;
  assign n3946 = n3945 ^ n3943 ;
  assign n3947 = n3941 & n3946 ;
  assign n3948 = n3947 ^ n3941 ;
  assign n3949 = n3948 ^ n3946 ;
  assign n3950 = x134 & ~n3949 ;
  assign n3966 = n3965 ^ n3950 ;
  assign n3976 = n279 & ~n2494 ;
  assign n3975 = n185 & ~n2548 ;
  assign n3977 = n3976 ^ n3975 ;
  assign n3981 = n136 & n2512 ;
  assign n3982 = n3981 ^ x133 ;
  assign n3978 = n254 & ~n2502 ;
  assign n3979 = ~n2499 & n3978 ;
  assign n3980 = n3979 ^ x132 ;
  assign n3983 = n3982 ^ n3980 ;
  assign n3984 = ~n3977 & ~n3983 ;
  assign n3985 = ~x134 & n3984 ;
  assign n3968 = n185 & ~n2486 ;
  assign n3967 = n136 & ~n2531 ;
  assign n3969 = n3968 ^ n3967 ;
  assign n3971 = n279 & ~n2540 ;
  assign n3970 = n254 & ~n2523 ;
  assign n3972 = n3971 ^ n3970 ;
  assign n3973 = ~n3969 & ~n3972 ;
  assign n3974 = x134 & n3973 ;
  assign n3986 = n3985 ^ n3974 ;
  assign n4003 = n279 & ~n2581 ;
  assign n4004 = n4003 ^ n279 ;
  assign n4001 = n185 & ~n2674 ;
  assign n4002 = n4001 ^ n185 ;
  assign n4005 = n4004 ^ n4002 ;
  assign n4008 = n254 & ~n2607 ;
  assign n4009 = ~n2604 & n4008 ;
  assign n4010 = n4009 ^ n254 ;
  assign n4006 = n136 & ~n2597 ;
  assign n4007 = n4006 ^ n136 ;
  assign n4011 = n4010 ^ n4007 ;
  assign n4012 = n4005 & n4011 ;
  assign n4013 = n4012 ^ n4005 ;
  assign n4014 = n4013 ^ n4011 ;
  assign n4015 = x134 & ~n4014 ;
  assign n4016 = n4015 ^ n4014 ;
  assign n3989 = n185 & ~n2566 ;
  assign n3990 = n3989 ^ n185 ;
  assign n3987 = n136 & ~n2643 ;
  assign n3988 = n3987 ^ n136 ;
  assign n3991 = n3990 ^ n3988 ;
  assign n3994 = n279 & ~n2659 ;
  assign n3995 = n3994 ^ n279 ;
  assign n3992 = n254 & ~n2628 ;
  assign n3993 = n3992 ^ n254 ;
  assign n3996 = n3995 ^ n3993 ;
  assign n3997 = n3991 & n3996 ;
  assign n3998 = n3997 ^ n3991 ;
  assign n3999 = n3998 ^ n3996 ;
  assign n4000 = x134 & ~n3999 ;
  assign n4017 = n4016 ^ n4000 ;
  assign n4027 = n279 & ~n2698 ;
  assign n4026 = n185 & ~n2751 ;
  assign n4028 = n4027 ^ n4026 ;
  assign n4030 = n254 & ~n2715 ;
  assign n4029 = n136 & ~n2707 ;
  assign n4031 = n4030 ^ n4029 ;
  assign n4032 = ~n4028 & ~n4031 ;
  assign n4033 = ~x134 & n4032 ;
  assign n4019 = n185 & ~n2690 ;
  assign n4018 = n136 & ~n2734 ;
  assign n4020 = n4019 ^ n4018 ;
  assign n4022 = n279 & ~n2743 ;
  assign n4021 = n254 & ~n2726 ;
  assign n4023 = n4022 ^ n4021 ;
  assign n4024 = ~n4020 & ~n4023 ;
  assign n4025 = x134 & n4024 ;
  assign n4034 = n4033 ^ n4025 ;
  assign n4051 = n279 & ~n2784 ;
  assign n4052 = n4051 ^ n279 ;
  assign n4049 = n185 & ~n2880 ;
  assign n4050 = n4049 ^ n185 ;
  assign n4053 = n4052 ^ n4050 ;
  assign n4056 = n254 & ~n2814 ;
  assign n4057 = n4056 ^ n254 ;
  assign n4054 = n136 & ~n2800 ;
  assign n4055 = n4054 ^ n136 ;
  assign n4058 = n4057 ^ n4055 ;
  assign n4059 = n4053 & n4058 ;
  assign n4060 = n4059 ^ n4053 ;
  assign n4061 = n4060 ^ n4058 ;
  assign n4062 = x134 & ~n4061 ;
  assign n4063 = n4062 ^ n4061 ;
  assign n4037 = n185 & ~n2769 ;
  assign n4038 = n4037 ^ n185 ;
  assign n4035 = n136 & ~n2849 ;
  assign n4036 = n4035 ^ n136 ;
  assign n4039 = n4038 ^ n4036 ;
  assign n4042 = n279 & ~n2865 ;
  assign n4043 = n4042 ^ n279 ;
  assign n4040 = n254 & ~n2834 ;
  assign n4041 = n4040 ^ n254 ;
  assign n4044 = n4043 ^ n4041 ;
  assign n4045 = n4039 & n4044 ;
  assign n4046 = n4045 ^ n4039 ;
  assign n4047 = n4046 ^ n4044 ;
  assign n4048 = x134 & ~n4047 ;
  assign n4064 = n4063 ^ n4048 ;
  assign n4066 = ~x134 & n325 ;
  assign n4065 = x134 & n505 ;
  assign n4067 = n4066 ^ n4065 ;
  assign n4068 = n813 ^ n812 ;
  assign n4069 = n4068 ^ n1135 ;
  assign n4071 = ~x134 & n1226 ;
  assign n4070 = x134 & n1310 ;
  assign n4072 = n4071 ^ n4070 ;
  assign n4073 = n1488 ^ n1487 ;
  assign n4074 = n4073 ^ n1650 ;
  assign n4076 = ~x134 & n1688 ;
  assign n4075 = x134 & n1724 ;
  assign n4077 = n4076 ^ n4075 ;
  assign n4078 = n1793 ^ n1792 ;
  assign n4079 = n4078 ^ n1859 ;
  assign n4081 = ~x134 & n1896 ;
  assign n4080 = x134 & n1932 ;
  assign n4082 = n4081 ^ n4080 ;
  assign n4083 = n1999 ^ n1998 ;
  assign n4084 = n4083 ^ n2065 ;
  assign n4086 = ~x134 & n2103 ;
  assign n4085 = x134 & n2139 ;
  assign n4087 = n4086 ^ n4085 ;
  assign n4088 = n2205 ^ n2204 ;
  assign n4089 = n4088 ^ n2271 ;
  assign n4091 = ~x134 & n2308 ;
  assign n4090 = x134 & n2344 ;
  assign n4092 = n4091 ^ n4090 ;
  assign n4093 = n2411 ^ n2410 ;
  assign n4094 = n4093 ^ n2477 ;
  assign n4096 = ~x134 & n2515 ;
  assign n4095 = x134 & n2551 ;
  assign n4097 = n4096 ^ n4095 ;
  assign n4098 = n2615 ^ n2614 ;
  assign n4099 = n4098 ^ n2681 ;
  assign n4101 = ~x134 & n2718 ;
  assign n4100 = x134 & n2754 ;
  assign n4102 = n4101 ^ n4100 ;
  assign n4103 = n2821 ^ n2820 ;
  assign n4104 = n4103 ^ n2887 ;
  assign n4106 = ~x134 & n2899 ;
  assign n4105 = x134 & n2907 ;
  assign n4107 = n4106 ^ n4105 ;
  assign n4108 = n2923 ^ n2922 ;
  assign n4109 = n4108 ^ n2937 ;
  assign n4111 = ~x134 & n2946 ;
  assign n4110 = x134 & n2954 ;
  assign n4112 = n4111 ^ n4110 ;
  assign n4113 = n2970 ^ n2969 ;
  assign n4114 = n4113 ^ n2984 ;
  assign n4116 = ~x134 & n2995 ;
  assign n4115 = x134 & n3003 ;
  assign n4117 = n4116 ^ n4115 ;
  assign n4118 = n3024 ^ n3023 ;
  assign n4119 = n4118 ^ n3038 ;
  assign n4121 = ~x134 & n3047 ;
  assign n4120 = x134 & n3055 ;
  assign n4122 = n4121 ^ n4120 ;
  assign n4123 = n3071 ^ n3070 ;
  assign n4124 = n4123 ^ n3085 ;
  assign n4126 = ~x134 & n3097 ;
  assign n4125 = x134 & n3105 ;
  assign n4127 = n4126 ^ n4125 ;
  assign n4128 = n3121 ^ n3120 ;
  assign n4129 = n4128 ^ n3135 ;
  assign n4131 = ~x134 & n3144 ;
  assign n4130 = x134 & n3152 ;
  assign n4132 = n4131 ^ n4130 ;
  assign n4133 = n3168 ^ n3167 ;
  assign n4134 = n4133 ^ n3182 ;
  assign n4136 = ~x134 & n3194 ;
  assign n4135 = x134 & n3202 ;
  assign n4137 = n4136 ^ n4135 ;
  assign n4138 = n3219 ^ n3218 ;
  assign n4139 = n4138 ^ n3233 ;
  assign n4141 = ~x134 & n3242 ;
  assign n4140 = x134 & n3250 ;
  assign n4142 = n4141 ^ n4140 ;
  assign n4143 = n3266 ^ n3265 ;
  assign n4144 = n4143 ^ n3280 ;
  assign n4146 = ~x134 & n3291 ;
  assign n4145 = x134 & n3299 ;
  assign n4147 = n4146 ^ n4145 ;
  assign n4148 = n3315 ^ n3314 ;
  assign n4149 = n4148 ^ n3329 ;
  assign n4151 = ~x134 & n3338 ;
  assign n4150 = x134 & n3346 ;
  assign n4152 = n4151 ^ n4150 ;
  assign n4153 = n3362 ^ n3361 ;
  assign n4154 = n4153 ^ n3376 ;
  assign n4156 = ~x134 & n3387 ;
  assign n4155 = x134 & n3395 ;
  assign n4157 = n4156 ^ n4155 ;
  assign n4158 = n3416 ^ n3415 ;
  assign n4159 = n4158 ^ n3430 ;
  assign n4161 = ~x134 & n3439 ;
  assign n4160 = x134 & n3447 ;
  assign n4162 = n4161 ^ n4160 ;
  assign n4163 = n3463 ^ n3462 ;
  assign n4164 = n4163 ^ n3477 ;
  assign n4166 = ~x134 & n3486 ;
  assign n4165 = x134 & n3496 ;
  assign n4167 = n4166 ^ n4165 ;
  assign n4168 = n3512 ^ n3511 ;
  assign n4169 = n4168 ^ n3526 ;
  assign n4171 = ~x134 & n3535 ;
  assign n4170 = x134 & n3543 ;
  assign n4172 = n4171 ^ n4170 ;
  assign n4173 = n3559 ^ n3558 ;
  assign n4174 = n4173 ^ n3573 ;
  assign n4176 = ~x134 & n3582 ;
  assign n4175 = x134 & n3592 ;
  assign n4177 = n4176 ^ n4175 ;
  assign n4178 = n3608 ^ n3607 ;
  assign n4179 = n4178 ^ n3623 ;
  assign n4181 = ~x134 & n3632 ;
  assign n4180 = x134 & n3640 ;
  assign n4182 = n4181 ^ n4180 ;
  assign n4183 = n3656 ^ n3655 ;
  assign n4184 = n4183 ^ n3670 ;
  assign n4186 = ~x134 & n3679 ;
  assign n4185 = x134 & n3689 ;
  assign n4187 = n4186 ^ n4185 ;
  assign n4188 = n3705 ^ n3704 ;
  assign n4189 = n4188 ^ n3719 ;
  assign n4191 = ~x134 & n3728 ;
  assign n4190 = x134 & n3736 ;
  assign n4192 = n4191 ^ n4190 ;
  assign n4193 = n3752 ^ n3751 ;
  assign n4194 = n4193 ^ n3766 ;
  assign n4196 = ~x134 & n3775 ;
  assign n4195 = x134 & n3786 ;
  assign n4197 = n4196 ^ n4195 ;
  assign n4198 = n3802 ^ n3801 ;
  assign n4199 = n4198 ^ n3821 ;
  assign n4201 = ~x134 & n3830 ;
  assign n4200 = x134 & n3838 ;
  assign n4202 = n4201 ^ n4200 ;
  assign n4203 = n3854 ^ n3853 ;
  assign n4204 = n4203 ^ n3868 ;
  assign n4206 = ~x134 & n3877 ;
  assign n4205 = x134 & n3887 ;
  assign n4207 = n4206 ^ n4205 ;
  assign n4208 = n3903 ^ n3902 ;
  assign n4209 = n4208 ^ n3917 ;
  assign n4211 = ~x134 & n3926 ;
  assign n4210 = x134 & n3934 ;
  assign n4212 = n4211 ^ n4210 ;
  assign n4213 = n3950 ^ n3949 ;
  assign n4214 = n4213 ^ n3964 ;
  assign n4216 = ~x134 & n3973 ;
  assign n4215 = x134 & n3984 ;
  assign n4217 = n4216 ^ n4215 ;
  assign n4218 = n4000 ^ n3999 ;
  assign n4219 = n4218 ^ n4015 ;
  assign n4221 = ~x134 & n4024 ;
  assign n4220 = x134 & n4032 ;
  assign n4222 = n4221 ^ n4220 ;
  assign n4223 = n4048 ^ n4047 ;
  assign n4224 = n4223 ^ n4062 ;
  assign y0 = ~n507 ;
  assign y1 = n1137 ;
  assign y2 = ~n1312 ;
  assign y3 = n1652 ;
  assign y4 = ~n1726 ;
  assign y5 = n1861 ;
  assign y6 = ~n1934 ;
  assign y7 = n2067 ;
  assign y8 = ~n2141 ;
  assign y9 = n2273 ;
  assign y10 = ~n2346 ;
  assign y11 = n2479 ;
  assign y12 = ~n2553 ;
  assign y13 = n2683 ;
  assign y14 = ~n2756 ;
  assign y15 = n2889 ;
  assign y16 = ~n2909 ;
  assign y17 = n2939 ;
  assign y18 = ~n2956 ;
  assign y19 = n2986 ;
  assign y20 = ~n3005 ;
  assign y21 = n3040 ;
  assign y22 = ~n3057 ;
  assign y23 = n3087 ;
  assign y24 = ~n3107 ;
  assign y25 = n3137 ;
  assign y26 = ~n3154 ;
  assign y27 = n3184 ;
  assign y28 = ~n3204 ;
  assign y29 = n3235 ;
  assign y30 = ~n3252 ;
  assign y31 = n3282 ;
  assign y32 = ~n3301 ;
  assign y33 = n3331 ;
  assign y34 = ~n3348 ;
  assign y35 = n3378 ;
  assign y36 = ~n3397 ;
  assign y37 = n3432 ;
  assign y38 = ~n3449 ;
  assign y39 = n3479 ;
  assign y40 = ~n3498 ;
  assign y41 = n3528 ;
  assign y42 = ~n3545 ;
  assign y43 = n3575 ;
  assign y44 = ~n3594 ;
  assign y45 = n3625 ;
  assign y46 = ~n3642 ;
  assign y47 = n3672 ;
  assign y48 = ~n3691 ;
  assign y49 = n3721 ;
  assign y50 = ~n3738 ;
  assign y51 = n3768 ;
  assign y52 = ~n3788 ;
  assign y53 = n3823 ;
  assign y54 = ~n3840 ;
  assign y55 = n3870 ;
  assign y56 = ~n3889 ;
  assign y57 = n3919 ;
  assign y58 = ~n3936 ;
  assign y59 = n3966 ;
  assign y60 = ~n3986 ;
  assign y61 = n4017 ;
  assign y62 = ~n4034 ;
  assign y63 = n4064 ;
  assign y64 = ~n4067 ;
  assign y65 = n4069 ;
  assign y66 = ~n4072 ;
  assign y67 = n4074 ;
  assign y68 = ~n4077 ;
  assign y69 = n4079 ;
  assign y70 = ~n4082 ;
  assign y71 = n4084 ;
  assign y72 = ~n4087 ;
  assign y73 = n4089 ;
  assign y74 = ~n4092 ;
  assign y75 = n4094 ;
  assign y76 = ~n4097 ;
  assign y77 = n4099 ;
  assign y78 = ~n4102 ;
  assign y79 = n4104 ;
  assign y80 = ~n4107 ;
  assign y81 = n4109 ;
  assign y82 = ~n4112 ;
  assign y83 = n4114 ;
  assign y84 = ~n4117 ;
  assign y85 = n4119 ;
  assign y86 = ~n4122 ;
  assign y87 = n4124 ;
  assign y88 = ~n4127 ;
  assign y89 = n4129 ;
  assign y90 = ~n4132 ;
  assign y91 = n4134 ;
  assign y92 = ~n4137 ;
  assign y93 = n4139 ;
  assign y94 = ~n4142 ;
  assign y95 = n4144 ;
  assign y96 = ~n4147 ;
  assign y97 = n4149 ;
  assign y98 = ~n4152 ;
  assign y99 = n4154 ;
  assign y100 = ~n4157 ;
  assign y101 = n4159 ;
  assign y102 = ~n4162 ;
  assign y103 = n4164 ;
  assign y104 = ~n4167 ;
  assign y105 = n4169 ;
  assign y106 = ~n4172 ;
  assign y107 = n4174 ;
  assign y108 = ~n4177 ;
  assign y109 = n4179 ;
  assign y110 = ~n4182 ;
  assign y111 = n4184 ;
  assign y112 = ~n4187 ;
  assign y113 = n4189 ;
  assign y114 = ~n4192 ;
  assign y115 = n4194 ;
  assign y116 = ~n4197 ;
  assign y117 = n4199 ;
  assign y118 = ~n4202 ;
  assign y119 = n4204 ;
  assign y120 = ~n4207 ;
  assign y121 = n4209 ;
  assign y122 = ~n4212 ;
  assign y123 = n4214 ;
  assign y124 = ~n4217 ;
  assign y125 = n4219 ;
  assign y126 = ~n4222 ;
  assign y127 = n4224 ;
endmodule
