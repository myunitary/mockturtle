// eight parties, each holding 16-bit data
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 ;
  assign n132 = ~x79 & ~x95 ;
  assign n133 = ~x111 & ~x127 ;
  assign n134 = n132 & n133 ;
  assign n129 = ~x15 & ~x31 ;
  assign n130 = ~x47 & ~x63 ;
  assign n131 = n129 & n130 ;
  assign n135 = n134 ^ n131 ;
  assign n467 = x94 ^ x78 ;
  assign n468 = x95 ^ x79 ;
  assign n525 = x94 ^ x77 ;
  assign n469 = x92 ^ x76 ;
  assign n517 = x92 ^ x75 ;
  assign n470 = x90 ^ x74 ;
  assign n509 = x90 ^ x73 ;
  assign n471 = x88 ^ x72 ;
  assign n501 = x88 ^ x71 ;
  assign n472 = x86 ^ x70 ;
  assign n493 = x86 ^ x69 ;
  assign n473 = x84 ^ x68 ;
  assign n485 = x84 ^ x67 ;
  assign n474 = x82 ^ x66 ;
  assign n477 = x82 ^ x65 ;
  assign n475 = x64 & ~x80 ;
  assign n476 = n475 ^ x82 ;
  assign n478 = n477 ^ n476 ;
  assign n479 = x81 ^ x65 ;
  assign n480 = n478 & ~n479 ;
  assign n481 = n480 ^ n477 ;
  assign n482 = ~n474 & n481 ;
  assign n483 = n482 ^ x66 ;
  assign n484 = n483 ^ x84 ;
  assign n486 = n485 ^ n484 ;
  assign n487 = x83 ^ x67 ;
  assign n488 = n486 & ~n487 ;
  assign n489 = n488 ^ n485 ;
  assign n490 = ~n473 & n489 ;
  assign n491 = n490 ^ x68 ;
  assign n492 = n491 ^ x86 ;
  assign n494 = n493 ^ n492 ;
  assign n495 = x85 ^ x69 ;
  assign n496 = n494 & ~n495 ;
  assign n497 = n496 ^ n493 ;
  assign n498 = ~n472 & n497 ;
  assign n499 = n498 ^ x70 ;
  assign n500 = n499 ^ x88 ;
  assign n502 = n501 ^ n500 ;
  assign n503 = x87 ^ x71 ;
  assign n504 = n502 & ~n503 ;
  assign n505 = n504 ^ n501 ;
  assign n506 = ~n471 & n505 ;
  assign n507 = n506 ^ x72 ;
  assign n508 = n507 ^ x90 ;
  assign n510 = n509 ^ n508 ;
  assign n511 = x89 ^ x73 ;
  assign n512 = n510 & ~n511 ;
  assign n513 = n512 ^ n509 ;
  assign n514 = ~n470 & n513 ;
  assign n515 = n514 ^ x74 ;
  assign n516 = n515 ^ x92 ;
  assign n518 = n517 ^ n516 ;
  assign n519 = x91 ^ x75 ;
  assign n520 = n518 & ~n519 ;
  assign n521 = n520 ^ n517 ;
  assign n522 = ~n469 & n521 ;
  assign n523 = n522 ^ x76 ;
  assign n524 = n523 ^ x94 ;
  assign n526 = n525 ^ n524 ;
  assign n527 = x93 ^ x77 ;
  assign n528 = n526 & ~n527 ;
  assign n529 = n528 ^ n525 ;
  assign n530 = ~n467 & n529 ;
  assign n531 = n530 ^ x78 ;
  assign n532 = n531 ^ x95 ;
  assign n533 = ~n468 & n532 ;
  assign n534 = n533 ^ x79 ;
  assign n535 = n467 & ~n534 ;
  assign n536 = n535 ^ x78 ;
  assign n397 = x126 ^ x110 ;
  assign n398 = x127 ^ x111 ;
  assign n455 = x126 ^ x109 ;
  assign n399 = x124 ^ x108 ;
  assign n447 = x124 ^ x107 ;
  assign n400 = x122 ^ x106 ;
  assign n439 = x122 ^ x105 ;
  assign n401 = x120 ^ x104 ;
  assign n431 = x120 ^ x103 ;
  assign n402 = x118 ^ x102 ;
  assign n423 = x118 ^ x101 ;
  assign n403 = x116 ^ x100 ;
  assign n415 = x116 ^ x99 ;
  assign n404 = x114 ^ x98 ;
  assign n407 = x114 ^ x97 ;
  assign n405 = x96 & ~x112 ;
  assign n406 = n405 ^ x114 ;
  assign n408 = n407 ^ n406 ;
  assign n409 = x113 ^ x97 ;
  assign n410 = n408 & ~n409 ;
  assign n411 = n410 ^ n407 ;
  assign n412 = ~n404 & n411 ;
  assign n413 = n412 ^ x98 ;
  assign n414 = n413 ^ x116 ;
  assign n416 = n415 ^ n414 ;
  assign n417 = x115 ^ x99 ;
  assign n418 = n416 & ~n417 ;
  assign n419 = n418 ^ n415 ;
  assign n420 = ~n403 & n419 ;
  assign n421 = n420 ^ x100 ;
  assign n422 = n421 ^ x118 ;
  assign n424 = n423 ^ n422 ;
  assign n425 = x117 ^ x101 ;
  assign n426 = n424 & ~n425 ;
  assign n427 = n426 ^ n423 ;
  assign n428 = ~n402 & n427 ;
  assign n429 = n428 ^ x102 ;
  assign n430 = n429 ^ x120 ;
  assign n432 = n431 ^ n430 ;
  assign n433 = x119 ^ x103 ;
  assign n434 = n432 & ~n433 ;
  assign n435 = n434 ^ n431 ;
  assign n436 = ~n401 & n435 ;
  assign n437 = n436 ^ x104 ;
  assign n438 = n437 ^ x122 ;
  assign n440 = n439 ^ n438 ;
  assign n441 = x121 ^ x105 ;
  assign n442 = n440 & ~n441 ;
  assign n443 = n442 ^ n439 ;
  assign n444 = ~n400 & n443 ;
  assign n445 = n444 ^ x106 ;
  assign n446 = n445 ^ x124 ;
  assign n448 = n447 ^ n446 ;
  assign n449 = x123 ^ x107 ;
  assign n450 = n448 & ~n449 ;
  assign n451 = n450 ^ n447 ;
  assign n452 = ~n399 & n451 ;
  assign n453 = n452 ^ x108 ;
  assign n454 = n453 ^ x126 ;
  assign n456 = n455 ^ n454 ;
  assign n457 = x125 ^ x109 ;
  assign n458 = n456 & ~n457 ;
  assign n459 = n458 ^ n455 ;
  assign n460 = ~n397 & n459 ;
  assign n461 = n460 ^ x110 ;
  assign n462 = n461 ^ x127 ;
  assign n463 = ~n398 & n462 ;
  assign n464 = n463 ^ x111 ;
  assign n465 = n397 & ~n464 ;
  assign n466 = n465 ^ x110 ;
  assign n537 = n536 ^ n466 ;
  assign n538 = n133 ^ n132 ;
  assign n541 = n457 & ~n464 ;
  assign n542 = n541 ^ x109 ;
  assign n539 = n527 & ~n534 ;
  assign n540 = n539 ^ x77 ;
  assign n543 = n542 ^ n540 ;
  assign n546 = n399 & ~n464 ;
  assign n547 = n546 ^ x108 ;
  assign n544 = n469 & ~n534 ;
  assign n545 = n544 ^ x76 ;
  assign n548 = n547 ^ n545 ;
  assign n551 = n519 & ~n534 ;
  assign n552 = n551 ^ x75 ;
  assign n549 = n449 & ~n464 ;
  assign n550 = n549 ^ x107 ;
  assign n553 = n552 ^ n550 ;
  assign n556 = n470 & ~n534 ;
  assign n557 = n556 ^ x74 ;
  assign n554 = n400 & ~n464 ;
  assign n555 = n554 ^ x106 ;
  assign n558 = n557 ^ n555 ;
  assign n561 = n441 & ~n464 ;
  assign n562 = n561 ^ x105 ;
  assign n559 = n511 & ~n534 ;
  assign n560 = n559 ^ x73 ;
  assign n563 = n562 ^ n560 ;
  assign n566 = n471 & ~n534 ;
  assign n567 = n566 ^ x72 ;
  assign n564 = n401 & ~n464 ;
  assign n565 = n564 ^ x104 ;
  assign n568 = n567 ^ n565 ;
  assign n571 = n433 & ~n464 ;
  assign n572 = n571 ^ x103 ;
  assign n569 = n503 & ~n534 ;
  assign n570 = n569 ^ x71 ;
  assign n573 = n572 ^ n570 ;
  assign n576 = n402 & ~n464 ;
  assign n577 = n576 ^ x102 ;
  assign n574 = n472 & ~n534 ;
  assign n575 = n574 ^ x70 ;
  assign n578 = n577 ^ n575 ;
  assign n581 = n425 & ~n464 ;
  assign n582 = n581 ^ x101 ;
  assign n579 = n495 & ~n534 ;
  assign n580 = n579 ^ x69 ;
  assign n583 = n582 ^ n580 ;
  assign n586 = n403 & ~n464 ;
  assign n587 = n586 ^ x100 ;
  assign n584 = n473 & ~n534 ;
  assign n585 = n584 ^ x68 ;
  assign n588 = n587 ^ n585 ;
  assign n591 = n487 & ~n534 ;
  assign n592 = n591 ^ x67 ;
  assign n589 = n417 & ~n464 ;
  assign n590 = n589 ^ x99 ;
  assign n593 = n592 ^ n590 ;
  assign n596 = n404 & ~n464 ;
  assign n597 = n596 ^ x98 ;
  assign n594 = n474 & ~n534 ;
  assign n595 = n594 ^ x66 ;
  assign n598 = n597 ^ n595 ;
  assign n601 = n479 & ~n534 ;
  assign n602 = n601 ^ x65 ;
  assign n599 = n409 & ~n464 ;
  assign n600 = n599 ^ x97 ;
  assign n603 = n602 ^ n600 ;
  assign n604 = x112 ^ x96 ;
  assign n605 = ~n464 & n604 ;
  assign n606 = n605 ^ x96 ;
  assign n607 = x80 ^ x64 ;
  assign n608 = ~n534 & n607 ;
  assign n609 = n608 ^ x64 ;
  assign n610 = ~n606 & n609 ;
  assign n611 = n610 ^ n600 ;
  assign n612 = ~n603 & ~n611 ;
  assign n613 = n612 ^ n600 ;
  assign n614 = n613 ^ n597 ;
  assign n615 = ~n598 & n614 ;
  assign n616 = n615 ^ n597 ;
  assign n617 = n616 ^ n590 ;
  assign n618 = ~n593 & n617 ;
  assign n619 = n618 ^ n590 ;
  assign n620 = n619 ^ n587 ;
  assign n621 = ~n588 & n620 ;
  assign n622 = n621 ^ n587 ;
  assign n623 = n622 ^ n580 ;
  assign n624 = ~n583 & ~n623 ;
  assign n625 = n624 ^ n580 ;
  assign n626 = n625 ^ n577 ;
  assign n627 = ~n578 & ~n626 ;
  assign n628 = n627 ^ n577 ;
  assign n629 = n628 ^ n570 ;
  assign n630 = ~n573 & ~n629 ;
  assign n631 = n630 ^ n570 ;
  assign n632 = n631 ^ n567 ;
  assign n633 = ~n568 & n632 ;
  assign n634 = n633 ^ n567 ;
  assign n635 = n634 ^ n560 ;
  assign n636 = ~n563 & n635 ;
  assign n637 = n636 ^ n560 ;
  assign n638 = n637 ^ n557 ;
  assign n639 = ~n558 & n638 ;
  assign n640 = n639 ^ n557 ;
  assign n641 = n640 ^ n550 ;
  assign n642 = ~n553 & ~n641 ;
  assign n643 = n642 ^ n550 ;
  assign n644 = n643 ^ n545 ;
  assign n645 = ~n548 & ~n644 ;
  assign n646 = n645 ^ n545 ;
  assign n647 = n646 ^ n540 ;
  assign n648 = ~n543 & ~n647 ;
  assign n649 = n648 ^ n542 ;
  assign n650 = n649 ^ n466 ;
  assign n651 = ~n537 & ~n650 ;
  assign n652 = n651 ^ n536 ;
  assign n653 = n652 ^ n133 ;
  assign n654 = ~n538 & ~n653 ;
  assign n655 = n654 ^ n132 ;
  assign n656 = n537 & n655 ;
  assign n657 = n656 ^ n536 ;
  assign n206 = x62 ^ x46 ;
  assign n207 = x63 ^ x47 ;
  assign n264 = x62 ^ x45 ;
  assign n208 = x60 ^ x44 ;
  assign n256 = x60 ^ x43 ;
  assign n209 = x58 ^ x42 ;
  assign n248 = x58 ^ x41 ;
  assign n210 = x56 ^ x40 ;
  assign n240 = x56 ^ x39 ;
  assign n211 = x54 ^ x38 ;
  assign n232 = x54 ^ x37 ;
  assign n212 = x52 ^ x36 ;
  assign n224 = x52 ^ x35 ;
  assign n213 = x50 ^ x34 ;
  assign n216 = x50 ^ x33 ;
  assign n214 = x32 & ~x48 ;
  assign n215 = n214 ^ x50 ;
  assign n217 = n216 ^ n215 ;
  assign n218 = x49 ^ x33 ;
  assign n219 = n217 & ~n218 ;
  assign n220 = n219 ^ n216 ;
  assign n221 = ~n213 & n220 ;
  assign n222 = n221 ^ x34 ;
  assign n223 = n222 ^ x52 ;
  assign n225 = n224 ^ n223 ;
  assign n226 = x51 ^ x35 ;
  assign n227 = n225 & ~n226 ;
  assign n228 = n227 ^ n224 ;
  assign n229 = ~n212 & n228 ;
  assign n230 = n229 ^ x36 ;
  assign n231 = n230 ^ x54 ;
  assign n233 = n232 ^ n231 ;
  assign n234 = x53 ^ x37 ;
  assign n235 = n233 & ~n234 ;
  assign n236 = n235 ^ n232 ;
  assign n237 = ~n211 & n236 ;
  assign n238 = n237 ^ x38 ;
  assign n239 = n238 ^ x56 ;
  assign n241 = n240 ^ n239 ;
  assign n242 = x55 ^ x39 ;
  assign n243 = n241 & ~n242 ;
  assign n244 = n243 ^ n240 ;
  assign n245 = ~n210 & n244 ;
  assign n246 = n245 ^ x40 ;
  assign n247 = n246 ^ x58 ;
  assign n249 = n248 ^ n247 ;
  assign n250 = x57 ^ x41 ;
  assign n251 = n249 & ~n250 ;
  assign n252 = n251 ^ n248 ;
  assign n253 = ~n209 & n252 ;
  assign n254 = n253 ^ x42 ;
  assign n255 = n254 ^ x60 ;
  assign n257 = n256 ^ n255 ;
  assign n258 = x59 ^ x43 ;
  assign n259 = n257 & ~n258 ;
  assign n260 = n259 ^ n256 ;
  assign n261 = ~n208 & n260 ;
  assign n262 = n261 ^ x44 ;
  assign n263 = n262 ^ x62 ;
  assign n265 = n264 ^ n263 ;
  assign n266 = x61 ^ x45 ;
  assign n267 = n265 & ~n266 ;
  assign n268 = n267 ^ n264 ;
  assign n269 = ~n206 & n268 ;
  assign n270 = n269 ^ x46 ;
  assign n271 = n270 ^ x63 ;
  assign n272 = ~n207 & n271 ;
  assign n273 = n272 ^ x47 ;
  assign n274 = n206 & ~n273 ;
  assign n275 = n274 ^ x46 ;
  assign n136 = x30 ^ x14 ;
  assign n137 = x31 ^ x15 ;
  assign n194 = x30 ^ x13 ;
  assign n138 = x28 ^ x12 ;
  assign n186 = x28 ^ x11 ;
  assign n139 = x26 ^ x10 ;
  assign n178 = x26 ^ x9 ;
  assign n140 = x24 ^ x8 ;
  assign n170 = x24 ^ x7 ;
  assign n141 = x22 ^ x6 ;
  assign n162 = x22 ^ x5 ;
  assign n142 = x20 ^ x4 ;
  assign n154 = x20 ^ x3 ;
  assign n143 = x18 ^ x2 ;
  assign n146 = x18 ^ x1 ;
  assign n144 = x0 & ~x16 ;
  assign n145 = n144 ^ x18 ;
  assign n147 = n146 ^ n145 ;
  assign n148 = x17 ^ x1 ;
  assign n149 = n147 & ~n148 ;
  assign n150 = n149 ^ n146 ;
  assign n151 = ~n143 & n150 ;
  assign n152 = n151 ^ x2 ;
  assign n153 = n152 ^ x20 ;
  assign n155 = n154 ^ n153 ;
  assign n156 = x19 ^ x3 ;
  assign n157 = n155 & ~n156 ;
  assign n158 = n157 ^ n154 ;
  assign n159 = ~n142 & n158 ;
  assign n160 = n159 ^ x4 ;
  assign n161 = n160 ^ x22 ;
  assign n163 = n162 ^ n161 ;
  assign n164 = x21 ^ x5 ;
  assign n165 = n163 & ~n164 ;
  assign n166 = n165 ^ n162 ;
  assign n167 = ~n141 & n166 ;
  assign n168 = n167 ^ x6 ;
  assign n169 = n168 ^ x24 ;
  assign n171 = n170 ^ n169 ;
  assign n172 = x23 ^ x7 ;
  assign n173 = n171 & ~n172 ;
  assign n174 = n173 ^ n170 ;
  assign n175 = ~n140 & n174 ;
  assign n176 = n175 ^ x8 ;
  assign n177 = n176 ^ x26 ;
  assign n179 = n178 ^ n177 ;
  assign n180 = x25 ^ x9 ;
  assign n181 = n179 & ~n180 ;
  assign n182 = n181 ^ n178 ;
  assign n183 = ~n139 & n182 ;
  assign n184 = n183 ^ x10 ;
  assign n185 = n184 ^ x28 ;
  assign n187 = n186 ^ n185 ;
  assign n188 = x27 ^ x11 ;
  assign n189 = n187 & ~n188 ;
  assign n190 = n189 ^ n186 ;
  assign n191 = ~n138 & n190 ;
  assign n192 = n191 ^ x12 ;
  assign n193 = n192 ^ x30 ;
  assign n195 = n194 ^ n193 ;
  assign n196 = x29 ^ x13 ;
  assign n197 = n195 & ~n196 ;
  assign n198 = n197 ^ n194 ;
  assign n199 = ~n136 & n198 ;
  assign n200 = n199 ^ x14 ;
  assign n201 = n200 ^ x31 ;
  assign n202 = ~n137 & n201 ;
  assign n203 = n202 ^ x15 ;
  assign n204 = n136 & ~n203 ;
  assign n205 = n204 ^ x14 ;
  assign n276 = n275 ^ n205 ;
  assign n277 = n130 ^ n129 ;
  assign n280 = n266 & ~n273 ;
  assign n281 = n280 ^ x45 ;
  assign n278 = n196 & ~n203 ;
  assign n279 = n278 ^ x13 ;
  assign n282 = n281 ^ n279 ;
  assign n285 = n138 & ~n203 ;
  assign n286 = n285 ^ x12 ;
  assign n283 = n208 & ~n273 ;
  assign n284 = n283 ^ x44 ;
  assign n287 = n286 ^ n284 ;
  assign n290 = n258 & ~n273 ;
  assign n291 = n290 ^ x43 ;
  assign n288 = n188 & ~n203 ;
  assign n289 = n288 ^ x11 ;
  assign n292 = n291 ^ n289 ;
  assign n295 = n139 & ~n203 ;
  assign n296 = n295 ^ x10 ;
  assign n293 = n209 & ~n273 ;
  assign n294 = n293 ^ x42 ;
  assign n297 = n296 ^ n294 ;
  assign n300 = n250 & ~n273 ;
  assign n301 = n300 ^ x41 ;
  assign n298 = n180 & ~n203 ;
  assign n299 = n298 ^ x9 ;
  assign n302 = n301 ^ n299 ;
  assign n305 = n210 & ~n273 ;
  assign n306 = n305 ^ x40 ;
  assign n303 = n140 & ~n203 ;
  assign n304 = n303 ^ x8 ;
  assign n307 = n306 ^ n304 ;
  assign n310 = n242 & ~n273 ;
  assign n311 = n310 ^ x39 ;
  assign n308 = n172 & ~n203 ;
  assign n309 = n308 ^ x7 ;
  assign n312 = n311 ^ n309 ;
  assign n315 = n141 & ~n203 ;
  assign n316 = n315 ^ x6 ;
  assign n313 = n211 & ~n273 ;
  assign n314 = n313 ^ x38 ;
  assign n317 = n316 ^ n314 ;
  assign n320 = n234 & ~n273 ;
  assign n321 = n320 ^ x37 ;
  assign n318 = n164 & ~n203 ;
  assign n319 = n318 ^ x5 ;
  assign n322 = n321 ^ n319 ;
  assign n325 = n142 & ~n203 ;
  assign n326 = n325 ^ x4 ;
  assign n323 = n212 & ~n273 ;
  assign n324 = n323 ^ x36 ;
  assign n327 = n326 ^ n324 ;
  assign n330 = n226 & ~n273 ;
  assign n331 = n330 ^ x35 ;
  assign n328 = n156 & ~n203 ;
  assign n329 = n328 ^ x3 ;
  assign n332 = n331 ^ n329 ;
  assign n335 = n213 & ~n273 ;
  assign n336 = n335 ^ x34 ;
  assign n333 = n143 & ~n203 ;
  assign n334 = n333 ^ x2 ;
  assign n337 = n336 ^ n334 ;
  assign n340 = n148 & ~n203 ;
  assign n341 = n340 ^ x1 ;
  assign n338 = n218 & ~n273 ;
  assign n339 = n338 ^ x33 ;
  assign n342 = n341 ^ n339 ;
  assign n343 = x48 ^ x32 ;
  assign n344 = ~n273 & n343 ;
  assign n345 = n344 ^ x32 ;
  assign n346 = x16 ^ x0 ;
  assign n347 = ~n203 & n346 ;
  assign n348 = n347 ^ x0 ;
  assign n349 = ~n345 & n348 ;
  assign n350 = n349 ^ n339 ;
  assign n351 = ~n342 & ~n350 ;
  assign n352 = n351 ^ n339 ;
  assign n353 = n352 ^ n334 ;
  assign n354 = ~n337 & ~n353 ;
  assign n355 = n354 ^ n334 ;
  assign n356 = n355 ^ n329 ;
  assign n357 = ~n332 & n356 ;
  assign n358 = n357 ^ n329 ;
  assign n359 = n358 ^ n326 ;
  assign n360 = ~n327 & n359 ;
  assign n361 = n360 ^ n326 ;
  assign n362 = n361 ^ n319 ;
  assign n363 = ~n322 & n362 ;
  assign n364 = n363 ^ n319 ;
  assign n365 = n364 ^ n316 ;
  assign n366 = ~n317 & n365 ;
  assign n367 = n366 ^ n316 ;
  assign n368 = n367 ^ n309 ;
  assign n369 = ~n312 & n368 ;
  assign n370 = n369 ^ n309 ;
  assign n371 = n370 ^ n306 ;
  assign n372 = ~n307 & ~n371 ;
  assign n373 = n372 ^ n306 ;
  assign n374 = n373 ^ n299 ;
  assign n375 = ~n302 & ~n374 ;
  assign n376 = n375 ^ n299 ;
  assign n377 = n376 ^ n296 ;
  assign n378 = ~n297 & n377 ;
  assign n379 = n378 ^ n296 ;
  assign n380 = n379 ^ n289 ;
  assign n381 = ~n292 & n380 ;
  assign n382 = n381 ^ n289 ;
  assign n383 = n382 ^ n284 ;
  assign n384 = ~n287 & ~n383 ;
  assign n385 = n384 ^ n284 ;
  assign n386 = n385 ^ n279 ;
  assign n387 = ~n282 & n386 ;
  assign n388 = n387 ^ n281 ;
  assign n389 = n388 ^ n205 ;
  assign n390 = ~n276 & n389 ;
  assign n391 = n390 ^ n275 ;
  assign n392 = n391 ^ n130 ;
  assign n393 = ~n277 & n392 ;
  assign n394 = n393 ^ n129 ;
  assign n395 = n276 & ~n394 ;
  assign n396 = n395 ^ n275 ;
  assign n658 = n657 ^ n396 ;
  assign n661 = n543 & n655 ;
  assign n662 = n661 ^ n540 ;
  assign n659 = n282 & n394 ;
  assign n660 = n659 ^ n279 ;
  assign n663 = n662 ^ n660 ;
  assign n666 = n287 & ~n394 ;
  assign n667 = n666 ^ n284 ;
  assign n664 = n548 & n655 ;
  assign n665 = n664 ^ n545 ;
  assign n668 = n667 ^ n665 ;
  assign n671 = n553 & ~n655 ;
  assign n672 = n671 ^ n550 ;
  assign n669 = n292 & n394 ;
  assign n670 = n669 ^ n289 ;
  assign n673 = n672 ^ n670 ;
  assign n676 = n558 & n655 ;
  assign n677 = n676 ^ n557 ;
  assign n674 = n297 & n394 ;
  assign n675 = n674 ^ n296 ;
  assign n678 = n677 ^ n675 ;
  assign n681 = n302 & ~n394 ;
  assign n682 = n681 ^ n301 ;
  assign n679 = n563 & ~n655 ;
  assign n680 = n679 ^ n562 ;
  assign n683 = n682 ^ n680 ;
  assign n686 = n568 & ~n655 ;
  assign n687 = n686 ^ n565 ;
  assign n684 = n307 & n394 ;
  assign n685 = n684 ^ n304 ;
  assign n688 = n687 ^ n685 ;
  assign n691 = n573 & n655 ;
  assign n692 = n691 ^ n570 ;
  assign n689 = n312 & n394 ;
  assign n690 = n689 ^ n309 ;
  assign n693 = n692 ^ n690 ;
  assign n696 = n317 & n394 ;
  assign n697 = n696 ^ n316 ;
  assign n694 = n578 & ~n655 ;
  assign n695 = n694 ^ n577 ;
  assign n698 = n697 ^ n695 ;
  assign n701 = n322 & ~n394 ;
  assign n702 = n701 ^ n321 ;
  assign n699 = n583 & ~n655 ;
  assign n700 = n699 ^ n582 ;
  assign n703 = n702 ^ n700 ;
  assign n706 = n327 & ~n394 ;
  assign n707 = n706 ^ n324 ;
  assign n704 = n588 & n655 ;
  assign n705 = n704 ^ n585 ;
  assign n708 = n707 ^ n705 ;
  assign n711 = n593 & ~n655 ;
  assign n712 = n711 ^ n590 ;
  assign n709 = n332 & n394 ;
  assign n710 = n709 ^ n329 ;
  assign n713 = n712 ^ n710 ;
  assign n716 = n598 & ~n655 ;
  assign n717 = n716 ^ n597 ;
  assign n714 = n337 & ~n394 ;
  assign n715 = n714 ^ n336 ;
  assign n718 = n717 ^ n715 ;
  assign n721 = n342 & n394 ;
  assign n722 = n721 ^ n341 ;
  assign n719 = n603 & n655 ;
  assign n720 = n719 ^ n602 ;
  assign n723 = n722 ^ n720 ;
  assign n724 = n609 ^ n606 ;
  assign n725 = ~n655 & n724 ;
  assign n726 = n725 ^ n606 ;
  assign n727 = n348 ^ n345 ;
  assign n728 = ~n394 & n727 ;
  assign n729 = n728 ^ n345 ;
  assign n730 = ~n726 & n729 ;
  assign n731 = n730 ^ n720 ;
  assign n732 = ~n723 & ~n731 ;
  assign n733 = n732 ^ n720 ;
  assign n734 = n733 ^ n717 ;
  assign n735 = ~n718 & n734 ;
  assign n736 = n735 ^ n717 ;
  assign n737 = n736 ^ n710 ;
  assign n738 = ~n713 & ~n737 ;
  assign n739 = n738 ^ n710 ;
  assign n740 = n739 ^ n707 ;
  assign n741 = ~n708 & n740 ;
  assign n742 = n741 ^ n707 ;
  assign n743 = n742 ^ n700 ;
  assign n744 = ~n703 & ~n743 ;
  assign n745 = n744 ^ n700 ;
  assign n746 = n745 ^ n697 ;
  assign n747 = ~n698 & ~n746 ;
  assign n748 = n747 ^ n697 ;
  assign n749 = n748 ^ n690 ;
  assign n750 = ~n693 & n749 ;
  assign n751 = n750 ^ n690 ;
  assign n752 = n751 ^ n687 ;
  assign n753 = ~n688 & ~n752 ;
  assign n754 = n753 ^ n687 ;
  assign n755 = n754 ^ n680 ;
  assign n756 = ~n683 & n755 ;
  assign n757 = n756 ^ n680 ;
  assign n758 = n757 ^ n677 ;
  assign n759 = ~n678 & n758 ;
  assign n760 = n759 ^ n677 ;
  assign n761 = n760 ^ n670 ;
  assign n762 = ~n673 & ~n761 ;
  assign n763 = n762 ^ n670 ;
  assign n764 = n763 ^ n667 ;
  assign n765 = ~n668 & n764 ;
  assign n766 = n765 ^ n667 ;
  assign n767 = n766 ^ n662 ;
  assign n768 = ~n663 & ~n767 ;
  assign n769 = n768 ^ n662 ;
  assign n770 = n769 ^ n657 ;
  assign n771 = ~n658 & ~n770 ;
  assign n772 = n771 ^ n396 ;
  assign n773 = n772 ^ n131 ;
  assign n774 = ~n135 & n773 ;
  assign n775 = n774 ^ n134 ;
  assign n776 = n655 ^ n394 ;
  assign n777 = ~n775 & n776 ;
  assign n778 = n777 ^ n394 ;
  assign n782 = n534 & ~n778 ;
  assign n783 = n464 & n655 ;
  assign n784 = ~n782 & ~n783 ;
  assign n779 = n203 & ~n778 ;
  assign n780 = n273 & n394 ;
  assign n781 = ~n779 & ~n780 ;
  assign n785 = n784 ^ n781 ;
  assign n786 = n775 & n785 ;
  assign n787 = n786 ^ n784 ;
  assign n788 = n729 ^ n726 ;
  assign n789 = n775 & n788 ;
  assign n790 = n789 ^ n726 ;
  assign n791 = n723 & ~n775 ;
  assign n792 = n791 ^ n722 ;
  assign n793 = n718 & n775 ;
  assign n794 = n793 ^ n717 ;
  assign n795 = n713 & ~n775 ;
  assign n796 = n795 ^ n710 ;
  assign n797 = n708 & n775 ;
  assign n798 = n797 ^ n705 ;
  assign n799 = n703 & ~n775 ;
  assign n800 = n799 ^ n702 ;
  assign n801 = n698 & ~n775 ;
  assign n802 = n801 ^ n697 ;
  assign n803 = n693 & ~n775 ;
  assign n804 = n803 ^ n690 ;
  assign n805 = n688 & ~n775 ;
  assign n806 = n805 ^ n685 ;
  assign n807 = n683 & ~n775 ;
  assign n808 = n807 ^ n682 ;
  assign n809 = n678 & n775 ;
  assign n810 = n809 ^ n677 ;
  assign n811 = n673 & ~n775 ;
  assign n812 = n811 ^ n670 ;
  assign n813 = n668 & n775 ;
  assign n814 = n813 ^ n665 ;
  assign n815 = n663 & n775 ;
  assign n816 = n815 ^ n662 ;
  assign n817 = n658 & n775 ;
  assign n818 = n817 ^ n657 ;
  assign n819 = n131 & n134 ;
  assign y0 = n787 ;
  assign y1 = n778 ;
  assign y2 = ~n775 ;
  assign y3 = n790 ;
  assign y4 = n792 ;
  assign y5 = n794 ;
  assign y6 = n796 ;
  assign y7 = n798 ;
  assign y8 = n800 ;
  assign y9 = n802 ;
  assign y10 = n804 ;
  assign y11 = n806 ;
  assign y12 = n808 ;
  assign y13 = n810 ;
  assign y14 = n812 ;
  assign y15 = n814 ;
  assign y16 = n816 ;
  assign y17 = n818 ;
  assign y18 = ~n819 ;
endmodule
