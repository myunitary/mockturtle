// eight parties, each holding 32-bit data
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 ;
  assign n260 = ~x159 & ~x191 ;
  assign n261 = ~x223 & ~x255 ;
  assign n262 = n260 & n261 ;
  assign n257 = ~x31 & ~x63 ;
  assign n258 = ~x95 & ~x127 ;
  assign n259 = n257 & n258 ;
  assign n263 = n262 ^ n259 ;
  assign n939 = x190 ^ x158 ;
  assign n940 = x191 ^ x159 ;
  assign n1069 = x190 ^ x157 ;
  assign n941 = x188 ^ x156 ;
  assign n1061 = x188 ^ x155 ;
  assign n942 = x186 ^ x154 ;
  assign n1053 = x186 ^ x153 ;
  assign n943 = x184 ^ x152 ;
  assign n1045 = x184 ^ x151 ;
  assign n944 = x182 ^ x150 ;
  assign n1037 = x182 ^ x149 ;
  assign n945 = x180 ^ x148 ;
  assign n1029 = x180 ^ x147 ;
  assign n946 = x178 ^ x146 ;
  assign n1021 = x178 ^ x145 ;
  assign n947 = x176 ^ x144 ;
  assign n1013 = x176 ^ x143 ;
  assign n948 = x174 ^ x142 ;
  assign n1005 = x174 ^ x141 ;
  assign n949 = x172 ^ x140 ;
  assign n997 = x172 ^ x139 ;
  assign n950 = x170 ^ x138 ;
  assign n989 = x170 ^ x137 ;
  assign n951 = x168 ^ x136 ;
  assign n981 = x168 ^ x135 ;
  assign n952 = x166 ^ x134 ;
  assign n973 = x166 ^ x133 ;
  assign n953 = x164 ^ x132 ;
  assign n965 = x164 ^ x131 ;
  assign n954 = x162 ^ x130 ;
  assign n957 = x162 ^ x129 ;
  assign n955 = x128 & ~x160 ;
  assign n956 = n955 ^ x162 ;
  assign n958 = n957 ^ n956 ;
  assign n959 = x161 ^ x129 ;
  assign n960 = n958 & ~n959 ;
  assign n961 = n960 ^ n957 ;
  assign n962 = ~n954 & n961 ;
  assign n963 = n962 ^ x130 ;
  assign n964 = n963 ^ x164 ;
  assign n966 = n965 ^ n964 ;
  assign n967 = x163 ^ x131 ;
  assign n968 = n966 & ~n967 ;
  assign n969 = n968 ^ n965 ;
  assign n970 = ~n953 & n969 ;
  assign n971 = n970 ^ x132 ;
  assign n972 = n971 ^ x166 ;
  assign n974 = n973 ^ n972 ;
  assign n975 = x165 ^ x133 ;
  assign n976 = n974 & ~n975 ;
  assign n977 = n976 ^ n973 ;
  assign n978 = ~n952 & n977 ;
  assign n979 = n978 ^ x134 ;
  assign n980 = n979 ^ x168 ;
  assign n982 = n981 ^ n980 ;
  assign n983 = x167 ^ x135 ;
  assign n984 = n982 & ~n983 ;
  assign n985 = n984 ^ n981 ;
  assign n986 = ~n951 & n985 ;
  assign n987 = n986 ^ x136 ;
  assign n988 = n987 ^ x170 ;
  assign n990 = n989 ^ n988 ;
  assign n991 = x169 ^ x137 ;
  assign n992 = n990 & ~n991 ;
  assign n993 = n992 ^ n989 ;
  assign n994 = ~n950 & n993 ;
  assign n995 = n994 ^ x138 ;
  assign n996 = n995 ^ x172 ;
  assign n998 = n997 ^ n996 ;
  assign n999 = x171 ^ x139 ;
  assign n1000 = n998 & ~n999 ;
  assign n1001 = n1000 ^ n997 ;
  assign n1002 = ~n949 & n1001 ;
  assign n1003 = n1002 ^ x140 ;
  assign n1004 = n1003 ^ x174 ;
  assign n1006 = n1005 ^ n1004 ;
  assign n1007 = x173 ^ x141 ;
  assign n1008 = n1006 & ~n1007 ;
  assign n1009 = n1008 ^ n1005 ;
  assign n1010 = ~n948 & n1009 ;
  assign n1011 = n1010 ^ x142 ;
  assign n1012 = n1011 ^ x176 ;
  assign n1014 = n1013 ^ n1012 ;
  assign n1015 = x175 ^ x143 ;
  assign n1016 = n1014 & ~n1015 ;
  assign n1017 = n1016 ^ n1013 ;
  assign n1018 = ~n947 & n1017 ;
  assign n1019 = n1018 ^ x144 ;
  assign n1020 = n1019 ^ x178 ;
  assign n1022 = n1021 ^ n1020 ;
  assign n1023 = x177 ^ x145 ;
  assign n1024 = n1022 & ~n1023 ;
  assign n1025 = n1024 ^ n1021 ;
  assign n1026 = ~n946 & n1025 ;
  assign n1027 = n1026 ^ x146 ;
  assign n1028 = n1027 ^ x180 ;
  assign n1030 = n1029 ^ n1028 ;
  assign n1031 = x179 ^ x147 ;
  assign n1032 = n1030 & ~n1031 ;
  assign n1033 = n1032 ^ n1029 ;
  assign n1034 = ~n945 & n1033 ;
  assign n1035 = n1034 ^ x148 ;
  assign n1036 = n1035 ^ x182 ;
  assign n1038 = n1037 ^ n1036 ;
  assign n1039 = x181 ^ x149 ;
  assign n1040 = n1038 & ~n1039 ;
  assign n1041 = n1040 ^ n1037 ;
  assign n1042 = ~n944 & n1041 ;
  assign n1043 = n1042 ^ x150 ;
  assign n1044 = n1043 ^ x184 ;
  assign n1046 = n1045 ^ n1044 ;
  assign n1047 = x183 ^ x151 ;
  assign n1048 = n1046 & ~n1047 ;
  assign n1049 = n1048 ^ n1045 ;
  assign n1050 = ~n943 & n1049 ;
  assign n1051 = n1050 ^ x152 ;
  assign n1052 = n1051 ^ x186 ;
  assign n1054 = n1053 ^ n1052 ;
  assign n1055 = x185 ^ x153 ;
  assign n1056 = n1054 & ~n1055 ;
  assign n1057 = n1056 ^ n1053 ;
  assign n1058 = ~n942 & n1057 ;
  assign n1059 = n1058 ^ x154 ;
  assign n1060 = n1059 ^ x188 ;
  assign n1062 = n1061 ^ n1060 ;
  assign n1063 = x187 ^ x155 ;
  assign n1064 = n1062 & ~n1063 ;
  assign n1065 = n1064 ^ n1061 ;
  assign n1066 = ~n941 & n1065 ;
  assign n1067 = n1066 ^ x156 ;
  assign n1068 = n1067 ^ x190 ;
  assign n1070 = n1069 ^ n1068 ;
  assign n1071 = x189 ^ x157 ;
  assign n1072 = n1070 & ~n1071 ;
  assign n1073 = n1072 ^ n1069 ;
  assign n1074 = ~n939 & n1073 ;
  assign n1075 = n1074 ^ x158 ;
  assign n1076 = n1075 ^ x191 ;
  assign n1077 = ~n940 & n1076 ;
  assign n1078 = n1077 ^ x159 ;
  assign n1079 = n939 & ~n1078 ;
  assign n1080 = n1079 ^ x158 ;
  assign n797 = x254 ^ x222 ;
  assign n798 = x255 ^ x223 ;
  assign n927 = x254 ^ x221 ;
  assign n799 = x252 ^ x220 ;
  assign n919 = x252 ^ x219 ;
  assign n800 = x250 ^ x218 ;
  assign n911 = x250 ^ x217 ;
  assign n801 = x248 ^ x216 ;
  assign n903 = x248 ^ x215 ;
  assign n802 = x246 ^ x214 ;
  assign n895 = x246 ^ x213 ;
  assign n803 = x244 ^ x212 ;
  assign n887 = x244 ^ x211 ;
  assign n804 = x242 ^ x210 ;
  assign n879 = x242 ^ x209 ;
  assign n805 = x240 ^ x208 ;
  assign n871 = x240 ^ x207 ;
  assign n806 = x238 ^ x206 ;
  assign n863 = x238 ^ x205 ;
  assign n807 = x236 ^ x204 ;
  assign n855 = x236 ^ x203 ;
  assign n808 = x234 ^ x202 ;
  assign n847 = x234 ^ x201 ;
  assign n809 = x232 ^ x200 ;
  assign n839 = x232 ^ x199 ;
  assign n810 = x230 ^ x198 ;
  assign n831 = x230 ^ x197 ;
  assign n811 = x228 ^ x196 ;
  assign n823 = x228 ^ x195 ;
  assign n812 = x226 ^ x194 ;
  assign n815 = x226 ^ x193 ;
  assign n813 = x192 & ~x224 ;
  assign n814 = n813 ^ x226 ;
  assign n816 = n815 ^ n814 ;
  assign n817 = x225 ^ x193 ;
  assign n818 = n816 & ~n817 ;
  assign n819 = n818 ^ n815 ;
  assign n820 = ~n812 & n819 ;
  assign n821 = n820 ^ x194 ;
  assign n822 = n821 ^ x228 ;
  assign n824 = n823 ^ n822 ;
  assign n825 = x227 ^ x195 ;
  assign n826 = n824 & ~n825 ;
  assign n827 = n826 ^ n823 ;
  assign n828 = ~n811 & n827 ;
  assign n829 = n828 ^ x196 ;
  assign n830 = n829 ^ x230 ;
  assign n832 = n831 ^ n830 ;
  assign n833 = x229 ^ x197 ;
  assign n834 = n832 & ~n833 ;
  assign n835 = n834 ^ n831 ;
  assign n836 = ~n810 & n835 ;
  assign n837 = n836 ^ x198 ;
  assign n838 = n837 ^ x232 ;
  assign n840 = n839 ^ n838 ;
  assign n841 = x231 ^ x199 ;
  assign n842 = n840 & ~n841 ;
  assign n843 = n842 ^ n839 ;
  assign n844 = ~n809 & n843 ;
  assign n845 = n844 ^ x200 ;
  assign n846 = n845 ^ x234 ;
  assign n848 = n847 ^ n846 ;
  assign n849 = x233 ^ x201 ;
  assign n850 = n848 & ~n849 ;
  assign n851 = n850 ^ n847 ;
  assign n852 = ~n808 & n851 ;
  assign n853 = n852 ^ x202 ;
  assign n854 = n853 ^ x236 ;
  assign n856 = n855 ^ n854 ;
  assign n857 = x235 ^ x203 ;
  assign n858 = n856 & ~n857 ;
  assign n859 = n858 ^ n855 ;
  assign n860 = ~n807 & n859 ;
  assign n861 = n860 ^ x204 ;
  assign n862 = n861 ^ x238 ;
  assign n864 = n863 ^ n862 ;
  assign n865 = x237 ^ x205 ;
  assign n866 = n864 & ~n865 ;
  assign n867 = n866 ^ n863 ;
  assign n868 = ~n806 & n867 ;
  assign n869 = n868 ^ x206 ;
  assign n870 = n869 ^ x240 ;
  assign n872 = n871 ^ n870 ;
  assign n873 = x239 ^ x207 ;
  assign n874 = n872 & ~n873 ;
  assign n875 = n874 ^ n871 ;
  assign n876 = ~n805 & n875 ;
  assign n877 = n876 ^ x208 ;
  assign n878 = n877 ^ x242 ;
  assign n880 = n879 ^ n878 ;
  assign n881 = x241 ^ x209 ;
  assign n882 = n880 & ~n881 ;
  assign n883 = n882 ^ n879 ;
  assign n884 = ~n804 & n883 ;
  assign n885 = n884 ^ x210 ;
  assign n886 = n885 ^ x244 ;
  assign n888 = n887 ^ n886 ;
  assign n889 = x243 ^ x211 ;
  assign n890 = n888 & ~n889 ;
  assign n891 = n890 ^ n887 ;
  assign n892 = ~n803 & n891 ;
  assign n893 = n892 ^ x212 ;
  assign n894 = n893 ^ x246 ;
  assign n896 = n895 ^ n894 ;
  assign n897 = x245 ^ x213 ;
  assign n898 = n896 & ~n897 ;
  assign n899 = n898 ^ n895 ;
  assign n900 = ~n802 & n899 ;
  assign n901 = n900 ^ x214 ;
  assign n902 = n901 ^ x248 ;
  assign n904 = n903 ^ n902 ;
  assign n905 = x247 ^ x215 ;
  assign n906 = n904 & ~n905 ;
  assign n907 = n906 ^ n903 ;
  assign n908 = ~n801 & n907 ;
  assign n909 = n908 ^ x216 ;
  assign n910 = n909 ^ x250 ;
  assign n912 = n911 ^ n910 ;
  assign n913 = x249 ^ x217 ;
  assign n914 = n912 & ~n913 ;
  assign n915 = n914 ^ n911 ;
  assign n916 = ~n800 & n915 ;
  assign n917 = n916 ^ x218 ;
  assign n918 = n917 ^ x252 ;
  assign n920 = n919 ^ n918 ;
  assign n921 = x251 ^ x219 ;
  assign n922 = n920 & ~n921 ;
  assign n923 = n922 ^ n919 ;
  assign n924 = ~n799 & n923 ;
  assign n925 = n924 ^ x220 ;
  assign n926 = n925 ^ x254 ;
  assign n928 = n927 ^ n926 ;
  assign n929 = x253 ^ x221 ;
  assign n930 = n928 & ~n929 ;
  assign n931 = n930 ^ n927 ;
  assign n932 = ~n797 & n931 ;
  assign n933 = n932 ^ x222 ;
  assign n934 = n933 ^ x255 ;
  assign n935 = ~n798 & n934 ;
  assign n936 = n935 ^ x223 ;
  assign n937 = n797 & ~n936 ;
  assign n938 = n937 ^ x222 ;
  assign n1081 = n1080 ^ n938 ;
  assign n1082 = n261 ^ n260 ;
  assign n1085 = n929 & ~n936 ;
  assign n1086 = n1085 ^ x221 ;
  assign n1083 = n1071 & ~n1078 ;
  assign n1084 = n1083 ^ x157 ;
  assign n1087 = n1086 ^ n1084 ;
  assign n1090 = n799 & ~n936 ;
  assign n1091 = n1090 ^ x220 ;
  assign n1088 = n941 & ~n1078 ;
  assign n1089 = n1088 ^ x156 ;
  assign n1092 = n1091 ^ n1089 ;
  assign n1095 = n1063 & ~n1078 ;
  assign n1096 = n1095 ^ x155 ;
  assign n1093 = n921 & ~n936 ;
  assign n1094 = n1093 ^ x219 ;
  assign n1097 = n1096 ^ n1094 ;
  assign n1100 = n942 & ~n1078 ;
  assign n1101 = n1100 ^ x154 ;
  assign n1098 = n800 & ~n936 ;
  assign n1099 = n1098 ^ x218 ;
  assign n1102 = n1101 ^ n1099 ;
  assign n1105 = n913 & ~n936 ;
  assign n1106 = n1105 ^ x217 ;
  assign n1103 = n1055 & ~n1078 ;
  assign n1104 = n1103 ^ x153 ;
  assign n1107 = n1106 ^ n1104 ;
  assign n1110 = n943 & ~n1078 ;
  assign n1111 = n1110 ^ x152 ;
  assign n1108 = n801 & ~n936 ;
  assign n1109 = n1108 ^ x216 ;
  assign n1112 = n1111 ^ n1109 ;
  assign n1115 = n905 & ~n936 ;
  assign n1116 = n1115 ^ x215 ;
  assign n1113 = n1047 & ~n1078 ;
  assign n1114 = n1113 ^ x151 ;
  assign n1117 = n1116 ^ n1114 ;
  assign n1120 = n944 & ~n1078 ;
  assign n1121 = n1120 ^ x150 ;
  assign n1118 = n802 & ~n936 ;
  assign n1119 = n1118 ^ x214 ;
  assign n1122 = n1121 ^ n1119 ;
  assign n1125 = n897 & ~n936 ;
  assign n1126 = n1125 ^ x213 ;
  assign n1123 = n1039 & ~n1078 ;
  assign n1124 = n1123 ^ x149 ;
  assign n1127 = n1126 ^ n1124 ;
  assign n1130 = n945 & ~n1078 ;
  assign n1131 = n1130 ^ x148 ;
  assign n1128 = n803 & ~n936 ;
  assign n1129 = n1128 ^ x212 ;
  assign n1132 = n1131 ^ n1129 ;
  assign n1135 = n889 & ~n936 ;
  assign n1136 = n1135 ^ x211 ;
  assign n1133 = n1031 & ~n1078 ;
  assign n1134 = n1133 ^ x147 ;
  assign n1137 = n1136 ^ n1134 ;
  assign n1140 = n946 & ~n1078 ;
  assign n1141 = n1140 ^ x146 ;
  assign n1138 = n804 & ~n936 ;
  assign n1139 = n1138 ^ x210 ;
  assign n1142 = n1141 ^ n1139 ;
  assign n1145 = n881 & ~n936 ;
  assign n1146 = n1145 ^ x209 ;
  assign n1143 = n1023 & ~n1078 ;
  assign n1144 = n1143 ^ x145 ;
  assign n1147 = n1146 ^ n1144 ;
  assign n1150 = n947 & ~n1078 ;
  assign n1151 = n1150 ^ x144 ;
  assign n1148 = n805 & ~n936 ;
  assign n1149 = n1148 ^ x208 ;
  assign n1152 = n1151 ^ n1149 ;
  assign n1155 = n873 & ~n936 ;
  assign n1156 = n1155 ^ x207 ;
  assign n1153 = n1015 & ~n1078 ;
  assign n1154 = n1153 ^ x143 ;
  assign n1157 = n1156 ^ n1154 ;
  assign n1160 = n948 & ~n1078 ;
  assign n1161 = n1160 ^ x142 ;
  assign n1158 = n806 & ~n936 ;
  assign n1159 = n1158 ^ x206 ;
  assign n1162 = n1161 ^ n1159 ;
  assign n1165 = n865 & ~n936 ;
  assign n1166 = n1165 ^ x205 ;
  assign n1163 = n1007 & ~n1078 ;
  assign n1164 = n1163 ^ x141 ;
  assign n1167 = n1166 ^ n1164 ;
  assign n1170 = n949 & ~n1078 ;
  assign n1171 = n1170 ^ x140 ;
  assign n1168 = n807 & ~n936 ;
  assign n1169 = n1168 ^ x204 ;
  assign n1172 = n1171 ^ n1169 ;
  assign n1175 = n857 & ~n936 ;
  assign n1176 = n1175 ^ x203 ;
  assign n1173 = n999 & ~n1078 ;
  assign n1174 = n1173 ^ x139 ;
  assign n1177 = n1176 ^ n1174 ;
  assign n1180 = n950 & ~n1078 ;
  assign n1181 = n1180 ^ x138 ;
  assign n1178 = n808 & ~n936 ;
  assign n1179 = n1178 ^ x202 ;
  assign n1182 = n1181 ^ n1179 ;
  assign n1185 = n849 & ~n936 ;
  assign n1186 = n1185 ^ x201 ;
  assign n1183 = n991 & ~n1078 ;
  assign n1184 = n1183 ^ x137 ;
  assign n1187 = n1186 ^ n1184 ;
  assign n1190 = n951 & ~n1078 ;
  assign n1191 = n1190 ^ x136 ;
  assign n1188 = n809 & ~n936 ;
  assign n1189 = n1188 ^ x200 ;
  assign n1192 = n1191 ^ n1189 ;
  assign n1195 = n841 & ~n936 ;
  assign n1196 = n1195 ^ x199 ;
  assign n1193 = n983 & ~n1078 ;
  assign n1194 = n1193 ^ x135 ;
  assign n1197 = n1196 ^ n1194 ;
  assign n1200 = n810 & ~n936 ;
  assign n1201 = n1200 ^ x198 ;
  assign n1198 = n952 & ~n1078 ;
  assign n1199 = n1198 ^ x134 ;
  assign n1202 = n1201 ^ n1199 ;
  assign n1205 = n833 & ~n936 ;
  assign n1206 = n1205 ^ x197 ;
  assign n1203 = n975 & ~n1078 ;
  assign n1204 = n1203 ^ x133 ;
  assign n1207 = n1206 ^ n1204 ;
  assign n1210 = n811 & ~n936 ;
  assign n1211 = n1210 ^ x196 ;
  assign n1208 = n953 & ~n1078 ;
  assign n1209 = n1208 ^ x132 ;
  assign n1212 = n1211 ^ n1209 ;
  assign n1215 = n967 & ~n1078 ;
  assign n1216 = n1215 ^ x131 ;
  assign n1213 = n825 & ~n936 ;
  assign n1214 = n1213 ^ x195 ;
  assign n1217 = n1216 ^ n1214 ;
  assign n1220 = n812 & ~n936 ;
  assign n1221 = n1220 ^ x194 ;
  assign n1218 = n954 & ~n1078 ;
  assign n1219 = n1218 ^ x130 ;
  assign n1222 = n1221 ^ n1219 ;
  assign n1225 = n959 & ~n1078 ;
  assign n1226 = n1225 ^ x129 ;
  assign n1223 = n817 & ~n936 ;
  assign n1224 = n1223 ^ x193 ;
  assign n1227 = n1226 ^ n1224 ;
  assign n1228 = x224 ^ x192 ;
  assign n1229 = ~n936 & n1228 ;
  assign n1230 = n1229 ^ x192 ;
  assign n1231 = x160 ^ x128 ;
  assign n1232 = ~n1078 & n1231 ;
  assign n1233 = n1232 ^ x128 ;
  assign n1234 = ~n1230 & n1233 ;
  assign n1235 = n1234 ^ n1224 ;
  assign n1236 = ~n1227 & ~n1235 ;
  assign n1237 = n1236 ^ n1224 ;
  assign n1238 = n1237 ^ n1221 ;
  assign n1239 = ~n1222 & n1238 ;
  assign n1240 = n1239 ^ n1221 ;
  assign n1241 = n1240 ^ n1214 ;
  assign n1242 = ~n1217 & n1241 ;
  assign n1243 = n1242 ^ n1214 ;
  assign n1244 = n1243 ^ n1211 ;
  assign n1245 = ~n1212 & n1244 ;
  assign n1246 = n1245 ^ n1211 ;
  assign n1247 = n1246 ^ n1204 ;
  assign n1248 = ~n1207 & ~n1247 ;
  assign n1249 = n1248 ^ n1204 ;
  assign n1250 = n1249 ^ n1201 ;
  assign n1251 = ~n1202 & ~n1250 ;
  assign n1252 = n1251 ^ n1201 ;
  assign n1253 = n1252 ^ n1194 ;
  assign n1254 = ~n1197 & ~n1253 ;
  assign n1255 = n1254 ^ n1194 ;
  assign n1256 = n1255 ^ n1191 ;
  assign n1257 = ~n1192 & n1256 ;
  assign n1258 = n1257 ^ n1191 ;
  assign n1259 = n1258 ^ n1184 ;
  assign n1260 = ~n1187 & n1259 ;
  assign n1261 = n1260 ^ n1184 ;
  assign n1262 = n1261 ^ n1181 ;
  assign n1263 = ~n1182 & n1262 ;
  assign n1264 = n1263 ^ n1181 ;
  assign n1265 = n1264 ^ n1174 ;
  assign n1266 = ~n1177 & n1265 ;
  assign n1267 = n1266 ^ n1174 ;
  assign n1268 = n1267 ^ n1171 ;
  assign n1269 = ~n1172 & n1268 ;
  assign n1270 = n1269 ^ n1171 ;
  assign n1271 = n1270 ^ n1164 ;
  assign n1272 = ~n1167 & n1271 ;
  assign n1273 = n1272 ^ n1164 ;
  assign n1274 = n1273 ^ n1161 ;
  assign n1275 = ~n1162 & n1274 ;
  assign n1276 = n1275 ^ n1161 ;
  assign n1277 = n1276 ^ n1154 ;
  assign n1278 = ~n1157 & n1277 ;
  assign n1279 = n1278 ^ n1154 ;
  assign n1280 = n1279 ^ n1151 ;
  assign n1281 = ~n1152 & n1280 ;
  assign n1282 = n1281 ^ n1151 ;
  assign n1283 = n1282 ^ n1144 ;
  assign n1284 = ~n1147 & n1283 ;
  assign n1285 = n1284 ^ n1144 ;
  assign n1286 = n1285 ^ n1141 ;
  assign n1287 = ~n1142 & n1286 ;
  assign n1288 = n1287 ^ n1141 ;
  assign n1289 = n1288 ^ n1134 ;
  assign n1290 = ~n1137 & n1289 ;
  assign n1291 = n1290 ^ n1134 ;
  assign n1292 = n1291 ^ n1131 ;
  assign n1293 = ~n1132 & n1292 ;
  assign n1294 = n1293 ^ n1131 ;
  assign n1295 = n1294 ^ n1124 ;
  assign n1296 = ~n1127 & n1295 ;
  assign n1297 = n1296 ^ n1124 ;
  assign n1298 = n1297 ^ n1121 ;
  assign n1299 = ~n1122 & n1298 ;
  assign n1300 = n1299 ^ n1121 ;
  assign n1301 = n1300 ^ n1114 ;
  assign n1302 = ~n1117 & n1301 ;
  assign n1303 = n1302 ^ n1114 ;
  assign n1304 = n1303 ^ n1111 ;
  assign n1305 = ~n1112 & n1304 ;
  assign n1306 = n1305 ^ n1111 ;
  assign n1307 = n1306 ^ n1104 ;
  assign n1308 = ~n1107 & n1307 ;
  assign n1309 = n1308 ^ n1104 ;
  assign n1310 = n1309 ^ n1101 ;
  assign n1311 = ~n1102 & n1310 ;
  assign n1312 = n1311 ^ n1101 ;
  assign n1313 = n1312 ^ n1094 ;
  assign n1314 = ~n1097 & ~n1313 ;
  assign n1315 = n1314 ^ n1094 ;
  assign n1316 = n1315 ^ n1089 ;
  assign n1317 = ~n1092 & ~n1316 ;
  assign n1318 = n1317 ^ n1089 ;
  assign n1319 = n1318 ^ n1084 ;
  assign n1320 = ~n1087 & ~n1319 ;
  assign n1321 = n1320 ^ n1086 ;
  assign n1322 = n1321 ^ n938 ;
  assign n1323 = ~n1081 & ~n1322 ;
  assign n1324 = n1323 ^ n1080 ;
  assign n1325 = n1324 ^ n261 ;
  assign n1326 = ~n1082 & ~n1325 ;
  assign n1327 = n1326 ^ n260 ;
  assign n1328 = n1081 & n1327 ;
  assign n1329 = n1328 ^ n1080 ;
  assign n406 = x126 ^ x94 ;
  assign n407 = x127 ^ x95 ;
  assign n536 = x126 ^ x93 ;
  assign n408 = x124 ^ x92 ;
  assign n528 = x124 ^ x91 ;
  assign n409 = x122 ^ x90 ;
  assign n520 = x122 ^ x89 ;
  assign n410 = x120 ^ x88 ;
  assign n512 = x120 ^ x87 ;
  assign n411 = x118 ^ x86 ;
  assign n504 = x118 ^ x85 ;
  assign n412 = x116 ^ x84 ;
  assign n496 = x116 ^ x83 ;
  assign n413 = x114 ^ x82 ;
  assign n488 = x114 ^ x81 ;
  assign n414 = x112 ^ x80 ;
  assign n480 = x112 ^ x79 ;
  assign n415 = x110 ^ x78 ;
  assign n472 = x110 ^ x77 ;
  assign n416 = x108 ^ x76 ;
  assign n464 = x108 ^ x75 ;
  assign n417 = x106 ^ x74 ;
  assign n456 = x106 ^ x73 ;
  assign n418 = x104 ^ x72 ;
  assign n448 = x104 ^ x71 ;
  assign n419 = x102 ^ x70 ;
  assign n440 = x102 ^ x69 ;
  assign n420 = x100 ^ x68 ;
  assign n432 = x100 ^ x67 ;
  assign n421 = x98 ^ x66 ;
  assign n424 = x98 ^ x65 ;
  assign n422 = x64 & ~x96 ;
  assign n423 = n422 ^ x98 ;
  assign n425 = n424 ^ n423 ;
  assign n426 = x97 ^ x65 ;
  assign n427 = n425 & ~n426 ;
  assign n428 = n427 ^ n424 ;
  assign n429 = ~n421 & n428 ;
  assign n430 = n429 ^ x66 ;
  assign n431 = n430 ^ x100 ;
  assign n433 = n432 ^ n431 ;
  assign n434 = x99 ^ x67 ;
  assign n435 = n433 & ~n434 ;
  assign n436 = n435 ^ n432 ;
  assign n437 = ~n420 & n436 ;
  assign n438 = n437 ^ x68 ;
  assign n439 = n438 ^ x102 ;
  assign n441 = n440 ^ n439 ;
  assign n442 = x101 ^ x69 ;
  assign n443 = n441 & ~n442 ;
  assign n444 = n443 ^ n440 ;
  assign n445 = ~n419 & n444 ;
  assign n446 = n445 ^ x70 ;
  assign n447 = n446 ^ x104 ;
  assign n449 = n448 ^ n447 ;
  assign n450 = x103 ^ x71 ;
  assign n451 = n449 & ~n450 ;
  assign n452 = n451 ^ n448 ;
  assign n453 = ~n418 & n452 ;
  assign n454 = n453 ^ x72 ;
  assign n455 = n454 ^ x106 ;
  assign n457 = n456 ^ n455 ;
  assign n458 = x105 ^ x73 ;
  assign n459 = n457 & ~n458 ;
  assign n460 = n459 ^ n456 ;
  assign n461 = ~n417 & n460 ;
  assign n462 = n461 ^ x74 ;
  assign n463 = n462 ^ x108 ;
  assign n465 = n464 ^ n463 ;
  assign n466 = x107 ^ x75 ;
  assign n467 = n465 & ~n466 ;
  assign n468 = n467 ^ n464 ;
  assign n469 = ~n416 & n468 ;
  assign n470 = n469 ^ x76 ;
  assign n471 = n470 ^ x110 ;
  assign n473 = n472 ^ n471 ;
  assign n474 = x109 ^ x77 ;
  assign n475 = n473 & ~n474 ;
  assign n476 = n475 ^ n472 ;
  assign n477 = ~n415 & n476 ;
  assign n478 = n477 ^ x78 ;
  assign n479 = n478 ^ x112 ;
  assign n481 = n480 ^ n479 ;
  assign n482 = x111 ^ x79 ;
  assign n483 = n481 & ~n482 ;
  assign n484 = n483 ^ n480 ;
  assign n485 = ~n414 & n484 ;
  assign n486 = n485 ^ x80 ;
  assign n487 = n486 ^ x114 ;
  assign n489 = n488 ^ n487 ;
  assign n490 = x113 ^ x81 ;
  assign n491 = n489 & ~n490 ;
  assign n492 = n491 ^ n488 ;
  assign n493 = ~n413 & n492 ;
  assign n494 = n493 ^ x82 ;
  assign n495 = n494 ^ x116 ;
  assign n497 = n496 ^ n495 ;
  assign n498 = x115 ^ x83 ;
  assign n499 = n497 & ~n498 ;
  assign n500 = n499 ^ n496 ;
  assign n501 = ~n412 & n500 ;
  assign n502 = n501 ^ x84 ;
  assign n503 = n502 ^ x118 ;
  assign n505 = n504 ^ n503 ;
  assign n506 = x117 ^ x85 ;
  assign n507 = n505 & ~n506 ;
  assign n508 = n507 ^ n504 ;
  assign n509 = ~n411 & n508 ;
  assign n510 = n509 ^ x86 ;
  assign n511 = n510 ^ x120 ;
  assign n513 = n512 ^ n511 ;
  assign n514 = x119 ^ x87 ;
  assign n515 = n513 & ~n514 ;
  assign n516 = n515 ^ n512 ;
  assign n517 = ~n410 & n516 ;
  assign n518 = n517 ^ x88 ;
  assign n519 = n518 ^ x122 ;
  assign n521 = n520 ^ n519 ;
  assign n522 = x121 ^ x89 ;
  assign n523 = n521 & ~n522 ;
  assign n524 = n523 ^ n520 ;
  assign n525 = ~n409 & n524 ;
  assign n526 = n525 ^ x90 ;
  assign n527 = n526 ^ x124 ;
  assign n529 = n528 ^ n527 ;
  assign n530 = x123 ^ x91 ;
  assign n531 = n529 & ~n530 ;
  assign n532 = n531 ^ n528 ;
  assign n533 = ~n408 & n532 ;
  assign n534 = n533 ^ x92 ;
  assign n535 = n534 ^ x126 ;
  assign n537 = n536 ^ n535 ;
  assign n538 = x125 ^ x93 ;
  assign n539 = n537 & ~n538 ;
  assign n540 = n539 ^ n536 ;
  assign n541 = ~n406 & n540 ;
  assign n542 = n541 ^ x94 ;
  assign n543 = n542 ^ x127 ;
  assign n544 = ~n407 & n543 ;
  assign n545 = n544 ^ x95 ;
  assign n546 = n406 & ~n545 ;
  assign n547 = n546 ^ x94 ;
  assign n264 = x62 ^ x30 ;
  assign n265 = x63 ^ x31 ;
  assign n394 = x62 ^ x29 ;
  assign n266 = x60 ^ x28 ;
  assign n386 = x60 ^ x27 ;
  assign n267 = x58 ^ x26 ;
  assign n378 = x58 ^ x25 ;
  assign n268 = x56 ^ x24 ;
  assign n370 = x56 ^ x23 ;
  assign n269 = x54 ^ x22 ;
  assign n362 = x54 ^ x21 ;
  assign n270 = x52 ^ x20 ;
  assign n354 = x52 ^ x19 ;
  assign n271 = x50 ^ x18 ;
  assign n346 = x50 ^ x17 ;
  assign n272 = x48 ^ x16 ;
  assign n338 = x48 ^ x15 ;
  assign n273 = x46 ^ x14 ;
  assign n330 = x46 ^ x13 ;
  assign n274 = x44 ^ x12 ;
  assign n322 = x44 ^ x11 ;
  assign n275 = x42 ^ x10 ;
  assign n314 = x42 ^ x9 ;
  assign n276 = x40 ^ x8 ;
  assign n306 = x40 ^ x7 ;
  assign n277 = x38 ^ x6 ;
  assign n298 = x38 ^ x5 ;
  assign n278 = x36 ^ x4 ;
  assign n290 = x36 ^ x3 ;
  assign n279 = x34 ^ x2 ;
  assign n282 = x34 ^ x1 ;
  assign n280 = x0 & ~x32 ;
  assign n281 = n280 ^ x34 ;
  assign n283 = n282 ^ n281 ;
  assign n284 = x33 ^ x1 ;
  assign n285 = n283 & ~n284 ;
  assign n286 = n285 ^ n282 ;
  assign n287 = ~n279 & n286 ;
  assign n288 = n287 ^ x2 ;
  assign n289 = n288 ^ x36 ;
  assign n291 = n290 ^ n289 ;
  assign n292 = x35 ^ x3 ;
  assign n293 = n291 & ~n292 ;
  assign n294 = n293 ^ n290 ;
  assign n295 = ~n278 & n294 ;
  assign n296 = n295 ^ x4 ;
  assign n297 = n296 ^ x38 ;
  assign n299 = n298 ^ n297 ;
  assign n300 = x37 ^ x5 ;
  assign n301 = n299 & ~n300 ;
  assign n302 = n301 ^ n298 ;
  assign n303 = ~n277 & n302 ;
  assign n304 = n303 ^ x6 ;
  assign n305 = n304 ^ x40 ;
  assign n307 = n306 ^ n305 ;
  assign n308 = x39 ^ x7 ;
  assign n309 = n307 & ~n308 ;
  assign n310 = n309 ^ n306 ;
  assign n311 = ~n276 & n310 ;
  assign n312 = n311 ^ x8 ;
  assign n313 = n312 ^ x42 ;
  assign n315 = n314 ^ n313 ;
  assign n316 = x41 ^ x9 ;
  assign n317 = n315 & ~n316 ;
  assign n318 = n317 ^ n314 ;
  assign n319 = ~n275 & n318 ;
  assign n320 = n319 ^ x10 ;
  assign n321 = n320 ^ x44 ;
  assign n323 = n322 ^ n321 ;
  assign n324 = x43 ^ x11 ;
  assign n325 = n323 & ~n324 ;
  assign n326 = n325 ^ n322 ;
  assign n327 = ~n274 & n326 ;
  assign n328 = n327 ^ x12 ;
  assign n329 = n328 ^ x46 ;
  assign n331 = n330 ^ n329 ;
  assign n332 = x45 ^ x13 ;
  assign n333 = n331 & ~n332 ;
  assign n334 = n333 ^ n330 ;
  assign n335 = ~n273 & n334 ;
  assign n336 = n335 ^ x14 ;
  assign n337 = n336 ^ x48 ;
  assign n339 = n338 ^ n337 ;
  assign n340 = x47 ^ x15 ;
  assign n341 = n339 & ~n340 ;
  assign n342 = n341 ^ n338 ;
  assign n343 = ~n272 & n342 ;
  assign n344 = n343 ^ x16 ;
  assign n345 = n344 ^ x50 ;
  assign n347 = n346 ^ n345 ;
  assign n348 = x49 ^ x17 ;
  assign n349 = n347 & ~n348 ;
  assign n350 = n349 ^ n346 ;
  assign n351 = ~n271 & n350 ;
  assign n352 = n351 ^ x18 ;
  assign n353 = n352 ^ x52 ;
  assign n355 = n354 ^ n353 ;
  assign n356 = x51 ^ x19 ;
  assign n357 = n355 & ~n356 ;
  assign n358 = n357 ^ n354 ;
  assign n359 = ~n270 & n358 ;
  assign n360 = n359 ^ x20 ;
  assign n361 = n360 ^ x54 ;
  assign n363 = n362 ^ n361 ;
  assign n364 = x53 ^ x21 ;
  assign n365 = n363 & ~n364 ;
  assign n366 = n365 ^ n362 ;
  assign n367 = ~n269 & n366 ;
  assign n368 = n367 ^ x22 ;
  assign n369 = n368 ^ x56 ;
  assign n371 = n370 ^ n369 ;
  assign n372 = x55 ^ x23 ;
  assign n373 = n371 & ~n372 ;
  assign n374 = n373 ^ n370 ;
  assign n375 = ~n268 & n374 ;
  assign n376 = n375 ^ x24 ;
  assign n377 = n376 ^ x58 ;
  assign n379 = n378 ^ n377 ;
  assign n380 = x57 ^ x25 ;
  assign n381 = n379 & ~n380 ;
  assign n382 = n381 ^ n378 ;
  assign n383 = ~n267 & n382 ;
  assign n384 = n383 ^ x26 ;
  assign n385 = n384 ^ x60 ;
  assign n387 = n386 ^ n385 ;
  assign n388 = x59 ^ x27 ;
  assign n389 = n387 & ~n388 ;
  assign n390 = n389 ^ n386 ;
  assign n391 = ~n266 & n390 ;
  assign n392 = n391 ^ x28 ;
  assign n393 = n392 ^ x62 ;
  assign n395 = n394 ^ n393 ;
  assign n396 = x61 ^ x29 ;
  assign n397 = n395 & ~n396 ;
  assign n398 = n397 ^ n394 ;
  assign n399 = ~n264 & n398 ;
  assign n400 = n399 ^ x30 ;
  assign n401 = n400 ^ x63 ;
  assign n402 = ~n265 & n401 ;
  assign n403 = n402 ^ x31 ;
  assign n404 = n264 & ~n403 ;
  assign n405 = n404 ^ x30 ;
  assign n548 = n547 ^ n405 ;
  assign n549 = n258 ^ n257 ;
  assign n552 = n538 & ~n545 ;
  assign n553 = n552 ^ x93 ;
  assign n550 = n396 & ~n403 ;
  assign n551 = n550 ^ x29 ;
  assign n554 = n553 ^ n551 ;
  assign n557 = n266 & ~n403 ;
  assign n558 = n557 ^ x28 ;
  assign n555 = n408 & ~n545 ;
  assign n556 = n555 ^ x92 ;
  assign n559 = n558 ^ n556 ;
  assign n562 = n530 & ~n545 ;
  assign n563 = n562 ^ x91 ;
  assign n560 = n388 & ~n403 ;
  assign n561 = n560 ^ x27 ;
  assign n564 = n563 ^ n561 ;
  assign n567 = n267 & ~n403 ;
  assign n568 = n567 ^ x26 ;
  assign n565 = n409 & ~n545 ;
  assign n566 = n565 ^ x90 ;
  assign n569 = n568 ^ n566 ;
  assign n572 = n522 & ~n545 ;
  assign n573 = n572 ^ x89 ;
  assign n570 = n380 & ~n403 ;
  assign n571 = n570 ^ x25 ;
  assign n574 = n573 ^ n571 ;
  assign n577 = n410 & ~n545 ;
  assign n578 = n577 ^ x88 ;
  assign n575 = n268 & ~n403 ;
  assign n576 = n575 ^ x24 ;
  assign n579 = n578 ^ n576 ;
  assign n582 = n514 & ~n545 ;
  assign n583 = n582 ^ x87 ;
  assign n580 = n372 & ~n403 ;
  assign n581 = n580 ^ x23 ;
  assign n584 = n583 ^ n581 ;
  assign n587 = n269 & ~n403 ;
  assign n588 = n587 ^ x22 ;
  assign n585 = n411 & ~n545 ;
  assign n586 = n585 ^ x86 ;
  assign n589 = n588 ^ n586 ;
  assign n592 = n506 & ~n545 ;
  assign n593 = n592 ^ x85 ;
  assign n590 = n364 & ~n403 ;
  assign n591 = n590 ^ x21 ;
  assign n594 = n593 ^ n591 ;
  assign n597 = n270 & ~n403 ;
  assign n598 = n597 ^ x20 ;
  assign n595 = n412 & ~n545 ;
  assign n596 = n595 ^ x84 ;
  assign n599 = n598 ^ n596 ;
  assign n602 = n498 & ~n545 ;
  assign n603 = n602 ^ x83 ;
  assign n600 = n356 & ~n403 ;
  assign n601 = n600 ^ x19 ;
  assign n604 = n603 ^ n601 ;
  assign n607 = n271 & ~n403 ;
  assign n608 = n607 ^ x18 ;
  assign n605 = n413 & ~n545 ;
  assign n606 = n605 ^ x82 ;
  assign n609 = n608 ^ n606 ;
  assign n612 = n490 & ~n545 ;
  assign n613 = n612 ^ x81 ;
  assign n610 = n348 & ~n403 ;
  assign n611 = n610 ^ x17 ;
  assign n614 = n613 ^ n611 ;
  assign n617 = n272 & ~n403 ;
  assign n618 = n617 ^ x16 ;
  assign n615 = n414 & ~n545 ;
  assign n616 = n615 ^ x80 ;
  assign n619 = n618 ^ n616 ;
  assign n622 = n482 & ~n545 ;
  assign n623 = n622 ^ x79 ;
  assign n620 = n340 & ~n403 ;
  assign n621 = n620 ^ x15 ;
  assign n624 = n623 ^ n621 ;
  assign n627 = n273 & ~n403 ;
  assign n628 = n627 ^ x14 ;
  assign n625 = n415 & ~n545 ;
  assign n626 = n625 ^ x78 ;
  assign n629 = n628 ^ n626 ;
  assign n632 = n474 & ~n545 ;
  assign n633 = n632 ^ x77 ;
  assign n630 = n332 & ~n403 ;
  assign n631 = n630 ^ x13 ;
  assign n634 = n633 ^ n631 ;
  assign n637 = n274 & ~n403 ;
  assign n638 = n637 ^ x12 ;
  assign n635 = n416 & ~n545 ;
  assign n636 = n635 ^ x76 ;
  assign n639 = n638 ^ n636 ;
  assign n642 = n466 & ~n545 ;
  assign n643 = n642 ^ x75 ;
  assign n640 = n324 & ~n403 ;
  assign n641 = n640 ^ x11 ;
  assign n644 = n643 ^ n641 ;
  assign n647 = n275 & ~n403 ;
  assign n648 = n647 ^ x10 ;
  assign n645 = n417 & ~n545 ;
  assign n646 = n645 ^ x74 ;
  assign n649 = n648 ^ n646 ;
  assign n652 = n458 & ~n545 ;
  assign n653 = n652 ^ x73 ;
  assign n650 = n316 & ~n403 ;
  assign n651 = n650 ^ x9 ;
  assign n654 = n653 ^ n651 ;
  assign n657 = n276 & ~n403 ;
  assign n658 = n657 ^ x8 ;
  assign n655 = n418 & ~n545 ;
  assign n656 = n655 ^ x72 ;
  assign n659 = n658 ^ n656 ;
  assign n662 = n450 & ~n545 ;
  assign n663 = n662 ^ x71 ;
  assign n660 = n308 & ~n403 ;
  assign n661 = n660 ^ x7 ;
  assign n664 = n663 ^ n661 ;
  assign n667 = n277 & ~n403 ;
  assign n668 = n667 ^ x6 ;
  assign n665 = n419 & ~n545 ;
  assign n666 = n665 ^ x70 ;
  assign n669 = n668 ^ n666 ;
  assign n672 = n442 & ~n545 ;
  assign n673 = n672 ^ x69 ;
  assign n670 = n300 & ~n403 ;
  assign n671 = n670 ^ x5 ;
  assign n674 = n673 ^ n671 ;
  assign n677 = n278 & ~n403 ;
  assign n678 = n677 ^ x4 ;
  assign n675 = n420 & ~n545 ;
  assign n676 = n675 ^ x68 ;
  assign n679 = n678 ^ n676 ;
  assign n682 = n434 & ~n545 ;
  assign n683 = n682 ^ x67 ;
  assign n680 = n292 & ~n403 ;
  assign n681 = n680 ^ x3 ;
  assign n684 = n683 ^ n681 ;
  assign n687 = n421 & ~n545 ;
  assign n688 = n687 ^ x66 ;
  assign n685 = n279 & ~n403 ;
  assign n686 = n685 ^ x2 ;
  assign n689 = n688 ^ n686 ;
  assign n692 = n284 & ~n403 ;
  assign n693 = n692 ^ x1 ;
  assign n690 = n426 & ~n545 ;
  assign n691 = n690 ^ x65 ;
  assign n694 = n693 ^ n691 ;
  assign n695 = x96 ^ x64 ;
  assign n696 = ~n545 & n695 ;
  assign n697 = n696 ^ x64 ;
  assign n698 = x32 ^ x0 ;
  assign n699 = ~n403 & n698 ;
  assign n700 = n699 ^ x0 ;
  assign n701 = ~n697 & n700 ;
  assign n702 = n701 ^ n691 ;
  assign n703 = ~n694 & ~n702 ;
  assign n704 = n703 ^ n691 ;
  assign n705 = n704 ^ n686 ;
  assign n706 = ~n689 & ~n705 ;
  assign n707 = n706 ^ n686 ;
  assign n708 = n707 ^ n681 ;
  assign n709 = ~n684 & n708 ;
  assign n710 = n709 ^ n681 ;
  assign n711 = n710 ^ n678 ;
  assign n712 = ~n679 & n711 ;
  assign n713 = n712 ^ n678 ;
  assign n714 = n713 ^ n671 ;
  assign n715 = ~n674 & n714 ;
  assign n716 = n715 ^ n671 ;
  assign n717 = n716 ^ n668 ;
  assign n718 = ~n669 & n717 ;
  assign n719 = n718 ^ n668 ;
  assign n720 = n719 ^ n661 ;
  assign n721 = ~n664 & n720 ;
  assign n722 = n721 ^ n661 ;
  assign n723 = n722 ^ n658 ;
  assign n724 = ~n659 & n723 ;
  assign n725 = n724 ^ n658 ;
  assign n726 = n725 ^ n651 ;
  assign n727 = ~n654 & n726 ;
  assign n728 = n727 ^ n651 ;
  assign n729 = n728 ^ n648 ;
  assign n730 = ~n649 & n729 ;
  assign n731 = n730 ^ n648 ;
  assign n732 = n731 ^ n641 ;
  assign n733 = ~n644 & n732 ;
  assign n734 = n733 ^ n641 ;
  assign n735 = n734 ^ n638 ;
  assign n736 = ~n639 & n735 ;
  assign n737 = n736 ^ n638 ;
  assign n738 = n737 ^ n631 ;
  assign n739 = ~n634 & n738 ;
  assign n740 = n739 ^ n631 ;
  assign n741 = n740 ^ n628 ;
  assign n742 = ~n629 & n741 ;
  assign n743 = n742 ^ n628 ;
  assign n744 = n743 ^ n621 ;
  assign n745 = ~n624 & n744 ;
  assign n746 = n745 ^ n621 ;
  assign n747 = n746 ^ n618 ;
  assign n748 = ~n619 & n747 ;
  assign n749 = n748 ^ n618 ;
  assign n750 = n749 ^ n611 ;
  assign n751 = ~n614 & n750 ;
  assign n752 = n751 ^ n611 ;
  assign n753 = n752 ^ n608 ;
  assign n754 = ~n609 & n753 ;
  assign n755 = n754 ^ n608 ;
  assign n756 = n755 ^ n601 ;
  assign n757 = ~n604 & n756 ;
  assign n758 = n757 ^ n601 ;
  assign n759 = n758 ^ n598 ;
  assign n760 = ~n599 & n759 ;
  assign n761 = n760 ^ n598 ;
  assign n762 = n761 ^ n591 ;
  assign n763 = ~n594 & n762 ;
  assign n764 = n763 ^ n591 ;
  assign n765 = n764 ^ n588 ;
  assign n766 = ~n589 & n765 ;
  assign n767 = n766 ^ n588 ;
  assign n768 = n767 ^ n581 ;
  assign n769 = ~n584 & n768 ;
  assign n770 = n769 ^ n581 ;
  assign n771 = n770 ^ n578 ;
  assign n772 = ~n579 & ~n771 ;
  assign n773 = n772 ^ n578 ;
  assign n774 = n773 ^ n571 ;
  assign n775 = ~n574 & ~n774 ;
  assign n776 = n775 ^ n571 ;
  assign n777 = n776 ^ n568 ;
  assign n778 = ~n569 & n777 ;
  assign n779 = n778 ^ n568 ;
  assign n780 = n779 ^ n561 ;
  assign n781 = ~n564 & n780 ;
  assign n782 = n781 ^ n561 ;
  assign n783 = n782 ^ n556 ;
  assign n784 = ~n559 & ~n783 ;
  assign n785 = n784 ^ n556 ;
  assign n786 = n785 ^ n551 ;
  assign n787 = ~n554 & n786 ;
  assign n788 = n787 ^ n553 ;
  assign n789 = n788 ^ n405 ;
  assign n790 = ~n548 & n789 ;
  assign n791 = n790 ^ n547 ;
  assign n792 = n791 ^ n258 ;
  assign n793 = ~n549 & n792 ;
  assign n794 = n793 ^ n257 ;
  assign n795 = n548 & ~n794 ;
  assign n796 = n795 ^ n547 ;
  assign n1330 = n1329 ^ n796 ;
  assign n1333 = n1087 & n1327 ;
  assign n1334 = n1333 ^ n1084 ;
  assign n1331 = n554 & n794 ;
  assign n1332 = n1331 ^ n551 ;
  assign n1335 = n1334 ^ n1332 ;
  assign n1338 = n559 & ~n794 ;
  assign n1339 = n1338 ^ n556 ;
  assign n1336 = n1092 & n1327 ;
  assign n1337 = n1336 ^ n1089 ;
  assign n1340 = n1339 ^ n1337 ;
  assign n1343 = n1097 & ~n1327 ;
  assign n1344 = n1343 ^ n1094 ;
  assign n1341 = n564 & n794 ;
  assign n1342 = n1341 ^ n561 ;
  assign n1345 = n1344 ^ n1342 ;
  assign n1348 = n1102 & n1327 ;
  assign n1349 = n1348 ^ n1101 ;
  assign n1346 = n569 & n794 ;
  assign n1347 = n1346 ^ n568 ;
  assign n1350 = n1349 ^ n1347 ;
  assign n1353 = n574 & ~n794 ;
  assign n1354 = n1353 ^ n573 ;
  assign n1351 = n1107 & ~n1327 ;
  assign n1352 = n1351 ^ n1106 ;
  assign n1355 = n1354 ^ n1352 ;
  assign n1358 = n1112 & ~n1327 ;
  assign n1359 = n1358 ^ n1109 ;
  assign n1356 = n579 & n794 ;
  assign n1357 = n1356 ^ n576 ;
  assign n1360 = n1359 ^ n1357 ;
  assign n1363 = n1117 & n1327 ;
  assign n1364 = n1363 ^ n1114 ;
  assign n1361 = n584 & n794 ;
  assign n1362 = n1361 ^ n581 ;
  assign n1365 = n1364 ^ n1362 ;
  assign n1368 = n1122 & n1327 ;
  assign n1369 = n1368 ^ n1121 ;
  assign n1366 = n589 & n794 ;
  assign n1367 = n1366 ^ n588 ;
  assign n1370 = n1369 ^ n1367 ;
  assign n1373 = n594 & ~n794 ;
  assign n1374 = n1373 ^ n593 ;
  assign n1371 = n1127 & ~n1327 ;
  assign n1372 = n1371 ^ n1126 ;
  assign n1375 = n1374 ^ n1372 ;
  assign n1378 = n599 & ~n794 ;
  assign n1379 = n1378 ^ n596 ;
  assign n1376 = n1132 & ~n1327 ;
  assign n1377 = n1376 ^ n1129 ;
  assign n1380 = n1379 ^ n1377 ;
  assign n1383 = n1137 & n1327 ;
  assign n1384 = n1383 ^ n1134 ;
  assign n1381 = n604 & n794 ;
  assign n1382 = n1381 ^ n601 ;
  assign n1385 = n1384 ^ n1382 ;
  assign n1388 = n1142 & n1327 ;
  assign n1389 = n1388 ^ n1141 ;
  assign n1386 = n609 & n794 ;
  assign n1387 = n1386 ^ n608 ;
  assign n1390 = n1389 ^ n1387 ;
  assign n1393 = n614 & ~n794 ;
  assign n1394 = n1393 ^ n613 ;
  assign n1391 = n1147 & ~n1327 ;
  assign n1392 = n1391 ^ n1146 ;
  assign n1395 = n1394 ^ n1392 ;
  assign n1398 = n619 & ~n794 ;
  assign n1399 = n1398 ^ n616 ;
  assign n1396 = n1152 & ~n1327 ;
  assign n1397 = n1396 ^ n1149 ;
  assign n1400 = n1399 ^ n1397 ;
  assign n1403 = n1157 & n1327 ;
  assign n1404 = n1403 ^ n1154 ;
  assign n1401 = n624 & n794 ;
  assign n1402 = n1401 ^ n621 ;
  assign n1405 = n1404 ^ n1402 ;
  assign n1408 = n1162 & n1327 ;
  assign n1409 = n1408 ^ n1161 ;
  assign n1406 = n629 & n794 ;
  assign n1407 = n1406 ^ n628 ;
  assign n1410 = n1409 ^ n1407 ;
  assign n1413 = n634 & ~n794 ;
  assign n1414 = n1413 ^ n633 ;
  assign n1411 = n1167 & ~n1327 ;
  assign n1412 = n1411 ^ n1166 ;
  assign n1415 = n1414 ^ n1412 ;
  assign n1418 = n639 & ~n794 ;
  assign n1419 = n1418 ^ n636 ;
  assign n1416 = n1172 & ~n1327 ;
  assign n1417 = n1416 ^ n1169 ;
  assign n1420 = n1419 ^ n1417 ;
  assign n1423 = n1177 & n1327 ;
  assign n1424 = n1423 ^ n1174 ;
  assign n1421 = n644 & n794 ;
  assign n1422 = n1421 ^ n641 ;
  assign n1425 = n1424 ^ n1422 ;
  assign n1428 = n1182 & n1327 ;
  assign n1429 = n1428 ^ n1181 ;
  assign n1426 = n649 & n794 ;
  assign n1427 = n1426 ^ n648 ;
  assign n1430 = n1429 ^ n1427 ;
  assign n1433 = n654 & ~n794 ;
  assign n1434 = n1433 ^ n653 ;
  assign n1431 = n1187 & ~n1327 ;
  assign n1432 = n1431 ^ n1186 ;
  assign n1435 = n1434 ^ n1432 ;
  assign n1438 = n659 & ~n794 ;
  assign n1439 = n1438 ^ n656 ;
  assign n1436 = n1192 & ~n1327 ;
  assign n1437 = n1436 ^ n1189 ;
  assign n1440 = n1439 ^ n1437 ;
  assign n1443 = n1197 & n1327 ;
  assign n1444 = n1443 ^ n1194 ;
  assign n1441 = n664 & n794 ;
  assign n1442 = n1441 ^ n661 ;
  assign n1445 = n1444 ^ n1442 ;
  assign n1448 = n669 & n794 ;
  assign n1449 = n1448 ^ n668 ;
  assign n1446 = n1202 & ~n1327 ;
  assign n1447 = n1446 ^ n1201 ;
  assign n1450 = n1449 ^ n1447 ;
  assign n1453 = n674 & ~n794 ;
  assign n1454 = n1453 ^ n673 ;
  assign n1451 = n1207 & ~n1327 ;
  assign n1452 = n1451 ^ n1206 ;
  assign n1455 = n1454 ^ n1452 ;
  assign n1458 = n679 & ~n794 ;
  assign n1459 = n1458 ^ n676 ;
  assign n1456 = n1212 & n1327 ;
  assign n1457 = n1456 ^ n1209 ;
  assign n1460 = n1459 ^ n1457 ;
  assign n1463 = n1217 & ~n1327 ;
  assign n1464 = n1463 ^ n1214 ;
  assign n1461 = n684 & n794 ;
  assign n1462 = n1461 ^ n681 ;
  assign n1465 = n1464 ^ n1462 ;
  assign n1468 = n1222 & ~n1327 ;
  assign n1469 = n1468 ^ n1221 ;
  assign n1466 = n689 & ~n794 ;
  assign n1467 = n1466 ^ n688 ;
  assign n1470 = n1469 ^ n1467 ;
  assign n1473 = n694 & n794 ;
  assign n1474 = n1473 ^ n693 ;
  assign n1471 = n1227 & n1327 ;
  assign n1472 = n1471 ^ n1226 ;
  assign n1475 = n1474 ^ n1472 ;
  assign n1476 = n1233 ^ n1230 ;
  assign n1477 = ~n1327 & n1476 ;
  assign n1478 = n1477 ^ n1230 ;
  assign n1479 = n700 ^ n697 ;
  assign n1480 = ~n794 & n1479 ;
  assign n1481 = n1480 ^ n697 ;
  assign n1482 = ~n1478 & n1481 ;
  assign n1483 = n1482 ^ n1472 ;
  assign n1484 = ~n1475 & ~n1483 ;
  assign n1485 = n1484 ^ n1472 ;
  assign n1486 = n1485 ^ n1469 ;
  assign n1487 = ~n1470 & n1486 ;
  assign n1488 = n1487 ^ n1469 ;
  assign n1489 = n1488 ^ n1462 ;
  assign n1490 = ~n1465 & ~n1489 ;
  assign n1491 = n1490 ^ n1462 ;
  assign n1492 = n1491 ^ n1459 ;
  assign n1493 = ~n1460 & n1492 ;
  assign n1494 = n1493 ^ n1459 ;
  assign n1495 = n1494 ^ n1452 ;
  assign n1496 = ~n1455 & ~n1495 ;
  assign n1497 = n1496 ^ n1452 ;
  assign n1498 = n1497 ^ n1449 ;
  assign n1499 = ~n1450 & ~n1498 ;
  assign n1500 = n1499 ^ n1449 ;
  assign n1501 = n1500 ^ n1442 ;
  assign n1502 = ~n1445 & n1501 ;
  assign n1503 = n1502 ^ n1442 ;
  assign n1504 = n1503 ^ n1439 ;
  assign n1505 = ~n1440 & n1504 ;
  assign n1506 = n1505 ^ n1439 ;
  assign n1507 = n1506 ^ n1432 ;
  assign n1508 = ~n1435 & ~n1507 ;
  assign n1509 = n1508 ^ n1432 ;
  assign n1510 = n1509 ^ n1429 ;
  assign n1511 = ~n1430 & n1510 ;
  assign n1512 = n1511 ^ n1429 ;
  assign n1513 = n1512 ^ n1422 ;
  assign n1514 = ~n1425 & ~n1513 ;
  assign n1515 = n1514 ^ n1422 ;
  assign n1516 = n1515 ^ n1419 ;
  assign n1517 = ~n1420 & n1516 ;
  assign n1518 = n1517 ^ n1419 ;
  assign n1519 = n1518 ^ n1412 ;
  assign n1520 = ~n1415 & ~n1519 ;
  assign n1521 = n1520 ^ n1412 ;
  assign n1522 = n1521 ^ n1409 ;
  assign n1523 = ~n1410 & n1522 ;
  assign n1524 = n1523 ^ n1409 ;
  assign n1525 = n1524 ^ n1402 ;
  assign n1526 = ~n1405 & ~n1525 ;
  assign n1527 = n1526 ^ n1402 ;
  assign n1528 = n1527 ^ n1399 ;
  assign n1529 = ~n1400 & n1528 ;
  assign n1530 = n1529 ^ n1399 ;
  assign n1531 = n1530 ^ n1392 ;
  assign n1532 = ~n1395 & ~n1531 ;
  assign n1533 = n1532 ^ n1392 ;
  assign n1534 = n1533 ^ n1389 ;
  assign n1535 = ~n1390 & n1534 ;
  assign n1536 = n1535 ^ n1389 ;
  assign n1537 = n1536 ^ n1382 ;
  assign n1538 = ~n1385 & ~n1537 ;
  assign n1539 = n1538 ^ n1382 ;
  assign n1540 = n1539 ^ n1379 ;
  assign n1541 = ~n1380 & n1540 ;
  assign n1542 = n1541 ^ n1379 ;
  assign n1543 = n1542 ^ n1372 ;
  assign n1544 = ~n1375 & ~n1543 ;
  assign n1545 = n1544 ^ n1372 ;
  assign n1546 = n1545 ^ n1369 ;
  assign n1547 = ~n1370 & n1546 ;
  assign n1548 = n1547 ^ n1369 ;
  assign n1549 = n1548 ^ n1362 ;
  assign n1550 = ~n1365 & ~n1549 ;
  assign n1551 = n1550 ^ n1362 ;
  assign n1552 = n1551 ^ n1359 ;
  assign n1553 = ~n1360 & ~n1552 ;
  assign n1554 = n1553 ^ n1359 ;
  assign n1555 = n1554 ^ n1352 ;
  assign n1556 = ~n1355 & n1555 ;
  assign n1557 = n1556 ^ n1352 ;
  assign n1558 = n1557 ^ n1349 ;
  assign n1559 = ~n1350 & n1558 ;
  assign n1560 = n1559 ^ n1349 ;
  assign n1561 = n1560 ^ n1342 ;
  assign n1562 = ~n1345 & ~n1561 ;
  assign n1563 = n1562 ^ n1342 ;
  assign n1564 = n1563 ^ n1339 ;
  assign n1565 = ~n1340 & n1564 ;
  assign n1566 = n1565 ^ n1339 ;
  assign n1567 = n1566 ^ n1334 ;
  assign n1568 = ~n1335 & ~n1567 ;
  assign n1569 = n1568 ^ n1334 ;
  assign n1570 = n1569 ^ n1329 ;
  assign n1571 = ~n1330 & ~n1570 ;
  assign n1572 = n1571 ^ n796 ;
  assign n1573 = n1572 ^ n259 ;
  assign n1574 = ~n263 & n1573 ;
  assign n1575 = n1574 ^ n262 ;
  assign n1576 = n1327 ^ n794 ;
  assign n1577 = ~n1575 & n1576 ;
  assign n1578 = n1577 ^ n794 ;
  assign n1582 = n1078 & ~n1578 ;
  assign n1583 = n936 & n1327 ;
  assign n1584 = ~n1582 & ~n1583 ;
  assign n1579 = n403 & ~n1578 ;
  assign n1580 = n545 & n794 ;
  assign n1581 = ~n1579 & ~n1580 ;
  assign n1585 = n1584 ^ n1581 ;
  assign n1586 = n1575 & n1585 ;
  assign n1587 = n1586 ^ n1584 ;
  assign n1588 = n1481 ^ n1478 ;
  assign n1589 = n1575 & n1588 ;
  assign n1590 = n1589 ^ n1478 ;
  assign n1591 = n1475 & ~n1575 ;
  assign n1592 = n1591 ^ n1474 ;
  assign n1593 = n1470 & n1575 ;
  assign n1594 = n1593 ^ n1469 ;
  assign n1595 = n1465 & ~n1575 ;
  assign n1596 = n1595 ^ n1462 ;
  assign n1597 = n1460 & n1575 ;
  assign n1598 = n1597 ^ n1457 ;
  assign n1599 = n1455 & ~n1575 ;
  assign n1600 = n1599 ^ n1454 ;
  assign n1601 = n1450 & ~n1575 ;
  assign n1602 = n1601 ^ n1449 ;
  assign n1603 = n1445 & ~n1575 ;
  assign n1604 = n1603 ^ n1442 ;
  assign n1605 = n1440 & n1575 ;
  assign n1606 = n1605 ^ n1437 ;
  assign n1607 = n1435 & ~n1575 ;
  assign n1608 = n1607 ^ n1434 ;
  assign n1609 = n1430 & n1575 ;
  assign n1610 = n1609 ^ n1429 ;
  assign n1611 = n1425 & ~n1575 ;
  assign n1612 = n1611 ^ n1422 ;
  assign n1613 = n1420 & n1575 ;
  assign n1614 = n1613 ^ n1417 ;
  assign n1615 = n1415 & ~n1575 ;
  assign n1616 = n1615 ^ n1414 ;
  assign n1617 = n1410 & n1575 ;
  assign n1618 = n1617 ^ n1409 ;
  assign n1619 = n1405 & ~n1575 ;
  assign n1620 = n1619 ^ n1402 ;
  assign n1621 = n1400 & n1575 ;
  assign n1622 = n1621 ^ n1397 ;
  assign n1623 = n1395 & ~n1575 ;
  assign n1624 = n1623 ^ n1394 ;
  assign n1625 = n1390 & n1575 ;
  assign n1626 = n1625 ^ n1389 ;
  assign n1627 = n1385 & ~n1575 ;
  assign n1628 = n1627 ^ n1382 ;
  assign n1629 = n1380 & n1575 ;
  assign n1630 = n1629 ^ n1377 ;
  assign n1631 = n1375 & ~n1575 ;
  assign n1632 = n1631 ^ n1374 ;
  assign n1633 = n1370 & n1575 ;
  assign n1634 = n1633 ^ n1369 ;
  assign n1635 = n1365 & ~n1575 ;
  assign n1636 = n1635 ^ n1362 ;
  assign n1637 = n1360 & ~n1575 ;
  assign n1638 = n1637 ^ n1357 ;
  assign n1639 = n1355 & ~n1575 ;
  assign n1640 = n1639 ^ n1354 ;
  assign n1641 = n1350 & n1575 ;
  assign n1642 = n1641 ^ n1349 ;
  assign n1643 = n1345 & ~n1575 ;
  assign n1644 = n1643 ^ n1342 ;
  assign n1645 = n1340 & n1575 ;
  assign n1646 = n1645 ^ n1337 ;
  assign n1647 = n1335 & n1575 ;
  assign n1648 = n1647 ^ n1334 ;
  assign n1649 = n1330 & n1575 ;
  assign n1650 = n1649 ^ n1329 ;
  assign n1651 = n259 & n262 ;
  assign y0 = n1587 ;
  assign y1 = n1578 ;
  assign y2 = ~n1575 ;
  assign y3 = n1590 ;
  assign y4 = n1592 ;
  assign y5 = n1594 ;
  assign y6 = n1596 ;
  assign y7 = n1598 ;
  assign y8 = n1600 ;
  assign y9 = n1602 ;
  assign y10 = n1604 ;
  assign y11 = n1606 ;
  assign y12 = n1608 ;
  assign y13 = n1610 ;
  assign y14 = n1612 ;
  assign y15 = n1614 ;
  assign y16 = n1616 ;
  assign y17 = n1618 ;
  assign y18 = n1620 ;
  assign y19 = n1622 ;
  assign y20 = n1624 ;
  assign y21 = n1626 ;
  assign y22 = n1628 ;
  assign y23 = n1630 ;
  assign y24 = n1632 ;
  assign y25 = n1634 ;
  assign y26 = n1636 ;
  assign y27 = n1638 ;
  assign y28 = n1640 ;
  assign y29 = n1642 ;
  assign y30 = n1644 ;
  assign y31 = n1646 ;
  assign y32 = n1648 ;
  assign y33 = n1650 ;
  assign y34 = ~n1651 ;
endmodule
