// Benchmark "bitonic_sort_inc" written by ABC on Wed Jul  9 17:56:52 2025

module bitonic_sort_inc_4 ( 
    \in_array[0] , \in_array[1] , \in_array[2] , \in_array[3] ,
    \in_array[4] , \in_array[5] , \in_array[6] , \in_array[7] ,
    \in_array[8] , \in_array[9] , \in_array[10] , \in_array[11] ,
    \in_array[12] , \in_array[13] , \in_array[14] , \in_array[15] ,
    \in_array[16] , \in_array[17] , \in_array[18] , \in_array[19] ,
    \in_array[20] , \in_array[21] , \in_array[22] , \in_array[23] ,
    \in_array[24] , \in_array[25] , \in_array[26] , \in_array[27] ,
    \in_array[28] , \in_array[29] , \in_array[30] , \in_array[31] ,
    \out_array[0] , \out_array[1] , \out_array[2] , \out_array[3] ,
    \out_array[4] , \out_array[5] , \out_array[6] , \out_array[7] ,
    \out_array[8] , \out_array[9] , \out_array[10] , \out_array[11] ,
    \out_array[12] , \out_array[13] , \out_array[14] , \out_array[15] ,
    \out_array[16] , \out_array[17] , \out_array[18] , \out_array[19] ,
    \out_array[20] , \out_array[21] , \out_array[22] , \out_array[23] ,
    \out_array[24] , \out_array[25] , \out_array[26] , \out_array[27] ,
    \out_array[28] , \out_array[29] , \out_array[30] , \out_array[31]   );
  input  \in_array[0] , \in_array[1] , \in_array[2] , \in_array[3] ,
    \in_array[4] , \in_array[5] , \in_array[6] , \in_array[7] ,
    \in_array[8] , \in_array[9] , \in_array[10] , \in_array[11] ,
    \in_array[12] , \in_array[13] , \in_array[14] , \in_array[15] ,
    \in_array[16] , \in_array[17] , \in_array[18] , \in_array[19] ,
    \in_array[20] , \in_array[21] , \in_array[22] , \in_array[23] ,
    \in_array[24] , \in_array[25] , \in_array[26] , \in_array[27] ,
    \in_array[28] , \in_array[29] , \in_array[30] , \in_array[31] ;
  output \out_array[0] , \out_array[1] , \out_array[2] , \out_array[3] ,
    \out_array[4] , \out_array[5] , \out_array[6] , \out_array[7] ,
    \out_array[8] , \out_array[9] , \out_array[10] , \out_array[11] ,
    \out_array[12] , \out_array[13] , \out_array[14] , \out_array[15] ,
    \out_array[16] , \out_array[17] , \out_array[18] , \out_array[19] ,
    \out_array[20] , \out_array[21] , \out_array[22] , \out_array[23] ,
    \out_array[24] , \out_array[25] , \out_array[26] , \out_array[27] ,
    \out_array[28] , \out_array[29] , \out_array[30] , \out_array[31] ;
  wire new__0550_, new__0561_, new__0569_, new__0576_, new__0587_,
    new__0598_, new__0608_, new__0615_, new__0622_, new__0633_, new__0644_,
    new__0655_, new__0666_, new__0677_, new__0688_, new__0699_, new__0710_,
    new__0721_, new__0730_, new__0737_, new__0747_, new__0758_, new__0769_,
    new__0776_, new__0783_, new__0784_, new__0785_, new__0786_, new__0787_,
    new__0788_, new__0789_, new__0790_, new__0791_, new__0792_, new__0793_,
    new__0000_, new__0001_, new__0002_, new__0003_, new__0004_, new__0005_,
    new__0006_, new__0007__neg, new__0007_, new__0008_, new__0009_,
    new__0010_, new__0011_, new__0012_, new__0013_, new__0014_, new__0015_,
    new__0016_, new__0017_, new__0018_, new__0019_, new__0020_, new__0021_,
    new__0022_, new__0023_, new__0024_, new__0025_, new__0026_, new__0027_,
    new__0028_, new__0029_, new__0030_, new__0031_, new__0032_, new__0033_,
    new__0034_, new__0035_, new__0036_, new__0037_, new__0038_, new__0039_,
    new__0040_, new__0041_, new__0042_, new__0043_, new__0044_, new__0045_,
    new__0046_, new__0047_, new__0048__neg, new__0048_, new__0049_,
    new__0050_, new__0051_, new__0052_, new__0053_, new__0054_, new__0055_,
    new__0056_, new__0057_, new__0058_, new__0059_, new__0060_, new__0061_,
    new__0062_, new__0063_, new__0064_, new__0065_, new__0066_, new__0067_,
    new__0068_, new__0069_, new__0070_, new__0071__neg, new__0071_,
    new__0072__neg, new__0072_, new__0073_, new__0074_, new__0075_,
    new__0076__neg, new__0076_, new__0077_, new__0078_, new__0079_,
    new__0080__neg, new__0080_, new__0081_, new__0082_, new__0083_,
    new__0084_, new__0085__neg, new__0085_, new__0086_, new__0087_,
    new__0088_, new__0089_, new__0090_, new__0091_, new__0092_, new__0093_,
    new__0094_, new__0095_, new__0096_, new__0097__neg, new__0097_,
    new__0098_, new__0099_, new__0100_, new__0101_, new__0102__neg,
    new__0102_, new__0103_, new__0104_, new__0105_, new__0106_, new__0107_,
    new__0108_, new__0109_, new__0110_, new__0111_, new__0112_, new__0113_,
    new__0114_, new__0115_, new__0116_, new__0117_, new__0118_, new__0119_,
    new__0120_, new__0121_, new__0122_, new__0123_, new__0124_, new__0125_,
    new__0126_, new__0127_, new__0128_, new__0129_, new__0130_, new__0131_,
    new__0132_, new__0133_, new__0134_, new__0135_, new__0136_, new__0137_,
    new__0138_, new__0139_, new__0140_, new__0141_, new__0142_, new__0143_,
    new__0144_, new__0145_, new__0146_, new__0147_, new__0148_, new__0149_,
    new__0150_, new__0151_, new__0152_, new__0153__neg, new__0153_,
    new__0154_, new__0155_, new__0156_, new__0157_, new__0158_, new__0159_,
    new__0160_, new__0161_, new__0162_, new__0163_, new__0164_, new__0165_,
    new__0166_, new__0167_, new__0168_, new__0169_, new__0170_, new__0171_,
    new__0172_, new__0173_, new__0174_, new__0175_, new__0176_, new__0177_,
    new__0178_, new__0179_, new__0180_, new__0181_, new__0182_, new__0183_,
    new__0184_, new__0185_, new__0186_, new__0187_, new__0188_, new__0189_,
    new__0190_, new__0191_, new__0192__neg, new__0192_, new__0193_,
    new__0194_, new__0195_, new__0196_, new__0197_, new__0198_, new__0199_,
    new__0200_, new__0201_, new__0202_, new__0203_, new__0204_, new__0205_,
    new__0206_, new__0207_, new__0208_, new__0209_, new__0210_, new__0211_,
    new__0212_, new__0213_, new__0214_, new__0215_, new__0216__neg,
    new__0216_, new__0217__neg, new__0217_, new__0218_, new__0219_,
    new__0220_, new__0221__neg, new__0221_, new__0222_, new__0223_,
    new__0224_, new__0225__neg, new__0225_, new__0226_, new__0227_,
    new__0228_, new__0229_, new__0230__neg, new__0230_, new__0231_,
    new__0232_, new__0233_, new__0234_, new__0235_, new__0236_, new__0237_,
    new__0238_, new__0239_, new__0240__neg, new__0240_, new__0241_,
    new__0242_, new__0243_, new__0244_, new__0245_, new__0246__neg,
    new__0246_, new__0247_, new__0248_, new__0249_, new__0250_, new__0251_,
    new__0252_, new__0253_, new__0254__neg, new__0254_, new__0255__neg,
    new__0255_, new__0256_, new__0257_, new__0258_, new__0259__neg,
    new__0259_, new__0260_, new__0261_, new__0262_, new__0263__neg,
    new__0263_, new__0264_, new__0265_, new__0266_, new__0267_,
    new__0268__neg, new__0268_, new__0269_, new__0270_, new__0271_,
    new__0272_, new__0273_, new__0274_, new__0275_, new__0276_, new__0277_,
    new__0278_, new__0279_, new__0280_, new__0281_, new__0282_, new__0283_,
    new__0284_, new__0285_, new__0286_, new__0287_, new__0288_, new__0289_,
    new__0290_, new__0291_, new__0292_, new__0293_, new__0294_,
    new__0295__neg, new__0295_, new__0296_, new__0297_, new__0298_,
    new__0299_, new__0300_, new__0301_, new__0302_, new__0303_, new__0304_,
    new__0305_, new__0306_, new__0307_, new__0308_, new__0309_, new__0310_,
    new__0311_, new__0312_, new__0313_, new__0314_, new__0315_, new__0316_,
    new__0317_, new__0318_, new__0319_, new__0320_, new__0321_, new__0322_,
    new__0323_, new__0324_, new__0325__neg, new__0325_, new__0326_,
    new__0327_, new__0328_, new__0329_, new__0330_, new__0331_, new__0332_,
    new__0333_, new__0334_, new__0335_, new__0336_, new__0337_, new__0338_,
    new__0339_, new__0340_, new__0341_, new__0342_, new__0343_, new__0344_,
    new__0345_, new__0346_, new__0347_, new__0348_, new__0349_, new__0350_,
    new__0351_, new__0352__neg, new__0352_, new__0353__neg, new__0353_,
    new__0354_, new__0355_, new__0356_, new__0357__neg, new__0357_,
    new__0358_, new__0359_, new__0360_, new__0361__neg, new__0361_,
    new__0362_, new__0363_, new__0364_, new__0365_, new__0366__neg,
    new__0366_, new__0367_, new__0368_, new__0369_, new__0370_, new__0371_,
    new__0372_, new__0373_, new__0374_, new__0375_, new__0376_, new__0377_,
    new__0378_, new__0379_, new__0380_, new__0381_, new__0382_, new__0383_,
    new__0384_, new__0385_, new__0386_, new__0387_, new__0388_, new__0389_,
    new__0390__neg, new__0390_, new__0391__neg, new__0391_, new__0392_,
    new__0393_, new__0394_, new__0395__neg, new__0395_, new__0396_,
    new__0397_, new__0398_, new__0399__neg, new__0399_, new__0400_,
    new__0401_, new__0402_, new__0403_, new__0404__neg, new__0404_,
    new__0405_, new__0406_, new__0407_, new__0408_, new__0409_, new__0410_,
    new__0411_, new__0412_, new__0413_, new__0414_, new__0415_, new__0416_,
    new__0417_, new__0418_, new__0419_, new__0420_, new__0421_, new__0422_,
    new__0423_, new__0424_, new__0425_, new__0426_, new__0427_, new__0428_,
    new__0429_, new__0430_, new__0431_, new__0432__neg, new__0432_,
    new__0433_, new__0434_, new__0435_, new__0436_, new__0437_, new__0438_,
    new__0439_, new__0440_, new__0441_, new__0442_, new__0443_, new__0444_,
    new__0445_, new__0446_, new__0447_, new__0448_, new__0449_, new__0450_,
    new__0451_, new__0452_, new__0453_, new__0454_, new__0455_, new__0456_,
    new__0457_, new__0458_, new__0459_, new__0460_, new__0461_,
    new__0462__neg, new__0462_, new__0463_, new__0464_, new__0465_,
    new__0466_, new__0467_, new__0468_, new__0469_, new__0470_, new__0471_,
    new__0472_, new__0473_, new__0474_, new__0475_, new__0476_, new__0477_,
    new__0478_, new__0479_, new__0480_, new__0481_, new__0482_, new__0483_,
    new__0484_, new__0485_, new__0486_, new__0487_, new__0488__neg,
    new__0488_, new__0489__neg, new__0489_, new__0490_, new__0491_,
    new__0492_, new__0493__neg, new__0493_, new__0494_, new__0495_,
    new__0496_, new__0497__neg, new__0497_, new__0498_, new__0499_,
    new__0500_, new__0501_, new__0502__neg, new__0502_, new__0503_,
    new__0504_, new__0505_, new__0506_, new__0507_, new__0508_, new__0509_,
    new__0510_, new__0511_, new__0512_, new__0513_, new__0514_, new__0515_,
    new__0516_, new__0517_, new__0518_, new__0519_, new__0520_, new__0521_,
    new__0522_, new__0523_, new__0524_, new__0525_, new__0526__neg,
    new__0526_, new__0527_, new__0528__neg, new__0528_, new__0529_,
    new__0530_, new__0531__neg, new__0531_, new__0532_, new__0533_,
    new__0534_, new__0535_, new__0536__neg, new__0536_, new__0537_,
    new__0538_, new__0539_, new__0540__neg, new__0540_, new__0541_,
    new__0542_, new__0543_, new__0544_, new__0545_, new__0546_, new__0547_,
    new__0548_, new__0549_, new__0551_, new__0552_, new__0553_, new__0554_,
    new__0555_, new__0556_, new__0557_, new__0558_, new__0559_, new__0560_,
    new__0562_, new__0563_, new__0564_, new__0565__neg, new__0565_,
    new__0566_, new__0567__neg, new__0567_, new__0568_, new__0570_,
    new__0571_, new__0572_, new__0573_, new__0574_, new__0575_, new__0577_,
    new__0578_, new__0579_, new__0580__neg, new__0580_, new__0581_,
    new__0582_, new__0583_, new__0584_, new__0585_, new__0586_, new__0588_,
    new__0589_, new__0590_, new__0591_, new__0592_, new__0593_, new__0594_,
    new__0595_, new__0596_, new__0597_, new__0599_, new__0600_, new__0601_,
    new__0602_, new__0603_, new__0604_, new__0605_, new__0606_,
    new__0607__neg, new__0607_, new__0609_, new__0610__neg, new__0610_,
    new__0611_, new__0612_, new__0613_, new__0614_, new__0616_, new__0617_,
    new__0618_, new__0619_, new__0620_, new__0621_, new__0623_, new__0624_,
    new__0625__neg, new__0625_, new__0626_, new__0627_, new__0628_,
    new__0629_, new__0630_, new__0631_, new__0632_, new__0634_, new__0635_,
    new__0636_, new__0637_, new__0638_, new__0639_, new__0640_, new__0641_,
    new__0642_, new__0643_, new__0645_, new__0646_, new__0647_, new__0648_,
    new__0649_, new__0650_, new__0651_, new__0652_, new__0653_, new__0654_,
    new__0656_, new__0657_, new__0658__neg, new__0658_, new__0659_,
    new__0660_, new__0661_, new__0662_, new__0663_, new__0664_, new__0665_,
    new__0667_, new__0668_, new__0669_, new__0670_, new__0671_, new__0672_,
    new__0673_, new__0674_, new__0675_, new__0676_, new__0678_, new__0679_,
    new__0680_, new__0681_, new__0682_, new__0683_, new__0684_, new__0685_,
    new__0686__neg, new__0686_, new__0687_, new__0689__neg, new__0689_,
    new__0690_, new__0691_, new__0692__neg, new__0692_, new__0693_,
    new__0694_, new__0695_, new__0696_, new__0697__neg, new__0697_,
    new__0698_, new__0700_, new__0701_, new__0702__neg, new__0702_,
    new__0703_, new__0704_, new__0705_, new__0706_, new__0707_, new__0708_,
    new__0709_, new__0711_, new__0712_, new__0713_, new__0714_, new__0715_,
    new__0716_, new__0717_, new__0718_, new__0719_, new__0720_, new__0722_,
    new__0723_, new__0724_, new__0725_, new__0726_, new__0727__neg,
    new__0727_, new__0728_, new__0729__neg, new__0729_, new__0731_,
    new__0732_, new__0733_, new__0734_, new__0735_, new__0736_, new__0738_,
    new__0739_, new__0740_, new__0741_, new__0742__neg, new__0742_,
    new__0743_, new__0744_, new__0745_, new__0746_, new__0748_, new__0749_,
    new__0750_, new__0751_, new__0752_, new__0753_, new__0754_, new__0755_,
    new__0756_, new__0757_, new__0759_, new__0760_, new__0761_, new__0762_,
    new__0763_, new__0764_, new__0765_, new__0766_, new__0767_, new__0768_,
    new__0770__neg, new__0770_, new__0771_, new__0772__neg, new__0772_,
    new__0773_, new__0774_, new__0775_, new__0777_, new__0778_, new__0779_,
    new__0780_, new__0781_, new__0782_;
  assign new__0550_ = ~\in_array[6] ;
  assign new__0561_ = ~\in_array[2]  ^ ~\in_array[6] ;
  assign new__0569_ = ~\in_array[0] ;
  assign new__0576_ = \in_array[4]  & new__0569_;
  assign new__0587_ = ~\in_array[1] ;
  assign new__0598_ = ~new__0576_ ^ ~new__0587_;
  assign new__0608_ = ~new__0576_ ^ ~\in_array[5] ;
  assign new__0615_ = new__0608_ & new__0598_;
  assign new__0622_ = ~new__0615_ ^ ~new__0576_;
  assign new__0633_ = ~\in_array[2] ;
  assign new__0644_ = ~new__0622_ ^ ~new__0633_;
  assign new__0655_ = ~new__0622_ ^ ~\in_array[6] ;
  assign new__0666_ = new__0655_ & new__0644_;
  assign new__0677_ = ~new__0666_ ^ ~new__0622_;
  assign new__0688_ = ~new__0677_;
  assign new__0699_ = ~\in_array[3] ;
  assign new__0710_ = ~new__0677_ ^ ~new__0699_;
  assign new__0721_ = ~new__0677_ ^ ~\in_array[7] ;
  assign new__0730_ = new__0721_ & new__0710_;
  assign new__0737_ = ~new__0730_ ^ ~new__0688_;
  assign new__0747_ = new__0737_ & new__0561_;
  assign new__0758_ = ~new__0747_ ^ ~new__0550_;
  assign new__0769_ = ~\in_array[10]  ^ ~\in_array[14] ;
  assign new__0776_ = ~\in_array[8] ;
  assign new__0783_ = \in_array[12]  & new__0776_;
  assign new__0784_ = ~\in_array[9] ;
  assign new__0785_ = ~new__0783_ ^ ~new__0784_;
  assign new__0786_ = ~new__0783_ ^ ~\in_array[13] ;
  assign new__0787_ = new__0786_ & new__0785_;
  assign new__0788_ = ~new__0787_ ^ ~new__0783_;
  assign new__0789_ = ~\in_array[10] ;
  assign new__0790_ = ~new__0788_ ^ ~new__0789_;
  assign new__0791_ = ~new__0788_ ^ ~\in_array[14] ;
  assign new__0792_ = new__0791_ & new__0790_;
  assign new__0793_ = ~new__0792_ ^ ~new__0788_;
  assign new__0000_ = ~\in_array[11] ;
  assign new__0001_ = ~new__0793_ ^ ~new__0000_;
  assign new__0002_ = ~new__0793_ ^ ~\in_array[15] ;
  assign new__0003_ = new__0002_ & new__0001_;
  assign new__0004_ = ~new__0003_ ^ ~new__0793_;
  assign new__0005_ = new__0004_ & new__0769_;
  assign new__0006_ = ~new__0005_ ^ ~\in_array[14] ;
  assign new__0007__neg = ~new__0006_ ^ ~new__0758_;
  assign new__0007_ = ~new__0007__neg;
  assign new__0008_ = ~\in_array[4] ;
  assign new__0009_ = ~\in_array[4]  ^ ~\in_array[0] ;
  assign new__0010_ = new__0009_ & new__0737_;
  assign new__0011_ = ~new__0010_ ^ ~new__0008_;
  assign new__0012_ = ~\in_array[12]  ^ ~\in_array[8] ;
  assign new__0013_ = new__0012_ & new__0004_;
  assign new__0014_ = ~new__0013_ ^ ~\in_array[12] ;
  assign new__0015_ = new__0014_ & new__0011_;
  assign new__0016_ = ~\in_array[5] ;
  assign new__0017_ = ~\in_array[1]  ^ ~\in_array[5] ;
  assign new__0018_ = new__0017_ & new__0737_;
  assign new__0019_ = ~new__0018_ ^ ~new__0016_;
  assign new__0020_ = ~new__0019_ ^ ~new__0015_;
  assign new__0021_ = ~\in_array[9]  ^ ~\in_array[13] ;
  assign new__0022_ = new__0021_ & new__0004_;
  assign new__0023_ = ~new__0022_ ^ ~\in_array[13] ;
  assign new__0024_ = ~new__0023_ ^ ~new__0015_;
  assign new__0025_ = new__0024_ & new__0020_;
  assign new__0026_ = ~new__0025_ ^ ~new__0015_;
  assign new__0027_ = ~new__0026_;
  assign new__0028_ = ~new__0026_ ^ ~new__0758_;
  assign new__0029_ = ~new__0026_ ^ ~new__0006_;
  assign new__0030_ = new__0029_ & new__0028_;
  assign new__0031_ = ~new__0030_ ^ ~new__0027_;
  assign new__0032_ = ~\in_array[7] ;
  assign new__0033_ = \in_array[3]  & new__0032_;
  assign new__0034_ = ~new__0033_ ^ ~new__0032_;
  assign new__0035_ = ~new__0034_;
  assign new__0036_ = ~new__0035_ ^ ~new__0031_;
  assign new__0037_ = new__0000_ & \in_array[15] ;
  assign new__0038_ = ~new__0037_ ^ ~\in_array[15] ;
  assign new__0039_ = ~new__0038_;
  assign new__0040_ = ~new__0039_ ^ ~new__0031_;
  assign new__0041_ = new__0040_ & new__0036_;
  assign new__0042_ = ~new__0041_ ^ ~new__0031_;
  assign new__0043_ = new__0042_ & new__0007_;
  assign new__0044_ = ~new__0043_ ^ ~new__0758_;
  assign new__0045_ = ~new__0747_ ^ ~new__0633_;
  assign new__0046_ = ~new__0045_;
  assign new__0047_ = ~new__0005_ ^ ~\in_array[10] ;
  assign new__0048__neg = ~new__0047_ ^ ~new__0045_;
  assign new__0048_ = ~new__0048__neg;
  assign new__0049_ = ~new__0010_ ^ ~new__0569_;
  assign new__0050_ = ~new__0013_ ^ ~\in_array[8] ;
  assign new__0051_ = new__0050_ & new__0049_;
  assign new__0052_ = ~new__0018_ ^ ~new__0587_;
  assign new__0053_ = ~new__0052_ ^ ~new__0051_;
  assign new__0054_ = ~new__0022_ ^ ~\in_array[9] ;
  assign new__0055_ = ~new__0054_ ^ ~new__0051_;
  assign new__0056_ = new__0055_ & new__0053_;
  assign new__0057_ = ~new__0056_ ^ ~new__0051_;
  assign new__0058_ = ~new__0057_;
  assign new__0059_ = ~new__0057_ ^ ~new__0045_;
  assign new__0060_ = ~new__0057_ ^ ~new__0047_;
  assign new__0061_ = new__0060_ & new__0059_;
  assign new__0062_ = ~new__0061_ ^ ~new__0058_;
  assign new__0063_ = ~new__0033_ ^ ~\in_array[3] ;
  assign new__0064_ = ~new__0063_ ^ ~new__0062_;
  assign new__0065_ = ~new__0037_ ^ ~new__0000_;
  assign new__0066_ = ~new__0065_ ^ ~new__0062_;
  assign new__0067_ = new__0066_ & new__0064_;
  assign new__0068_ = ~new__0067_ ^ ~new__0062_;
  assign new__0069_ = new__0068_ & new__0048_;
  assign new__0070_ = ~new__0069_ ^ ~new__0046_;
  assign new__0071__neg = ~new__0070_ ^ ~new__0044_;
  assign new__0071_ = ~new__0071__neg;
  assign new__0072__neg = ~new__0014_ ^ ~new__0011_;
  assign new__0072_ = ~new__0072__neg;
  assign new__0073_ = new__0072_ & new__0042_;
  assign new__0074_ = ~new__0073_ ^ ~new__0011_;
  assign new__0075_ = ~new__0049_;
  assign new__0076__neg = ~new__0050_ ^ ~new__0049_;
  assign new__0076_ = ~new__0076__neg;
  assign new__0077_ = new__0076_ & new__0068_;
  assign new__0078_ = ~new__0077_ ^ ~new__0075_;
  assign new__0079_ = new__0078_ & new__0074_;
  assign new__0080__neg = ~new__0023_ ^ ~new__0019_;
  assign new__0080_ = ~new__0080__neg;
  assign new__0081_ = new__0080_ & new__0042_;
  assign new__0082_ = ~new__0081_ ^ ~new__0019_;
  assign new__0083_ = ~new__0082_ ^ ~new__0079_;
  assign new__0084_ = ~new__0052_;
  assign new__0085__neg = ~new__0054_ ^ ~new__0052_;
  assign new__0085_ = ~new__0085__neg;
  assign new__0086_ = new__0085_ & new__0068_;
  assign new__0087_ = ~new__0086_ ^ ~new__0084_;
  assign new__0088_ = ~new__0087_ ^ ~new__0079_;
  assign new__0089_ = new__0088_ & new__0083_;
  assign new__0090_ = ~new__0089_ ^ ~new__0079_;
  assign new__0091_ = ~new__0090_;
  assign new__0092_ = ~new__0090_ ^ ~new__0044_;
  assign new__0093_ = ~new__0090_ ^ ~new__0070_;
  assign new__0094_ = new__0093_ & new__0092_;
  assign new__0095_ = ~new__0094_ ^ ~new__0091_;
  assign new__0096_ = ~new__0094_ ^ ~new__0090_;
  assign new__0097__neg = ~new__0038_ ^ ~new__0034_;
  assign new__0097_ = ~new__0097__neg;
  assign new__0098_ = new__0097_ & new__0042_;
  assign new__0099_ = ~new__0098_ ^ ~new__0034_;
  assign new__0100_ = ~new__0099_ ^ ~new__0096_;
  assign new__0101_ = ~new__0063_;
  assign new__0102__neg = ~new__0065_ ^ ~new__0063_;
  assign new__0102_ = ~new__0102__neg;
  assign new__0103_ = new__0102_ & new__0068_;
  assign new__0104_ = ~new__0103_ ^ ~new__0101_;
  assign new__0105_ = ~new__0104_ ^ ~new__0095_;
  assign new__0106_ = new__0105_ & new__0100_;
  assign new__0107_ = ~new__0106_ ^ ~new__0095_;
  assign new__0108_ = new__0107_ & new__0071_;
  assign new__0109_ = ~new__0108_ ^ ~new__0044_;
  assign new__0110_ = ~new__0109_;
  assign new__0111_ = ~\in_array[22] ;
  assign new__0112_ = ~\in_array[18]  ^ ~\in_array[22] ;
  assign new__0113_ = ~\in_array[16] ;
  assign new__0114_ = \in_array[20]  & new__0113_;
  assign new__0115_ = ~\in_array[17] ;
  assign new__0116_ = ~new__0114_ ^ ~new__0115_;
  assign new__0117_ = ~new__0114_ ^ ~\in_array[21] ;
  assign new__0118_ = new__0117_ & new__0116_;
  assign new__0119_ = ~new__0118_ ^ ~new__0114_;
  assign new__0120_ = ~\in_array[18] ;
  assign new__0121_ = ~new__0119_ ^ ~new__0120_;
  assign new__0122_ = ~new__0119_ ^ ~\in_array[22] ;
  assign new__0123_ = new__0122_ & new__0121_;
  assign new__0124_ = ~new__0123_ ^ ~new__0119_;
  assign new__0125_ = ~new__0124_;
  assign new__0126_ = ~\in_array[19] ;
  assign new__0127_ = ~new__0124_ ^ ~new__0126_;
  assign new__0128_ = ~new__0124_ ^ ~\in_array[23] ;
  assign new__0129_ = new__0128_ & new__0127_;
  assign new__0130_ = ~new__0129_ ^ ~new__0125_;
  assign new__0131_ = new__0130_ & new__0112_;
  assign new__0132_ = ~new__0131_ ^ ~new__0111_;
  assign new__0133_ = ~\in_array[26]  ^ ~\in_array[30] ;
  assign new__0134_ = ~\in_array[24] ;
  assign new__0135_ = \in_array[28]  & new__0134_;
  assign new__0136_ = ~\in_array[25] ;
  assign new__0137_ = ~new__0135_ ^ ~new__0136_;
  assign new__0138_ = ~new__0135_ ^ ~\in_array[29] ;
  assign new__0139_ = new__0138_ & new__0137_;
  assign new__0140_ = ~new__0139_ ^ ~new__0135_;
  assign new__0141_ = ~\in_array[26] ;
  assign new__0142_ = ~new__0140_ ^ ~new__0141_;
  assign new__0143_ = ~new__0140_ ^ ~\in_array[30] ;
  assign new__0144_ = new__0143_ & new__0142_;
  assign new__0145_ = ~new__0144_ ^ ~new__0140_;
  assign new__0146_ = ~\in_array[27] ;
  assign new__0147_ = ~new__0145_ ^ ~new__0146_;
  assign new__0148_ = ~new__0145_ ^ ~\in_array[31] ;
  assign new__0149_ = new__0148_ & new__0147_;
  assign new__0150_ = ~new__0149_ ^ ~new__0145_;
  assign new__0151_ = new__0150_ & new__0133_;
  assign new__0152_ = ~new__0151_ ^ ~\in_array[30] ;
  assign new__0153__neg = ~new__0152_ ^ ~new__0132_;
  assign new__0153_ = ~new__0153__neg;
  assign new__0154_ = ~\in_array[20] ;
  assign new__0155_ = ~\in_array[20]  ^ ~\in_array[16] ;
  assign new__0156_ = new__0155_ & new__0130_;
  assign new__0157_ = ~new__0156_ ^ ~new__0154_;
  assign new__0158_ = ~\in_array[28]  ^ ~\in_array[24] ;
  assign new__0159_ = new__0158_ & new__0150_;
  assign new__0160_ = ~new__0159_ ^ ~\in_array[28] ;
  assign new__0161_ = new__0160_ & new__0157_;
  assign new__0162_ = ~\in_array[21] ;
  assign new__0163_ = ~\in_array[17]  ^ ~\in_array[21] ;
  assign new__0164_ = new__0163_ & new__0130_;
  assign new__0165_ = ~new__0164_ ^ ~new__0162_;
  assign new__0166_ = ~new__0165_ ^ ~new__0161_;
  assign new__0167_ = ~\in_array[25]  ^ ~\in_array[29] ;
  assign new__0168_ = new__0167_ & new__0150_;
  assign new__0169_ = ~new__0168_ ^ ~\in_array[29] ;
  assign new__0170_ = ~new__0169_ ^ ~new__0161_;
  assign new__0171_ = new__0170_ & new__0166_;
  assign new__0172_ = ~new__0171_ ^ ~new__0161_;
  assign new__0173_ = ~new__0172_ ^ ~new__0132_;
  assign new__0174_ = ~new__0172_ ^ ~new__0152_;
  assign new__0175_ = new__0174_ & new__0173_;
  assign new__0176_ = ~new__0175_ ^ ~new__0172_;
  assign new__0177_ = ~\in_array[23] ;
  assign new__0178_ = \in_array[19]  & new__0177_;
  assign new__0179_ = ~new__0178_ ^ ~new__0177_;
  assign new__0180_ = ~new__0179_ ^ ~new__0176_;
  assign new__0181_ = new__0146_ & \in_array[31] ;
  assign new__0182_ = ~new__0181_ ^ ~\in_array[31] ;
  assign new__0183_ = ~new__0182_ ^ ~new__0176_;
  assign new__0184_ = new__0183_ & new__0180_;
  assign new__0185_ = ~new__0184_ ^ ~new__0176_;
  assign new__0186_ = new__0185_ & new__0153_;
  assign new__0187_ = ~new__0186_ ^ ~new__0132_;
  assign new__0188_ = ~new__0187_;
  assign new__0189_ = ~new__0131_ ^ ~new__0120_;
  assign new__0190_ = ~new__0189_;
  assign new__0191_ = ~new__0151_ ^ ~\in_array[26] ;
  assign new__0192__neg = ~new__0191_ ^ ~new__0189_;
  assign new__0192_ = ~new__0192__neg;
  assign new__0193_ = ~new__0156_ ^ ~new__0113_;
  assign new__0194_ = ~new__0159_ ^ ~\in_array[24] ;
  assign new__0195_ = new__0194_ & new__0193_;
  assign new__0196_ = ~new__0164_ ^ ~new__0115_;
  assign new__0197_ = ~new__0196_ ^ ~new__0195_;
  assign new__0198_ = ~new__0168_ ^ ~\in_array[25] ;
  assign new__0199_ = ~new__0198_ ^ ~new__0195_;
  assign new__0200_ = new__0199_ & new__0197_;
  assign new__0201_ = ~new__0200_ ^ ~new__0195_;
  assign new__0202_ = ~new__0201_ ^ ~new__0189_;
  assign new__0203_ = ~new__0201_ ^ ~new__0191_;
  assign new__0204_ = new__0203_ & new__0202_;
  assign new__0205_ = ~new__0204_ ^ ~new__0201_;
  assign new__0206_ = ~new__0178_ ^ ~\in_array[19] ;
  assign new__0207_ = ~new__0206_;
  assign new__0208_ = ~new__0207_ ^ ~new__0205_;
  assign new__0209_ = ~new__0181_ ^ ~new__0146_;
  assign new__0210_ = ~new__0209_;
  assign new__0211_ = ~new__0210_ ^ ~new__0205_;
  assign new__0212_ = new__0211_ & new__0208_;
  assign new__0213_ = ~new__0212_ ^ ~new__0205_;
  assign new__0214_ = new__0213_ & new__0192_;
  assign new__0215_ = ~new__0214_ ^ ~new__0190_;
  assign new__0216__neg = ~new__0215_ ^ ~new__0187_;
  assign new__0216_ = ~new__0216__neg;
  assign new__0217__neg = ~new__0160_ ^ ~new__0157_;
  assign new__0217_ = ~new__0217__neg;
  assign new__0218_ = new__0217_ & new__0185_;
  assign new__0219_ = ~new__0218_ ^ ~new__0157_;
  assign new__0220_ = ~new__0193_;
  assign new__0221__neg = ~new__0194_ ^ ~new__0193_;
  assign new__0221_ = ~new__0221__neg;
  assign new__0222_ = new__0221_ & new__0213_;
  assign new__0223_ = ~new__0222_ ^ ~new__0220_;
  assign new__0224_ = new__0223_ & new__0219_;
  assign new__0225__neg = ~new__0169_ ^ ~new__0165_;
  assign new__0225_ = ~new__0225__neg;
  assign new__0226_ = new__0225_ & new__0185_;
  assign new__0227_ = ~new__0226_ ^ ~new__0165_;
  assign new__0228_ = ~new__0227_ ^ ~new__0224_;
  assign new__0229_ = ~new__0196_;
  assign new__0230__neg = ~new__0198_ ^ ~new__0196_;
  assign new__0230_ = ~new__0230__neg;
  assign new__0231_ = new__0230_ & new__0213_;
  assign new__0232_ = ~new__0231_ ^ ~new__0229_;
  assign new__0233_ = ~new__0232_ ^ ~new__0224_;
  assign new__0234_ = new__0233_ & new__0228_;
  assign new__0235_ = ~new__0234_ ^ ~new__0224_;
  assign new__0236_ = ~new__0235_ ^ ~new__0187_;
  assign new__0237_ = ~new__0235_ ^ ~new__0215_;
  assign new__0238_ = new__0237_ & new__0236_;
  assign new__0239_ = ~new__0238_ ^ ~new__0235_;
  assign new__0240__neg = ~new__0182_ ^ ~new__0179_;
  assign new__0240_ = ~new__0240__neg;
  assign new__0241_ = new__0240_ & new__0185_;
  assign new__0242_ = ~new__0241_ ^ ~new__0179_;
  assign new__0243_ = ~new__0242_ ^ ~new__0239_;
  assign new__0244_ = ~new__0235_;
  assign new__0245_ = ~new__0238_ ^ ~new__0244_;
  assign new__0246__neg = ~new__0209_ ^ ~new__0206_;
  assign new__0246_ = ~new__0246__neg;
  assign new__0247_ = new__0246_ & new__0213_;
  assign new__0248_ = ~new__0247_ ^ ~new__0207_;
  assign new__0249_ = ~new__0248_ ^ ~new__0245_;
  assign new__0250_ = new__0249_ & new__0243_;
  assign new__0251_ = ~new__0250_ ^ ~new__0239_;
  assign new__0252_ = new__0251_ & new__0216_;
  assign new__0253_ = ~new__0252_ ^ ~new__0188_;
  assign new__0254__neg = ~new__0253_ ^ ~new__0109_;
  assign new__0254_ = ~new__0254__neg;
  assign new__0255__neg = ~new__0078_ ^ ~new__0074_;
  assign new__0255_ = ~new__0255__neg;
  assign new__0256_ = new__0255_ & new__0107_;
  assign new__0257_ = ~new__0256_ ^ ~new__0074_;
  assign new__0258_ = ~new__0219_;
  assign new__0259__neg = ~new__0223_ ^ ~new__0219_;
  assign new__0259_ = ~new__0259__neg;
  assign new__0260_ = new__0259_ & new__0251_;
  assign new__0261_ = ~new__0260_ ^ ~new__0258_;
  assign new__0262_ = new__0261_ & new__0257_;
  assign new__0263__neg = ~new__0087_ ^ ~new__0082_;
  assign new__0263_ = ~new__0263__neg;
  assign new__0264_ = new__0263_ & new__0107_;
  assign new__0265_ = ~new__0264_ ^ ~new__0082_;
  assign new__0266_ = ~new__0265_ ^ ~new__0262_;
  assign new__0267_ = ~new__0227_;
  assign new__0268__neg = ~new__0232_ ^ ~new__0227_;
  assign new__0268_ = ~new__0268__neg;
  assign new__0269_ = new__0268_ & new__0251_;
  assign new__0270_ = ~new__0269_ ^ ~new__0267_;
  assign new__0271_ = ~new__0270_ ^ ~new__0262_;
  assign new__0272_ = new__0271_ & new__0266_;
  assign new__0273_ = ~new__0272_ ^ ~new__0262_;
  assign new__0274_ = ~new__0273_;
  assign new__0275_ = ~new__0273_ ^ ~new__0109_;
  assign new__0276_ = ~new__0273_ ^ ~new__0253_;
  assign new__0277_ = new__0276_ & new__0275_;
  assign new__0278_ = ~new__0277_ ^ ~new__0274_;
  assign new__0279_ = ~new__0277_ ^ ~new__0273_;
  assign new__0280_ = ~new__0104_ ^ ~new__0099_;
  assign new__0281_ = new__0280_ & new__0107_;
  assign new__0282_ = ~new__0281_ ^ ~new__0099_;
  assign new__0283_ = ~new__0282_ ^ ~new__0279_;
  assign new__0284_ = ~new__0248_ ^ ~new__0242_;
  assign new__0285_ = new__0284_ & new__0251_;
  assign new__0286_ = ~new__0285_ ^ ~new__0242_;
  assign new__0287_ = ~new__0286_ ^ ~new__0278_;
  assign new__0288_ = new__0287_ & new__0283_;
  assign new__0289_ = ~new__0288_ ^ ~new__0278_;
  assign new__0290_ = new__0289_ & new__0254_;
  assign new__0291_ = ~new__0290_ ^ ~new__0110_;
  assign new__0292_ = ~new__0006_;
  assign new__0293_ = ~new__0043_ ^ ~new__0292_;
  assign new__0294_ = ~new__0069_ ^ ~new__0047_;
  assign new__0295__neg = ~new__0294_ ^ ~new__0293_;
  assign new__0295_ = ~new__0295__neg;
  assign new__0296_ = ~new__0014_;
  assign new__0297_ = ~new__0073_ ^ ~new__0296_;
  assign new__0298_ = ~new__0077_ ^ ~new__0050_;
  assign new__0299_ = new__0298_ & new__0297_;
  assign new__0300_ = ~new__0023_;
  assign new__0301_ = ~new__0081_ ^ ~new__0300_;
  assign new__0302_ = ~new__0301_ ^ ~new__0299_;
  assign new__0303_ = ~new__0086_ ^ ~new__0054_;
  assign new__0304_ = ~new__0303_ ^ ~new__0299_;
  assign new__0305_ = new__0304_ & new__0302_;
  assign new__0306_ = ~new__0305_ ^ ~new__0299_;
  assign new__0307_ = ~new__0306_;
  assign new__0308_ = ~new__0306_ ^ ~new__0293_;
  assign new__0309_ = ~new__0306_ ^ ~new__0294_;
  assign new__0310_ = new__0309_ & new__0308_;
  assign new__0311_ = ~new__0310_ ^ ~new__0307_;
  assign new__0312_ = ~new__0310_ ^ ~new__0306_;
  assign new__0313_ = ~new__0098_ ^ ~new__0039_;
  assign new__0314_ = ~new__0313_ ^ ~new__0312_;
  assign new__0315_ = ~new__0103_ ^ ~new__0065_;
  assign new__0316_ = ~new__0315_ ^ ~new__0311_;
  assign new__0317_ = new__0316_ & new__0314_;
  assign new__0318_ = ~new__0317_ ^ ~new__0311_;
  assign new__0319_ = new__0318_ & new__0295_;
  assign new__0320_ = ~new__0319_ ^ ~new__0293_;
  assign new__0321_ = ~new__0152_;
  assign new__0322_ = ~new__0186_ ^ ~new__0321_;
  assign new__0323_ = ~new__0322_;
  assign new__0324_ = ~new__0214_ ^ ~new__0191_;
  assign new__0325__neg = ~new__0324_ ^ ~new__0322_;
  assign new__0325_ = ~new__0325__neg;
  assign new__0326_ = ~new__0160_;
  assign new__0327_ = ~new__0218_ ^ ~new__0326_;
  assign new__0328_ = ~new__0222_ ^ ~new__0194_;
  assign new__0329_ = new__0328_ & new__0327_;
  assign new__0330_ = ~new__0169_;
  assign new__0331_ = ~new__0226_ ^ ~new__0330_;
  assign new__0332_ = ~new__0331_ ^ ~new__0329_;
  assign new__0333_ = ~new__0231_ ^ ~new__0198_;
  assign new__0334_ = ~new__0333_ ^ ~new__0329_;
  assign new__0335_ = new__0334_ & new__0332_;
  assign new__0336_ = ~new__0335_ ^ ~new__0329_;
  assign new__0337_ = ~new__0336_ ^ ~new__0322_;
  assign new__0338_ = ~new__0336_ ^ ~new__0324_;
  assign new__0339_ = new__0338_ & new__0337_;
  assign new__0340_ = ~new__0339_ ^ ~new__0336_;
  assign new__0341_ = ~new__0182_;
  assign new__0342_ = ~new__0241_ ^ ~new__0341_;
  assign new__0343_ = ~new__0342_ ^ ~new__0340_;
  assign new__0344_ = ~new__0336_;
  assign new__0345_ = ~new__0339_ ^ ~new__0344_;
  assign new__0346_ = ~new__0247_ ^ ~new__0209_;
  assign new__0347_ = ~new__0346_ ^ ~new__0345_;
  assign new__0348_ = new__0347_ & new__0343_;
  assign new__0349_ = ~new__0348_ ^ ~new__0340_;
  assign new__0350_ = new__0349_ & new__0325_;
  assign new__0351_ = ~new__0350_ ^ ~new__0323_;
  assign new__0352__neg = ~new__0351_ ^ ~new__0320_;
  assign new__0352_ = ~new__0352__neg;
  assign new__0353__neg = ~new__0298_ ^ ~new__0297_;
  assign new__0353_ = ~new__0353__neg;
  assign new__0354_ = new__0353_ & new__0318_;
  assign new__0355_ = ~new__0354_ ^ ~new__0297_;
  assign new__0356_ = ~new__0327_;
  assign new__0357__neg = ~new__0328_ ^ ~new__0327_;
  assign new__0357_ = ~new__0357__neg;
  assign new__0358_ = new__0357_ & new__0349_;
  assign new__0359_ = ~new__0358_ ^ ~new__0356_;
  assign new__0360_ = new__0359_ & new__0355_;
  assign new__0361__neg = ~new__0303_ ^ ~new__0301_;
  assign new__0361_ = ~new__0361__neg;
  assign new__0362_ = new__0361_ & new__0318_;
  assign new__0363_ = ~new__0362_ ^ ~new__0301_;
  assign new__0364_ = ~new__0363_ ^ ~new__0360_;
  assign new__0365_ = ~new__0331_;
  assign new__0366__neg = ~new__0333_ ^ ~new__0331_;
  assign new__0366_ = ~new__0366__neg;
  assign new__0367_ = new__0366_ & new__0349_;
  assign new__0368_ = ~new__0367_ ^ ~new__0365_;
  assign new__0369_ = ~new__0368_ ^ ~new__0360_;
  assign new__0370_ = new__0369_ & new__0364_;
  assign new__0371_ = ~new__0370_ ^ ~new__0360_;
  assign new__0372_ = ~new__0371_;
  assign new__0373_ = ~new__0371_ ^ ~new__0320_;
  assign new__0374_ = ~new__0371_ ^ ~new__0351_;
  assign new__0375_ = new__0374_ & new__0373_;
  assign new__0376_ = ~new__0375_ ^ ~new__0372_;
  assign new__0377_ = ~new__0375_ ^ ~new__0371_;
  assign new__0378_ = ~new__0315_ ^ ~new__0313_;
  assign new__0379_ = new__0378_ & new__0318_;
  assign new__0380_ = ~new__0379_ ^ ~new__0313_;
  assign new__0381_ = ~new__0380_ ^ ~new__0377_;
  assign new__0382_ = ~new__0346_ ^ ~new__0342_;
  assign new__0383_ = new__0382_ & new__0349_;
  assign new__0384_ = ~new__0383_ ^ ~new__0342_;
  assign new__0385_ = ~new__0384_ ^ ~new__0376_;
  assign new__0386_ = new__0385_ & new__0381_;
  assign new__0387_ = ~new__0386_ ^ ~new__0376_;
  assign new__0388_ = new__0387_ & new__0352_;
  assign new__0389_ = ~new__0388_ ^ ~new__0320_;
  assign new__0390__neg = ~new__0389_ ^ ~new__0291_;
  assign new__0390_ = ~new__0390__neg;
  assign new__0391__neg = ~new__0359_ ^ ~new__0355_;
  assign new__0391_ = ~new__0391__neg;
  assign new__0392_ = new__0391_ & new__0387_;
  assign new__0393_ = ~new__0392_ ^ ~new__0355_;
  assign new__0394_ = ~new__0257_;
  assign new__0395__neg = ~new__0261_ ^ ~new__0257_;
  assign new__0395_ = ~new__0395__neg;
  assign new__0396_ = new__0395_ & new__0289_;
  assign new__0397_ = ~new__0396_ ^ ~new__0394_;
  assign new__0398_ = new__0397_ & new__0393_;
  assign new__0399__neg = ~new__0368_ ^ ~new__0363_;
  assign new__0399_ = ~new__0399__neg;
  assign new__0400_ = new__0399_ & new__0387_;
  assign new__0401_ = ~new__0400_ ^ ~new__0363_;
  assign new__0402_ = ~new__0401_ ^ ~new__0398_;
  assign new__0403_ = ~new__0265_;
  assign new__0404__neg = ~new__0270_ ^ ~new__0265_;
  assign new__0404_ = ~new__0404__neg;
  assign new__0405_ = new__0404_ & new__0289_;
  assign new__0406_ = ~new__0405_ ^ ~new__0403_;
  assign new__0407_ = ~new__0406_ ^ ~new__0398_;
  assign new__0408_ = new__0407_ & new__0402_;
  assign new__0409_ = ~new__0408_ ^ ~new__0398_;
  assign new__0410_ = ~new__0409_;
  assign new__0411_ = ~new__0409_ ^ ~new__0389_;
  assign new__0412_ = ~new__0409_ ^ ~new__0291_;
  assign new__0413_ = new__0412_ & new__0411_;
  assign new__0414_ = ~new__0413_ ^ ~new__0410_;
  assign new__0415_ = ~new__0413_ ^ ~new__0409_;
  assign new__0416_ = ~new__0384_ ^ ~new__0380_;
  assign new__0417_ = new__0416_ & new__0387_;
  assign new__0418_ = ~new__0417_ ^ ~new__0380_;
  assign new__0419_ = ~new__0418_ ^ ~new__0415_;
  assign new__0420_ = ~new__0286_ ^ ~new__0282_;
  assign new__0421_ = new__0420_ & new__0289_;
  assign new__0422_ = ~new__0421_ ^ ~new__0282_;
  assign new__0423_ = ~new__0422_ ^ ~new__0414_;
  assign new__0424_ = new__0423_ & new__0419_;
  assign new__0425_ = ~new__0424_ ^ ~new__0414_;
  assign new__0426_ = new__0425_ & new__0390_;
  assign new__0427_ = ~new__0426_ ^ ~new__0291_;
  assign new__0428_ = ~new__0070_;
  assign new__0429_ = ~new__0108_ ^ ~new__0428_;
  assign new__0430_ = ~new__0429_;
  assign new__0431_ = ~new__0252_ ^ ~new__0215_;
  assign new__0432__neg = ~new__0431_ ^ ~new__0429_;
  assign new__0432_ = ~new__0432__neg;
  assign new__0433_ = ~new__0078_;
  assign new__0434_ = ~new__0256_ ^ ~new__0433_;
  assign new__0435_ = ~new__0260_ ^ ~new__0223_;
  assign new__0436_ = new__0435_ & new__0434_;
  assign new__0437_ = ~new__0087_;
  assign new__0438_ = ~new__0264_ ^ ~new__0437_;
  assign new__0439_ = ~new__0438_ ^ ~new__0436_;
  assign new__0440_ = ~new__0269_ ^ ~new__0232_;
  assign new__0441_ = ~new__0440_ ^ ~new__0436_;
  assign new__0442_ = new__0441_ & new__0439_;
  assign new__0443_ = ~new__0442_ ^ ~new__0436_;
  assign new__0444_ = ~new__0443_;
  assign new__0445_ = ~new__0443_ ^ ~new__0429_;
  assign new__0446_ = ~new__0443_ ^ ~new__0431_;
  assign new__0447_ = new__0446_ & new__0445_;
  assign new__0448_ = ~new__0447_ ^ ~new__0444_;
  assign new__0449_ = ~new__0447_ ^ ~new__0443_;
  assign new__0450_ = ~new__0281_ ^ ~new__0104_;
  assign new__0451_ = ~new__0450_ ^ ~new__0449_;
  assign new__0452_ = ~new__0285_ ^ ~new__0248_;
  assign new__0453_ = ~new__0452_ ^ ~new__0448_;
  assign new__0454_ = new__0453_ & new__0451_;
  assign new__0455_ = ~new__0454_ ^ ~new__0448_;
  assign new__0456_ = new__0455_ & new__0432_;
  assign new__0457_ = ~new__0456_ ^ ~new__0430_;
  assign new__0458_ = ~new__0457_;
  assign new__0459_ = ~new__0294_;
  assign new__0460_ = ~new__0319_ ^ ~new__0459_;
  assign new__0461_ = ~new__0350_ ^ ~new__0324_;
  assign new__0462__neg = ~new__0461_ ^ ~new__0460_;
  assign new__0462_ = ~new__0462__neg;
  assign new__0463_ = ~new__0298_;
  assign new__0464_ = ~new__0354_ ^ ~new__0463_;
  assign new__0465_ = ~new__0358_ ^ ~new__0328_;
  assign new__0466_ = new__0465_ & new__0464_;
  assign new__0467_ = ~new__0303_;
  assign new__0468_ = ~new__0362_ ^ ~new__0467_;
  assign new__0469_ = ~new__0468_ ^ ~new__0466_;
  assign new__0470_ = ~new__0367_ ^ ~new__0333_;
  assign new__0471_ = ~new__0470_ ^ ~new__0466_;
  assign new__0472_ = new__0471_ & new__0469_;
  assign new__0473_ = ~new__0472_ ^ ~new__0466_;
  assign new__0474_ = ~new__0473_;
  assign new__0475_ = ~new__0473_ ^ ~new__0460_;
  assign new__0476_ = ~new__0473_ ^ ~new__0461_;
  assign new__0477_ = new__0476_ & new__0475_;
  assign new__0478_ = ~new__0477_ ^ ~new__0474_;
  assign new__0479_ = ~new__0477_ ^ ~new__0473_;
  assign new__0480_ = ~new__0379_ ^ ~new__0315_;
  assign new__0481_ = ~new__0480_ ^ ~new__0479_;
  assign new__0482_ = ~new__0383_ ^ ~new__0346_;
  assign new__0483_ = ~new__0482_ ^ ~new__0478_;
  assign new__0484_ = new__0483_ & new__0481_;
  assign new__0485_ = ~new__0484_ ^ ~new__0478_;
  assign new__0486_ = new__0485_ & new__0462_;
  assign new__0487_ = ~new__0486_ ^ ~new__0460_;
  assign new__0488__neg = ~new__0487_ ^ ~new__0457_;
  assign new__0488_ = ~new__0488__neg;
  assign new__0489__neg = ~new__0465_ ^ ~new__0464_;
  assign new__0489_ = ~new__0489__neg;
  assign new__0490_ = new__0489_ & new__0485_;
  assign new__0491_ = ~new__0490_ ^ ~new__0464_;
  assign new__0492_ = ~new__0434_;
  assign new__0493__neg = ~new__0435_ ^ ~new__0434_;
  assign new__0493_ = ~new__0493__neg;
  assign new__0494_ = new__0493_ & new__0455_;
  assign new__0495_ = ~new__0494_ ^ ~new__0492_;
  assign new__0496_ = new__0495_ & new__0491_;
  assign new__0497__neg = ~new__0470_ ^ ~new__0468_;
  assign new__0497_ = ~new__0497__neg;
  assign new__0498_ = new__0497_ & new__0485_;
  assign new__0499_ = ~new__0498_ ^ ~new__0468_;
  assign new__0500_ = ~new__0499_ ^ ~new__0496_;
  assign new__0501_ = ~new__0438_;
  assign new__0502__neg = ~new__0440_ ^ ~new__0438_;
  assign new__0502_ = ~new__0502__neg;
  assign new__0503_ = new__0502_ & new__0455_;
  assign new__0504_ = ~new__0503_ ^ ~new__0501_;
  assign new__0505_ = ~new__0504_ ^ ~new__0496_;
  assign new__0506_ = new__0505_ & new__0500_;
  assign new__0507_ = ~new__0506_ ^ ~new__0496_;
  assign new__0508_ = ~new__0507_;
  assign new__0509_ = ~new__0507_ ^ ~new__0487_;
  assign new__0510_ = ~new__0507_ ^ ~new__0457_;
  assign new__0511_ = new__0510_ & new__0509_;
  assign new__0512_ = ~new__0511_ ^ ~new__0508_;
  assign new__0513_ = ~new__0511_ ^ ~new__0507_;
  assign new__0514_ = ~new__0482_ ^ ~new__0480_;
  assign new__0515_ = new__0514_ & new__0485_;
  assign new__0516_ = ~new__0515_ ^ ~new__0480_;
  assign new__0517_ = ~new__0516_ ^ ~new__0513_;
  assign new__0518_ = ~new__0452_ ^ ~new__0450_;
  assign new__0519_ = new__0518_ & new__0455_;
  assign new__0520_ = ~new__0519_ ^ ~new__0450_;
  assign new__0521_ = ~new__0520_ ^ ~new__0512_;
  assign new__0522_ = new__0521_ & new__0517_;
  assign new__0523_ = ~new__0522_ ^ ~new__0512_;
  assign new__0524_ = new__0523_ & new__0488_;
  assign new__0525_ = ~new__0524_ ^ ~new__0458_;
  assign new__0526__neg = ~new__0525_ ^ ~new__0427_;
  assign new__0526_ = ~new__0526__neg;
  assign new__0527_ = ~new__0495_;
  assign new__0528__neg = ~new__0495_ ^ ~new__0491_;
  assign new__0528_ = ~new__0528__neg;
  assign new__0529_ = new__0528_ & new__0523_;
  assign new__0530_ = ~new__0529_ ^ ~new__0527_;
  assign new__0531__neg = ~new__0397_ ^ ~new__0393_;
  assign new__0531_ = ~new__0531__neg;
  assign new__0532_ = new__0531_ & new__0425_;
  assign new__0533_ = ~new__0532_ ^ ~new__0397_;
  assign new__0534_ = new__0533_ & new__0530_;
  assign new__0535_ = ~new__0504_;
  assign new__0536__neg = ~new__0504_ ^ ~new__0499_;
  assign new__0536_ = ~new__0536__neg;
  assign new__0537_ = new__0536_ & new__0523_;
  assign new__0538_ = ~new__0537_ ^ ~new__0535_;
  assign new__0539_ = ~new__0538_ ^ ~new__0534_;
  assign new__0540__neg = ~new__0406_ ^ ~new__0401_;
  assign new__0540_ = ~new__0540__neg;
  assign new__0541_ = new__0540_ & new__0425_;
  assign new__0542_ = ~new__0541_ ^ ~new__0406_;
  assign new__0543_ = ~new__0542_ ^ ~new__0534_;
  assign new__0544_ = new__0543_ & new__0539_;
  assign new__0545_ = ~new__0544_ ^ ~new__0534_;
  assign new__0546_ = ~new__0545_;
  assign new__0547_ = ~new__0545_ ^ ~new__0525_;
  assign new__0548_ = ~new__0545_ ^ ~new__0427_;
  assign new__0549_ = new__0548_ & new__0547_;
  assign new__0551_ = ~new__0549_ ^ ~new__0546_;
  assign new__0552_ = ~new__0549_ ^ ~new__0545_;
  assign new__0553_ = ~new__0520_ ^ ~new__0516_;
  assign new__0554_ = new__0553_ & new__0523_;
  assign new__0555_ = ~new__0554_ ^ ~new__0520_;
  assign new__0556_ = ~new__0555_ ^ ~new__0552_;
  assign new__0557_ = ~new__0422_ ^ ~new__0418_;
  assign new__0558_ = new__0557_ & new__0425_;
  assign new__0559_ = ~new__0558_ ^ ~new__0422_;
  assign new__0560_ = ~new__0559_ ^ ~new__0551_;
  assign new__0562_ = new__0560_ & new__0556_;
  assign new__0563_ = ~new__0562_ ^ ~new__0551_;
  assign new__0564_ = new__0563_ & new__0526_;
  assign \out_array[18]  = ~new__0564_ ^ ~new__0427_;
  assign new__0565__neg = ~new__0542_ ^ ~new__0538_;
  assign new__0565_ = ~new__0565__neg;
  assign new__0566_ = new__0565_ & new__0563_;
  assign \out_array[17]  = ~new__0566_ ^ ~new__0542_;
  assign new__0567__neg = ~new__0533_ ^ ~new__0530_;
  assign new__0567_ = ~new__0567__neg;
  assign new__0568_ = new__0567_ & new__0563_;
  assign \out_array[16]  = ~new__0568_ ^ ~new__0533_;
  assign new__0570_ = ~new__0525_;
  assign \out_array[22]  = ~new__0564_ ^ ~new__0570_;
  assign new__0571_ = ~new__0538_;
  assign \out_array[21]  = ~new__0566_ ^ ~new__0571_;
  assign new__0572_ = ~new__0530_;
  assign \out_array[20]  = ~new__0568_ ^ ~new__0572_;
  assign new__0573_ = ~new__0559_;
  assign new__0574_ = ~new__0559_ ^ ~new__0555_;
  assign new__0575_ = new__0574_ & new__0563_;
  assign \out_array[19]  = ~new__0575_ ^ ~new__0573_;
  assign new__0577_ = ~new__0389_;
  assign new__0578_ = ~new__0426_ ^ ~new__0577_;
  assign new__0579_ = ~new__0524_ ^ ~new__0487_;
  assign new__0580__neg = ~new__0579_ ^ ~new__0578_;
  assign new__0580_ = ~new__0580__neg;
  assign new__0581_ = ~new__0529_ ^ ~new__0491_;
  assign new__0582_ = ~new__0393_;
  assign new__0583_ = ~new__0532_ ^ ~new__0582_;
  assign new__0584_ = new__0583_ & new__0581_;
  assign new__0585_ = ~new__0537_ ^ ~new__0499_;
  assign new__0586_ = ~new__0585_ ^ ~new__0584_;
  assign new__0588_ = ~new__0401_;
  assign new__0589_ = ~new__0541_ ^ ~new__0588_;
  assign new__0590_ = ~new__0589_ ^ ~new__0584_;
  assign new__0591_ = new__0590_ & new__0586_;
  assign new__0592_ = ~new__0591_ ^ ~new__0584_;
  assign new__0593_ = ~new__0592_;
  assign new__0594_ = ~new__0592_ ^ ~new__0579_;
  assign new__0595_ = ~new__0592_ ^ ~new__0578_;
  assign new__0596_ = new__0595_ & new__0594_;
  assign new__0597_ = ~new__0596_ ^ ~new__0593_;
  assign new__0599_ = ~new__0596_ ^ ~new__0592_;
  assign new__0600_ = ~new__0554_ ^ ~new__0516_;
  assign new__0601_ = ~new__0600_ ^ ~new__0599_;
  assign new__0602_ = ~new__0558_ ^ ~new__0418_;
  assign new__0603_ = ~new__0602_ ^ ~new__0597_;
  assign new__0604_ = new__0603_ & new__0601_;
  assign new__0605_ = ~new__0604_ ^ ~new__0597_;
  assign new__0606_ = new__0605_ & new__0580_;
  assign \out_array[26]  = ~new__0606_ ^ ~new__0578_;
  assign new__0607__neg = ~new__0589_ ^ ~new__0585_;
  assign new__0607_ = ~new__0607__neg;
  assign new__0609_ = new__0607_ & new__0605_;
  assign \out_array[25]  = ~new__0609_ ^ ~new__0589_;
  assign new__0610__neg = ~new__0583_ ^ ~new__0581_;
  assign new__0610_ = ~new__0610__neg;
  assign new__0611_ = new__0610_ & new__0605_;
  assign \out_array[24]  = ~new__0611_ ^ ~new__0583_;
  assign new__0612_ = ~new__0579_;
  assign \out_array[30]  = ~new__0606_ ^ ~new__0612_;
  assign new__0613_ = ~new__0585_;
  assign \out_array[29]  = ~new__0609_ ^ ~new__0613_;
  assign new__0614_ = ~new__0581_;
  assign \out_array[28]  = ~new__0611_ ^ ~new__0614_;
  assign new__0616_ = ~new__0602_;
  assign new__0617_ = ~new__0602_ ^ ~new__0600_;
  assign new__0618_ = new__0617_ & new__0605_;
  assign \out_array[27]  = ~new__0618_ ^ ~new__0616_;
  assign new__0619_ = ~new__0555_;
  assign \out_array[23]  = ~new__0575_ ^ ~new__0619_;
  assign new__0620_ = ~new__0600_;
  assign \out_array[31]  = ~new__0618_ ^ ~new__0620_;
  assign new__0621_ = ~new__0290_ ^ ~new__0253_;
  assign new__0623_ = ~new__0351_;
  assign new__0624_ = ~new__0388_ ^ ~new__0623_;
  assign new__0625__neg = ~new__0624_ ^ ~new__0621_;
  assign new__0625_ = ~new__0625__neg;
  assign new__0626_ = ~new__0359_;
  assign new__0627_ = ~new__0392_ ^ ~new__0626_;
  assign new__0628_ = ~new__0396_ ^ ~new__0261_;
  assign new__0629_ = new__0628_ & new__0627_;
  assign new__0630_ = ~new__0368_;
  assign new__0631_ = ~new__0400_ ^ ~new__0630_;
  assign new__0632_ = ~new__0631_ ^ ~new__0629_;
  assign new__0634_ = ~new__0405_ ^ ~new__0270_;
  assign new__0635_ = ~new__0634_ ^ ~new__0629_;
  assign new__0636_ = new__0635_ & new__0632_;
  assign new__0637_ = ~new__0636_ ^ ~new__0629_;
  assign new__0638_ = ~new__0637_;
  assign new__0639_ = ~new__0637_ ^ ~new__0624_;
  assign new__0640_ = ~new__0637_ ^ ~new__0621_;
  assign new__0641_ = new__0640_ & new__0639_;
  assign new__0642_ = ~new__0641_ ^ ~new__0638_;
  assign new__0643_ = ~new__0641_ ^ ~new__0637_;
  assign new__0645_ = ~new__0417_ ^ ~new__0384_;
  assign new__0646_ = ~new__0645_ ^ ~new__0643_;
  assign new__0647_ = ~new__0421_ ^ ~new__0286_;
  assign new__0648_ = ~new__0647_ ^ ~new__0642_;
  assign new__0649_ = new__0648_ & new__0646_;
  assign new__0650_ = ~new__0649_ ^ ~new__0642_;
  assign new__0651_ = new__0650_ & new__0625_;
  assign new__0652_ = ~new__0651_ ^ ~new__0621_;
  assign new__0653_ = ~new__0456_ ^ ~new__0431_;
  assign new__0654_ = ~new__0653_;
  assign new__0656_ = ~new__0461_;
  assign new__0657_ = ~new__0486_ ^ ~new__0656_;
  assign new__0658__neg = ~new__0657_ ^ ~new__0653_;
  assign new__0658_ = ~new__0658__neg;
  assign new__0659_ = ~new__0465_;
  assign new__0660_ = ~new__0490_ ^ ~new__0659_;
  assign new__0661_ = ~new__0494_ ^ ~new__0435_;
  assign new__0662_ = new__0661_ & new__0660_;
  assign new__0663_ = ~new__0470_;
  assign new__0664_ = ~new__0498_ ^ ~new__0663_;
  assign new__0665_ = ~new__0664_ ^ ~new__0662_;
  assign new__0667_ = ~new__0503_ ^ ~new__0440_;
  assign new__0668_ = ~new__0667_ ^ ~new__0662_;
  assign new__0669_ = new__0668_ & new__0665_;
  assign new__0670_ = ~new__0669_ ^ ~new__0662_;
  assign new__0671_ = ~new__0670_;
  assign new__0672_ = ~new__0670_ ^ ~new__0657_;
  assign new__0673_ = ~new__0670_ ^ ~new__0653_;
  assign new__0674_ = new__0673_ & new__0672_;
  assign new__0675_ = ~new__0674_ ^ ~new__0671_;
  assign new__0676_ = ~new__0674_ ^ ~new__0670_;
  assign new__0678_ = ~new__0515_ ^ ~new__0482_;
  assign new__0679_ = ~new__0678_ ^ ~new__0676_;
  assign new__0680_ = ~new__0519_ ^ ~new__0452_;
  assign new__0681_ = ~new__0680_ ^ ~new__0675_;
  assign new__0682_ = new__0681_ & new__0679_;
  assign new__0683_ = ~new__0682_ ^ ~new__0675_;
  assign new__0684_ = new__0683_ & new__0658_;
  assign new__0685_ = ~new__0684_ ^ ~new__0654_;
  assign new__0686__neg = ~new__0685_ ^ ~new__0652_;
  assign new__0686_ = ~new__0686__neg;
  assign new__0687_ = ~new__0661_;
  assign new__0689__neg = ~new__0661_ ^ ~new__0660_;
  assign new__0689_ = ~new__0689__neg;
  assign new__0690_ = new__0689_ & new__0683_;
  assign new__0691_ = ~new__0690_ ^ ~new__0687_;
  assign new__0692__neg = ~new__0628_ ^ ~new__0627_;
  assign new__0692_ = ~new__0692__neg;
  assign new__0693_ = new__0692_ & new__0650_;
  assign new__0694_ = ~new__0693_ ^ ~new__0628_;
  assign new__0695_ = new__0694_ & new__0691_;
  assign new__0696_ = ~new__0667_;
  assign new__0697__neg = ~new__0667_ ^ ~new__0664_;
  assign new__0697_ = ~new__0697__neg;
  assign new__0698_ = new__0697_ & new__0683_;
  assign new__0700_ = ~new__0698_ ^ ~new__0696_;
  assign new__0701_ = ~new__0700_ ^ ~new__0695_;
  assign new__0702__neg = ~new__0634_ ^ ~new__0631_;
  assign new__0702_ = ~new__0702__neg;
  assign new__0703_ = new__0702_ & new__0650_;
  assign new__0704_ = ~new__0703_ ^ ~new__0634_;
  assign new__0705_ = ~new__0704_ ^ ~new__0695_;
  assign new__0706_ = new__0705_ & new__0701_;
  assign new__0707_ = ~new__0706_ ^ ~new__0695_;
  assign new__0708_ = ~new__0707_;
  assign new__0709_ = ~new__0707_ ^ ~new__0685_;
  assign new__0711_ = ~new__0707_ ^ ~new__0652_;
  assign new__0712_ = new__0711_ & new__0709_;
  assign new__0713_ = ~new__0712_ ^ ~new__0708_;
  assign new__0714_ = ~new__0712_ ^ ~new__0707_;
  assign new__0715_ = ~new__0680_ ^ ~new__0678_;
  assign new__0716_ = new__0715_ & new__0683_;
  assign new__0717_ = ~new__0716_ ^ ~new__0680_;
  assign new__0718_ = ~new__0717_ ^ ~new__0714_;
  assign new__0719_ = ~new__0647_ ^ ~new__0645_;
  assign new__0720_ = new__0719_ & new__0650_;
  assign new__0722_ = ~new__0720_ ^ ~new__0647_;
  assign new__0723_ = ~new__0722_ ^ ~new__0713_;
  assign new__0724_ = new__0723_ & new__0718_;
  assign new__0725_ = ~new__0724_ ^ ~new__0713_;
  assign new__0726_ = new__0725_ & new__0686_;
  assign \out_array[2]  = ~new__0726_ ^ ~new__0652_;
  assign new__0727__neg = ~new__0704_ ^ ~new__0700_;
  assign new__0727_ = ~new__0727__neg;
  assign new__0728_ = new__0727_ & new__0725_;
  assign \out_array[1]  = ~new__0728_ ^ ~new__0704_;
  assign new__0729__neg = ~new__0694_ ^ ~new__0691_;
  assign new__0729_ = ~new__0729__neg;
  assign new__0731_ = new__0729_ & new__0725_;
  assign \out_array[0]  = ~new__0731_ ^ ~new__0694_;
  assign new__0732_ = ~new__0685_;
  assign \out_array[6]  = ~new__0726_ ^ ~new__0732_;
  assign new__0733_ = ~new__0700_;
  assign \out_array[5]  = ~new__0728_ ^ ~new__0733_;
  assign new__0734_ = ~new__0691_;
  assign \out_array[4]  = ~new__0731_ ^ ~new__0734_;
  assign new__0735_ = ~new__0722_;
  assign new__0736_ = ~new__0722_ ^ ~new__0717_;
  assign new__0738_ = new__0736_ & new__0725_;
  assign \out_array[3]  = ~new__0738_ ^ ~new__0735_;
  assign new__0739_ = ~new__0624_;
  assign new__0740_ = ~new__0651_ ^ ~new__0739_;
  assign new__0741_ = ~new__0684_ ^ ~new__0657_;
  assign new__0742__neg = ~new__0741_ ^ ~new__0740_;
  assign new__0742_ = ~new__0742__neg;
  assign new__0743_ = ~new__0690_ ^ ~new__0660_;
  assign new__0744_ = ~new__0627_;
  assign new__0745_ = ~new__0693_ ^ ~new__0744_;
  assign new__0746_ = new__0745_ & new__0743_;
  assign new__0748_ = ~new__0698_ ^ ~new__0664_;
  assign new__0749_ = ~new__0748_ ^ ~new__0746_;
  assign new__0750_ = ~new__0631_;
  assign new__0751_ = ~new__0703_ ^ ~new__0750_;
  assign new__0752_ = ~new__0751_ ^ ~new__0746_;
  assign new__0753_ = new__0752_ & new__0749_;
  assign new__0754_ = ~new__0753_ ^ ~new__0746_;
  assign new__0755_ = ~new__0754_;
  assign new__0756_ = ~new__0754_ ^ ~new__0741_;
  assign new__0757_ = ~new__0754_ ^ ~new__0740_;
  assign new__0759_ = new__0757_ & new__0756_;
  assign new__0760_ = ~new__0759_ ^ ~new__0755_;
  assign new__0761_ = ~new__0759_ ^ ~new__0754_;
  assign new__0762_ = ~new__0716_ ^ ~new__0678_;
  assign new__0763_ = ~new__0762_ ^ ~new__0761_;
  assign new__0764_ = ~new__0720_ ^ ~new__0645_;
  assign new__0765_ = ~new__0764_ ^ ~new__0760_;
  assign new__0766_ = new__0765_ & new__0763_;
  assign new__0767_ = ~new__0766_ ^ ~new__0760_;
  assign new__0768_ = new__0767_ & new__0742_;
  assign \out_array[10]  = ~new__0768_ ^ ~new__0740_;
  assign new__0770__neg = ~new__0751_ ^ ~new__0748_;
  assign new__0770_ = ~new__0770__neg;
  assign new__0771_ = new__0770_ & new__0767_;
  assign \out_array[9]  = ~new__0771_ ^ ~new__0751_;
  assign new__0772__neg = ~new__0745_ ^ ~new__0743_;
  assign new__0772_ = ~new__0772__neg;
  assign new__0773_ = new__0772_ & new__0767_;
  assign \out_array[8]  = ~new__0773_ ^ ~new__0745_;
  assign new__0774_ = ~new__0741_;
  assign \out_array[14]  = ~new__0768_ ^ ~new__0774_;
  assign new__0775_ = ~new__0748_;
  assign \out_array[13]  = ~new__0771_ ^ ~new__0775_;
  assign new__0777_ = ~new__0743_;
  assign \out_array[12]  = ~new__0773_ ^ ~new__0777_;
  assign new__0778_ = ~new__0764_;
  assign new__0779_ = ~new__0764_ ^ ~new__0762_;
  assign new__0780_ = new__0779_ & new__0767_;
  assign \out_array[11]  = ~new__0780_ ^ ~new__0778_;
  assign new__0781_ = ~new__0717_;
  assign \out_array[7]  = ~new__0738_ ^ ~new__0781_;
  assign new__0782_ = ~new__0762_;
  assign \out_array[15]  = ~new__0780_ ^ ~new__0782_;
endmodule


