module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 ;
  assign n70 = x2 & ~x8 ;
  assign n71 = x9 & n70 ;
  assign n33 = x2 & x6 ;
  assign n58 = n33 ^ x6 ;
  assign n59 = x3 & n58 ;
  assign n60 = n59 ^ x3 ;
  assign n61 = x1 & x8 ;
  assign n62 = n61 ^ x1 ;
  assign n63 = n62 ^ x8 ;
  assign n64 = x9 & n63 ;
  assign n65 = n64 ^ x9 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = n60 & n66 ;
  assign n68 = n67 ^ n60 ;
  assign n69 = n68 ^ n66 ;
  assign n72 = n71 ^ n69 ;
  assign n79 = x2 & x3 ;
  assign n80 = n79 ^ x2 ;
  assign n81 = x1 & x9 ;
  assign n82 = n81 ^ x9 ;
  assign n83 = n80 & n82 ;
  assign n73 = x0 & x5 ;
  assign n74 = n73 ^ x0 ;
  assign n84 = n74 ^ x5 ;
  assign n85 = n62 & n84 ;
  assign n86 = n85 ^ n62 ;
  assign n87 = n86 ^ n84 ;
  assign n88 = n83 & n87 ;
  assign n89 = n88 ^ n83 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = n72 & n90 ;
  assign n92 = n91 ^ n72 ;
  assign n93 = n92 ^ n90 ;
  assign n94 = n93 ^ n90 ;
  assign n75 = n72 & n74 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = n77 ^ x5 ;
  assign n95 = n94 ^ n78 ;
  assign n101 = n81 ^ x1 ;
  assign n102 = n101 ^ x9 ;
  assign n103 = x8 & n102 ;
  assign n104 = n103 ^ x8 ;
  assign n105 = n104 ^ n102 ;
  assign n106 = n80 ^ x3 ;
  assign n107 = x0 & n106 ;
  assign n108 = n107 ^ x0 ;
  assign n109 = n108 ^ n106 ;
  assign n110 = n105 & ~n109 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = n95 & ~n111 ;
  assign n113 = n112 ^ n95 ;
  assign n11 = x1 & x3 ;
  assign n12 = n11 ^ x1 ;
  assign n23 = x0 & x9 ;
  assign n29 = n23 ^ x9 ;
  assign n30 = n12 & n29 ;
  assign n31 = n30 ^ n12 ;
  assign n24 = n23 ^ x0 ;
  assign n25 = x2 & n24 ;
  assign n26 = n25 ^ x2 ;
  assign n27 = n26 ^ n24 ;
  assign n15 = x9 ^ x2 ;
  assign n16 = n15 ^ x9 ;
  assign n13 = x9 ^ x0 ;
  assign n14 = n13 ^ x9 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n14 ^ x9 ;
  assign n19 = n17 & ~n18 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = n12 & ~n20 ;
  assign n22 = n21 ^ n12 ;
  assign n28 = n27 ^ n22 ;
  assign n32 = n31 ^ n28 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n34 ^ x6 ;
  assign n36 = n24 & ~n35 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = n37 ^ x6 ;
  assign n39 = x5 & ~n38 ;
  assign n40 = n39 ^ x5 ;
  assign n41 = n40 ^ x5 ;
  assign n42 = n32 & n41 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = ~x1 & ~x2 ;
  assign n46 = ~x9 & n45 ;
  assign n47 = n46 ^ x2 ;
  assign n48 = n47 ^ x9 ;
  assign n49 = x0 & x3 ;
  assign n50 = n49 ^ x0 ;
  assign n51 = n50 ^ x3 ;
  assign n52 = x6 & ~n51 ;
  assign n53 = n48 & n52 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = n44 & n54 ;
  assign n56 = n55 ^ n44 ;
  assign n57 = n56 ^ n54 ;
  assign n96 = x8 & ~n95 ;
  assign n97 = n96 ^ x8 ;
  assign n98 = n57 & n97 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = n99 ^ n97 ;
  assign n114 = n113 ^ n100 ;
  assign n119 = x0 & x2 ;
  assign n120 = n119 ^ x0 ;
  assign n121 = n120 ^ x2 ;
  assign n122 = n82 & n121 ;
  assign n123 = n122 ^ n82 ;
  assign n124 = x5 & x6 ;
  assign n125 = n124 ^ x6 ;
  assign n126 = n123 & n125 ;
  assign n127 = n126 ^ n125 ;
  assign n128 = n127 ^ x6 ;
  assign n129 = n128 ^ x8 ;
  assign n130 = x1 & x5 ;
  assign n131 = x2 & ~n13 ;
  assign n132 = n130 & n131 ;
  assign n133 = n132 ^ x8 ;
  assign n134 = n132 & ~n133 ;
  assign n135 = n134 ^ x8 ;
  assign n136 = ~n129 & ~n135 ;
  assign n137 = n136 ^ n134 ;
  assign n138 = n137 ^ n128 ;
  assign n139 = n138 ^ x8 ;
  assign n140 = n29 & ~n63 ;
  assign n141 = n140 ^ n63 ;
  assign n142 = n141 ^ x8 ;
  assign n143 = x1 & x2 ;
  assign n144 = n143 ^ x2 ;
  assign n145 = n24 & n144 ;
  assign n146 = ~n142 & n145 ;
  assign n147 = n146 ^ n145 ;
  assign n148 = n147 ^ n142 ;
  assign n149 = n148 ^ n145 ;
  assign n150 = x5 & ~n149 ;
  assign n151 = n150 ^ x5 ;
  assign n152 = n151 ^ n149 ;
  assign n153 = x3 & ~x7 ;
  assign n154 = ~n152 & n153 ;
  assign n155 = n154 ^ n153 ;
  assign n156 = n155 ^ n153 ;
  assign n157 = ~n139 & n156 ;
  assign n158 = n157 ^ n156 ;
  assign n159 = ~n114 & n158 ;
  assign n160 = n159 ^ n158 ;
  assign n115 = ~x3 & ~x7 ;
  assign n116 = ~n114 & n115 ;
  assign n117 = n116 ^ n115 ;
  assign n118 = n117 ^ x7 ;
  assign n161 = n160 ^ n118 ;
  assign n190 = x1 & n29 ;
  assign n191 = n190 ^ x1 ;
  assign n192 = x3 & x5 ;
  assign n193 = n192 ^ x3 ;
  assign n194 = n193 ^ x5 ;
  assign n195 = n82 & n194 ;
  assign n196 = n195 ^ n82 ;
  assign n197 = n196 ^ n194 ;
  assign n198 = n191 & n197 ;
  assign n199 = n198 ^ n191 ;
  assign n200 = n199 ^ n197 ;
  assign n206 = x7 & n101 ;
  assign n207 = n206 ^ x7 ;
  assign n208 = n207 ^ n101 ;
  assign n201 = x1 & x7 ;
  assign n202 = n201 ^ x1 ;
  assign n203 = n202 ^ x7 ;
  assign n204 = n24 & ~n203 ;
  assign n205 = n204 ^ n203 ;
  assign n209 = n208 ^ n205 ;
  assign n213 = n200 & ~n209 ;
  assign n214 = n213 ^ n200 ;
  assign n215 = n214 ^ n209 ;
  assign n216 = n215 ^ n200 ;
  assign n217 = n216 ^ n209 ;
  assign n210 = x2 & ~n209 ;
  assign n211 = n200 & n210 ;
  assign n212 = n211 ^ x2 ;
  assign n218 = n217 ^ n212 ;
  assign n219 = ~x7 & ~x9 ;
  assign n224 = x0 & x1 ;
  assign n225 = n224 ^ x0 ;
  assign n226 = n225 ^ x1 ;
  assign n220 = x3 & x9 ;
  assign n227 = n220 ^ x3 ;
  assign n228 = n226 & n227 ;
  assign n229 = n228 ^ n227 ;
  assign n230 = n229 ^ x3 ;
  assign n221 = n220 ^ x9 ;
  assign n222 = n144 & n221 ;
  assign n223 = n222 ^ x1 ;
  assign n231 = n230 ^ n223 ;
  assign n232 = n219 & n231 ;
  assign n233 = n232 ^ n219 ;
  assign n239 = x2 ^ x0 ;
  assign n234 = x5 ^ x1 ;
  assign n235 = n234 ^ x5 ;
  assign n236 = n235 ^ x5 ;
  assign n270 = x5 ^ x2 ;
  assign n271 = n270 ^ n235 ;
  assign n272 = n236 & n271 ;
  assign n273 = n272 ^ n271 ;
  assign n274 = n273 ^ n236 ;
  assign n275 = n274 ^ n235 ;
  assign n276 = n239 & ~n275 ;
  assign n277 = n276 ^ n239 ;
  assign n278 = n277 ^ n275 ;
  assign n279 = n278 ^ x2 ;
  assign n280 = n279 ^ x5 ;
  assign n281 = n280 ^ x5 ;
  assign n282 = n233 & n281 ;
  assign n283 = n282 ^ n233 ;
  assign n284 = n283 ^ n233 ;
  assign n268 = x7 & n231 ;
  assign n269 = n268 ^ n231 ;
  assign n285 = n284 ^ n269 ;
  assign n264 = ~x7 & x8 ;
  assign n265 = n231 & n264 ;
  assign n240 = n239 ^ x2 ;
  assign n255 = n240 ^ x8 ;
  assign n242 = n240 ^ x2 ;
  assign n247 = n242 ^ x8 ;
  assign n248 = n242 & n247 ;
  assign n257 = n248 ^ n235 ;
  assign n256 = n236 ^ x8 ;
  assign n258 = n257 ^ n256 ;
  assign n259 = ~n255 & ~n258 ;
  assign n251 = n242 ^ n240 ;
  assign n241 = n240 ^ n236 ;
  assign n243 = n242 ^ n241 ;
  assign n244 = n242 ^ n236 ;
  assign n245 = n244 ^ x8 ;
  assign n246 = n243 & ~n245 ;
  assign n249 = n248 ^ n246 ;
  assign n250 = n249 ^ n235 ;
  assign n252 = n251 ^ n250 ;
  assign n253 = n246 ^ n235 ;
  assign n254 = ~n252 & n253 ;
  assign n260 = n259 ^ n254 ;
  assign n261 = n260 ^ n248 ;
  assign n237 = n236 ^ n235 ;
  assign n238 = n237 ^ x8 ;
  assign n262 = n261 ^ n238 ;
  assign n263 = n233 & ~n262 ;
  assign n266 = n265 ^ n263 ;
  assign n267 = n266 ^ x8 ;
  assign n286 = n285 ^ n267 ;
  assign n287 = ~n218 & n286 ;
  assign n288 = n287 ^ n218 ;
  assign n289 = n288 ^ n286 ;
  assign n290 = n289 ^ x8 ;
  assign n305 = x9 ^ x7 ;
  assign n303 = x9 ^ x5 ;
  assign n304 = n303 ^ x9 ;
  assign n306 = n305 ^ n304 ;
  assign n308 = n306 ^ x9 ;
  assign n310 = n308 ^ n306 ;
  assign n307 = n306 ^ n304 ;
  assign n311 = n307 ^ n306 ;
  assign n312 = ~n310 & n311 ;
  assign n313 = n312 ^ n306 ;
  assign n316 = n312 ^ n307 ;
  assign n314 = n303 ^ x1 ;
  assign n315 = n314 ^ n308 ;
  assign n317 = n316 ^ n315 ;
  assign n318 = ~n313 & n317 ;
  assign n319 = n318 ^ n312 ;
  assign n309 = n308 ^ n307 ;
  assign n320 = n319 ^ n309 ;
  assign n323 = n316 ^ n308 ;
  assign n324 = n314 ^ n307 ;
  assign n321 = n306 ^ x8 ;
  assign n325 = n324 ^ n321 ;
  assign n326 = ~n323 & n325 ;
  assign n327 = n326 ^ n318 ;
  assign n328 = n327 ^ n312 ;
  assign n322 = n321 ^ n307 ;
  assign n329 = n328 ^ n322 ;
  assign n330 = ~n320 & ~n329 ;
  assign n331 = n330 ^ n318 ;
  assign n332 = n331 ^ n306 ;
  assign n333 = n332 ^ n303 ;
  assign n334 = n333 ^ x9 ;
  assign n335 = n334 ^ n314 ;
  assign n336 = n335 ^ n308 ;
  assign n337 = n336 ^ n307 ;
  assign n338 = n337 ^ n306 ;
  assign n291 = x5 & x7 ;
  assign n292 = n291 ^ x7 ;
  assign n293 = x8 & n292 ;
  assign n294 = x2 & x9 ;
  assign n295 = n294 ^ x2 ;
  assign n296 = n226 & n295 ;
  assign n297 = n296 ^ n295 ;
  assign n298 = n293 & n297 ;
  assign n339 = ~x3 & n120 ;
  assign n340 = n298 & n339 ;
  assign n341 = n340 ^ n339 ;
  assign n342 = n338 & n341 ;
  assign n343 = n342 ^ n341 ;
  assign n344 = n343 ^ n341 ;
  assign n345 = ~n290 & n344 ;
  assign n346 = n345 ^ n344 ;
  assign n299 = ~x3 & n298 ;
  assign n300 = ~n290 & n299 ;
  assign n301 = n300 ^ n299 ;
  assign n302 = n301 ^ n290 ;
  assign n347 = n346 ^ n302 ;
  assign n162 = x6 ^ x5 ;
  assign n163 = n162 ^ x8 ;
  assign n164 = n163 ^ x8 ;
  assign n165 = n164 ^ n163 ;
  assign n166 = x5 ^ x4 ;
  assign n167 = n166 ^ x6 ;
  assign n168 = n167 ^ n163 ;
  assign n169 = n168 ^ n164 ;
  assign n170 = ~x9 & n169 ;
  assign n171 = n170 ^ n164 ;
  assign n172 = ~n165 & ~n171 ;
  assign n173 = n172 ^ n169 ;
  assign n174 = x6 & ~n164 ;
  assign n175 = n174 ^ n165 ;
  assign n176 = n173 & ~n175 ;
  assign n177 = n176 ^ n174 ;
  assign n178 = n177 ^ x8 ;
  assign n179 = n178 ^ n162 ;
  assign n180 = n179 ^ n164 ;
  assign n181 = n12 ^ x3 ;
  assign n182 = ~x7 & ~n121 ;
  assign n183 = ~n181 & n182 ;
  assign n184 = n180 & n183 ;
  assign n185 = n184 ^ n183 ;
  assign n348 = ~x4 & ~x6 ;
  assign n349 = n185 & n348 ;
  assign n350 = n349 ^ n348 ;
  assign n351 = ~n347 & n350 ;
  assign n352 = n351 ^ n350 ;
  assign n353 = n352 ^ n350 ;
  assign n354 = n161 & n353 ;
  assign n186 = ~x4 & ~n185 ;
  assign n187 = n161 & n186 ;
  assign n188 = n187 ^ n186 ;
  assign n189 = n188 ^ n185 ;
  assign n355 = n354 ^ n189 ;
  assign n356 = x2 & x8 ;
  assign n369 = n356 ^ x8 ;
  assign n370 = n369 ^ x0 ;
  assign n371 = x5 ^ x0 ;
  assign n372 = n371 ^ x0 ;
  assign n373 = n371 & n372 ;
  assign n374 = n373 ^ n371 ;
  assign n375 = n374 ^ n369 ;
  assign n376 = n370 & n375 ;
  assign n377 = n376 ^ n373 ;
  assign n378 = n377 ^ n369 ;
  assign n381 = n378 ^ x1 ;
  assign n357 = n356 ^ x2 ;
  assign n358 = n357 ^ x8 ;
  assign n359 = x5 & n358 ;
  assign n360 = n359 ^ x5 ;
  assign n361 = x5 ^ x3 ;
  assign n362 = x8 & n361 ;
  assign n363 = n362 ^ n361 ;
  assign n364 = n363 ^ x5 ;
  assign n365 = x0 & n364 ;
  assign n366 = n360 & n365 ;
  assign n367 = n366 ^ n360 ;
  assign n368 = n367 ^ n365 ;
  assign n379 = n378 ^ n368 ;
  assign n380 = n379 ^ n378 ;
  assign n382 = n381 ^ n380 ;
  assign n383 = n380 ^ n378 ;
  assign n384 = ~n382 & ~n383 ;
  assign n385 = n384 ^ n382 ;
  assign n386 = n385 ^ n380 ;
  assign n387 = ~x0 & ~x2 ;
  assign n388 = x3 & x8 ;
  assign n389 = n387 & ~n388 ;
  assign n390 = n389 ^ x0 ;
  assign n391 = x6 & ~n390 ;
  assign n392 = n391 ^ x6 ;
  assign n393 = n392 ^ n390 ;
  assign n394 = n386 & n393 ;
  assign n395 = n394 ^ x6 ;
  assign n396 = ~x5 & ~x9 ;
  assign n397 = x8 ^ x2 ;
  assign n398 = n397 ^ x8 ;
  assign n399 = n398 ^ x1 ;
  assign n402 = n399 ^ n398 ;
  assign n400 = n399 ^ x8 ;
  assign n403 = n402 ^ n400 ;
  assign n404 = n402 ^ x6 ;
  assign n405 = n403 ^ x3 ;
  assign n406 = n404 & n405 ;
  assign n407 = n406 ^ x6 ;
  assign n408 = n407 ^ n403 ;
  assign n409 = n403 & n408 ;
  assign n410 = n409 ^ n403 ;
  assign n411 = n410 ^ n406 ;
  assign n412 = n411 ^ x6 ;
  assign n401 = n400 ^ n399 ;
  assign n413 = n412 ^ n401 ;
  assign n414 = n402 ^ n399 ;
  assign n416 = n400 ^ x6 ;
  assign n415 = n402 ^ x3 ;
  assign n417 = n416 ^ n415 ;
  assign n418 = ~n414 & ~n417 ;
  assign n419 = n418 ^ n410 ;
  assign n420 = n419 ^ n406 ;
  assign n421 = n413 & n420 ;
  assign n422 = x0 & x8 ;
  assign n423 = n422 ^ x8 ;
  assign n424 = x2 & n423 ;
  assign n425 = n424 ^ x2 ;
  assign n426 = n425 ^ n423 ;
  assign n427 = x6 ^ x0 ;
  assign n428 = x1 & n427 ;
  assign n429 = n428 ^ x1 ;
  assign n430 = n429 ^ x6 ;
  assign n431 = ~n426 & n430 ;
  assign n432 = n421 & n431 ;
  assign n433 = n432 ^ n421 ;
  assign n434 = n433 ^ n431 ;
  assign n435 = n396 & n434 ;
  assign n436 = n435 ^ x9 ;
  assign n437 = n395 & n436 ;
  assign n438 = n437 ^ n395 ;
  assign n439 = n438 ^ n436 ;
  assign n440 = n439 ^ n436 ;
  assign n452 = n11 ^ x3 ;
  assign n453 = n358 & n452 ;
  assign n454 = n453 ^ n452 ;
  assign n455 = x0 & n130 ;
  assign n456 = n455 ^ x0 ;
  assign n457 = n454 & n456 ;
  assign n458 = n457 ^ n456 ;
  assign n459 = n458 ^ x0 ;
  assign n460 = n459 ^ x6 ;
  assign n464 = n143 & n193 ;
  assign n465 = n464 ^ x5 ;
  assign n461 = ~x2 & ~x3 ;
  assign n462 = ~x5 & n461 ;
  assign n463 = n462 ^ n106 ;
  assign n466 = n465 ^ n463 ;
  assign n467 = n466 ^ x6 ;
  assign n468 = ~n466 & n467 ;
  assign n469 = n468 ^ x6 ;
  assign n470 = ~n460 & ~n469 ;
  assign n471 = n470 ^ n468 ;
  assign n472 = n471 ^ n459 ;
  assign n473 = n472 ^ x6 ;
  assign n443 = x3 & n143 ;
  assign n441 = x5 & x8 ;
  assign n442 = n441 ^ x5 ;
  assign n444 = n443 ^ n442 ;
  assign n445 = n442 ^ x9 ;
  assign n446 = ~x9 & ~n445 ;
  assign n447 = n446 ^ x9 ;
  assign n448 = n447 ^ n443 ;
  assign n449 = n444 & ~n448 ;
  assign n450 = n449 ^ n446 ;
  assign n451 = n450 ^ n443 ;
  assign n474 = n473 ^ n451 ;
  assign n475 = n451 ^ x4 ;
  assign n476 = x4 & ~n475 ;
  assign n477 = n476 ^ x4 ;
  assign n478 = n477 ^ n473 ;
  assign n479 = n474 & ~n478 ;
  assign n480 = n479 ^ n474 ;
  assign n481 = n480 ^ n478 ;
  assign n482 = n481 ^ n476 ;
  assign n483 = n482 ^ n473 ;
  assign n484 = ~n440 & ~n483 ;
  assign n485 = n484 ^ n483 ;
  assign n486 = n485 ^ n483 ;
  assign n493 = x0 & x6 ;
  assign n538 = n493 ^ x6 ;
  assign n539 = x2 & n538 ;
  assign n540 = n539 ^ x2 ;
  assign n541 = n540 ^ n538 ;
  assign n542 = n441 ^ x8 ;
  assign n550 = n541 & n542 ;
  assign n526 = x6 & x8 ;
  assign n545 = n526 ^ x6 ;
  assign n546 = n545 ^ x8 ;
  assign n551 = n550 ^ n546 ;
  assign n547 = x9 & n546 ;
  assign n543 = x9 & n542 ;
  assign n544 = n541 & n543 ;
  assign n548 = n547 ^ n544 ;
  assign n549 = n548 ^ x9 ;
  assign n552 = n551 ^ n549 ;
  assign n561 = x8 ^ x0 ;
  assign n557 = x9 ^ x8 ;
  assign n553 = x9 ^ x6 ;
  assign n559 = n557 ^ n553 ;
  assign n554 = n553 ^ n303 ;
  assign n555 = n554 ^ x8 ;
  assign n556 = n555 ^ x9 ;
  assign n558 = n557 ^ n556 ;
  assign n560 = n559 ^ n558 ;
  assign n562 = n561 ^ n560 ;
  assign n563 = n562 ^ n560 ;
  assign n564 = n562 ^ n559 ;
  assign n565 = n563 & n564 ;
  assign n566 = n565 ^ n562 ;
  assign n574 = n564 ^ n563 ;
  assign n575 = n574 ^ n562 ;
  assign n567 = n562 ^ n557 ;
  assign n568 = n567 ^ n564 ;
  assign n569 = n568 ^ n563 ;
  assign n570 = n562 ^ x9 ;
  assign n571 = n570 ^ n564 ;
  assign n572 = n571 ^ n563 ;
  assign n573 = n569 & n572 ;
  assign n576 = n575 ^ n573 ;
  assign n577 = n566 & n576 ;
  assign n578 = n577 ^ n562 ;
  assign n579 = n578 ^ n562 ;
  assign n583 = x2 & n579 ;
  assign n584 = n583 ^ x2 ;
  assign n585 = n584 ^ x2 ;
  assign n586 = n585 ^ n579 ;
  assign n532 = x1 & ~x4 ;
  assign n580 = ~x2 & ~n532 ;
  assign n581 = n579 & n580 ;
  assign n582 = n581 ^ n532 ;
  assign n587 = n586 ^ n582 ;
  assign n588 = n552 & ~n587 ;
  assign n589 = n588 ^ n552 ;
  assign n487 = x6 & n84 ;
  assign n488 = n487 ^ x6 ;
  assign n489 = n488 ^ n84 ;
  assign n490 = x8 & x9 ;
  assign n521 = n144 & n490 ;
  assign n522 = ~n489 & n521 ;
  assign n496 = ~x6 & x9 ;
  assign n494 = n490 ^ x9 ;
  assign n495 = n493 & n494 ;
  assign n497 = n496 ^ n495 ;
  assign n519 = n144 & n497 ;
  assign n501 = x5 & ~x9 ;
  assign n499 = n490 ^ x8 ;
  assign n500 = n74 & n499 ;
  assign n502 = n501 ^ n500 ;
  assign n518 = n144 & n502 ;
  assign n520 = n519 ^ n518 ;
  assign n523 = n522 ^ n520 ;
  assign n524 = n523 ^ n144 ;
  assign n505 = n24 ^ x9 ;
  assign n506 = n358 & n505 ;
  assign n507 = n506 ^ n358 ;
  assign n508 = n507 ^ n505 ;
  assign n504 = n294 & n422 ;
  assign n509 = n508 ^ n504 ;
  assign n515 = ~x1 & x5 ;
  assign n516 = ~n509 & n515 ;
  assign n491 = n489 & n490 ;
  assign n492 = n491 ^ n490 ;
  assign n498 = n497 ^ n492 ;
  assign n503 = n502 ^ n498 ;
  assign n510 = x5 & n144 ;
  assign n511 = n509 & n510 ;
  assign n512 = n511 ^ n510 ;
  assign n513 = n503 & n512 ;
  assign n514 = n513 ^ n512 ;
  assign n517 = n516 ^ n514 ;
  assign n525 = n524 ^ n517 ;
  assign n527 = n526 ^ x8 ;
  assign n528 = n295 & n527 ;
  assign n534 = n525 & n528 ;
  assign n535 = n534 ^ n528 ;
  assign n536 = n535 ^ n525 ;
  assign n590 = n589 ^ n536 ;
  assign n591 = n590 ^ n586 ;
  assign n592 = n589 ^ n532 ;
  assign n593 = n591 & n592 ;
  assign n594 = n593 ^ n591 ;
  assign n595 = n594 ^ n592 ;
  assign n596 = n595 ^ n589 ;
  assign n597 = n596 ^ n582 ;
  assign n529 = ~x4 & ~n528 ;
  assign n530 = ~n525 & n529 ;
  assign n531 = n530 ^ x4 ;
  assign n533 = n532 ^ n531 ;
  assign n537 = n536 ^ n533 ;
  assign n598 = n597 ^ n537 ;
  assign n599 = x6 & x9 ;
  assign n600 = n599 ^ x6 ;
  assign n601 = n600 ^ x9 ;
  assign n602 = x8 & n166 ;
  assign n603 = n602 ^ x5 ;
  assign n604 = ~n601 & ~n603 ;
  assign n605 = n604 ^ n601 ;
  assign n606 = x4 & n599 ;
  assign n607 = ~n605 & n606 ;
  assign n608 = n607 ^ n605 ;
  assign n609 = n608 ^ n606 ;
  assign n610 = ~x2 & ~n226 ;
  assign n611 = ~x3 & n610 ;
  assign n612 = ~n609 & n611 ;
  assign n613 = n612 ^ x3 ;
  assign n653 = n598 & n613 ;
  assign n654 = n653 ^ n598 ;
  assign n655 = n654 ^ n613 ;
  assign n656 = n655 ^ n613 ;
  assign n657 = n656 ^ x3 ;
  assign n651 = x3 & x7 ;
  assign n649 = x7 & ~n613 ;
  assign n650 = n598 & n649 ;
  assign n652 = n651 ^ n650 ;
  assign n658 = n657 ^ n652 ;
  assign n659 = n486 & ~n658 ;
  assign n660 = n659 ^ n486 ;
  assign n661 = n660 ^ n658 ;
  assign n662 = n661 ^ x7 ;
  assign n629 = x2 ^ x1 ;
  assign n630 = n629 ^ x8 ;
  assign n631 = n630 ^ n239 ;
  assign n625 = n239 ^ x8 ;
  assign n632 = n631 ^ n625 ;
  assign n624 = n295 ^ x9 ;
  assign n626 = n625 ^ n624 ;
  assign n627 = n624 ^ n239 ;
  assign n628 = n626 & n627 ;
  assign n633 = n632 ^ n628 ;
  assign n634 = ~n239 & ~n632 ;
  assign n635 = n634 ^ n626 ;
  assign n636 = ~n633 & n635 ;
  assign n637 = n636 ^ n624 ;
  assign n638 = n637 ^ x8 ;
  assign n639 = n638 ^ x8 ;
  assign n640 = n639 ^ n239 ;
  assign n641 = n640 ^ n625 ;
  assign n642 = n641 ^ n632 ;
  assign n643 = x7 & ~n297 ;
  assign n644 = ~n642 & n643 ;
  assign n645 = n644 ^ n297 ;
  assign n614 = ~x6 & ~n194 ;
  assign n615 = ~x4 & n614 ;
  assign n646 = x7 & n615 ;
  assign n647 = n645 & n646 ;
  assign n616 = ~x7 & n297 ;
  assign n617 = n615 & n616 ;
  assign n620 = x3 & n617 ;
  assign n618 = ~n613 & n617 ;
  assign n619 = n598 & n618 ;
  assign n621 = n620 ^ n619 ;
  assign n622 = n486 & n621 ;
  assign n623 = n622 ^ n621 ;
  assign n648 = n647 ^ n623 ;
  assign n663 = n662 ^ n648 ;
  assign n664 = n143 & ~n527 ;
  assign n665 = n664 ^ x1 ;
  assign n666 = ~x2 & x5 ;
  assign n667 = ~n388 & n666 ;
  assign n668 = n667 ^ x5 ;
  assign n669 = n665 & n668 ;
  assign n670 = n669 ^ n668 ;
  assign n671 = x9 ^ x3 ;
  assign n672 = ~x6 & ~n671 ;
  assign n675 = n557 ^ x9 ;
  assign n673 = x8 ^ x1 ;
  assign n674 = n673 ^ n557 ;
  assign n676 = n675 ^ n674 ;
  assign n677 = n675 ^ n557 ;
  assign n678 = ~n676 & ~n677 ;
  assign n679 = n678 ^ n675 ;
  assign n680 = n672 & ~n679 ;
  assign n681 = x1 & n221 ;
  assign n682 = x4 & n545 ;
  assign n683 = n682 ^ n545 ;
  assign n684 = n681 & n683 ;
  assign n685 = n684 ^ x4 ;
  assign n686 = n680 & n685 ;
  assign n687 = n686 ^ n680 ;
  assign n688 = n687 ^ n685 ;
  assign n689 = n670 & ~n688 ;
  assign n690 = n689 ^ n688 ;
  assign n695 = ~x5 & ~x8 ;
  assign n693 = ~x2 & x3 ;
  assign n694 = x8 & n693 ;
  assign n696 = n695 ^ n694 ;
  assign n697 = n696 ^ n192 ;
  assign n698 = n101 & ~n697 ;
  assign n691 = ~x3 & n125 ;
  assign n692 = ~n66 & n691 ;
  assign n699 = n698 ^ n692 ;
  assign n711 = ~x8 & n82 ;
  assign n704 = n61 & ~n601 ;
  assign n705 = n704 ^ n601 ;
  assign n702 = x9 & n61 ;
  assign n703 = n702 ^ n61 ;
  assign n706 = n705 ^ n703 ;
  assign n707 = x2 & ~n706 ;
  assign n708 = n707 ^ x2 ;
  assign n709 = n708 ^ n706 ;
  assign n700 = ~x8 & x9 ;
  assign n701 = n45 & n700 ;
  assign n710 = n709 ^ n701 ;
  assign n712 = n711 ^ n710 ;
  assign n713 = x3 & n712 ;
  assign n714 = n699 & n713 ;
  assign n715 = n714 ^ n699 ;
  assign n716 = n715 ^ n713 ;
  assign n717 = ~n690 & ~n716 ;
  assign n718 = x8 & n553 ;
  assign n719 = n718 ^ n553 ;
  assign n720 = n719 ^ x9 ;
  assign n721 = x5 & ~n720 ;
  assign n722 = n721 ^ x5 ;
  assign n723 = n722 ^ n720 ;
  assign n724 = ~x3 & x4 ;
  assign n725 = n45 & n724 ;
  assign n726 = ~n723 & n725 ;
  assign n727 = n726 ^ x4 ;
  assign n728 = x0 & n727 ;
  assign n729 = n728 ^ x0 ;
  assign n730 = n729 ^ n727 ;
  assign n731 = n717 & ~n730 ;
  assign n732 = n731 ^ n730 ;
  assign n808 = n499 ^ x9 ;
  assign n809 = x5 & n808 ;
  assign n810 = n809 ^ x5 ;
  assign n811 = n810 ^ x5 ;
  assign n806 = x5 & x9 ;
  assign n807 = n422 & n806 ;
  assign n812 = n811 ^ n807 ;
  assign n813 = n130 ^ x1 ;
  assign n814 = n294 & n813 ;
  assign n815 = n814 ^ n813 ;
  assign n816 = n815 ^ x1 ;
  assign n817 = n812 & n816 ;
  assign n818 = n817 ^ n816 ;
  assign n819 = x2 & n557 ;
  assign n820 = n819 ^ x2 ;
  assign n821 = n102 & n820 ;
  assign n822 = n821 ^ x2 ;
  assign n823 = x3 & n822 ;
  assign n824 = n823 ^ x3 ;
  assign n825 = n824 ^ n822 ;
  assign n826 = n818 & ~n825 ;
  assign n827 = n826 ^ n825 ;
  assign n828 = n827 ^ x3 ;
  assign n829 = x5 & n452 ;
  assign n830 = n829 ^ x5 ;
  assign n842 = ~x8 & ~x9 ;
  assign n843 = x0 & ~x2 ;
  assign n844 = n842 & n843 ;
  assign n845 = ~n830 & n844 ;
  assign n831 = x2 & n808 ;
  assign n832 = n831 ^ x2 ;
  assign n833 = n832 ^ n808 ;
  assign n834 = n830 & ~n833 ;
  assign n835 = n834 ^ n833 ;
  assign n836 = x9 & n106 ;
  assign n837 = n61 ^ x8 ;
  assign n838 = x0 & n837 ;
  assign n839 = n836 & n838 ;
  assign n840 = ~n835 & n839 ;
  assign n841 = n840 ^ n839 ;
  assign n846 = n845 ^ n841 ;
  assign n847 = ~n828 & n846 ;
  assign n848 = n847 ^ n846 ;
  assign n849 = n848 ^ n828 ;
  assign n850 = n849 ^ n846 ;
  assign n733 = x9 ^ x1 ;
  assign n734 = n733 ^ x9 ;
  assign n736 = n734 ^ n675 ;
  assign n735 = n734 ^ n553 ;
  assign n737 = n736 ^ n735 ;
  assign n741 = n736 & n737 ;
  assign n742 = n741 ^ n736 ;
  assign n739 = n734 ^ x9 ;
  assign n740 = n739 ^ x2 ;
  assign n743 = n742 ^ n740 ;
  assign n756 = x2 & ~n553 ;
  assign n757 = n743 & n756 ;
  assign n754 = n553 & ~n734 ;
  assign n753 = x2 & ~n734 ;
  assign n755 = n754 ^ n753 ;
  assign n758 = n757 ^ n755 ;
  assign n744 = x2 & n743 ;
  assign n745 = n744 ^ x2 ;
  assign n747 = n745 ^ n735 ;
  assign n748 = n747 ^ x2 ;
  assign n749 = n741 ^ n734 ;
  assign n750 = n749 ^ n737 ;
  assign n751 = n748 & n750 ;
  assign n752 = n751 ^ n748 ;
  assign n759 = n758 ^ n752 ;
  assign n746 = n745 ^ n741 ;
  assign n760 = n759 ^ n746 ;
  assign n738 = n737 ^ x2 ;
  assign n761 = n760 ^ n738 ;
  assign n762 = n761 ^ x2 ;
  assign n763 = n762 ^ n557 ;
  assign n764 = n763 ^ x9 ;
  assign n798 = ~x3 & n74 ;
  assign n799 = n764 & n798 ;
  assign n766 = x6 ^ x3 ;
  assign n767 = n766 ^ x9 ;
  assign n768 = n767 ^ x9 ;
  assign n769 = n768 ^ n553 ;
  assign n778 = ~x8 & n769 ;
  assign n765 = n733 ^ x8 ;
  assign n770 = n553 ^ x9 ;
  assign n771 = n770 ^ n769 ;
  assign n772 = x8 & n771 ;
  assign n773 = n772 ^ n771 ;
  assign n774 = n773 ^ n553 ;
  assign n775 = n765 & n774 ;
  assign n776 = n775 ^ n774 ;
  assign n777 = n776 ^ n773 ;
  assign n779 = n778 ^ n777 ;
  assign n780 = n779 ^ n733 ;
  assign n781 = n780 ^ x8 ;
  assign n782 = n781 ^ x9 ;
  assign n783 = n782 ^ n553 ;
  assign n793 = n74 & n106 ;
  assign n794 = n793 ^ n74 ;
  assign n795 = n783 & n794 ;
  assign n796 = n795 ^ n794 ;
  assign n797 = n764 & n796 ;
  assign n800 = n799 ^ n797 ;
  assign n790 = n74 & n764 ;
  assign n791 = n790 ^ n74 ;
  assign n784 = x2 & n74 ;
  assign n785 = n784 ^ n74 ;
  assign n786 = n783 & n785 ;
  assign n787 = n786 ^ n785 ;
  assign n788 = n764 & n787 ;
  assign n789 = n788 ^ n787 ;
  assign n792 = n791 ^ n789 ;
  assign n801 = n800 ^ n792 ;
  assign n802 = n801 ^ n74 ;
  assign n851 = ~x7 & n348 ;
  assign n852 = n802 & n851 ;
  assign n853 = n852 ^ n851 ;
  assign n854 = ~n850 & n853 ;
  assign n855 = n854 ^ n853 ;
  assign n803 = ~x4 & ~x7 ;
  assign n804 = n802 & n803 ;
  assign n805 = n804 ^ x7 ;
  assign n856 = n855 ^ n805 ;
  assign n894 = ~n732 & n856 ;
  assign n895 = n894 ^ n732 ;
  assign n896 = n895 ^ n856 ;
  assign n897 = n896 ^ x7 ;
  assign n857 = n557 ^ x1 ;
  assign n859 = n857 ^ n675 ;
  assign n860 = n675 ^ x7 ;
  assign n861 = x1 ^ x0 ;
  assign n862 = n861 ^ x1 ;
  assign n863 = n862 ^ x1 ;
  assign n864 = n863 ^ x9 ;
  assign n865 = n864 ^ n859 ;
  assign n866 = ~n860 & n865 ;
  assign n867 = n866 ^ x7 ;
  assign n868 = n867 ^ n859 ;
  assign n869 = n859 & ~n868 ;
  assign n870 = n869 ^ n866 ;
  assign n871 = n870 ^ x7 ;
  assign n858 = n857 ^ n557 ;
  assign n872 = n871 ^ n858 ;
  assign n874 = n857 ^ x7 ;
  assign n873 = n864 ^ n675 ;
  assign n875 = n874 ^ n873 ;
  assign n876 = ~n677 & ~n875 ;
  assign n877 = n876 ^ n869 ;
  assign n878 = n877 ^ n866 ;
  assign n879 = n872 & n878 ;
  assign n880 = n879 ^ n862 ;
  assign n881 = n880 ^ x1 ;
  assign n882 = n881 ^ n863 ;
  assign n883 = ~x5 & ~x6 ;
  assign n884 = ~x4 & ~n106 ;
  assign n885 = n883 & n884 ;
  assign n886 = ~n882 & n885 ;
  assign n887 = n886 ^ n885 ;
  assign n892 = ~x7 & n887 ;
  assign n888 = n856 & n887 ;
  assign n889 = n888 ^ n887 ;
  assign n890 = ~n732 & n889 ;
  assign n891 = n890 ^ n889 ;
  assign n893 = n892 ^ n891 ;
  assign n898 = n897 ^ n893 ;
  assign n899 = n898 ^ n887 ;
  assign n900 = n192 ^ x5 ;
  assign n901 = n494 & n900 ;
  assign n902 = n901 ^ x3 ;
  assign n903 = x2 & n902 ;
  assign n904 = n903 ^ x2 ;
  assign n905 = n904 ^ x2 ;
  assign n906 = n905 ^ n902 ;
  assign n910 = n388 ^ x3 ;
  assign n911 = x6 & n910 ;
  assign n912 = n911 ^ x6 ;
  assign n913 = n912 ^ n910 ;
  assign n907 = ~x6 & x8 ;
  assign n908 = n193 & n907 ;
  assign n909 = n908 ^ n193 ;
  assign n914 = n913 ^ n909 ;
  assign n915 = n906 & n914 ;
  assign n916 = n915 ^ n906 ;
  assign n917 = n916 ^ n914 ;
  assign n918 = n270 ^ x5 ;
  assign n919 = n361 ^ n270 ;
  assign n920 = n918 & n919 ;
  assign n921 = n920 ^ n270 ;
  assign n922 = x8 & n921 ;
  assign n923 = n922 ^ n921 ;
  assign n924 = n923 ^ x2 ;
  assign n925 = n924 ^ x5 ;
  assign n926 = n101 & n925 ;
  assign n927 = n926 ^ x1 ;
  assign n928 = n917 & n927 ;
  assign n929 = n928 ^ n927 ;
  assign n930 = n929 ^ x1 ;
  assign n931 = n930 ^ x0 ;
  assign n932 = x0 & ~x9 ;
  assign n933 = n361 ^ x6 ;
  assign n934 = n933 ^ n766 ;
  assign n940 = x6 & n933 ;
  assign n935 = x1 & x6 ;
  assign n936 = n935 ^ x1 ;
  assign n937 = n936 ^ x6 ;
  assign n938 = n358 & ~n937 ;
  assign n939 = n938 ^ n937 ;
  assign n941 = n940 ^ n939 ;
  assign n942 = n934 & ~n941 ;
  assign n943 = n942 ^ n940 ;
  assign n944 = n932 & n943 ;
  assign n945 = n944 ^ x0 ;
  assign n946 = n931 & n945 ;
  assign n947 = n946 ^ n931 ;
  assign n948 = n947 ^ n945 ;
  assign n949 = n948 ^ n944 ;
  assign n950 = n949 ^ n930 ;
  assign n951 = n950 ^ x0 ;
  assign n952 = x9 & n125 ;
  assign n953 = n952 ^ n125 ;
  assign n954 = n61 & n953 ;
  assign n963 = n806 ^ x5 ;
  assign n964 = n963 ^ x9 ;
  assign n965 = n546 & n964 ;
  assign n966 = n965 ^ n964 ;
  assign n967 = n966 ^ n546 ;
  assign n968 = n967 ^ n964 ;
  assign n969 = n968 ^ n546 ;
  assign n970 = x2 & n969 ;
  assign n971 = n970 ^ x2 ;
  assign n972 = n971 ^ x2 ;
  assign n973 = n972 ^ x2 ;
  assign n974 = n973 ^ n969 ;
  assign n955 = x6 & n303 ;
  assign n956 = n955 ^ n303 ;
  assign n957 = n673 ^ x8 ;
  assign n958 = n957 ^ n557 ;
  assign n959 = n557 ^ x8 ;
  assign n960 = n958 & n959 ;
  assign n961 = n960 ^ n557 ;
  assign n962 = n956 & n961 ;
  assign n975 = n974 ^ n962 ;
  assign n976 = n962 ^ x3 ;
  assign n977 = x3 & n976 ;
  assign n978 = n977 ^ n976 ;
  assign n979 = n978 ^ x3 ;
  assign n980 = n979 ^ n974 ;
  assign n981 = n975 & n980 ;
  assign n982 = n981 ^ n975 ;
  assign n983 = n982 ^ n980 ;
  assign n984 = n983 ^ n978 ;
  assign n985 = n984 ^ n974 ;
  assign n986 = n954 & ~n985 ;
  assign n987 = n986 ^ n954 ;
  assign n988 = n987 ^ n954 ;
  assign n989 = n988 ^ n985 ;
  assign n992 = n766 ^ x5 ;
  assign n990 = x6 ^ x2 ;
  assign n991 = n990 ^ n766 ;
  assign n993 = n992 ^ n991 ;
  assign n995 = n993 ^ x6 ;
  assign n994 = n993 ^ n991 ;
  assign n996 = n995 ^ n994 ;
  assign n997 = n993 ^ n766 ;
  assign n998 = n997 ^ n995 ;
  assign n999 = n996 & n998 ;
  assign n1000 = n999 ^ n996 ;
  assign n1001 = n993 & n995 ;
  assign n1002 = n1001 ^ n995 ;
  assign n1003 = n1000 & n1002 ;
  assign n1004 = n1003 ^ n1000 ;
  assign n1005 = n1004 ^ n1002 ;
  assign n1006 = n1005 ^ x6 ;
  assign n1007 = n1006 ^ n990 ;
  assign n1008 = n1007 ^ n993 ;
  assign n1009 = n1008 ^ n995 ;
  assign n1010 = x9 & n1009 ;
  assign n1011 = n1010 ^ x9 ;
  assign n1012 = n1011 ^ x9 ;
  assign n1020 = n361 ^ x9 ;
  assign n1022 = n1020 ^ x5 ;
  assign n1021 = n1020 ^ x9 ;
  assign n1023 = n1022 ^ n1021 ;
  assign n1024 = n1021 ^ n1020 ;
  assign n1025 = n1023 & n1024 ;
  assign n1026 = n1025 ^ n1021 ;
  assign n1027 = x6 & n1026 ;
  assign n1028 = n1027 ^ n1020 ;
  assign n1029 = n1028 ^ x5 ;
  assign n1030 = n1029 ^ x6 ;
  assign n1031 = n1030 ^ x9 ;
  assign n1014 = x3 & x6 ;
  assign n1015 = n1014 ^ x3 ;
  assign n1016 = x8 & n1015 ;
  assign n1013 = n125 & n499 ;
  assign n1017 = n1016 ^ n1013 ;
  assign n1018 = n1017 ^ x8 ;
  assign n1019 = n1018 ^ x8 ;
  assign n1032 = n1031 ^ n1019 ;
  assign n1040 = n1012 & n1032 ;
  assign n1041 = n1040 ^ n1012 ;
  assign n1042 = n1041 ^ n1032 ;
  assign n1033 = x1 & n1032 ;
  assign n1034 = n1033 ^ x1 ;
  assign n1035 = n1012 & n1034 ;
  assign n1036 = n1035 ^ n1034 ;
  assign n1037 = n1036 ^ x1 ;
  assign n1038 = n1037 ^ x1 ;
  assign n1039 = n1038 ^ x1 ;
  assign n1043 = n1042 ^ n1039 ;
  assign n1052 = ~n989 & n1043 ;
  assign n1053 = n1052 ^ n1043 ;
  assign n1054 = n1053 ^ n1043 ;
  assign n1055 = n1054 ^ n989 ;
  assign n1056 = n951 & ~n1055 ;
  assign n1057 = n1056 ^ n951 ;
  assign n1058 = n1057 ^ n1055 ;
  assign n1059 = n1058 ^ n951 ;
  assign n1060 = n1059 ^ n1055 ;
  assign n1061 = n1060 ^ n1055 ;
  assign n1044 = x4 & n1043 ;
  assign n1045 = n1044 ^ x4 ;
  assign n1046 = ~n989 & n1045 ;
  assign n1047 = n951 & n1046 ;
  assign n1048 = n1047 ^ n1046 ;
  assign n1049 = n1048 ^ x4 ;
  assign n1050 = n1049 ^ x4 ;
  assign n1051 = n1050 ^ x4 ;
  assign n1062 = n1061 ^ n1051 ;
  assign n1070 = n553 ^ x2 ;
  assign n1071 = n304 ^ x2 ;
  assign n1072 = n1070 & n1071 ;
  assign n1073 = n1072 ^ n1070 ;
  assign n1074 = n557 & n1073 ;
  assign n1075 = n1074 ^ n1073 ;
  assign n1085 = n1075 ^ n1073 ;
  assign n1067 = n557 ^ n303 ;
  assign n1068 = n1067 ^ x2 ;
  assign n1069 = n1067 & n1068 ;
  assign n1076 = n1075 ^ n1069 ;
  assign n1077 = n1076 ^ n1073 ;
  assign n1078 = n1077 ^ n1068 ;
  assign n1080 = n1073 ^ n1069 ;
  assign n1079 = n303 ^ x2 ;
  assign n1081 = n1080 ^ n1079 ;
  assign n1082 = n1078 & n1081 ;
  assign n1083 = n1082 ^ n1078 ;
  assign n1084 = n1083 ^ n1069 ;
  assign n1086 = n1085 ^ n1084 ;
  assign n1087 = n1086 ^ n1068 ;
  assign n1089 = x8 ^ x5 ;
  assign n1088 = x8 ^ x3 ;
  assign n1090 = n1089 ^ n1088 ;
  assign n1092 = x8 ^ x6 ;
  assign n1093 = n1092 ^ x8 ;
  assign n1091 = n1089 ^ x8 ;
  assign n1094 = n1093 ^ n1091 ;
  assign n1095 = n1091 ^ x8 ;
  assign n1096 = n1094 & ~n1095 ;
  assign n1097 = n1096 ^ n1091 ;
  assign n1098 = ~n1090 & ~n1097 ;
  assign n1099 = n1098 ^ n1089 ;
  assign n1100 = n1099 ^ x8 ;
  assign n1108 = n1087 & n1100 ;
  assign n1109 = n1108 ^ n1087 ;
  assign n1110 = n1109 ^ n1087 ;
  assign n1111 = n1110 ^ n1100 ;
  assign n1103 = x6 & n106 ;
  assign n1104 = ~n227 & ~n1103 ;
  assign n1112 = n1111 ^ n1104 ;
  assign n1113 = n1112 ^ n1104 ;
  assign n1116 = n1113 ^ n1104 ;
  assign n1107 = n1104 ^ x1 ;
  assign n1114 = n1113 ^ n1107 ;
  assign n1105 = ~x1 & n1104 ;
  assign n1101 = ~x1 & n1100 ;
  assign n1102 = ~n1087 & n1101 ;
  assign n1106 = n1105 ^ n1102 ;
  assign n1115 = n1114 ^ n1106 ;
  assign n1117 = n1116 ^ n1115 ;
  assign n1118 = n1117 ^ n1114 ;
  assign n1119 = n1118 ^ n1116 ;
  assign n1120 = n1119 ^ n1113 ;
  assign n1063 = x2 & n125 ;
  assign n1064 = ~x4 & ~n1063 ;
  assign n1065 = n1064 ^ x4 ;
  assign n1121 = n1120 ^ n1065 ;
  assign n1066 = n1065 ^ n1064 ;
  assign n1122 = n1121 ^ n1066 ;
  assign n1123 = n1121 ^ n1065 ;
  assign n1124 = ~n1122 & ~n1123 ;
  assign n1125 = n1124 ^ n1121 ;
  assign n1127 = ~x5 & ~n490 ;
  assign n1128 = n725 & ~n1127 ;
  assign n1129 = ~n162 & n1128 ;
  assign n1148 = x0 & ~n1129 ;
  assign n1149 = ~n1125 & n1148 ;
  assign n1150 = n1149 ^ x0 ;
  assign n1141 = n1064 & ~n1120 ;
  assign n1142 = n1141 ^ n1064 ;
  assign n1143 = n1142 ^ x4 ;
  assign n1137 = x4 & ~n162 ;
  assign n1138 = n1128 & n1137 ;
  assign n1133 = ~x4 & ~n162 ;
  assign n1134 = ~n1063 & n1133 ;
  assign n1135 = n1128 & n1134 ;
  assign n1136 = n1120 & n1135 ;
  assign n1139 = n1138 ^ n1136 ;
  assign n1140 = n1139 ^ n1129 ;
  assign n1144 = n1143 ^ n1140 ;
  assign n1145 = n1144 ^ n1129 ;
  assign n1151 = n1150 ^ n1145 ;
  assign n1146 = x7 & n1145 ;
  assign n1126 = x0 & x7 ;
  assign n1130 = n1126 & ~n1129 ;
  assign n1131 = ~n1125 & n1130 ;
  assign n1132 = n1131 ^ n1126 ;
  assign n1147 = n1146 ^ n1132 ;
  assign n1152 = n1151 ^ n1147 ;
  assign n1153 = n1062 & n1152 ;
  assign n1154 = n1153 ^ n1152 ;
  assign n1155 = n1154 ^ x7 ;
  assign n1156 = x2 & ~n226 ;
  assign n1157 = n1156 ^ x2 ;
  assign n1158 = ~x4 & n1157 ;
  assign n1159 = x4 ^ x3 ;
  assign n1160 = n610 & n1159 ;
  assign n1161 = ~n1158 & ~n1160 ;
  assign n1162 = ~x7 & n124 ;
  assign n1163 = ~n1161 & n1162 ;
  assign n1164 = x3 & ~x4 ;
  assign n1165 = ~n610 & n1164 ;
  assign n1166 = n610 & n724 ;
  assign n1167 = ~n1165 & ~n1166 ;
  assign n1168 = n1162 & ~n1167 ;
  assign n1287 = n675 ^ n15 ;
  assign n1289 = n1287 ^ n16 ;
  assign n1290 = n16 ^ x7 ;
  assign n1291 = n629 ^ x9 ;
  assign n1292 = n1291 ^ x9 ;
  assign n1293 = n1292 ^ n1289 ;
  assign n1294 = n1290 & n1293 ;
  assign n1295 = n1294 ^ n1290 ;
  assign n1296 = n1295 ^ x7 ;
  assign n1297 = n1296 ^ n1289 ;
  assign n1298 = n1289 & n1297 ;
  assign n1299 = n1298 ^ n1289 ;
  assign n1300 = n1299 ^ n1297 ;
  assign n1301 = n1300 ^ n1295 ;
  assign n1302 = n1301 ^ x7 ;
  assign n1288 = n1287 ^ n15 ;
  assign n1303 = n1302 ^ n1288 ;
  assign n1304 = n16 ^ n15 ;
  assign n1306 = n1287 ^ x7 ;
  assign n1305 = n1292 ^ n16 ;
  assign n1307 = n1306 ^ n1305 ;
  assign n1308 = n1304 & ~n1307 ;
  assign n1309 = n1308 ^ n1300 ;
  assign n1310 = n1309 ^ n1295 ;
  assign n1311 = ~n1303 & ~n1310 ;
  assign n1312 = n1311 ^ n1310 ;
  assign n1313 = n1312 ^ x9 ;
  assign n1314 = n1313 ^ n1291 ;
  assign n1315 = x0 & ~n1314 ;
  assign n1316 = n1315 ^ x0 ;
  assign n1317 = n1316 ^ x0 ;
  assign n1318 = n1317 ^ n1314 ;
  assign n1411 = n1318 ^ n883 ;
  assign n1383 = ~x3 & x7 ;
  assign n1169 = n13 ^ x2 ;
  assign n1327 = n1169 ^ n239 ;
  assign n1328 = x2 & ~n1169 ;
  assign n1329 = n1328 ^ n63 ;
  assign n1330 = ~n1327 & ~n1329 ;
  assign n1331 = n1330 ^ n1328 ;
  assign n1332 = x6 & n557 ;
  assign n1333 = n1332 ^ x6 ;
  assign n1334 = n397 & n1333 ;
  assign n1335 = n1334 ^ n1333 ;
  assign n1336 = x5 & ~x7 ;
  assign n1337 = n1335 & n1336 ;
  assign n1338 = n1337 ^ n1336 ;
  assign n1339 = n1331 & n1338 ;
  assign n1340 = n1339 ^ n1338 ;
  assign n1341 = n1340 ^ n1338 ;
  assign n1353 = x9 & n130 ;
  assign n1354 = n422 & n1353 ;
  assign n1346 = n813 ^ x5 ;
  assign n1347 = x2 & n1346 ;
  assign n1348 = n1347 ^ x2 ;
  assign n1349 = n1348 ^ x2 ;
  assign n1350 = n422 & ~n601 ;
  assign n1351 = n1349 & n1350 ;
  assign n1352 = n1351 ^ n1350 ;
  assign n1355 = n1354 ^ n1352 ;
  assign n1275 = n119 ^ x2 ;
  assign n1342 = n964 & n1275 ;
  assign n1343 = n1342 ^ n1275 ;
  assign n1344 = n1343 ^ n1275 ;
  assign n1345 = x8 & n1344 ;
  assign n1356 = n1355 ^ n1345 ;
  assign n1371 = n1341 & n1356 ;
  assign n1372 = n1371 ^ n1341 ;
  assign n1360 = ~x7 & ~n397 ;
  assign n1361 = n1333 & n1360 ;
  assign n1362 = n1361 ^ x7 ;
  assign n1363 = n1356 & ~n1362 ;
  assign n1364 = n1363 ^ n1362 ;
  assign n1365 = n1364 ^ x7 ;
  assign n1373 = n1372 ^ n1365 ;
  assign n1391 = n1383 ^ n1373 ;
  assign n1412 = n1411 ^ n1391 ;
  assign n1384 = n1383 ^ n883 ;
  assign n1396 = n1384 ^ n1373 ;
  assign n1385 = n1383 ^ n1318 ;
  assign n1386 = n1384 & ~n1385 ;
  assign n1387 = n1386 ^ n1384 ;
  assign n1388 = n1387 ^ n1318 ;
  assign n1319 = n81 & n422 ;
  assign n1320 = ~x2 & x7 ;
  assign n1321 = n808 & n1320 ;
  assign n1322 = ~n1319 & n1321 ;
  assign n1323 = n1322 ^ n1320 ;
  assign n1389 = n1388 ^ n1323 ;
  assign n1397 = n1396 ^ n1389 ;
  assign n1398 = n1323 ^ n883 ;
  assign n1399 = n1398 ^ n1388 ;
  assign n1400 = n1397 & ~n1399 ;
  assign n1390 = n1388 ^ n883 ;
  assign n1392 = n1391 ^ n1390 ;
  assign n1393 = ~n1389 & n1392 ;
  assign n1394 = n1393 ^ n1389 ;
  assign n1401 = n1400 ^ n1394 ;
  assign n1402 = n1401 ^ n1388 ;
  assign n1403 = n1402 ^ n1396 ;
  assign n1404 = n1394 ^ n1323 ;
  assign n1405 = n1404 ^ n1373 ;
  assign n1406 = ~n1403 & n1405 ;
  assign n1407 = n1406 ^ n1403 ;
  assign n1408 = n1407 ^ n1405 ;
  assign n1409 = n1408 ^ n1400 ;
  assign n1395 = n1394 ^ n1387 ;
  assign n1410 = n1409 ^ n1395 ;
  assign n1413 = n1412 ^ n1410 ;
  assign n1414 = n1413 ^ n1383 ;
  assign n1415 = n1414 ^ x7 ;
  assign n1324 = ~n1318 & n1323 ;
  assign n1325 = n1324 ^ n1318 ;
  assign n1326 = n1325 ^ n1323 ;
  assign n1366 = n883 & ~n1365 ;
  assign n1357 = n883 & n1356 ;
  assign n1358 = n1357 ^ n883 ;
  assign n1359 = n1341 & n1358 ;
  assign n1367 = n1366 ^ n1359 ;
  assign n1368 = ~n1326 & n1367 ;
  assign n1369 = n1368 ^ n1367 ;
  assign n1370 = n1369 ^ n1367 ;
  assign n1374 = n1373 ^ n1370 ;
  assign n1229 = n29 & n356 ;
  assign n1230 = ~x0 & ~n545 ;
  assign n1231 = ~n441 & ~n624 ;
  assign n1232 = ~n1230 & n1231 ;
  assign n1233 = ~n1229 & ~n1232 ;
  assign n1378 = ~x1 & n115 ;
  assign n1379 = n1233 & n1378 ;
  assign n1185 = n270 ^ x6 ;
  assign n1170 = n1169 ^ x5 ;
  assign n1171 = n1170 ^ x2 ;
  assign n1174 = n1171 ^ x5 ;
  assign n1175 = n1174 ^ x9 ;
  assign n1176 = n1175 ^ x6 ;
  assign n1177 = x9 & n1176 ;
  assign n1178 = n1177 ^ x6 ;
  assign n1179 = n1178 ^ x9 ;
  assign n1180 = x6 & n1179 ;
  assign n1181 = n1180 ^ x6 ;
  assign n1182 = n1181 ^ n1179 ;
  assign n1172 = n1171 ^ n270 ;
  assign n1173 = n270 & n1172 ;
  assign n1183 = n1182 ^ n1173 ;
  assign n1184 = n1183 ^ n1177 ;
  assign n1186 = n1185 ^ n1184 ;
  assign n1188 = n1182 ^ x6 ;
  assign n1187 = n1175 ^ x9 ;
  assign n1189 = n1188 ^ n1187 ;
  assign n1190 = ~n1186 & ~n1189 ;
  assign n1191 = n1190 ^ n1189 ;
  assign n1192 = n1191 ^ n1182 ;
  assign n1193 = n1192 ^ n1178 ;
  assign n1194 = n1193 ^ n13 ;
  assign n1195 = n1194 ^ x2 ;
  assign n1196 = n1195 ^ x5 ;
  assign n1197 = n1196 ^ n1170 ;
  assign n1198 = x8 & n1197 ;
  assign n1199 = n1198 ^ x8 ;
  assign n1200 = n1199 ^ n1197 ;
  assign n1219 = n16 ^ x6 ;
  assign n1205 = n16 ^ x9 ;
  assign n1212 = n1205 ^ x6 ;
  assign n1213 = ~n1205 & ~n1212 ;
  assign n1221 = n1213 ^ n422 ;
  assign n1201 = n423 ^ n422 ;
  assign n1202 = n1201 ^ n422 ;
  assign n1220 = n1202 ^ x6 ;
  assign n1222 = n1221 ^ n1220 ;
  assign n1223 = n1219 & ~n1222 ;
  assign n1207 = n1202 ^ n16 ;
  assign n1208 = n1207 ^ n1205 ;
  assign n1209 = n1205 ^ n1202 ;
  assign n1210 = n1209 ^ x6 ;
  assign n1211 = n1208 & n1210 ;
  assign n1214 = n1213 ^ n1211 ;
  assign n1215 = n1214 ^ n422 ;
  assign n1206 = n1205 ^ n16 ;
  assign n1216 = n1215 ^ n1206 ;
  assign n1217 = n1211 ^ n422 ;
  assign n1218 = ~n1216 & n1217 ;
  assign n1224 = n1223 ^ n1218 ;
  assign n1225 = n1224 ^ n1213 ;
  assign n1203 = n1202 ^ n422 ;
  assign n1204 = n1203 ^ x6 ;
  assign n1226 = n1225 ^ n1204 ;
  assign n1375 = x1 & n115 ;
  assign n1376 = n1226 & n1375 ;
  assign n1377 = n1200 & n1376 ;
  assign n1380 = n1379 ^ n1377 ;
  assign n1381 = ~n1374 & n1380 ;
  assign n1236 = n1200 & ~n1226 ;
  assign n1237 = n1236 ^ n1226 ;
  assign n1238 = n1237 ^ n1200 ;
  assign n1239 = n1238 ^ n1226 ;
  assign n1240 = n1239 ^ n1233 ;
  assign n1234 = x1 & n1233 ;
  assign n1227 = x1 & n1226 ;
  assign n1228 = n1200 & n1227 ;
  assign n1235 = n1234 ^ n1228 ;
  assign n1241 = n1240 ^ n1235 ;
  assign n1242 = n1241 ^ n1239 ;
  assign n1243 = n493 ^ x0 ;
  assign n1244 = n1243 ^ x6 ;
  assign n1245 = n63 & n1244 ;
  assign n1246 = n1245 ^ n63 ;
  assign n1247 = n1246 ^ n1244 ;
  assign n1248 = n1247 ^ n1244 ;
  assign n1249 = n143 & n733 ;
  assign n1250 = n1249 ^ n733 ;
  assign n1251 = ~n1248 & n1250 ;
  assign n1252 = n1251 ^ n733 ;
  assign n1256 = ~x9 & n224 ;
  assign n1254 = n225 & n808 ;
  assign n1255 = n1254 ^ x0 ;
  assign n1257 = n1256 ^ n1255 ;
  assign n1265 = n1252 & n1257 ;
  assign n1266 = n1265 ^ n1252 ;
  assign n1267 = n1266 ^ n1257 ;
  assign n1253 = n1252 ^ x5 ;
  assign n1258 = n1257 ^ x5 ;
  assign n1259 = n1257 & ~n1258 ;
  assign n1260 = n1259 ^ x5 ;
  assign n1261 = ~n1253 & ~n1260 ;
  assign n1262 = n1261 ^ n1259 ;
  assign n1263 = n1262 ^ n1252 ;
  assign n1264 = n1263 ^ x5 ;
  assign n1268 = n1267 ^ n1264 ;
  assign n1269 = n1268 ^ n153 ;
  assign n1274 = x1 & ~x8 ;
  assign n1276 = n1274 & ~n1275 ;
  assign n1273 = n120 & n526 ;
  assign n1277 = n1276 ^ n1273 ;
  assign n1278 = x9 & n1277 ;
  assign n1270 = ~x0 & ~x8 ;
  assign n1271 = ~n74 & n101 ;
  assign n1272 = ~n1270 & n1271 ;
  assign n1279 = n1278 ^ n1272 ;
  assign n1280 = n1279 ^ n153 ;
  assign n1281 = n1279 & ~n1280 ;
  assign n1282 = n1281 ^ n153 ;
  assign n1283 = n1269 & ~n1282 ;
  assign n1284 = n1283 ^ n1281 ;
  assign n1285 = n1284 ^ n1268 ;
  assign n1286 = n1242 & n1285 ;
  assign n1382 = n1381 ^ n1286 ;
  assign n1416 = n1415 ^ n1382 ;
  assign n1417 = x4 & ~n226 ;
  assign n1418 = ~n106 & n1417 ;
  assign n1419 = ~n124 & ~n1418 ;
  assign n1420 = ~x7 & ~n1419 ;
  assign n1421 = ~x4 & ~n1420 ;
  assign n1422 = ~n1416 & n1421 ;
  assign n1423 = n1422 ^ n1421 ;
  assign n1424 = n1423 ^ n1421 ;
  assign n1425 = n1424 ^ n1420 ;
  assign n1459 = n84 & n499 ;
  assign n1460 = n1459 ^ n499 ;
  assign n1461 = n1460 ^ n499 ;
  assign n1456 = x2 & x5 ;
  assign n1457 = n494 & n1456 ;
  assign n1455 = x8 & n120 ;
  assign n1458 = n1457 ^ n1455 ;
  assign n1462 = n1461 ^ n1458 ;
  assign n1463 = x3 & n1462 ;
  assign n1464 = n1463 ^ n1462 ;
  assign n1465 = n192 & n624 ;
  assign n1466 = n1465 ^ n192 ;
  assign n1477 = ~n1464 & ~n1466 ;
  assign n1441 = n239 ^ x9 ;
  assign n1442 = ~x0 & n1441 ;
  assign n1443 = n1442 ^ x9 ;
  assign n1444 = n1443 ^ x0 ;
  assign n1445 = x9 & ~n1444 ;
  assign n1440 = x5 & n361 ;
  assign n1446 = n1445 ^ n1440 ;
  assign n1447 = n1446 ^ n1442 ;
  assign n1448 = n1447 ^ n303 ;
  assign n1450 = n1445 ^ x9 ;
  assign n1449 = n239 ^ x0 ;
  assign n1451 = n1450 ^ n1449 ;
  assign n1452 = n1448 & ~n1451 ;
  assign n1453 = n1452 ^ n1445 ;
  assign n1454 = n1453 ^ n1443 ;
  assign n1467 = x8 & n1466 ;
  assign n1468 = n1467 ^ x8 ;
  assign n1469 = n1468 ^ n1466 ;
  assign n1470 = n1464 & n1469 ;
  assign n1471 = n1470 ^ n1464 ;
  assign n1472 = n1471 ^ n1469 ;
  assign n1473 = n1454 & n1472 ;
  assign n1474 = n1473 ^ n1454 ;
  assign n1475 = n1474 ^ n1472 ;
  assign n1476 = n1475 ^ n1472 ;
  assign n1478 = n1477 ^ n1476 ;
  assign n1436 = x8 & n806 ;
  assign n1437 = n79 & n1436 ;
  assign n1479 = x1 & ~x6 ;
  assign n1480 = ~n1437 & n1479 ;
  assign n1481 = ~n1478 & n1480 ;
  assign n1482 = n1481 ^ n1480 ;
  assign n1426 = x2 & ~n808 ;
  assign n1427 = n49 & n1426 ;
  assign n1428 = ~n79 & n557 ;
  assign n1429 = ~n49 & n666 ;
  assign n1430 = n1429 ^ x5 ;
  assign n1431 = n1428 & n1430 ;
  assign n1432 = n1431 ^ n1430 ;
  assign n1433 = n1427 & n1432 ;
  assign n1434 = n1433 ^ n1427 ;
  assign n1435 = n1434 ^ n1432 ;
  assign n1438 = ~n937 & ~n1437 ;
  assign n1439 = ~n1435 & n1438 ;
  assign n1483 = n1482 ^ n1439 ;
  assign n1484 = n1483 ^ x6 ;
  assign n1510 = ~n181 & n883 ;
  assign n1494 = n1449 ^ n557 ;
  assign n1487 = ~n1441 & n1449 ;
  assign n1488 = n1487 ^ x9 ;
  assign n1489 = n1488 ^ x7 ;
  assign n1495 = n1494 ^ n1489 ;
  assign n1496 = x7 ^ x0 ;
  assign n1497 = n1496 ^ n1488 ;
  assign n1498 = ~n1495 & ~n1497 ;
  assign n1490 = n1488 ^ x0 ;
  assign n1485 = n557 ^ n239 ;
  assign n1491 = n1490 ^ n1485 ;
  assign n1492 = ~n1489 & ~n1491 ;
  assign n1499 = n1498 ^ n1492 ;
  assign n1500 = n1499 ^ n1488 ;
  assign n1501 = n1500 ^ n1494 ;
  assign n1502 = n1492 ^ x7 ;
  assign n1503 = n1502 ^ n557 ;
  assign n1504 = ~n1501 & n1503 ;
  assign n1505 = n1504 ^ n1498 ;
  assign n1493 = n1492 ^ n1487 ;
  assign n1506 = n1505 ^ n1493 ;
  assign n1486 = n1485 ^ n13 ;
  assign n1507 = n1506 ^ n1486 ;
  assign n1508 = n1507 ^ n557 ;
  assign n1509 = n1508 ^ n557 ;
  assign n1511 = n1510 ^ n1509 ;
  assign n1512 = n1510 ^ n803 ;
  assign n1513 = ~n803 & ~n1512 ;
  assign n1514 = n1513 ^ n803 ;
  assign n1515 = n1514 ^ n1509 ;
  assign n1516 = ~n1511 & n1515 ;
  assign n1517 = n1516 ^ n1513 ;
  assign n1518 = n1517 ^ n1509 ;
  assign n1519 = n1484 & n1518 ;
  assign n1589 = ~x3 & ~x6 ;
  assign n1590 = x8 & n1589 ;
  assign n1591 = n1590 ^ x6 ;
  assign n1587 = ~x9 & n545 ;
  assign n1585 = x9 & n423 ;
  assign n1583 = ~x6 & ~n51 ;
  assign n1584 = n499 & n1583 ;
  assign n1586 = n1585 ^ n1584 ;
  assign n1588 = n1587 ^ n1586 ;
  assign n1592 = n1591 ^ n1588 ;
  assign n1542 = n910 ^ x8 ;
  assign n1593 = ~n601 & n1542 ;
  assign n1594 = n1593 ^ n601 ;
  assign n1595 = ~x2 & n1594 ;
  assign n1596 = ~n1592 & n1595 ;
  assign n1558 = x3 & n490 ;
  assign n1559 = n1558 ^ x3 ;
  assign n1560 = ~x6 & ~n422 ;
  assign n1561 = ~n1559 & n1560 ;
  assign n1562 = n1561 ^ x6 ;
  assign n1567 = n557 ^ x3 ;
  assign n1568 = n1567 ^ x2 ;
  assign n1569 = n1567 & n1568 ;
  assign n1563 = n671 ^ x2 ;
  assign n1564 = ~n1070 & n1563 ;
  assign n1565 = ~n557 & n1564 ;
  assign n1570 = n1569 ^ n1565 ;
  assign n1571 = n1570 ^ n1564 ;
  assign n1572 = n1571 ^ n1568 ;
  assign n1574 = x3 ^ x2 ;
  assign n1573 = n1569 ^ n1564 ;
  assign n1575 = n1574 ^ n1573 ;
  assign n1576 = n1572 & ~n1575 ;
  assign n1577 = n1576 ^ n1569 ;
  assign n1566 = n1565 ^ n1564 ;
  assign n1578 = n1577 ^ n1566 ;
  assign n1579 = n1578 ^ n1568 ;
  assign n1580 = n1579 ^ x2 ;
  assign n1581 = ~n1562 & n1580 ;
  assign n1582 = n1581 ^ n1580 ;
  assign n1597 = n1596 ^ n1582 ;
  assign n1553 = x3 & ~n358 ;
  assign n1554 = n600 & n1553 ;
  assign n1598 = n813 & ~n1554 ;
  assign n1599 = n1597 & n1598 ;
  assign n1520 = n538 & n557 ;
  assign n1521 = n1520 ^ n538 ;
  assign n1522 = n561 ^ n557 ;
  assign n1523 = n1522 ^ n675 ;
  assign n1524 = n677 & n1523 ;
  assign n1525 = n1524 ^ n1523 ;
  assign n1526 = n1525 ^ n675 ;
  assign n1527 = ~n35 & n1526 ;
  assign n1528 = n1527 ^ n35 ;
  assign n1529 = n1521 & ~n1528 ;
  assign n1530 = n1529 ^ n1521 ;
  assign n1531 = n1530 ^ n1528 ;
  assign n1532 = x3 & ~n1531 ;
  assign n1533 = n1532 ^ x3 ;
  assign n1534 = n1533 ^ x3 ;
  assign n1535 = ~x9 & ~n561 ;
  assign n1536 = n990 ^ x6 ;
  assign n1537 = n1536 ^ x6 ;
  assign n1538 = n1536 ^ n1092 ;
  assign n1539 = ~n1537 & n1538 ;
  assign n1540 = n1539 ^ n1536 ;
  assign n1541 = n1535 & ~n1540 ;
  assign n1543 = x6 & n1542 ;
  assign n1544 = n1543 ^ n1542 ;
  assign n1545 = n831 & n1544 ;
  assign n1546 = n1545 ^ n831 ;
  assign n1547 = n1541 & n1546 ;
  assign n1548 = n1547 ^ n1541 ;
  assign n1549 = n1548 ^ n1546 ;
  assign n1550 = n1534 & n1549 ;
  assign n1551 = n1550 ^ n1534 ;
  assign n1552 = n1551 ^ n1549 ;
  assign n1555 = ~n1346 & ~n1554 ;
  assign n1556 = n1552 & n1555 ;
  assign n1557 = n1556 ^ n1555 ;
  assign n1600 = n1599 ^ n1557 ;
  assign n1601 = n1600 ^ x5 ;
  assign n1614 = n1519 & n1601 ;
  assign n1607 = ~x4 & x7 ;
  assign n1608 = n1509 & n1510 ;
  assign n1609 = n1608 ^ n1510 ;
  assign n1610 = n1607 & ~n1609 ;
  assign n1611 = n1610 ^ x4 ;
  assign n1615 = n1614 ^ n1611 ;
  assign n1602 = ~x5 & ~x7 ;
  assign n1603 = n1166 & n1602 ;
  assign n1604 = ~x6 & n1603 ;
  assign n1612 = n1604 & n1611 ;
  assign n1605 = n1601 & n1604 ;
  assign n1606 = n1519 & n1605 ;
  assign n1613 = n1612 ^ n1606 ;
  assign n1616 = n1615 ^ n1613 ;
  assign n1716 = n1603 ^ n615 ;
  assign n1718 = n557 ^ x2 ;
  assign n1717 = n629 ^ n557 ;
  assign n1719 = n1718 ^ n1717 ;
  assign n1721 = n1719 ^ x9 ;
  assign n1720 = n1719 ^ n1717 ;
  assign n1722 = n1721 ^ n1720 ;
  assign n1729 = n1722 ^ n1721 ;
  assign n1726 = n629 ^ x0 ;
  assign n1727 = n1726 ^ n557 ;
  assign n1724 = n1719 ^ n557 ;
  assign n1725 = n1724 ^ n1721 ;
  assign n1728 = n1727 ^ n1725 ;
  assign n1730 = n1729 ^ n1728 ;
  assign n1731 = n1725 ^ n1722 ;
  assign n1732 = n1725 ^ n1719 ;
  assign n1733 = ~n1731 & ~n1732 ;
  assign n1734 = n1733 ^ n1721 ;
  assign n1735 = n1734 ^ n1732 ;
  assign n1736 = n1730 & ~n1735 ;
  assign n1737 = n1736 ^ n1733 ;
  assign n1723 = n1722 ^ n1719 ;
  assign n1738 = n1737 ^ n1723 ;
  assign n1739 = n1721 ^ n1719 ;
  assign n1740 = n1739 ^ n1722 ;
  assign n1741 = n1740 ^ n1728 ;
  assign n1742 = ~n1727 & n1741 ;
  assign n1743 = n1742 ^ n1736 ;
  assign n1744 = n1743 ^ n1721 ;
  assign n1745 = n1744 ^ n1731 ;
  assign n1746 = n1738 & ~n1745 ;
  assign n1747 = n1746 ^ n1736 ;
  assign n1748 = n1747 ^ n1721 ;
  assign n1749 = n1748 ^ n1731 ;
  assign n1750 = n1749 ^ n629 ;
  assign n1751 = n1750 ^ n629 ;
  assign n1752 = n1751 ^ n1727 ;
  assign n1753 = n1752 ^ n615 ;
  assign n1754 = ~n1752 & n1753 ;
  assign n1755 = n1754 ^ n615 ;
  assign n1756 = ~n1716 & ~n1755 ;
  assign n1757 = n1756 ^ n1754 ;
  assign n1758 = n1757 ^ n1603 ;
  assign n1761 = x7 & ~n1758 ;
  assign n1652 = n143 & n192 ;
  assign n1653 = n1652 ^ n143 ;
  assign n1654 = x8 & n1653 ;
  assign n1655 = n1654 ^ x8 ;
  assign n1663 = ~x3 & ~x5 ;
  assign n1664 = n843 & n1663 ;
  assign n1656 = ~x1 & n270 ;
  assign n1657 = n371 ^ x5 ;
  assign n1658 = n1657 ^ n361 ;
  assign n1659 = n1657 ^ x5 ;
  assign n1660 = ~n1658 & n1659 ;
  assign n1661 = n1660 ^ n1657 ;
  assign n1662 = n1656 & n1661 ;
  assign n1665 = n1664 ^ n1662 ;
  assign n1679 = n1655 & n1665 ;
  assign n1680 = n1679 ^ n1655 ;
  assign n1668 = x8 & n74 ;
  assign n1669 = n1653 & n1668 ;
  assign n1677 = n1665 & n1669 ;
  assign n1678 = n1677 ^ n1669 ;
  assign n1681 = n1680 ^ n1678 ;
  assign n1672 = n442 & n1653 ;
  assign n1673 = n1672 ^ x8 ;
  assign n1682 = n1681 ^ n1673 ;
  assign n1674 = x9 & n1673 ;
  assign n1666 = x9 & ~n1665 ;
  assign n1670 = n1666 & ~n1669 ;
  assign n1667 = ~n1655 & n1666 ;
  assign n1671 = n1670 ^ n1667 ;
  assign n1675 = n1674 ^ n1671 ;
  assign n1676 = n1675 ^ x9 ;
  assign n1683 = n1682 ^ n1676 ;
  assign n1638 = n1456 ^ x2 ;
  assign n1639 = ~n192 & ~n1638 ;
  assign n1640 = n11 & ~n369 ;
  assign n1641 = n1640 ^ x1 ;
  assign n1642 = n1639 & n1641 ;
  assign n1643 = n1642 ^ n1641 ;
  assign n1644 = n73 ^ x5 ;
  assign n1645 = n369 & n1644 ;
  assign n1646 = n1645 ^ n369 ;
  assign n1647 = x9 & n452 ;
  assign n1648 = n1646 & n1647 ;
  assign n1649 = n1648 ^ x9 ;
  assign n1650 = n1643 & n1649 ;
  assign n1651 = n1650 ^ n1649 ;
  assign n1684 = n1683 ^ n1651 ;
  assign n1689 = ~x6 & n1684 ;
  assign n1617 = n515 ^ n194 ;
  assign n1618 = ~x2 & n102 ;
  assign n1619 = ~n221 & n1618 ;
  assign n1620 = ~n1617 & n1619 ;
  assign n1621 = n1456 ^ x5 ;
  assign n1624 = n1621 ^ x9 ;
  assign n1622 = n1621 ^ x3 ;
  assign n1623 = n1622 ^ n1621 ;
  assign n1625 = n1624 ^ n1623 ;
  assign n1626 = n1623 ^ n1621 ;
  assign n1627 = ~n1625 & ~n1626 ;
  assign n1628 = n1627 ^ n1623 ;
  assign n1629 = ~x0 & ~n733 ;
  assign n1630 = ~n1628 & n1629 ;
  assign n1631 = n733 & n1346 ;
  assign n1632 = n80 & ~n1631 ;
  assign n1633 = n1630 & n1632 ;
  assign n1634 = n1633 ^ n1630 ;
  assign n1635 = n1634 ^ n1632 ;
  assign n1636 = n1620 & ~n1635 ;
  assign n1637 = n1636 ^ n1635 ;
  assign n1685 = n546 & ~n1684 ;
  assign n1686 = n1685 ^ n1684 ;
  assign n1687 = ~n1637 & ~n1686 ;
  assign n1688 = n1687 ^ n1686 ;
  assign n1690 = n1689 ^ n1688 ;
  assign n1691 = ~x2 & x6 ;
  assign n1694 = n423 ^ x9 ;
  assign n1695 = n1694 ^ n423 ;
  assign n1692 = n423 ^ x1 ;
  assign n1693 = n1692 ^ n423 ;
  assign n1696 = n1695 ^ n1693 ;
  assign n1697 = n1693 ^ n423 ;
  assign n1698 = ~n1696 & ~n1697 ;
  assign n1699 = n1698 ^ n1693 ;
  assign n1700 = n1691 & n1699 ;
  assign n1701 = n1700 ^ x2 ;
  assign n1702 = n193 & ~n1701 ;
  assign n1703 = n1702 ^ n193 ;
  assign n1704 = ~x6 & ~n62 ;
  assign n1705 = ~n1255 & n1704 ;
  assign n1706 = ~x7 & ~n1705 ;
  assign n1707 = n1703 & n1706 ;
  assign n1708 = n1707 ^ x7 ;
  assign n1759 = ~n1708 & ~n1758 ;
  assign n1760 = n1690 & n1759 ;
  assign n1762 = n1761 ^ n1760 ;
  assign n1709 = ~x4 & ~n1603 ;
  assign n1712 = x7 & n1709 ;
  assign n1710 = ~n1708 & n1709 ;
  assign n1711 = n1690 & n1710 ;
  assign n1713 = n1712 ^ n1711 ;
  assign n1714 = n1713 ^ n1709 ;
  assign n1715 = n1714 ^ n1603 ;
  assign n1763 = n1762 ^ n1715 ;
  assign n1764 = x1 & n808 ;
  assign n1765 = n1764 ^ n808 ;
  assign n1766 = x2 & n1015 ;
  assign n1767 = ~x7 & n74 ;
  assign n1768 = n1766 & n1767 ;
  assign n1769 = n1768 ^ x7 ;
  assign n1770 = n1765 & ~n1769 ;
  assign n1771 = n1770 ^ n1765 ;
  assign n1772 = n1771 ^ n1769 ;
  assign n1773 = ~x2 & ~x7 ;
  assign n1774 = ~n181 & n1773 ;
  assign n1775 = n1774 ^ x7 ;
  assign n1776 = x0 & ~n1775 ;
  assign n1777 = n1776 ^ x0 ;
  assign n1778 = ~x5 & x6 ;
  assign n1779 = ~n80 & n1778 ;
  assign n1780 = n1779 ^ x6 ;
  assign n1781 = x2 & x4 ;
  assign n1782 = n1781 ^ x4 ;
  assign n1783 = n181 & n1782 ;
  assign n1784 = n1783 ^ n1782 ;
  assign n1785 = n1784 ^ x4 ;
  assign n1786 = x7 & n80 ;
  assign n1787 = n1786 ^ x7 ;
  assign n1788 = n1785 & n1787 ;
  assign n1789 = n1788 ^ n1785 ;
  assign n1790 = n1789 ^ n1787 ;
  assign n1791 = n1780 & n1790 ;
  assign n1792 = n1791 ^ n1780 ;
  assign n1793 = n1792 ^ n1790 ;
  assign n1794 = n1777 & n1793 ;
  assign n1795 = n1794 ^ n1777 ;
  assign n1796 = n1795 ^ n1793 ;
  assign n1797 = n1772 & n1796 ;
  assign n1798 = n1797 ^ n1772 ;
  assign n1799 = n1798 ^ n1796 ;
  assign n1844 = n1127 & n1766 ;
  assign n1845 = n806 & n907 ;
  assign n1846 = n1845 ^ x6 ;
  assign n1847 = x3 & ~n1846 ;
  assign n1848 = n1847 ^ x3 ;
  assign n1849 = n1848 ^ n1846 ;
  assign n1850 = n1844 & n1849 ;
  assign n1851 = n1850 ^ n1844 ;
  assign n1852 = n1851 ^ n1849 ;
  assign n1858 = n423 ^ x3 ;
  assign n1859 = n1858 ^ n423 ;
  assign n1874 = n1859 ^ x2 ;
  assign n1860 = n1859 ^ n423 ;
  assign n1867 = n1860 ^ x2 ;
  assign n1868 = n1860 & ~n1867 ;
  assign n1876 = n1868 ^ n599 ;
  assign n1853 = n964 ^ n599 ;
  assign n1854 = n1853 ^ n599 ;
  assign n1855 = n1854 ^ n599 ;
  assign n1875 = n1855 ^ x2 ;
  assign n1877 = n1876 ^ n1875 ;
  assign n1878 = n1874 & n1877 ;
  assign n1862 = n1859 ^ n1855 ;
  assign n1863 = n1862 ^ n1860 ;
  assign n1864 = n1860 ^ n1855 ;
  assign n1865 = n1864 ^ x2 ;
  assign n1866 = n1863 & n1865 ;
  assign n1869 = n1868 ^ n1866 ;
  assign n1870 = n1869 ^ n599 ;
  assign n1861 = n1860 ^ n1859 ;
  assign n1871 = n1870 ^ n1861 ;
  assign n1872 = n1866 ^ n599 ;
  assign n1873 = ~n1871 & n1872 ;
  assign n1879 = n1878 ^ n1873 ;
  assign n1880 = n1879 ^ n1868 ;
  assign n1856 = n1855 ^ n599 ;
  assign n1857 = n1856 ^ x2 ;
  assign n1881 = n1880 ^ n1857 ;
  assign n1882 = x1 & ~n1881 ;
  assign n1883 = ~n1852 & n1882 ;
  assign n1884 = n1883 ^ x1 ;
  assign n1887 = n1799 & n1884 ;
  assign n1888 = n1887 ^ n1884 ;
  assign n1889 = n1888 ^ n1799 ;
  assign n1807 = n423 ^ x6 ;
  assign n1808 = n1807 ^ n423 ;
  assign n1823 = n1808 ^ x3 ;
  assign n1809 = n1808 ^ n423 ;
  assign n1816 = n1809 ^ x3 ;
  assign n1817 = ~n1809 & ~n1816 ;
  assign n1825 = n1817 ^ n806 ;
  assign n1802 = n806 ^ x9 ;
  assign n1803 = n1802 ^ n806 ;
  assign n1804 = n1803 ^ n806 ;
  assign n1824 = n1804 ^ x3 ;
  assign n1826 = n1825 ^ n1824 ;
  assign n1827 = n1823 & ~n1826 ;
  assign n1811 = n1808 ^ n1804 ;
  assign n1812 = n1811 ^ n1809 ;
  assign n1813 = n1809 ^ n1804 ;
  assign n1814 = n1813 ^ x3 ;
  assign n1815 = n1812 & n1814 ;
  assign n1818 = n1817 ^ n1815 ;
  assign n1819 = n1818 ^ n806 ;
  assign n1810 = n1809 ^ n1808 ;
  assign n1820 = n1819 ^ n1810 ;
  assign n1821 = n1815 ^ n806 ;
  assign n1822 = ~n1820 & n1821 ;
  assign n1828 = n1827 ^ n1822 ;
  assign n1829 = n1828 ^ n1817 ;
  assign n1805 = n1804 ^ n806 ;
  assign n1806 = n1805 ^ x3 ;
  assign n1830 = n1829 ^ n1806 ;
  assign n1831 = n1830 ^ x3 ;
  assign n1832 = n724 & ~n883 ;
  assign n1833 = ~x2 & ~n1832 ;
  assign n1834 = ~n1831 & n1833 ;
  assign n1835 = n1834 ^ n1833 ;
  assign n1800 = n80 & n808 ;
  assign n1801 = ~n1127 & n1800 ;
  assign n1836 = n1835 ^ n1801 ;
  assign n1837 = n1801 ^ x1 ;
  assign n1838 = x1 & ~n1837 ;
  assign n1839 = n1838 ^ x1 ;
  assign n1840 = n1839 ^ n1835 ;
  assign n1841 = n1836 & ~n1840 ;
  assign n1842 = n1841 ^ n1838 ;
  assign n1843 = n1842 ^ n1835 ;
  assign n1885 = n1843 & ~n1884 ;
  assign n1886 = ~n1799 & n1885 ;
  assign n1890 = n1889 ^ n1886 ;
  assign n1891 = ~x7 & n883 ;
  assign n1892 = x8 & ~n191 ;
  assign n1893 = x1 & n24 ;
  assign n1894 = n1893 ^ x1 ;
  assign n1895 = n1894 ^ n24 ;
  assign n1896 = x2 & n1164 ;
  assign n1897 = n1895 & n1896 ;
  assign n1898 = ~n1892 & n1897 ;
  assign n1899 = ~n1166 & ~n1898 ;
  assign n1900 = n1891 & ~n1899 ;
  assign y0 = n355 ;
  assign y1 = ~n663 ;
  assign y2 = ~n899 ;
  assign y3 = ~n1155 ;
  assign y4 = n1163 ;
  assign y5 = n1168 ;
  assign y6 = ~n1425 ;
  assign y7 = n1616 ;
  assign y8 = ~n1763 ;
  assign y9 = ~n1890 ;
  assign y10 = n1900 ;
endmodule
