module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 ;
  assign n33 = x29 & x30 ;
  assign n34 = x27 & x28 ;
  assign n35 = n33 & n34 ;
  assign n36 = x26 & x27 ;
  assign n37 = n35 & n36 ;
  assign n38 = x22 & x23 ;
  assign n39 = x23 & x24 ;
  assign n40 = n38 & n39 ;
  assign n41 = x25 & x26 ;
  assign n42 = x24 & x25 ;
  assign n43 = n41 & n42 ;
  assign n44 = n40 & n43 ;
  assign n45 = ~n37 & ~n44 ;
  assign n46 = n34 & n36 ;
  assign n47 = n43 & n46 ;
  assign n48 = ~n45 & n47 ;
  assign n49 = x28 & x29 ;
  assign n50 = x30 & x31 ;
  assign n51 = n49 & n50 ;
  assign n52 = n34 & n51 ;
  assign n53 = n36 & n41 ;
  assign n54 = n39 & n42 ;
  assign n55 = n53 & n54 ;
  assign n56 = n52 & n55 ;
  assign n57 = n56 ^ n52 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n34 & n49 ;
  assign n60 = n53 & n59 ;
  assign n61 = ~n58 & n60 ;
  assign n62 = n61 ^ n60 ;
  assign n63 = n48 & n62 ;
  assign n64 = x10 & x11 ;
  assign n65 = x17 & x18 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = x12 & x13 ;
  assign n68 = x13 & x14 ;
  assign n69 = n67 & n68 ;
  assign n70 = x14 & x15 ;
  assign n71 = x15 & x16 ;
  assign n72 = n70 & n71 ;
  assign n73 = n69 & n72 ;
  assign n74 = n66 & n73 ;
  assign n75 = n74 ^ n73 ;
  assign n76 = x16 & x17 ;
  assign n77 = n71 & n76 ;
  assign n78 = x19 & x20 ;
  assign n79 = n65 & n78 ;
  assign n80 = n77 & n79 ;
  assign n81 = n75 & n80 ;
  assign n82 = n81 ^ n75 ;
  assign n83 = n82 ^ n80 ;
  assign n84 = x18 & x19 ;
  assign n85 = x11 & x12 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = n68 & n70 ;
  assign n88 = n77 & n87 ;
  assign n89 = n86 & n88 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = ~n83 & n90 ;
  assign n92 = n91 ^ n90 ;
  assign n93 = x21 & x22 ;
  assign n94 = ~n70 & ~n93 ;
  assign n95 = n78 & n84 ;
  assign n96 = n65 & n76 ;
  assign n97 = n95 & n96 ;
  assign n98 = n94 & n97 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = n65 & n84 ;
  assign n101 = n77 & n100 ;
  assign n102 = x20 & x21 ;
  assign n103 = n84 & n102 ;
  assign n104 = n96 & n103 ;
  assign n105 = n101 & n104 ;
  assign n106 = n99 & n105 ;
  assign n107 = n92 & n106 ;
  assign n108 = n107 ^ n92 ;
  assign n109 = n108 ^ n106 ;
  assign n110 = n63 & ~n109 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = n78 & n93 ;
  assign n113 = n95 & n112 ;
  assign n114 = n38 & n102 ;
  assign n115 = n113 & n114 ;
  assign n116 = n65 & n103 ;
  assign n117 = n115 & n116 ;
  assign n118 = ~n39 & ~n76 ;
  assign n119 = n117 & ~n118 ;
  assign n120 = ~n41 & ~n84 ;
  assign n121 = n39 & n93 ;
  assign n122 = n102 & n121 ;
  assign n123 = ~n120 & n122 ;
  assign n124 = n34 & n41 ;
  assign n125 = n54 & n124 ;
  assign n126 = ~n123 & ~n125 ;
  assign n127 = ~n36 & ~n78 ;
  assign n128 = n38 & n93 ;
  assign n129 = n54 & n128 ;
  assign n130 = ~n127 & n129 ;
  assign n131 = ~n126 & n130 ;
  assign n132 = ~n119 & ~n131 ;
  assign n133 = ~n111 & n132 ;
  assign n155 = n68 & n71 ;
  assign n156 = n67 & n85 ;
  assign n157 = n155 & n156 ;
  assign n134 = x8 & x9 ;
  assign n135 = x7 & n134 ;
  assign n136 = x9 & x10 ;
  assign n137 = n85 & n136 ;
  assign n138 = n135 & n137 ;
  assign n139 = x7 & x8 ;
  assign n140 = n136 & n139 ;
  assign n141 = x6 & x7 ;
  assign n142 = n139 & n141 ;
  assign n143 = n140 & n142 ;
  assign n144 = n138 & n143 ;
  assign n145 = n64 & n136 ;
  assign n146 = n68 & n85 ;
  assign n147 = n145 & n146 ;
  assign n148 = n134 & n136 ;
  assign n149 = n64 & n85 ;
  assign n150 = n148 & n149 ;
  assign n151 = n147 & n150 ;
  assign n152 = n144 & n151 ;
  assign n153 = n152 ^ n144 ;
  assign n154 = n153 ^ n151 ;
  assign n158 = n157 ^ n154 ;
  assign n159 = n145 & n156 ;
  assign n160 = ~n70 & ~n139 ;
  assign n161 = n159 & n160 ;
  assign n162 = n161 ^ n159 ;
  assign n163 = n162 ^ n157 ;
  assign n164 = ~n162 & n163 ;
  assign n165 = n164 ^ n162 ;
  assign n166 = n165 ^ n154 ;
  assign n167 = n158 & n166 ;
  assign n168 = n167 ^ n164 ;
  assign n169 = n168 ^ n154 ;
  assign n170 = x4 & x5 ;
  assign n171 = x3 & x4 ;
  assign n172 = n170 & n171 ;
  assign n173 = x5 & x6 ;
  assign n174 = n139 & n173 ;
  assign n175 = n172 & n174 ;
  assign n176 = n170 & n173 ;
  assign n177 = x2 & x3 ;
  assign n178 = n171 & n177 ;
  assign n179 = n176 & n178 ;
  assign n180 = n175 & n179 ;
  assign n181 = n134 & n141 ;
  assign n182 = n173 & n181 ;
  assign n183 = n140 & n182 ;
  assign n184 = n170 & n177 ;
  assign n185 = x1 & x2 ;
  assign n186 = n171 & n185 ;
  assign n187 = x0 & x1 ;
  assign n188 = n186 & n187 ;
  assign n189 = n184 & n188 ;
  assign n190 = n183 & n189 ;
  assign n191 = n190 ^ n183 ;
  assign n192 = n191 ^ n189 ;
  assign n193 = n180 & ~n192 ;
  assign n194 = n193 ^ n192 ;
  assign n195 = n141 & n173 ;
  assign n196 = n172 & n195 ;
  assign n197 = n176 & n181 ;
  assign n198 = n196 & n197 ;
  assign n199 = n177 & n185 ;
  assign n200 = n172 & n199 ;
  assign n201 = n141 & n170 ;
  assign n202 = n178 & n201 ;
  assign n203 = n200 & n202 ;
  assign n204 = n198 & n203 ;
  assign n205 = n204 ^ n198 ;
  assign n206 = n205 ^ n203 ;
  assign n207 = ~n194 & ~n206 ;
  assign n208 = n207 ^ n194 ;
  assign n209 = n208 ^ n206 ;
  assign n210 = n142 & n176 ;
  assign n211 = n183 & n210 ;
  assign n212 = n144 & n211 ;
  assign n213 = n212 ^ n144 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = n64 & n134 ;
  assign n216 = n143 & n215 ;
  assign n217 = n182 & n216 ;
  assign n218 = ~n214 & n217 ;
  assign n219 = n218 ^ n217 ;
  assign n220 = ~n209 & n219 ;
  assign n221 = n220 ^ n209 ;
  assign n222 = n221 ^ n219 ;
  assign n223 = n169 & n222 ;
  assign n224 = n223 ^ n222 ;
  assign n225 = n133 & n224 ;
  assign n527 = ~n48 & ~n62 ;
  assign n528 = ~n117 & n527 ;
  assign n529 = ~n206 & n211 ;
  assign n530 = n529 ^ n206 ;
  assign n531 = ~n154 & n217 ;
  assign n532 = n531 ^ n154 ;
  assign n533 = ~n530 & ~n532 ;
  assign n357 = n171 & n173 ;
  assign n465 = n199 & n357 ;
  assign n534 = n188 & n465 ;
  assign n535 = ~n105 & ~n123 ;
  assign n536 = ~n534 & n535 ;
  assign n537 = n90 & n99 ;
  assign n538 = n537 ^ n90 ;
  assign n539 = n538 ^ n99 ;
  assign n540 = n130 & ~n539 ;
  assign n541 = n540 ^ n539 ;
  assign n542 = n75 & n162 ;
  assign n543 = n542 ^ n75 ;
  assign n544 = n543 ^ n162 ;
  assign n545 = n180 & ~n544 ;
  assign n546 = n545 ^ n544 ;
  assign n547 = ~n541 & ~n546 ;
  assign n548 = n536 & n547 ;
  assign n549 = n533 & n548 ;
  assign n550 = n528 & n549 ;
  assign n466 = n125 & n465 ;
  assign n467 = n466 ^ n125 ;
  assign n468 = n467 ^ n465 ;
  assign n383 = n36 & n42 ;
  assign n469 = n40 & n383 ;
  assign n375 = n67 & n70 ;
  assign n470 = n149 & n375 ;
  assign n471 = n469 & n470 ;
  assign n472 = n471 ^ n469 ;
  assign n473 = n472 ^ n470 ;
  assign n474 = ~n468 & ~n473 ;
  assign n475 = n147 & n157 ;
  assign n476 = n475 ^ n147 ;
  assign n477 = n476 ^ n157 ;
  assign n478 = n80 & n104 ;
  assign n479 = n478 ^ n80 ;
  assign n480 = n479 ^ n104 ;
  assign n481 = ~n477 & ~n480 ;
  assign n482 = n474 & n481 ;
  assign n271 = ~x20 & ~x26 ;
  assign n483 = n129 & n271 ;
  assign n484 = n483 ^ n129 ;
  assign n444 = n72 & n96 ;
  assign n485 = ~x13 & ~x19 ;
  assign n486 = n444 & n485 ;
  assign n487 = n486 ^ n444 ;
  assign n488 = n484 & n487 ;
  assign n489 = n488 ^ n484 ;
  assign n490 = n489 ^ n487 ;
  assign n309 = x19 & n102 ;
  assign n491 = n121 & n309 ;
  assign n492 = n35 & n53 ;
  assign n493 = n491 & n492 ;
  assign n494 = n493 ^ n491 ;
  assign n495 = n494 ^ n492 ;
  assign n496 = ~n490 & ~n495 ;
  assign n497 = ~n192 & n496 ;
  assign n498 = n482 & n497 ;
  assign n499 = n112 & n116 ;
  assign n384 = n51 & n383 ;
  assign n385 = n384 ^ n51 ;
  assign n386 = n385 ^ n383 ;
  assign n398 = n36 & n49 ;
  assign n500 = ~n386 & n398 ;
  assign n501 = n500 ^ n398 ;
  assign n399 = n70 & n76 ;
  assign n502 = n399 ^ n67 ;
  assign n503 = ~n67 & n502 ;
  assign n504 = n503 ^ n67 ;
  assign n505 = n504 ^ n150 ;
  assign n506 = n399 ^ n150 ;
  assign n507 = n505 & n506 ;
  assign n508 = n507 ^ n503 ;
  assign n509 = n508 ^ n150 ;
  assign n510 = n501 & n509 ;
  assign n511 = n510 ^ n501 ;
  assign n512 = n511 ^ n509 ;
  assign n513 = n499 & ~n512 ;
  assign n514 = n513 ^ n512 ;
  assign n515 = n175 & n197 ;
  assign n516 = n515 ^ n175 ;
  assign n517 = n516 ^ n197 ;
  assign n518 = n138 & n202 ;
  assign n519 = n518 ^ n138 ;
  assign n520 = n519 ^ n202 ;
  assign n521 = ~n517 & ~n520 ;
  assign n522 = ~n115 & ~n216 ;
  assign n523 = n521 & n522 ;
  assign n524 = ~n514 & n523 ;
  assign n525 = n498 & n524 ;
  assign n415 = n179 & n196 ;
  assign n416 = n415 ^ n196 ;
  assign n417 = n416 ^ n179 ;
  assign n418 = n182 & ~n417 ;
  assign n419 = n418 ^ n417 ;
  assign n420 = ~n143 & ~n188 ;
  assign n421 = ~n419 & n420 ;
  assign n422 = n87 & n156 ;
  assign n423 = n150 & n422 ;
  assign n424 = n423 ^ n150 ;
  assign n425 = n424 ^ n422 ;
  assign n426 = n47 & n60 ;
  assign n427 = n426 ^ n47 ;
  assign n428 = n427 ^ n60 ;
  assign n429 = ~n425 & ~n428 ;
  assign n430 = n135 & n145 ;
  assign n431 = n200 & n430 ;
  assign n432 = n431 ^ n430 ;
  assign n433 = n432 ^ n200 ;
  assign n434 = n159 & n210 ;
  assign n435 = n434 ^ n159 ;
  assign n436 = n435 ^ n210 ;
  assign n437 = ~n433 & ~n436 ;
  assign n438 = n429 & n437 ;
  assign n439 = n421 & n438 ;
  assign n440 = n69 & n149 ;
  assign n441 = n129 & n440 ;
  assign n442 = n441 ^ n129 ;
  assign n443 = n442 ^ n440 ;
  assign n445 = n128 & n309 ;
  assign n446 = n444 & n445 ;
  assign n447 = n446 ^ n444 ;
  assign n448 = n447 ^ n445 ;
  assign n449 = ~n443 & ~n448 ;
  assign n450 = n73 & n101 ;
  assign n451 = n450 ^ n73 ;
  assign n452 = n451 ^ n101 ;
  assign n453 = n88 & n97 ;
  assign n454 = n453 ^ n88 ;
  assign n455 = n454 ^ n97 ;
  assign n456 = ~n452 & ~n455 ;
  assign n457 = n449 & n456 ;
  assign n458 = n45 & ~n58 ;
  assign n459 = ~n113 & ~n116 ;
  assign n460 = ~n122 & n459 ;
  assign n461 = n458 & n460 ;
  assign n462 = n457 & n461 ;
  assign n463 = n439 & n462 ;
  assign n346 = n38 & n42 ;
  assign n347 = n177 & n187 ;
  assign n348 = n346 & n347 ;
  assign n349 = n348 ^ n346 ;
  assign n350 = n349 ^ n347 ;
  assign n351 = n65 & n71 ;
  assign n352 = n64 & n67 ;
  assign n353 = n351 & n352 ;
  assign n354 = n353 ^ n352 ;
  assign n355 = n354 ^ n351 ;
  assign n356 = ~n350 & ~n355 ;
  assign n358 = n146 & n357 ;
  assign n359 = n358 ^ n357 ;
  assign n360 = n359 ^ n146 ;
  assign n361 = n124 & n174 ;
  assign n362 = n361 ^ n174 ;
  assign n363 = n362 ^ n124 ;
  assign n364 = ~n360 & ~n363 ;
  assign n365 = n356 & n364 ;
  assign n366 = n76 & n84 ;
  assign n367 = n201 & n366 ;
  assign n368 = n367 ^ n201 ;
  assign n369 = n368 ^ n366 ;
  assign n370 = n79 & ~n369 ;
  assign n371 = n370 ^ n369 ;
  assign n372 = n137 & n155 ;
  assign n373 = n372 ^ n155 ;
  assign n374 = n373 ^ n137 ;
  assign n376 = n39 & n41 ;
  assign n377 = n375 & n376 ;
  assign n378 = n377 ^ n376 ;
  assign n379 = n378 ^ n375 ;
  assign n380 = ~n374 & ~n379 ;
  assign n381 = ~n371 & n380 ;
  assign n382 = n365 & n381 ;
  assign n387 = n140 & n181 ;
  assign n388 = n387 ^ n140 ;
  assign n389 = n388 ^ n181 ;
  assign n390 = n184 & n186 ;
  assign n391 = n390 ^ n186 ;
  assign n392 = n391 ^ n184 ;
  assign n393 = ~n389 & ~n392 ;
  assign n394 = ~n386 & n393 ;
  assign n395 = n103 & n121 ;
  assign n396 = n395 ^ n103 ;
  assign n397 = n396 ^ n121 ;
  assign n400 = n398 & n399 ;
  assign n401 = n400 ^ n398 ;
  assign n402 = n401 ^ n399 ;
  assign n403 = ~n397 & ~n402 ;
  assign n404 = n35 & n215 ;
  assign n405 = n404 ^ n35 ;
  assign n406 = n405 ^ n215 ;
  assign n407 = n112 & n114 ;
  assign n408 = n407 ^ n112 ;
  assign n409 = n408 ^ n114 ;
  assign n410 = ~n406 & ~n409 ;
  assign n411 = n403 & n410 ;
  assign n412 = n394 & n411 ;
  assign n413 = n382 & n412 ;
  assign n285 = n44 ^ n40 ;
  assign n286 = n285 ^ n43 ;
  assign n287 = n33 & n50 ;
  assign n288 = n46 & n287 ;
  assign n289 = n288 ^ n46 ;
  assign n290 = n289 ^ n287 ;
  assign n291 = ~n286 & ~n290 ;
  assign n292 = n87 & n148 ;
  assign n293 = n292 ^ n87 ;
  assign n294 = n293 ^ n148 ;
  assign n295 = n33 & n49 ;
  assign n296 = n72 & n295 ;
  assign n297 = n296 ^ n72 ;
  assign n298 = n297 ^ n295 ;
  assign n299 = ~n294 & ~n298 ;
  assign n300 = n291 & n299 ;
  assign n272 = ~x0 & ~x3 ;
  assign n301 = n185 & ~n272 ;
  assign n302 = ~x15 & x16 ;
  assign n303 = x17 & ~x18 ;
  assign n304 = n302 & n303 ;
  assign n305 = n304 ^ n76 ;
  assign n306 = ~n301 & ~n305 ;
  assign n307 = n55 ^ n53 ;
  assign n308 = n307 ^ n54 ;
  assign n310 = n59 & n309 ;
  assign n311 = n310 ^ n59 ;
  assign n312 = n311 ^ n309 ;
  assign n313 = ~n308 & ~n312 ;
  assign n314 = n306 & n313 ;
  assign n315 = n300 & n314 ;
  assign n241 = ~n38 & ~n102 ;
  assign n316 = n93 & ~n241 ;
  assign n317 = ~x17 & x18 ;
  assign n318 = x19 & ~x20 ;
  assign n319 = n317 & n318 ;
  assign n320 = n319 ^ n84 ;
  assign n321 = n196 ^ n195 ;
  assign n322 = n321 ^ n172 ;
  assign n323 = n320 & ~n322 ;
  assign n324 = n323 ^ n322 ;
  assign n325 = n316 & ~n324 ;
  assign n326 = n325 ^ n324 ;
  assign n327 = ~x9 & x10 ;
  assign n328 = x11 & ~x12 ;
  assign n329 = n327 & n328 ;
  assign n330 = n329 ^ n64 ;
  assign n331 = ~x11 & x12 ;
  assign n332 = x13 & ~x14 ;
  assign n333 = n331 & n332 ;
  assign n334 = n333 ^ n67 ;
  assign n335 = ~n330 & ~n334 ;
  assign n336 = n210 ^ n142 ;
  assign n337 = n336 ^ n176 ;
  assign n338 = n135 & n178 ;
  assign n339 = n338 ^ n135 ;
  assign n340 = n339 ^ n178 ;
  assign n341 = ~n337 & ~n340 ;
  assign n342 = n335 & n341 ;
  assign n343 = ~n326 & n342 ;
  assign n344 = n315 & n343 ;
  assign n253 = ~x18 & ~x19 ;
  assign n254 = ~x21 & ~x22 ;
  assign n255 = n253 & n254 ;
  assign n256 = ~x14 & ~x15 ;
  assign n257 = ~x16 & ~x17 ;
  assign n258 = n256 & n257 ;
  assign n259 = n255 & n258 ;
  assign n260 = ~x28 & ~x29 ;
  assign n261 = ~x30 & ~x31 ;
  assign n262 = n260 & n261 ;
  assign n263 = ~x23 & ~x24 ;
  assign n264 = ~x25 & ~x27 ;
  assign n265 = n263 & n264 ;
  assign n266 = n262 & n265 ;
  assign n267 = n259 & n266 ;
  assign n268 = ~x1 & ~x2 ;
  assign n269 = ~x4 & ~x5 ;
  assign n270 = n268 & n269 ;
  assign n273 = n271 & n272 ;
  assign n274 = n270 & n273 ;
  assign n275 = ~x10 & ~x11 ;
  assign n276 = ~x12 & ~x13 ;
  assign n277 = n275 & n276 ;
  assign n278 = ~x6 & ~x7 ;
  assign n279 = ~x8 & ~x9 ;
  assign n280 = n278 & n279 ;
  assign n281 = n277 & n280 ;
  assign n282 = n274 & n281 ;
  assign n283 = n267 & n282 ;
  assign n226 = ~n71 & ~n177 ;
  assign n227 = ~n33 & ~n49 ;
  assign n228 = n226 & n227 ;
  assign n229 = ~n64 & ~n85 ;
  assign n230 = ~n67 & ~n68 ;
  assign n231 = n229 & n230 ;
  assign n232 = n228 & n231 ;
  assign n233 = ~n50 & ~n93 ;
  assign n234 = ~n42 & n233 ;
  assign n235 = ~n34 & ~n36 ;
  assign n236 = n120 & n235 ;
  assign n237 = n234 & n236 ;
  assign n238 = n232 & n237 ;
  assign n239 = ~n141 & ~n173 ;
  assign n240 = n118 & n239 ;
  assign n242 = ~n65 & ~n78 ;
  assign n243 = n241 & n242 ;
  assign n244 = n240 & n243 ;
  assign n245 = ~n134 & ~n136 ;
  assign n246 = ~n185 & ~n187 ;
  assign n247 = n245 & n246 ;
  assign n248 = ~n170 & ~n171 ;
  assign n249 = n160 & n248 ;
  assign n250 = n247 & n249 ;
  assign n251 = n244 & n250 ;
  assign n252 = n238 & n251 ;
  assign n284 = n283 ^ n252 ;
  assign n345 = n344 ^ n284 ;
  assign n414 = n413 ^ n345 ;
  assign n464 = n463 ^ n414 ;
  assign n526 = n525 ^ n464 ;
  assign n551 = n550 ^ n526 ;
  assign n552 = n225 & n551 ;
  assign n553 = n552 ^ n225 ;
  assign n554 = n553 ^ n551 ;
  assign n569 = ~n463 & n525 ;
  assign n568 = n414 & n525 ;
  assign n570 = n569 ^ n568 ;
  assign n566 = ~n414 & n463 ;
  assign n561 = ~n252 & n283 ;
  assign n562 = n344 & n561 ;
  assign n560 = ~n344 & ~n413 ;
  assign n563 = n562 ^ n560 ;
  assign n558 = n252 & ~n283 ;
  assign n559 = ~n344 & n558 ;
  assign n564 = n563 ^ n559 ;
  assign n556 = ~n252 & n413 ;
  assign n555 = ~n283 & ~n413 ;
  assign n557 = n556 ^ n555 ;
  assign n565 = n564 ^ n557 ;
  assign n567 = n566 ^ n565 ;
  assign n571 = n570 ^ n567 ;
  assign n572 = ~n554 & n571 ;
  assign n573 = n572 ^ n554 ;
  assign n575 = n439 & n460 ;
  assign n576 = n457 & n458 ;
  assign n579 = n345 & n576 ;
  assign n580 = n575 & n579 ;
  assign n577 = n413 & n576 ;
  assign n578 = n575 & n577 ;
  assign n581 = n580 ^ n578 ;
  assign n582 = n581 ^ n413 ;
  assign n574 = n565 ^ n345 ;
  assign n583 = n582 ^ n574 ;
  assign n588 = n464 & n583 ;
  assign n589 = n588 ^ n583 ;
  assign n590 = n550 & n589 ;
  assign n591 = n590 ^ n589 ;
  assign n584 = n525 & n583 ;
  assign n585 = n584 ^ n583 ;
  assign n586 = n550 & n585 ;
  assign n587 = n586 ^ n585 ;
  assign n592 = n591 ^ n587 ;
  assign n596 = n252 & n344 ;
  assign n595 = n283 & ~n344 ;
  assign n597 = n596 ^ n595 ;
  assign n598 = n597 ^ n561 ;
  assign n604 = n592 & n598 ;
  assign n605 = n604 ^ n598 ;
  assign n593 = n414 & n463 ;
  assign n594 = n593 ^ n414 ;
  assign n599 = n565 & ~n598 ;
  assign n600 = n594 & n599 ;
  assign n601 = n600 ^ n599 ;
  assign n602 = n592 & n601 ;
  assign n603 = n602 ^ n601 ;
  assign n606 = n605 ^ n603 ;
  assign n607 = ~n573 & n606 ;
  assign n608 = n607 ^ n573 ;
  assign n609 = n565 ^ n464 ;
  assign n610 = ~n565 & ~n609 ;
  assign n611 = n610 ^ n464 ;
  assign n612 = n611 ^ n525 ;
  assign n613 = n525 & n612 ;
  assign n614 = n613 ^ n610 ;
  assign n615 = n614 ^ n464 ;
  assign n634 = n615 ^ n601 ;
  assign n635 = n634 ^ n598 ;
  assign n624 = n464 & n525 ;
  assign n625 = n624 ^ n525 ;
  assign n626 = n625 ^ n464 ;
  assign n627 = n583 ^ n565 ;
  assign n628 = ~n626 & n627 ;
  assign n629 = n628 ^ n583 ;
  assign n630 = n629 ^ n626 ;
  assign n631 = ~n554 & ~n630 ;
  assign n632 = n631 ^ n592 ;
  assign n616 = n615 ^ n592 ;
  assign n617 = n601 ^ n598 ;
  assign n618 = ~n615 & n617 ;
  assign n619 = n618 ^ n592 ;
  assign n620 = n619 ^ n615 ;
  assign n621 = n620 ^ n617 ;
  assign n622 = ~n616 & ~n621 ;
  assign n623 = n622 ^ n618 ;
  assign n633 = n632 ^ n623 ;
  assign n636 = n635 ^ n633 ;
  assign n637 = n526 & ~n550 ;
  assign n638 = n554 & ~n637 ;
  assign n639 = n638 ^ n571 ;
  assign n640 = n551 ^ n225 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = 1'b0 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = ~n608 ;
  assign y29 = n636 ;
  assign y30 = n639 ;
  assign y31 = n640 ;
endmodule
