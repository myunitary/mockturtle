module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 ;
  assign n33 = ~x12 & ~x13 ;
  assign n34 = ~x14 & ~x15 ;
  assign n35 = n33 & n34 ;
  assign n36 = ~x8 & ~x9 ;
  assign n37 = ~x10 & ~x11 ;
  assign n38 = n36 & n37 ;
  assign n39 = n35 & n38 ;
  assign n40 = ~x4 & ~x5 ;
  assign n41 = ~x6 & ~x7 ;
  assign n42 = n40 & n41 ;
  assign n43 = ~x0 & ~x1 ;
  assign n44 = ~x2 & ~x3 ;
  assign n45 = n43 & n44 ;
  assign n46 = n42 & n45 ;
  assign n47 = ~n39 & ~n46 ;
  assign n48 = ~x28 & ~x29 ;
  assign n49 = ~x30 & ~x31 ;
  assign n50 = n48 & n49 ;
  assign n51 = ~x24 & ~x25 ;
  assign n52 = ~x26 & ~x27 ;
  assign n53 = n51 & n52 ;
  assign n54 = n50 & n53 ;
  assign n55 = ~x20 & ~x21 ;
  assign n56 = ~x22 & ~x23 ;
  assign n57 = n55 & n56 ;
  assign n58 = ~x16 & ~x17 ;
  assign n59 = ~x18 & ~x19 ;
  assign n60 = n58 & n59 ;
  assign n61 = n57 & n60 ;
  assign n62 = ~n54 & ~n61 ;
  assign n63 = n47 & n62 ;
  assign n64 = n54 & ~n61 ;
  assign n65 = n64 ^ n61 ;
  assign n66 = n47 & n65 ;
  assign n67 = n47 & ~n64 ;
  assign n68 = n67 ^ n46 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = 1'b0 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = n63 ;
  assign y30 = n66 ;
  assign y31 = ~n68 ;
endmodule
