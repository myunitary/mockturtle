module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 ;
  assign n49 = x4 & x5 ;
  assign n50 = n49 ^ x5 ;
  assign n51 = x8 & n50 ;
  assign n54 = n51 ^ x5 ;
  assign n33 = x2 & x7 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n34 ^ x7 ;
  assign n36 = x1 & x5 ;
  assign n37 = ~n35 & n36 ;
  assign n16 = ~x4 & x7 ;
  assign n38 = x3 & ~n16 ;
  assign n39 = ~n37 & n38 ;
  assign n40 = n39 ^ x3 ;
  assign n19 = x3 & x4 ;
  assign n31 = n19 ^ x4 ;
  assign n32 = x7 & n31 ;
  assign n41 = n40 ^ n32 ;
  assign n42 = n32 ^ x8 ;
  assign n43 = x8 & ~n42 ;
  assign n44 = n43 ^ x8 ;
  assign n45 = n44 ^ n40 ;
  assign n46 = n41 & ~n45 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = n47 ^ n40 ;
  assign n71 = n54 ^ n48 ;
  assign n58 = x1 & x4 ;
  assign n59 = ~x4 & x8 ;
  assign n60 = ~n58 & ~n59 ;
  assign n61 = x0 & ~n60 ;
  assign n62 = ~x0 & ~n58 ;
  assign n63 = ~x6 & ~x7 ;
  assign n64 = ~n62 & n63 ;
  assign n65 = ~n61 & n64 ;
  assign n20 = x4 & x8 ;
  assign n55 = n51 ^ n20 ;
  assign n56 = n54 & n55 ;
  assign n57 = n56 ^ n20 ;
  assign n66 = n65 ^ n57 ;
  assign n72 = n71 ^ n66 ;
  assign n73 = n65 ^ x5 ;
  assign n74 = n73 ^ n57 ;
  assign n75 = ~n72 & ~n74 ;
  assign n67 = n57 ^ x5 ;
  assign n52 = n51 ^ n48 ;
  assign n68 = n67 ^ n52 ;
  assign n69 = n66 & n68 ;
  assign n76 = n75 ^ n69 ;
  assign n77 = n76 ^ n57 ;
  assign n78 = n77 ^ n71 ;
  assign n79 = n69 ^ n65 ;
  assign n80 = n79 ^ n48 ;
  assign n81 = n78 & n80 ;
  assign n82 = n81 ^ n75 ;
  assign n70 = n69 ^ n56 ;
  assign n83 = n82 ^ n70 ;
  assign n30 = n20 ^ x5 ;
  assign n53 = n52 ^ n30 ;
  assign n84 = n83 ^ n53 ;
  assign n85 = x9 & n84 ;
  assign n86 = n85 ^ x9 ;
  assign n87 = n86 ^ n84 ;
  assign n12 = x5 & x6 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = x9 & n13 ;
  assign n15 = n12 ^ x5 ;
  assign n17 = x1 & ~x2 ;
  assign n18 = ~n16 & n17 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = n18 & n21 ;
  assign n23 = ~x7 & ~x8 ;
  assign n24 = ~x1 & x2 ;
  assign n25 = n23 & n24 ;
  assign n26 = ~x9 & ~n25 ;
  assign n27 = ~n22 & n26 ;
  assign n28 = n15 & ~n27 ;
  assign n29 = ~n14 & ~n28 ;
  assign n88 = n87 ^ n29 ;
  assign n89 = n29 ^ x10 ;
  assign n90 = x10 & n89 ;
  assign n91 = n90 ^ x10 ;
  assign n92 = n91 ^ n87 ;
  assign n93 = n88 & n92 ;
  assign n94 = n93 ^ n90 ;
  assign n95 = n94 ^ n87 ;
  assign n96 = ~x6 & x7 ;
  assign n97 = x10 & n96 ;
  assign n98 = x3 ^ x2 ;
  assign n99 = x8 & x9 ;
  assign n100 = n99 ^ x8 ;
  assign n101 = n100 ^ x9 ;
  assign n102 = n98 & ~n101 ;
  assign n103 = ~x10 & ~n102 ;
  assign n104 = ~x7 & ~n103 ;
  assign n105 = x8 & x10 ;
  assign n106 = x9 & n105 ;
  assign n107 = ~n104 & ~n106 ;
  assign n108 = x6 & ~n107 ;
  assign n109 = ~n97 & ~n108 ;
  assign n110 = ~n95 & n109 ;
  assign n111 = n110 ^ n109 ;
  assign n116 = x1 & x2 ;
  assign n117 = x0 & ~n116 ;
  assign n118 = ~x0 & x2 ;
  assign n119 = x4 & ~x7 ;
  assign n120 = ~n118 & n119 ;
  assign n121 = ~n117 & n120 ;
  assign n122 = x4 & x9 ;
  assign n123 = n122 ^ x4 ;
  assign n124 = n123 ^ x9 ;
  assign n125 = n35 & ~n124 ;
  assign n126 = n125 ^ n35 ;
  assign n127 = x8 & ~x9 ;
  assign n128 = ~x1 & ~n127 ;
  assign n129 = ~n126 & n128 ;
  assign n130 = n129 ^ n127 ;
  assign n131 = n121 & ~n130 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = x6 & ~n132 ;
  assign n134 = n133 ^ x6 ;
  assign n135 = n134 ^ n132 ;
  assign n112 = ~x7 & x9 ;
  assign n113 = x7 & ~n101 ;
  assign n114 = ~n19 & n113 ;
  assign n115 = ~n112 & ~n114 ;
  assign n136 = n135 ^ n115 ;
  assign n137 = n115 ^ x5 ;
  assign n138 = x5 & n137 ;
  assign n139 = n138 ^ x5 ;
  assign n140 = n139 ^ n135 ;
  assign n141 = ~n136 & ~n140 ;
  assign n142 = n141 ^ n138 ;
  assign n143 = n142 ^ n135 ;
  assign n144 = x4 & x6 ;
  assign n145 = n144 ^ x4 ;
  assign n146 = n145 ^ x6 ;
  assign n147 = x7 & n116 ;
  assign n148 = n147 ^ n116 ;
  assign n149 = ~n146 & n148 ;
  assign n150 = n147 ^ x7 ;
  assign n151 = n150 ^ n116 ;
  assign n152 = x4 & ~n101 ;
  assign n153 = ~n151 & n152 ;
  assign n154 = n153 ^ n152 ;
  assign n155 = n149 & n154 ;
  assign n156 = n155 ^ n149 ;
  assign n157 = n156 ^ n154 ;
  assign n158 = n157 ^ x3 ;
  assign n159 = x6 & n101 ;
  assign n160 = ~n112 & n124 ;
  assign n161 = n159 & n160 ;
  assign n162 = n161 ^ x3 ;
  assign n163 = n161 & n162 ;
  assign n164 = n163 ^ n161 ;
  assign n165 = n164 ^ n157 ;
  assign n166 = n158 & n165 ;
  assign n167 = n166 ^ n163 ;
  assign n168 = n167 ^ n157 ;
  assign n169 = n168 ^ x5 ;
  assign n170 = ~x9 & n59 ;
  assign n171 = ~n112 & ~n170 ;
  assign n172 = ~x6 & ~n171 ;
  assign n173 = n172 ^ x5 ;
  assign n174 = n172 & n173 ;
  assign n175 = n174 ^ n172 ;
  assign n176 = n175 ^ n168 ;
  assign n177 = n169 & n176 ;
  assign n178 = n177 ^ n174 ;
  assign n179 = n178 ^ n168 ;
  assign n180 = n143 & ~n179 ;
  assign n181 = n180 ^ n179 ;
  assign n182 = x10 & ~n181 ;
  assign n183 = n182 ^ x10 ;
  assign n184 = n183 ^ n181 ;
  assign n186 = x6 & x7 ;
  assign n189 = ~x8 & ~n186 ;
  assign n192 = n189 ^ x10 ;
  assign n187 = ~x9 & n186 ;
  assign n188 = n105 & n187 ;
  assign n228 = n192 ^ n188 ;
  assign n196 = x6 & x9 ;
  assign n197 = n196 ^ x6 ;
  assign n198 = x4 & n197 ;
  assign n199 = n198 ^ n197 ;
  assign n200 = x1 & n15 ;
  assign n201 = n200 ^ n15 ;
  assign n202 = ~n199 & ~n201 ;
  assign n203 = ~x3 & ~n202 ;
  assign n205 = x6 ^ x3 ;
  assign n206 = n205 ^ x5 ;
  assign n204 = x5 ^ x3 ;
  assign n207 = n206 ^ n204 ;
  assign n209 = ~x4 & ~x9 ;
  assign n208 = x5 & n206 ;
  assign n210 = n209 ^ n208 ;
  assign n211 = n207 & n210 ;
  assign n212 = n211 ^ n208 ;
  assign n213 = x2 & ~n212 ;
  assign n214 = n213 ^ x2 ;
  assign n215 = n214 ^ n212 ;
  assign n216 = x2 & n19 ;
  assign n217 = n197 & n216 ;
  assign n218 = n215 & n217 ;
  assign n219 = n218 ^ n215 ;
  assign n220 = n219 ^ n217 ;
  assign n221 = n203 & ~n220 ;
  assign n222 = n221 ^ n220 ;
  assign n193 = n189 ^ x7 ;
  assign n194 = ~n192 & ~n193 ;
  assign n195 = n194 ^ x7 ;
  assign n223 = n222 ^ n195 ;
  assign n229 = n228 ^ n223 ;
  assign n230 = n222 ^ x10 ;
  assign n231 = n230 ^ n195 ;
  assign n232 = ~n229 & n231 ;
  assign n224 = n195 ^ x10 ;
  assign n190 = n189 ^ n188 ;
  assign n225 = n224 ^ n190 ;
  assign n226 = ~n223 & ~n225 ;
  assign n233 = n232 ^ n226 ;
  assign n234 = n233 ^ n195 ;
  assign n235 = n234 ^ n228 ;
  assign n236 = n226 ^ n222 ;
  assign n237 = n236 ^ n188 ;
  assign n238 = ~n235 & ~n237 ;
  assign n239 = n238 ^ n232 ;
  assign n227 = n226 ^ n194 ;
  assign n240 = n239 ^ n227 ;
  assign n185 = x10 ^ x7 ;
  assign n191 = n190 ^ n185 ;
  assign n241 = n240 ^ n191 ;
  assign n242 = n241 ^ n188 ;
  assign n243 = n184 & n242 ;
  assign n244 = n243 ^ n242 ;
  assign n245 = x6 & ~x7 ;
  assign n246 = n49 & n245 ;
  assign n247 = ~n96 & ~n246 ;
  assign n248 = x8 & ~n247 ;
  assign n363 = n248 ^ x9 ;
  assign n249 = x5 & ~x8 ;
  assign n250 = x9 & n249 ;
  assign n251 = ~n105 & ~n250 ;
  assign n252 = n186 & ~n251 ;
  assign n253 = x5 & x7 ;
  assign n254 = x8 & ~n253 ;
  assign n255 = ~x10 & ~n254 ;
  assign n256 = x9 & ~n255 ;
  assign n257 = ~n252 & ~n256 ;
  assign n342 = n257 ^ x10 ;
  assign n364 = n363 ^ n342 ;
  assign n258 = n257 ^ n248 ;
  assign n348 = n258 ^ x10 ;
  assign n287 = x0 & x6 ;
  assign n288 = n287 ^ x0 ;
  assign n289 = n288 ^ x4 ;
  assign n290 = n289 ^ x5 ;
  assign n291 = x4 & n290 ;
  assign n292 = n291 ^ n290 ;
  assign n293 = n292 ^ x4 ;
  assign n294 = n293 ^ n289 ;
  assign n295 = x4 ^ x3 ;
  assign n296 = x1 & n295 ;
  assign n297 = ~n294 & n296 ;
  assign n298 = n297 ^ n296 ;
  assign n299 = x0 & x1 ;
  assign n300 = n19 & n299 ;
  assign n301 = n300 ^ n19 ;
  assign n302 = x5 & ~n146 ;
  assign n303 = n302 ^ x5 ;
  assign n304 = n303 ^ n146 ;
  assign n305 = n301 & n304 ;
  assign n306 = n305 ^ n304 ;
  assign n307 = n306 ^ x5 ;
  assign n308 = n298 & n307 ;
  assign n309 = n308 ^ n298 ;
  assign n310 = n309 ^ n298 ;
  assign n311 = n310 ^ n307 ;
  assign n312 = x2 & n311 ;
  assign n313 = n312 ^ x2 ;
  assign n262 = x6 ^ x5 ;
  assign n277 = n262 ^ x2 ;
  assign n276 = n262 ^ x6 ;
  assign n278 = n277 ^ n276 ;
  assign n279 = n276 ^ n262 ;
  assign n280 = ~n278 & ~n279 ;
  assign n281 = n280 ^ n276 ;
  assign n282 = x3 & n281 ;
  assign n283 = n282 ^ n262 ;
  assign n284 = n283 ^ x6 ;
  assign n285 = x4 & ~n284 ;
  assign n286 = n285 ^ x4 ;
  assign n314 = n313 ^ n286 ;
  assign n315 = x4 & x7 ;
  assign n316 = n284 & n315 ;
  assign n317 = n316 ^ x7 ;
  assign n318 = n317 ^ n313 ;
  assign n319 = n314 & n318 ;
  assign n320 = n319 ^ n314 ;
  assign n321 = n320 ^ n316 ;
  assign n322 = n321 ^ n313 ;
  assign n265 = x6 ^ x2 ;
  assign n263 = x2 ^ x1 ;
  assign n264 = n263 ^ x2 ;
  assign n266 = n265 ^ n264 ;
  assign n267 = n265 ^ x2 ;
  assign n268 = n266 & ~n267 ;
  assign n269 = n268 ^ n265 ;
  assign n270 = n262 & ~n269 ;
  assign n271 = n270 ^ n12 ;
  assign n272 = n19 & ~n271 ;
  assign n273 = n272 ^ n19 ;
  assign n274 = n273 ^ n271 ;
  assign n275 = n274 ^ n270 ;
  assign n323 = n322 ^ n275 ;
  assign n324 = n275 ^ x8 ;
  assign n325 = x8 & ~n324 ;
  assign n326 = n325 ^ x8 ;
  assign n327 = n326 ^ n322 ;
  assign n328 = ~n323 & n327 ;
  assign n329 = n328 ^ n323 ;
  assign n330 = n329 ^ n327 ;
  assign n331 = n330 ^ n325 ;
  assign n332 = n331 ^ n322 ;
  assign n333 = ~n49 & n186 ;
  assign n334 = x3 & n96 ;
  assign n335 = ~x2 & n245 ;
  assign n336 = ~n334 & ~n335 ;
  assign n337 = n49 & ~n336 ;
  assign n338 = ~n333 & ~n337 ;
  assign n339 = n332 & n338 ;
  assign n340 = n339 ^ n338 ;
  assign n259 = n257 ^ x9 ;
  assign n260 = ~n258 & ~n259 ;
  assign n261 = n260 ^ x9 ;
  assign n341 = n340 ^ n261 ;
  assign n349 = n348 ^ n341 ;
  assign n350 = n340 ^ n248 ;
  assign n351 = n350 ^ n261 ;
  assign n352 = n349 & n351 ;
  assign n353 = n352 ^ n349 ;
  assign n343 = n261 ^ n248 ;
  assign n344 = n343 ^ n342 ;
  assign n345 = n341 & n344 ;
  assign n346 = n345 ^ n341 ;
  assign n354 = n353 ^ n346 ;
  assign n355 = n354 ^ n261 ;
  assign n356 = n355 ^ n348 ;
  assign n357 = n346 ^ n340 ;
  assign n358 = n357 ^ x10 ;
  assign n359 = n356 & n358 ;
  assign n360 = n359 ^ n358 ;
  assign n361 = n360 ^ n353 ;
  assign n347 = n346 ^ n260 ;
  assign n362 = n361 ^ n347 ;
  assign n365 = n364 ^ n362 ;
  assign n366 = n365 ^ n257 ;
  assign n367 = x7 & n12 ;
  assign n368 = ~x2 & n20 ;
  assign n369 = n367 & n368 ;
  assign n370 = ~x5 & ~x6 ;
  assign n371 = ~x4 & ~x7 ;
  assign n372 = ~x8 & n371 ;
  assign n373 = n370 & n372 ;
  assign n374 = ~n369 & ~n373 ;
  assign n375 = ~x9 & ~x10 ;
  assign n376 = ~x3 & n375 ;
  assign n377 = ~n374 & n376 ;
  assign n390 = n148 ^ n12 ;
  assign n391 = n12 ^ x3 ;
  assign n392 = ~x3 & n391 ;
  assign n393 = n392 ^ x3 ;
  assign n394 = n393 ^ n148 ;
  assign n395 = n390 & n394 ;
  assign n396 = n395 ^ n392 ;
  assign n397 = n396 ^ n148 ;
  assign n398 = ~x5 & ~x7 ;
  assign n399 = n397 & n398 ;
  assign n400 = n399 ^ n397 ;
  assign n401 = n400 ^ n398 ;
  assign n402 = x4 & ~n245 ;
  assign n403 = n401 & n402 ;
  assign n404 = n403 ^ n245 ;
  assign n386 = x2 & x3 ;
  assign n387 = n299 & n370 ;
  assign n388 = ~n246 & ~n387 ;
  assign n389 = n386 & ~n388 ;
  assign n405 = n404 ^ n389 ;
  assign n406 = n389 ^ x8 ;
  assign n407 = x8 & ~n406 ;
  assign n408 = n407 ^ x8 ;
  assign n409 = n408 ^ n404 ;
  assign n410 = ~n405 & n409 ;
  assign n411 = n410 ^ n407 ;
  assign n412 = n411 ^ n404 ;
  assign n378 = x8 & n367 ;
  assign n379 = x9 & ~n378 ;
  assign n380 = x2 & ~x3 ;
  assign n381 = x3 & x8 ;
  assign n382 = ~n380 & ~n381 ;
  assign n383 = n49 & n187 ;
  assign n384 = ~n382 & n383 ;
  assign n385 = ~n379 & ~n384 ;
  assign n413 = n412 ^ n385 ;
  assign n414 = n385 ^ x10 ;
  assign n415 = x10 & n414 ;
  assign n416 = n415 ^ x10 ;
  assign n417 = n416 ^ n412 ;
  assign n418 = n413 & n417 ;
  assign n419 = n418 ^ n415 ;
  assign n420 = n419 ^ n412 ;
  assign n421 = x3 & ~x8 ;
  assign n422 = n299 & n421 ;
  assign n423 = n398 & n422 ;
  assign n424 = ~n378 & ~n423 ;
  assign n425 = x2 & ~n424 ;
  assign n426 = n367 & n381 ;
  assign n427 = ~n425 & ~n426 ;
  assign n428 = x4 & ~n427 ;
  assign n429 = n12 & n216 ;
  assign n430 = n23 & ~n370 ;
  assign n431 = ~n429 & n430 ;
  assign n432 = n375 & ~n431 ;
  assign n433 = ~n428 & n432 ;
  assign n434 = n23 & n375 ;
  assign n435 = ~n429 & n434 ;
  assign y0 = ~n111 ;
  assign y1 = n244 ;
  assign y2 = n366 ;
  assign y3 = ~n377 ;
  assign y4 = n420 ;
  assign y5 = ~n433 ;
  assign y6 = ~n435 ;
endmodule
