module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 ;
  assign n8 = x2 ^ x1 ;
  assign n9 = n8 ^ x4 ;
  assign n12 = n9 ^ x4 ;
  assign n10 = n9 ^ x2 ;
  assign n13 = n12 ^ n10 ;
  assign n14 = n12 ^ x0 ;
  assign n15 = x4 ^ x3 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = ~n14 & n16 ;
  assign n18 = n17 ^ x0 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = ~n13 & ~n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ x0 ;
  assign n11 = n10 ^ n9 ;
  assign n23 = n22 ^ n11 ;
  assign n24 = n12 ^ n9 ;
  assign n26 = n10 ^ x0 ;
  assign n25 = n15 ^ n12 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = ~n24 & n27 ;
  assign n29 = n28 ^ n20 ;
  assign n30 = n29 ^ n17 ;
  assign n31 = n23 & n30 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = n32 ^ x2 ;
  assign n34 = n33 ^ x3 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = n35 ^ n8 ;
  assign n38 = x3 ^ x1 ;
  assign n41 = n38 ^ x3 ;
  assign n37 = x4 ^ x2 ;
  assign n50 = n41 ^ n37 ;
  assign n42 = n38 ^ x4 ;
  assign n43 = n41 & n42 ;
  assign n44 = n43 ^ x4 ;
  assign n45 = n44 ^ x0 ;
  assign n51 = n50 ^ n45 ;
  assign n52 = x3 ^ x0 ;
  assign n53 = n52 ^ n44 ;
  assign n54 = ~n51 & ~n53 ;
  assign n46 = n44 ^ x3 ;
  assign n39 = n38 ^ n37 ;
  assign n47 = n46 ^ n39 ;
  assign n48 = ~n45 & n47 ;
  assign n55 = n54 ^ n48 ;
  assign n56 = n55 ^ n44 ;
  assign n57 = n56 ^ n50 ;
  assign n58 = n48 ^ x0 ;
  assign n59 = n58 ^ n37 ;
  assign n60 = n57 & ~n59 ;
  assign n61 = n60 ^ n54 ;
  assign n49 = n48 ^ n43 ;
  assign n62 = n61 ^ n49 ;
  assign n40 = n39 ^ n15 ;
  assign n63 = n62 ^ n40 ;
  assign n64 = n63 ^ n37 ;
  assign n65 = n64 ^ n37 ;
  assign n66 = ~x2 & ~n42 ;
  assign n67 = n52 ^ x3 ;
  assign n68 = n67 ^ n15 ;
  assign n69 = n15 ^ x3 ;
  assign n70 = ~n68 & n69 ;
  assign n71 = n70 ^ n15 ;
  assign n72 = n66 & n71 ;
  assign n73 = x3 & x4 ;
  assign n74 = x0 & n73 ;
  assign n75 = x1 & x2 ;
  assign n76 = n75 ^ x1 ;
  assign n77 = n76 ^ x2 ;
  assign n78 = n77 ^ x4 ;
  assign n79 = x3 & ~n78 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n74 & n81 ;
  assign n83 = n82 ^ n81 ;
  assign n89 = x5 ^ x0 ;
  assign n90 = n89 ^ x4 ;
  assign n91 = n90 ^ x5 ;
  assign n92 = n91 ^ x4 ;
  assign n95 = n92 ^ n91 ;
  assign n93 = n92 ^ x5 ;
  assign n96 = n95 ^ n93 ;
  assign n97 = n95 ^ x6 ;
  assign n98 = n96 ^ x3 ;
  assign n99 = n97 & n98 ;
  assign n100 = n99 ^ n97 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = n101 ^ x6 ;
  assign n103 = n102 ^ n96 ;
  assign n104 = n96 & n103 ;
  assign n105 = n104 ^ n96 ;
  assign n106 = n105 ^ n103 ;
  assign n107 = n106 ^ n101 ;
  assign n108 = n107 ^ x6 ;
  assign n94 = n93 ^ n92 ;
  assign n109 = n108 ^ n94 ;
  assign n110 = n95 ^ n92 ;
  assign n112 = n93 ^ x6 ;
  assign n111 = n95 ^ x3 ;
  assign n113 = n112 ^ n111 ;
  assign n114 = n110 & n113 ;
  assign n115 = n114 ^ n106 ;
  assign n116 = n115 ^ n101 ;
  assign n117 = n109 & n116 ;
  assign n118 = n117 ^ x3 ;
  assign n119 = n118 ^ x3 ;
  assign n120 = x1 & ~x2 ;
  assign n121 = n119 & n120 ;
  assign n122 = n121 ^ x2 ;
  assign n84 = ~x0 & x2 ;
  assign n85 = n73 ^ x4 ;
  assign n86 = x2 & n85 ;
  assign n87 = n86 ^ x2 ;
  assign n88 = ~n84 & ~n87 ;
  assign n123 = n122 ^ n88 ;
  assign n124 = x4 & x6 ;
  assign n125 = n124 ^ x4 ;
  assign n126 = ~x2 & x3 ;
  assign n127 = ~n125 & n126 ;
  assign n128 = n127 ^ x2 ;
  assign n129 = n75 & ~n85 ;
  assign n130 = n129 ^ x1 ;
  assign n131 = ~n128 & n130 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = x0 & x1 ;
  assign n134 = n73 & n133 ;
  assign n135 = n134 ^ n73 ;
  assign n136 = n135 ^ x2 ;
  assign n137 = n15 & n37 ;
  assign n138 = n137 ^ n15 ;
  assign n139 = n138 ^ x4 ;
  assign n140 = n139 ^ x2 ;
  assign n141 = ~n139 & n140 ;
  assign n142 = n141 ^ n139 ;
  assign n143 = n142 ^ n135 ;
  assign n144 = ~n136 & ~n143 ;
  assign n145 = n144 ^ n141 ;
  assign n146 = n145 ^ n135 ;
  assign n147 = x4 ^ x1 ;
  assign n149 = n147 ^ n37 ;
  assign n148 = n147 ^ x0 ;
  assign n150 = n149 ^ n148 ;
  assign n152 = n150 ^ x4 ;
  assign n151 = n150 ^ n149 ;
  assign n153 = n152 ^ n151 ;
  assign n158 = n153 ^ n152 ;
  assign n155 = n150 ^ n147 ;
  assign n156 = n155 ^ n152 ;
  assign n157 = n156 ^ n15 ;
  assign n159 = n158 ^ n157 ;
  assign n160 = n156 ^ n153 ;
  assign n161 = n156 ^ n150 ;
  assign n162 = ~n160 & ~n161 ;
  assign n163 = n162 ^ n152 ;
  assign n164 = n163 ^ n161 ;
  assign n165 = n159 & ~n164 ;
  assign n166 = n165 ^ n162 ;
  assign n154 = n153 ^ n150 ;
  assign n167 = n166 ^ n154 ;
  assign n168 = n152 ^ n150 ;
  assign n169 = n168 ^ n153 ;
  assign n170 = n169 ^ n157 ;
  assign n171 = ~n15 & ~n170 ;
  assign n172 = n171 ^ n165 ;
  assign n173 = n172 ^ n152 ;
  assign n174 = n173 ^ n160 ;
  assign n175 = n167 & ~n174 ;
  assign n176 = n175 ^ n165 ;
  assign n177 = n176 ^ n152 ;
  assign n178 = n177 ^ n160 ;
  assign n179 = n178 ^ n15 ;
  assign n180 = n15 ^ x2 ;
  assign n184 = n180 ^ n15 ;
  assign n193 = n184 ^ x1 ;
  assign n185 = n180 ^ x4 ;
  assign n186 = n184 & n185 ;
  assign n187 = n186 ^ x4 ;
  assign n188 = n187 ^ x0 ;
  assign n194 = n193 ^ n188 ;
  assign n195 = n15 ^ x0 ;
  assign n196 = n195 ^ n187 ;
  assign n197 = ~n194 & ~n196 ;
  assign n189 = n187 ^ n15 ;
  assign n181 = n180 ^ x1 ;
  assign n190 = n189 ^ n181 ;
  assign n191 = ~n188 & n190 ;
  assign n198 = n197 ^ n191 ;
  assign n199 = n198 ^ n187 ;
  assign n200 = n199 ^ n193 ;
  assign n201 = n191 ^ x0 ;
  assign n202 = n201 ^ x1 ;
  assign n203 = n200 & ~n202 ;
  assign n204 = n203 ^ n197 ;
  assign n192 = n191 ^ n186 ;
  assign n205 = n204 ^ n192 ;
  assign n182 = n15 ^ x4 ;
  assign n183 = n182 ^ n181 ;
  assign n206 = n205 ^ n183 ;
  assign n207 = n206 ^ x1 ;
  assign n208 = n207 ^ x1 ;
  assign n209 = n147 ^ n15 ;
  assign n212 = n209 ^ n15 ;
  assign n221 = n212 ^ n37 ;
  assign n213 = n209 ^ x4 ;
  assign n214 = n212 & n213 ;
  assign n215 = n214 ^ x4 ;
  assign n216 = n215 ^ x0 ;
  assign n222 = n221 ^ n216 ;
  assign n223 = n215 ^ n195 ;
  assign n224 = ~n222 & ~n223 ;
  assign n217 = n215 ^ n15 ;
  assign n210 = n209 ^ n37 ;
  assign n218 = n217 ^ n210 ;
  assign n219 = ~n216 & n218 ;
  assign n225 = n224 ^ n219 ;
  assign n226 = n225 ^ n215 ;
  assign n227 = n226 ^ n221 ;
  assign n228 = n219 ^ x0 ;
  assign n229 = n228 ^ n37 ;
  assign n230 = n227 & ~n229 ;
  assign n231 = n230 ^ n224 ;
  assign n220 = n219 ^ n214 ;
  assign n232 = n231 ^ n220 ;
  assign n211 = n210 ^ n182 ;
  assign n233 = n232 ^ n211 ;
  assign n234 = n233 ^ n37 ;
  assign n235 = n234 ^ n37 ;
  assign n240 = x3 ^ x2 ;
  assign n243 = n240 ^ n182 ;
  assign n244 = ~n182 & n243 ;
  assign n255 = n244 ^ n240 ;
  assign n236 = ~x1 & x4 ;
  assign n256 = n244 ^ n236 ;
  assign n237 = n236 ^ n15 ;
  assign n238 = n237 ^ n236 ;
  assign n257 = n256 ^ n238 ;
  assign n258 = ~n255 & ~n257 ;
  assign n242 = n133 ^ x1 ;
  assign n245 = n244 ^ n242 ;
  assign n246 = n245 ^ n238 ;
  assign n247 = n246 ^ n243 ;
  assign n248 = n244 ^ n238 ;
  assign n249 = n248 ^ n240 ;
  assign n250 = ~n247 & ~n249 ;
  assign n251 = n250 ^ n242 ;
  assign n252 = n251 ^ n243 ;
  assign n253 = n251 ^ n238 ;
  assign n254 = ~n252 & ~n253 ;
  assign n259 = n258 ^ n254 ;
  assign n260 = n259 ^ n251 ;
  assign n239 = n238 ^ n182 ;
  assign n241 = n240 ^ n239 ;
  assign n261 = n260 ^ n241 ;
  assign n262 = n261 ^ n236 ;
  assign n263 = n73 ^ x3 ;
  assign n264 = n263 ^ x4 ;
  assign n265 = ~x0 & ~n264 ;
  assign n266 = ~n77 & n265 ;
  assign n269 = ~x3 & x4 ;
  assign n270 = n133 ^ x0 ;
  assign n271 = n270 ^ x1 ;
  assign n272 = n269 & n271 ;
  assign n273 = n272 ^ x3 ;
  assign n267 = x1 & ~x3 ;
  assign n268 = ~x4 & ~n267 ;
  assign n274 = n273 ^ n268 ;
  assign n275 = x2 & ~n274 ;
  assign n276 = n275 ^ n274 ;
  assign n277 = n276 ^ n268 ;
  assign n278 = x2 & ~n264 ;
  assign n279 = x0 & n278 ;
  assign n280 = n84 & ~n264 ;
  assign n281 = x1 & n263 ;
  assign n282 = n281 ^ n263 ;
  assign n283 = n84 & n282 ;
  assign n284 = n263 & n270 ;
  assign n285 = x2 & n284 ;
  assign n286 = x2 & n263 ;
  assign n287 = n133 & n286 ;
  assign n288 = n242 & n286 ;
  assign n291 = x4 & x5 ;
  assign n292 = n291 ^ x4 ;
  assign n293 = x3 & n292 ;
  assign n294 = n293 ^ x3 ;
  assign n295 = n133 & n294 ;
  assign n296 = n285 ^ x2 ;
  assign n297 = n296 ^ n284 ;
  assign n298 = n295 & n297 ;
  assign n299 = n298 ^ n295 ;
  assign n300 = n299 ^ n297 ;
  assign n289 = x2 & n135 ;
  assign n290 = n289 ^ x2 ;
  assign n301 = n300 ^ n290 ;
  assign n302 = x0 & ~x2 ;
  assign n329 = x6 ^ x4 ;
  assign n310 = n147 ^ x3 ;
  assign n330 = n329 ^ n310 ;
  assign n303 = n147 ^ x4 ;
  assign n315 = n303 ^ x3 ;
  assign n304 = n147 ^ x6 ;
  assign n305 = n303 & n304 ;
  assign n306 = n305 ^ n304 ;
  assign n307 = n306 ^ x6 ;
  assign n308 = n307 ^ x5 ;
  assign n316 = n315 ^ n308 ;
  assign n317 = x5 ^ x4 ;
  assign n318 = n317 ^ n307 ;
  assign n319 = n316 & n318 ;
  assign n320 = n319 ^ n316 ;
  assign n309 = n307 ^ x4 ;
  assign n311 = n310 ^ n309 ;
  assign n312 = n308 & n311 ;
  assign n313 = n312 ^ n311 ;
  assign n321 = n320 ^ n313 ;
  assign n322 = n321 ^ n307 ;
  assign n323 = n322 ^ n315 ;
  assign n324 = n313 ^ x5 ;
  assign n325 = n324 ^ x3 ;
  assign n326 = n323 & n325 ;
  assign n327 = n326 ^ n320 ;
  assign n314 = n313 ^ n306 ;
  assign n328 = n327 ^ n314 ;
  assign n331 = n330 ^ n328 ;
  assign n332 = n331 ^ x3 ;
  assign n333 = n332 ^ x3 ;
  assign n334 = n302 & n333 ;
  assign n335 = n334 ^ n302 ;
  assign n336 = n335 ^ n302 ;
  assign n337 = x2 & n133 ;
  assign n338 = n337 ^ n133 ;
  assign n342 = x3 & n125 ;
  assign n343 = n342 ^ x3 ;
  assign n339 = x5 & x6 ;
  assign n340 = n339 ^ x6 ;
  assign n341 = n73 & n340 ;
  assign n344 = n343 ^ n341 ;
  assign n345 = n338 & n344 ;
  assign n346 = n345 ^ x2 ;
  assign n347 = n346 ^ n290 ;
  assign n348 = x1 ^ x0 ;
  assign n349 = ~x2 & n85 ;
  assign n350 = ~n348 & n349 ;
  assign n351 = ~x1 & n85 ;
  assign n352 = n302 & n351 ;
  assign y0 = ~n36 ;
  assign y1 = n65 ;
  assign y2 = n72 ;
  assign y3 = n83 ;
  assign y4 = ~n123 ;
  assign y5 = n132 ;
  assign y6 = ~n146 ;
  assign y7 = n179 ;
  assign y8 = n208 ;
  assign y9 = n235 ;
  assign y10 = n262 ;
  assign y11 = n266 ;
  assign y12 = n277 ;
  assign y13 = n279 ;
  assign y14 = n280 ;
  assign y15 = n283 ;
  assign y16 = n285 ;
  assign y17 = n287 ;
  assign y18 = n288 ;
  assign y19 = n278 ;
  assign y20 = n301 ;
  assign y21 = n336 ;
  assign y22 = n347 ;
  assign y23 = ~1'b0 ;
  assign y24 = n350 ;
  assign y25 = n352 ;
endmodule
