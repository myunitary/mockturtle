module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 ;
  assign n8 = x2 ^ x1 ;
  assign n9 = n8 ^ x4 ;
  assign n11 = n9 ^ x2 ;
  assign n22 = n11 ^ n9 ;
  assign n10 = n9 ^ x4 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n10 ^ x0 ;
  assign n14 = x4 ^ x3 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = ~n13 & n15 ;
  assign n17 = n16 ^ x0 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = ~n12 & ~n18 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n20 ^ x0 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n10 ^ n9 ;
  assign n26 = n14 ^ n10 ;
  assign n25 = n11 ^ x0 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = ~n24 & n27 ;
  assign n29 = n28 ^ n19 ;
  assign n30 = n29 ^ n16 ;
  assign n31 = n23 & n30 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = n32 ^ x2 ;
  assign n34 = n33 ^ x3 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = n35 ^ n8 ;
  assign n40 = x3 & x4 ;
  assign n45 = n40 ^ x3 ;
  assign n46 = n45 ^ x4 ;
  assign n47 = x1 & ~n46 ;
  assign n48 = x2 & n47 ;
  assign n41 = n40 ^ x4 ;
  assign n42 = x1 & n41 ;
  assign n37 = ~x0 & x3 ;
  assign n38 = ~x1 & x4 ;
  assign n39 = n37 & n38 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = ~x2 & n43 ;
  assign n49 = n48 ^ n44 ;
  assign n50 = x3 ^ x1 ;
  assign n51 = n50 ^ x4 ;
  assign n52 = ~x2 & ~n51 ;
  assign n53 = x3 ^ x0 ;
  assign n54 = n53 ^ x3 ;
  assign n55 = n54 ^ n14 ;
  assign n56 = n14 ^ x3 ;
  assign n57 = ~n55 & n56 ;
  assign n58 = n57 ^ n14 ;
  assign n59 = n52 & n58 ;
  assign n60 = x0 & n40 ;
  assign n61 = ~x1 & ~x2 ;
  assign n62 = x3 & ~n61 ;
  assign n63 = n46 & ~n62 ;
  assign n64 = ~n60 & n63 ;
  assign n98 = ~x0 & x2 ;
  assign n99 = x2 & ~n41 ;
  assign n100 = ~n98 & ~n99 ;
  assign n65 = x1 & ~x2 ;
  assign n66 = x5 ^ x0 ;
  assign n67 = n66 ^ x4 ;
  assign n68 = n67 ^ x5 ;
  assign n69 = n68 ^ x4 ;
  assign n71 = n69 ^ x5 ;
  assign n84 = n71 ^ n69 ;
  assign n70 = n69 ^ n68 ;
  assign n72 = n71 ^ n70 ;
  assign n73 = n70 ^ x6 ;
  assign n74 = n72 ^ x3 ;
  assign n75 = n73 & n74 ;
  assign n76 = n75 ^ n73 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = n77 ^ x6 ;
  assign n79 = n78 ^ n72 ;
  assign n80 = n72 & ~n79 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = n81 ^ n77 ;
  assign n83 = n82 ^ x6 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = n70 ^ n69 ;
  assign n88 = n70 ^ x3 ;
  assign n87 = n71 ^ x6 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = n86 & n89 ;
  assign n91 = n90 ^ n81 ;
  assign n92 = n91 ^ n77 ;
  assign n93 = n85 & n92 ;
  assign n94 = n93 ^ x3 ;
  assign n95 = n94 ^ x3 ;
  assign n96 = n65 & n95 ;
  assign n97 = n96 ^ x2 ;
  assign n101 = n100 ^ n97 ;
  assign n102 = x4 & x6 ;
  assign n103 = n102 ^ x4 ;
  assign n104 = x3 & n103 ;
  assign n105 = n104 ^ x3 ;
  assign n106 = ~x2 & ~n105 ;
  assign n107 = x1 & ~n99 ;
  assign n108 = ~n106 & n107 ;
  assign n109 = x0 & x1 ;
  assign n110 = n40 & ~n109 ;
  assign n111 = ~x2 & n110 ;
  assign n112 = x2 & n40 ;
  assign n113 = n112 ^ x2 ;
  assign n114 = n46 & ~n113 ;
  assign n115 = ~n111 & n114 ;
  assign n117 = x4 ^ x1 ;
  assign n119 = n117 ^ x0 ;
  assign n116 = x4 ^ x2 ;
  assign n118 = n117 ^ n116 ;
  assign n120 = n119 ^ n118 ;
  assign n122 = n120 ^ n118 ;
  assign n121 = n120 ^ x4 ;
  assign n123 = n122 ^ n121 ;
  assign n136 = n123 ^ n120 ;
  assign n125 = n120 ^ n117 ;
  assign n126 = n125 ^ n121 ;
  assign n127 = n126 ^ n14 ;
  assign n124 = n123 ^ n121 ;
  assign n128 = n127 ^ n124 ;
  assign n129 = n126 ^ n123 ;
  assign n130 = n126 ^ n120 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = n131 ^ n121 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = n128 & ~n133 ;
  assign n135 = n134 ^ n131 ;
  assign n137 = n136 ^ n135 ;
  assign n138 = n121 ^ n120 ;
  assign n139 = n138 ^ n123 ;
  assign n140 = n139 ^ n127 ;
  assign n141 = ~n14 & ~n140 ;
  assign n142 = n141 ^ n134 ;
  assign n143 = n142 ^ n121 ;
  assign n144 = n143 ^ n129 ;
  assign n145 = n137 & ~n144 ;
  assign n146 = n145 ^ n134 ;
  assign n147 = n146 ^ n121 ;
  assign n148 = n147 ^ n129 ;
  assign n149 = n148 ^ n14 ;
  assign n174 = n14 ^ x4 ;
  assign n150 = n14 ^ x2 ;
  assign n162 = n150 ^ x1 ;
  assign n175 = n174 ^ n162 ;
  assign n151 = n150 ^ n14 ;
  assign n153 = n150 ^ x4 ;
  assign n154 = n151 & n153 ;
  assign n155 = n154 ^ x4 ;
  assign n156 = n155 ^ x0 ;
  assign n161 = n155 ^ n14 ;
  assign n163 = n162 ^ n161 ;
  assign n164 = ~n156 & n163 ;
  assign n172 = n164 ^ n154 ;
  assign n152 = n151 ^ x1 ;
  assign n157 = n156 ^ n152 ;
  assign n158 = n14 ^ x0 ;
  assign n159 = n158 ^ n155 ;
  assign n160 = ~n157 & ~n159 ;
  assign n165 = n164 ^ n160 ;
  assign n166 = n165 ^ n155 ;
  assign n167 = n166 ^ n152 ;
  assign n168 = n164 ^ x0 ;
  assign n169 = n168 ^ x1 ;
  assign n170 = n167 & ~n169 ;
  assign n171 = n170 ^ n160 ;
  assign n173 = n172 ^ n171 ;
  assign n176 = n175 ^ n173 ;
  assign n177 = n176 ^ x1 ;
  assign n178 = n177 ^ x1 ;
  assign n179 = n117 ^ n14 ;
  assign n190 = n179 ^ n116 ;
  assign n202 = n190 ^ n174 ;
  assign n180 = n179 ^ n14 ;
  assign n182 = n179 ^ x4 ;
  assign n183 = n180 & n182 ;
  assign n184 = n183 ^ x4 ;
  assign n185 = n184 ^ x0 ;
  assign n189 = n184 ^ n14 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = ~n185 & n191 ;
  assign n200 = n192 ^ n183 ;
  assign n181 = n180 ^ n116 ;
  assign n186 = n185 ^ n181 ;
  assign n187 = n184 ^ n158 ;
  assign n188 = ~n186 & ~n187 ;
  assign n193 = n192 ^ n188 ;
  assign n194 = n193 ^ n184 ;
  assign n195 = n194 ^ n181 ;
  assign n196 = n192 ^ x0 ;
  assign n197 = n196 ^ n116 ;
  assign n198 = n195 & ~n197 ;
  assign n199 = n198 ^ n188 ;
  assign n201 = n200 ^ n199 ;
  assign n203 = n202 ^ n201 ;
  assign n204 = n203 ^ n116 ;
  assign n205 = n204 ^ n116 ;
  assign n211 = n38 ^ n14 ;
  assign n212 = n211 ^ n38 ;
  assign n228 = n212 ^ n174 ;
  assign n206 = x3 ^ x2 ;
  assign n229 = n228 ^ n206 ;
  assign n215 = n109 ^ x1 ;
  assign n207 = n206 ^ n174 ;
  assign n208 = ~n174 & n207 ;
  assign n216 = n215 ^ n208 ;
  assign n217 = n216 ^ n212 ;
  assign n218 = n217 ^ n207 ;
  assign n219 = n212 ^ n208 ;
  assign n220 = n219 ^ n206 ;
  assign n221 = ~n218 & ~n220 ;
  assign n222 = n221 ^ n215 ;
  assign n223 = n222 ^ n207 ;
  assign n224 = n222 ^ n212 ;
  assign n225 = ~n223 & ~n224 ;
  assign n209 = n208 ^ n206 ;
  assign n210 = n208 ^ n38 ;
  assign n213 = n212 ^ n210 ;
  assign n214 = ~n209 & ~n213 ;
  assign n226 = n225 ^ n214 ;
  assign n227 = n226 ^ n222 ;
  assign n230 = n229 ^ n227 ;
  assign n231 = n230 ^ n38 ;
  assign n232 = ~x0 & ~n46 ;
  assign n233 = n61 & n232 ;
  assign n239 = x1 & ~x3 ;
  assign n240 = ~x4 & ~n239 ;
  assign n234 = n109 ^ x0 ;
  assign n235 = n234 ^ x1 ;
  assign n236 = ~x3 & x4 ;
  assign n237 = n235 & n236 ;
  assign n238 = n237 ^ x3 ;
  assign n241 = n240 ^ n238 ;
  assign n242 = x2 & ~n241 ;
  assign n243 = n242 ^ n241 ;
  assign n244 = n243 ^ n240 ;
  assign n245 = x2 & ~n46 ;
  assign n246 = x0 & n245 ;
  assign n247 = ~n46 & n98 ;
  assign n248 = x3 & ~x4 ;
  assign n249 = ~x1 & n248 ;
  assign n250 = n98 & n249 ;
  assign n251 = x0 & ~x1 ;
  assign n252 = n248 & n251 ;
  assign n253 = x2 & n252 ;
  assign n254 = x2 & n248 ;
  assign n255 = n109 & n254 ;
  assign n256 = n215 & n254 ;
  assign n257 = x2 & ~n110 ;
  assign n263 = ~x2 & n248 ;
  assign n264 = n251 & n263 ;
  assign n265 = n264 ^ x2 ;
  assign n258 = x4 & x5 ;
  assign n259 = n258 ^ x4 ;
  assign n260 = x3 & ~n259 ;
  assign n261 = ~x2 & n109 ;
  assign n262 = n260 & n261 ;
  assign n266 = n265 ^ n262 ;
  assign n267 = ~n257 & n266 ;
  assign n268 = x0 & ~x2 ;
  assign n292 = x6 ^ x4 ;
  assign n280 = n117 ^ x3 ;
  assign n293 = n292 ^ n280 ;
  assign n269 = n117 ^ x4 ;
  assign n271 = n117 ^ x6 ;
  assign n272 = ~n269 & n271 ;
  assign n273 = n272 ^ x6 ;
  assign n274 = n273 ^ x5 ;
  assign n279 = n273 ^ x4 ;
  assign n281 = n280 ^ n279 ;
  assign n282 = ~n274 & n281 ;
  assign n290 = n282 ^ n272 ;
  assign n270 = n269 ^ x3 ;
  assign n275 = n274 ^ n270 ;
  assign n276 = x5 ^ x4 ;
  assign n277 = n276 ^ n273 ;
  assign n278 = n275 & ~n277 ;
  assign n283 = n282 ^ n278 ;
  assign n284 = n283 ^ n273 ;
  assign n285 = n284 ^ n270 ;
  assign n286 = n282 ^ x5 ;
  assign n287 = n286 ^ x3 ;
  assign n288 = n285 & n287 ;
  assign n289 = n288 ^ n278 ;
  assign n291 = n290 ^ n289 ;
  assign n294 = n293 ^ n291 ;
  assign n295 = n294 ^ x3 ;
  assign n296 = n295 ^ x3 ;
  assign n297 = n268 & ~n296 ;
  assign n298 = n297 ^ n268 ;
  assign n300 = x3 & x6 ;
  assign n301 = n259 & n300 ;
  assign n302 = n301 ^ n105 ;
  assign n303 = n261 & n302 ;
  assign n299 = x2 & n110 ;
  assign n304 = n303 ^ n299 ;
  assign n305 = x1 ^ x0 ;
  assign n306 = ~x2 & n41 ;
  assign n307 = ~n305 & n306 ;
  assign n308 = ~x1 & n41 ;
  assign n309 = n268 & n308 ;
  assign y0 = ~n36 ;
  assign y1 = n49 ;
  assign y2 = n59 ;
  assign y3 = n64 ;
  assign y4 = ~n101 ;
  assign y5 = n108 ;
  assign y6 = n115 ;
  assign y7 = n149 ;
  assign y8 = n178 ;
  assign y9 = n205 ;
  assign y10 = n231 ;
  assign y11 = n233 ;
  assign y12 = n244 ;
  assign y13 = n246 ;
  assign y14 = n247 ;
  assign y15 = n250 ;
  assign y16 = n253 ;
  assign y17 = n255 ;
  assign y18 = n256 ;
  assign y19 = n245 ;
  assign y20 = n267 ;
  assign y21 = n298 ;
  assign y22 = n304 ;
  assign y23 = ~1'b0 ;
  assign y24 = n307 ;
  assign y25 = n309 ;
endmodule
