module bitonic_sort_inc_2_8 (in_array_0, in_array_1, in_array_2, in_array_3, in_array_4, in_array_5, in_array_6, in_array_7, in_array_8, in_array_9, in_array_10, in_array_11, in_array_12, in_array_13, in_array_14, in_array_15, out_array_0, out_array_1, out_array_2, out_array_3, out_array_4, out_array_5, out_array_6, out_array_7, out_array_8, out_array_9, out_array_10, out_array_11, out_array_12, out_array_13, out_array_14, out_array_15);
input in_array_0, in_array_1, in_array_2, in_array_3, in_array_4, in_array_5, in_array_6, in_array_7, in_array_8, in_array_9, in_array_10, in_array_11, in_array_12, in_array_13, in_array_14, in_array_15;
output out_array_0, out_array_1, out_array_2, out_array_3, out_array_4, out_array_5, out_array_6, out_array_7, out_array_8, out_array_9, out_array_10, out_array_11, out_array_12, out_array_13, out_array_14, out_array_15;
wire _000_, _001_, _002_, _003_, _004_, _005_, _006_, _007_, _008_, _009_, _010_, _011_, _012_, _013_, _014_, _015_, _016_, _017_, _018_, _019_, _020_, _021_, _022_, _023_, _023__neg, _024_, _025_, _026_, _027_, _028_, _029_, _030_, _031_, _032_, _033_, _034_, _035_, _036_, _037_, _038_, _039_, _040_, _040__neg, _041_, _042_, _043_, _044_, _045_, _046_, _047_, _048_, _049_, _050_, _051_, _052_, _052__neg, _053_, _054_, _054__neg, _055_, _056_, _057_, _058_, _058__neg, _059_, _060_, _061_, _062_, _063_, _064_, _065_, _066_, _066__neg, _067_, _068_, _069_, _070_, _071_, _072_, _073_, _074_, _075_, _076_, _077_, _078_, _079_, _079__neg, _080_, _081_, _082_, _083_, _084_, _085_, _086_, _087_, _088_, _088__neg, _089_, _090_, _091_, _092_, _093_, _094_, _095_, _096_, _097_, _098_, _099_, _100_, _101_, _102_, _103_, _104_, _104__neg, _105_, _106_, _107_, _108_, _109_, _110_, _111_, _112_, _113_, _114_, _115_, _115__neg, _116_, _117_, _118_, _119_, _120_, _121_, _122_, _123_, _124_, _125_, _126_, _126__neg, _127_, _128_, _129_, _130_, _131_, _132_, _132__neg, _133_, _134_, _135_, _135__neg, _136_, _137_, _138_, _139_, _140_, _140__neg, _141_, _142_, _143_, _144_, _145_, _146_, _147_, _148_, _149_, _150_, _151_, _152_, _152__neg, _153_, _154_, _155_, _156_, _157_, _158_, _159_, _160_, _161_, _162_, _163_, _164_, _165_, _166_, _167_, _168_, _168__neg, _169_, _170_, _171_, _172_, _173_, _174_, _175_, _176_, _177_, _178_, _179_, _180_, _180__neg, _181_, _182_, _183_, _183__neg, _184_, _185_, _186_, _187_, _188_, _188__neg, _189_, _190_, _191_, _192_, _193_, _194_, _195_, _196_, _196__neg, _197_, _198_, _199_, _200_, _200__neg, _201_, _202_, _203_, _204_, _204__neg, _205_, _206_, _207_, _208_, _209_, _210_, _211_, _212_, _212__neg, _213_, _214_, _215_, _216_, _217_, _217__neg, _218_, _219_, _220_, _221_, _222_, _223_, _224_, _225_, _226_, _227_, _228_, _229_, _230_, _230__neg, _231_, _232_, _233_, _234_, _235_, _236_, _237_, _238_, _238__neg, _239_, _240_, _241_, _242_, _243_, _244_, _245_, _246_, _247_, _248_, _249_, _250_, _251_, _252_, _253_, _254_, _255_, _256_, _256__neg, _257_, _258_, _259_, _260_, _261_, _262_, _263_, _264_, _265_, _266_, _267_, _268_, _269_, _269__neg, _270_, _271_, _272_, _273_, _273__neg, _274_, _275_, _276_, _277_, _278_, _278__neg, _279_, _280_, _281_, _282_, _283_, _284_, _285_, _286_, _287_, _287__neg, _288_, _289_, _290_, _291_, _292_, _292__neg, _293_, _294_, _295_, _296_, _297_, _298_, _299_, _300_, _301_, _302_, _303_, _304_, _305_, _306_, _306__neg, _307_, _308_, _309_, _310_, _311_, _312_, _313_, _314_, _315_, _316_, _317_, _318_, _319_, _320_, _321_, _322_, _323_, _323__neg, _324_, _325_, _326_, _327_, _328_, _329_, _330_, _331_, _332_, _333_, _334_, _335_, _336_, _337_, _338_, _339_, _340_, _340__neg, _341_, _342_, _343_, _344_, _345_, _346_, _347_, _348_, _349_, _350_, _351_, _352_, _353_, _353__neg, _354_, _355_, _356_, _356__neg, _357_, _358_, _359_, _360_, _360__neg, _361_, _362_, _363_, _364_, _365_, _366_, _367_;
assign _347_ = ~_346_;
assign _348_ = _347_ ^ _341_;
assign _349_ = _348_ & _345_;
assign _350_ = _349_ ^ _342_;
assign _351_ = _350_ & _340_;
assign _352_ = _351_ ^ _338_;
assign _353__neg = _352_ ^ _336_;
assign _353_ = ~_353__neg;
assign _354_ = _352_ & _336_;
assign _355_ = ~_354_;
assign _356__neg = _331_ ^ _328_;
assign _356_ = ~_356__neg;
assign _357_ = _356_ & _334_;
assign _358_ = _357_ ^ _328_;
assign _359_ = _358_ ^ _354_;
assign _360__neg = _346_ ^ _343_;
assign _360_ = ~_360__neg;
assign _361_ = _360_ & _350_;
assign _362_ = _361_ ^ _343_;
assign _363_ = _362_ ^ _354_;
assign _364_ = _363_ & _359_;
assign _365_ = _364_ ^ _355_;
assign _366_ = _365_ & _353_;
assign _367_ = _366_ ^ _336_;
assign _000_ = ~_367_;
assign _001_ = ~in_array_10;
assign _002_ = in_array_10 ^ in_array_8;
assign _003_ = ~in_array_8;
assign _004_ = in_array_10 & _003_;
assign _005_ = ~_004_;
assign _006_ = ~in_array_9;
assign _007_ = _004_ ^ _006_;
assign _008_ = _004_ ^ in_array_11;
assign _009_ = _008_ & _007_;
assign _010_ = _009_ ^ _005_;
assign _011_ = _010_ & _002_;
assign _012_ = _011_ ^ _001_;
assign _013_ = in_array_14 ^ in_array_12;
assign _014_ = ~in_array_12;
assign _015_ = in_array_14 & _014_;
assign _016_ = ~in_array_13;
assign _017_ = _015_ ^ _016_;
assign _018_ = _015_ ^ in_array_15;
assign _019_ = _018_ & _017_;
assign _020_ = _019_ ^ _015_;
assign _021_ = _020_ & _013_;
assign _022_ = _021_ ^ in_array_14;
assign _023__neg = _022_ ^ _012_;
assign _023_ = ~_023__neg;
assign _024_ = _022_ & _012_;
assign _025_ = ~in_array_11;
assign _026_ = in_array_9 & _025_;
assign _027_ = _026_ ^ _025_;
assign _028_ = _027_ ^ _024_;
assign _029_ = _016_ & in_array_15;
assign _030_ = _029_ ^ in_array_15;
assign _031_ = _030_ ^ _024_;
assign _032_ = _031_ & _028_;
assign _033_ = _032_ ^ _024_;
assign _034_ = _033_ & _023_;
assign _035_ = _034_ ^ _012_;
assign _036_ = ~_035_;
assign _037_ = _011_ ^ _003_;
assign _038_ = ~_037_;
assign _039_ = _021_ ^ in_array_12;
assign _040__neg = _039_ ^ _037_;
assign _040_ = ~_040__neg;
assign _041_ = _039_ & _037_;
assign _042_ = _026_ ^ in_array_9;
assign _043_ = ~_042_;
assign _044_ = _043_ ^ _041_;
assign _045_ = _029_ ^ _016_;
assign _046_ = ~_045_;
assign _047_ = _046_ ^ _041_;
assign _048_ = _047_ & _044_;
assign _049_ = _048_ ^ _041_;
assign _050_ = _049_ & _040_;
assign _051_ = _050_ ^ _038_;
assign _052__neg = _051_ ^ _035_;
assign _052_ = ~_052__neg;
assign _053_ = _051_ & _035_;
assign _054__neg = _030_ ^ _027_;
assign _054_ = ~_054__neg;
assign _055_ = _054_ & _033_;
assign _056_ = _055_ ^ _027_;
assign _057_ = _056_ ^ _053_;
assign _058__neg = _045_ ^ _042_;
assign _058_ = ~_058__neg;
assign _059_ = _058_ & _049_;
assign _060_ = _059_ ^ _042_;
assign _061_ = _060_ ^ _053_;
assign _062_ = _061_ & _057_;
assign _063_ = _062_ ^ _053_;
assign _064_ = _063_ & _052_;
assign _065_ = _064_ ^ _036_;
assign _066__neg = _065_ ^ _367_;
assign _066_ = ~_066__neg;
assign _067_ = _065_ & _367_;
assign _068_ = ~_067_;
assign _069_ = ~_328_;
assign _070_ = _357_ ^ _069_;
assign _071_ = _362_ ^ _070_;
assign _072_ = _071_ & _365_;
assign _073_ = _072_ ^ _358_;
assign _074_ = _073_ ^ _067_;
assign _075_ = ~_027_;
assign _076_ = _055_ ^ _075_;
assign _077_ = _060_ ^ _076_;
assign _078_ = _077_ & _063_;
assign _079__neg = _078_ ^ _056_;
assign _079_ = ~_079__neg;
assign _080_ = _079_ ^ _067_;
assign _081_ = _080_ & _074_;
assign _082_ = _081_ ^ _068_;
assign _083_ = _082_ & _066_;
assign _084_ = _083_ ^ _000_;
assign _085_ = ~_322_;
assign _086_ = _335_ ^ _085_;
assign _087_ = _351_ ^ _339_;
assign _088__neg = _087_ ^ _086_;
assign _088_ = ~_088__neg;
assign _089_ = _087_ & _086_;
assign _090_ = ~_089_;
assign _091_ = ~_331_;
assign _092_ = _357_ ^ _091_;
assign _093_ = _092_ ^ _089_;
assign _094_ = _361_ ^ _347_;
assign _095_ = _094_ ^ _089_;
assign _096_ = _095_ & _093_;
assign _097_ = _096_ ^ _090_;
assign _098_ = _097_ & _088_;
assign _099_ = _098_ ^ _086_;
assign _100_ = ~_022_;
assign _101_ = _034_ ^ _100_;
assign _102_ = ~_101_;
assign _103_ = _050_ ^ _039_;
assign _104__neg = _103_ ^ _101_;
assign _104_ = ~_104__neg;
assign _105_ = _103_ & _101_;
assign _106_ = ~_030_;
assign _107_ = _055_ ^ _106_;
assign _108_ = _107_ ^ _105_;
assign _109_ = _059_ ^ _046_;
assign _110_ = _109_ ^ _105_;
assign _111_ = _110_ & _108_;
assign _112_ = _111_ ^ _105_;
assign _113_ = _112_ & _104_;
assign _114_ = _113_ ^ _102_;
assign _115__neg = _114_ ^ _099_;
assign _115_ = ~_115__neg;
assign _116_ = _114_ & _099_;
assign _117_ = ~_116_;
assign _118_ = _357_ ^ _331_;
assign _119_ = _094_ ^ _118_;
assign _120_ = _119_ & _097_;
assign _121_ = _120_ ^ _092_;
assign _122_ = _121_ ^ _116_;
assign _123_ = _055_ ^ _030_;
assign _124_ = _109_ ^ _123_;
assign _125_ = _124_ & _112_;
assign _126__neg = _125_ ^ _107_;
assign _126_ = ~_126__neg;
assign _127_ = _126_ ^ _116_;
assign _128_ = _127_ & _122_;
assign _129_ = _128_ ^ _117_;
assign _130_ = _129_ & _115_;
assign _131_ = _130_ ^ _099_;
assign _132__neg = _131_ ^ _084_;
assign _132_ = ~_132__neg;
assign _133_ = _131_ & _084_;
assign _134_ = ~_133_;
assign _135__neg = _126_ ^ _121_;
assign _135_ = ~_135__neg;
assign _136_ = _135_ & _129_;
assign _137_ = _136_ ^ _121_;
assign _138_ = _137_ ^ _133_;
assign _139_ = ~_073_;
assign _140__neg = _079_ ^ _073_;
assign _140_ = ~_140__neg;
assign _141_ = _140_ & _082_;
assign _142_ = _141_ ^ _139_;
assign _143_ = _142_ ^ _133_;
assign _144_ = _143_ & _138_;
assign _145_ = _144_ ^ _134_;
assign _146_ = _145_ & _132_;
assign _147_ = _146_ ^ _084_;
assign _148_ = ~_352_;
assign _149_ = _366_ ^ _148_;
assign _150_ = ~_149_;
assign _151_ = _064_ ^ _051_;
assign _152__neg = _151_ ^ _149_;
assign _152_ = ~_152__neg;
assign _153_ = _151_ & _149_;
assign _154_ = ~_153_;
assign _155_ = ~_362_;
assign _156_ = _072_ ^ _155_;
assign _157_ = _156_ ^ _153_;
assign _158_ = _078_ ^ _060_;
assign _159_ = _158_ ^ _153_;
assign _160_ = _159_ & _157_;
assign _161_ = _160_ ^ _154_;
assign _162_ = _161_ & _152_;
assign _163_ = _162_ ^ _150_;
assign _164_ = ~_163_;
assign _165_ = ~_087_;
assign _166_ = _098_ ^ _165_;
assign _167_ = _113_ ^ _103_;
assign _168__neg = _167_ ^ _166_;
assign _168_ = ~_168__neg;
assign _169_ = _167_ & _166_;
assign _170_ = ~_169_;
assign _171_ = ~_094_;
assign _172_ = _120_ ^ _171_;
assign _173_ = _172_ ^ _169_;
assign _174_ = _125_ ^ _109_;
assign _175_ = _174_ ^ _169_;
assign _176_ = _175_ & _173_;
assign _177_ = _176_ ^ _170_;
assign _178_ = _177_ & _168_;
assign _179_ = _178_ ^ _166_;
assign _180__neg = _179_ ^ _163_;
assign _180_ = ~_180__neg;
assign _181_ = _179_ & _163_;
assign _182_ = ~_181_;
assign _183__neg = _174_ ^ _172_;
assign _183_ = ~_183__neg;
assign _184_ = _183_ & _177_;
assign _185_ = _184_ ^ _172_;
assign _186_ = _185_ ^ _181_;
assign _187_ = ~_156_;
assign _188__neg = _158_ ^ _156_;
assign _188_ = ~_188__neg;
assign _189_ = _188_ & _161_;
assign _190_ = _189_ ^ _187_;
assign _191_ = _190_ ^ _181_;
assign _192_ = _191_ & _186_;
assign _193_ = _192_ ^ _182_;
assign _194_ = _193_ & _180_;
assign _195_ = _194_ ^ _164_;
assign _196__neg = _195_ ^ _147_;
assign _196_ = ~_196__neg;
assign _197_ = _195_ & _147_;
assign _198_ = ~_197_;
assign _199_ = ~_190_;
assign _200__neg = _190_ ^ _185_;
assign _200_ = ~_200__neg;
assign _201_ = _200_ & _193_;
assign _202_ = _201_ ^ _199_;
assign _203_ = _202_ ^ _197_;
assign _204__neg = _142_ ^ _137_;
assign _204_ = ~_204__neg;
assign _205_ = _204_ & _145_;
assign _206_ = _205_ ^ _142_;
assign _207_ = _206_ ^ _197_;
assign _208_ = _207_ & _203_;
assign _209_ = _208_ ^ _198_;
assign _210_ = _209_ & _196_;
assign out_array_8 = _210_ ^ _147_;
assign _211_ = ~_195_;
assign out_array_10 = _210_ ^ _211_;
assign _212__neg = _206_ ^ _202_;
assign _212_ = ~_212__neg;
assign _213_ = _212_ & _209_;
assign out_array_9 = _213_ ^ _206_;
assign _214_ = ~_131_;
assign _215_ = _146_ ^ _214_;
assign _216_ = _194_ ^ _179_;
assign _217__neg = _216_ ^ _215_;
assign _217_ = ~_217__neg;
assign _218_ = _216_ & _215_;
assign _219_ = ~_218_;
assign _220_ = _201_ ^ _185_;
assign _221_ = _220_ ^ _218_;
assign _222_ = ~_137_;
assign _223_ = _205_ ^ _222_;
assign _224_ = _223_ ^ _218_;
assign _225_ = _224_ & _221_;
assign _226_ = _225_ ^ _219_;
assign _228_ = _226_ & _217_;
assign out_array_12 = _228_ ^ _215_;
assign _229_ = ~_216_;
assign out_array_14 = _228_ ^ _229_;
assign _230__neg = _223_ ^ _220_;
assign _230_ = ~_230__neg;
assign _231_ = _230_ & _226_;
assign out_array_13 = _231_ ^ _223_;
assign _232_ = ~_202_;
assign out_array_11 = _213_ ^ _232_;
assign _233_ = ~_220_;
assign out_array_15 = _231_ ^ _233_;
assign _235_ = _083_ ^ _065_;
assign _236_ = ~_114_;
assign _237_ = _130_ ^ _236_;
assign _238__neg = _237_ ^ _235_;
assign _238_ = ~_238__neg;
assign _239_ = _237_ & _235_;
assign _240_ = ~_239_;
assign _241_ = ~_126_;
assign _242_ = _136_ ^ _241_;
assign _243_ = _242_ ^ _239_;
assign _245_ = _141_ ^ _079_;
assign _246_ = _245_ ^ _239_;
assign _247_ = _246_ & _243_;
assign _248_ = _247_ ^ _240_;
assign _249_ = _248_ & _238_;
assign _250_ = _249_ ^ _235_;
assign _251_ = _162_ ^ _151_;
assign _252_ = ~_251_;
assign _253_ = ~_167_;
assign _254_ = _178_ ^ _253_;
assign _256__neg = _254_ ^ _251_;
assign _256_ = ~_256__neg;
assign _257_ = _254_ & _251_;
assign _258_ = ~_257_;
assign _259_ = ~_174_;
assign _260_ = _184_ ^ _259_;
assign _261_ = _260_ ^ _257_;
assign _262_ = _189_ ^ _158_;
assign _263_ = _262_ ^ _257_;
assign _264_ = _263_ & _261_;
assign _265_ = _264_ ^ _258_;
assign _267_ = _265_ & _256_;
assign _268_ = _267_ ^ _252_;
assign _269__neg = _268_ ^ _250_;
assign _269_ = ~_269__neg;
assign _270_ = _268_ & _250_;
assign _271_ = ~_270_;
assign _272_ = ~_262_;
assign _273__neg = _262_ ^ _260_;
assign _273_ = ~_273__neg;
assign _274_ = _273_ & _265_;
assign _275_ = _274_ ^ _272_;
assign _276_ = _275_ ^ _270_;
assign _278__neg = _245_ ^ _242_;
assign _278_ = ~_278__neg;
assign _279_ = _278_ & _248_;
assign _280_ = _279_ ^ _245_;
assign _281_ = _280_ ^ _270_;
assign _282_ = _281_ & _276_;
assign _283_ = _282_ ^ _271_;
assign _284_ = _283_ & _269_;
assign out_array_0 = _284_ ^ _250_;
assign _285_ = ~_268_;
assign out_array_2 = _284_ ^ _285_;
assign _287__neg = _280_ ^ _275_;
assign _287_ = ~_287__neg;
assign _288_ = _287_ & _283_;
assign out_array_1 = _288_ ^ _280_;
assign _289_ = ~_237_;
assign _290_ = _249_ ^ _289_;
assign _291_ = _267_ ^ _254_;
assign _292__neg = _291_ ^ _290_;
assign _292_ = ~_292__neg;
assign _293_ = _291_ & _290_;
assign _294_ = ~_293_;
assign _295_ = _274_ ^ _260_;
assign _297_ = _295_ ^ _293_;
assign _298_ = ~_242_;
assign _299_ = _279_ ^ _298_;
assign _300_ = _299_ ^ _293_;
assign _301_ = _300_ & _297_;
assign _302_ = _301_ ^ _294_;
assign _303_ = _302_ & _292_;
assign out_array_4 = _303_ ^ _290_;
assign _304_ = ~_291_;
assign out_array_6 = _303_ ^ _304_;
assign _306__neg = _299_ ^ _295_;
assign _306_ = ~_306__neg;
assign _307_ = _306_ & _302_;
assign out_array_5 = _307_ ^ _299_;
assign _308_ = ~_275_;
assign out_array_3 = _288_ ^ _308_;
assign _309_ = ~_295_;
assign out_array_7 = _307_ ^ _309_;
assign _227_ = ~in_array_2;
assign _234_ = in_array_2 ^ in_array_0;
assign _244_ = ~in_array_0;
assign _255_ = in_array_2 & _244_;
assign _266_ = ~_255_;
assign _277_ = ~in_array_1;
assign _286_ = _255_ ^ _277_;
assign _296_ = _255_ ^ in_array_3;
assign _305_ = _296_ & _286_;
assign _310_ = _305_ ^ _266_;
assign _311_ = _310_ & _234_;
assign _312_ = _311_ ^ _227_;
assign _313_ = in_array_6 ^ in_array_4;
assign _314_ = ~in_array_4;
assign _315_ = in_array_6 & _314_;
assign _316_ = ~in_array_5;
assign _317_ = _315_ ^ _316_;
assign _318_ = _315_ ^ in_array_7;
assign _319_ = _318_ & _317_;
assign _320_ = _319_ ^ _315_;
assign _321_ = _320_ & _313_;
assign _322_ = _321_ ^ in_array_6;
assign _323__neg = _322_ ^ _312_;
assign _323_ = ~_323__neg;
assign _324_ = _322_ & _312_;
assign _325_ = ~_324_;
assign _326_ = ~in_array_3;
assign _327_ = in_array_1 & _326_;
assign _328_ = _327_ ^ _326_;
assign _329_ = _328_ ^ _324_;
assign _330_ = _316_ & in_array_7;
assign _331_ = _330_ ^ in_array_7;
assign _332_ = _331_ ^ _324_;
assign _333_ = _332_ & _329_;
assign _334_ = _333_ ^ _325_;
assign _335_ = _334_ & _323_;
assign _336_ = _335_ ^ _312_;
assign _337_ = _311_ ^ _244_;
assign _338_ = ~_337_;
assign _339_ = _321_ ^ in_array_4;
assign _340__neg = _339_ ^ _337_;
assign _340_ = ~_340__neg;
assign _341_ = _339_ & _337_;
assign _342_ = ~_341_;
assign _343_ = _327_ ^ in_array_1;
assign _344_ = ~_343_;
assign _345_ = _344_ ^ _341_;
assign _346_ = _330_ ^ _316_;
endmodule
