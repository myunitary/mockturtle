// Benchmark "/tmp/tmp" written by ABC on Wed Nov 12 17:42:45 2025

module max_opt ( 
    n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
    n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127, po128, po129  );
  input  n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
    n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
    n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127, po128, po129;
  wire new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1364, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1374, new_n1375, new_n1376, new_n1377, new_n1378, new_n1379,
    new_n1380, new_n1381, new_n1382, new_n1383, new_n1384, new_n1385,
    new_n1386, new_n1387, new_n1388, new_n1389, new_n1390, new_n1391,
    new_n1392, new_n1393, new_n1394, new_n1395, new_n1396, new_n1397,
    new_n1398, new_n1399, new_n1400, new_n1401, new_n1402, new_n1403,
    new_n1404, new_n1405, new_n1406, new_n1407, new_n1408, new_n1409,
    new_n1410, new_n1411, new_n1412, new_n1413, new_n1414, new_n1415,
    new_n1416, new_n1417, new_n1418, new_n1419, new_n1420, new_n1421,
    new_n1422, new_n1423, new_n1424, new_n1425, new_n1426, new_n1427,
    new_n1428, new_n1429, new_n1430, new_n1431, new_n1432, new_n1433,
    new_n1434, new_n1435, new_n1436, new_n1437, new_n1438, new_n1439,
    new_n1440, new_n1441, new_n1442, new_n1443, new_n1444, new_n1445,
    new_n1446, new_n1447, new_n1448, new_n1449, new_n1450, new_n1451,
    new_n1452, new_n1453, new_n1454, new_n1455, new_n1456, new_n1457,
    new_n1458, new_n1459, new_n1460, new_n1461, new_n1462, new_n1463,
    new_n1464, new_n1465, new_n1466, new_n1467, new_n1468, new_n1469,
    new_n1470, new_n1471, new_n1472, new_n1473, new_n1474, new_n1475,
    new_n1476, new_n1477, new_n1478, new_n1479, new_n1480, new_n1481,
    new_n1482, new_n1483, new_n1484, new_n1485, new_n1486, new_n1487,
    new_n1488, new_n1489, new_n1490, new_n1491, new_n1492, new_n1493,
    new_n1494, new_n1495, new_n1496, new_n1497, new_n1498, new_n1499,
    new_n1500, new_n1501, new_n1502, new_n1503, new_n1504, new_n1505,
    new_n1506, new_n1507, new_n1508, new_n1509, new_n1510, new_n1511,
    new_n1512, new_n1513, new_n1514, new_n1515, new_n1516, new_n1517,
    new_n1518, new_n1519, new_n1520, new_n1521, new_n1522, new_n1523,
    new_n1524, new_n1525, new_n1526, new_n1527, new_n1528, new_n1529,
    new_n1530, new_n1531, new_n1532, new_n1533, new_n1534, new_n1535,
    new_n1536, new_n1537, new_n1538, new_n1539, new_n1540, new_n1541,
    new_n1542, new_n1543, new_n1544, new_n1545, new_n1546, new_n1547,
    new_n1548, new_n1549, new_n1550, new_n1551, new_n1552, new_n1553,
    new_n1554, new_n1555, new_n1556, new_n1557, new_n1558, new_n1559,
    new_n1560, new_n1561, new_n1562, new_n1563, new_n1564, new_n1565,
    new_n1566, new_n1567, new_n1568, new_n1569, new_n1570, new_n1571,
    new_n1572, new_n1573, new_n1574, new_n1575, new_n1576, new_n1577,
    new_n1578, new_n1579, new_n1580, new_n1581, new_n1582, new_n1583,
    new_n1584, new_n1585, new_n1586, new_n1587, new_n1588, new_n1589,
    new_n1590, new_n1591, new_n1592, new_n1593, new_n1594, new_n1595,
    new_n1596, new_n1597, new_n1598, new_n1599, new_n1600, new_n1601,
    new_n1602, new_n1603, new_n1604, new_n1605, new_n1606, new_n1607,
    new_n1608, new_n1609, new_n1610, new_n1611, new_n1612, new_n1613,
    new_n1614, new_n1615, new_n1616, new_n1617, new_n1618, new_n1619,
    new_n1620, new_n1621, new_n1622, new_n1623, new_n1624, new_n1625,
    new_n1626, new_n1627, new_n1628, new_n1629, new_n1630, new_n1631,
    new_n1632, new_n1633, new_n1634, new_n1635, new_n1636, new_n1637,
    new_n1638, new_n1639, new_n1640, new_n1641, new_n1642, new_n1643,
    new_n1644, new_n1645, new_n1646, new_n1647, new_n1648, new_n1649,
    new_n1650, new_n1651, new_n1652, new_n1653, new_n1654, new_n1655,
    new_n1656, new_n1657, new_n1658, new_n1659, new_n1660, new_n1661,
    new_n1662, new_n1663, new_n1664, new_n1665, new_n1666, new_n1667,
    new_n1668, new_n1669, new_n1670, new_n1671, new_n1672, new_n1673,
    new_n1674, new_n1675, new_n1676, new_n1677, new_n1678, new_n1679,
    new_n1680, new_n1681, new_n1682, new_n1683, new_n1684, new_n1685,
    new_n1686, new_n1687, new_n1688, new_n1689, new_n1690, new_n1691,
    new_n1692, new_n1693, new_n1694, new_n1695, new_n1696, new_n1697,
    new_n1698, new_n1699, new_n1700, new_n1701, new_n1702, new_n1703,
    new_n1704, new_n1705, new_n1706, new_n1707, new_n1708, new_n1709,
    new_n1710, new_n1711, new_n1712, new_n1713, new_n1714, new_n1715,
    new_n1716, new_n1717, new_n1718, new_n1719, new_n1720, new_n1721,
    new_n1722, new_n1723, new_n1724, new_n1725, new_n1726, new_n1727,
    new_n1728, new_n1729, new_n1730, new_n1731, new_n1732, new_n1733,
    new_n1734, new_n1735, new_n1736, new_n1737, new_n1738, new_n1739,
    new_n1740, new_n1741, new_n1742, new_n1743, new_n1744, new_n1745,
    new_n1746, new_n1747, new_n1748, new_n1749, new_n1750, new_n1751,
    new_n1752, new_n1753, new_n1754, new_n1755, new_n1756, new_n1757,
    new_n1758, new_n1759, new_n1760, new_n1761, new_n1762, new_n1763,
    new_n1764, new_n1765, new_n1766, new_n1767, new_n1768, new_n1769,
    new_n1770, new_n1771, new_n1772, new_n1773, new_n1774, new_n1775,
    new_n1776, new_n1777, new_n1778, new_n1779, new_n1780, new_n1781,
    new_n1782, new_n1783, new_n1784, new_n1785, new_n1786, new_n1787,
    new_n1788, new_n1789, new_n1790, new_n1791, new_n1792, new_n1793,
    new_n1794, new_n1795, new_n1796, new_n1797, new_n1798, new_n1799,
    new_n1800, new_n1801, new_n1802, new_n1803, new_n1804, new_n1805,
    new_n1806, new_n1807, new_n1808, new_n1809, new_n1810, new_n1811,
    new_n1812, new_n1813, new_n1814, new_n1815, new_n1816, new_n1817,
    new_n1818, new_n1819, new_n1820, new_n1821, new_n1822, new_n1823,
    new_n1824, new_n1825, new_n1826, new_n1827, new_n1828, new_n1829,
    new_n1830, new_n1831, new_n1832, new_n1833, new_n1834, new_n1835,
    new_n1836, new_n1837, new_n1838, new_n1839, new_n1840, new_n1841,
    new_n1842, new_n1843, new_n1844, new_n1845, new_n1846, new_n1847,
    new_n1848, new_n1849, new_n1850, new_n1851, new_n1852, new_n1853,
    new_n1854, new_n1855, new_n1856, new_n1857, new_n1858, new_n1859,
    new_n1860, new_n1861, new_n1862, new_n1863, new_n1864, new_n1865,
    new_n1866, new_n1867, new_n1868, new_n1869, new_n1870, new_n1871,
    new_n1872, new_n1873, new_n1874, new_n1875, new_n1876, new_n1877,
    new_n1878, new_n1879, new_n1880, new_n1881, new_n1882, new_n1883,
    new_n1884, new_n1885, new_n1886, new_n1887, new_n1888, new_n1889,
    new_n1890, new_n1891, new_n1892, new_n1893, new_n1894, new_n1895,
    new_n1896, new_n1897, new_n1898, new_n1899, new_n1900, new_n1901,
    new_n1902, new_n1903, new_n1904, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1909, new_n1910, new_n1911, new_n1912, new_n1913,
    new_n1914, new_n1915, new_n1916, new_n1917, new_n1918, new_n1919,
    new_n1920, new_n1921, new_n1922, new_n1923, new_n1924, new_n1925,
    new_n1926, new_n1927, new_n1928, new_n1929, new_n1930, new_n1931,
    new_n1932, new_n1933, new_n1934, new_n1935, new_n1936, new_n1937,
    new_n1938, new_n1939, new_n1940, new_n1941, new_n1942, new_n1943,
    new_n1944, new_n1945, new_n1946, new_n1947, new_n1948, new_n1949,
    new_n1950, new_n1951, new_n1952, new_n1953, new_n1954, new_n1955,
    new_n1956, new_n1957, new_n1958, new_n1959, new_n1960, new_n1961,
    new_n1962, new_n1963, new_n1964, new_n1965, new_n1966, new_n1967,
    new_n1968, new_n1969, new_n1970, new_n1971, new_n1972, new_n1973,
    new_n1974, new_n1975, new_n1976, new_n1977, new_n1978, new_n1979,
    new_n1980, new_n1981, new_n1982, new_n1983, new_n1984, new_n1985,
    new_n1986, new_n1987, new_n1988, new_n1989, new_n1990, new_n1991,
    new_n1992, new_n1993, new_n1994, new_n1995, new_n1996, new_n1997,
    new_n1998, new_n1999, new_n2000, new_n2001, new_n2002, new_n2003,
    new_n2004, new_n2005, new_n2006, new_n2007, new_n2008, new_n2009,
    new_n2010, new_n2011, new_n2012, new_n2013, new_n2014, new_n2015,
    new_n2016, new_n2017, new_n2018, new_n2019, new_n2020, new_n2021,
    new_n2022, new_n2023, new_n2024, new_n2025, new_n2026, new_n2027,
    new_n2028, new_n2029, new_n2030, new_n2031, new_n2032, new_n2033,
    new_n2034, new_n2035, new_n2036, new_n2037, new_n2038, new_n2039,
    new_n2040, new_n2041, new_n2042, new_n2043, new_n2044, new_n2045,
    new_n2046, new_n2047, new_n2048, new_n2049, new_n2050, new_n2051,
    new_n2052, new_n2053, new_n2054, new_n2055, new_n2056, new_n2057,
    new_n2058, new_n2059, new_n2060, new_n2061, new_n2062, new_n2063,
    new_n2064, new_n2065, new_n2066, new_n2067, new_n2068, new_n2069,
    new_n2070, new_n2071, new_n2072, new_n2073, new_n2074, new_n2075,
    new_n2076, new_n2077, new_n2078, new_n2079, new_n2080, new_n2081,
    new_n2082, new_n2083, new_n2084, new_n2085, new_n2086, new_n2087,
    new_n2088, new_n2089, new_n2090, new_n2091, new_n2092, new_n2093,
    new_n2094, new_n2095, new_n2096, new_n2097, new_n2098, new_n2099,
    new_n2100, new_n2101, new_n2102, new_n2103, new_n2104, new_n2105,
    new_n2106, new_n2107, new_n2108, new_n2109, new_n2110, new_n2111,
    new_n2112, new_n2113, new_n2114, new_n2115, new_n2116, new_n2117,
    new_n2118, new_n2119, new_n2120, new_n2121, new_n2122, new_n2123,
    new_n2124, new_n2125, new_n2126, new_n2127, new_n2128, new_n2129,
    new_n2130, new_n2131, new_n2132, new_n2133, new_n2134, new_n2135,
    new_n2136, new_n2137, new_n2138, new_n2139, new_n2140, new_n2141,
    new_n2142, new_n2143, new_n2144, new_n2145, new_n2146, new_n2147,
    new_n2148, new_n2149, new_n2150, new_n2151, new_n2152, new_n2153,
    new_n2154, new_n2155, new_n2156, new_n2157, new_n2158, new_n2159,
    new_n2160, new_n2161, new_n2162, new_n2163, new_n2164, new_n2165,
    new_n2166, new_n2167, new_n2168, new_n2169, new_n2170, new_n2171,
    new_n2172, new_n2173, new_n2174, new_n2175, new_n2176, new_n2177,
    new_n2178, new_n2179, new_n2180, new_n2181, new_n2182, new_n2183,
    new_n2184, new_n2185, new_n2186, new_n2187, new_n2188, new_n2189,
    new_n2190, new_n2191, new_n2192, new_n2193, new_n2194, new_n2195,
    new_n2196, new_n2197, new_n2198, new_n2199, new_n2200, new_n2201,
    new_n2202, new_n2203, new_n2204, new_n2205, new_n2206, new_n2207,
    new_n2208, new_n2209, new_n2210, new_n2211, new_n2212, new_n2213,
    new_n2214, new_n2215, new_n2216, new_n2217, new_n2218, new_n2219,
    new_n2220, new_n2221, new_n2222, new_n2223, new_n2224, new_n2225,
    new_n2226, new_n2227, new_n2228, new_n2229, new_n2230, new_n2231,
    new_n2232, new_n2233, new_n2234, new_n2235, new_n2236, new_n2237,
    new_n2238, new_n2239, new_n2240, new_n2241, new_n2242, new_n2243,
    new_n2244, new_n2245, new_n2246, new_n2247, new_n2248, new_n2249,
    new_n2250, new_n2251, new_n2252, new_n2253, new_n2254, new_n2255,
    new_n2256, new_n2257, new_n2258, new_n2259, new_n2260, new_n2261,
    new_n2262, new_n2263, new_n2264, new_n2265, new_n2266, new_n2267,
    new_n2268, new_n2269, new_n2270, new_n2271, new_n2272, new_n2273,
    new_n2274, new_n2275, new_n2276, new_n2277, new_n2278, new_n2279,
    new_n2280, new_n2281, new_n2282, new_n2283, new_n2284, new_n2285,
    new_n2286, new_n2287, new_n2288, new_n2289, new_n2290, new_n2291,
    new_n2292, new_n2293, new_n2294, new_n2295, new_n2296, new_n2297,
    new_n2298, new_n2299, new_n2300, new_n2301, new_n2302, new_n2303,
    new_n2304, new_n2305, new_n2306, new_n2307, new_n2308, new_n2309,
    new_n2310, new_n2311, new_n2312, new_n2313, new_n2314, new_n2315,
    new_n2316, new_n2317, new_n2318, new_n2319, new_n2320, new_n2321,
    new_n2322, new_n2323, new_n2324, new_n2325, new_n2326, new_n2327,
    new_n2328, new_n2329, new_n2330, new_n2331, new_n2332, new_n2333,
    new_n2334, new_n2335, new_n2336, new_n2337, new_n2338, new_n2339,
    new_n2340, new_n2341, new_n2342, new_n2343, new_n2344, new_n2345,
    new_n2346, new_n2347, new_n2348, new_n2349, new_n2350, new_n2351,
    new_n2352, new_n2353, new_n2354, new_n2355, new_n2356, new_n2357,
    new_n2358, new_n2359, new_n2360, new_n2361, new_n2362, new_n2363,
    new_n2364, new_n2365, new_n2366, new_n2367, new_n2368, new_n2369,
    new_n2370, new_n2371, new_n2372, new_n2373, new_n2374, new_n2375,
    new_n2376, new_n2377, new_n2378, new_n2379, new_n2380, new_n2381,
    new_n2382, new_n2383, new_n2384, new_n2385, new_n2386, new_n2387,
    new_n2388, new_n2389, new_n2390, new_n2391, new_n2392, new_n2393,
    new_n2394, new_n2395, new_n2396, new_n2397, new_n2398, new_n2399,
    new_n2400, new_n2401, new_n2402, new_n2403, new_n2404, new_n2405,
    new_n2406, new_n2407, new_n2408, new_n2409, new_n2410, new_n2411,
    new_n2412, new_n2413, new_n2414, new_n2415, new_n2416, new_n2417,
    new_n2418, new_n2419, new_n2420, new_n2421, new_n2422, new_n2423,
    new_n2424, new_n2425, new_n2426, new_n2427, new_n2428, new_n2429,
    new_n2430, new_n2431, new_n2432, new_n2433, new_n2434, new_n2435,
    new_n2436, new_n2437, new_n2438, new_n2439, new_n2440, new_n2441,
    new_n2442, new_n2443, new_n2444, new_n2445, new_n2446, new_n2447,
    new_n2448, new_n2449, new_n2450, new_n2451, new_n2452, new_n2453,
    new_n2454, new_n2455, new_n2456, new_n2457, new_n2458, new_n2459,
    new_n2460, new_n2461, new_n2462, new_n2463, new_n2464, new_n2465,
    new_n2466, new_n2467, new_n2468, new_n2469, new_n2470, new_n2471,
    new_n2472, new_n2473, new_n2474, new_n2475, new_n2476, new_n2477,
    new_n2478, new_n2479, new_n2480, new_n2481, new_n2482, new_n2483,
    new_n2484, new_n2485, new_n2486, new_n2487, new_n2488, new_n2489,
    new_n2490, new_n2491, new_n2492, new_n2493, new_n2494, new_n2495,
    new_n2496, new_n2497, new_n2498, new_n2499, new_n2500, new_n2501,
    new_n2502, new_n2503, new_n2504, new_n2505, new_n2506, new_n2507,
    new_n2508, new_n2509, new_n2510, new_n2511, new_n2512, new_n2513,
    new_n2514, new_n2515, new_n2516, new_n2517, new_n2518, new_n2519,
    new_n2520, new_n2521, new_n2522, new_n2523, new_n2524, new_n2525,
    new_n2526, new_n2527, new_n2528, new_n2529, new_n2530, new_n2531,
    new_n2532, new_n2533, new_n2534, new_n2535, new_n2536, new_n2537,
    new_n2538, new_n2539, new_n2540, new_n2541, new_n2542, new_n2543,
    new_n2544, new_n2545, new_n2546, new_n2547, new_n2548, new_n2549,
    new_n2550, new_n2551, new_n2552, new_n2553, new_n2554, new_n2555,
    new_n2556, new_n2557, new_n2558, new_n2559, new_n2560, new_n2561,
    new_n2562, new_n2563, new_n2564, new_n2565, new_n2566, new_n2567,
    new_n2568, new_n2569, new_n2570, new_n2571, new_n2572, new_n2573,
    new_n2574, new_n2575, new_n2576, new_n2577, new_n2578, new_n2579,
    new_n2580, new_n2581, new_n2582, new_n2583, new_n2584, new_n2585,
    new_n2586, new_n2587, new_n2588, new_n2589, new_n2590, new_n2591,
    new_n2592, new_n2593, new_n2594, new_n2595, new_n2596, new_n2597,
    new_n2598, new_n2599, new_n2600, new_n2601, new_n2602, new_n2603,
    new_n2604, new_n2605, new_n2606, new_n2607, new_n2608, new_n2609,
    new_n2610, new_n2611, new_n2612, new_n2613, new_n2614, new_n2615,
    new_n2616, new_n2617, new_n2618, new_n2619, new_n2620, new_n2621,
    new_n2622, new_n2623, new_n2624, new_n2625, new_n2626, new_n2627,
    new_n2628, new_n2629, new_n2630, new_n2631, new_n2632, new_n2633,
    new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639,
    new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2645,
    new_n2646, new_n2647, new_n2648, new_n2649, new_n2650, new_n2651,
    new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657,
    new_n2658, new_n2659, new_n2660, new_n2661, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2670, new_n2671, new_n2672, new_n2673, new_n2674, new_n2675,
    new_n2676, new_n2677, new_n2678, new_n2679, new_n2680, new_n2681,
    new_n2682, new_n2683, new_n2684, new_n2685, new_n2686, new_n2687,
    new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693,
    new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699,
    new_n2700, new_n2701, new_n2702, new_n2703, new_n2704, new_n2705,
    new_n2706, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779, new_n2780, new_n2781, new_n2782, new_n2783,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2848, new_n2849,
    new_n2850, new_n2851, new_n2852, new_n2853, new_n2854, new_n2855,
    new_n2856, new_n2857, new_n2858, new_n2859, new_n2860, new_n2861,
    new_n2862, new_n2863, new_n2864, new_n2865, new_n2866, new_n2867,
    new_n2868, new_n2869, new_n2870, new_n2871, new_n2872, new_n2873,
    new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879,
    new_n2880, new_n2881, new_n2882, new_n2883, new_n2884, new_n2885,
    new_n2886, new_n2887, new_n2888, new_n2889, new_n2890, new_n2891,
    new_n2892, new_n2893, new_n2894, new_n2895, new_n2896, new_n2897,
    new_n2898, new_n2899, new_n2900, new_n2901, new_n2902, new_n2903,
    new_n2904, new_n2905, new_n2906, new_n2907, new_n2908, new_n2909,
    new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915,
    new_n2916, new_n2917, new_n2918, new_n2919, new_n2920, new_n2921,
    new_n2922;
  assign new_n513 = n128 & n256;
  assign new_n514 = n384 & n512;
  assign new_n515 = new_n514 ^ new_n513;
  assign new_n516 = n255 ^ n127;
  assign new_n517 = n256 ^ n128;
  assign new_n518 = n254 ^ n126;
  assign new_n519 = n253 ^ n125;
  assign new_n520 = ~n125 & n253;
  assign new_n521 = new_n520 ^ new_n519;
  assign new_n522 = new_n521 ^ n254;
  assign new_n523 = ~new_n518 & ~new_n522;
  assign new_n524 = new_n523 ^ n254;
  assign new_n525 = new_n524 ^ n255;
  assign new_n526 = ~new_n516 & new_n525;
  assign new_n527 = new_n526 ^ n255;
  assign new_n528 = new_n527 ^ n256;
  assign new_n529 = new_n528 ^ n256;
  assign new_n530 = ~n126 & n254;
  assign new_n531 = ~n127 & n255;
  assign new_n532 = ~new_n530 & ~new_n531;
  assign new_n533 = n252 ^ n124;
  assign new_n534 = ~n252 & n124;
  assign new_n535 = new_n534 ^ new_n533;
  assign new_n536 = ~new_n520 & ~new_n535;
  assign new_n537 = new_n532 & new_n536;
  assign new_n538 = n251 ^ n123;
  assign new_n539 = n250 ^ n122;
  assign new_n540 = n249 ^ n121;
  assign new_n541 = n248 ^ n120;
  assign new_n542 = n247 ^ n119;
  assign new_n543 = n246 ^ n118;
  assign new_n544 = n245 ^ n117;
  assign new_n545 = n244 ^ n116;
  assign new_n546 = n243 ^ n115;
  assign new_n547 = n242 ^ n114;
  assign new_n548 = n241 ^ n113;
  assign new_n549 = n240 ^ n112;
  assign new_n550 = n239 ^ n111;
  assign new_n551 = n238 ^ n110;
  assign new_n552 = n237 ^ n109;
  assign new_n553 = n236 ^ n108;
  assign new_n554 = n235 ^ n107;
  assign new_n555 = n234 ^ n106;
  assign new_n556 = n233 ^ n105;
  assign new_n557 = n232 ^ n104;
  assign new_n558 = n231 ^ n103;
  assign new_n559 = n230 ^ n102;
  assign new_n560 = n229 ^ n101;
  assign new_n561 = n228 ^ n100;
  assign new_n562 = n227 ^ n99;
  assign new_n563 = n226 ^ n98;
  assign new_n564 = n225 ^ n97;
  assign new_n565 = n224 ^ n96;
  assign new_n566 = n223 ^ n95;
  assign new_n567 = n222 ^ n94;
  assign new_n568 = n221 ^ n93;
  assign new_n569 = n220 ^ n92;
  assign new_n570 = n219 ^ n91;
  assign new_n571 = n218 ^ n90;
  assign new_n572 = n217 ^ n89;
  assign new_n573 = n216 ^ n88;
  assign new_n574 = n215 ^ n87;
  assign new_n575 = n214 ^ n86;
  assign new_n576 = n213 ^ n85;
  assign new_n577 = n212 ^ n84;
  assign new_n578 = n211 ^ n83;
  assign new_n579 = n210 ^ n82;
  assign new_n580 = n209 ^ n81;
  assign new_n581 = ~n81 & n209;
  assign new_n582 = new_n581 ^ new_n580;
  assign new_n583 = new_n582 ^ n210;
  assign new_n584 = new_n583 ^ n210;
  assign new_n585 = ~n71 & n199;
  assign new_n586 = ~n70 & n198;
  assign new_n587 = ~new_n585 & ~new_n586;
  assign new_n588 = n197 ^ n69;
  assign new_n589 = ~n197 & n69;
  assign new_n590 = new_n589 ^ new_n588;
  assign new_n591 = ~new_n590 & new_n587;
  assign new_n592 = n196 ^ n68;
  assign new_n593 = n195 ^ n67;
  assign new_n594 = n194 ^ n66;
  assign new_n595 = n193 ^ n65;
  assign new_n596 = n192 ^ n64;
  assign new_n597 = ~n192 & n64;
  assign new_n598 = new_n597 ^ new_n596;
  assign new_n599 = new_n598 ^ n193;
  assign new_n600 = new_n599 ^ n193;
  assign new_n601 = ~n63 & n191;
  assign new_n602 = ~n62 & n190;
  assign new_n603 = ~new_n601 & ~new_n602;
  assign new_n604 = n188 ^ n60;
  assign new_n605 = ~n188 & n60;
  assign new_n606 = new_n605 ^ new_n604;
  assign new_n607 = n189 ^ n61;
  assign new_n608 = ~n189 & n61;
  assign new_n609 = new_n608 ^ new_n607;
  assign new_n610 = ~new_n606 & ~new_n609;
  assign new_n611 = new_n603 & new_n610;
  assign new_n612 = n187 ^ n59;
  assign new_n613 = n186 ^ n58;
  assign new_n614 = n185 ^ n57;
  assign new_n615 = n184 ^ n56;
  assign new_n616 = n183 ^ n55;
  assign new_n617 = n182 ^ n54;
  assign new_n618 = n181 ^ n53;
  assign new_n619 = n180 ^ n52;
  assign new_n620 = n179 ^ n51;
  assign new_n621 = n178 ^ n50;
  assign new_n622 = n177 ^ n49;
  assign new_n623 = ~n49 & n177;
  assign new_n624 = new_n623 ^ new_n622;
  assign new_n625 = new_n624 ^ n178;
  assign new_n626 = new_n625 ^ n178;
  assign new_n627 = n167 ^ n39;
  assign new_n628 = n166 ^ n38;
  assign new_n629 = n165 ^ n37;
  assign new_n630 = n164 ^ n36;
  assign new_n631 = n163 ^ n35;
  assign new_n632 = n162 ^ n34;
  assign new_n633 = n161 ^ n33;
  assign new_n634 = n160 ^ n32;
  assign new_n635 = n159 ^ n31;
  assign new_n636 = n158 ^ n30;
  assign new_n637 = n157 ^ n29;
  assign new_n638 = n156 ^ n28;
  assign new_n639 = n155 ^ n27;
  assign new_n640 = n154 ^ n26;
  assign new_n641 = n153 ^ n25;
  assign new_n642 = n152 ^ n24;
  assign new_n643 = n151 ^ n23;
  assign new_n644 = n150 ^ n22;
  assign new_n645 = n149 ^ n21;
  assign new_n646 = n148 ^ n20;
  assign new_n647 = n147 ^ n19;
  assign new_n648 = n146 ^ n18;
  assign new_n649 = n145 ^ n17;
  assign new_n650 = n144 ^ n16;
  assign new_n651 = n143 ^ n15;
  assign new_n652 = n142 ^ n14;
  assign new_n653 = n141 ^ n13;
  assign new_n654 = n140 ^ n12;
  assign new_n655 = n139 ^ n11;
  assign new_n656 = n138 ^ n10;
  assign new_n657 = n137 ^ n9;
  assign new_n658 = n136 ^ n8;
  assign new_n659 = n135 ^ n7;
  assign new_n660 = n134 ^ n6;
  assign new_n661 = n133 ^ n5;
  assign new_n662 = n132 ^ n4;
  assign new_n663 = n131 ^ n3;
  assign new_n664 = n130 ^ n2;
  assign new_n665 = ~n129 & n1;
  assign new_n666 = new_n665 ^ n130;
  assign new_n667 = ~new_n664 & ~new_n666;
  assign new_n668 = new_n667 ^ n130;
  assign new_n669 = new_n668 ^ n131;
  assign new_n670 = ~new_n663 & new_n669;
  assign new_n671 = new_n670 ^ n131;
  assign new_n672 = new_n671 ^ n132;
  assign new_n673 = ~new_n662 & new_n672;
  assign new_n674 = new_n673 ^ n132;
  assign new_n675 = new_n674 ^ n133;
  assign new_n676 = ~new_n661 & ~new_n675;
  assign new_n677 = new_n676 ^ n5;
  assign new_n678 = new_n677 ^ n134;
  assign new_n679 = ~new_n660 & new_n678;
  assign new_n680 = new_n679 ^ n6;
  assign new_n681 = new_n680 ^ n135;
  assign new_n682 = ~new_n659 & ~new_n681;
  assign new_n683 = new_n682 ^ n135;
  assign new_n684 = new_n683 ^ n136;
  assign new_n685 = ~new_n658 & ~new_n684;
  assign new_n686 = new_n685 ^ n8;
  assign new_n687 = new_n686 ^ n137;
  assign new_n688 = ~new_n657 & new_n687;
  assign new_n689 = new_n688 ^ n9;
  assign new_n690 = new_n689 ^ n138;
  assign new_n691 = ~new_n656 & ~new_n690;
  assign new_n692 = new_n691 ^ n138;
  assign new_n693 = new_n692 ^ n139;
  assign new_n694 = ~new_n655 & ~new_n693;
  assign new_n695 = new_n694 ^ n11;
  assign new_n696 = new_n695 ^ n140;
  assign new_n697 = ~new_n654 & new_n696;
  assign new_n698 = new_n697 ^ n12;
  assign new_n699 = new_n698 ^ n141;
  assign new_n700 = ~new_n653 & new_n699;
  assign new_n701 = new_n700 ^ n13;
  assign new_n702 = new_n701 ^ n142;
  assign new_n703 = ~new_n652 & new_n702;
  assign new_n704 = new_n703 ^ n14;
  assign new_n705 = new_n704 ^ n143;
  assign new_n706 = ~new_n651 & new_n705;
  assign new_n707 = new_n706 ^ n15;
  assign new_n708 = new_n707 ^ n144;
  assign new_n709 = ~new_n650 & new_n708;
  assign new_n710 = new_n709 ^ n16;
  assign new_n711 = new_n710 ^ n145;
  assign new_n712 = ~new_n649 & ~new_n711;
  assign new_n713 = new_n712 ^ n145;
  assign new_n714 = new_n713 ^ n146;
  assign new_n715 = ~new_n648 & ~new_n714;
  assign new_n716 = new_n715 ^ n18;
  assign new_n717 = new_n716 ^ n147;
  assign new_n718 = ~new_n647 & new_n717;
  assign new_n719 = new_n718 ^ n19;
  assign new_n720 = new_n719 ^ n148;
  assign new_n721 = ~new_n646 & ~new_n720;
  assign new_n722 = new_n721 ^ n148;
  assign new_n723 = new_n722 ^ n149;
  assign new_n724 = ~new_n645 & new_n723;
  assign new_n725 = new_n724 ^ n149;
  assign new_n726 = new_n725 ^ n150;
  assign new_n727 = ~new_n644 & new_n726;
  assign new_n728 = new_n727 ^ n150;
  assign new_n729 = new_n728 ^ n151;
  assign new_n730 = ~new_n643 & new_n729;
  assign new_n731 = new_n730 ^ n151;
  assign new_n732 = new_n731 ^ n152;
  assign new_n733 = ~new_n642 & new_n732;
  assign new_n734 = new_n733 ^ n152;
  assign new_n735 = new_n734 ^ n153;
  assign new_n736 = ~new_n641 & new_n735;
  assign new_n737 = new_n736 ^ n153;
  assign new_n738 = new_n737 ^ n154;
  assign new_n739 = ~new_n640 & ~new_n738;
  assign new_n740 = new_n739 ^ n26;
  assign new_n741 = new_n740 ^ n155;
  assign new_n742 = ~new_n639 & new_n741;
  assign new_n743 = new_n742 ^ n27;
  assign new_n744 = new_n743 ^ n156;
  assign new_n745 = ~new_n638 & ~new_n744;
  assign new_n746 = new_n745 ^ n156;
  assign new_n747 = new_n746 ^ n157;
  assign new_n748 = ~new_n637 & ~new_n747;
  assign new_n749 = new_n748 ^ n29;
  assign new_n750 = new_n749 ^ n158;
  assign new_n751 = ~new_n636 & new_n750;
  assign new_n752 = new_n751 ^ n30;
  assign new_n753 = new_n752 ^ n159;
  assign new_n754 = ~new_n635 & ~new_n753;
  assign new_n755 = new_n754 ^ n159;
  assign new_n756 = new_n755 ^ n160;
  assign new_n757 = ~new_n634 & ~new_n756;
  assign new_n758 = new_n757 ^ n32;
  assign new_n759 = new_n758 ^ n161;
  assign new_n760 = ~new_n633 & new_n759;
  assign new_n761 = new_n760 ^ n33;
  assign new_n762 = new_n761 ^ n162;
  assign new_n763 = ~new_n632 & ~new_n762;
  assign new_n764 = new_n763 ^ n162;
  assign new_n765 = new_n764 ^ n163;
  assign new_n766 = ~new_n631 & new_n765;
  assign new_n767 = new_n766 ^ n163;
  assign new_n768 = new_n767 ^ n164;
  assign new_n769 = ~new_n630 & new_n768;
  assign new_n770 = new_n769 ^ n164;
  assign new_n771 = new_n770 ^ n165;
  assign new_n772 = ~new_n629 & new_n771;
  assign new_n773 = new_n772 ^ n165;
  assign new_n774 = new_n773 ^ n166;
  assign new_n775 = ~new_n628 & ~new_n774;
  assign new_n776 = new_n775 ^ n38;
  assign new_n777 = new_n776 ^ n167;
  assign new_n778 = ~new_n627 & new_n777;
  assign new_n779 = new_n778 ^ n39;
  assign new_n780 = n168 ^ n40;
  assign new_n781 = ~n40 & n168;
  assign new_n782 = new_n781 ^ new_n780;
  assign new_n783 = ~new_n779 & ~new_n782;
  assign new_n784 = ~n42 & n170;
  assign new_n785 = ~n43 & n171;
  assign new_n786 = ~new_n784 & ~new_n785;
  assign new_n787 = n169 ^ n41;
  assign new_n788 = ~n169 & n41;
  assign new_n789 = new_n788 ^ new_n787;
  assign new_n790 = ~new_n781 & ~new_n789;
  assign new_n791 = new_n786 & new_n790;
  assign new_n792 = ~new_n783 & new_n791;
  assign new_n793 = n171 ^ n43;
  assign new_n794 = n170 ^ n42;
  assign new_n795 = new_n788 ^ n170;
  assign new_n796 = ~new_n794 & ~new_n795;
  assign new_n797 = new_n796 ^ n170;
  assign new_n798 = new_n797 ^ n171;
  assign new_n799 = ~new_n793 & new_n798;
  assign new_n800 = new_n799 ^ n171;
  assign new_n801 = n172 ^ n44;
  assign new_n802 = ~n44 & n172;
  assign new_n803 = new_n802 ^ new_n801;
  assign new_n804 = ~new_n803 & new_n800;
  assign new_n805 = ~new_n792 & new_n804;
  assign new_n806 = ~n47 & n175;
  assign new_n807 = ~n46 & n174;
  assign new_n808 = ~new_n806 & ~new_n807;
  assign new_n809 = n173 ^ n45;
  assign new_n810 = ~n173 & n45;
  assign new_n811 = new_n810 ^ new_n809;
  assign new_n812 = ~new_n802 & ~new_n811;
  assign new_n813 = new_n808 & new_n812;
  assign new_n814 = ~new_n805 & new_n813;
  assign new_n815 = n175 ^ n47;
  assign new_n816 = n174 ^ n46;
  assign new_n817 = new_n810 ^ n174;
  assign new_n818 = ~new_n816 & ~new_n817;
  assign new_n819 = new_n818 ^ n174;
  assign new_n820 = new_n819 ^ n175;
  assign new_n821 = ~new_n815 & new_n820;
  assign new_n822 = new_n821 ^ n175;
  assign new_n823 = n176 ^ n48;
  assign new_n824 = ~n48 & n176;
  assign new_n825 = new_n824 ^ new_n823;
  assign new_n826 = ~new_n825 & new_n822;
  assign new_n827 = ~new_n814 & new_n826;
  assign new_n828 = ~new_n623 & ~new_n824;
  assign new_n829 = ~new_n827 & new_n828;
  assign new_n830 = new_n829 ^ n178;
  assign new_n831 = new_n830 ^ n178;
  assign new_n832 = ~new_n626 & ~new_n831;
  assign new_n833 = new_n832 ^ n178;
  assign new_n834 = ~new_n621 & ~new_n833;
  assign new_n835 = new_n834 ^ n50;
  assign new_n836 = new_n835 ^ n179;
  assign new_n837 = ~new_n620 & ~new_n836;
  assign new_n838 = new_n837 ^ n179;
  assign new_n839 = new_n838 ^ n180;
  assign new_n840 = ~new_n619 & new_n839;
  assign new_n841 = new_n840 ^ n180;
  assign new_n842 = new_n841 ^ n181;
  assign new_n843 = ~new_n618 & new_n842;
  assign new_n844 = new_n843 ^ n181;
  assign new_n845 = new_n844 ^ n182;
  assign new_n846 = ~new_n617 & new_n845;
  assign new_n847 = new_n846 ^ n182;
  assign new_n848 = new_n847 ^ n183;
  assign new_n849 = ~new_n616 & new_n848;
  assign new_n850 = new_n849 ^ n183;
  assign new_n851 = new_n850 ^ n184;
  assign new_n852 = ~new_n615 & ~new_n851;
  assign new_n853 = new_n852 ^ n56;
  assign new_n854 = new_n853 ^ n185;
  assign new_n855 = ~new_n614 & new_n854;
  assign new_n856 = new_n855 ^ n57;
  assign new_n857 = new_n856 ^ n186;
  assign new_n858 = ~new_n613 & ~new_n857;
  assign new_n859 = new_n858 ^ n186;
  assign new_n860 = new_n859 ^ n187;
  assign new_n861 = ~new_n612 & new_n860;
  assign new_n862 = new_n861 ^ n187;
  assign new_n863 = ~new_n605 & new_n862;
  assign new_n864 = ~new_n863 & new_n611;
  assign new_n865 = n191 ^ n63;
  assign new_n866 = n190 ^ n62;
  assign new_n867 = new_n608 ^ n190;
  assign new_n868 = ~new_n866 & ~new_n867;
  assign new_n869 = new_n868 ^ n190;
  assign new_n870 = new_n869 ^ n191;
  assign new_n871 = ~new_n865 & new_n870;
  assign new_n872 = new_n871 ^ n191;
  assign new_n873 = ~new_n597 & new_n872;
  assign new_n874 = ~new_n864 & new_n873;
  assign new_n875 = new_n874 ^ n193;
  assign new_n876 = new_n875 ^ n193;
  assign new_n877 = ~new_n600 & ~new_n876;
  assign new_n878 = new_n877 ^ n193;
  assign new_n879 = ~new_n595 & new_n878;
  assign new_n880 = new_n879 ^ n65;
  assign new_n881 = new_n880 ^ n194;
  assign new_n882 = ~new_n594 & ~new_n881;
  assign new_n883 = new_n882 ^ n194;
  assign new_n884 = new_n883 ^ n195;
  assign new_n885 = ~new_n593 & ~new_n884;
  assign new_n886 = new_n885 ^ n67;
  assign new_n887 = new_n886 ^ n196;
  assign new_n888 = ~new_n592 & new_n887;
  assign new_n889 = new_n888 ^ n68;
  assign new_n890 = new_n591 & new_n889;
  assign new_n891 = n199 ^ n71;
  assign new_n892 = n198 ^ n70;
  assign new_n893 = new_n589 ^ n198;
  assign new_n894 = ~new_n892 & ~new_n893;
  assign new_n895 = new_n894 ^ n198;
  assign new_n896 = new_n895 ^ n199;
  assign new_n897 = ~new_n891 & new_n896;
  assign new_n898 = new_n897 ^ n199;
  assign new_n899 = n200 ^ n72;
  assign new_n900 = ~n72 & n200;
  assign new_n901 = new_n900 ^ new_n899;
  assign new_n902 = ~new_n901 & new_n898;
  assign new_n903 = ~new_n890 & new_n902;
  assign new_n904 = n201 ^ n73;
  assign new_n905 = ~n201 & n73;
  assign new_n906 = new_n905 ^ new_n904;
  assign new_n907 = ~new_n900 & ~new_n906;
  assign new_n908 = ~new_n903 & new_n907;
  assign new_n909 = n202 ^ n74;
  assign new_n910 = ~n74 & n202;
  assign new_n911 = new_n910 ^ new_n909;
  assign new_n912 = ~new_n905 & ~new_n911;
  assign new_n913 = ~new_n908 & new_n912;
  assign new_n914 = n203 ^ n75;
  assign new_n915 = ~n203 & n75;
  assign new_n916 = new_n915 ^ new_n914;
  assign new_n917 = ~new_n910 & ~new_n916;
  assign new_n918 = ~new_n913 & new_n917;
  assign new_n919 = n204 ^ n76;
  assign new_n920 = ~n76 & n204;
  assign new_n921 = new_n920 ^ new_n919;
  assign new_n922 = ~new_n915 & ~new_n921;
  assign new_n923 = ~new_n918 & new_n922;
  assign new_n924 = n205 ^ n77;
  assign new_n925 = ~n205 & n77;
  assign new_n926 = new_n925 ^ new_n924;
  assign new_n927 = ~new_n920 & ~new_n926;
  assign new_n928 = ~new_n923 & new_n927;
  assign new_n929 = n206 ^ n78;
  assign new_n930 = ~n78 & n206;
  assign new_n931 = new_n930 ^ new_n929;
  assign new_n932 = ~new_n925 & ~new_n931;
  assign new_n933 = ~new_n928 & new_n932;
  assign new_n934 = n207 ^ n79;
  assign new_n935 = ~n207 & n79;
  assign new_n936 = new_n935 ^ new_n934;
  assign new_n937 = ~new_n930 & ~new_n936;
  assign new_n938 = ~new_n933 & new_n937;
  assign new_n939 = n208 ^ n80;
  assign new_n940 = ~n80 & n208;
  assign new_n941 = new_n940 ^ new_n939;
  assign new_n942 = ~new_n935 & ~new_n941;
  assign new_n943 = ~new_n938 & new_n942;
  assign new_n944 = ~new_n581 & ~new_n940;
  assign new_n945 = ~new_n943 & new_n944;
  assign new_n946 = new_n945 ^ n210;
  assign new_n947 = new_n946 ^ n210;
  assign new_n948 = ~new_n584 & ~new_n947;
  assign new_n949 = new_n948 ^ n210;
  assign new_n950 = ~new_n579 & ~new_n949;
  assign new_n951 = new_n950 ^ n82;
  assign new_n952 = new_n951 ^ n211;
  assign new_n953 = ~new_n578 & ~new_n952;
  assign new_n954 = new_n953 ^ n211;
  assign new_n955 = new_n954 ^ n212;
  assign new_n956 = ~new_n577 & new_n955;
  assign new_n957 = new_n956 ^ n212;
  assign new_n958 = new_n957 ^ n213;
  assign new_n959 = ~new_n576 & new_n958;
  assign new_n960 = new_n959 ^ n213;
  assign new_n961 = new_n960 ^ n214;
  assign new_n962 = ~new_n575 & new_n961;
  assign new_n963 = new_n962 ^ n214;
  assign new_n964 = new_n963 ^ n215;
  assign new_n965 = ~new_n574 & new_n964;
  assign new_n966 = new_n965 ^ n215;
  assign new_n967 = new_n966 ^ n216;
  assign new_n968 = ~new_n573 & new_n967;
  assign new_n969 = new_n968 ^ n216;
  assign new_n970 = new_n969 ^ n217;
  assign new_n971 = ~new_n572 & new_n970;
  assign new_n972 = new_n971 ^ n217;
  assign new_n973 = new_n972 ^ n218;
  assign new_n974 = ~new_n571 & ~new_n973;
  assign new_n975 = new_n974 ^ n90;
  assign new_n976 = new_n975 ^ n219;
  assign new_n977 = ~new_n570 & new_n976;
  assign new_n978 = new_n977 ^ n91;
  assign new_n979 = new_n978 ^ n220;
  assign new_n980 = ~new_n569 & new_n979;
  assign new_n981 = new_n980 ^ n92;
  assign new_n982 = new_n981 ^ n221;
  assign new_n983 = ~new_n568 & new_n982;
  assign new_n984 = new_n983 ^ n93;
  assign new_n985 = new_n984 ^ n222;
  assign new_n986 = ~new_n567 & new_n985;
  assign new_n987 = new_n986 ^ n94;
  assign new_n988 = new_n987 ^ n223;
  assign new_n989 = ~new_n566 & new_n988;
  assign new_n990 = new_n989 ^ n95;
  assign new_n991 = new_n990 ^ n224;
  assign new_n992 = ~new_n565 & ~new_n991;
  assign new_n993 = new_n992 ^ n224;
  assign new_n994 = new_n993 ^ n225;
  assign new_n995 = ~new_n564 & ~new_n994;
  assign new_n996 = new_n995 ^ n97;
  assign new_n997 = new_n996 ^ n226;
  assign new_n998 = ~new_n563 & new_n997;
  assign new_n999 = new_n998 ^ n98;
  assign new_n1000 = new_n999 ^ n227;
  assign new_n1001 = ~new_n562 & ~new_n1000;
  assign new_n1002 = new_n1001 ^ n227;
  assign new_n1003 = new_n1002 ^ n228;
  assign new_n1004 = ~new_n561 & new_n1003;
  assign new_n1005 = new_n1004 ^ n228;
  assign new_n1006 = new_n1005 ^ n229;
  assign new_n1007 = ~new_n560 & ~new_n1006;
  assign new_n1008 = new_n1007 ^ n101;
  assign new_n1009 = new_n1008 ^ n230;
  assign new_n1010 = ~new_n559 & new_n1009;
  assign new_n1011 = new_n1010 ^ n102;
  assign new_n1012 = new_n1011 ^ n231;
  assign new_n1013 = ~new_n558 & ~new_n1012;
  assign new_n1014 = new_n1013 ^ n231;
  assign new_n1015 = new_n1014 ^ n232;
  assign new_n1016 = ~new_n557 & new_n1015;
  assign new_n1017 = new_n1016 ^ n232;
  assign new_n1018 = new_n1017 ^ n233;
  assign new_n1019 = ~new_n556 & ~new_n1018;
  assign new_n1020 = new_n1019 ^ n105;
  assign new_n1021 = new_n1020 ^ n234;
  assign new_n1022 = ~new_n555 & new_n1021;
  assign new_n1023 = new_n1022 ^ n106;
  assign new_n1024 = new_n1023 ^ n235;
  assign new_n1025 = ~new_n554 & ~new_n1024;
  assign new_n1026 = new_n1025 ^ n235;
  assign new_n1027 = new_n1026 ^ n236;
  assign new_n1028 = ~new_n553 & new_n1027;
  assign new_n1029 = new_n1028 ^ n236;
  assign new_n1030 = new_n1029 ^ n237;
  assign new_n1031 = ~new_n552 & ~new_n1030;
  assign new_n1032 = new_n1031 ^ n109;
  assign new_n1033 = new_n1032 ^ n238;
  assign new_n1034 = ~new_n551 & new_n1033;
  assign new_n1035 = new_n1034 ^ n110;
  assign new_n1036 = new_n1035 ^ n239;
  assign new_n1037 = ~new_n550 & ~new_n1036;
  assign new_n1038 = new_n1037 ^ n239;
  assign new_n1039 = new_n1038 ^ n240;
  assign new_n1040 = ~new_n549 & new_n1039;
  assign new_n1041 = new_n1040 ^ n240;
  assign new_n1042 = new_n1041 ^ n241;
  assign new_n1043 = ~new_n548 & ~new_n1042;
  assign new_n1044 = new_n1043 ^ n113;
  assign new_n1045 = new_n1044 ^ n242;
  assign new_n1046 = ~new_n547 & new_n1045;
  assign new_n1047 = new_n1046 ^ n114;
  assign new_n1048 = new_n1047 ^ n243;
  assign new_n1049 = ~new_n546 & ~new_n1048;
  assign new_n1050 = new_n1049 ^ n243;
  assign new_n1051 = new_n1050 ^ n244;
  assign new_n1052 = ~new_n545 & ~new_n1051;
  assign new_n1053 = new_n1052 ^ n116;
  assign new_n1054 = new_n1053 ^ n245;
  assign new_n1055 = ~new_n544 & new_n1054;
  assign new_n1056 = new_n1055 ^ n117;
  assign new_n1057 = new_n1056 ^ n246;
  assign new_n1058 = ~new_n543 & ~new_n1057;
  assign new_n1059 = new_n1058 ^ n246;
  assign new_n1060 = new_n1059 ^ n247;
  assign new_n1061 = ~new_n542 & ~new_n1060;
  assign new_n1062 = new_n1061 ^ n119;
  assign new_n1063 = new_n1062 ^ n248;
  assign new_n1064 = ~new_n541 & new_n1063;
  assign new_n1065 = new_n1064 ^ n120;
  assign new_n1066 = new_n1065 ^ n249;
  assign new_n1067 = ~new_n540 & new_n1066;
  assign new_n1068 = new_n1067 ^ n121;
  assign new_n1069 = new_n1068 ^ n250;
  assign new_n1070 = ~new_n539 & new_n1069;
  assign new_n1071 = new_n1070 ^ n122;
  assign new_n1072 = new_n1071 ^ n251;
  assign new_n1073 = ~new_n538 & ~new_n1072;
  assign new_n1074 = new_n1073 ^ n251;
  assign new_n1075 = ~new_n534 & new_n1074;
  assign new_n1076 = ~new_n1075 & new_n537;
  assign new_n1077 = new_n1076 ^ n256;
  assign new_n1078 = new_n1077 ^ n256;
  assign new_n1079 = ~new_n1078 & new_n529;
  assign new_n1080 = new_n1079 ^ n256;
  assign new_n1081 = ~new_n517 & new_n1080;
  assign new_n1082 = new_n1081 ^ n128;
  assign new_n1083 = new_n516 & new_n1082;
  assign new_n1084 = new_n1083 ^ n127;
  assign new_n1085 = n511 ^ n383;
  assign new_n1086 = n512 ^ n384;
  assign new_n1087 = n510 ^ n382;
  assign new_n1088 = n509 ^ n381;
  assign new_n1089 = ~n381 & n509;
  assign new_n1090 = new_n1089 ^ new_n1088;
  assign new_n1091 = new_n1090 ^ n510;
  assign new_n1092 = ~new_n1087 & ~new_n1091;
  assign new_n1093 = new_n1092 ^ n510;
  assign new_n1094 = new_n1093 ^ n511;
  assign new_n1095 = ~new_n1085 & new_n1094;
  assign new_n1096 = new_n1095 ^ n511;
  assign new_n1097 = new_n1096 ^ n512;
  assign new_n1098 = new_n1097 ^ n512;
  assign new_n1099 = ~n382 & n510;
  assign new_n1100 = ~n383 & n511;
  assign new_n1101 = ~new_n1099 & ~new_n1100;
  assign new_n1102 = n508 ^ n380;
  assign new_n1103 = ~n508 & n380;
  assign new_n1104 = new_n1103 ^ new_n1102;
  assign new_n1105 = ~new_n1089 & ~new_n1104;
  assign new_n1106 = new_n1101 & new_n1105;
  assign new_n1107 = n507 ^ n379;
  assign new_n1108 = n506 ^ n378;
  assign new_n1109 = n505 ^ n377;
  assign new_n1110 = n504 ^ n376;
  assign new_n1111 = n503 ^ n375;
  assign new_n1112 = n502 ^ n374;
  assign new_n1113 = n501 ^ n373;
  assign new_n1114 = n500 ^ n372;
  assign new_n1115 = n499 ^ n371;
  assign new_n1116 = n498 ^ n370;
  assign new_n1117 = n497 ^ n369;
  assign new_n1118 = n496 ^ n368;
  assign new_n1119 = n495 ^ n367;
  assign new_n1120 = n494 ^ n366;
  assign new_n1121 = n493 ^ n365;
  assign new_n1122 = n492 ^ n364;
  assign new_n1123 = n491 ^ n363;
  assign new_n1124 = n490 ^ n362;
  assign new_n1125 = n489 ^ n361;
  assign new_n1126 = n488 ^ n360;
  assign new_n1127 = n487 ^ n359;
  assign new_n1128 = n486 ^ n358;
  assign new_n1129 = n485 ^ n357;
  assign new_n1130 = n484 ^ n356;
  assign new_n1131 = n483 ^ n355;
  assign new_n1132 = n482 ^ n354;
  assign new_n1133 = n481 ^ n353;
  assign new_n1134 = n480 ^ n352;
  assign new_n1135 = n479 ^ n351;
  assign new_n1136 = n478 ^ n350;
  assign new_n1137 = n477 ^ n349;
  assign new_n1138 = n476 ^ n348;
  assign new_n1139 = n475 ^ n347;
  assign new_n1140 = n474 ^ n346;
  assign new_n1141 = n473 ^ n345;
  assign new_n1142 = n472 ^ n344;
  assign new_n1143 = n471 ^ n343;
  assign new_n1144 = n470 ^ n342;
  assign new_n1145 = n469 ^ n341;
  assign new_n1146 = n468 ^ n340;
  assign new_n1147 = n467 ^ n339;
  assign new_n1148 = n466 ^ n338;
  assign new_n1149 = n465 ^ n337;
  assign new_n1150 = n464 ^ n336;
  assign new_n1151 = n463 ^ n335;
  assign new_n1152 = n462 ^ n334;
  assign new_n1153 = n461 ^ n333;
  assign new_n1154 = n460 ^ n332;
  assign new_n1155 = n459 ^ n331;
  assign new_n1156 = n458 ^ n330;
  assign new_n1157 = n457 ^ n329;
  assign new_n1158 = n456 ^ n328;
  assign new_n1159 = ~n456 & n328;
  assign new_n1160 = new_n1159 ^ new_n1158;
  assign new_n1161 = new_n1160 ^ n457;
  assign new_n1162 = new_n1161 ^ n457;
  assign new_n1163 = ~n326 & n454;
  assign new_n1164 = ~n327 & n455;
  assign new_n1165 = ~new_n1163 & ~new_n1164;
  assign new_n1166 = n452 ^ n324;
  assign new_n1167 = ~n452 & n324;
  assign new_n1168 = new_n1167 ^ new_n1166;
  assign new_n1169 = n453 ^ n325;
  assign new_n1170 = ~n453 & n325;
  assign new_n1171 = new_n1170 ^ new_n1169;
  assign new_n1172 = ~new_n1168 & ~new_n1171;
  assign new_n1173 = new_n1165 & new_n1172;
  assign new_n1174 = n451 ^ n323;
  assign new_n1175 = n450 ^ n322;
  assign new_n1176 = n449 ^ n321;
  assign new_n1177 = ~n449 & n321;
  assign new_n1178 = new_n1177 ^ new_n1176;
  assign new_n1179 = new_n1178 ^ n450;
  assign new_n1180 = new_n1179 ^ n450;
  assign new_n1181 = n443 ^ n315;
  assign new_n1182 = n442 ^ n314;
  assign new_n1183 = n441 ^ n313;
  assign new_n1184 = n440 ^ n312;
  assign new_n1185 = n439 ^ n311;
  assign new_n1186 = n438 ^ n310;
  assign new_n1187 = n437 ^ n309;
  assign new_n1188 = n436 ^ n308;
  assign new_n1189 = ~n436 & n308;
  assign new_n1190 = new_n1189 ^ new_n1188;
  assign new_n1191 = new_n1190 ^ n437;
  assign new_n1192 = new_n1191 ^ n437;
  assign new_n1193 = ~n298 & n426;
  assign new_n1194 = ~n299 & n427;
  assign new_n1195 = ~new_n1193 & ~new_n1194;
  assign new_n1196 = n424 ^ n296;
  assign new_n1197 = ~n424 & n296;
  assign new_n1198 = new_n1197 ^ new_n1196;
  assign new_n1199 = n425 ^ n297;
  assign new_n1200 = ~n425 & n297;
  assign new_n1201 = new_n1200 ^ new_n1199;
  assign new_n1202 = ~new_n1198 & ~new_n1201;
  assign new_n1203 = new_n1195 & new_n1202;
  assign new_n1204 = n423 ^ n295;
  assign new_n1205 = n422 ^ n294;
  assign new_n1206 = n421 ^ n293;
  assign new_n1207 = n420 ^ n292;
  assign new_n1208 = n419 ^ n291;
  assign new_n1209 = n418 ^ n290;
  assign new_n1210 = n417 ^ n289;
  assign new_n1211 = n416 ^ n288;
  assign new_n1212 = n415 ^ n287;
  assign new_n1213 = n414 ^ n286;
  assign new_n1214 = n413 ^ n285;
  assign new_n1215 = n412 ^ n284;
  assign new_n1216 = n411 ^ n283;
  assign new_n1217 = n410 ^ n282;
  assign new_n1218 = n409 ^ n281;
  assign new_n1219 = n408 ^ n280;
  assign new_n1220 = n407 ^ n279;
  assign new_n1221 = n406 ^ n278;
  assign new_n1222 = n405 ^ n277;
  assign new_n1223 = n404 ^ n276;
  assign new_n1224 = n403 ^ n275;
  assign new_n1225 = n402 ^ n274;
  assign new_n1226 = n401 ^ n273;
  assign new_n1227 = n400 ^ n272;
  assign new_n1228 = n399 ^ n271;
  assign new_n1229 = n398 ^ n270;
  assign new_n1230 = n397 ^ n269;
  assign new_n1231 = n396 ^ n268;
  assign new_n1232 = n395 ^ n267;
  assign new_n1233 = n394 ^ n266;
  assign new_n1234 = n393 ^ n265;
  assign new_n1235 = n392 ^ n264;
  assign new_n1236 = n391 ^ n263;
  assign new_n1237 = n390 ^ n262;
  assign new_n1238 = n389 ^ n261;
  assign new_n1239 = n388 ^ n260;
  assign new_n1240 = n387 ^ n259;
  assign new_n1241 = n386 ^ n258;
  assign new_n1242 = ~n385 & n257;
  assign new_n1243 = new_n1242 ^ n386;
  assign new_n1244 = ~new_n1241 & ~new_n1243;
  assign new_n1245 = new_n1244 ^ n386;
  assign new_n1246 = new_n1245 ^ n387;
  assign new_n1247 = ~new_n1240 & new_n1246;
  assign new_n1248 = new_n1247 ^ n387;
  assign new_n1249 = new_n1248 ^ n388;
  assign new_n1250 = ~new_n1239 & ~new_n1249;
  assign new_n1251 = new_n1250 ^ n260;
  assign new_n1252 = new_n1251 ^ n389;
  assign new_n1253 = ~new_n1238 & new_n1252;
  assign new_n1254 = new_n1253 ^ n261;
  assign new_n1255 = new_n1254 ^ n390;
  assign new_n1256 = ~new_n1237 & ~new_n1255;
  assign new_n1257 = new_n1256 ^ n390;
  assign new_n1258 = new_n1257 ^ n391;
  assign new_n1259 = ~new_n1236 & new_n1258;
  assign new_n1260 = new_n1259 ^ n391;
  assign new_n1261 = new_n1260 ^ n392;
  assign new_n1262 = ~new_n1235 & new_n1261;
  assign new_n1263 = new_n1262 ^ n392;
  assign new_n1264 = new_n1263 ^ n393;
  assign new_n1265 = ~new_n1234 & new_n1264;
  assign new_n1266 = new_n1265 ^ n393;
  assign new_n1267 = new_n1266 ^ n394;
  assign new_n1268 = ~new_n1233 & new_n1267;
  assign new_n1269 = new_n1268 ^ n394;
  assign new_n1270 = new_n1269 ^ n395;
  assign new_n1271 = ~new_n1232 & ~new_n1270;
  assign new_n1272 = new_n1271 ^ n267;
  assign new_n1273 = new_n1272 ^ n396;
  assign new_n1274 = ~new_n1231 & new_n1273;
  assign new_n1275 = new_n1274 ^ n268;
  assign new_n1276 = new_n1275 ^ n397;
  assign new_n1277 = ~new_n1230 & new_n1276;
  assign new_n1278 = new_n1277 ^ n269;
  assign new_n1279 = new_n1278 ^ n398;
  assign new_n1280 = ~new_n1229 & new_n1279;
  assign new_n1281 = new_n1280 ^ n270;
  assign new_n1282 = new_n1281 ^ n399;
  assign new_n1283 = ~new_n1228 & new_n1282;
  assign new_n1284 = new_n1283 ^ n271;
  assign new_n1285 = new_n1284 ^ n400;
  assign new_n1286 = ~new_n1227 & new_n1285;
  assign new_n1287 = new_n1286 ^ n272;
  assign new_n1288 = new_n1287 ^ n401;
  assign new_n1289 = ~new_n1226 & new_n1288;
  assign new_n1290 = new_n1289 ^ n273;
  assign new_n1291 = new_n1290 ^ n402;
  assign new_n1292 = ~new_n1225 & new_n1291;
  assign new_n1293 = new_n1292 ^ n274;
  assign new_n1294 = new_n1293 ^ n403;
  assign new_n1295 = ~new_n1224 & ~new_n1294;
  assign new_n1296 = new_n1295 ^ n403;
  assign new_n1297 = new_n1296 ^ n404;
  assign new_n1298 = ~new_n1223 & ~new_n1297;
  assign new_n1299 = new_n1298 ^ n276;
  assign new_n1300 = new_n1299 ^ n405;
  assign new_n1301 = ~new_n1222 & new_n1300;
  assign new_n1302 = new_n1301 ^ n277;
  assign new_n1303 = new_n1302 ^ n406;
  assign new_n1304 = ~new_n1221 & ~new_n1303;
  assign new_n1305 = new_n1304 ^ n406;
  assign new_n1306 = new_n1305 ^ n407;
  assign new_n1307 = ~new_n1220 & new_n1306;
  assign new_n1308 = new_n1307 ^ n407;
  assign new_n1309 = new_n1308 ^ n408;
  assign new_n1310 = ~new_n1219 & new_n1309;
  assign new_n1311 = new_n1310 ^ n408;
  assign new_n1312 = new_n1311 ^ n409;
  assign new_n1313 = ~new_n1218 & new_n1312;
  assign new_n1314 = new_n1313 ^ n409;
  assign new_n1315 = new_n1314 ^ n410;
  assign new_n1316 = ~new_n1217 & ~new_n1315;
  assign new_n1317 = new_n1316 ^ n282;
  assign new_n1318 = new_n1317 ^ n411;
  assign new_n1319 = ~new_n1216 & new_n1318;
  assign new_n1320 = new_n1319 ^ n283;
  assign new_n1321 = new_n1320 ^ n412;
  assign new_n1322 = ~new_n1215 & ~new_n1321;
  assign new_n1323 = new_n1322 ^ n412;
  assign new_n1324 = new_n1323 ^ n413;
  assign new_n1325 = ~new_n1214 & new_n1324;
  assign new_n1326 = new_n1325 ^ n413;
  assign new_n1327 = new_n1326 ^ n414;
  assign new_n1328 = ~new_n1213 & ~new_n1327;
  assign new_n1329 = new_n1328 ^ n286;
  assign new_n1330 = new_n1329 ^ n415;
  assign new_n1331 = ~new_n1212 & new_n1330;
  assign new_n1332 = new_n1331 ^ n287;
  assign new_n1333 = new_n1332 ^ n416;
  assign new_n1334 = ~new_n1211 & ~new_n1333;
  assign new_n1335 = new_n1334 ^ n416;
  assign new_n1336 = new_n1335 ^ n417;
  assign new_n1337 = ~new_n1210 & new_n1336;
  assign new_n1338 = new_n1337 ^ n417;
  assign new_n1339 = new_n1338 ^ n418;
  assign new_n1340 = ~new_n1209 & new_n1339;
  assign new_n1341 = new_n1340 ^ n418;
  assign new_n1342 = new_n1341 ^ n419;
  assign new_n1343 = ~new_n1208 & ~new_n1342;
  assign new_n1344 = new_n1343 ^ n291;
  assign new_n1345 = new_n1344 ^ n420;
  assign new_n1346 = ~new_n1207 & new_n1345;
  assign new_n1347 = new_n1346 ^ n292;
  assign new_n1348 = new_n1347 ^ n421;
  assign new_n1349 = ~new_n1206 & new_n1348;
  assign new_n1350 = new_n1349 ^ n293;
  assign new_n1351 = new_n1350 ^ n422;
  assign new_n1352 = ~new_n1205 & new_n1351;
  assign new_n1353 = new_n1352 ^ n294;
  assign new_n1354 = new_n1353 ^ n423;
  assign new_n1355 = ~new_n1204 & ~new_n1354;
  assign new_n1356 = new_n1355 ^ n423;
  assign new_n1357 = ~new_n1197 & new_n1356;
  assign new_n1358 = ~new_n1357 & new_n1203;
  assign new_n1359 = n427 ^ n299;
  assign new_n1360 = n426 ^ n298;
  assign new_n1361 = new_n1200 ^ n426;
  assign new_n1362 = ~new_n1360 & ~new_n1361;
  assign new_n1363 = new_n1362 ^ n426;
  assign new_n1364 = new_n1363 ^ n427;
  assign new_n1365 = ~new_n1359 & new_n1364;
  assign new_n1366 = new_n1365 ^ n427;
  assign new_n1367 = n428 ^ n300;
  assign new_n1368 = ~n300 & n428;
  assign new_n1369 = new_n1368 ^ new_n1367;
  assign new_n1370 = ~new_n1369 & new_n1366;
  assign new_n1371 = ~new_n1358 & new_n1370;
  assign new_n1372 = ~n303 & n431;
  assign new_n1373 = ~n302 & n430;
  assign new_n1374 = ~new_n1372 & ~new_n1373;
  assign new_n1375 = n429 ^ n301;
  assign new_n1376 = ~n429 & n301;
  assign new_n1377 = new_n1376 ^ new_n1375;
  assign new_n1378 = ~new_n1368 & ~new_n1377;
  assign new_n1379 = new_n1374 & new_n1378;
  assign new_n1380 = ~new_n1371 & new_n1379;
  assign new_n1381 = n431 ^ n303;
  assign new_n1382 = n430 ^ n302;
  assign new_n1383 = new_n1376 ^ n430;
  assign new_n1384 = ~new_n1382 & ~new_n1383;
  assign new_n1385 = new_n1384 ^ n430;
  assign new_n1386 = new_n1385 ^ n431;
  assign new_n1387 = ~new_n1381 & new_n1386;
  assign new_n1388 = new_n1387 ^ n431;
  assign new_n1389 = n432 ^ n304;
  assign new_n1390 = ~n304 & n432;
  assign new_n1391 = new_n1390 ^ new_n1389;
  assign new_n1392 = ~new_n1391 & new_n1388;
  assign new_n1393 = ~new_n1380 & new_n1392;
  assign new_n1394 = n433 ^ n305;
  assign new_n1395 = ~n433 & n305;
  assign new_n1396 = new_n1395 ^ new_n1394;
  assign new_n1397 = ~new_n1390 & ~new_n1396;
  assign new_n1398 = ~new_n1393 & new_n1397;
  assign new_n1399 = n434 ^ n306;
  assign new_n1400 = ~n306 & n434;
  assign new_n1401 = new_n1400 ^ new_n1399;
  assign new_n1402 = ~new_n1395 & ~new_n1401;
  assign new_n1403 = ~new_n1398 & new_n1402;
  assign new_n1404 = n435 ^ n307;
  assign new_n1405 = ~n435 & n307;
  assign new_n1406 = new_n1405 ^ new_n1404;
  assign new_n1407 = ~new_n1400 & ~new_n1406;
  assign new_n1408 = ~new_n1403 & new_n1407;
  assign new_n1409 = ~new_n1189 & ~new_n1405;
  assign new_n1410 = ~new_n1408 & new_n1409;
  assign new_n1411 = new_n1410 ^ n437;
  assign new_n1412 = new_n1411 ^ n437;
  assign new_n1413 = ~new_n1192 & ~new_n1412;
  assign new_n1414 = new_n1413 ^ n437;
  assign new_n1415 = ~new_n1187 & new_n1414;
  assign new_n1416 = new_n1415 ^ n309;
  assign new_n1417 = new_n1416 ^ n438;
  assign new_n1418 = ~new_n1186 & ~new_n1417;
  assign new_n1419 = new_n1418 ^ n438;
  assign new_n1420 = new_n1419 ^ n439;
  assign new_n1421 = ~new_n1185 & new_n1420;
  assign new_n1422 = new_n1421 ^ n439;
  assign new_n1423 = new_n1422 ^ n440;
  assign new_n1424 = ~new_n1184 & new_n1423;
  assign new_n1425 = new_n1424 ^ n440;
  assign new_n1426 = new_n1425 ^ n441;
  assign new_n1427 = ~new_n1183 & new_n1426;
  assign new_n1428 = new_n1427 ^ n441;
  assign new_n1429 = new_n1428 ^ n442;
  assign new_n1430 = ~new_n1182 & ~new_n1429;
  assign new_n1431 = new_n1430 ^ n314;
  assign new_n1432 = new_n1431 ^ n443;
  assign new_n1433 = ~new_n1181 & new_n1432;
  assign new_n1434 = new_n1433 ^ n315;
  assign new_n1435 = n444 ^ n316;
  assign new_n1436 = ~n316 & n444;
  assign new_n1437 = new_n1436 ^ new_n1435;
  assign new_n1438 = ~new_n1434 & ~new_n1437;
  assign new_n1439 = n445 ^ n317;
  assign new_n1440 = ~n445 & n317;
  assign new_n1441 = new_n1440 ^ new_n1439;
  assign new_n1442 = ~new_n1436 & ~new_n1441;
  assign new_n1443 = n447 ^ n319;
  assign new_n1444 = ~n447 & n319;
  assign new_n1445 = new_n1444 ^ new_n1443;
  assign new_n1446 = n446 ^ n318;
  assign new_n1447 = ~n446 & n318;
  assign new_n1448 = new_n1447 ^ new_n1446;
  assign new_n1449 = ~new_n1445 & ~new_n1448;
  assign new_n1450 = ~n320 & n448;
  assign new_n1451 = ~new_n1450 & new_n1449;
  assign new_n1452 = new_n1442 & new_n1451;
  assign new_n1453 = ~new_n1438 & new_n1452;
  assign new_n1454 = ~new_n1440 & ~new_n1447;
  assign new_n1455 = ~new_n1454 & new_n1451;
  assign new_n1456 = n448 ^ n320;
  assign new_n1457 = new_n1444 ^ n448;
  assign new_n1458 = ~new_n1456 & new_n1457;
  assign new_n1459 = new_n1458 ^ n320;
  assign new_n1460 = ~new_n1177 & ~new_n1459;
  assign new_n1461 = ~new_n1455 & new_n1460;
  assign new_n1462 = ~new_n1453 & new_n1461;
  assign new_n1463 = new_n1462 ^ n450;
  assign new_n1464 = new_n1463 ^ n450;
  assign new_n1465 = ~new_n1180 & ~new_n1464;
  assign new_n1466 = new_n1465 ^ n450;
  assign new_n1467 = ~new_n1175 & new_n1466;
  assign new_n1468 = new_n1467 ^ n322;
  assign new_n1469 = new_n1468 ^ n451;
  assign new_n1470 = ~new_n1174 & ~new_n1469;
  assign new_n1471 = new_n1470 ^ n451;
  assign new_n1472 = ~new_n1167 & new_n1471;
  assign new_n1473 = ~new_n1472 & new_n1173;
  assign new_n1474 = n455 ^ n327;
  assign new_n1475 = n454 ^ n326;
  assign new_n1476 = new_n1170 ^ n454;
  assign new_n1477 = ~new_n1475 & ~new_n1476;
  assign new_n1478 = new_n1477 ^ n454;
  assign new_n1479 = new_n1478 ^ n455;
  assign new_n1480 = ~new_n1474 & new_n1479;
  assign new_n1481 = new_n1480 ^ n455;
  assign new_n1482 = ~new_n1159 & new_n1481;
  assign new_n1483 = ~new_n1473 & new_n1482;
  assign new_n1484 = new_n1483 ^ n457;
  assign new_n1485 = new_n1484 ^ n457;
  assign new_n1486 = ~new_n1162 & ~new_n1485;
  assign new_n1487 = new_n1486 ^ n457;
  assign new_n1488 = ~new_n1157 & new_n1487;
  assign new_n1489 = new_n1488 ^ n329;
  assign new_n1490 = new_n1489 ^ n458;
  assign new_n1491 = ~new_n1156 & ~new_n1490;
  assign new_n1492 = new_n1491 ^ n458;
  assign new_n1493 = new_n1492 ^ n459;
  assign new_n1494 = ~new_n1155 & ~new_n1493;
  assign new_n1495 = new_n1494 ^ n331;
  assign new_n1496 = new_n1495 ^ n460;
  assign new_n1497 = ~new_n1154 & new_n1496;
  assign new_n1498 = new_n1497 ^ n332;
  assign new_n1499 = new_n1498 ^ n461;
  assign new_n1500 = ~new_n1153 & ~new_n1499;
  assign new_n1501 = new_n1500 ^ n461;
  assign new_n1502 = new_n1501 ^ n462;
  assign new_n1503 = ~new_n1152 & ~new_n1502;
  assign new_n1504 = new_n1503 ^ n334;
  assign new_n1505 = new_n1504 ^ n463;
  assign new_n1506 = ~new_n1151 & new_n1505;
  assign new_n1507 = new_n1506 ^ n335;
  assign new_n1508 = new_n1507 ^ n464;
  assign new_n1509 = ~new_n1150 & ~new_n1508;
  assign new_n1510 = new_n1509 ^ n464;
  assign new_n1511 = new_n1510 ^ n465;
  assign new_n1512 = ~new_n1149 & new_n1511;
  assign new_n1513 = new_n1512 ^ n465;
  assign new_n1514 = new_n1513 ^ n466;
  assign new_n1515 = ~new_n1148 & ~new_n1514;
  assign new_n1516 = new_n1515 ^ n338;
  assign new_n1517 = new_n1516 ^ n467;
  assign new_n1518 = ~new_n1147 & new_n1517;
  assign new_n1519 = new_n1518 ^ n339;
  assign new_n1520 = new_n1519 ^ n468;
  assign new_n1521 = ~new_n1146 & ~new_n1520;
  assign new_n1522 = new_n1521 ^ n468;
  assign new_n1523 = new_n1522 ^ n469;
  assign new_n1524 = ~new_n1145 & new_n1523;
  assign new_n1525 = new_n1524 ^ n469;
  assign new_n1526 = new_n1525 ^ n470;
  assign new_n1527 = ~new_n1144 & new_n1526;
  assign new_n1528 = new_n1527 ^ n470;
  assign new_n1529 = new_n1528 ^ n471;
  assign new_n1530 = ~new_n1143 & ~new_n1529;
  assign new_n1531 = new_n1530 ^ n343;
  assign new_n1532 = new_n1531 ^ n472;
  assign new_n1533 = ~new_n1142 & new_n1532;
  assign new_n1534 = new_n1533 ^ n344;
  assign new_n1535 = new_n1534 ^ n473;
  assign new_n1536 = ~new_n1141 & new_n1535;
  assign new_n1537 = new_n1536 ^ n345;
  assign new_n1538 = new_n1537 ^ n474;
  assign new_n1539 = ~new_n1140 & new_n1538;
  assign new_n1540 = new_n1539 ^ n346;
  assign new_n1541 = new_n1540 ^ n475;
  assign new_n1542 = ~new_n1139 & ~new_n1541;
  assign new_n1543 = new_n1542 ^ n475;
  assign new_n1544 = new_n1543 ^ n476;
  assign new_n1545 = ~new_n1138 & ~new_n1544;
  assign new_n1546 = new_n1545 ^ n348;
  assign new_n1547 = new_n1546 ^ n477;
  assign new_n1548 = ~new_n1137 & new_n1547;
  assign new_n1549 = new_n1548 ^ n349;
  assign new_n1550 = new_n1549 ^ n478;
  assign new_n1551 = ~new_n1136 & ~new_n1550;
  assign new_n1552 = new_n1551 ^ n478;
  assign new_n1553 = new_n1552 ^ n479;
  assign new_n1554 = ~new_n1135 & new_n1553;
  assign new_n1555 = new_n1554 ^ n479;
  assign new_n1556 = new_n1555 ^ n480;
  assign new_n1557 = ~new_n1134 & new_n1556;
  assign new_n1558 = new_n1557 ^ n480;
  assign new_n1559 = new_n1558 ^ n481;
  assign new_n1560 = ~new_n1133 & new_n1559;
  assign new_n1561 = new_n1560 ^ n481;
  assign new_n1562 = new_n1561 ^ n482;
  assign new_n1563 = ~new_n1132 & ~new_n1562;
  assign new_n1564 = new_n1563 ^ n354;
  assign new_n1565 = new_n1564 ^ n483;
  assign new_n1566 = ~new_n1131 & new_n1565;
  assign new_n1567 = new_n1566 ^ n355;
  assign new_n1568 = new_n1567 ^ n484;
  assign new_n1569 = ~new_n1130 & ~new_n1568;
  assign new_n1570 = new_n1569 ^ n484;
  assign new_n1571 = new_n1570 ^ n485;
  assign new_n1572 = ~new_n1129 & new_n1571;
  assign new_n1573 = new_n1572 ^ n485;
  assign new_n1574 = new_n1573 ^ n486;
  assign new_n1575 = ~new_n1128 & new_n1574;
  assign new_n1576 = new_n1575 ^ n486;
  assign new_n1577 = new_n1576 ^ n487;
  assign new_n1578 = ~new_n1127 & ~new_n1577;
  assign new_n1579 = new_n1578 ^ n359;
  assign new_n1580 = new_n1579 ^ n488;
  assign new_n1581 = ~new_n1126 & new_n1580;
  assign new_n1582 = new_n1581 ^ n360;
  assign new_n1583 = new_n1582 ^ n489;
  assign new_n1584 = ~new_n1125 & new_n1583;
  assign new_n1585 = new_n1584 ^ n361;
  assign new_n1586 = new_n1585 ^ n490;
  assign new_n1587 = ~new_n1124 & new_n1586;
  assign new_n1588 = new_n1587 ^ n362;
  assign new_n1589 = new_n1588 ^ n491;
  assign new_n1590 = ~new_n1123 & new_n1589;
  assign new_n1591 = new_n1590 ^ n363;
  assign new_n1592 = new_n1591 ^ n492;
  assign new_n1593 = ~new_n1122 & new_n1592;
  assign new_n1594 = new_n1593 ^ n364;
  assign new_n1595 = new_n1594 ^ n493;
  assign new_n1596 = ~new_n1121 & ~new_n1595;
  assign new_n1597 = new_n1596 ^ n493;
  assign new_n1598 = new_n1597 ^ n494;
  assign new_n1599 = ~new_n1120 & ~new_n1598;
  assign new_n1600 = new_n1599 ^ n366;
  assign new_n1601 = new_n1600 ^ n495;
  assign new_n1602 = ~new_n1119 & new_n1601;
  assign new_n1603 = new_n1602 ^ n367;
  assign new_n1604 = new_n1603 ^ n496;
  assign new_n1605 = ~new_n1118 & ~new_n1604;
  assign new_n1606 = new_n1605 ^ n496;
  assign new_n1607 = new_n1606 ^ n497;
  assign new_n1608 = ~new_n1117 & new_n1607;
  assign new_n1609 = new_n1608 ^ n497;
  assign new_n1610 = new_n1609 ^ n498;
  assign new_n1611 = ~new_n1116 & new_n1610;
  assign new_n1612 = new_n1611 ^ n498;
  assign new_n1613 = new_n1612 ^ n499;
  assign new_n1614 = ~new_n1115 & new_n1613;
  assign new_n1615 = new_n1614 ^ n499;
  assign new_n1616 = new_n1615 ^ n500;
  assign new_n1617 = ~new_n1114 & ~new_n1616;
  assign new_n1618 = new_n1617 ^ n372;
  assign new_n1619 = new_n1618 ^ n501;
  assign new_n1620 = ~new_n1113 & new_n1619;
  assign new_n1621 = new_n1620 ^ n373;
  assign new_n1622 = new_n1621 ^ n502;
  assign new_n1623 = ~new_n1112 & ~new_n1622;
  assign new_n1624 = new_n1623 ^ n502;
  assign new_n1625 = new_n1624 ^ n503;
  assign new_n1626 = ~new_n1111 & ~new_n1625;
  assign new_n1627 = new_n1626 ^ n375;
  assign new_n1628 = new_n1627 ^ n504;
  assign new_n1629 = ~new_n1110 & new_n1628;
  assign new_n1630 = new_n1629 ^ n376;
  assign new_n1631 = new_n1630 ^ n505;
  assign new_n1632 = ~new_n1109 & ~new_n1631;
  assign new_n1633 = new_n1632 ^ n505;
  assign new_n1634 = new_n1633 ^ n506;
  assign new_n1635 = ~new_n1108 & new_n1634;
  assign new_n1636 = new_n1635 ^ n506;
  assign new_n1637 = new_n1636 ^ n507;
  assign new_n1638 = ~new_n1107 & new_n1637;
  assign new_n1639 = new_n1638 ^ n507;
  assign new_n1640 = ~new_n1103 & new_n1639;
  assign new_n1641 = ~new_n1640 & new_n1106;
  assign new_n1642 = new_n1641 ^ n512;
  assign new_n1643 = new_n1642 ^ n512;
  assign new_n1644 = ~new_n1643 & new_n1098;
  assign new_n1645 = new_n1644 ^ n512;
  assign new_n1646 = ~new_n1086 & new_n1645;
  assign new_n1647 = new_n1646 ^ n384;
  assign new_n1648 = new_n1085 & new_n1647;
  assign new_n1649 = new_n1648 ^ n383;
  assign new_n1650 = new_n1649 ^ new_n1084;
  assign new_n1651 = new_n1087 & new_n1647;
  assign new_n1652 = new_n1651 ^ n382;
  assign new_n1653 = new_n518 & new_n1082;
  assign new_n1654 = new_n1653 ^ n126;
  assign new_n1655 = new_n1654 ^ new_n1652;
  assign new_n1656 = new_n1088 & new_n1647;
  assign new_n1657 = new_n1656 ^ n381;
  assign new_n1658 = new_n519 & new_n1082;
  assign new_n1659 = new_n1658 ^ n125;
  assign new_n1660 = new_n1659 ^ new_n1657;
  assign new_n1661 = new_n1102 & new_n1647;
  assign new_n1662 = new_n1661 ^ n380;
  assign new_n1663 = new_n533 & new_n1082;
  assign new_n1664 = new_n1663 ^ n124;
  assign new_n1665 = new_n1664 ^ new_n1662;
  assign new_n1666 = new_n1107 & new_n1647;
  assign new_n1667 = new_n1666 ^ n379;
  assign new_n1668 = new_n538 & new_n1082;
  assign new_n1669 = new_n1668 ^ n123;
  assign new_n1670 = new_n1669 ^ new_n1667;
  assign new_n1671 = new_n1108 & new_n1647;
  assign new_n1672 = new_n1671 ^ n378;
  assign new_n1673 = new_n539 & new_n1082;
  assign new_n1674 = new_n1673 ^ n122;
  assign new_n1675 = new_n1674 ^ new_n1672;
  assign new_n1676 = new_n540 & new_n1082;
  assign new_n1677 = new_n1676 ^ n121;
  assign new_n1678 = new_n1109 & new_n1647;
  assign new_n1679 = new_n1678 ^ n377;
  assign new_n1680 = new_n1679 ^ new_n1677;
  assign new_n1681 = new_n1110 & new_n1647;
  assign new_n1682 = new_n1681 ^ n376;
  assign new_n1683 = new_n541 & new_n1082;
  assign new_n1684 = new_n1683 ^ n120;
  assign new_n1685 = new_n1684 ^ new_n1682;
  assign new_n1686 = new_n1111 & new_n1647;
  assign new_n1687 = new_n1686 ^ n375;
  assign new_n1688 = new_n542 & new_n1082;
  assign new_n1689 = new_n1688 ^ n119;
  assign new_n1690 = new_n1689 ^ new_n1687;
  assign new_n1691 = new_n1112 & new_n1647;
  assign new_n1692 = new_n1691 ^ n374;
  assign new_n1693 = new_n543 & new_n1082;
  assign new_n1694 = new_n1693 ^ n118;
  assign new_n1695 = new_n1694 ^ new_n1692;
  assign new_n1696 = new_n544 & new_n1082;
  assign new_n1697 = new_n1696 ^ n117;
  assign new_n1698 = new_n1113 & new_n1647;
  assign new_n1699 = new_n1698 ^ n373;
  assign new_n1700 = new_n1699 ^ new_n1697;
  assign new_n1701 = new_n545 & new_n1082;
  assign new_n1702 = new_n1701 ^ n116;
  assign new_n1703 = new_n1114 & new_n1647;
  assign new_n1704 = new_n1703 ^ n372;
  assign new_n1705 = new_n1704 ^ new_n1702;
  assign new_n1706 = new_n1115 & new_n1647;
  assign new_n1707 = new_n1706 ^ n371;
  assign new_n1708 = new_n546 & new_n1082;
  assign new_n1709 = new_n1708 ^ n115;
  assign new_n1710 = new_n1709 ^ new_n1707;
  assign new_n1711 = new_n1116 & new_n1647;
  assign new_n1712 = new_n1711 ^ n370;
  assign new_n1713 = new_n547 & new_n1082;
  assign new_n1714 = new_n1713 ^ n114;
  assign new_n1715 = new_n1714 ^ new_n1712;
  assign new_n1716 = new_n1117 & new_n1647;
  assign new_n1717 = new_n1716 ^ n369;
  assign new_n1718 = new_n548 & new_n1082;
  assign new_n1719 = new_n1718 ^ n113;
  assign new_n1720 = new_n1719 ^ new_n1717;
  assign new_n1721 = new_n1118 & new_n1647;
  assign new_n1722 = new_n1721 ^ n368;
  assign new_n1723 = new_n549 & new_n1082;
  assign new_n1724 = new_n1723 ^ n112;
  assign new_n1725 = new_n1724 ^ new_n1722;
  assign new_n1726 = new_n550 & new_n1082;
  assign new_n1727 = new_n1726 ^ n111;
  assign new_n1728 = new_n1119 & new_n1647;
  assign new_n1729 = new_n1728 ^ n367;
  assign new_n1730 = new_n1729 ^ new_n1727;
  assign new_n1731 = new_n551 & new_n1082;
  assign new_n1732 = new_n1731 ^ n110;
  assign new_n1733 = new_n1120 & new_n1647;
  assign new_n1734 = new_n1733 ^ n366;
  assign new_n1735 = new_n1734 ^ new_n1732;
  assign new_n1736 = new_n552 & new_n1082;
  assign new_n1737 = new_n1736 ^ n109;
  assign new_n1738 = new_n1121 & new_n1647;
  assign new_n1739 = new_n1738 ^ n365;
  assign new_n1740 = new_n1739 ^ new_n1737;
  assign new_n1741 = new_n1122 & new_n1647;
  assign new_n1742 = new_n1741 ^ n364;
  assign new_n1743 = new_n553 & new_n1082;
  assign new_n1744 = new_n1743 ^ n108;
  assign new_n1745 = new_n1744 ^ new_n1742;
  assign new_n1746 = new_n1123 & new_n1647;
  assign new_n1747 = new_n1746 ^ n363;
  assign new_n1748 = new_n554 & new_n1082;
  assign new_n1749 = new_n1748 ^ n107;
  assign new_n1750 = new_n1749 ^ new_n1747;
  assign new_n1751 = new_n1124 & new_n1647;
  assign new_n1752 = new_n1751 ^ n362;
  assign new_n1753 = new_n555 & new_n1082;
  assign new_n1754 = new_n1753 ^ n106;
  assign new_n1755 = new_n1754 ^ new_n1752;
  assign new_n1756 = new_n556 & new_n1082;
  assign new_n1757 = new_n1756 ^ n105;
  assign new_n1758 = new_n1125 & new_n1647;
  assign new_n1759 = new_n1758 ^ n361;
  assign new_n1760 = new_n1759 ^ new_n1757;
  assign new_n1761 = new_n557 & new_n1082;
  assign new_n1762 = new_n1761 ^ n104;
  assign new_n1763 = new_n1126 & new_n1647;
  assign new_n1764 = new_n1763 ^ n360;
  assign new_n1765 = new_n1764 ^ new_n1762;
  assign new_n1766 = new_n1127 & new_n1647;
  assign new_n1767 = new_n1766 ^ n359;
  assign new_n1768 = new_n558 & new_n1082;
  assign new_n1769 = new_n1768 ^ n103;
  assign new_n1770 = new_n1769 ^ new_n1767;
  assign new_n1771 = new_n559 & new_n1082;
  assign new_n1772 = new_n1771 ^ n102;
  assign new_n1773 = new_n1128 & new_n1647;
  assign new_n1774 = new_n1773 ^ n358;
  assign new_n1775 = new_n1774 ^ new_n1772;
  assign new_n1776 = new_n560 & new_n1082;
  assign new_n1777 = new_n1776 ^ n101;
  assign new_n1778 = new_n1129 & new_n1647;
  assign new_n1779 = new_n1778 ^ n357;
  assign new_n1780 = new_n1779 ^ new_n1777;
  assign new_n1781 = new_n1130 & new_n1647;
  assign new_n1782 = new_n1781 ^ n356;
  assign new_n1783 = new_n561 & new_n1082;
  assign new_n1784 = new_n1783 ^ n100;
  assign new_n1785 = new_n1784 ^ new_n1782;
  assign new_n1786 = new_n1131 & new_n1647;
  assign new_n1787 = new_n1786 ^ n355;
  assign new_n1788 = new_n562 & new_n1082;
  assign new_n1789 = new_n1788 ^ n99;
  assign new_n1790 = new_n1789 ^ new_n1787;
  assign new_n1791 = new_n563 & new_n1082;
  assign new_n1792 = new_n1791 ^ n98;
  assign new_n1793 = new_n1132 & new_n1647;
  assign new_n1794 = new_n1793 ^ n354;
  assign new_n1795 = new_n1794 ^ new_n1792;
  assign new_n1796 = new_n1133 & new_n1647;
  assign new_n1797 = new_n1796 ^ n353;
  assign new_n1798 = new_n564 & new_n1082;
  assign new_n1799 = new_n1798 ^ n97;
  assign new_n1800 = new_n1799 ^ new_n1797;
  assign new_n1801 = new_n1134 & new_n1647;
  assign new_n1802 = new_n1801 ^ n352;
  assign new_n1803 = new_n565 & new_n1082;
  assign new_n1804 = new_n1803 ^ n96;
  assign new_n1805 = new_n1804 ^ new_n1802;
  assign new_n1806 = new_n1135 & new_n1647;
  assign new_n1807 = new_n1806 ^ n351;
  assign new_n1808 = new_n566 & new_n1082;
  assign new_n1809 = new_n1808 ^ n95;
  assign new_n1810 = new_n1809 ^ new_n1807;
  assign new_n1811 = new_n1136 & new_n1647;
  assign new_n1812 = new_n1811 ^ n350;
  assign new_n1813 = new_n567 & new_n1082;
  assign new_n1814 = new_n1813 ^ n94;
  assign new_n1815 = new_n1814 ^ new_n1812;
  assign new_n1816 = new_n568 & new_n1082;
  assign new_n1817 = new_n1816 ^ n93;
  assign new_n1818 = new_n1137 & new_n1647;
  assign new_n1819 = new_n1818 ^ n349;
  assign new_n1820 = new_n1819 ^ new_n1817;
  assign new_n1821 = new_n569 & new_n1082;
  assign new_n1822 = new_n1821 ^ n92;
  assign new_n1823 = new_n1138 & new_n1647;
  assign new_n1824 = new_n1823 ^ n348;
  assign new_n1825 = new_n1824 ^ new_n1822;
  assign new_n1826 = new_n570 & new_n1082;
  assign new_n1827 = new_n1826 ^ n91;
  assign new_n1828 = new_n1139 & new_n1647;
  assign new_n1829 = new_n1828 ^ n347;
  assign new_n1830 = new_n1829 ^ new_n1827;
  assign new_n1831 = new_n1140 & new_n1647;
  assign new_n1832 = new_n1831 ^ n346;
  assign new_n1833 = new_n571 & new_n1082;
  assign new_n1834 = new_n1833 ^ n90;
  assign new_n1835 = new_n1834 ^ new_n1832;
  assign new_n1836 = new_n572 & new_n1082;
  assign new_n1837 = new_n1836 ^ n89;
  assign new_n1838 = new_n1141 & new_n1647;
  assign new_n1839 = new_n1838 ^ n345;
  assign new_n1840 = new_n1839 ^ new_n1837;
  assign new_n1841 = new_n573 & new_n1082;
  assign new_n1842 = new_n1841 ^ n88;
  assign new_n1843 = new_n1142 & new_n1647;
  assign new_n1844 = new_n1843 ^ n344;
  assign new_n1845 = new_n1844 ^ new_n1842;
  assign new_n1846 = new_n574 & new_n1082;
  assign new_n1847 = new_n1846 ^ n87;
  assign new_n1848 = new_n1143 & new_n1647;
  assign new_n1849 = new_n1848 ^ n343;
  assign new_n1850 = new_n1849 ^ new_n1847;
  assign new_n1851 = new_n575 & new_n1082;
  assign new_n1852 = new_n1851 ^ n86;
  assign new_n1853 = new_n1144 & new_n1647;
  assign new_n1854 = new_n1853 ^ n342;
  assign new_n1855 = new_n1854 ^ new_n1852;
  assign new_n1856 = new_n1145 & new_n1647;
  assign new_n1857 = new_n1856 ^ n341;
  assign new_n1858 = new_n576 & new_n1082;
  assign new_n1859 = new_n1858 ^ n85;
  assign new_n1860 = new_n1859 ^ new_n1857;
  assign new_n1861 = new_n577 & new_n1082;
  assign new_n1862 = new_n1861 ^ n84;
  assign new_n1863 = new_n1146 & new_n1647;
  assign new_n1864 = new_n1863 ^ n340;
  assign new_n1865 = new_n1864 ^ new_n1862;
  assign new_n1866 = new_n1147 & new_n1647;
  assign new_n1867 = new_n1866 ^ n339;
  assign new_n1868 = new_n578 & new_n1082;
  assign new_n1869 = new_n1868 ^ n83;
  assign new_n1870 = new_n1869 ^ new_n1867;
  assign new_n1871 = new_n579 & new_n1082;
  assign new_n1872 = new_n1871 ^ n82;
  assign new_n1873 = new_n1148 & new_n1647;
  assign new_n1874 = new_n1873 ^ n338;
  assign new_n1875 = new_n1874 ^ new_n1872;
  assign new_n1876 = new_n580 & new_n1082;
  assign new_n1877 = new_n1876 ^ n81;
  assign new_n1878 = new_n1149 & new_n1647;
  assign new_n1879 = new_n1878 ^ n337;
  assign new_n1880 = new_n1879 ^ new_n1877;
  assign new_n1881 = new_n939 & new_n1082;
  assign new_n1882 = new_n1881 ^ n80;
  assign new_n1883 = new_n1150 & new_n1647;
  assign new_n1884 = new_n1883 ^ n336;
  assign new_n1885 = new_n1884 ^ new_n1882;
  assign new_n1886 = new_n1151 & new_n1647;
  assign new_n1887 = new_n1886 ^ n335;
  assign new_n1888 = new_n934 & new_n1082;
  assign new_n1889 = new_n1888 ^ n79;
  assign new_n1890 = new_n1889 ^ new_n1887;
  assign new_n1891 = new_n929 & new_n1082;
  assign new_n1892 = new_n1891 ^ n78;
  assign new_n1893 = new_n1152 & new_n1647;
  assign new_n1894 = new_n1893 ^ n334;
  assign new_n1895 = new_n1894 ^ new_n1892;
  assign new_n1896 = new_n1153 & new_n1647;
  assign new_n1897 = new_n1896 ^ n333;
  assign new_n1898 = new_n924 & new_n1082;
  assign new_n1899 = new_n1898 ^ n77;
  assign new_n1900 = new_n1899 ^ new_n1897;
  assign new_n1901 = new_n1154 & new_n1647;
  assign new_n1902 = new_n1901 ^ n332;
  assign new_n1903 = new_n919 & new_n1082;
  assign new_n1904 = new_n1903 ^ n76;
  assign new_n1905 = new_n1904 ^ new_n1902;
  assign new_n1906 = new_n1155 & new_n1647;
  assign new_n1907 = new_n1906 ^ n331;
  assign new_n1908 = new_n914 & new_n1082;
  assign new_n1909 = new_n1908 ^ n75;
  assign new_n1910 = new_n1909 ^ new_n1907;
  assign new_n1911 = new_n1156 & new_n1647;
  assign new_n1912 = new_n1911 ^ n330;
  assign new_n1913 = new_n909 & new_n1082;
  assign new_n1914 = new_n1913 ^ n74;
  assign new_n1915 = new_n1914 ^ new_n1912;
  assign new_n1916 = new_n904 & new_n1082;
  assign new_n1917 = new_n1916 ^ n73;
  assign new_n1918 = new_n1157 & new_n1647;
  assign new_n1919 = new_n1918 ^ n329;
  assign new_n1920 = new_n1919 ^ new_n1917;
  assign new_n1921 = new_n899 & new_n1082;
  assign new_n1922 = new_n1921 ^ n72;
  assign new_n1923 = new_n1158 & new_n1647;
  assign new_n1924 = new_n1923 ^ n328;
  assign new_n1925 = new_n1924 ^ new_n1922;
  assign new_n1926 = new_n1474 & new_n1647;
  assign new_n1927 = new_n1926 ^ n327;
  assign new_n1928 = new_n891 & new_n1082;
  assign new_n1929 = new_n1928 ^ n71;
  assign new_n1930 = new_n1929 ^ new_n1927;
  assign new_n1931 = new_n892 & new_n1082;
  assign new_n1932 = new_n1931 ^ n70;
  assign new_n1933 = new_n1475 & new_n1647;
  assign new_n1934 = new_n1933 ^ n326;
  assign new_n1935 = new_n1934 ^ new_n1932;
  assign new_n1936 = new_n1169 & new_n1647;
  assign new_n1937 = new_n1936 ^ n325;
  assign new_n1938 = new_n588 & new_n1082;
  assign new_n1939 = new_n1938 ^ n69;
  assign new_n1940 = new_n1939 ^ new_n1937;
  assign new_n1941 = new_n592 & new_n1082;
  assign new_n1942 = new_n1941 ^ n68;
  assign new_n1943 = new_n1166 & new_n1647;
  assign new_n1944 = new_n1943 ^ n324;
  assign new_n1945 = new_n1944 ^ new_n1942;
  assign new_n1946 = new_n593 & new_n1082;
  assign new_n1947 = new_n1946 ^ n67;
  assign new_n1948 = new_n1174 & new_n1647;
  assign new_n1949 = new_n1948 ^ n323;
  assign new_n1950 = new_n1949 ^ new_n1947;
  assign new_n1951 = new_n1175 & new_n1647;
  assign new_n1952 = new_n1951 ^ n322;
  assign new_n1953 = new_n594 & new_n1082;
  assign new_n1954 = new_n1953 ^ n66;
  assign new_n1955 = new_n1954 ^ new_n1952;
  assign new_n1956 = new_n595 & new_n1082;
  assign new_n1957 = new_n1956 ^ n65;
  assign new_n1958 = new_n1176 & new_n1647;
  assign new_n1959 = new_n1958 ^ n321;
  assign new_n1960 = new_n1959 ^ new_n1957;
  assign new_n1961 = new_n1456 & new_n1647;
  assign new_n1962 = new_n1961 ^ n320;
  assign new_n1963 = new_n596 & new_n1082;
  assign new_n1964 = new_n1963 ^ n64;
  assign new_n1965 = new_n1964 ^ new_n1962;
  assign new_n1966 = new_n865 & new_n1082;
  assign new_n1967 = new_n1966 ^ n63;
  assign new_n1968 = new_n1443 & new_n1647;
  assign new_n1969 = new_n1968 ^ n319;
  assign new_n1970 = new_n1969 ^ new_n1967;
  assign new_n1971 = new_n866 & new_n1082;
  assign new_n1972 = new_n1971 ^ n62;
  assign new_n1973 = new_n1446 & new_n1647;
  assign new_n1974 = new_n1973 ^ n318;
  assign new_n1975 = new_n1974 ^ new_n1972;
  assign new_n1976 = new_n607 & new_n1082;
  assign new_n1977 = new_n1976 ^ n61;
  assign new_n1978 = new_n1439 & new_n1647;
  assign new_n1979 = new_n1978 ^ n317;
  assign new_n1980 = new_n1979 ^ new_n1977;
  assign new_n1981 = new_n604 & new_n1082;
  assign new_n1982 = new_n1981 ^ n60;
  assign new_n1983 = new_n1435 & new_n1647;
  assign new_n1984 = new_n1983 ^ n316;
  assign new_n1985 = new_n1984 ^ new_n1982;
  assign new_n1986 = new_n1181 & new_n1647;
  assign new_n1987 = new_n1986 ^ n315;
  assign new_n1988 = new_n612 & new_n1082;
  assign new_n1989 = new_n1988 ^ n59;
  assign new_n1990 = new_n1989 ^ new_n1987;
  assign new_n1991 = new_n1182 & new_n1647;
  assign new_n1992 = new_n1991 ^ n314;
  assign new_n1993 = new_n613 & new_n1082;
  assign new_n1994 = new_n1993 ^ n58;
  assign new_n1995 = new_n1994 ^ new_n1992;
  assign new_n1996 = new_n614 & new_n1082;
  assign new_n1997 = new_n1996 ^ n57;
  assign new_n1998 = new_n1183 & new_n1647;
  assign new_n1999 = new_n1998 ^ n313;
  assign new_n2000 = new_n1999 ^ new_n1997;
  assign new_n2001 = new_n615 & new_n1082;
  assign new_n2002 = new_n2001 ^ n56;
  assign new_n2003 = new_n1184 & new_n1647;
  assign new_n2004 = new_n2003 ^ n312;
  assign new_n2005 = new_n2004 ^ new_n2002;
  assign new_n2006 = new_n616 & new_n1082;
  assign new_n2007 = new_n2006 ^ n55;
  assign new_n2008 = new_n1185 & new_n1647;
  assign new_n2009 = new_n2008 ^ n311;
  assign new_n2010 = new_n2009 ^ new_n2007;
  assign new_n2011 = new_n1186 & new_n1647;
  assign new_n2012 = new_n2011 ^ n310;
  assign new_n2013 = new_n617 & new_n1082;
  assign new_n2014 = new_n2013 ^ n54;
  assign new_n2015 = new_n2014 ^ new_n2012;
  assign new_n2016 = new_n618 & new_n1082;
  assign new_n2017 = new_n2016 ^ n53;
  assign new_n2018 = new_n1187 & new_n1647;
  assign new_n2019 = new_n2018 ^ n309;
  assign new_n2020 = new_n2019 ^ new_n2017;
  assign new_n2021 = new_n1188 & new_n1647;
  assign new_n2022 = new_n2021 ^ n308;
  assign new_n2023 = new_n619 & new_n1082;
  assign new_n2024 = new_n2023 ^ n52;
  assign new_n2025 = new_n2024 ^ new_n2022;
  assign new_n2026 = new_n620 & new_n1082;
  assign new_n2027 = new_n2026 ^ n51;
  assign new_n2028 = new_n1404 & new_n1647;
  assign new_n2029 = new_n2028 ^ n307;
  assign new_n2030 = new_n2029 ^ new_n2027;
  assign new_n2031 = new_n621 & new_n1082;
  assign new_n2032 = new_n2031 ^ n50;
  assign new_n2033 = new_n1399 & new_n1647;
  assign new_n2034 = new_n2033 ^ n306;
  assign new_n2035 = new_n2034 ^ new_n2032;
  assign new_n2036 = new_n1394 & new_n1647;
  assign new_n2037 = new_n2036 ^ n305;
  assign new_n2038 = new_n622 & new_n1082;
  assign new_n2039 = new_n2038 ^ n49;
  assign new_n2040 = new_n2039 ^ new_n2037;
  assign new_n2041 = new_n823 & new_n1082;
  assign new_n2042 = new_n2041 ^ n48;
  assign new_n2043 = new_n1389 & new_n1647;
  assign new_n2044 = new_n2043 ^ n304;
  assign new_n2045 = new_n2044 ^ new_n2042;
  assign new_n2046 = new_n815 & new_n1082;
  assign new_n2047 = new_n2046 ^ n47;
  assign new_n2048 = new_n1381 & new_n1647;
  assign new_n2049 = new_n2048 ^ n303;
  assign new_n2050 = new_n2049 ^ new_n2047;
  assign new_n2051 = new_n816 & new_n1082;
  assign new_n2052 = new_n2051 ^ n46;
  assign new_n2053 = new_n1382 & new_n1647;
  assign new_n2054 = new_n2053 ^ n302;
  assign new_n2055 = new_n2054 ^ new_n2052;
  assign new_n2056 = new_n809 & new_n1082;
  assign new_n2057 = new_n2056 ^ n45;
  assign new_n2058 = new_n1375 & new_n1647;
  assign new_n2059 = new_n2058 ^ n301;
  assign new_n2060 = new_n2059 ^ new_n2057;
  assign new_n2061 = new_n1367 & new_n1647;
  assign new_n2062 = new_n2061 ^ n300;
  assign new_n2063 = new_n801 & new_n1082;
  assign new_n2064 = new_n2063 ^ n44;
  assign new_n2065 = new_n2064 ^ new_n2062;
  assign new_n2066 = new_n793 & new_n1082;
  assign new_n2067 = new_n2066 ^ n43;
  assign new_n2068 = new_n1359 & new_n1647;
  assign new_n2069 = new_n2068 ^ n299;
  assign new_n2070 = new_n2069 ^ new_n2067;
  assign new_n2071 = new_n794 & new_n1082;
  assign new_n2072 = new_n2071 ^ n42;
  assign new_n2073 = new_n1360 & new_n1647;
  assign new_n2074 = new_n2073 ^ n298;
  assign new_n2075 = new_n2074 ^ new_n2072;
  assign new_n2076 = new_n787 & new_n1082;
  assign new_n2077 = new_n2076 ^ n41;
  assign new_n2078 = new_n1199 & new_n1647;
  assign new_n2079 = new_n2078 ^ n297;
  assign new_n2080 = new_n2079 ^ new_n2077;
  assign new_n2081 = new_n780 & new_n1082;
  assign new_n2082 = new_n2081 ^ n40;
  assign new_n2083 = new_n1196 & new_n1647;
  assign new_n2084 = new_n2083 ^ n296;
  assign new_n2085 = new_n2084 ^ new_n2082;
  assign new_n2086 = new_n627 & new_n1082;
  assign new_n2087 = new_n2086 ^ n39;
  assign new_n2088 = new_n1204 & new_n1647;
  assign new_n2089 = new_n2088 ^ n295;
  assign new_n2090 = new_n2089 ^ new_n2087;
  assign new_n2091 = new_n1205 & new_n1647;
  assign new_n2092 = new_n2091 ^ n294;
  assign new_n2093 = new_n628 & new_n1082;
  assign new_n2094 = new_n2093 ^ n38;
  assign new_n2095 = new_n2094 ^ new_n2092;
  assign new_n2096 = new_n629 & new_n1082;
  assign new_n2097 = new_n2096 ^ n37;
  assign new_n2098 = new_n1206 & new_n1647;
  assign new_n2099 = new_n2098 ^ n293;
  assign new_n2100 = new_n2099 ^ new_n2097;
  assign new_n2101 = new_n1207 & new_n1647;
  assign new_n2102 = new_n2101 ^ n292;
  assign new_n2103 = new_n630 & new_n1082;
  assign new_n2104 = new_n2103 ^ n36;
  assign new_n2105 = new_n2104 ^ new_n2102;
  assign new_n2106 = new_n1208 & new_n1647;
  assign new_n2107 = new_n2106 ^ n291;
  assign new_n2108 = new_n631 & new_n1082;
  assign new_n2109 = new_n2108 ^ n35;
  assign new_n2110 = new_n2109 ^ new_n2107;
  assign new_n2111 = new_n632 & new_n1082;
  assign new_n2112 = new_n2111 ^ n34;
  assign new_n2113 = new_n1209 & new_n1647;
  assign new_n2114 = new_n2113 ^ n290;
  assign new_n2115 = new_n2114 ^ new_n2112;
  assign new_n2116 = new_n633 & new_n1082;
  assign new_n2117 = new_n2116 ^ n33;
  assign new_n2118 = new_n1210 & new_n1647;
  assign new_n2119 = new_n2118 ^ n289;
  assign new_n2120 = new_n2119 ^ new_n2117;
  assign new_n2121 = new_n634 & new_n1082;
  assign new_n2122 = new_n2121 ^ n32;
  assign new_n2123 = new_n1211 & new_n1647;
  assign new_n2124 = new_n2123 ^ n288;
  assign new_n2125 = new_n2124 ^ new_n2122;
  assign new_n2126 = new_n1212 & new_n1647;
  assign new_n2127 = new_n2126 ^ n287;
  assign new_n2128 = new_n635 & new_n1082;
  assign new_n2129 = new_n2128 ^ n31;
  assign new_n2130 = new_n2129 ^ new_n2127;
  assign new_n2131 = new_n636 & new_n1082;
  assign new_n2132 = new_n2131 ^ n30;
  assign new_n2133 = new_n1213 & new_n1647;
  assign new_n2134 = new_n2133 ^ n286;
  assign new_n2135 = new_n2134 ^ new_n2132;
  assign new_n2136 = new_n637 & new_n1082;
  assign new_n2137 = new_n2136 ^ n29;
  assign new_n2138 = new_n1214 & new_n1647;
  assign new_n2139 = new_n2138 ^ n285;
  assign new_n2140 = new_n2139 ^ new_n2137;
  assign new_n2141 = new_n1215 & new_n1647;
  assign new_n2142 = new_n2141 ^ n284;
  assign new_n2143 = new_n638 & new_n1082;
  assign new_n2144 = new_n2143 ^ n28;
  assign new_n2145 = new_n2144 ^ new_n2142;
  assign new_n2146 = new_n639 & new_n1082;
  assign new_n2147 = new_n2146 ^ n27;
  assign new_n2148 = new_n1216 & new_n1647;
  assign new_n2149 = new_n2148 ^ n283;
  assign new_n2150 = new_n2149 ^ new_n2147;
  assign new_n2151 = new_n640 & new_n1082;
  assign new_n2152 = new_n2151 ^ n26;
  assign new_n2153 = new_n1217 & new_n1647;
  assign new_n2154 = new_n2153 ^ n282;
  assign new_n2155 = new_n2154 ^ new_n2152;
  assign new_n2156 = new_n641 & new_n1082;
  assign new_n2157 = new_n2156 ^ n25;
  assign new_n2158 = new_n1218 & new_n1647;
  assign new_n2159 = new_n2158 ^ n281;
  assign new_n2160 = new_n2159 ^ new_n2157;
  assign new_n2161 = new_n642 & new_n1082;
  assign new_n2162 = new_n2161 ^ n24;
  assign new_n2163 = new_n1219 & new_n1647;
  assign new_n2164 = new_n2163 ^ n280;
  assign new_n2165 = new_n2164 ^ new_n2162;
  assign new_n2166 = new_n1220 & new_n1647;
  assign new_n2167 = new_n2166 ^ n279;
  assign new_n2168 = new_n643 & new_n1082;
  assign new_n2169 = new_n2168 ^ n23;
  assign new_n2170 = new_n2169 ^ new_n2167;
  assign new_n2171 = new_n1221 & new_n1647;
  assign new_n2172 = new_n2171 ^ n278;
  assign new_n2173 = new_n644 & new_n1082;
  assign new_n2174 = new_n2173 ^ n22;
  assign new_n2175 = new_n2174 ^ new_n2172;
  assign new_n2176 = new_n645 & new_n1082;
  assign new_n2177 = new_n2176 ^ n21;
  assign new_n2178 = new_n1222 & new_n1647;
  assign new_n2179 = new_n2178 ^ n277;
  assign new_n2180 = new_n2179 ^ new_n2177;
  assign new_n2181 = new_n1223 & new_n1647;
  assign new_n2182 = new_n2181 ^ n276;
  assign new_n2183 = new_n646 & new_n1082;
  assign new_n2184 = new_n2183 ^ n20;
  assign new_n2185 = new_n2184 ^ new_n2182;
  assign new_n2186 = new_n647 & new_n1082;
  assign new_n2187 = new_n2186 ^ n19;
  assign new_n2188 = new_n1224 & new_n1647;
  assign new_n2189 = new_n2188 ^ n275;
  assign new_n2190 = new_n2189 ^ new_n2187;
  assign new_n2191 = new_n648 & new_n1082;
  assign new_n2192 = new_n2191 ^ n18;
  assign new_n2193 = new_n1225 & new_n1647;
  assign new_n2194 = new_n2193 ^ n274;
  assign new_n2195 = new_n2194 ^ new_n2192;
  assign new_n2196 = new_n1226 & new_n1647;
  assign new_n2197 = new_n2196 ^ n273;
  assign new_n2198 = new_n649 & new_n1082;
  assign new_n2199 = new_n2198 ^ n17;
  assign new_n2200 = new_n2199 ^ new_n2197;
  assign new_n2201 = new_n650 & new_n1082;
  assign new_n2202 = new_n2201 ^ n16;
  assign new_n2203 = new_n1227 & new_n1647;
  assign new_n2204 = new_n2203 ^ n272;
  assign new_n2205 = new_n2204 ^ new_n2202;
  assign new_n2206 = new_n651 & new_n1082;
  assign new_n2207 = new_n2206 ^ n15;
  assign new_n2208 = new_n1228 & new_n1647;
  assign new_n2209 = new_n2208 ^ n271;
  assign new_n2210 = new_n2209 ^ new_n2207;
  assign new_n2211 = new_n1229 & new_n1647;
  assign new_n2212 = new_n2211 ^ n270;
  assign new_n2213 = new_n652 & new_n1082;
  assign new_n2214 = new_n2213 ^ n14;
  assign new_n2215 = new_n2214 ^ new_n2212;
  assign new_n2216 = new_n1230 & new_n1647;
  assign new_n2217 = new_n2216 ^ n269;
  assign new_n2218 = new_n653 & new_n1082;
  assign new_n2219 = new_n2218 ^ n13;
  assign new_n2220 = new_n2219 ^ new_n2217;
  assign new_n2221 = new_n654 & new_n1082;
  assign new_n2222 = new_n2221 ^ n12;
  assign new_n2223 = new_n1231 & new_n1647;
  assign new_n2224 = new_n2223 ^ n268;
  assign new_n2225 = new_n2224 ^ new_n2222;
  assign new_n2226 = new_n1232 & new_n1647;
  assign new_n2227 = new_n2226 ^ n267;
  assign new_n2228 = new_n655 & new_n1082;
  assign new_n2229 = new_n2228 ^ n11;
  assign new_n2230 = new_n2229 ^ new_n2227;
  assign new_n2231 = new_n1233 & new_n1647;
  assign new_n2232 = new_n2231 ^ n266;
  assign new_n2233 = new_n656 & new_n1082;
  assign new_n2234 = new_n2233 ^ n10;
  assign new_n2235 = new_n2234 ^ new_n2232;
  assign new_n2236 = new_n1234 & new_n1647;
  assign new_n2237 = new_n2236 ^ n265;
  assign new_n2238 = new_n657 & new_n1082;
  assign new_n2239 = new_n2238 ^ n9;
  assign new_n2240 = new_n2239 ^ new_n2237;
  assign new_n2241 = new_n658 & new_n1082;
  assign new_n2242 = new_n2241 ^ n8;
  assign new_n2243 = new_n1235 & new_n1647;
  assign new_n2244 = new_n2243 ^ n264;
  assign new_n2245 = new_n2244 ^ new_n2242;
  assign new_n2246 = new_n1236 & new_n1647;
  assign new_n2247 = new_n2246 ^ n263;
  assign new_n2248 = new_n659 & new_n1082;
  assign new_n2249 = new_n2248 ^ n7;
  assign new_n2250 = new_n2249 ^ new_n2247;
  assign new_n2251 = new_n660 & new_n1082;
  assign new_n2252 = new_n2251 ^ n6;
  assign new_n2253 = new_n1237 & new_n1647;
  assign new_n2254 = new_n2253 ^ n262;
  assign new_n2255 = new_n2254 ^ new_n2252;
  assign new_n2256 = new_n661 & new_n1082;
  assign new_n2257 = new_n2256 ^ n5;
  assign new_n2258 = new_n1238 & new_n1647;
  assign new_n2259 = new_n2258 ^ n261;
  assign new_n2260 = new_n2259 ^ new_n2257;
  assign new_n2261 = new_n662 & new_n1082;
  assign new_n2262 = new_n2261 ^ n4;
  assign new_n2263 = new_n1239 & new_n1647;
  assign new_n2264 = new_n2263 ^ n260;
  assign new_n2265 = new_n2264 ^ new_n2262;
  assign new_n2266 = new_n1240 & new_n1647;
  assign new_n2267 = new_n2266 ^ n259;
  assign new_n2268 = new_n663 & new_n1082;
  assign new_n2269 = new_n2268 ^ n3;
  assign new_n2270 = new_n2269 ^ new_n2267;
  assign new_n2271 = new_n1241 & new_n1647;
  assign new_n2272 = new_n2271 ^ n258;
  assign new_n2273 = new_n664 & new_n1082;
  assign new_n2274 = new_n2273 ^ n2;
  assign new_n2275 = new_n2274 ^ new_n2272;
  assign new_n2276 = n385 ^ n257;
  assign new_n2277 = new_n1647 & new_n2276;
  assign new_n2278 = new_n2277 ^ n257;
  assign new_n2279 = n129 ^ n1;
  assign new_n2280 = new_n1082 & new_n2279;
  assign new_n2281 = new_n2280 ^ n1;
  assign new_n2282 = ~new_n2278 & new_n2281;
  assign new_n2283 = new_n2282 ^ new_n2274;
  assign new_n2284 = ~new_n2275 & new_n2283;
  assign new_n2285 = new_n2284 ^ new_n2274;
  assign new_n2286 = new_n2285 ^ new_n2269;
  assign new_n2287 = ~new_n2270 & new_n2286;
  assign new_n2288 = new_n2287 ^ new_n2269;
  assign new_n2289 = new_n2288 ^ new_n2262;
  assign new_n2290 = ~new_n2265 & ~new_n2289;
  assign new_n2291 = new_n2290 ^ new_n2264;
  assign new_n2292 = new_n2291 ^ new_n2259;
  assign new_n2293 = ~new_n2260 & ~new_n2292;
  assign new_n2294 = new_n2293 ^ new_n2257;
  assign new_n2295 = new_n2294 ^ new_n2254;
  assign new_n2296 = ~new_n2255 & ~new_n2295;
  assign new_n2297 = new_n2296 ^ new_n2254;
  assign new_n2298 = new_n2297 ^ new_n2249;
  assign new_n2299 = ~new_n2250 & new_n2298;
  assign new_n2300 = new_n2299 ^ new_n2247;
  assign new_n2301 = new_n2300 ^ new_n2244;
  assign new_n2302 = ~new_n2245 & ~new_n2301;
  assign new_n2303 = new_n2302 ^ new_n2242;
  assign new_n2304 = new_n2303 ^ new_n2239;
  assign new_n2305 = ~new_n2240 & new_n2304;
  assign new_n2306 = new_n2305 ^ new_n2239;
  assign new_n2307 = new_n2306 ^ new_n2234;
  assign new_n2308 = ~new_n2235 & new_n2307;
  assign new_n2309 = new_n2308 ^ new_n2234;
  assign new_n2310 = new_n2309 ^ new_n2227;
  assign new_n2311 = ~new_n2230 & ~new_n2310;
  assign new_n2312 = new_n2311 ^ new_n2227;
  assign new_n2313 = new_n2312 ^ new_n2224;
  assign new_n2314 = ~new_n2225 & new_n2313;
  assign new_n2315 = new_n2314 ^ new_n2224;
  assign new_n2316 = new_n2315 ^ new_n2217;
  assign new_n2317 = ~new_n2220 & new_n2316;
  assign new_n2318 = new_n2317 ^ new_n2217;
  assign new_n2319 = new_n2318 ^ new_n2214;
  assign new_n2320 = ~new_n2215 & ~new_n2319;
  assign new_n2321 = new_n2320 ^ new_n2214;
  assign new_n2322 = new_n2321 ^ new_n2207;
  assign new_n2323 = ~new_n2210 & ~new_n2322;
  assign new_n2324 = new_n2323 ^ new_n2209;
  assign new_n2325 = new_n2324 ^ new_n2204;
  assign new_n2326 = ~new_n2205 & ~new_n2325;
  assign new_n2327 = new_n2326 ^ new_n2202;
  assign new_n2328 = new_n2327 ^ new_n2199;
  assign new_n2329 = ~new_n2200 & new_n2328;
  assign new_n2330 = new_n2329 ^ new_n2199;
  assign new_n2331 = new_n2330 ^ new_n2194;
  assign new_n2332 = ~new_n2195 & new_n2331;
  assign new_n2333 = new_n2332 ^ new_n2192;
  assign new_n2334 = new_n2333 ^ new_n2189;
  assign new_n2335 = ~new_n2190 & ~new_n2334;
  assign new_n2336 = new_n2335 ^ new_n2189;
  assign new_n2337 = new_n2336 ^ new_n2184;
  assign new_n2338 = ~new_n2185 & new_n2337;
  assign new_n2339 = new_n2338 ^ new_n2182;
  assign new_n2340 = new_n2339 ^ new_n2179;
  assign new_n2341 = ~new_n2180 & ~new_n2340;
  assign new_n2342 = new_n2341 ^ new_n2177;
  assign new_n2343 = new_n2342 ^ new_n2174;
  assign new_n2344 = ~new_n2175 & new_n2343;
  assign new_n2345 = new_n2344 ^ new_n2174;
  assign new_n2346 = new_n2345 ^ new_n2169;
  assign new_n2347 = ~new_n2170 & new_n2346;
  assign new_n2348 = new_n2347 ^ new_n2169;
  assign new_n2349 = new_n2348 ^ new_n2162;
  assign new_n2350 = ~new_n2165 & ~new_n2349;
  assign new_n2351 = new_n2350 ^ new_n2164;
  assign new_n2352 = new_n2351 ^ new_n2159;
  assign new_n2353 = ~new_n2160 & ~new_n2352;
  assign new_n2354 = new_n2353 ^ new_n2157;
  assign new_n2355 = new_n2354 ^ new_n2154;
  assign new_n2356 = ~new_n2155 & ~new_n2355;
  assign new_n2357 = new_n2356 ^ new_n2154;
  assign new_n2358 = new_n2357 ^ new_n2149;
  assign new_n2359 = ~new_n2150 & ~new_n2358;
  assign new_n2360 = new_n2359 ^ new_n2147;
  assign new_n2361 = new_n2360 ^ new_n2144;
  assign new_n2362 = ~new_n2145 & new_n2361;
  assign new_n2363 = new_n2362 ^ new_n2144;
  assign new_n2364 = new_n2363 ^ new_n2139;
  assign new_n2365 = ~new_n2140 & new_n2364;
  assign new_n2366 = new_n2365 ^ new_n2137;
  assign new_n2367 = new_n2366 ^ new_n2134;
  assign new_n2368 = ~new_n2135 & new_n2367;
  assign new_n2369 = new_n2368 ^ new_n2132;
  assign new_n2370 = new_n2369 ^ new_n2129;
  assign new_n2371 = ~new_n2130 & new_n2370;
  assign new_n2372 = new_n2371 ^ new_n2129;
  assign new_n2373 = new_n2372 ^ new_n2124;
  assign new_n2374 = ~new_n2125 & new_n2373;
  assign new_n2375 = new_n2374 ^ new_n2122;
  assign new_n2376 = new_n2375 ^ new_n2119;
  assign new_n2377 = ~new_n2120 & ~new_n2376;
  assign new_n2378 = new_n2377 ^ new_n2119;
  assign new_n2379 = new_n2378 ^ new_n2114;
  assign new_n2380 = ~new_n2115 & ~new_n2379;
  assign new_n2381 = new_n2380 ^ new_n2112;
  assign new_n2382 = new_n2381 ^ new_n2109;
  assign new_n2383 = ~new_n2110 & new_n2382;
  assign new_n2384 = new_n2383 ^ new_n2109;
  assign new_n2385 = new_n2384 ^ new_n2102;
  assign new_n2386 = ~new_n2105 & new_n2385;
  assign new_n2387 = new_n2386 ^ new_n2104;
  assign new_n2388 = new_n2387 ^ new_n2099;
  assign new_n2389 = ~new_n2100 & new_n2388;
  assign new_n2390 = new_n2389 ^ new_n2097;
  assign new_n2391 = new_n2390 ^ new_n2094;
  assign new_n2392 = ~new_n2095 & new_n2391;
  assign new_n2393 = new_n2392 ^ new_n2094;
  assign new_n2394 = new_n2393 ^ new_n2089;
  assign new_n2395 = ~new_n2090 & new_n2394;
  assign new_n2396 = new_n2395 ^ new_n2087;
  assign new_n2397 = new_n2396 ^ new_n2084;
  assign new_n2398 = ~new_n2085 & ~new_n2397;
  assign new_n2399 = new_n2398 ^ new_n2084;
  assign new_n2400 = new_n2399 ^ new_n2079;
  assign new_n2401 = ~new_n2080 & ~new_n2400;
  assign new_n2402 = new_n2401 ^ new_n2077;
  assign new_n2403 = new_n2402 ^ new_n2074;
  assign new_n2404 = ~new_n2075 & new_n2403;
  assign new_n2405 = new_n2404 ^ new_n2072;
  assign new_n2406 = new_n2405 ^ new_n2069;
  assign new_n2407 = ~new_n2070 & ~new_n2406;
  assign new_n2408 = new_n2407 ^ new_n2069;
  assign new_n2409 = new_n2408 ^ new_n2064;
  assign new_n2410 = ~new_n2065 & ~new_n2409;
  assign new_n2411 = new_n2410 ^ new_n2064;
  assign new_n2412 = new_n2411 ^ new_n2057;
  assign new_n2413 = ~new_n2060 & ~new_n2412;
  assign new_n2414 = new_n2413 ^ new_n2059;
  assign new_n2415 = new_n2414 ^ new_n2054;
  assign new_n2416 = ~new_n2055 & ~new_n2415;
  assign new_n2417 = new_n2416 ^ new_n2052;
  assign new_n2418 = new_n2417 ^ new_n2049;
  assign new_n2419 = ~new_n2050 & ~new_n2418;
  assign new_n2420 = new_n2419 ^ new_n2049;
  assign new_n2421 = new_n2420 ^ new_n2044;
  assign new_n2422 = ~new_n2045 & ~new_n2421;
  assign new_n2423 = new_n2422 ^ new_n2042;
  assign new_n2424 = new_n2423 ^ new_n2039;
  assign new_n2425 = ~new_n2040 & new_n2424;
  assign new_n2426 = new_n2425 ^ new_n2039;
  assign new_n2427 = new_n2426 ^ new_n2034;
  assign new_n2428 = ~new_n2035 & ~new_n2427;
  assign new_n2429 = new_n2428 ^ new_n2034;
  assign new_n2430 = new_n2429 ^ new_n2027;
  assign new_n2431 = ~new_n2030 & ~new_n2430;
  assign new_n2432 = new_n2431 ^ new_n2027;
  assign new_n2433 = new_n2432 ^ new_n2024;
  assign new_n2434 = ~new_n2025 & ~new_n2433;
  assign new_n2435 = new_n2434 ^ new_n2022;
  assign new_n2436 = new_n2435 ^ new_n2019;
  assign new_n2437 = ~new_n2020 & ~new_n2436;
  assign new_n2438 = new_n2437 ^ new_n2017;
  assign new_n2439 = new_n2438 ^ new_n2014;
  assign new_n2440 = ~new_n2015 & new_n2439;
  assign new_n2441 = new_n2440 ^ new_n2014;
  assign new_n2442 = new_n2441 ^ new_n2009;
  assign new_n2443 = ~new_n2010 & ~new_n2442;
  assign new_n2444 = new_n2443 ^ new_n2009;
  assign new_n2445 = new_n2444 ^ new_n2002;
  assign new_n2446 = ~new_n2005 & new_n2445;
  assign new_n2447 = new_n2446 ^ new_n2004;
  assign new_n2448 = new_n2447 ^ new_n1999;
  assign new_n2449 = ~new_n2000 & ~new_n2448;
  assign new_n2450 = new_n2449 ^ new_n1997;
  assign new_n2451 = new_n2450 ^ new_n1994;
  assign new_n2452 = ~new_n1995 & new_n2451;
  assign new_n2453 = new_n2452 ^ new_n1994;
  assign new_n2454 = new_n2453 ^ new_n1989;
  assign new_n2455 = ~new_n1990 & new_n2454;
  assign new_n2456 = new_n2455 ^ new_n1989;
  assign new_n2457 = new_n2456 ^ new_n1982;
  assign new_n2458 = ~new_n1985 & new_n2457;
  assign new_n2459 = new_n2458 ^ new_n1982;
  assign new_n2460 = new_n2459 ^ new_n1979;
  assign new_n2461 = ~new_n1980 & ~new_n2460;
  assign new_n2462 = new_n2461 ^ new_n1979;
  assign new_n2463 = new_n2462 ^ new_n1972;
  assign new_n2464 = ~new_n1975 & ~new_n2463;
  assign new_n2465 = new_n2464 ^ new_n1972;
  assign new_n2466 = new_n2465 ^ new_n1969;
  assign new_n2467 = ~new_n1970 & ~new_n2466;
  assign new_n2468 = new_n2467 ^ new_n1969;
  assign new_n2469 = new_n2468 ^ new_n1962;
  assign new_n2470 = ~new_n1965 & new_n2469;
  assign new_n2471 = new_n2470 ^ new_n1962;
  assign new_n2472 = new_n2471 ^ new_n1959;
  assign new_n2473 = ~new_n1960 & new_n2472;
  assign new_n2474 = new_n2473 ^ new_n1959;
  assign new_n2475 = new_n2474 ^ new_n1952;
  assign new_n2476 = ~new_n1955 & new_n2475;
  assign new_n2477 = new_n2476 ^ new_n1952;
  assign new_n2478 = new_n2477 ^ new_n1949;
  assign new_n2479 = ~new_n1950 & ~new_n2478;
  assign new_n2480 = new_n2479 ^ new_n1947;
  assign new_n2481 = new_n2480 ^ new_n1944;
  assign new_n2482 = ~new_n1945 & new_n2481;
  assign new_n2483 = new_n2482 ^ new_n1942;
  assign new_n2484 = new_n2483 ^ new_n1939;
  assign new_n2485 = ~new_n1940 & new_n2484;
  assign new_n2486 = new_n2485 ^ new_n1939;
  assign new_n2487 = new_n2486 ^ new_n1934;
  assign new_n2488 = ~new_n1935 & ~new_n2487;
  assign new_n2489 = new_n2488 ^ new_n1934;
  assign new_n2490 = new_n2489 ^ new_n1927;
  assign new_n2491 = ~new_n1930 & ~new_n2490;
  assign new_n2492 = new_n2491 ^ new_n1929;
  assign new_n2493 = new_n2492 ^ new_n1924;
  assign new_n2494 = ~new_n1925 & new_n2493;
  assign new_n2495 = new_n2494 ^ new_n1922;
  assign new_n2496 = new_n2495 ^ new_n1919;
  assign new_n2497 = ~new_n1920 & ~new_n2496;
  assign new_n2498 = new_n2497 ^ new_n1919;
  assign new_n2499 = new_n2498 ^ new_n1914;
  assign new_n2500 = ~new_n1915 & ~new_n2499;
  assign new_n2501 = new_n2500 ^ new_n1914;
  assign new_n2502 = new_n2501 ^ new_n1909;
  assign new_n2503 = ~new_n1910 & new_n2502;
  assign new_n2504 = new_n2503 ^ new_n1909;
  assign new_n2505 = new_n2504 ^ new_n1902;
  assign new_n2506 = ~new_n1905 & ~new_n2505;
  assign new_n2507 = new_n2506 ^ new_n1902;
  assign new_n2508 = new_n2507 ^ new_n1899;
  assign new_n2509 = ~new_n1900 & ~new_n2508;
  assign new_n2510 = new_n2509 ^ new_n1899;
  assign new_n2511 = new_n2510 ^ new_n1892;
  assign new_n2512 = ~new_n1895 & ~new_n2511;
  assign new_n2513 = new_n2512 ^ new_n1894;
  assign new_n2514 = new_n2513 ^ new_n1889;
  assign new_n2515 = ~new_n1890 & new_n2514;
  assign new_n2516 = new_n2515 ^ new_n1887;
  assign new_n2517 = new_n2516 ^ new_n1882;
  assign new_n2518 = ~new_n1885 & ~new_n2517;
  assign new_n2519 = new_n2518 ^ new_n1882;
  assign new_n2520 = new_n2519 ^ new_n1879;
  assign new_n2521 = ~new_n1880 & new_n2520;
  assign new_n2522 = new_n2521 ^ new_n1877;
  assign new_n2523 = new_n2522 ^ new_n1874;
  assign new_n2524 = ~new_n1875 & new_n2523;
  assign new_n2525 = new_n2524 ^ new_n1872;
  assign new_n2526 = new_n2525 ^ new_n1867;
  assign new_n2527 = ~new_n1870 & ~new_n2526;
  assign new_n2528 = new_n2527 ^ new_n1867;
  assign new_n2529 = new_n2528 ^ new_n1862;
  assign new_n2530 = ~new_n1865 & ~new_n2529;
  assign new_n2531 = new_n2530 ^ new_n1862;
  assign new_n2532 = new_n2531 ^ new_n1859;
  assign new_n2533 = ~new_n1860 & new_n2532;
  assign new_n2534 = new_n2533 ^ new_n1859;
  assign new_n2535 = new_n2534 ^ new_n1852;
  assign new_n2536 = ~new_n1855 & new_n2535;
  assign new_n2537 = new_n2536 ^ new_n1852;
  assign new_n2538 = new_n2537 ^ new_n1847;
  assign new_n2539 = ~new_n1850 & new_n2538;
  assign new_n2540 = new_n2539 ^ new_n1847;
  assign new_n2541 = new_n2540 ^ new_n1842;
  assign new_n2542 = ~new_n1845 & new_n2541;
  assign new_n2543 = new_n2542 ^ new_n1842;
  assign new_n2544 = new_n2543 ^ new_n1839;
  assign new_n2545 = ~new_n1840 & ~new_n2544;
  assign new_n2546 = new_n2545 ^ new_n1839;
  assign new_n2547 = new_n2546 ^ new_n1832;
  assign new_n2548 = ~new_n1835 & new_n2547;
  assign new_n2549 = new_n2548 ^ new_n1832;
  assign new_n2550 = new_n2549 ^ new_n1829;
  assign new_n2551 = ~new_n1830 & new_n2550;
  assign new_n2552 = new_n2551 ^ new_n1829;
  assign new_n2553 = new_n2552 ^ new_n1822;
  assign new_n2554 = ~new_n1825 & ~new_n2553;
  assign new_n2555 = new_n2554 ^ new_n1822;
  assign new_n2556 = new_n2555 ^ new_n1817;
  assign new_n2557 = ~new_n1820 & ~new_n2556;
  assign new_n2558 = new_n2557 ^ new_n1819;
  assign new_n2559 = new_n2558 ^ new_n1814;
  assign new_n2560 = ~new_n1815 & new_n2559;
  assign new_n2561 = new_n2560 ^ new_n1812;
  assign new_n2562 = new_n2561 ^ new_n1807;
  assign new_n2563 = ~new_n1810 & new_n2562;
  assign new_n2564 = new_n2563 ^ new_n1807;
  assign new_n2565 = new_n2564 ^ new_n1802;
  assign new_n2566 = ~new_n1805 & new_n2565;
  assign new_n2567 = new_n2566 ^ new_n1802;
  assign new_n2568 = new_n2567 ^ new_n1797;
  assign new_n2569 = ~new_n1800 & ~new_n2568;
  assign new_n2570 = new_n2569 ^ new_n1799;
  assign new_n2571 = new_n2570 ^ new_n1794;
  assign new_n2572 = ~new_n1795 & new_n2571;
  assign new_n2573 = new_n2572 ^ new_n1792;
  assign new_n2574 = new_n2573 ^ new_n1787;
  assign new_n2575 = ~new_n1790 & ~new_n2574;
  assign new_n2576 = new_n2575 ^ new_n1787;
  assign new_n2577 = new_n2576 ^ new_n1782;
  assign new_n2578 = ~new_n1785 & new_n2577;
  assign new_n2579 = new_n2578 ^ new_n1782;
  assign new_n2580 = new_n2579 ^ new_n1779;
  assign new_n2581 = ~new_n1780 & ~new_n2580;
  assign new_n2582 = new_n2581 ^ new_n1777;
  assign new_n2583 = new_n2582 ^ new_n1774;
  assign new_n2584 = ~new_n1775 & new_n2583;
  assign new_n2585 = new_n2584 ^ new_n1772;
  assign new_n2586 = new_n2585 ^ new_n1767;
  assign new_n2587 = ~new_n1770 & ~new_n2586;
  assign new_n2588 = new_n2587 ^ new_n1767;
  assign new_n2589 = new_n2588 ^ new_n1762;
  assign new_n2590 = ~new_n1765 & new_n2589;
  assign new_n2591 = new_n2590 ^ new_n1764;
  assign new_n2592 = new_n2591 ^ new_n1759;
  assign new_n2593 = ~new_n1760 & ~new_n2592;
  assign new_n2594 = new_n2593 ^ new_n1757;
  assign new_n2595 = new_n2594 ^ new_n1752;
  assign new_n2596 = ~new_n1755 & ~new_n2595;
  assign new_n2597 = new_n2596 ^ new_n1752;
  assign new_n2598 = new_n2597 ^ new_n1749;
  assign new_n2599 = ~new_n1750 & new_n2598;
  assign new_n2600 = new_n2599 ^ new_n1747;
  assign new_n2601 = new_n2600 ^ new_n1744;
  assign new_n2602 = ~new_n1745 & new_n2601;
  assign new_n2603 = new_n2602 ^ new_n1742;
  assign new_n2604 = new_n2603 ^ new_n1739;
  assign new_n2605 = ~new_n1740 & new_n2604;
  assign new_n2606 = new_n2605 ^ new_n1739;
  assign new_n2607 = new_n2606 ^ new_n1734;
  assign new_n2608 = ~new_n1735 & ~new_n2607;
  assign new_n2609 = new_n2608 ^ new_n1732;
  assign new_n2610 = new_n2609 ^ new_n1729;
  assign new_n2611 = ~new_n1730 & new_n2610;
  assign new_n2612 = new_n2611 ^ new_n1727;
  assign new_n2613 = new_n2612 ^ new_n1722;
  assign new_n2614 = ~new_n1725 & ~new_n2613;
  assign new_n2615 = new_n2614 ^ new_n1722;
  assign new_n2616 = new_n2615 ^ new_n1717;
  assign new_n2617 = ~new_n1720 & new_n2616;
  assign new_n2618 = new_n2617 ^ new_n1717;
  assign new_n2619 = new_n2618 ^ new_n1714;
  assign new_n2620 = ~new_n1715 & ~new_n2619;
  assign new_n2621 = new_n2620 ^ new_n1714;
  assign new_n2622 = new_n2621 ^ new_n1707;
  assign new_n2623 = ~new_n1710 & ~new_n2622;
  assign new_n2624 = new_n2623 ^ new_n1707;
  assign new_n2625 = new_n2624 ^ new_n1704;
  assign new_n2626 = ~new_n1705 & new_n2625;
  assign new_n2627 = new_n2626 ^ new_n1704;
  assign new_n2628 = new_n2627 ^ new_n1697;
  assign new_n2629 = ~new_n1700 & ~new_n2628;
  assign new_n2630 = new_n2629 ^ new_n1697;
  assign new_n2631 = new_n2630 ^ new_n1694;
  assign new_n2632 = ~new_n1695 & new_n2631;
  assign new_n2633 = new_n2632 ^ new_n1694;
  assign new_n2634 = new_n2633 ^ new_n1689;
  assign new_n2635 = ~new_n1690 & ~new_n2634;
  assign new_n2636 = new_n2635 ^ new_n1687;
  assign new_n2637 = new_n2636 ^ new_n1684;
  assign new_n2638 = ~new_n1685 & new_n2637;
  assign new_n2639 = new_n2638 ^ new_n1682;
  assign new_n2640 = new_n2639 ^ new_n1679;
  assign new_n2641 = ~new_n1680 & new_n2640;
  assign new_n2642 = new_n2641 ^ new_n1679;
  assign new_n2643 = new_n2642 ^ new_n1672;
  assign new_n2644 = ~new_n1675 & ~new_n2643;
  assign new_n2645 = new_n2644 ^ new_n1674;
  assign new_n2646 = new_n2645 ^ new_n1669;
  assign new_n2647 = ~new_n1670 & ~new_n2646;
  assign new_n2648 = new_n2647 ^ new_n1667;
  assign new_n2649 = new_n2648 ^ new_n1662;
  assign new_n2650 = ~new_n1665 & new_n2649;
  assign new_n2651 = new_n2650 ^ new_n1662;
  assign new_n2652 = new_n2651 ^ new_n1657;
  assign new_n2653 = ~new_n1660 & new_n2652;
  assign new_n2654 = new_n2653 ^ new_n1657;
  assign new_n2655 = new_n2654 ^ new_n1654;
  assign new_n2656 = ~new_n1655 & ~new_n2655;
  assign new_n2657 = new_n2656 ^ new_n1654;
  assign new_n2658 = new_n2657 ^ new_n1084;
  assign new_n2659 = ~new_n1650 & ~new_n2658;
  assign new_n2660 = new_n1649 ^ new_n514;
  assign new_n2661 = new_n2660 ^ new_n2659;
  assign new_n2662 = ~new_n515 & new_n2661;
  assign new_n2663 = new_n2662 ^ new_n513;
  assign new_n2664 = new_n2281 ^ new_n2278;
  assign new_n2665 = ~new_n2663 & new_n2664;
  assign new_n2666 = new_n2665 ^ new_n2278;
  assign new_n2667 = ~new_n2663 & new_n2275;
  assign new_n2668 = new_n2667 ^ new_n2272;
  assign new_n2669 = ~new_n2663 & new_n2270;
  assign new_n2670 = new_n2669 ^ new_n2267;
  assign new_n2671 = ~new_n2663 & new_n2265;
  assign new_n2672 = new_n2671 ^ new_n2264;
  assign new_n2673 = new_n2260 & new_n2663;
  assign new_n2674 = new_n2673 ^ new_n2257;
  assign new_n2675 = new_n2255 & new_n2663;
  assign new_n2676 = new_n2675 ^ new_n2252;
  assign new_n2677 = ~new_n2663 & new_n2250;
  assign new_n2678 = new_n2677 ^ new_n2247;
  assign new_n2679 = new_n2245 & new_n2663;
  assign new_n2680 = new_n2679 ^ new_n2242;
  assign new_n2681 = ~new_n2663 & new_n2240;
  assign new_n2682 = new_n2681 ^ new_n2237;
  assign new_n2683 = ~new_n2663 & new_n2235;
  assign new_n2684 = new_n2683 ^ new_n2232;
  assign new_n2685 = new_n2230 & new_n2663;
  assign new_n2686 = new_n2685 ^ new_n2229;
  assign new_n2687 = new_n2225 & new_n2663;
  assign new_n2688 = new_n2687 ^ new_n2222;
  assign new_n2689 = new_n2220 & new_n2663;
  assign new_n2690 = new_n2689 ^ new_n2219;
  assign new_n2691 = ~new_n2663 & new_n2215;
  assign new_n2692 = new_n2691 ^ new_n2212;
  assign new_n2693 = ~new_n2663 & new_n2210;
  assign new_n2694 = new_n2693 ^ new_n2209;
  assign new_n2695 = new_n2205 & new_n2663;
  assign new_n2696 = new_n2695 ^ new_n2202;
  assign new_n2697 = ~new_n2663 & new_n2200;
  assign new_n2698 = new_n2697 ^ new_n2197;
  assign new_n2699 = new_n2195 & new_n2663;
  assign new_n2700 = new_n2699 ^ new_n2192;
  assign new_n2701 = new_n2190 & new_n2663;
  assign new_n2702 = new_n2701 ^ new_n2187;
  assign new_n2703 = ~new_n2663 & new_n2185;
  assign new_n2704 = new_n2703 ^ new_n2182;
  assign new_n2705 = new_n2180 & new_n2663;
  assign new_n2706 = new_n2705 ^ new_n2177;
  assign new_n2707 = ~new_n2663 & new_n2175;
  assign new_n2708 = new_n2707 ^ new_n2172;
  assign new_n2709 = ~new_n2663 & new_n2170;
  assign new_n2710 = new_n2709 ^ new_n2167;
  assign new_n2711 = ~new_n2663 & new_n2165;
  assign new_n2712 = new_n2711 ^ new_n2164;
  assign new_n2713 = new_n2160 & new_n2663;
  assign new_n2714 = new_n2713 ^ new_n2157;
  assign new_n2715 = new_n2155 & new_n2663;
  assign new_n2716 = new_n2715 ^ new_n2152;
  assign new_n2717 = new_n2150 & new_n2663;
  assign new_n2718 = new_n2717 ^ new_n2147;
  assign new_n2719 = ~new_n2663 & new_n2145;
  assign new_n2720 = new_n2719 ^ new_n2142;
  assign new_n2721 = new_n2140 & new_n2663;
  assign new_n2722 = new_n2721 ^ new_n2137;
  assign new_n2723 = new_n2135 & new_n2663;
  assign new_n2724 = new_n2723 ^ new_n2132;
  assign new_n2725 = ~new_n2663 & new_n2130;
  assign new_n2726 = new_n2725 ^ new_n2127;
  assign new_n2727 = new_n2125 & new_n2663;
  assign new_n2728 = new_n2727 ^ new_n2122;
  assign new_n2729 = new_n2120 & new_n2663;
  assign new_n2730 = new_n2729 ^ new_n2117;
  assign new_n2731 = new_n2115 & new_n2663;
  assign new_n2732 = new_n2731 ^ new_n2112;
  assign new_n2733 = ~new_n2663 & new_n2110;
  assign new_n2734 = new_n2733 ^ new_n2107;
  assign new_n2735 = new_n2105 & new_n2663;
  assign new_n2736 = new_n2735 ^ new_n2104;
  assign new_n2737 = new_n2100 & new_n2663;
  assign new_n2738 = new_n2737 ^ new_n2097;
  assign new_n2739 = ~new_n2663 & new_n2095;
  assign new_n2740 = new_n2739 ^ new_n2092;
  assign new_n2741 = new_n2090 & new_n2663;
  assign new_n2742 = new_n2741 ^ new_n2087;
  assign new_n2743 = new_n2085 & new_n2663;
  assign new_n2744 = new_n2743 ^ new_n2082;
  assign new_n2745 = new_n2080 & new_n2663;
  assign new_n2746 = new_n2745 ^ new_n2077;
  assign new_n2747 = new_n2075 & new_n2663;
  assign new_n2748 = new_n2747 ^ new_n2072;
  assign new_n2749 = new_n2070 & new_n2663;
  assign new_n2750 = new_n2749 ^ new_n2067;
  assign new_n2751 = ~new_n2663 & new_n2065;
  assign new_n2752 = new_n2751 ^ new_n2062;
  assign new_n2753 = ~new_n2663 & new_n2060;
  assign new_n2754 = new_n2753 ^ new_n2059;
  assign new_n2755 = new_n2055 & new_n2663;
  assign new_n2756 = new_n2755 ^ new_n2052;
  assign new_n2757 = new_n2050 & new_n2663;
  assign new_n2758 = new_n2757 ^ new_n2047;
  assign new_n2759 = new_n2045 & new_n2663;
  assign new_n2760 = new_n2759 ^ new_n2042;
  assign new_n2761 = ~new_n2663 & new_n2040;
  assign new_n2762 = new_n2761 ^ new_n2037;
  assign new_n2763 = new_n2035 & new_n2663;
  assign new_n2764 = new_n2763 ^ new_n2032;
  assign new_n2765 = ~new_n2663 & new_n2030;
  assign new_n2766 = new_n2765 ^ new_n2029;
  assign new_n2767 = ~new_n2663 & new_n2025;
  assign new_n2768 = new_n2767 ^ new_n2022;
  assign new_n2769 = new_n2020 & new_n2663;
  assign new_n2770 = new_n2769 ^ new_n2017;
  assign new_n2771 = ~new_n2663 & new_n2015;
  assign new_n2772 = new_n2771 ^ new_n2012;
  assign new_n2773 = new_n2010 & new_n2663;
  assign new_n2774 = new_n2773 ^ new_n2007;
  assign new_n2775 = ~new_n2663 & new_n2005;
  assign new_n2776 = new_n2775 ^ new_n2004;
  assign new_n2777 = new_n2000 & new_n2663;
  assign new_n2778 = new_n2777 ^ new_n1997;
  assign new_n2779 = ~new_n2663 & new_n1995;
  assign new_n2780 = new_n2779 ^ new_n1992;
  assign new_n2781 = ~new_n2663 & new_n1990;
  assign new_n2782 = new_n2781 ^ new_n1987;
  assign new_n2783 = ~new_n2663 & new_n1985;
  assign new_n2784 = new_n2783 ^ new_n1984;
  assign new_n2785 = new_n1980 & new_n2663;
  assign new_n2786 = new_n2785 ^ new_n1977;
  assign new_n2787 = ~new_n2663 & new_n1975;
  assign new_n2788 = new_n2787 ^ new_n1974;
  assign new_n2789 = new_n1970 & new_n2663;
  assign new_n2790 = new_n2789 ^ new_n1967;
  assign new_n2791 = new_n1965 & new_n2663;
  assign new_n2792 = new_n2791 ^ new_n1964;
  assign new_n2793 = new_n1960 & new_n2663;
  assign new_n2794 = new_n2793 ^ new_n1957;
  assign new_n2795 = new_n1955 & new_n2663;
  assign new_n2796 = new_n2795 ^ new_n1954;
  assign new_n2797 = new_n1950 & new_n2663;
  assign new_n2798 = new_n2797 ^ new_n1947;
  assign new_n2799 = new_n1945 & new_n2663;
  assign new_n2800 = new_n2799 ^ new_n1942;
  assign new_n2801 = ~new_n2663 & new_n1940;
  assign new_n2802 = new_n2801 ^ new_n1937;
  assign new_n2803 = new_n1935 & new_n2663;
  assign new_n2804 = new_n2803 ^ new_n1932;
  assign new_n2805 = new_n1930 & new_n2663;
  assign new_n2806 = new_n2805 ^ new_n1929;
  assign new_n2807 = new_n1925 & new_n2663;
  assign new_n2808 = new_n2807 ^ new_n1922;
  assign new_n2809 = new_n1920 & new_n2663;
  assign new_n2810 = new_n2809 ^ new_n1917;
  assign new_n2811 = ~new_n2663 & new_n1915;
  assign new_n2812 = new_n2811 ^ new_n1912;
  assign new_n2813 = new_n1910 & new_n2663;
  assign new_n2814 = new_n2813 ^ new_n1909;
  assign new_n2815 = ~new_n2663 & new_n1905;
  assign new_n2816 = new_n2815 ^ new_n1902;
  assign new_n2817 = new_n1900 & new_n2663;
  assign new_n2818 = new_n2817 ^ new_n1899;
  assign new_n2819 = ~new_n2663 & new_n1895;
  assign new_n2820 = new_n2819 ^ new_n1894;
  assign new_n2821 = ~new_n2663 & new_n1890;
  assign new_n2822 = new_n2821 ^ new_n1887;
  assign new_n2823 = new_n1885 & new_n2663;
  assign new_n2824 = new_n2823 ^ new_n1882;
  assign new_n2825 = new_n1880 & new_n2663;
  assign new_n2826 = new_n2825 ^ new_n1877;
  assign new_n2827 = new_n1875 & new_n2663;
  assign new_n2828 = new_n2827 ^ new_n1872;
  assign new_n2829 = ~new_n2663 & new_n1870;
  assign new_n2830 = new_n2829 ^ new_n1867;
  assign new_n2831 = new_n1865 & new_n2663;
  assign new_n2832 = new_n2831 ^ new_n1862;
  assign new_n2833 = new_n1860 & new_n2663;
  assign new_n2834 = new_n2833 ^ new_n1859;
  assign new_n2835 = new_n1855 & new_n2663;
  assign new_n2836 = new_n2835 ^ new_n1852;
  assign new_n2837 = ~new_n2663 & new_n1850;
  assign new_n2838 = new_n2837 ^ new_n1849;
  assign new_n2839 = new_n1845 & new_n2663;
  assign new_n2840 = new_n2839 ^ new_n1842;
  assign new_n2841 = ~new_n2663 & new_n1840;
  assign new_n2842 = new_n2841 ^ new_n1839;
  assign new_n2843 = ~new_n2663 & new_n1835;
  assign new_n2844 = new_n2843 ^ new_n1832;
  assign new_n2845 = ~new_n2663 & new_n1830;
  assign new_n2846 = new_n2845 ^ new_n1829;
  assign new_n2847 = new_n1825 & new_n2663;
  assign new_n2848 = new_n2847 ^ new_n1822;
  assign new_n2849 = ~new_n2663 & new_n1820;
  assign new_n2850 = new_n2849 ^ new_n1819;
  assign new_n2851 = ~new_n2663 & new_n1815;
  assign new_n2852 = new_n2851 ^ new_n1812;
  assign new_n2853 = ~new_n2663 & new_n1810;
  assign new_n2854 = new_n2853 ^ new_n1807;
  assign new_n2855 = ~new_n2663 & new_n1805;
  assign new_n2856 = new_n2855 ^ new_n1802;
  assign new_n2857 = new_n1800 & new_n2663;
  assign new_n2858 = new_n2857 ^ new_n1799;
  assign new_n2859 = new_n1795 & new_n2663;
  assign new_n2860 = new_n2859 ^ new_n1792;
  assign new_n2861 = ~new_n2663 & new_n1790;
  assign new_n2862 = new_n2861 ^ new_n1787;
  assign new_n2863 = ~new_n2663 & new_n1785;
  assign new_n2864 = new_n2863 ^ new_n1782;
  assign new_n2865 = new_n1780 & new_n2663;
  assign new_n2866 = new_n2865 ^ new_n1777;
  assign new_n2867 = new_n1775 & new_n2663;
  assign new_n2868 = new_n2867 ^ new_n1772;
  assign new_n2869 = ~new_n2663 & new_n1770;
  assign new_n2870 = new_n2869 ^ new_n1767;
  assign new_n2871 = ~new_n2663 & new_n1765;
  assign new_n2872 = new_n2871 ^ new_n1764;
  assign new_n2873 = new_n1760 & new_n2663;
  assign new_n2874 = new_n2873 ^ new_n1757;
  assign new_n2875 = ~new_n2663 & new_n1755;
  assign new_n2876 = new_n2875 ^ new_n1752;
  assign new_n2877 = ~new_n2663 & new_n1750;
  assign new_n2878 = new_n2877 ^ new_n1747;
  assign new_n2879 = ~new_n2663 & new_n1745;
  assign new_n2880 = new_n2879 ^ new_n1742;
  assign new_n2881 = new_n1740 & new_n2663;
  assign new_n2882 = new_n2881 ^ new_n1737;
  assign new_n2883 = new_n1735 & new_n2663;
  assign new_n2884 = new_n2883 ^ new_n1732;
  assign new_n2885 = new_n1730 & new_n2663;
  assign new_n2886 = new_n2885 ^ new_n1727;
  assign new_n2887 = ~new_n2663 & new_n1725;
  assign new_n2888 = new_n2887 ^ new_n1722;
  assign new_n2889 = ~new_n2663 & new_n1720;
  assign new_n2890 = new_n2889 ^ new_n1717;
  assign new_n2891 = new_n1715 & new_n2663;
  assign new_n2892 = new_n2891 ^ new_n1714;
  assign new_n2893 = ~new_n2663 & new_n1710;
  assign new_n2894 = new_n2893 ^ new_n1707;
  assign new_n2895 = ~new_n2663 & new_n1705;
  assign new_n2896 = new_n2895 ^ new_n1704;
  assign new_n2897 = new_n1700 & new_n2663;
  assign new_n2898 = new_n2897 ^ new_n1697;
  assign new_n2899 = new_n1695 & new_n2663;
  assign new_n2900 = new_n2899 ^ new_n1694;
  assign new_n2901 = ~new_n2663 & new_n1690;
  assign new_n2902 = new_n2901 ^ new_n1687;
  assign new_n2903 = ~new_n2663 & new_n1685;
  assign new_n2904 = new_n2903 ^ new_n1682;
  assign new_n2905 = new_n1680 & new_n2663;
  assign new_n2906 = new_n2905 ^ new_n1677;
  assign new_n2907 = new_n1675 & new_n2663;
  assign new_n2908 = new_n2907 ^ new_n1674;
  assign new_n2909 = ~new_n2663 & new_n1670;
  assign new_n2910 = new_n2909 ^ new_n1667;
  assign new_n2911 = ~new_n2663 & new_n1665;
  assign new_n2912 = new_n2911 ^ new_n1662;
  assign new_n2913 = ~new_n2663 & new_n1660;
  assign new_n2914 = new_n2913 ^ new_n1657;
  assign new_n2915 = new_n1655 & new_n2663;
  assign new_n2916 = new_n2915 ^ new_n1654;
  assign new_n2917 = ~new_n2663 & new_n1650;
  assign new_n2918 = new_n2917 ^ new_n1649;
  assign new_n2919 = new_n513 & new_n514;
  assign new_n2920 = new_n1647 ^ new_n1082;
  assign new_n2921 = ~new_n2663 & new_n2920;
  assign new_n2922 = new_n2921 ^ new_n1647;
  assign po0 = new_n2666;
  assign po1 = new_n2668;
  assign po2 = new_n2670;
  assign po3 = new_n2672;
  assign po4 = new_n2674;
  assign po5 = new_n2676;
  assign po6 = new_n2678;
  assign po7 = new_n2680;
  assign po8 = new_n2682;
  assign po9 = new_n2684;
  assign po10 = new_n2686;
  assign po11 = new_n2688;
  assign po12 = new_n2690;
  assign po13 = new_n2692;
  assign po14 = new_n2694;
  assign po15 = new_n2696;
  assign po16 = new_n2698;
  assign po17 = new_n2700;
  assign po18 = new_n2702;
  assign po19 = new_n2704;
  assign po20 = new_n2706;
  assign po21 = new_n2708;
  assign po22 = new_n2710;
  assign po23 = new_n2712;
  assign po24 = new_n2714;
  assign po25 = new_n2716;
  assign po26 = new_n2718;
  assign po27 = new_n2720;
  assign po28 = new_n2722;
  assign po29 = new_n2724;
  assign po30 = new_n2726;
  assign po31 = new_n2728;
  assign po32 = new_n2730;
  assign po33 = new_n2732;
  assign po34 = new_n2734;
  assign po35 = new_n2736;
  assign po36 = new_n2738;
  assign po37 = new_n2740;
  assign po38 = new_n2742;
  assign po39 = new_n2744;
  assign po40 = new_n2746;
  assign po41 = new_n2748;
  assign po42 = new_n2750;
  assign po43 = new_n2752;
  assign po44 = new_n2754;
  assign po45 = new_n2756;
  assign po46 = new_n2758;
  assign po47 = new_n2760;
  assign po48 = new_n2762;
  assign po49 = new_n2764;
  assign po50 = new_n2766;
  assign po51 = new_n2768;
  assign po52 = new_n2770;
  assign po53 = new_n2772;
  assign po54 = new_n2774;
  assign po55 = new_n2776;
  assign po56 = new_n2778;
  assign po57 = new_n2780;
  assign po58 = new_n2782;
  assign po59 = new_n2784;
  assign po60 = new_n2786;
  assign po61 = new_n2788;
  assign po62 = new_n2790;
  assign po63 = new_n2792;
  assign po64 = new_n2794;
  assign po65 = new_n2796;
  assign po66 = new_n2798;
  assign po67 = new_n2800;
  assign po68 = new_n2802;
  assign po69 = new_n2804;
  assign po70 = new_n2806;
  assign po71 = new_n2808;
  assign po72 = new_n2810;
  assign po73 = new_n2812;
  assign po74 = new_n2814;
  assign po75 = new_n2816;
  assign po76 = new_n2818;
  assign po77 = new_n2820;
  assign po78 = new_n2822;
  assign po79 = new_n2824;
  assign po80 = new_n2826;
  assign po81 = new_n2828;
  assign po82 = new_n2830;
  assign po83 = new_n2832;
  assign po84 = new_n2834;
  assign po85 = new_n2836;
  assign po86 = new_n2838;
  assign po87 = new_n2840;
  assign po88 = new_n2842;
  assign po89 = new_n2844;
  assign po90 = new_n2846;
  assign po91 = new_n2848;
  assign po92 = new_n2850;
  assign po93 = new_n2852;
  assign po94 = new_n2854;
  assign po95 = new_n2856;
  assign po96 = new_n2858;
  assign po97 = new_n2860;
  assign po98 = new_n2862;
  assign po99 = new_n2864;
  assign po100 = new_n2866;
  assign po101 = new_n2868;
  assign po102 = new_n2870;
  assign po103 = new_n2872;
  assign po104 = new_n2874;
  assign po105 = new_n2876;
  assign po106 = new_n2878;
  assign po107 = new_n2880;
  assign po108 = new_n2882;
  assign po109 = new_n2884;
  assign po110 = new_n2886;
  assign po111 = new_n2888;
  assign po112 = new_n2890;
  assign po113 = new_n2892;
  assign po114 = new_n2894;
  assign po115 = new_n2896;
  assign po116 = new_n2898;
  assign po117 = new_n2900;
  assign po118 = new_n2902;
  assign po119 = new_n2904;
  assign po120 = new_n2906;
  assign po121 = new_n2908;
  assign po122 = new_n2910;
  assign po123 = new_n2912;
  assign po124 = new_n2914;
  assign po125 = new_n2916;
  assign po126 = new_n2918;
  assign po127 = new_n2919;
  assign po128 = new_n2922;
  assign po129 = new_n2663;
endmodule


