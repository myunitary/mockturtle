module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n9 = x0 & x1 ;
  assign n10 = n9 ^ x0 ;
  assign n11 = x2 & n10 ;
  assign n12 = x2 ^ x0 ;
  assign n13 = x1 & n12 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = x3 & n16 ;
  assign n18 = x4 ^ x2 ;
  assign n19 = x3 & n18 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n16 & n22 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n16 ;
  assign n26 = x4 & n25 ;
  assign n27 = x5 & n25 ;
  assign n28 = x6 & n16 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = x4 & x5 ;
  assign n31 = n30 ^ x4 ;
  assign n32 = n22 & n31 ;
  assign n33 = n32 ^ n22 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n29 & ~n34 ;
  assign n36 = n35 ^ x6 ;
  assign n38 = n31 ^ x5 ;
  assign n37 = x5 & x6 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = x7 & ~n39 ;
  assign n41 = n25 & n40 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n42 ^ x7 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = n11 ;
  assign y3 = n17 ;
  assign y4 = n26 ;
  assign y5 = n27 ;
  assign y6 = n36 ;
  assign y7 = n43 ;
endmodule
