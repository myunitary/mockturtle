// Benchmark "/tmp/tmp" written by ABC on Wed Nov 12 17:26:00 2025

module aes_1cc_firstframe ( 
    n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
    n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127  );
  input  n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
    n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
    n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127;
  wire new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1456, new_n1457, new_n1458, new_n1459, new_n1460,
    new_n1461, new_n1462, new_n1463, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1469, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1474, new_n1475, new_n1476, new_n1477, new_n1478,
    new_n1479, new_n1480, new_n1481, new_n1482, new_n1483, new_n1484,
    new_n1485, new_n1486, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1557, new_n1558, new_n1559, new_n1560, new_n1561, new_n1562,
    new_n1563, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1580,
    new_n1581, new_n1582, new_n1583, new_n1584, new_n1585, new_n1586,
    new_n1587, new_n1588, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1692, new_n1693, new_n1694,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1725, new_n1726, new_n1727, new_n1728, new_n1729, new_n1730,
    new_n1731, new_n1732, new_n1733, new_n1734, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1746, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1775, new_n1776, new_n1777, new_n1778,
    new_n1779, new_n1780, new_n1781, new_n1782, new_n1783, new_n1784,
    new_n1785, new_n1786, new_n1787, new_n1788, new_n1789, new_n1790,
    new_n1791, new_n1792, new_n1793, new_n1794, new_n1795, new_n1796,
    new_n1797, new_n1798, new_n1799, new_n1800, new_n1801, new_n1802,
    new_n1803, new_n1804, new_n1805, new_n1806, new_n1807, new_n1808,
    new_n1809, new_n1810, new_n1811, new_n1812, new_n1813, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1818, new_n1819, new_n1820,
    new_n1821, new_n1822, new_n1823, new_n1824, new_n1825, new_n1826,
    new_n1827, new_n1828, new_n1829, new_n1830, new_n1831, new_n1832,
    new_n1833, new_n1834, new_n1835, new_n1836, new_n1837, new_n1838,
    new_n1839, new_n1840, new_n1841, new_n1842, new_n1843, new_n1844,
    new_n1845, new_n1846, new_n1847, new_n1848, new_n1849, new_n1850,
    new_n1851, new_n1852, new_n1853, new_n1854, new_n1855, new_n1856,
    new_n1857, new_n1858, new_n1859, new_n1860, new_n1861, new_n1862,
    new_n1863, new_n1864, new_n1865, new_n1866, new_n1867, new_n1868,
    new_n1869, new_n1870, new_n1871, new_n1872, new_n1873, new_n1874,
    new_n1875, new_n1876, new_n1877, new_n1878, new_n1879, new_n1880,
    new_n1881, new_n1882, new_n1883, new_n1884, new_n1885, new_n1886,
    new_n1887, new_n1888, new_n1889, new_n1890, new_n1891, new_n1892,
    new_n1893, new_n1894, new_n1895, new_n1896, new_n1897, new_n1898,
    new_n1899, new_n1900, new_n1901, new_n1902, new_n1903, new_n1904,
    new_n1905, new_n1906, new_n1907, new_n1908, new_n1909, new_n1910,
    new_n1911, new_n1912, new_n1913, new_n1914, new_n1915, new_n1916,
    new_n1917, new_n1918, new_n1919, new_n1920, new_n1921, new_n1922,
    new_n1923, new_n1924, new_n1925, new_n1926, new_n1927, new_n1928,
    new_n1929, new_n1930, new_n1931, new_n1932, new_n1933, new_n1934,
    new_n1935, new_n1936, new_n1937, new_n1938, new_n1939, new_n1940,
    new_n1941, new_n1942, new_n1943, new_n1944, new_n1945, new_n1946,
    new_n1947, new_n1948, new_n1949, new_n1950, new_n1951, new_n1952,
    new_n1953, new_n1954, new_n1955, new_n1956, new_n1957, new_n1958,
    new_n1959, new_n1960, new_n1961, new_n1962, new_n1963, new_n1964,
    new_n1965, new_n1966, new_n1967, new_n1968, new_n1969, new_n1970,
    new_n1971, new_n1972, new_n1973, new_n1974, new_n1975, new_n1976,
    new_n1977, new_n1978, new_n1979, new_n1980, new_n1981, new_n1982,
    new_n1983, new_n1984, new_n1985, new_n1986, new_n1987, new_n1988,
    new_n1989, new_n1990, new_n1991, new_n1992, new_n1993, new_n1994,
    new_n1995, new_n1996, new_n1997, new_n1998, new_n1999, new_n2000,
    new_n2001, new_n2002, new_n2003, new_n2004, new_n2005, new_n2006,
    new_n2007, new_n2008, new_n2009, new_n2010, new_n2011, new_n2012,
    new_n2013, new_n2014, new_n2015, new_n2016, new_n2017, new_n2018,
    new_n2019, new_n2020, new_n2021, new_n2022, new_n2023, new_n2024,
    new_n2025, new_n2026, new_n2027, new_n2028, new_n2029, new_n2030,
    new_n2031, new_n2032, new_n2033, new_n2034, new_n2035, new_n2036,
    new_n2037, new_n2038, new_n2039, new_n2040, new_n2041, new_n2042,
    new_n2043, new_n2044, new_n2045, new_n2046, new_n2047, new_n2048,
    new_n2049, new_n2050, new_n2051, new_n2052, new_n2053, new_n2054,
    new_n2055, new_n2056, new_n2057, new_n2058, new_n2059, new_n2060,
    new_n2061, new_n2062, new_n2063, new_n2064, new_n2065, new_n2066,
    new_n2067, new_n2068, new_n2069, new_n2070, new_n2071, new_n2072,
    new_n2073, new_n2074, new_n2075, new_n2076, new_n2077, new_n2078,
    new_n2079, new_n2080, new_n2081, new_n2082, new_n2083, new_n2084,
    new_n2085, new_n2086, new_n2087, new_n2088, new_n2089, new_n2090,
    new_n2091, new_n2092, new_n2093, new_n2094, new_n2095, new_n2096,
    new_n2097, new_n2098, new_n2099, new_n2100, new_n2101, new_n2102,
    new_n2103, new_n2104, new_n2105, new_n2106, new_n2107, new_n2108,
    new_n2109, new_n2110, new_n2111, new_n2112, new_n2113, new_n2114,
    new_n2115, new_n2116, new_n2117, new_n2118, new_n2119, new_n2120,
    new_n2121, new_n2122, new_n2123, new_n2124, new_n2125, new_n2126,
    new_n2127, new_n2128, new_n2129, new_n2130, new_n2131, new_n2132,
    new_n2133, new_n2134, new_n2135, new_n2136, new_n2137, new_n2138,
    new_n2139, new_n2140, new_n2141, new_n2142, new_n2143, new_n2144,
    new_n2145, new_n2146, new_n2147, new_n2148, new_n2149, new_n2150,
    new_n2151, new_n2152, new_n2153, new_n2154, new_n2155, new_n2156,
    new_n2157, new_n2158, new_n2159, new_n2160, new_n2161, new_n2162,
    new_n2163, new_n2164, new_n2165, new_n2166, new_n2167, new_n2168,
    new_n2169, new_n2170, new_n2171, new_n2172, new_n2173, new_n2174,
    new_n2175, new_n2176, new_n2177, new_n2178, new_n2179, new_n2180,
    new_n2181, new_n2182, new_n2183, new_n2184, new_n2185, new_n2186,
    new_n2187, new_n2188, new_n2189, new_n2190, new_n2191, new_n2192,
    new_n2193, new_n2194, new_n2195, new_n2196, new_n2197, new_n2198,
    new_n2199, new_n2200, new_n2201, new_n2202, new_n2203, new_n2204,
    new_n2205, new_n2206, new_n2207, new_n2208, new_n2209, new_n2210,
    new_n2211, new_n2212, new_n2213, new_n2214, new_n2215, new_n2216,
    new_n2217, new_n2218, new_n2219, new_n2220, new_n2221, new_n2222,
    new_n2223, new_n2224, new_n2225, new_n2226, new_n2227, new_n2228,
    new_n2229, new_n2230, new_n2231, new_n2232, new_n2233, new_n2234,
    new_n2235, new_n2236, new_n2237, new_n2238, new_n2239, new_n2240,
    new_n2241, new_n2242, new_n2243, new_n2244, new_n2245, new_n2246,
    new_n2247, new_n2248, new_n2249, new_n2250, new_n2251, new_n2252,
    new_n2253, new_n2254, new_n2255, new_n2256, new_n2257, new_n2258,
    new_n2259, new_n2260, new_n2261, new_n2262, new_n2263, new_n2264,
    new_n2265, new_n2266, new_n2267, new_n2268, new_n2269, new_n2270,
    new_n2271, new_n2272, new_n2273, new_n2274, new_n2275, new_n2276,
    new_n2277, new_n2278, new_n2279, new_n2280, new_n2281, new_n2282,
    new_n2283, new_n2284, new_n2285, new_n2286, new_n2287, new_n2288,
    new_n2289, new_n2290, new_n2291, new_n2292, new_n2293, new_n2294,
    new_n2295, new_n2296, new_n2297, new_n2298, new_n2299, new_n2300,
    new_n2301, new_n2302, new_n2303, new_n2304, new_n2305, new_n2306,
    new_n2307, new_n2308, new_n2309, new_n2310, new_n2311, new_n2312,
    new_n2313, new_n2314, new_n2315, new_n2316, new_n2317, new_n2318,
    new_n2319, new_n2320, new_n2321, new_n2322, new_n2323, new_n2324,
    new_n2325, new_n2326, new_n2327, new_n2328, new_n2329, new_n2330,
    new_n2331, new_n2332, new_n2333, new_n2334, new_n2335, new_n2336,
    new_n2337, new_n2338, new_n2339, new_n2340, new_n2341, new_n2342,
    new_n2343, new_n2344, new_n2345, new_n2346, new_n2347, new_n2348,
    new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2362, new_n2363, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513, new_n2514, new_n2515, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2551, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577, new_n2578, new_n2579, new_n2580, new_n2581, new_n2582,
    new_n2583, new_n2584, new_n2585, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726,
    new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732,
    new_n2733, new_n2734, new_n2735, new_n2736, new_n2737, new_n2738,
    new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802, new_n2803, new_n2804,
    new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870,
    new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2879, new_n2880, new_n2881, new_n2882,
    new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902, new_n2903, new_n2904, new_n2905, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912,
    new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918,
    new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924,
    new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930,
    new_n2931, new_n2932, new_n2933, new_n2934, new_n2935, new_n2936,
    new_n2937, new_n2938, new_n2939, new_n2940, new_n2941, new_n2942,
    new_n2943, new_n2944, new_n2945, new_n2946, new_n2947, new_n2948,
    new_n2949, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954,
    new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2960,
    new_n2961, new_n2962, new_n2963, new_n2964, new_n2965, new_n2966,
    new_n2967, new_n2968, new_n2969, new_n2970, new_n2971, new_n2972,
    new_n2973, new_n2974, new_n2975, new_n2976, new_n2977, new_n2978,
    new_n2979, new_n2980, new_n2981, new_n2982, new_n2983, new_n2984,
    new_n2985, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990,
    new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996,
    new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3002,
    new_n3003, new_n3004, new_n3005, new_n3006, new_n3007, new_n3008,
    new_n3009, new_n3010, new_n3011, new_n3012, new_n3013, new_n3014,
    new_n3015, new_n3016, new_n3017, new_n3018, new_n3019, new_n3020,
    new_n3021, new_n3022, new_n3023, new_n3024, new_n3025, new_n3026,
    new_n3027, new_n3028, new_n3029, new_n3030, new_n3031, new_n3032,
    new_n3033, new_n3034, new_n3035, new_n3036, new_n3037, new_n3038,
    new_n3039, new_n3040, new_n3041, new_n3042, new_n3043, new_n3044,
    new_n3045, new_n3046, new_n3047, new_n3048, new_n3049, new_n3050,
    new_n3051, new_n3052, new_n3053, new_n3054, new_n3055, new_n3056,
    new_n3057, new_n3058, new_n3059, new_n3060, new_n3061, new_n3062,
    new_n3063, new_n3064, new_n3065, new_n3066, new_n3067, new_n3068,
    new_n3069, new_n3070, new_n3071, new_n3072, new_n3073, new_n3074,
    new_n3075, new_n3076, new_n3077, new_n3078, new_n3079, new_n3080,
    new_n3081, new_n3082, new_n3083, new_n3084, new_n3085, new_n3086,
    new_n3087, new_n3088, new_n3089, new_n3090, new_n3091, new_n3092,
    new_n3093, new_n3094, new_n3095, new_n3096, new_n3097, new_n3098,
    new_n3099, new_n3100, new_n3101, new_n3102, new_n3103, new_n3104,
    new_n3105, new_n3106, new_n3107, new_n3108, new_n3109, new_n3110,
    new_n3111, new_n3112, new_n3113, new_n3114, new_n3115, new_n3116,
    new_n3117, new_n3118, new_n3119, new_n3120, new_n3121, new_n3122,
    new_n3123, new_n3124, new_n3125, new_n3126, new_n3127, new_n3128,
    new_n3129, new_n3130, new_n3131, new_n3132, new_n3133, new_n3134,
    new_n3135, new_n3136, new_n3137, new_n3138, new_n3139, new_n3140,
    new_n3141, new_n3142, new_n3143, new_n3144, new_n3145, new_n3146,
    new_n3147, new_n3148, new_n3149, new_n3150, new_n3151, new_n3152,
    new_n3153, new_n3154, new_n3155, new_n3156, new_n3157, new_n3158,
    new_n3159, new_n3160, new_n3161, new_n3162, new_n3163, new_n3164,
    new_n3165, new_n3166, new_n3167, new_n3168, new_n3169, new_n3170,
    new_n3171, new_n3172, new_n3173, new_n3174, new_n3175, new_n3176,
    new_n3177, new_n3178, new_n3179, new_n3180, new_n3181, new_n3182,
    new_n3183, new_n3184, new_n3185, new_n3186, new_n3187, new_n3188,
    new_n3189, new_n3190, new_n3191, new_n3192, new_n3193, new_n3194,
    new_n3195, new_n3196, new_n3197, new_n3198, new_n3199, new_n3200,
    new_n3201, new_n3202, new_n3203, new_n3204, new_n3205, new_n3206,
    new_n3207, new_n3208, new_n3209, new_n3210, new_n3211, new_n3212,
    new_n3213, new_n3214, new_n3215, new_n3216, new_n3217, new_n3218,
    new_n3219, new_n3220, new_n3221, new_n3222, new_n3223, new_n3224,
    new_n3225, new_n3226, new_n3227, new_n3228, new_n3229, new_n3230,
    new_n3231, new_n3232, new_n3233, new_n3234, new_n3235, new_n3236,
    new_n3237, new_n3238, new_n3239, new_n3240, new_n3241, new_n3242,
    new_n3243, new_n3244, new_n3245, new_n3246, new_n3247, new_n3248,
    new_n3249, new_n3250, new_n3251, new_n3252, new_n3253, new_n3254,
    new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260,
    new_n3261, new_n3262, new_n3263, new_n3264, new_n3265, new_n3266,
    new_n3267, new_n3268, new_n3269, new_n3270, new_n3271, new_n3272,
    new_n3273, new_n3274, new_n3275, new_n3276, new_n3277, new_n3278,
    new_n3279, new_n3280, new_n3281, new_n3282, new_n3283, new_n3284,
    new_n3285, new_n3286, new_n3287, new_n3288, new_n3289, new_n3290,
    new_n3291, new_n3292, new_n3293, new_n3294, new_n3295, new_n3296,
    new_n3297, new_n3298, new_n3299, new_n3300, new_n3301, new_n3302,
    new_n3303, new_n3304, new_n3305, new_n3306, new_n3307, new_n3308,
    new_n3309, new_n3310, new_n3311, new_n3312, new_n3313, new_n3314,
    new_n3315, new_n3316, new_n3317, new_n3318, new_n3319, new_n3320,
    new_n3321, new_n3322, new_n3323, new_n3324, new_n3325, new_n3326,
    new_n3327, new_n3328, new_n3329, new_n3330, new_n3331, new_n3332,
    new_n3333, new_n3334, new_n3335, new_n3336, new_n3337, new_n3338,
    new_n3339, new_n3340, new_n3341, new_n3342, new_n3343, new_n3344,
    new_n3345, new_n3346, new_n3347, new_n3348, new_n3349, new_n3350,
    new_n3351, new_n3352, new_n3353, new_n3354, new_n3355, new_n3356,
    new_n3357, new_n3358, new_n3359, new_n3360, new_n3361, new_n3362,
    new_n3363, new_n3364, new_n3365, new_n3366, new_n3367, new_n3368,
    new_n3369, new_n3370, new_n3371, new_n3372, new_n3373, new_n3374,
    new_n3375, new_n3376, new_n3377, new_n3378, new_n3379, new_n3380,
    new_n3381, new_n3382, new_n3383, new_n3384, new_n3385, new_n3386,
    new_n3387, new_n3388, new_n3389, new_n3390, new_n3391, new_n3392,
    new_n3393, new_n3394, new_n3395, new_n3396, new_n3397, new_n3398,
    new_n3399, new_n3400, new_n3401, new_n3402, new_n3403, new_n3404,
    new_n3405, new_n3406, new_n3407, new_n3408, new_n3409, new_n3410,
    new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416,
    new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425, new_n3426, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458,
    new_n3459, new_n3460, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502, new_n3503, new_n3504, new_n3505, new_n3506,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561, new_n3562, new_n3563, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616, new_n3617, new_n3618, new_n3619, new_n3620,
    new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626,
    new_n3627, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649, new_n3650,
    new_n3651, new_n3652, new_n3653, new_n3654, new_n3655, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3724, new_n3725, new_n3726, new_n3727, new_n3728,
    new_n3729, new_n3730, new_n3731, new_n3732, new_n3733, new_n3734,
    new_n3735, new_n3736, new_n3737, new_n3738, new_n3739, new_n3740,
    new_n3741, new_n3742, new_n3743, new_n3744, new_n3745, new_n3746,
    new_n3747, new_n3748, new_n3749, new_n3750, new_n3751, new_n3752,
    new_n3753, new_n3754, new_n3755, new_n3756, new_n3757, new_n3758,
    new_n3759, new_n3760, new_n3761, new_n3762, new_n3763, new_n3764,
    new_n3765, new_n3766, new_n3767, new_n3768, new_n3769, new_n3770,
    new_n3771, new_n3772, new_n3773, new_n3774, new_n3775, new_n3776,
    new_n3777, new_n3778, new_n3779, new_n3780, new_n3781, new_n3782,
    new_n3783, new_n3784, new_n3785, new_n3786, new_n3787, new_n3788,
    new_n3789, new_n3790, new_n3791, new_n3792, new_n3793, new_n3794,
    new_n3795, new_n3796, new_n3797, new_n3798, new_n3799, new_n3800,
    new_n3801, new_n3802, new_n3803, new_n3804, new_n3805, new_n3806,
    new_n3807, new_n3808, new_n3809, new_n3810, new_n3811, new_n3812,
    new_n3813, new_n3814, new_n3815, new_n3816, new_n3817, new_n3818,
    new_n3819, new_n3820, new_n3821, new_n3822, new_n3823, new_n3824,
    new_n3825, new_n3826, new_n3827, new_n3828, new_n3829, new_n3830,
    new_n3831, new_n3832, new_n3833, new_n3834, new_n3835, new_n3836,
    new_n3837, new_n3838, new_n3839, new_n3840, new_n3841, new_n3842,
    new_n3843, new_n3844, new_n3845, new_n3846, new_n3847, new_n3848,
    new_n3849, new_n3850, new_n3851, new_n3852, new_n3853, new_n3854,
    new_n3855, new_n3856, new_n3857, new_n3858, new_n3859, new_n3860,
    new_n3861, new_n3862, new_n3863, new_n3864, new_n3865, new_n3866,
    new_n3867, new_n3868, new_n3869, new_n3870, new_n3871, new_n3872,
    new_n3873, new_n3874, new_n3875, new_n3876, new_n3877, new_n3878,
    new_n3879, new_n3880, new_n3881, new_n3882, new_n3883, new_n3884,
    new_n3885, new_n3886, new_n3887, new_n3888, new_n3889, new_n3890,
    new_n3891, new_n3892, new_n3893, new_n3894, new_n3895, new_n3896,
    new_n3897, new_n3898, new_n3899, new_n3900, new_n3901, new_n3902,
    new_n3903, new_n3904, new_n3905, new_n3906, new_n3907, new_n3908,
    new_n3909, new_n3910, new_n3911, new_n3912, new_n3913, new_n3914,
    new_n3915, new_n3916, new_n3917, new_n3918, new_n3919, new_n3920,
    new_n3921, new_n3922, new_n3923, new_n3924, new_n3925, new_n3926,
    new_n3927, new_n3928, new_n3929, new_n3930, new_n3931, new_n3932,
    new_n3933, new_n3934, new_n3935, new_n3936, new_n3937, new_n3938,
    new_n3939, new_n3940, new_n3941, new_n3942, new_n3943, new_n3944,
    new_n3945, new_n3946, new_n3947, new_n3948, new_n3949, new_n3950,
    new_n3951, new_n3952, new_n3953, new_n3954, new_n3955, new_n3956,
    new_n3957, new_n3958, new_n3959, new_n3960, new_n3961, new_n3962,
    new_n3963, new_n3964, new_n3965, new_n3966, new_n3967, new_n3968,
    new_n3969, new_n3970, new_n3971, new_n3972, new_n3973, new_n3974,
    new_n3975, new_n3976, new_n3977, new_n3978, new_n3979, new_n3980,
    new_n3981, new_n3982, new_n3983, new_n3984, new_n3985, new_n3986,
    new_n3987, new_n3988, new_n3989, new_n3990, new_n3991, new_n3992,
    new_n3993, new_n3994, new_n3995, new_n3996, new_n3997, new_n3998,
    new_n3999, new_n4000, new_n4001, new_n4002, new_n4003, new_n4004,
    new_n4005, new_n4006, new_n4007, new_n4008, new_n4009, new_n4010,
    new_n4011, new_n4012, new_n4013, new_n4014, new_n4015, new_n4016,
    new_n4017, new_n4018, new_n4019, new_n4020, new_n4021, new_n4022,
    new_n4023, new_n4024, new_n4025, new_n4026, new_n4027, new_n4028,
    new_n4029, new_n4030, new_n4031, new_n4032, new_n4033, new_n4034,
    new_n4035, new_n4036, new_n4037, new_n4038, new_n4039, new_n4040,
    new_n4041, new_n4042, new_n4043, new_n4044, new_n4045, new_n4046,
    new_n4047, new_n4048, new_n4049, new_n4050, new_n4051, new_n4052,
    new_n4053, new_n4054, new_n4055, new_n4056, new_n4057, new_n4058,
    new_n4059, new_n4060, new_n4061, new_n4062, new_n4063, new_n4064,
    new_n4065, new_n4066, new_n4067, new_n4068, new_n4069, new_n4070,
    new_n4071, new_n4072, new_n4073, new_n4074, new_n4075, new_n4076,
    new_n4077, new_n4078, new_n4079, new_n4080, new_n4081, new_n4082,
    new_n4083, new_n4084, new_n4085, new_n4086, new_n4087, new_n4088,
    new_n4089, new_n4090, new_n4091, new_n4092, new_n4093, new_n4094,
    new_n4095, new_n4096, new_n4097, new_n4098, new_n4099, new_n4100,
    new_n4101, new_n4102, new_n4103, new_n4104, new_n4105, new_n4106,
    new_n4107, new_n4108, new_n4109, new_n4110, new_n4111, new_n4112,
    new_n4113, new_n4114, new_n4115, new_n4116, new_n4117, new_n4118,
    new_n4119, new_n4120, new_n4121, new_n4122, new_n4123, new_n4124,
    new_n4125, new_n4126, new_n4127, new_n4128, new_n4129, new_n4130,
    new_n4131, new_n4132, new_n4133, new_n4134, new_n4135, new_n4136,
    new_n4137, new_n4138, new_n4139, new_n4140, new_n4141, new_n4142,
    new_n4143, new_n4144, new_n4145, new_n4146, new_n4147, new_n4148,
    new_n4149, new_n4150, new_n4151, new_n4152, new_n4153, new_n4154,
    new_n4155, new_n4156, new_n4157, new_n4158, new_n4159, new_n4160,
    new_n4161, new_n4162, new_n4163, new_n4164, new_n4165, new_n4166,
    new_n4167, new_n4168, new_n4169, new_n4170, new_n4171, new_n4172,
    new_n4173, new_n4174, new_n4175, new_n4176, new_n4177, new_n4178,
    new_n4179, new_n4180, new_n4181, new_n4182, new_n4183, new_n4184,
    new_n4185, new_n4186, new_n4187, new_n4188, new_n4189, new_n4190,
    new_n4191, new_n4192, new_n4193, new_n4194, new_n4195, new_n4196,
    new_n4197, new_n4198, new_n4199, new_n4200, new_n4201, new_n4202,
    new_n4203, new_n4204, new_n4205, new_n4206, new_n4207, new_n4208,
    new_n4209, new_n4210, new_n4211, new_n4212, new_n4213, new_n4214,
    new_n4215, new_n4216, new_n4217, new_n4218, new_n4219, new_n4220,
    new_n4221, new_n4222, new_n4223, new_n4224, new_n4225, new_n4226,
    new_n4227, new_n4228, new_n4229, new_n4230, new_n4231, new_n4232,
    new_n4233, new_n4234, new_n4235, new_n4236, new_n4237, new_n4238,
    new_n4239, new_n4240, new_n4241, new_n4242, new_n4243, new_n4244,
    new_n4245, new_n4246, new_n4247, new_n4248, new_n4249, new_n4250,
    new_n4251, new_n4252, new_n4253, new_n4254, new_n4255, new_n4256,
    new_n4257, new_n4258, new_n4259, new_n4260, new_n4261, new_n4262,
    new_n4263, new_n4264, new_n4265, new_n4266, new_n4267, new_n4268,
    new_n4269, new_n4270, new_n4271, new_n4272, new_n4273, new_n4274,
    new_n4275, new_n4276, new_n4277, new_n4278, new_n4279, new_n4280,
    new_n4281, new_n4282, new_n4283, new_n4284, new_n4285, new_n4286,
    new_n4287, new_n4288, new_n4289, new_n4290, new_n4291, new_n4292,
    new_n4293, new_n4294, new_n4295, new_n4296, new_n4297, new_n4298,
    new_n4299, new_n4300, new_n4301, new_n4302, new_n4303, new_n4304,
    new_n4305, new_n4306, new_n4307, new_n4308, new_n4309, new_n4310,
    new_n4311, new_n4312, new_n4313, new_n4314, new_n4315, new_n4316,
    new_n4317, new_n4318, new_n4319, new_n4320, new_n4321, new_n4322,
    new_n4323, new_n4324, new_n4325, new_n4326, new_n4327, new_n4328,
    new_n4329, new_n4330, new_n4331, new_n4332, new_n4333, new_n4334,
    new_n4335, new_n4336, new_n4337, new_n4338, new_n4339, new_n4340,
    new_n4341, new_n4342, new_n4343, new_n4344, new_n4345, new_n4346,
    new_n4347, new_n4348, new_n4349, new_n4350, new_n4351, new_n4352,
    new_n4353, new_n4354, new_n4355, new_n4356, new_n4357, new_n4358,
    new_n4359, new_n4360, new_n4361, new_n4362, new_n4363, new_n4364,
    new_n4365, new_n4366, new_n4367, new_n4368, new_n4369, new_n4370,
    new_n4371, new_n4372, new_n4373, new_n4374, new_n4375, new_n4376,
    new_n4377, new_n4378, new_n4379, new_n4380, new_n4381, new_n4382,
    new_n4383, new_n4384, new_n4385, new_n4386, new_n4387, new_n4388,
    new_n4389, new_n4390, new_n4391, new_n4392, new_n4393, new_n4394,
    new_n4395, new_n4396, new_n4397, new_n4398, new_n4399, new_n4400,
    new_n4401, new_n4402, new_n4403, new_n4404, new_n4405, new_n4406,
    new_n4407, new_n4408, new_n4409, new_n4410, new_n4411, new_n4412,
    new_n4413, new_n4414, new_n4415, new_n4416, new_n4417, new_n4418,
    new_n4419, new_n4420, new_n4421, new_n4422, new_n4423, new_n4424,
    new_n4425, new_n4426, new_n4427, new_n4428, new_n4429, new_n4430,
    new_n4431, new_n4432, new_n4433, new_n4434, new_n4435, new_n4436,
    new_n4437, new_n4438, new_n4439, new_n4440, new_n4441, new_n4442,
    new_n4443, new_n4444, new_n4445, new_n4446, new_n4447, new_n4448,
    new_n4449, new_n4450, new_n4451, new_n4452, new_n4453, new_n4454,
    new_n4455, new_n4456, new_n4457, new_n4458, new_n4459, new_n4460,
    new_n4461, new_n4462, new_n4463, new_n4464, new_n4465, new_n4466,
    new_n4467, new_n4468, new_n4469, new_n4470, new_n4471, new_n4472,
    new_n4473, new_n4474, new_n4475, new_n4476, new_n4477, new_n4478,
    new_n4479, new_n4480, new_n4481, new_n4482, new_n4483, new_n4484,
    new_n4485, new_n4486, new_n4487, new_n4488, new_n4489, new_n4490,
    new_n4491, new_n4492, new_n4493, new_n4494, new_n4495, new_n4496,
    new_n4497, new_n4498, new_n4499, new_n4500, new_n4501, new_n4502,
    new_n4503, new_n4504, new_n4505, new_n4506, new_n4507, new_n4508,
    new_n4509, new_n4510, new_n4511, new_n4512, new_n4513, new_n4514,
    new_n4515, new_n4516, new_n4517, new_n4518, new_n4519, new_n4520,
    new_n4521, new_n4522, new_n4523, new_n4524, new_n4525, new_n4526,
    new_n4527, new_n4528, new_n4529, new_n4530, new_n4531, new_n4532,
    new_n4533, new_n4534, new_n4535, new_n4536, new_n4537, new_n4538,
    new_n4539, new_n4540, new_n4541, new_n4542, new_n4543, new_n4544,
    new_n4545, new_n4546, new_n4547, new_n4548, new_n4549, new_n4550,
    new_n4551, new_n4552, new_n4553, new_n4554, new_n4555, new_n4556,
    new_n4557, new_n4558, new_n4559, new_n4560, new_n4561, new_n4562,
    new_n4563, new_n4564, new_n4565, new_n4566, new_n4567, new_n4568,
    new_n4569, new_n4570, new_n4571, new_n4572, new_n4573, new_n4574,
    new_n4575, new_n4576, new_n4577, new_n4578, new_n4579, new_n4580,
    new_n4581, new_n4582, new_n4583, new_n4584, new_n4585, new_n4586,
    new_n4587, new_n4588, new_n4589, new_n4590, new_n4591, new_n4592,
    new_n4593, new_n4594, new_n4595, new_n4596, new_n4597, new_n4598,
    new_n4599, new_n4600, new_n4601, new_n4602, new_n4603, new_n4604,
    new_n4605, new_n4606, new_n4607, new_n4608, new_n4609, new_n4610,
    new_n4611, new_n4612, new_n4613, new_n4614, new_n4615, new_n4616,
    new_n4617, new_n4618, new_n4619, new_n4620, new_n4621, new_n4622,
    new_n4623, new_n4624, new_n4625, new_n4626, new_n4627, new_n4628,
    new_n4629, new_n4630, new_n4631, new_n4632, new_n4633, new_n4634,
    new_n4635, new_n4636, new_n4637, new_n4638, new_n4639, new_n4640,
    new_n4641, new_n4642, new_n4643, new_n4644, new_n4645, new_n4646,
    new_n4647, new_n4648, new_n4649, new_n4650, new_n4651, new_n4652,
    new_n4653, new_n4654, new_n4655, new_n4656, new_n4657, new_n4658,
    new_n4659, new_n4660, new_n4661, new_n4662, new_n4663, new_n4664,
    new_n4665, new_n4666, new_n4667, new_n4668, new_n4669, new_n4670,
    new_n4671, new_n4672, new_n4673, new_n4674, new_n4675, new_n4676,
    new_n4677, new_n4678, new_n4679, new_n4680, new_n4681, new_n4682,
    new_n4683, new_n4684, new_n4685, new_n4686, new_n4687, new_n4688,
    new_n4689, new_n4690, new_n4691, new_n4692, new_n4693, new_n4694,
    new_n4695, new_n4696, new_n4697, new_n4698, new_n4699, new_n4700,
    new_n4701, new_n4702, new_n4703, new_n4704, new_n4705, new_n4706,
    new_n4707, new_n4708, new_n4709, new_n4710, new_n4711, new_n4712,
    new_n4713, new_n4714, new_n4715, new_n4716, new_n4717, new_n4718,
    new_n4719, new_n4720, new_n4721, new_n4722, new_n4723, new_n4724,
    new_n4725, new_n4726, new_n4727, new_n4728, new_n4729, new_n4730,
    new_n4731, new_n4732, new_n4733, new_n4734, new_n4735, new_n4736,
    new_n4737, new_n4738, new_n4739, new_n4740, new_n4741, new_n4742,
    new_n4743, new_n4744, new_n4745, new_n4746, new_n4747, new_n4748,
    new_n4749, new_n4750, new_n4751, new_n4752, new_n4753, new_n4754,
    new_n4755, new_n4756, new_n4757, new_n4758, new_n4759, new_n4760,
    new_n4761, new_n4762, new_n4763, new_n4764, new_n4765, new_n4766,
    new_n4767, new_n4768, new_n4769, new_n4770, new_n4771, new_n4772,
    new_n4773, new_n4774, new_n4775, new_n4776, new_n4777, new_n4778,
    new_n4779, new_n4780, new_n4781, new_n4782, new_n4783, new_n4784,
    new_n4785, new_n4786, new_n4787, new_n4788, new_n4789, new_n4790,
    new_n4791, new_n4792, new_n4793, new_n4794, new_n4795, new_n4796,
    new_n4797, new_n4798, new_n4799, new_n4800, new_n4801, new_n4802,
    new_n4803, new_n4804, new_n4805, new_n4806, new_n4807, new_n4808,
    new_n4809, new_n4810, new_n4811, new_n4812, new_n4813, new_n4814,
    new_n4815, new_n4816, new_n4817, new_n4818, new_n4819, new_n4820,
    new_n4821, new_n4822, new_n4823, new_n4824, new_n4825, new_n4826,
    new_n4827, new_n4828, new_n4829, new_n4830, new_n4831, new_n4832,
    new_n4833, new_n4834, new_n4835, new_n4836, new_n4837, new_n4838,
    new_n4839, new_n4840, new_n4841, new_n4842, new_n4843, new_n4844,
    new_n4845, new_n4846, new_n4847, new_n4848, new_n4849, new_n4850,
    new_n4851, new_n4852, new_n4853, new_n4854, new_n4855, new_n4856,
    new_n4857, new_n4858, new_n4859, new_n4860, new_n4861, new_n4862,
    new_n4863, new_n4864, new_n4865, new_n4866, new_n4867, new_n4868,
    new_n4869, new_n4870, new_n4871, new_n4872, new_n4873, new_n4874,
    new_n4875, new_n4876, new_n4877, new_n4878, new_n4879, new_n4880,
    new_n4881, new_n4882, new_n4883, new_n4884, new_n4885, new_n4886,
    new_n4887, new_n4888, new_n4889, new_n4890, new_n4891, new_n4892,
    new_n4893, new_n4894, new_n4895, new_n4896, new_n4897, new_n4898,
    new_n4899, new_n4900, new_n4901, new_n4902, new_n4903, new_n4904,
    new_n4905, new_n4906, new_n4907, new_n4908, new_n4909, new_n4910,
    new_n4911, new_n4912, new_n4913, new_n4914, new_n4915, new_n4916,
    new_n4917, new_n4918, new_n4919, new_n4920, new_n4921, new_n4922,
    new_n4923, new_n4924, new_n4925, new_n4926, new_n4927, new_n4928,
    new_n4929, new_n4930, new_n4931, new_n4932, new_n4933, new_n4934,
    new_n4935, new_n4936, new_n4937, new_n4938, new_n4939, new_n4940,
    new_n4941, new_n4942, new_n4943, new_n4944, new_n4945, new_n4946,
    new_n4947, new_n4948, new_n4949, new_n4950, new_n4951, new_n4952,
    new_n4953, new_n4954, new_n4955, new_n4956, new_n4957, new_n4958,
    new_n4959, new_n4960, new_n4961, new_n4962, new_n4963, new_n4964,
    new_n4965, new_n4966, new_n4967, new_n4968, new_n4969, new_n4970,
    new_n4971, new_n4972, new_n4973, new_n4974, new_n4975, new_n4976,
    new_n4977, new_n4978, new_n4979, new_n4980, new_n4981, new_n4982,
    new_n4983, new_n4984, new_n4985, new_n4986, new_n4987, new_n4988,
    new_n4989, new_n4990, new_n4991, new_n4992, new_n4993, new_n4994,
    new_n4995, new_n4996, new_n4997, new_n4998, new_n4999, new_n5000,
    new_n5001, new_n5002, new_n5003, new_n5004, new_n5005, new_n5006,
    new_n5007, new_n5008, new_n5009, new_n5010, new_n5011, new_n5012,
    new_n5013, new_n5014, new_n5015, new_n5016, new_n5017, new_n5018,
    new_n5019, new_n5020, new_n5021, new_n5022, new_n5023, new_n5024,
    new_n5025, new_n5026, new_n5027, new_n5028, new_n5029, new_n5030,
    new_n5031, new_n5032, new_n5033, new_n5034, new_n5035, new_n5036,
    new_n5037, new_n5038, new_n5039, new_n5040, new_n5041, new_n5042,
    new_n5043, new_n5044, new_n5045, new_n5046, new_n5047, new_n5048,
    new_n5049, new_n5050, new_n5051, new_n5052, new_n5053, new_n5054,
    new_n5055, new_n5056, new_n5057, new_n5058, new_n5059, new_n5060,
    new_n5061, new_n5062, new_n5063, new_n5064, new_n5065, new_n5066,
    new_n5067, new_n5068, new_n5069, new_n5070, new_n5071, new_n5072,
    new_n5073, new_n5074, new_n5075, new_n5076, new_n5077, new_n5078,
    new_n5079, new_n5080, new_n5081, new_n5082, new_n5083, new_n5084,
    new_n5085, new_n5086, new_n5087, new_n5088, new_n5089, new_n5090,
    new_n5091, new_n5092, new_n5093, new_n5094, new_n5095, new_n5096,
    new_n5097, new_n5098, new_n5099, new_n5100, new_n5101, new_n5102,
    new_n5103, new_n5104, new_n5105, new_n5106, new_n5107, new_n5108,
    new_n5109, new_n5110, new_n5111, new_n5112, new_n5113, new_n5114,
    new_n5115, new_n5116, new_n5117, new_n5118, new_n5119, new_n5120,
    new_n5121, new_n5122, new_n5123, new_n5124, new_n5125, new_n5126,
    new_n5127, new_n5128, new_n5129, new_n5130, new_n5131, new_n5132,
    new_n5133, new_n5134, new_n5135, new_n5136, new_n5137, new_n5138,
    new_n5139, new_n5140, new_n5141, new_n5142, new_n5143, new_n5144,
    new_n5145, new_n5146, new_n5147, new_n5148, new_n5149, new_n5150,
    new_n5151, new_n5152, new_n5153, new_n5154, new_n5155, new_n5156,
    new_n5157, new_n5158, new_n5159, new_n5160, new_n5161, new_n5162,
    new_n5163, new_n5164, new_n5165, new_n5166, new_n5167, new_n5168,
    new_n5169, new_n5170, new_n5171, new_n5172, new_n5173, new_n5174,
    new_n5175, new_n5176, new_n5177, new_n5178, new_n5179, new_n5180,
    new_n5181, new_n5182, new_n5183, new_n5184, new_n5185, new_n5186,
    new_n5187, new_n5188, new_n5189, new_n5190, new_n5191, new_n5192,
    new_n5193, new_n5194, new_n5195, new_n5196, new_n5197, new_n5198,
    new_n5199, new_n5200, new_n5201, new_n5202, new_n5203, new_n5204,
    new_n5205, new_n5206, new_n5207, new_n5208, new_n5209, new_n5210,
    new_n5211, new_n5212, new_n5213, new_n5214, new_n5215, new_n5216,
    new_n5217, new_n5218, new_n5219, new_n5220, new_n5221, new_n5222,
    new_n5223, new_n5224, new_n5225, new_n5226, new_n5227, new_n5228,
    new_n5229, new_n5230, new_n5231, new_n5232, new_n5233, new_n5234,
    new_n5235, new_n5236, new_n5237, new_n5238, new_n5239, new_n5240,
    new_n5241, new_n5242, new_n5243, new_n5244, new_n5245, new_n5246,
    new_n5247, new_n5248, new_n5249, new_n5250, new_n5251, new_n5252,
    new_n5253, new_n5254, new_n5255, new_n5256, new_n5257, new_n5258,
    new_n5259, new_n5260, new_n5261, new_n5262, new_n5263, new_n5264,
    new_n5265, new_n5266, new_n5267, new_n5268, new_n5269, new_n5270,
    new_n5271, new_n5272, new_n5273, new_n5274, new_n5275, new_n5276,
    new_n5277, new_n5278, new_n5279, new_n5280, new_n5281, new_n5282,
    new_n5283, new_n5284, new_n5285, new_n5286, new_n5287, new_n5288,
    new_n5289, new_n5290, new_n5291, new_n5292, new_n5293, new_n5294,
    new_n5295, new_n5296, new_n5297, new_n5298, new_n5299, new_n5300,
    new_n5301, new_n5302, new_n5303, new_n5304, new_n5305, new_n5306,
    new_n5307, new_n5308, new_n5309, new_n5310, new_n5311, new_n5312,
    new_n5313, new_n5314, new_n5315, new_n5316, new_n5317, new_n5318,
    new_n5319, new_n5320, new_n5321, new_n5322, new_n5323, new_n5324,
    new_n5325, new_n5326, new_n5327, new_n5328, new_n5329, new_n5330,
    new_n5331, new_n5332, new_n5333, new_n5334, new_n5335, new_n5336,
    new_n5337, new_n5338, new_n5339, new_n5340, new_n5341, new_n5342,
    new_n5343, new_n5344, new_n5345, new_n5346, new_n5347, new_n5348,
    new_n5349, new_n5350, new_n5351, new_n5352, new_n5353, new_n5354,
    new_n5355, new_n5356, new_n5357, new_n5358, new_n5359, new_n5360,
    new_n5361, new_n5362, new_n5363, new_n5364, new_n5365, new_n5366,
    new_n5367, new_n5368, new_n5369, new_n5370, new_n5371, new_n5372,
    new_n5373, new_n5374, new_n5375, new_n5376, new_n5377, new_n5378,
    new_n5379, new_n5380, new_n5381, new_n5382, new_n5383, new_n5384,
    new_n5385, new_n5386, new_n5387, new_n5388, new_n5389, new_n5390,
    new_n5391, new_n5392, new_n5393, new_n5394, new_n5395, new_n5396,
    new_n5397, new_n5398, new_n5399, new_n5400, new_n5401, new_n5402,
    new_n5403, new_n5404, new_n5405, new_n5406, new_n5407, new_n5408,
    new_n5409, new_n5410, new_n5411, new_n5412, new_n5413, new_n5414,
    new_n5415, new_n5416, new_n5417, new_n5418, new_n5419, new_n5420,
    new_n5421, new_n5422, new_n5423, new_n5424, new_n5425, new_n5426,
    new_n5427, new_n5428, new_n5429, new_n5430, new_n5431, new_n5432,
    new_n5433, new_n5434, new_n5435, new_n5436, new_n5437, new_n5438,
    new_n5439, new_n5440, new_n5441, new_n5442, new_n5443, new_n5444,
    new_n5445, new_n5446, new_n5447, new_n5448, new_n5449, new_n5450,
    new_n5451, new_n5452, new_n5453, new_n5454, new_n5455, new_n5456,
    new_n5457, new_n5458, new_n5459, new_n5460, new_n5461, new_n5462,
    new_n5463, new_n5464, new_n5465, new_n5466, new_n5467, new_n5468,
    new_n5469, new_n5470, new_n5471, new_n5472, new_n5473, new_n5474,
    new_n5475, new_n5476, new_n5477, new_n5478, new_n5479, new_n5480,
    new_n5481, new_n5482, new_n5483, new_n5484, new_n5485, new_n5486,
    new_n5487, new_n5488, new_n5489, new_n5490, new_n5491, new_n5492,
    new_n5493, new_n5494, new_n5495, new_n5496, new_n5497, new_n5498,
    new_n5499, new_n5500, new_n5501, new_n5502, new_n5503, new_n5504,
    new_n5505, new_n5506, new_n5507, new_n5508, new_n5509, new_n5510,
    new_n5511, new_n5512, new_n5513, new_n5514, new_n5515, new_n5516,
    new_n5517, new_n5518, new_n5519, new_n5520, new_n5521, new_n5522,
    new_n5523, new_n5524, new_n5525, new_n5526, new_n5527, new_n5528,
    new_n5529, new_n5530, new_n5531, new_n5532, new_n5533, new_n5534,
    new_n5535, new_n5536, new_n5537, new_n5538, new_n5539, new_n5540,
    new_n5541, new_n5542, new_n5543, new_n5544, new_n5545, new_n5546,
    new_n5547, new_n5548, new_n5549, new_n5550, new_n5551, new_n5552,
    new_n5553, new_n5554, new_n5555, new_n5556, new_n5557, new_n5558,
    new_n5559, new_n5560, new_n5561, new_n5562, new_n5563, new_n5564,
    new_n5565, new_n5566, new_n5567, new_n5568, new_n5569, new_n5570,
    new_n5571, new_n5572, new_n5573, new_n5574, new_n5575, new_n5576,
    new_n5577, new_n5578, new_n5579, new_n5580, new_n5581, new_n5582,
    new_n5583, new_n5584, new_n5585, new_n5586, new_n5587, new_n5588,
    new_n5589, new_n5590, new_n5591, new_n5592, new_n5593, new_n5594,
    new_n5595, new_n5596, new_n5597, new_n5598, new_n5599, new_n5600,
    new_n5601, new_n5602, new_n5603, new_n5604, new_n5605, new_n5606,
    new_n5607, new_n5608, new_n5609, new_n5610, new_n5611, new_n5612,
    new_n5613, new_n5614, new_n5615, new_n5616, new_n5617, new_n5618,
    new_n5619, new_n5620, new_n5621, new_n5622, new_n5623, new_n5624,
    new_n5625, new_n5626, new_n5627, new_n5628, new_n5629, new_n5630,
    new_n5631, new_n5632, new_n5633, new_n5634, new_n5635, new_n5636,
    new_n5637, new_n5638, new_n5639, new_n5640, new_n5641, new_n5642,
    new_n5643, new_n5644, new_n5645, new_n5646, new_n5647, new_n5648,
    new_n5649, new_n5650, new_n5651, new_n5652, new_n5653, new_n5654,
    new_n5655, new_n5656, new_n5657, new_n5658, new_n5659, new_n5660,
    new_n5661, new_n5662, new_n5663, new_n5664, new_n5665, new_n5666,
    new_n5667, new_n5668, new_n5669, new_n5670, new_n5671, new_n5672,
    new_n5673, new_n5674, new_n5675, new_n5676, new_n5677, new_n5678,
    new_n5679, new_n5680, new_n5681, new_n5682, new_n5683, new_n5684,
    new_n5685, new_n5686, new_n5687, new_n5688, new_n5689, new_n5690,
    new_n5691, new_n5692, new_n5693, new_n5694, new_n5695, new_n5696,
    new_n5697, new_n5698, new_n5699, new_n5700, new_n5701, new_n5702,
    new_n5703, new_n5704, new_n5705, new_n5706, new_n5707, new_n5708,
    new_n5709, new_n5710, new_n5711, new_n5712, new_n5713, new_n5714,
    new_n5715, new_n5716, new_n5717, new_n5718, new_n5719, new_n5720,
    new_n5721, new_n5722, new_n5723, new_n5724, new_n5725, new_n5726,
    new_n5727, new_n5728, new_n5729, new_n5730, new_n5731, new_n5732,
    new_n5733, new_n5734, new_n5735, new_n5736, new_n5737, new_n5738,
    new_n5739, new_n5740, new_n5741, new_n5742, new_n5743, new_n5744,
    new_n5745, new_n5746, new_n5747, new_n5748, new_n5749, new_n5750,
    new_n5751, new_n5752, new_n5753, new_n5754, new_n5755, new_n5756,
    new_n5757, new_n5758, new_n5759, new_n5760, new_n5761, new_n5762,
    new_n5763, new_n5764, new_n5765, new_n5766, new_n5767, new_n5768,
    new_n5769, new_n5770, new_n5771, new_n5772, new_n5773, new_n5774,
    new_n5775, new_n5776, new_n5777, new_n5778, new_n5779, new_n5780,
    new_n5781, new_n5782, new_n5783, new_n5784, new_n5785, new_n5786,
    new_n5787, new_n5788, new_n5789, new_n5790, new_n5791, new_n5792,
    new_n5793, new_n5794, new_n5795, new_n5796, new_n5797, new_n5798,
    new_n5799, new_n5800, new_n5801, new_n5802, new_n5803, new_n5804,
    new_n5805, new_n5806, new_n5807, new_n5808, new_n5809, new_n5810,
    new_n5811, new_n5812, new_n5813, new_n5814, new_n5815, new_n5816,
    new_n5817, new_n5818, new_n5819, new_n5820, new_n5821, new_n5822,
    new_n5823, new_n5824, new_n5825, new_n5826, new_n5827, new_n5828,
    new_n5829, new_n5830, new_n5831, new_n5832, new_n5833, new_n5834,
    new_n5835, new_n5836, new_n5837, new_n5838, new_n5839, new_n5840,
    new_n5841, new_n5842, new_n5843, new_n5844, new_n5845, new_n5846,
    new_n5847, new_n5848, new_n5849, new_n5850, new_n5851, new_n5852,
    new_n5853, new_n5854, new_n5855, new_n5856, new_n5857, new_n5858,
    new_n5859, new_n5860, new_n5861, new_n5862, new_n5863, new_n5864,
    new_n5865, new_n5866, new_n5867, new_n5868, new_n5869, new_n5870,
    new_n5871, new_n5872, new_n5873, new_n5874, new_n5875, new_n5876,
    new_n5877, new_n5878, new_n5879, new_n5880, new_n5881, new_n5882,
    new_n5883, new_n5884, new_n5885, new_n5886, new_n5887, new_n5888,
    new_n5889, new_n5890, new_n5891, new_n5892, new_n5893, new_n5894,
    new_n5895, new_n5896, new_n5897, new_n5898, new_n5899, new_n5900,
    new_n5901, new_n5902, new_n5903, new_n5904, new_n5905, new_n5906,
    new_n5907, new_n5908, new_n5909, new_n5910, new_n5911, new_n5912,
    new_n5913, new_n5914, new_n5915, new_n5916, new_n5917, new_n5918,
    new_n5919, new_n5920, new_n5921, new_n5922, new_n5923, new_n5924,
    new_n5925, new_n5926, new_n5927, new_n5928, new_n5929, new_n5930,
    new_n5931, new_n5932, new_n5933, new_n5934, new_n5935, new_n5936,
    new_n5937, new_n5938, new_n5939, new_n5940, new_n5941, new_n5942,
    new_n5943, new_n5944, new_n5945, new_n5946, new_n5947, new_n5948,
    new_n5949, new_n5950, new_n5951, new_n5952, new_n5953, new_n5954,
    new_n5955, new_n5956, new_n5957, new_n5958, new_n5959, new_n5960,
    new_n5961, new_n5962, new_n5963, new_n5964, new_n5965, new_n5966,
    new_n5967, new_n5968, new_n5969, new_n5970, new_n5971, new_n5972,
    new_n5973, new_n5974, new_n5975, new_n5976, new_n5977, new_n5978,
    new_n5979, new_n5980, new_n5981, new_n5982, new_n5983, new_n5984,
    new_n5985, new_n5986, new_n5987, new_n5988, new_n5989, new_n5990,
    new_n5991, new_n5992, new_n5993, new_n5994, new_n5995, new_n5996,
    new_n5997, new_n5998, new_n5999, new_n6000, new_n6001, new_n6002,
    new_n6003, new_n6004, new_n6005, new_n6006, new_n6007, new_n6008,
    new_n6009, new_n6010, new_n6011, new_n6012, new_n6013, new_n6014,
    new_n6015, new_n6016, new_n6017, new_n6018, new_n6019, new_n6020,
    new_n6021, new_n6022, new_n6023, new_n6024, new_n6025, new_n6026,
    new_n6027, new_n6028, new_n6029, new_n6030, new_n6031, new_n6032,
    new_n6033, new_n6034, new_n6035, new_n6036, new_n6037, new_n6038,
    new_n6039, new_n6040, new_n6041, new_n6042, new_n6043, new_n6044,
    new_n6045, new_n6046, new_n6047, new_n6048, new_n6049, new_n6050,
    new_n6051, new_n6052, new_n6053, new_n6054, new_n6055, new_n6056,
    new_n6057, new_n6058, new_n6059, new_n6060, new_n6061, new_n6062,
    new_n6063, new_n6064, new_n6065, new_n6066, new_n6067, new_n6068,
    new_n6069, new_n6070, new_n6071, new_n6072, new_n6073, new_n6074,
    new_n6075, new_n6076, new_n6077, new_n6078, new_n6079, new_n6080,
    new_n6081, new_n6082, new_n6083, new_n6084, new_n6085, new_n6086,
    new_n6087, new_n6088, new_n6089, new_n6090, new_n6091, new_n6092,
    new_n6093, new_n6094, new_n6095, new_n6096, new_n6097, new_n6098,
    new_n6099, new_n6100, new_n6101, new_n6102, new_n6103, new_n6104,
    new_n6105, new_n6106, new_n6107, new_n6108, new_n6109, new_n6110,
    new_n6111, new_n6112, new_n6113, new_n6114, new_n6115, new_n6116,
    new_n6117, new_n6118, new_n6119, new_n6120, new_n6121, new_n6122,
    new_n6123, new_n6124, new_n6125, new_n6126, new_n6127, new_n6128,
    new_n6129, new_n6130, new_n6131, new_n6132, new_n6133, new_n6134,
    new_n6135, new_n6136, new_n6137, new_n6138, new_n6139, new_n6140,
    new_n6141, new_n6142, new_n6143, new_n6144, new_n6145, new_n6146,
    new_n6147, new_n6148, new_n6149, new_n6150, new_n6151, new_n6152,
    new_n6153, new_n6154, new_n6155, new_n6156, new_n6157, new_n6158,
    new_n6159, new_n6160, new_n6161, new_n6162, new_n6163, new_n6164,
    new_n6165, new_n6166, new_n6167, new_n6168, new_n6169, new_n6170,
    new_n6171, new_n6172, new_n6173, new_n6174, new_n6175, new_n6176,
    new_n6177, new_n6178, new_n6179, new_n6180, new_n6181, new_n6182,
    new_n6183, new_n6184, new_n6185, new_n6186, new_n6187, new_n6188,
    new_n6189, new_n6190, new_n6191, new_n6192, new_n6193, new_n6194,
    new_n6195, new_n6196, new_n6197, new_n6198, new_n6199, new_n6200,
    new_n6201, new_n6202, new_n6203, new_n6204, new_n6205, new_n6206,
    new_n6207, new_n6208, new_n6209, new_n6210, new_n6211, new_n6212,
    new_n6213, new_n6214, new_n6215, new_n6216, new_n6217, new_n6218,
    new_n6219, new_n6220, new_n6221, new_n6222, new_n6223, new_n6224,
    new_n6225, new_n6226, new_n6227, new_n6228, new_n6229, new_n6230,
    new_n6231, new_n6232, new_n6233, new_n6234, new_n6235, new_n6236,
    new_n6237, new_n6238, new_n6239, new_n6240, new_n6241, new_n6242,
    new_n6243, new_n6244, new_n6245, new_n6246, new_n6247, new_n6248,
    new_n6249, new_n6250, new_n6251, new_n6252, new_n6253, new_n6254,
    new_n6255, new_n6256, new_n6257, new_n6258, new_n6259, new_n6260,
    new_n6261, new_n6262, new_n6263, new_n6264, new_n6265, new_n6266,
    new_n6267, new_n6268, new_n6269, new_n6270, new_n6271, new_n6272,
    new_n6273, new_n6274, new_n6275, new_n6276, new_n6277, new_n6278,
    new_n6279, new_n6280, new_n6281, new_n6282, new_n6283, new_n6284,
    new_n6285, new_n6286, new_n6287, new_n6288, new_n6289, new_n6290,
    new_n6291, new_n6292, new_n6293, new_n6294, new_n6295, new_n6296,
    new_n6297, new_n6298, new_n6299, new_n6300, new_n6301, new_n6302,
    new_n6303, new_n6304, new_n6305, new_n6306, new_n6307, new_n6308,
    new_n6309, new_n6310, new_n6311, new_n6312, new_n6313, new_n6314,
    new_n6315, new_n6316, new_n6317, new_n6318, new_n6319, new_n6320,
    new_n6321, new_n6322, new_n6323, new_n6324, new_n6325, new_n6326,
    new_n6327, new_n6328, new_n6329, new_n6330, new_n6331, new_n6332,
    new_n6333, new_n6334, new_n6335, new_n6336, new_n6337, new_n6338,
    new_n6339, new_n6340, new_n6341, new_n6342, new_n6343, new_n6344,
    new_n6345, new_n6346, new_n6347, new_n6348, new_n6349, new_n6350,
    new_n6351, new_n6352, new_n6353, new_n6354, new_n6355, new_n6356,
    new_n6357, new_n6358, new_n6359, new_n6360, new_n6361, new_n6362,
    new_n6363, new_n6364, new_n6365, new_n6366, new_n6367, new_n6368,
    new_n6369, new_n6370, new_n6371, new_n6372, new_n6373, new_n6374,
    new_n6375, new_n6376, new_n6377, new_n6378, new_n6379, new_n6380,
    new_n6381, new_n6382, new_n6383, new_n6384, new_n6385, new_n6386,
    new_n6387, new_n6388, new_n6389, new_n6390, new_n6391, new_n6392,
    new_n6393, new_n6394, new_n6395, new_n6396, new_n6397, new_n6398,
    new_n6399, new_n6400, new_n6401, new_n6402, new_n6403, new_n6404,
    new_n6405, new_n6406, new_n6407, new_n6408, new_n6409, new_n6410,
    new_n6411, new_n6412, new_n6413, new_n6414, new_n6415, new_n6416,
    new_n6417, new_n6418, new_n6419, new_n6420, new_n6421, new_n6422,
    new_n6423, new_n6424, new_n6425, new_n6426, new_n6427, new_n6428,
    new_n6429, new_n6430, new_n6431, new_n6432, new_n6433, new_n6434,
    new_n6435, new_n6436, new_n6437, new_n6438, new_n6439, new_n6440,
    new_n6441, new_n6442, new_n6443, new_n6444, new_n6445, new_n6446,
    new_n6447, new_n6448, new_n6449, new_n6450, new_n6451, new_n6452,
    new_n6453, new_n6454, new_n6455, new_n6456, new_n6457, new_n6458,
    new_n6459, new_n6460, new_n6461, new_n6462, new_n6463, new_n6464,
    new_n6465, new_n6466, new_n6467, new_n6468, new_n6469, new_n6470,
    new_n6471, new_n6472, new_n6473, new_n6474, new_n6475, new_n6476,
    new_n6477, new_n6478, new_n6479, new_n6480, new_n6481, new_n6482,
    new_n6483, new_n6484, new_n6485, new_n6486, new_n6487, new_n6488,
    new_n6489, new_n6490, new_n6491, new_n6492, new_n6493, new_n6494,
    new_n6495, new_n6496, new_n6497, new_n6498, new_n6499, new_n6500,
    new_n6501, new_n6502, new_n6503, new_n6504, new_n6505, new_n6506,
    new_n6507, new_n6508, new_n6509, new_n6510, new_n6511, new_n6512,
    new_n6513, new_n6514, new_n6515, new_n6516, new_n6517, new_n6518,
    new_n6519, new_n6520, new_n6521, new_n6522, new_n6523, new_n6524,
    new_n6525, new_n6526, new_n6527, new_n6528, new_n6529, new_n6530,
    new_n6531, new_n6532, new_n6533, new_n6534, new_n6535, new_n6536,
    new_n6537, new_n6538, new_n6539, new_n6540, new_n6541, new_n6542,
    new_n6543, new_n6544, new_n6545, new_n6546, new_n6547, new_n6548,
    new_n6549, new_n6550, new_n6551, new_n6552, new_n6553, new_n6554,
    new_n6555, new_n6556, new_n6557, new_n6558, new_n6559, new_n6560,
    new_n6561, new_n6562, new_n6563, new_n6564, new_n6565, new_n6566,
    new_n6567, new_n6568, new_n6569, new_n6570, new_n6571, new_n6572,
    new_n6573, new_n6574, new_n6575, new_n6576, new_n6577, new_n6578,
    new_n6579, new_n6580, new_n6581, new_n6582, new_n6583, new_n6584,
    new_n6585, new_n6586, new_n6587, new_n6588, new_n6589, new_n6590,
    new_n6591, new_n6592, new_n6593, new_n6594, new_n6595, new_n6596,
    new_n6597, new_n6598, new_n6599, new_n6600, new_n6601, new_n6602,
    new_n6603, new_n6604, new_n6605, new_n6606, new_n6607, new_n6608,
    new_n6609, new_n6610, new_n6611, new_n6612, new_n6613, new_n6614,
    new_n6615, new_n6616, new_n6617, new_n6618, new_n6619, new_n6620,
    new_n6621, new_n6622, new_n6623, new_n6624, new_n6625, new_n6626,
    new_n6627, new_n6628, new_n6629, new_n6630, new_n6631, new_n6632,
    new_n6633, new_n6634, new_n6635, new_n6636, new_n6637, new_n6638,
    new_n6639, new_n6640, new_n6641, new_n6642, new_n6643, new_n6644,
    new_n6645, new_n6646, new_n6647, new_n6648, new_n6649, new_n6650,
    new_n6651, new_n6652, new_n6653, new_n6654, new_n6655, new_n6656,
    new_n6657, new_n6658, new_n6659, new_n6660, new_n6661, new_n6662,
    new_n6663, new_n6664, new_n6665, new_n6666, new_n6667, new_n6668,
    new_n6669, new_n6670, new_n6671, new_n6672, new_n6673, new_n6674,
    new_n6675, new_n6676, new_n6677, new_n6678, new_n6679, new_n6680,
    new_n6681, new_n6682, new_n6683, new_n6684, new_n6685, new_n6686,
    new_n6687, new_n6688, new_n6689, new_n6690, new_n6691, new_n6692,
    new_n6693, new_n6694, new_n6695, new_n6696, new_n6697, new_n6698,
    new_n6699, new_n6700, new_n6701, new_n6702, new_n6703, new_n6704,
    new_n6705, new_n6706, new_n6707, new_n6708, new_n6709, new_n6710,
    new_n6711, new_n6712, new_n6713, new_n6714, new_n6715, new_n6716,
    new_n6717, new_n6718, new_n6719, new_n6720, new_n6721, new_n6722,
    new_n6723, new_n6724, new_n6725, new_n6726, new_n6727, new_n6728,
    new_n6729, new_n6730, new_n6731, new_n6732, new_n6733, new_n6734,
    new_n6735, new_n6736, new_n6737, new_n6738, new_n6739, new_n6740,
    new_n6741, new_n6742, new_n6743, new_n6744, new_n6745, new_n6746,
    new_n6747, new_n6748, new_n6749, new_n6750, new_n6751, new_n6752,
    new_n6753, new_n6754, new_n6755, new_n6756, new_n6757, new_n6758,
    new_n6759, new_n6760, new_n6761, new_n6762, new_n6763, new_n6764,
    new_n6765, new_n6766, new_n6767, new_n6768, new_n6769, new_n6770,
    new_n6771, new_n6772, new_n6773, new_n6774, new_n6775, new_n6776,
    new_n6777, new_n6778, new_n6779, new_n6780, new_n6781, new_n6782,
    new_n6783, new_n6784, new_n6785, new_n6786, new_n6787, new_n6788,
    new_n6789, new_n6790, new_n6791, new_n6792, new_n6793, new_n6794,
    new_n6795, new_n6796, new_n6797, new_n6798, new_n6799, new_n6800,
    new_n6801, new_n6802, new_n6803, new_n6804, new_n6805, new_n6806,
    new_n6807, new_n6808, new_n6809, new_n6810, new_n6811, new_n6812,
    new_n6813, new_n6814, new_n6815, new_n6816, new_n6817, new_n6818,
    new_n6819, new_n6820, new_n6821, new_n6822, new_n6823, new_n6824,
    new_n6825, new_n6826, new_n6827, new_n6828, new_n6829, new_n6830,
    new_n6831, new_n6832, new_n6833, new_n6834, new_n6835, new_n6836,
    new_n6837, new_n6838, new_n6839, new_n6840, new_n6841, new_n6842,
    new_n6843, new_n6844, new_n6845, new_n6846, new_n6847, new_n6848,
    new_n6849, new_n6850, new_n6851, new_n6852, new_n6853, new_n6854,
    new_n6855, new_n6856, new_n6857, new_n6858, new_n6859, new_n6860,
    new_n6861, new_n6862, new_n6863, new_n6864, new_n6865, new_n6866,
    new_n6867, new_n6868, new_n6869, new_n6870, new_n6871, new_n6872,
    new_n6873, new_n6874, new_n6875, new_n6876, new_n6877, new_n6878,
    new_n6879, new_n6880, new_n6881, new_n6882, new_n6883, new_n6884,
    new_n6885, new_n6886, new_n6887, new_n6888, new_n6889, new_n6890,
    new_n6891, new_n6892, new_n6893, new_n6894, new_n6895, new_n6896,
    new_n6897, new_n6898, new_n6899, new_n6900, new_n6901, new_n6902,
    new_n6903, new_n6904, new_n6905, new_n6906, new_n6907, new_n6908,
    new_n6909, new_n6910, new_n6911, new_n6912, new_n6913, new_n6914,
    new_n6915, new_n6916, new_n6917, new_n6918, new_n6919, new_n6920,
    new_n6921, new_n6922, new_n6923, new_n6924, new_n6925, new_n6926,
    new_n6927, new_n6928, new_n6929, new_n6930, new_n6931, new_n6932,
    new_n6933, new_n6934, new_n6935, new_n6936, new_n6937, new_n6938,
    new_n6939, new_n6940, new_n6941, new_n6942, new_n6943, new_n6944,
    new_n6945, new_n6946, new_n6947, new_n6948, new_n6949, new_n6950,
    new_n6951, new_n6952, new_n6953, new_n6954, new_n6955, new_n6956,
    new_n6957, new_n6958, new_n6959, new_n6960, new_n6961, new_n6962,
    new_n6963, new_n6964, new_n6965, new_n6966, new_n6967, new_n6968,
    new_n6969, new_n6970, new_n6971, new_n6972, new_n6973, new_n6974,
    new_n6975, new_n6976, new_n6977, new_n6978, new_n6979, new_n6980,
    new_n6981, new_n6982, new_n6983, new_n6984, new_n6985, new_n6986,
    new_n6987, new_n6988, new_n6989, new_n6990, new_n6991, new_n6992,
    new_n6993, new_n6994, new_n6995, new_n6996, new_n6997, new_n6998,
    new_n6999, new_n7000, new_n7001, new_n7002, new_n7003, new_n7004,
    new_n7005, new_n7006, new_n7007, new_n7008, new_n7009, new_n7010,
    new_n7011, new_n7012, new_n7013, new_n7014, new_n7015, new_n7016,
    new_n7017, new_n7018, new_n7019, new_n7020, new_n7021, new_n7022,
    new_n7023, new_n7024, new_n7025, new_n7026, new_n7027, new_n7028,
    new_n7029, new_n7030, new_n7031, new_n7032, new_n7033, new_n7034,
    new_n7035, new_n7036, new_n7037, new_n7038, new_n7039, new_n7040,
    new_n7041, new_n7042, new_n7043, new_n7044, new_n7045, new_n7046,
    new_n7047, new_n7048, new_n7049, new_n7050, new_n7051, new_n7052,
    new_n7053, new_n7054, new_n7055, new_n7056, new_n7057, new_n7058,
    new_n7059, new_n7060, new_n7061, new_n7062, new_n7063, new_n7064,
    new_n7065, new_n7066, new_n7067, new_n7068, new_n7069, new_n7070,
    new_n7071, new_n7072, new_n7073, new_n7074, new_n7075, new_n7076,
    new_n7077, new_n7078, new_n7079, new_n7080, new_n7081, new_n7082,
    new_n7083, new_n7084, new_n7085, new_n7086, new_n7087, new_n7088,
    new_n7089, new_n7090, new_n7091, new_n7092, new_n7093, new_n7094,
    new_n7095, new_n7096, new_n7097, new_n7098, new_n7099, new_n7100,
    new_n7101, new_n7102, new_n7103, new_n7104, new_n7105, new_n7106,
    new_n7107, new_n7108, new_n7109, new_n7110, new_n7111, new_n7112,
    new_n7113, new_n7114, new_n7115, new_n7116, new_n7117, new_n7118,
    new_n7119, new_n7120, new_n7121, new_n7122, new_n7123, new_n7124,
    new_n7125, new_n7126, new_n7127, new_n7128, new_n7129, new_n7130,
    new_n7131, new_n7132, new_n7133, new_n7134, new_n7135, new_n7136,
    new_n7137, new_n7138, new_n7139, new_n7140, new_n7141, new_n7142,
    new_n7143, new_n7144, new_n7145, new_n7146, new_n7147, new_n7148,
    new_n7149, new_n7150, new_n7151, new_n7152, new_n7153, new_n7154,
    new_n7155, new_n7156, new_n7157, new_n7158, new_n7159, new_n7160,
    new_n7161, new_n7162, new_n7163, new_n7164, new_n7165, new_n7166,
    new_n7167, new_n7168, new_n7169, new_n7170, new_n7171, new_n7172,
    new_n7173, new_n7174, new_n7175, new_n7176, new_n7177, new_n7178,
    new_n7179, new_n7180, new_n7181, new_n7182, new_n7183, new_n7184,
    new_n7185, new_n7186, new_n7187, new_n7188, new_n7189, new_n7190,
    new_n7191, new_n7192, new_n7193, new_n7194, new_n7195, new_n7196,
    new_n7197, new_n7198, new_n7199, new_n7200, new_n7201, new_n7202,
    new_n7203, new_n7204, new_n7205, new_n7206, new_n7207, new_n7208,
    new_n7209, new_n7210, new_n7211, new_n7212, new_n7213, new_n7214,
    new_n7215, new_n7216, new_n7217, new_n7218, new_n7219, new_n7220,
    new_n7221, new_n7222, new_n7223, new_n7224, new_n7225, new_n7226,
    new_n7227, new_n7228, new_n7229, new_n7230, new_n7231, new_n7232,
    new_n7233, new_n7234, new_n7235, new_n7236, new_n7237, new_n7238,
    new_n7239, new_n7240, new_n7241, new_n7242, new_n7243, new_n7244,
    new_n7245, new_n7246, new_n7247, new_n7248, new_n7249, new_n7250,
    new_n7251, new_n7252, new_n7253, new_n7254, new_n7255, new_n7256,
    new_n7257, new_n7258, new_n7259, new_n7260, new_n7261, new_n7262,
    new_n7263, new_n7264, new_n7265, new_n7266, new_n7267, new_n7268,
    new_n7269, new_n7270, new_n7271, new_n7272, new_n7273, new_n7274,
    new_n7275, new_n7276, new_n7277, new_n7278, new_n7279, new_n7280,
    new_n7281, new_n7282, new_n7283, new_n7284, new_n7285, new_n7286,
    new_n7287, new_n7288, new_n7289, new_n7290, new_n7291, new_n7292,
    new_n7293, new_n7294, new_n7295, new_n7296, new_n7297, new_n7298,
    new_n7299, new_n7300, new_n7301, new_n7302, new_n7303, new_n7304,
    new_n7305, new_n7306, new_n7307, new_n7308, new_n7309, new_n7310,
    new_n7311, new_n7312, new_n7313, new_n7314, new_n7315, new_n7316,
    new_n7317, new_n7318, new_n7319, new_n7320, new_n7321, new_n7322,
    new_n7323, new_n7324, new_n7325, new_n7326, new_n7327, new_n7328,
    new_n7329, new_n7330, new_n7331, new_n7332, new_n7333, new_n7334,
    new_n7335, new_n7336, new_n7337, new_n7338, new_n7339, new_n7340,
    new_n7341, new_n7342, new_n7343, new_n7344, new_n7345, new_n7346,
    new_n7347, new_n7348, new_n7349, new_n7350, new_n7351, new_n7352,
    new_n7353, new_n7354, new_n7355, new_n7356, new_n7357, new_n7358,
    new_n7359, new_n7360, new_n7361, new_n7362, new_n7363, new_n7364,
    new_n7365, new_n7366, new_n7367, new_n7368, new_n7369, new_n7370,
    new_n7371, new_n7372, new_n7373, new_n7374, new_n7375, new_n7376,
    new_n7377, new_n7378, new_n7379, new_n7380, new_n7381, new_n7382,
    new_n7383, new_n7384, new_n7385, new_n7386, new_n7387, new_n7388,
    new_n7389, new_n7390, new_n7391, new_n7392, new_n7393, new_n7394,
    new_n7395, new_n7396, new_n7397, new_n7398, new_n7399, new_n7400,
    new_n7401, new_n7402, new_n7403, new_n7404, new_n7405, new_n7406,
    new_n7407, new_n7408, new_n7409, new_n7410, new_n7411, new_n7412,
    new_n7413, new_n7414, new_n7415, new_n7416, new_n7417, new_n7418,
    new_n7419, new_n7420, new_n7421, new_n7422, new_n7423, new_n7424,
    new_n7425, new_n7426, new_n7427, new_n7428, new_n7429, new_n7430,
    new_n7431, new_n7432, new_n7433, new_n7434, new_n7435, new_n7436,
    new_n7437, new_n7438, new_n7439, new_n7440, new_n7441, new_n7442,
    new_n7443, new_n7444, new_n7445, new_n7446, new_n7447, new_n7448,
    new_n7449, new_n7450, new_n7451, new_n7452, new_n7453, new_n7454,
    new_n7455, new_n7456, new_n7457, new_n7458, new_n7459, new_n7460,
    new_n7461, new_n7462, new_n7463, new_n7464, new_n7465, new_n7466,
    new_n7467, new_n7468, new_n7469, new_n7470, new_n7471, new_n7472,
    new_n7473, new_n7474, new_n7475, new_n7476, new_n7477, new_n7478,
    new_n7479, new_n7480, new_n7481, new_n7482, new_n7483, new_n7484,
    new_n7485, new_n7486, new_n7487, new_n7488, new_n7489, new_n7490,
    new_n7491, new_n7492, new_n7493, new_n7494, new_n7495, new_n7496,
    new_n7497, new_n7498, new_n7499, new_n7500, new_n7501, new_n7502,
    new_n7503, new_n7504, new_n7505, new_n7506, new_n7507, new_n7508,
    new_n7509, new_n7510, new_n7511, new_n7512, new_n7513, new_n7514,
    new_n7515, new_n7516, new_n7517, new_n7518, new_n7519, new_n7520,
    new_n7521, new_n7522, new_n7523, new_n7524, new_n7525, new_n7526,
    new_n7527, new_n7528, new_n7529, new_n7530, new_n7531, new_n7532,
    new_n7533, new_n7534, new_n7535, new_n7536, new_n7537, new_n7538,
    new_n7539, new_n7540, new_n7541, new_n7542, new_n7543, new_n7544,
    new_n7545, new_n7546, new_n7547, new_n7548, new_n7549, new_n7550,
    new_n7551, new_n7552, new_n7553, new_n7554, new_n7555, new_n7556,
    new_n7557, new_n7558, new_n7559, new_n7560, new_n7561, new_n7562,
    new_n7563, new_n7564, new_n7565, new_n7566, new_n7567, new_n7568,
    new_n7569, new_n7570, new_n7571, new_n7572, new_n7573, new_n7574,
    new_n7575, new_n7576, new_n7577, new_n7578, new_n7579, new_n7580,
    new_n7581, new_n7582, new_n7583, new_n7584, new_n7585, new_n7586,
    new_n7587, new_n7588, new_n7589, new_n7590, new_n7591, new_n7592,
    new_n7593, new_n7594, new_n7595, new_n7596, new_n7597, new_n7598,
    new_n7599, new_n7600, new_n7601, new_n7602, new_n7603, new_n7604,
    new_n7605, new_n7606, new_n7607, new_n7608, new_n7609, new_n7610,
    new_n7611, new_n7612, new_n7613, new_n7614, new_n7615, new_n7616,
    new_n7617, new_n7618, new_n7619, new_n7620, new_n7621, new_n7622,
    new_n7623, new_n7624, new_n7625, new_n7626, new_n7627, new_n7628,
    new_n7629, new_n7630, new_n7631, new_n7632, new_n7633, new_n7634,
    new_n7635, new_n7636, new_n7637, new_n7638, new_n7639, new_n7640,
    new_n7641, new_n7642, new_n7643, new_n7644, new_n7645, new_n7646,
    new_n7647, new_n7648, new_n7649, new_n7650, new_n7651, new_n7652,
    new_n7653, new_n7654, new_n7655, new_n7656, new_n7657, new_n7658,
    new_n7659, new_n7660, new_n7661, new_n7662, new_n7663, new_n7664,
    new_n7665, new_n7666, new_n7667, new_n7668, new_n7669, new_n7670,
    new_n7671, new_n7672, new_n7673, new_n7674, new_n7675, new_n7676,
    new_n7677, new_n7678, new_n7679, new_n7680, new_n7681, new_n7682,
    new_n7683, new_n7684, new_n7685, new_n7686, new_n7687, new_n7688,
    new_n7689, new_n7690, new_n7691, new_n7692, new_n7693, new_n7694,
    new_n7695, new_n7696, new_n7697, new_n7698, new_n7699, new_n7700,
    new_n7701, new_n7702, new_n7703, new_n7704, new_n7705, new_n7706,
    new_n7707, new_n7708, new_n7709, new_n7710, new_n7711, new_n7712,
    new_n7713, new_n7714, new_n7715, new_n7716, new_n7717, new_n7718,
    new_n7719, new_n7720, new_n7721, new_n7722, new_n7723, new_n7724,
    new_n7725, new_n7726, new_n7727, new_n7728, new_n7729, new_n7730,
    new_n7731, new_n7732, new_n7733, new_n7734, new_n7735, new_n7736,
    new_n7737, new_n7738, new_n7739, new_n7740, new_n7741, new_n7742,
    new_n7743, new_n7744, new_n7745, new_n7746, new_n7747, new_n7748,
    new_n7749, new_n7750, new_n7751, new_n7752, new_n7753, new_n7754,
    new_n7755, new_n7756, new_n7757, new_n7758, new_n7759, new_n7760,
    new_n7761, new_n7762, new_n7763, new_n7764, new_n7765, new_n7766,
    new_n7767, new_n7768, new_n7769, new_n7770, new_n7771, new_n7772,
    new_n7773, new_n7774, new_n7775, new_n7776, new_n7777, new_n7778,
    new_n7779, new_n7780, new_n7781, new_n7782, new_n7783, new_n7784,
    new_n7785, new_n7786, new_n7787, new_n7788, new_n7789, new_n7790,
    new_n7791, new_n7792, new_n7793, new_n7794, new_n7795, new_n7796,
    new_n7797, new_n7798, new_n7799, new_n7800, new_n7801, new_n7802,
    new_n7803, new_n7804, new_n7805, new_n7806, new_n7807, new_n7808,
    new_n7809, new_n7810, new_n7811, new_n7812, new_n7813, new_n7814,
    new_n7815, new_n7816, new_n7817, new_n7818, new_n7819, new_n7820,
    new_n7821, new_n7822, new_n7823, new_n7824, new_n7825, new_n7826,
    new_n7827, new_n7828, new_n7829, new_n7830, new_n7831, new_n7832,
    new_n7833, new_n7834, new_n7835, new_n7836, new_n7837, new_n7838,
    new_n7839, new_n7840, new_n7841, new_n7842, new_n7843, new_n7844,
    new_n7845, new_n7846, new_n7847, new_n7848, new_n7849, new_n7850,
    new_n7851, new_n7852, new_n7853, new_n7854, new_n7855, new_n7856,
    new_n7857, new_n7858, new_n7859, new_n7860, new_n7861, new_n7862,
    new_n7863, new_n7864, new_n7865, new_n7866, new_n7867, new_n7868,
    new_n7869, new_n7870, new_n7871, new_n7872, new_n7873, new_n7874,
    new_n7875, new_n7876, new_n7877, new_n7878, new_n7879, new_n7880,
    new_n7881, new_n7882, new_n7883, new_n7884, new_n7885, new_n7886,
    new_n7887, new_n7888, new_n7889, new_n7890, new_n7891, new_n7892,
    new_n7893, new_n7894, new_n7895, new_n7896, new_n7897, new_n7898,
    new_n7899, new_n7900, new_n7901, new_n7902, new_n7903, new_n7904,
    new_n7905, new_n7906, new_n7907, new_n7908, new_n7909, new_n7910,
    new_n7911, new_n7912, new_n7913, new_n7914, new_n7915, new_n7916,
    new_n7917, new_n7918, new_n7919, new_n7920, new_n7921, new_n7922,
    new_n7923, new_n7924, new_n7925, new_n7926, new_n7927, new_n7928,
    new_n7929, new_n7930, new_n7931, new_n7932, new_n7933, new_n7934,
    new_n7935, new_n7936, new_n7937, new_n7938, new_n7939, new_n7940,
    new_n7941, new_n7942, new_n7943, new_n7944, new_n7945, new_n7946,
    new_n7947, new_n7948, new_n7949, new_n7950, new_n7951, new_n7952,
    new_n7953, new_n7954, new_n7955, new_n7956, new_n7957, new_n7958,
    new_n7959, new_n7960, new_n7961, new_n7962, new_n7963, new_n7964,
    new_n7965, new_n7966, new_n7967, new_n7968, new_n7969, new_n7970,
    new_n7971, new_n7972, new_n7973, new_n7974, new_n7975, new_n7976,
    new_n7977, new_n7978, new_n7979, new_n7980, new_n7981, new_n7982,
    new_n7983, new_n7984, new_n7985, new_n7986, new_n7987, new_n7988,
    new_n7989, new_n7990, new_n7991, new_n7992, new_n7993, new_n7994,
    new_n7995, new_n7996, new_n7997, new_n7998, new_n7999, new_n8000,
    new_n8001, new_n8002, new_n8003, new_n8004, new_n8005, new_n8006,
    new_n8007, new_n8008, new_n8009, new_n8010, new_n8011, new_n8012,
    new_n8013, new_n8014, new_n8015, new_n8016, new_n8017, new_n8018,
    new_n8019, new_n8020, new_n8021, new_n8022, new_n8023, new_n8024,
    new_n8025, new_n8026, new_n8027, new_n8028, new_n8029, new_n8030,
    new_n8031, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036,
    new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042,
    new_n8043, new_n8044, new_n8045, new_n8046, new_n8047, new_n8048,
    new_n8049, new_n8050, new_n8051, new_n8052, new_n8053, new_n8054,
    new_n8055, new_n8056, new_n8057, new_n8058, new_n8059, new_n8060,
    new_n8061, new_n8062, new_n8063, new_n8064, new_n8065, new_n8066,
    new_n8067, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120,
    new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127, new_n8128, new_n8129, new_n8130, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135, new_n8136, new_n8137, new_n8138,
    new_n8139, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148, new_n8149, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215, new_n8216,
    new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228,
    new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234,
    new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244, new_n8245, new_n8246,
    new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252,
    new_n8253, new_n8254, new_n8255, new_n8256, new_n8257, new_n8258,
    new_n8259, new_n8260, new_n8261, new_n8262, new_n8263, new_n8264,
    new_n8265, new_n8266, new_n8267, new_n8268, new_n8269, new_n8270,
    new_n8271, new_n8272, new_n8273, new_n8274, new_n8275, new_n8276,
    new_n8277, new_n8278, new_n8279, new_n8280, new_n8281, new_n8282,
    new_n8283, new_n8284, new_n8285, new_n8286, new_n8287, new_n8288,
    new_n8289, new_n8290, new_n8291, new_n8292, new_n8293, new_n8294,
    new_n8295, new_n8296, new_n8297, new_n8298, new_n8299, new_n8300,
    new_n8301, new_n8302, new_n8303, new_n8304, new_n8305, new_n8306,
    new_n8307, new_n8308, new_n8309, new_n8310, new_n8311, new_n8312,
    new_n8313, new_n8314, new_n8315, new_n8316, new_n8317, new_n8318,
    new_n8319, new_n8320, new_n8321, new_n8322, new_n8323, new_n8324,
    new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330,
    new_n8331, new_n8332, new_n8333, new_n8334, new_n8335, new_n8336,
    new_n8337, new_n8338, new_n8339, new_n8340, new_n8341, new_n8342,
    new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348,
    new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354,
    new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360,
    new_n8361, new_n8362, new_n8363, new_n8364, new_n8365, new_n8366,
    new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372,
    new_n8373, new_n8374, new_n8375, new_n8376, new_n8377, new_n8378,
    new_n8379, new_n8380, new_n8381, new_n8382, new_n8383, new_n8384,
    new_n8385, new_n8386, new_n8387, new_n8388, new_n8389, new_n8390,
    new_n8391, new_n8392, new_n8393, new_n8394, new_n8395, new_n8396,
    new_n8397, new_n8398, new_n8399, new_n8400, new_n8401, new_n8402,
    new_n8403, new_n8404, new_n8405, new_n8406, new_n8407, new_n8408,
    new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414,
    new_n8415, new_n8416, new_n8417, new_n8418, new_n8419, new_n8420,
    new_n8421, new_n8422, new_n8423, new_n8424, new_n8425, new_n8426,
    new_n8427, new_n8428, new_n8429, new_n8430, new_n8431, new_n8432,
    new_n8433, new_n8434, new_n8435, new_n8436, new_n8437, new_n8438,
    new_n8439, new_n8440, new_n8441, new_n8442, new_n8443, new_n8444,
    new_n8445, new_n8446, new_n8447, new_n8448, new_n8449, new_n8450,
    new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456,
    new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462,
    new_n8463, new_n8464, new_n8465, new_n8466, new_n8467, new_n8468,
    new_n8469, new_n8470, new_n8471, new_n8472, new_n8473, new_n8474,
    new_n8475, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8637, new_n8638, new_n8639, new_n8640, new_n8641, new_n8642,
    new_n8643, new_n8644, new_n8645, new_n8646, new_n8647, new_n8648,
    new_n8649, new_n8650, new_n8651, new_n8652, new_n8653, new_n8654,
    new_n8655, new_n8656, new_n8657, new_n8658, new_n8659, new_n8660,
    new_n8661, new_n8662, new_n8663, new_n8664, new_n8665, new_n8666,
    new_n8667, new_n8668, new_n8669, new_n8670, new_n8671, new_n8672,
    new_n8673, new_n8674, new_n8675, new_n8676, new_n8677, new_n8678,
    new_n8679, new_n8680, new_n8681, new_n8682, new_n8683, new_n8684,
    new_n8685, new_n8686, new_n8687, new_n8688, new_n8689, new_n8690,
    new_n8691, new_n8692, new_n8693, new_n8694, new_n8695, new_n8696,
    new_n8697, new_n8698, new_n8699, new_n8700, new_n8701, new_n8702,
    new_n8703, new_n8704, new_n8705, new_n8706, new_n8707, new_n8708,
    new_n8709, new_n8710, new_n8711, new_n8712, new_n8713, new_n8714,
    new_n8715, new_n8716, new_n8717, new_n8718, new_n8719, new_n8720,
    new_n8721, new_n8722, new_n8723, new_n8724, new_n8725, new_n8726,
    new_n8727, new_n8728, new_n8729, new_n8730, new_n8731, new_n8732,
    new_n8733, new_n8734, new_n8735, new_n8736, new_n8737, new_n8738,
    new_n8739, new_n8740, new_n8741, new_n8742, new_n8743, new_n8744,
    new_n8745, new_n8746, new_n8747, new_n8748, new_n8749, new_n8750,
    new_n8751, new_n8752, new_n8753, new_n8754, new_n8755, new_n8756,
    new_n8757, new_n8758, new_n8759, new_n8760, new_n8761, new_n8762,
    new_n8763, new_n8764, new_n8765, new_n8766, new_n8767, new_n8768,
    new_n8769, new_n8770, new_n8771, new_n8772, new_n8773, new_n8774,
    new_n8775, new_n8776, new_n8777, new_n8778, new_n8779, new_n8780,
    new_n8781, new_n8782, new_n8783, new_n8784, new_n8785, new_n8786,
    new_n8787, new_n8788, new_n8789, new_n8790, new_n8791, new_n8792,
    new_n8793, new_n8794, new_n8795, new_n8796, new_n8797, new_n8798,
    new_n8799, new_n8800, new_n8801, new_n8802, new_n8803, new_n8804,
    new_n8805, new_n8806, new_n8807, new_n8808, new_n8809, new_n8810,
    new_n8811, new_n8812, new_n8813, new_n8814, new_n8815, new_n8816,
    new_n8817, new_n8818, new_n8819, new_n8820, new_n8821, new_n8822,
    new_n8823, new_n8824, new_n8825, new_n8826, new_n8827, new_n8828,
    new_n8829, new_n8830, new_n8831, new_n8832, new_n8833, new_n8834,
    new_n8835, new_n8836, new_n8837, new_n8838, new_n8839, new_n8840,
    new_n8841, new_n8842, new_n8843, new_n8844, new_n8845, new_n8846,
    new_n8847, new_n8848, new_n8849, new_n8850, new_n8851, new_n8852,
    new_n8853, new_n8854, new_n8855, new_n8856, new_n8857, new_n8858,
    new_n8859, new_n8860, new_n8861, new_n8862, new_n8863, new_n8864,
    new_n8865, new_n8866, new_n8867, new_n8868, new_n8869, new_n8870,
    new_n8871, new_n8872, new_n8873, new_n8874, new_n8875, new_n8876,
    new_n8877, new_n8878, new_n8879, new_n8880, new_n8881, new_n8882,
    new_n8883, new_n8884, new_n8885, new_n8886, new_n8887, new_n8888,
    new_n8889, new_n8890, new_n8891, new_n8892, new_n8893, new_n8894,
    new_n8895, new_n8896, new_n8897, new_n8898, new_n8899, new_n8900,
    new_n8901, new_n8902, new_n8903, new_n8904, new_n8905, new_n8906,
    new_n8907, new_n8908, new_n8909, new_n8910, new_n8911, new_n8912,
    new_n8913, new_n8914, new_n8915, new_n8916, new_n8917, new_n8918,
    new_n8919, new_n8920, new_n8921, new_n8922, new_n8923, new_n8924,
    new_n8925, new_n8926, new_n8927, new_n8928, new_n8929, new_n8930,
    new_n8931, new_n8932, new_n8933, new_n8934, new_n8935, new_n8936,
    new_n8937, new_n8938, new_n8939, new_n8940, new_n8941, new_n8942,
    new_n8943, new_n8944, new_n8945, new_n8946, new_n8947, new_n8948,
    new_n8949, new_n8950, new_n8951, new_n8952, new_n8953, new_n8954,
    new_n8955, new_n8956, new_n8957, new_n8958, new_n8959, new_n8960,
    new_n8961, new_n8962, new_n8963, new_n8964, new_n8965, new_n8966,
    new_n8967, new_n8968, new_n8969, new_n8970, new_n8971, new_n8972,
    new_n8973, new_n8974, new_n8975, new_n8976, new_n8977, new_n8978,
    new_n8979, new_n8980, new_n8981, new_n8982, new_n8983, new_n8984,
    new_n8985, new_n8986, new_n8987, new_n8988, new_n8989, new_n8990,
    new_n8991, new_n8992, new_n8993, new_n8994, new_n8995, new_n8996,
    new_n8997, new_n8998, new_n8999, new_n9000, new_n9001, new_n9002,
    new_n9003, new_n9004, new_n9005, new_n9006, new_n9007, new_n9008,
    new_n9009, new_n9010, new_n9011, new_n9012, new_n9013, new_n9014,
    new_n9015, new_n9016, new_n9017, new_n9018, new_n9019, new_n9020,
    new_n9021, new_n9022, new_n9023, new_n9024, new_n9025, new_n9026,
    new_n9027, new_n9028, new_n9029, new_n9030, new_n9031, new_n9032,
    new_n9033, new_n9034, new_n9035, new_n9036, new_n9037, new_n9038,
    new_n9039, new_n9040, new_n9041, new_n9042, new_n9043, new_n9044,
    new_n9045, new_n9046, new_n9047, new_n9048, new_n9049, new_n9050,
    new_n9051, new_n9052, new_n9053, new_n9054, new_n9055, new_n9056,
    new_n9057, new_n9058, new_n9059, new_n9060, new_n9061, new_n9062,
    new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068,
    new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074,
    new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080,
    new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086,
    new_n9087, new_n9088, new_n9089, new_n9090, new_n9091, new_n9092,
    new_n9093, new_n9094, new_n9095, new_n9096, new_n9097, new_n9098,
    new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104,
    new_n9105, new_n9106, new_n9107, new_n9108, new_n9109, new_n9110,
    new_n9111, new_n9112, new_n9113, new_n9114, new_n9115, new_n9116,
    new_n9117, new_n9118, new_n9119, new_n9120, new_n9121, new_n9122,
    new_n9123, new_n9124, new_n9125, new_n9126, new_n9127, new_n9128,
    new_n9129, new_n9130, new_n9131, new_n9132, new_n9133, new_n9134,
    new_n9135, new_n9136, new_n9137, new_n9138, new_n9139, new_n9140,
    new_n9141, new_n9142, new_n9143, new_n9144, new_n9145, new_n9146,
    new_n9147, new_n9148, new_n9149, new_n9150, new_n9151, new_n9152,
    new_n9153, new_n9154, new_n9155, new_n9156, new_n9157, new_n9158,
    new_n9159, new_n9160, new_n9161, new_n9162, new_n9163, new_n9164,
    new_n9165, new_n9166, new_n9167, new_n9168, new_n9169, new_n9170,
    new_n9171, new_n9172, new_n9173, new_n9174, new_n9175, new_n9176,
    new_n9177, new_n9178, new_n9179, new_n9180, new_n9181, new_n9182,
    new_n9183, new_n9184, new_n9185, new_n9186, new_n9187, new_n9188,
    new_n9189, new_n9190, new_n9191, new_n9192, new_n9193, new_n9194,
    new_n9195, new_n9196, new_n9197, new_n9198, new_n9199, new_n9200,
    new_n9201, new_n9202, new_n9203, new_n9204, new_n9205, new_n9206,
    new_n9207, new_n9208, new_n9209, new_n9210, new_n9211, new_n9212,
    new_n9213, new_n9214, new_n9215, new_n9216, new_n9217, new_n9218,
    new_n9219, new_n9220, new_n9221, new_n9222, new_n9223, new_n9224,
    new_n9225, new_n9226, new_n9227, new_n9228, new_n9229, new_n9230,
    new_n9231, new_n9232, new_n9233, new_n9234, new_n9235, new_n9236,
    new_n9237, new_n9238, new_n9239, new_n9240, new_n9241, new_n9242,
    new_n9243, new_n9244, new_n9245, new_n9246, new_n9247, new_n9248,
    new_n9249, new_n9250, new_n9251, new_n9252, new_n9253, new_n9254,
    new_n9255, new_n9256, new_n9257, new_n9258, new_n9259, new_n9260,
    new_n9261, new_n9262, new_n9263, new_n9264, new_n9265, new_n9266,
    new_n9267, new_n9268, new_n9269, new_n9270, new_n9271, new_n9272,
    new_n9273, new_n9274, new_n9275, new_n9276, new_n9277, new_n9278,
    new_n9279, new_n9280, new_n9281, new_n9282, new_n9283, new_n9284,
    new_n9285, new_n9286, new_n9287, new_n9288, new_n9289, new_n9290,
    new_n9291, new_n9292, new_n9293, new_n9294, new_n9295, new_n9296,
    new_n9297, new_n9298, new_n9299, new_n9300, new_n9301, new_n9302,
    new_n9303, new_n9304, new_n9305, new_n9306, new_n9307, new_n9308,
    new_n9309, new_n9310, new_n9311, new_n9312, new_n9313, new_n9314,
    new_n9315, new_n9316, new_n9317, new_n9318, new_n9319, new_n9320,
    new_n9321, new_n9322, new_n9323, new_n9324, new_n9325, new_n9326,
    new_n9327, new_n9328, new_n9329, new_n9330, new_n9331, new_n9332,
    new_n9333, new_n9334, new_n9335, new_n9336, new_n9337, new_n9338,
    new_n9339, new_n9340, new_n9341, new_n9342, new_n9343, new_n9344,
    new_n9345, new_n9346, new_n9347, new_n9348, new_n9349, new_n9350,
    new_n9351, new_n9352, new_n9353, new_n9354, new_n9355, new_n9356,
    new_n9357, new_n9358, new_n9359, new_n9360, new_n9361, new_n9362,
    new_n9363, new_n9364, new_n9365, new_n9366, new_n9367, new_n9368,
    new_n9369, new_n9370, new_n9371, new_n9372, new_n9373, new_n9374,
    new_n9375, new_n9376, new_n9377, new_n9378, new_n9379, new_n9380,
    new_n9381, new_n9382, new_n9383, new_n9384, new_n9385, new_n9386,
    new_n9387, new_n9388, new_n9389, new_n9390, new_n9391, new_n9392,
    new_n9393, new_n9394, new_n9395, new_n9396, new_n9397, new_n9398,
    new_n9399, new_n9400, new_n9401, new_n9402, new_n9403, new_n9404,
    new_n9405, new_n9406, new_n9407, new_n9408, new_n9409, new_n9410,
    new_n9411, new_n9412, new_n9413, new_n9414, new_n9415, new_n9416,
    new_n9417, new_n9418, new_n9419, new_n9420, new_n9421, new_n9422,
    new_n9423, new_n9424, new_n9425, new_n9426, new_n9427, new_n9428,
    new_n9429, new_n9430, new_n9431, new_n9432, new_n9433, new_n9434,
    new_n9435, new_n9436, new_n9437, new_n9438, new_n9439, new_n9440,
    new_n9441, new_n9442, new_n9443, new_n9444, new_n9445, new_n9446,
    new_n9447, new_n9448, new_n9449, new_n9450, new_n9451, new_n9452,
    new_n9453, new_n9454, new_n9455, new_n9456, new_n9457, new_n9458,
    new_n9459, new_n9460, new_n9461, new_n9462, new_n9463, new_n9464,
    new_n9465, new_n9466, new_n9467, new_n9468, new_n9469, new_n9470,
    new_n9471, new_n9472, new_n9473, new_n9474, new_n9475, new_n9476,
    new_n9477, new_n9478, new_n9479, new_n9480, new_n9481, new_n9482,
    new_n9483, new_n9484, new_n9485, new_n9486, new_n9487, new_n9488,
    new_n9489, new_n9490, new_n9491, new_n9492, new_n9493, new_n9494,
    new_n9495, new_n9496, new_n9497, new_n9498, new_n9499, new_n9500,
    new_n9501, new_n9502, new_n9503, new_n9504, new_n9505, new_n9506,
    new_n9507, new_n9508, new_n9509, new_n9510, new_n9511, new_n9512,
    new_n9513, new_n9514, new_n9515, new_n9516, new_n9517, new_n9518,
    new_n9519, new_n9520, new_n9521, new_n9522, new_n9523, new_n9524,
    new_n9525, new_n9526, new_n9527, new_n9528, new_n9529, new_n9530,
    new_n9531, new_n9532, new_n9533, new_n9534, new_n9535, new_n9536,
    new_n9537, new_n9538, new_n9539, new_n9540, new_n9541, new_n9542,
    new_n9543, new_n9544, new_n9545, new_n9546, new_n9547, new_n9548,
    new_n9549, new_n9550, new_n9551, new_n9552, new_n9553, new_n9554,
    new_n9555, new_n9556, new_n9557, new_n9558, new_n9559, new_n9560,
    new_n9561, new_n9562, new_n9563, new_n9564, new_n9565, new_n9566,
    new_n9567, new_n9568, new_n9569, new_n9570, new_n9571, new_n9572,
    new_n9573, new_n9574, new_n9575, new_n9576, new_n9577, new_n9578,
    new_n9579, new_n9580, new_n9581, new_n9582, new_n9583, new_n9584,
    new_n9585, new_n9586, new_n9587, new_n9588, new_n9589, new_n9590,
    new_n9591, new_n9592, new_n9593, new_n9594, new_n9595, new_n9596,
    new_n9597, new_n9598, new_n9599, new_n9600, new_n9601, new_n9602,
    new_n9603, new_n9604, new_n9605, new_n9606, new_n9607, new_n9608,
    new_n9609, new_n9610, new_n9611, new_n9612, new_n9613, new_n9614,
    new_n9615, new_n9616, new_n9617, new_n9618, new_n9619, new_n9620,
    new_n9621, new_n9622, new_n9623, new_n9624, new_n9625, new_n9626,
    new_n9627, new_n9628, new_n9629, new_n9630, new_n9631, new_n9632,
    new_n9633, new_n9634, new_n9635, new_n9636, new_n9637, new_n9638,
    new_n9639, new_n9640, new_n9641, new_n9642, new_n9643, new_n9644,
    new_n9645, new_n9646, new_n9647, new_n9648, new_n9649, new_n9650,
    new_n9651, new_n9652, new_n9653, new_n9654, new_n9655, new_n9656,
    new_n9657, new_n9658, new_n9659, new_n9660, new_n9661, new_n9662,
    new_n9663, new_n9664, new_n9665, new_n9666, new_n9667, new_n9668,
    new_n9669, new_n9670, new_n9671, new_n9672, new_n9673, new_n9674,
    new_n9675, new_n9676, new_n9677, new_n9678, new_n9679, new_n9680,
    new_n9681, new_n9682, new_n9683, new_n9684, new_n9685, new_n9686,
    new_n9687, new_n9688, new_n9689, new_n9690, new_n9691, new_n9692,
    new_n9693, new_n9694, new_n9695, new_n9696, new_n9697, new_n9698,
    new_n9699, new_n9700, new_n9701, new_n9702, new_n9703, new_n9704,
    new_n9705, new_n9706, new_n9707, new_n9708, new_n9709, new_n9710,
    new_n9711, new_n9712, new_n9713, new_n9714, new_n9715, new_n9716,
    new_n9717, new_n9718, new_n9719, new_n9720, new_n9721, new_n9722,
    new_n9723, new_n9724, new_n9725, new_n9726, new_n9727, new_n9728,
    new_n9729, new_n9730, new_n9731, new_n9732, new_n9733, new_n9734,
    new_n9735, new_n9736, new_n9737, new_n9738, new_n9739, new_n9740,
    new_n9741, new_n9742, new_n9743, new_n9744, new_n9745, new_n9746,
    new_n9747, new_n9748, new_n9749, new_n9750, new_n9751, new_n9752,
    new_n9753, new_n9754, new_n9755, new_n9756, new_n9757, new_n9758,
    new_n9759, new_n9760, new_n9761, new_n9762, new_n9763, new_n9764,
    new_n9765, new_n9766, new_n9767, new_n9768, new_n9769, new_n9770,
    new_n9771, new_n9772, new_n9773, new_n9774, new_n9775, new_n9776,
    new_n9777, new_n9778, new_n9779, new_n9780, new_n9781, new_n9782,
    new_n9783, new_n9784, new_n9785, new_n9786, new_n9787, new_n9788,
    new_n9789, new_n9790, new_n9791, new_n9792, new_n9793, new_n9794,
    new_n9795, new_n9796, new_n9797, new_n9798, new_n9799, new_n9800,
    new_n9801, new_n9802, new_n9803, new_n9804, new_n9805, new_n9806,
    new_n9807, new_n9808, new_n9809, new_n9810, new_n9811, new_n9812,
    new_n9813, new_n9814, new_n9815, new_n9816, new_n9817, new_n9818,
    new_n9819, new_n9820, new_n9821, new_n9822, new_n9823, new_n9824,
    new_n9825, new_n9826, new_n9827, new_n9828, new_n9829, new_n9830,
    new_n9831, new_n9832, new_n9833, new_n9834, new_n9835, new_n9836,
    new_n9837, new_n9838, new_n9839, new_n9840, new_n9841, new_n9842,
    new_n9843, new_n9844, new_n9845, new_n9846, new_n9847, new_n9848,
    new_n9849, new_n9850, new_n9851, new_n9852, new_n9853, new_n9854,
    new_n9855, new_n9856, new_n9857, new_n9858, new_n9859, new_n9860,
    new_n9861, new_n9862, new_n9863, new_n9864, new_n9865, new_n9866,
    new_n9867, new_n9868, new_n9869, new_n9870, new_n9871, new_n9872,
    new_n9873, new_n9874, new_n9875, new_n9876, new_n9877, new_n9878,
    new_n9879, new_n9880, new_n9881, new_n9882, new_n9883, new_n9884,
    new_n9885, new_n9886, new_n9887, new_n9888, new_n9889, new_n9890,
    new_n9891, new_n9892, new_n9893, new_n9894, new_n9895, new_n9896,
    new_n9897, new_n9898, new_n9899, new_n9900, new_n9901, new_n9902,
    new_n9903, new_n9904, new_n9905, new_n9906, new_n9907, new_n9908,
    new_n9909, new_n9910, new_n9911, new_n9912, new_n9913, new_n9914,
    new_n9915, new_n9916, new_n9917, new_n9918, new_n9919, new_n9920,
    new_n9921, new_n9922, new_n9923, new_n9924, new_n9925, new_n9926,
    new_n9927, new_n9928, new_n9929, new_n9930, new_n9931, new_n9932,
    new_n9933, new_n9934, new_n9935, new_n9936, new_n9937, new_n9938,
    new_n9939, new_n9940, new_n9941, new_n9942, new_n9943, new_n9944,
    new_n9945, new_n9946, new_n9947, new_n9948, new_n9949, new_n9950,
    new_n9951, new_n9952, new_n9953, new_n9954, new_n9955, new_n9956,
    new_n9957, new_n9958, new_n9959, new_n9960, new_n9961, new_n9962,
    new_n9963, new_n9964, new_n9965, new_n9966, new_n9967, new_n9968,
    new_n9969, new_n9970, new_n9971, new_n9972, new_n9973, new_n9974,
    new_n9975, new_n9976, new_n9977, new_n9978, new_n9979, new_n9980,
    new_n9981, new_n9982, new_n9983, new_n9984, new_n9985, new_n9986,
    new_n9987, new_n9988, new_n9989, new_n9990, new_n9991, new_n9992,
    new_n9993, new_n9994, new_n9995, new_n9996, new_n9997, new_n9998,
    new_n9999, new_n10000, new_n10001, new_n10002, new_n10003, new_n10004,
    new_n10005, new_n10006, new_n10007, new_n10008, new_n10009, new_n10010,
    new_n10011, new_n10012, new_n10013, new_n10014, new_n10015, new_n10016,
    new_n10017, new_n10018, new_n10019, new_n10020, new_n10021, new_n10022,
    new_n10023, new_n10024, new_n10025, new_n10026, new_n10027, new_n10028,
    new_n10029, new_n10030, new_n10031, new_n10032, new_n10033, new_n10034,
    new_n10035, new_n10036, new_n10037, new_n10038, new_n10039, new_n10040,
    new_n10041, new_n10042, new_n10043, new_n10044, new_n10045, new_n10046,
    new_n10047, new_n10048, new_n10049, new_n10050, new_n10051, new_n10052,
    new_n10053, new_n10054, new_n10055, new_n10056, new_n10057, new_n10058,
    new_n10059, new_n10060, new_n10061, new_n10062, new_n10063, new_n10064,
    new_n10065, new_n10066, new_n10067, new_n10068, new_n10069, new_n10070,
    new_n10071, new_n10072, new_n10073, new_n10074, new_n10075, new_n10076,
    new_n10077, new_n10078, new_n10079, new_n10080, new_n10081, new_n10082,
    new_n10083, new_n10084, new_n10085, new_n10086, new_n10087, new_n10088,
    new_n10089, new_n10090, new_n10091, new_n10092, new_n10093, new_n10094,
    new_n10095, new_n10096, new_n10097, new_n10098, new_n10099, new_n10100,
    new_n10101, new_n10102, new_n10103, new_n10104, new_n10105, new_n10106,
    new_n10107, new_n10108, new_n10109, new_n10110, new_n10111, new_n10112,
    new_n10113, new_n10114, new_n10115, new_n10116, new_n10117, new_n10118,
    new_n10119, new_n10120, new_n10121, new_n10122, new_n10123, new_n10124,
    new_n10125, new_n10126, new_n10127, new_n10128, new_n10129, new_n10130,
    new_n10131, new_n10132, new_n10133, new_n10134, new_n10135, new_n10136,
    new_n10137, new_n10138, new_n10139, new_n10140, new_n10141, new_n10142,
    new_n10143, new_n10144, new_n10145, new_n10146, new_n10147, new_n10148,
    new_n10149, new_n10150, new_n10151, new_n10152, new_n10153, new_n10154,
    new_n10155, new_n10156, new_n10157, new_n10158, new_n10159, new_n10160,
    new_n10161, new_n10162, new_n10163, new_n10164, new_n10165, new_n10166,
    new_n10167, new_n10168, new_n10169, new_n10170, new_n10171, new_n10172,
    new_n10173, new_n10174, new_n10175, new_n10176, new_n10177, new_n10178,
    new_n10179, new_n10180, new_n10181, new_n10182, new_n10183, new_n10184,
    new_n10185, new_n10186, new_n10187, new_n10188, new_n10189, new_n10190,
    new_n10191, new_n10192, new_n10193, new_n10194, new_n10195, new_n10196,
    new_n10197, new_n10198, new_n10199, new_n10200, new_n10201, new_n10202,
    new_n10203, new_n10204, new_n10205, new_n10206, new_n10207, new_n10208,
    new_n10209, new_n10210, new_n10211, new_n10212, new_n10213, new_n10214,
    new_n10215, new_n10216, new_n10217, new_n10218, new_n10219, new_n10220,
    new_n10221, new_n10222, new_n10223, new_n10224, new_n10225, new_n10226,
    new_n10227, new_n10228, new_n10229, new_n10230, new_n10231, new_n10232,
    new_n10233, new_n10234, new_n10235, new_n10236, new_n10237, new_n10238,
    new_n10239, new_n10240, new_n10241, new_n10242, new_n10243, new_n10244,
    new_n10245, new_n10246, new_n10247, new_n10248, new_n10249, new_n10250,
    new_n10251, new_n10252, new_n10253, new_n10254, new_n10255, new_n10256,
    new_n10257, new_n10258, new_n10259, new_n10260, new_n10261, new_n10262,
    new_n10263, new_n10264, new_n10265, new_n10266, new_n10267, new_n10268,
    new_n10269, new_n10270, new_n10271, new_n10272, new_n10273, new_n10274,
    new_n10275, new_n10276, new_n10277, new_n10278, new_n10279, new_n10280,
    new_n10281, new_n10282, new_n10283, new_n10284, new_n10285, new_n10286,
    new_n10287, new_n10288, new_n10289, new_n10290, new_n10291, new_n10292,
    new_n10293, new_n10294, new_n10295, new_n10296, new_n10297, new_n10298,
    new_n10299, new_n10300, new_n10301, new_n10302, new_n10303, new_n10304,
    new_n10305, new_n10306, new_n10307, new_n10308, new_n10309, new_n10310,
    new_n10311, new_n10312, new_n10313, new_n10314, new_n10315, new_n10316,
    new_n10317, new_n10318, new_n10319, new_n10320, new_n10321, new_n10322,
    new_n10323, new_n10324, new_n10325, new_n10326, new_n10327, new_n10328,
    new_n10329, new_n10330, new_n10331, new_n10332, new_n10333, new_n10334,
    new_n10335, new_n10336, new_n10337, new_n10338, new_n10339, new_n10340,
    new_n10341, new_n10342, new_n10343, new_n10344, new_n10345, new_n10346,
    new_n10347, new_n10348, new_n10349, new_n10350, new_n10351, new_n10352,
    new_n10353, new_n10354, new_n10355, new_n10356, new_n10357, new_n10358,
    new_n10359, new_n10360, new_n10361, new_n10362, new_n10363, new_n10364,
    new_n10365, new_n10366, new_n10367, new_n10368, new_n10369, new_n10370,
    new_n10371, new_n10372, new_n10373, new_n10374, new_n10375, new_n10376,
    new_n10377, new_n10378, new_n10379, new_n10380, new_n10381, new_n10382,
    new_n10383, new_n10384, new_n10385, new_n10386, new_n10387, new_n10388,
    new_n10389, new_n10390, new_n10391, new_n10392, new_n10393, new_n10394,
    new_n10395, new_n10396, new_n10397, new_n10398, new_n10399, new_n10400,
    new_n10401, new_n10402, new_n10403, new_n10404, new_n10405, new_n10406,
    new_n10407, new_n10408, new_n10409, new_n10410, new_n10411, new_n10412,
    new_n10413, new_n10414, new_n10415, new_n10416, new_n10417, new_n10418,
    new_n10419, new_n10420, new_n10421, new_n10422, new_n10423, new_n10424,
    new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430,
    new_n10431, new_n10432, new_n10433, new_n10434, new_n10435, new_n10436,
    new_n10437, new_n10438, new_n10439, new_n10440, new_n10441, new_n10442,
    new_n10443, new_n10444, new_n10445, new_n10446, new_n10447, new_n10448,
    new_n10449, new_n10450, new_n10451, new_n10452, new_n10453, new_n10454,
    new_n10455, new_n10456, new_n10457, new_n10458, new_n10459, new_n10460,
    new_n10461, new_n10462, new_n10463, new_n10464, new_n10465, new_n10466,
    new_n10467, new_n10468, new_n10469, new_n10470, new_n10471, new_n10472,
    new_n10473, new_n10474, new_n10475, new_n10476, new_n10477, new_n10478,
    new_n10479, new_n10480, new_n10481, new_n10482, new_n10483, new_n10484,
    new_n10485, new_n10486, new_n10487, new_n10488, new_n10489, new_n10490,
    new_n10491, new_n10492, new_n10493, new_n10494, new_n10495, new_n10496,
    new_n10497, new_n10498, new_n10499, new_n10500, new_n10501, new_n10502,
    new_n10503, new_n10504, new_n10505, new_n10506, new_n10507, new_n10508,
    new_n10509, new_n10510, new_n10511, new_n10512, new_n10513, new_n10514,
    new_n10515, new_n10516, new_n10517, new_n10518, new_n10519, new_n10520,
    new_n10521, new_n10522, new_n10523, new_n10524, new_n10525, new_n10526,
    new_n10527, new_n10528, new_n10529, new_n10530, new_n10531, new_n10532,
    new_n10533, new_n10534, new_n10535, new_n10536, new_n10537, new_n10538,
    new_n10539, new_n10540, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545, new_n10546, new_n10547, new_n10548, new_n10549, new_n10550,
    new_n10551, new_n10552, new_n10553, new_n10554, new_n10555, new_n10556,
    new_n10557, new_n10558, new_n10559, new_n10560, new_n10561, new_n10562,
    new_n10563, new_n10564, new_n10565, new_n10566, new_n10567, new_n10568,
    new_n10569, new_n10570, new_n10571, new_n10572, new_n10573, new_n10574,
    new_n10575, new_n10576, new_n10577, new_n10578, new_n10579, new_n10580,
    new_n10581, new_n10582, new_n10583, new_n10584, new_n10585, new_n10586,
    new_n10587, new_n10588, new_n10589, new_n10590, new_n10591, new_n10592,
    new_n10593, new_n10594, new_n10595, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10606, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611, new_n10612, new_n10613, new_n10614, new_n10615, new_n10616,
    new_n10617, new_n10618, new_n10619, new_n10620, new_n10621, new_n10622,
    new_n10623, new_n10624, new_n10625, new_n10626, new_n10627, new_n10628,
    new_n10629, new_n10630, new_n10631, new_n10632, new_n10633, new_n10634,
    new_n10635, new_n10636, new_n10637, new_n10638, new_n10639, new_n10640,
    new_n10641, new_n10642, new_n10643, new_n10644, new_n10645, new_n10646,
    new_n10647, new_n10648, new_n10649, new_n10650, new_n10651, new_n10652,
    new_n10653, new_n10654, new_n10655, new_n10656, new_n10657, new_n10658,
    new_n10659, new_n10660, new_n10661, new_n10662, new_n10663, new_n10664,
    new_n10665, new_n10666, new_n10667, new_n10668, new_n10669, new_n10670,
    new_n10671, new_n10672, new_n10673, new_n10674, new_n10675, new_n10676,
    new_n10677, new_n10678, new_n10679, new_n10680, new_n10681, new_n10682,
    new_n10683, new_n10684, new_n10685, new_n10686, new_n10687, new_n10688,
    new_n10689, new_n10690, new_n10691, new_n10692, new_n10693, new_n10694,
    new_n10695, new_n10696, new_n10697, new_n10698, new_n10699, new_n10700,
    new_n10701, new_n10702, new_n10703, new_n10704, new_n10705, new_n10706,
    new_n10707, new_n10708, new_n10709, new_n10710, new_n10711, new_n10712,
    new_n10713, new_n10714, new_n10715, new_n10716, new_n10717, new_n10718,
    new_n10719, new_n10720, new_n10721, new_n10722, new_n10723, new_n10724,
    new_n10725, new_n10726, new_n10727, new_n10728, new_n10729, new_n10730,
    new_n10731, new_n10732, new_n10733, new_n10734, new_n10735, new_n10736,
    new_n10737, new_n10738, new_n10739, new_n10740, new_n10741, new_n10742,
    new_n10743, new_n10744, new_n10745, new_n10746, new_n10747, new_n10748,
    new_n10749, new_n10750, new_n10751, new_n10752, new_n10753, new_n10754,
    new_n10755, new_n10756, new_n10757, new_n10758, new_n10759, new_n10760,
    new_n10761, new_n10762, new_n10763, new_n10764, new_n10765, new_n10766,
    new_n10767, new_n10768, new_n10769, new_n10770, new_n10771, new_n10772,
    new_n10773, new_n10774, new_n10775, new_n10776, new_n10777, new_n10778,
    new_n10779, new_n10780, new_n10781, new_n10782, new_n10783, new_n10784,
    new_n10785, new_n10786, new_n10787, new_n10788, new_n10789, new_n10790,
    new_n10791, new_n10792, new_n10793, new_n10794, new_n10795, new_n10796,
    new_n10797, new_n10798, new_n10799, new_n10800, new_n10801, new_n10802,
    new_n10803, new_n10804, new_n10805, new_n10806, new_n10807, new_n10808,
    new_n10809, new_n10810, new_n10811, new_n10812, new_n10813, new_n10814,
    new_n10815, new_n10816, new_n10817, new_n10818, new_n10819, new_n10820,
    new_n10821, new_n10822, new_n10823, new_n10824, new_n10825, new_n10826,
    new_n10827, new_n10828, new_n10829, new_n10830, new_n10831, new_n10832,
    new_n10833, new_n10834, new_n10835, new_n10836, new_n10837, new_n10838,
    new_n10839, new_n10840, new_n10841, new_n10842, new_n10843, new_n10844,
    new_n10845, new_n10846, new_n10847, new_n10848, new_n10849, new_n10850,
    new_n10851, new_n10852, new_n10853, new_n10854, new_n10855, new_n10856,
    new_n10857, new_n10858, new_n10859, new_n10860, new_n10861, new_n10862,
    new_n10863, new_n10864, new_n10865, new_n10866, new_n10867, new_n10868,
    new_n10869, new_n10870, new_n10871, new_n10872, new_n10873, new_n10874,
    new_n10875, new_n10876, new_n10877, new_n10878, new_n10879, new_n10880,
    new_n10881, new_n10882, new_n10883, new_n10884, new_n10885, new_n10886,
    new_n10887, new_n10888, new_n10889, new_n10890, new_n10891, new_n10892,
    new_n10893, new_n10894, new_n10895, new_n10896, new_n10897, new_n10898,
    new_n10899, new_n10900, new_n10901, new_n10902, new_n10903, new_n10904,
    new_n10905, new_n10906, new_n10907, new_n10908, new_n10909, new_n10910,
    new_n10911, new_n10912, new_n10913, new_n10914, new_n10915, new_n10916,
    new_n10917, new_n10918, new_n10919, new_n10920, new_n10921, new_n10922,
    new_n10923, new_n10924, new_n10925, new_n10926, new_n10927, new_n10928,
    new_n10929, new_n10930, new_n10931, new_n10932, new_n10933, new_n10934,
    new_n10935, new_n10936, new_n10937, new_n10938, new_n10939, new_n10940,
    new_n10941, new_n10942, new_n10943, new_n10944, new_n10945, new_n10946,
    new_n10947, new_n10948, new_n10949, new_n10950, new_n10951, new_n10952,
    new_n10953, new_n10954, new_n10955, new_n10956, new_n10957, new_n10958,
    new_n10959, new_n10960, new_n10961, new_n10962, new_n10963, new_n10964,
    new_n10965, new_n10966, new_n10967, new_n10968, new_n10969, new_n10970,
    new_n10971, new_n10972, new_n10973, new_n10974, new_n10975, new_n10976,
    new_n10977, new_n10978, new_n10979, new_n10980, new_n10981, new_n10982,
    new_n10983, new_n10984, new_n10985, new_n10986, new_n10987, new_n10988,
    new_n10989, new_n10990, new_n10991, new_n10992, new_n10993, new_n10994,
    new_n10995, new_n10996, new_n10997, new_n10998, new_n10999, new_n11000,
    new_n11001, new_n11002, new_n11003, new_n11004, new_n11005, new_n11006,
    new_n11007, new_n11008, new_n11009, new_n11010, new_n11011, new_n11012,
    new_n11013, new_n11014, new_n11015, new_n11016, new_n11017, new_n11018,
    new_n11019, new_n11020, new_n11021, new_n11022, new_n11023, new_n11024,
    new_n11025, new_n11026, new_n11027, new_n11028, new_n11029, new_n11030,
    new_n11031, new_n11032, new_n11033, new_n11034, new_n11035, new_n11036,
    new_n11037, new_n11038, new_n11039, new_n11040, new_n11041, new_n11042,
    new_n11043, new_n11044, new_n11045, new_n11046, new_n11047, new_n11048,
    new_n11049, new_n11050, new_n11051, new_n11052, new_n11053, new_n11054,
    new_n11055, new_n11056, new_n11057, new_n11058, new_n11059, new_n11060,
    new_n11061, new_n11062, new_n11063, new_n11064, new_n11065, new_n11066,
    new_n11067, new_n11068, new_n11069, new_n11070, new_n11071, new_n11072,
    new_n11073, new_n11074, new_n11075, new_n11076, new_n11077, new_n11078,
    new_n11079, new_n11080, new_n11081, new_n11082, new_n11083, new_n11084,
    new_n11085, new_n11086, new_n11087, new_n11088, new_n11089, new_n11090,
    new_n11091, new_n11092, new_n11093, new_n11094, new_n11095, new_n11096,
    new_n11097, new_n11098, new_n11099, new_n11100, new_n11101, new_n11102,
    new_n11103, new_n11104, new_n11105, new_n11106, new_n11107, new_n11108,
    new_n11109, new_n11110, new_n11111, new_n11112, new_n11113, new_n11114,
    new_n11115, new_n11116, new_n11117, new_n11118, new_n11119, new_n11120,
    new_n11121, new_n11122, new_n11123, new_n11124, new_n11125, new_n11126,
    new_n11127, new_n11128, new_n11129, new_n11130, new_n11131, new_n11132,
    new_n11133, new_n11134, new_n11135, new_n11136, new_n11137, new_n11138,
    new_n11139, new_n11140, new_n11141, new_n11142, new_n11143, new_n11144,
    new_n11145, new_n11146, new_n11147, new_n11148, new_n11149, new_n11150,
    new_n11151, new_n11152, new_n11153, new_n11154, new_n11155, new_n11156,
    new_n11157, new_n11158, new_n11159, new_n11160, new_n11161, new_n11162,
    new_n11163, new_n11164, new_n11165, new_n11166, new_n11167, new_n11168,
    new_n11169, new_n11170, new_n11171, new_n11172, new_n11173, new_n11174,
    new_n11175, new_n11176, new_n11177, new_n11178, new_n11179, new_n11180,
    new_n11181, new_n11182, new_n11183, new_n11184, new_n11185, new_n11186,
    new_n11187, new_n11188, new_n11189, new_n11190, new_n11191, new_n11192,
    new_n11193, new_n11194, new_n11195, new_n11196, new_n11197, new_n11198,
    new_n11199, new_n11200, new_n11201, new_n11202, new_n11203, new_n11204,
    new_n11205, new_n11206, new_n11207, new_n11208, new_n11209, new_n11210,
    new_n11211, new_n11212, new_n11213, new_n11214, new_n11215, new_n11216,
    new_n11217, new_n11218, new_n11219, new_n11220, new_n11221, new_n11222,
    new_n11223, new_n11224, new_n11225, new_n11226, new_n11227, new_n11228,
    new_n11229, new_n11230, new_n11231, new_n11232, new_n11233, new_n11234,
    new_n11235, new_n11236, new_n11237, new_n11238, new_n11239, new_n11240,
    new_n11241, new_n11242, new_n11243, new_n11244, new_n11245, new_n11246,
    new_n11247, new_n11248, new_n11249, new_n11250, new_n11251, new_n11252,
    new_n11253, new_n11254, new_n11255, new_n11256, new_n11257, new_n11258,
    new_n11259, new_n11260, new_n11261, new_n11262, new_n11263, new_n11264,
    new_n11265, new_n11266, new_n11267, new_n11268, new_n11269, new_n11270,
    new_n11271, new_n11272, new_n11273, new_n11274, new_n11275, new_n11276,
    new_n11277, new_n11278, new_n11279, new_n11280, new_n11281, new_n11282,
    new_n11283, new_n11284, new_n11285, new_n11286, new_n11287, new_n11288,
    new_n11289, new_n11290, new_n11291, new_n11292, new_n11293, new_n11294,
    new_n11295, new_n11296, new_n11297, new_n11298, new_n11299, new_n11300,
    new_n11301, new_n11302, new_n11303, new_n11304, new_n11305, new_n11306,
    new_n11307, new_n11308, new_n11309, new_n11310, new_n11311, new_n11312,
    new_n11313, new_n11314, new_n11315, new_n11316, new_n11317, new_n11318,
    new_n11319, new_n11320, new_n11321, new_n11322, new_n11323, new_n11324,
    new_n11325, new_n11326, new_n11327, new_n11328, new_n11329, new_n11330,
    new_n11331, new_n11332, new_n11333, new_n11334, new_n11335, new_n11336,
    new_n11337, new_n11338, new_n11339, new_n11340, new_n11341, new_n11342,
    new_n11343, new_n11344, new_n11345, new_n11346, new_n11347, new_n11348,
    new_n11349, new_n11350, new_n11351, new_n11352, new_n11353, new_n11354,
    new_n11355, new_n11356, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375, new_n11376, new_n11377, new_n11378,
    new_n11379, new_n11380, new_n11381, new_n11382, new_n11383, new_n11384,
    new_n11385, new_n11386, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391, new_n11392, new_n11393, new_n11394, new_n11395, new_n11396,
    new_n11397, new_n11398, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403, new_n11404, new_n11405, new_n11406, new_n11407, new_n11408,
    new_n11409, new_n11410, new_n11411, new_n11412, new_n11413, new_n11414,
    new_n11415, new_n11416, new_n11417, new_n11418, new_n11419, new_n11420,
    new_n11421, new_n11422, new_n11423, new_n11424, new_n11425, new_n11426,
    new_n11427, new_n11428, new_n11429, new_n11430, new_n11431, new_n11432,
    new_n11433, new_n11434, new_n11435, new_n11436, new_n11437, new_n11438,
    new_n11439, new_n11440, new_n11441, new_n11442, new_n11443, new_n11444,
    new_n11445, new_n11446, new_n11447, new_n11448, new_n11449, new_n11450,
    new_n11451, new_n11452, new_n11453, new_n11454, new_n11455, new_n11456,
    new_n11457, new_n11458, new_n11459, new_n11460, new_n11461, new_n11462,
    new_n11463, new_n11464, new_n11465, new_n11466, new_n11467, new_n11468,
    new_n11469, new_n11470, new_n11471, new_n11472, new_n11473, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478, new_n11479, new_n11480,
    new_n11481, new_n11482, new_n11483, new_n11484, new_n11485, new_n11486,
    new_n11487, new_n11488, new_n11489, new_n11490, new_n11491, new_n11492,
    new_n11493, new_n11494, new_n11495, new_n11496, new_n11497, new_n11498,
    new_n11499, new_n11500, new_n11501, new_n11502, new_n11503, new_n11504,
    new_n11505, new_n11506, new_n11507, new_n11508, new_n11509, new_n11510,
    new_n11511, new_n11512, new_n11513, new_n11514, new_n11515, new_n11516,
    new_n11517, new_n11518, new_n11519, new_n11520, new_n11521, new_n11522,
    new_n11523, new_n11524, new_n11525, new_n11526, new_n11527, new_n11528,
    new_n11529, new_n11530, new_n11531, new_n11532, new_n11533, new_n11534,
    new_n11535, new_n11536, new_n11537, new_n11538, new_n11539, new_n11540,
    new_n11541, new_n11542, new_n11543, new_n11544, new_n11545, new_n11546,
    new_n11547, new_n11548, new_n11549, new_n11550, new_n11551, new_n11552,
    new_n11553, new_n11554, new_n11555, new_n11556, new_n11557, new_n11558,
    new_n11559, new_n11560, new_n11561, new_n11562, new_n11563, new_n11564,
    new_n11565, new_n11566, new_n11567, new_n11568, new_n11569, new_n11570,
    new_n11571, new_n11572, new_n11573, new_n11574, new_n11575, new_n11576,
    new_n11577, new_n11578, new_n11579, new_n11580, new_n11581, new_n11582,
    new_n11583, new_n11584, new_n11585, new_n11586, new_n11587, new_n11588,
    new_n11589, new_n11590, new_n11591, new_n11592, new_n11593, new_n11594,
    new_n11595, new_n11596, new_n11597, new_n11598, new_n11599, new_n11600,
    new_n11601, new_n11602, new_n11603, new_n11604, new_n11605, new_n11606,
    new_n11607, new_n11608, new_n11609, new_n11610, new_n11611, new_n11612,
    new_n11613, new_n11614, new_n11615, new_n11616, new_n11617, new_n11618,
    new_n11619, new_n11620, new_n11621, new_n11622, new_n11623, new_n11624,
    new_n11625, new_n11626, new_n11627, new_n11628, new_n11629, new_n11630,
    new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636,
    new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642,
    new_n11643, new_n11644, new_n11645, new_n11646, new_n11647, new_n11648,
    new_n11649, new_n11650, new_n11651, new_n11652, new_n11653, new_n11654,
    new_n11655, new_n11656, new_n11657, new_n11658, new_n11659, new_n11660,
    new_n11661, new_n11662, new_n11663, new_n11664, new_n11665, new_n11666,
    new_n11667, new_n11668, new_n11669, new_n11670, new_n11671, new_n11672,
    new_n11673, new_n11674, new_n11675, new_n11676, new_n11677, new_n11678,
    new_n11679, new_n11680, new_n11681, new_n11682, new_n11683, new_n11684,
    new_n11685, new_n11686, new_n11687, new_n11688, new_n11689, new_n11690,
    new_n11691, new_n11692, new_n11693, new_n11694, new_n11695, new_n11696,
    new_n11697, new_n11698, new_n11699, new_n11700, new_n11701, new_n11702,
    new_n11703, new_n11704, new_n11705, new_n11706, new_n11707, new_n11708,
    new_n11709, new_n11710, new_n11711, new_n11712, new_n11713, new_n11714,
    new_n11715, new_n11716, new_n11717, new_n11718, new_n11719, new_n11720,
    new_n11721, new_n11722, new_n11723, new_n11724, new_n11725, new_n11726,
    new_n11727, new_n11728, new_n11729, new_n11730, new_n11731, new_n11732,
    new_n11733, new_n11734, new_n11735, new_n11736, new_n11737, new_n11738,
    new_n11739, new_n11740, new_n11741, new_n11742, new_n11743, new_n11744,
    new_n11745, new_n11746, new_n11747, new_n11748, new_n11749, new_n11750,
    new_n11751, new_n11752, new_n11753, new_n11754, new_n11755, new_n11756,
    new_n11757, new_n11758, new_n11759, new_n11760, new_n11761, new_n11762,
    new_n11763, new_n11764, new_n11765, new_n11766, new_n11767, new_n11768,
    new_n11769, new_n11770, new_n11771, new_n11772, new_n11773, new_n11774,
    new_n11775, new_n11776, new_n11777, new_n11778, new_n11779, new_n11780,
    new_n11781, new_n11782, new_n11783, new_n11784, new_n11785, new_n11786,
    new_n11787, new_n11788, new_n11789, new_n11790, new_n11791, new_n11792,
    new_n11793, new_n11794, new_n11795, new_n11796, new_n11797, new_n11798,
    new_n11799, new_n11800, new_n11801, new_n11802, new_n11803, new_n11804,
    new_n11805, new_n11806, new_n11807, new_n11808, new_n11809, new_n11810,
    new_n11811, new_n11812, new_n11813, new_n11814, new_n11815, new_n11816,
    new_n11817, new_n11818, new_n11819, new_n11820, new_n11821, new_n11822,
    new_n11823, new_n11824, new_n11825, new_n11826, new_n11827, new_n11828,
    new_n11829, new_n11830, new_n11831, new_n11832, new_n11833, new_n11834,
    new_n11835, new_n11836, new_n11837, new_n11838, new_n11839, new_n11840,
    new_n11841, new_n11842, new_n11843, new_n11844, new_n11845, new_n11846,
    new_n11847, new_n11848, new_n11849, new_n11850, new_n11851, new_n11852,
    new_n11853, new_n11854, new_n11855, new_n11856, new_n11857, new_n11858,
    new_n11859, new_n11860, new_n11861, new_n11862, new_n11863, new_n11864,
    new_n11865, new_n11866, new_n11867, new_n11868, new_n11869, new_n11870,
    new_n11871, new_n11872, new_n11873, new_n11874, new_n11875, new_n11876,
    new_n11877, new_n11878, new_n11879, new_n11880, new_n11881, new_n11882,
    new_n11883, new_n11884, new_n11885, new_n11886, new_n11887, new_n11888,
    new_n11889, new_n11890, new_n11891, new_n11892, new_n11893, new_n11894,
    new_n11895, new_n11896, new_n11897, new_n11898, new_n11899, new_n11900,
    new_n11901, new_n11902, new_n11903, new_n11904, new_n11905, new_n11906,
    new_n11907, new_n11908, new_n11909, new_n11910, new_n11911, new_n11912,
    new_n11913, new_n11914, new_n11915, new_n11916, new_n11917, new_n11918,
    new_n11919, new_n11920, new_n11921, new_n11922, new_n11923, new_n11924,
    new_n11925, new_n11926, new_n11927, new_n11928, new_n11929, new_n11930,
    new_n11931, new_n11932, new_n11933, new_n11934, new_n11935, new_n11936,
    new_n11937, new_n11938, new_n11939, new_n11940, new_n11941, new_n11942,
    new_n11943, new_n11944, new_n11945, new_n11946, new_n11947, new_n11948,
    new_n11949, new_n11950, new_n11951, new_n11952, new_n11953, new_n11954,
    new_n11955, new_n11956, new_n11957, new_n11958, new_n11959, new_n11960,
    new_n11961, new_n11962, new_n11963, new_n11964, new_n11965, new_n11966,
    new_n11967, new_n11968, new_n11969, new_n11970, new_n11971, new_n11972,
    new_n11973, new_n11974, new_n11975, new_n11976, new_n11977, new_n11978,
    new_n11979, new_n11980, new_n11981, new_n11982, new_n11983, new_n11984,
    new_n11985, new_n11986, new_n11987, new_n11988, new_n11989, new_n11990,
    new_n11991, new_n11992, new_n11993, new_n11994, new_n11995, new_n11996,
    new_n11997, new_n11998, new_n11999, new_n12000, new_n12001, new_n12002,
    new_n12003, new_n12004, new_n12005, new_n12006, new_n12007, new_n12008,
    new_n12009, new_n12010, new_n12011, new_n12012, new_n12013, new_n12014,
    new_n12015, new_n12016, new_n12017, new_n12018, new_n12019, new_n12020,
    new_n12021, new_n12022, new_n12023, new_n12024, new_n12025, new_n12026,
    new_n12027, new_n12028, new_n12029, new_n12030, new_n12031, new_n12032,
    new_n12033, new_n12034, new_n12035, new_n12036, new_n12037, new_n12038,
    new_n12039, new_n12040, new_n12041, new_n12042, new_n12043, new_n12044,
    new_n12045, new_n12046, new_n12047, new_n12048, new_n12049, new_n12050,
    new_n12051, new_n12052, new_n12053, new_n12054, new_n12055, new_n12056,
    new_n12057, new_n12058, new_n12059, new_n12060, new_n12061, new_n12062,
    new_n12063, new_n12064, new_n12065, new_n12066, new_n12067, new_n12068,
    new_n12069, new_n12070, new_n12071, new_n12072, new_n12073, new_n12074,
    new_n12075, new_n12076, new_n12077, new_n12078, new_n12079, new_n12080,
    new_n12081, new_n12082, new_n12083, new_n12084, new_n12085, new_n12086,
    new_n12087, new_n12088, new_n12089, new_n12090, new_n12091, new_n12092,
    new_n12093, new_n12094, new_n12095, new_n12096, new_n12097, new_n12098,
    new_n12099, new_n12100, new_n12101, new_n12102, new_n12103, new_n12104,
    new_n12105, new_n12106, new_n12107, new_n12108, new_n12109, new_n12110,
    new_n12111, new_n12112, new_n12113, new_n12114, new_n12115, new_n12116,
    new_n12117, new_n12118, new_n12119, new_n12120, new_n12121, new_n12122,
    new_n12123, new_n12124, new_n12125, new_n12126, new_n12127, new_n12128,
    new_n12129, new_n12130, new_n12131, new_n12132, new_n12133, new_n12134,
    new_n12135, new_n12136, new_n12137, new_n12138, new_n12139, new_n12140,
    new_n12141, new_n12142, new_n12143, new_n12144, new_n12145, new_n12146,
    new_n12147, new_n12148, new_n12149, new_n12150, new_n12151, new_n12152,
    new_n12153, new_n12154, new_n12155, new_n12156, new_n12157, new_n12158,
    new_n12159, new_n12160, new_n12161, new_n12162, new_n12163, new_n12164,
    new_n12165, new_n12166, new_n12167, new_n12168, new_n12169, new_n12170,
    new_n12171, new_n12172, new_n12173, new_n12174, new_n12175, new_n12176,
    new_n12177, new_n12178, new_n12179, new_n12180, new_n12181, new_n12182,
    new_n12183, new_n12184, new_n12185, new_n12186, new_n12187, new_n12188,
    new_n12189, new_n12190, new_n12191, new_n12192, new_n12193, new_n12194,
    new_n12195, new_n12196, new_n12197, new_n12198, new_n12199, new_n12200,
    new_n12201, new_n12202, new_n12203, new_n12204, new_n12205, new_n12206,
    new_n12207, new_n12208, new_n12209, new_n12210, new_n12211, new_n12212,
    new_n12213, new_n12214, new_n12215, new_n12216, new_n12217, new_n12218,
    new_n12219, new_n12220, new_n12221, new_n12222, new_n12223, new_n12224,
    new_n12225, new_n12226, new_n12227, new_n12228, new_n12229, new_n12230,
    new_n12231, new_n12232, new_n12233, new_n12234, new_n12235, new_n12236,
    new_n12237, new_n12238, new_n12239, new_n12240, new_n12241, new_n12242,
    new_n12243, new_n12244, new_n12245, new_n12246, new_n12247, new_n12248,
    new_n12249, new_n12250, new_n12251, new_n12252, new_n12253, new_n12254,
    new_n12255, new_n12256, new_n12257, new_n12258, new_n12259, new_n12260,
    new_n12261, new_n12262, new_n12263, new_n12264, new_n12265, new_n12266,
    new_n12267, new_n12268, new_n12269, new_n12270, new_n12271, new_n12272,
    new_n12273, new_n12274, new_n12275, new_n12276, new_n12277, new_n12278,
    new_n12279, new_n12280, new_n12281, new_n12282, new_n12283, new_n12284,
    new_n12285, new_n12286, new_n12287, new_n12288, new_n12289, new_n12290,
    new_n12291, new_n12292, new_n12293, new_n12294, new_n12295, new_n12296,
    new_n12297, new_n12298, new_n12299, new_n12300, new_n12301, new_n12302,
    new_n12303, new_n12304, new_n12305, new_n12306, new_n12307, new_n12308,
    new_n12309, new_n12310, new_n12311, new_n12312, new_n12313, new_n12314,
    new_n12315, new_n12316, new_n12317, new_n12318, new_n12319, new_n12320,
    new_n12321, new_n12322, new_n12323, new_n12324, new_n12325, new_n12326,
    new_n12327, new_n12328, new_n12329, new_n12330, new_n12331, new_n12332,
    new_n12333, new_n12334, new_n12335, new_n12336, new_n12337, new_n12338,
    new_n12339, new_n12340, new_n12341, new_n12342, new_n12343, new_n12344,
    new_n12345, new_n12346, new_n12347, new_n12348, new_n12349, new_n12350,
    new_n12351, new_n12352, new_n12353, new_n12354, new_n12355, new_n12356,
    new_n12357, new_n12358, new_n12359, new_n12360, new_n12361, new_n12362,
    new_n12363, new_n12364, new_n12365, new_n12366, new_n12367, new_n12368,
    new_n12369, new_n12370, new_n12371, new_n12372, new_n12373, new_n12374,
    new_n12375, new_n12376, new_n12377, new_n12378, new_n12379, new_n12380,
    new_n12381, new_n12382, new_n12383, new_n12384, new_n12385, new_n12386,
    new_n12387, new_n12388, new_n12389, new_n12390, new_n12391, new_n12392,
    new_n12393, new_n12394, new_n12395, new_n12396, new_n12397, new_n12398,
    new_n12399, new_n12400, new_n12401, new_n12402, new_n12403, new_n12404,
    new_n12405, new_n12406, new_n12407, new_n12408, new_n12409, new_n12410,
    new_n12411, new_n12412, new_n12413, new_n12414, new_n12415, new_n12416,
    new_n12417, new_n12418, new_n12419, new_n12420, new_n12421, new_n12422,
    new_n12423, new_n12424, new_n12425, new_n12426, new_n12427, new_n12428,
    new_n12429, new_n12430, new_n12431, new_n12432, new_n12433, new_n12434,
    new_n12435, new_n12436, new_n12437, new_n12438, new_n12439, new_n12440,
    new_n12441, new_n12442, new_n12443, new_n12444, new_n12445, new_n12446,
    new_n12447, new_n12448, new_n12449, new_n12450, new_n12451, new_n12452,
    new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458,
    new_n12459, new_n12460, new_n12461, new_n12462, new_n12463, new_n12464,
    new_n12465, new_n12466, new_n12467, new_n12468, new_n12469, new_n12470,
    new_n12471, new_n12472, new_n12473, new_n12474, new_n12475, new_n12476,
    new_n12477, new_n12478, new_n12479, new_n12480, new_n12481, new_n12482,
    new_n12483, new_n12484, new_n12485, new_n12486, new_n12487, new_n12488,
    new_n12489, new_n12490, new_n12491, new_n12492, new_n12493, new_n12494,
    new_n12495, new_n12496, new_n12497, new_n12498, new_n12499, new_n12500,
    new_n12501, new_n12502, new_n12503, new_n12504, new_n12505, new_n12506,
    new_n12507, new_n12508, new_n12509, new_n12510, new_n12511, new_n12512,
    new_n12513, new_n12514, new_n12515, new_n12516, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12531, new_n12532, new_n12533, new_n12534, new_n12535, new_n12536,
    new_n12537, new_n12538, new_n12539, new_n12540, new_n12541, new_n12542,
    new_n12543, new_n12544, new_n12545, new_n12546, new_n12547, new_n12548,
    new_n12549, new_n12550, new_n12551, new_n12552, new_n12553, new_n12554,
    new_n12555, new_n12556, new_n12557, new_n12558, new_n12559, new_n12560,
    new_n12561, new_n12562, new_n12563, new_n12564, new_n12565, new_n12566,
    new_n12567, new_n12568, new_n12569, new_n12570, new_n12571, new_n12572,
    new_n12573, new_n12574, new_n12575, new_n12576, new_n12577, new_n12578,
    new_n12579, new_n12580, new_n12581, new_n12582, new_n12583, new_n12584,
    new_n12585, new_n12586, new_n12587, new_n12588, new_n12589, new_n12590,
    new_n12591, new_n12592, new_n12593, new_n12594, new_n12595, new_n12596,
    new_n12597, new_n12598, new_n12599, new_n12600, new_n12601, new_n12602,
    new_n12603, new_n12604, new_n12605, new_n12606, new_n12607, new_n12608,
    new_n12609, new_n12610, new_n12611, new_n12612, new_n12613, new_n12614,
    new_n12615, new_n12616, new_n12617, new_n12618, new_n12619, new_n12620,
    new_n12621, new_n12622, new_n12623, new_n12624, new_n12625, new_n12626,
    new_n12627, new_n12628, new_n12629, new_n12630, new_n12631, new_n12632,
    new_n12633, new_n12634, new_n12635, new_n12636, new_n12637, new_n12638,
    new_n12639, new_n12640, new_n12641, new_n12642, new_n12643, new_n12644,
    new_n12645, new_n12646, new_n12647, new_n12648, new_n12649, new_n12650,
    new_n12651, new_n12652, new_n12653, new_n12654, new_n12655, new_n12656,
    new_n12657, new_n12658, new_n12659, new_n12660, new_n12661, new_n12662,
    new_n12663, new_n12664, new_n12665, new_n12666, new_n12667, new_n12668,
    new_n12669, new_n12670, new_n12671, new_n12672, new_n12673, new_n12674,
    new_n12675, new_n12676, new_n12677, new_n12678, new_n12679, new_n12680,
    new_n12681, new_n12682, new_n12683, new_n12684, new_n12685, new_n12686,
    new_n12687, new_n12688, new_n12689, new_n12690, new_n12691, new_n12692,
    new_n12693, new_n12694, new_n12695, new_n12696, new_n12697, new_n12698,
    new_n12699, new_n12700, new_n12701, new_n12702, new_n12703, new_n12704,
    new_n12705, new_n12706, new_n12707, new_n12708, new_n12709, new_n12710,
    new_n12711, new_n12712, new_n12713, new_n12714, new_n12715, new_n12716,
    new_n12717, new_n12718, new_n12719, new_n12720, new_n12721, new_n12722,
    new_n12723, new_n12724, new_n12725, new_n12726, new_n12727, new_n12728,
    new_n12729, new_n12730, new_n12731, new_n12732, new_n12733, new_n12734,
    new_n12735, new_n12736, new_n12737, new_n12738, new_n12739, new_n12740,
    new_n12741, new_n12742, new_n12743, new_n12744, new_n12745, new_n12746,
    new_n12747, new_n12748, new_n12749, new_n12750, new_n12751, new_n12752,
    new_n12753, new_n12754, new_n12755, new_n12756, new_n12757, new_n12758,
    new_n12759, new_n12760, new_n12761, new_n12762, new_n12763, new_n12764,
    new_n12765, new_n12766, new_n12767, new_n12768, new_n12769, new_n12770,
    new_n12771, new_n12772, new_n12773, new_n12774, new_n12775, new_n12776,
    new_n12777, new_n12778, new_n12779, new_n12780, new_n12781, new_n12782,
    new_n12783, new_n12784, new_n12785, new_n12786, new_n12787, new_n12788,
    new_n12789, new_n12790, new_n12791, new_n12792, new_n12793, new_n12794,
    new_n12795, new_n12796, new_n12797, new_n12798, new_n12799, new_n12800,
    new_n12801, new_n12802, new_n12803, new_n12804, new_n12805, new_n12806,
    new_n12807, new_n12808, new_n12809, new_n12810, new_n12811, new_n12812,
    new_n12813, new_n12814, new_n12815, new_n12816, new_n12817, new_n12818,
    new_n12819, new_n12820, new_n12821, new_n12822, new_n12823, new_n12824,
    new_n12825, new_n12826, new_n12827, new_n12828, new_n12829, new_n12830,
    new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836,
    new_n12837, new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843, new_n12844, new_n12845, new_n12846, new_n12847, new_n12848,
    new_n12849, new_n12850, new_n12851, new_n12852, new_n12853, new_n12854,
    new_n12855, new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861, new_n12862, new_n12863, new_n12864, new_n12865, new_n12866,
    new_n12867, new_n12868, new_n12869, new_n12870, new_n12871, new_n12872,
    new_n12873, new_n12874, new_n12875, new_n12876, new_n12877, new_n12878,
    new_n12879, new_n12880, new_n12881, new_n12882, new_n12883, new_n12884,
    new_n12885, new_n12886, new_n12887, new_n12888, new_n12889, new_n12890,
    new_n12891, new_n12892, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900, new_n12901, new_n12902,
    new_n12903, new_n12904, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917, new_n12918, new_n12919, new_n12920,
    new_n12921, new_n12922, new_n12923, new_n12924, new_n12925, new_n12926,
    new_n12927, new_n12928, new_n12929, new_n12930, new_n12931, new_n12932,
    new_n12933, new_n12934, new_n12935, new_n12936, new_n12937, new_n12938,
    new_n12939, new_n12940, new_n12941, new_n12942, new_n12943, new_n12944,
    new_n12945, new_n12946, new_n12947, new_n12948, new_n12949, new_n12950,
    new_n12951, new_n12952, new_n12953, new_n12954, new_n12955, new_n12956,
    new_n12957, new_n12958, new_n12959, new_n12960, new_n12961, new_n12962,
    new_n12963, new_n12964, new_n12965, new_n12966, new_n12967, new_n12968,
    new_n12969, new_n12970, new_n12971, new_n12972, new_n12973, new_n12974,
    new_n12975, new_n12976, new_n12977, new_n12978, new_n12979, new_n12980,
    new_n12981, new_n12982, new_n12983, new_n12984, new_n12985, new_n12986,
    new_n12987, new_n12988, new_n12989, new_n12990, new_n12991, new_n12992,
    new_n12993, new_n12994, new_n12995, new_n12996, new_n12997, new_n12998,
    new_n12999, new_n13000, new_n13001, new_n13002, new_n13003, new_n13004,
    new_n13005, new_n13006, new_n13007, new_n13008, new_n13009, new_n13010,
    new_n13011, new_n13012, new_n13013, new_n13014, new_n13015, new_n13016,
    new_n13017, new_n13018, new_n13019, new_n13020, new_n13021, new_n13022,
    new_n13023, new_n13024, new_n13025, new_n13026, new_n13027, new_n13028,
    new_n13029, new_n13030, new_n13031, new_n13032, new_n13033, new_n13034,
    new_n13035, new_n13036, new_n13037, new_n13038, new_n13039, new_n13040,
    new_n13041, new_n13042, new_n13043, new_n13044, new_n13045, new_n13046,
    new_n13047, new_n13048, new_n13049, new_n13050, new_n13051, new_n13052,
    new_n13053, new_n13054, new_n13055, new_n13056, new_n13057, new_n13058,
    new_n13059, new_n13060, new_n13061, new_n13062, new_n13063, new_n13064,
    new_n13065, new_n13066, new_n13067, new_n13068, new_n13069, new_n13070,
    new_n13071, new_n13072, new_n13073, new_n13074, new_n13075, new_n13076,
    new_n13077, new_n13078, new_n13079, new_n13080, new_n13081, new_n13082,
    new_n13083, new_n13084, new_n13085, new_n13086, new_n13087, new_n13088,
    new_n13089, new_n13090, new_n13091, new_n13092, new_n13093, new_n13094,
    new_n13095, new_n13096, new_n13097, new_n13098, new_n13099, new_n13100,
    new_n13101, new_n13102, new_n13103, new_n13104, new_n13105, new_n13106,
    new_n13107, new_n13108, new_n13109, new_n13110, new_n13111, new_n13112,
    new_n13113, new_n13114, new_n13115, new_n13116, new_n13117, new_n13118,
    new_n13119, new_n13120, new_n13121, new_n13122, new_n13123, new_n13124,
    new_n13125, new_n13126, new_n13127, new_n13128, new_n13129, new_n13130,
    new_n13131, new_n13132, new_n13133, new_n13134, new_n13135, new_n13136,
    new_n13137, new_n13138, new_n13139, new_n13140, new_n13141, new_n13142,
    new_n13143, new_n13144, new_n13145, new_n13146, new_n13147, new_n13148,
    new_n13149, new_n13150, new_n13151, new_n13152, new_n13153, new_n13154,
    new_n13155, new_n13156, new_n13157, new_n13158, new_n13159, new_n13160,
    new_n13161, new_n13162, new_n13163, new_n13164, new_n13165, new_n13166,
    new_n13167, new_n13168, new_n13169, new_n13170, new_n13171, new_n13172,
    new_n13173, new_n13174, new_n13175, new_n13176, new_n13177, new_n13178,
    new_n13179, new_n13180, new_n13181, new_n13182, new_n13183, new_n13184,
    new_n13185, new_n13186, new_n13187, new_n13188, new_n13189, new_n13190,
    new_n13191, new_n13192, new_n13193, new_n13194, new_n13195, new_n13196,
    new_n13197, new_n13198, new_n13199, new_n13200, new_n13201, new_n13202,
    new_n13203, new_n13204, new_n13205, new_n13206, new_n13207, new_n13208,
    new_n13209, new_n13210, new_n13211, new_n13212, new_n13213, new_n13214,
    new_n13215, new_n13216, new_n13217, new_n13218, new_n13219, new_n13220,
    new_n13221, new_n13222, new_n13223, new_n13224, new_n13225, new_n13226,
    new_n13227, new_n13228, new_n13229, new_n13230, new_n13231, new_n13232,
    new_n13233, new_n13234, new_n13235, new_n13236, new_n13237, new_n13238,
    new_n13239, new_n13240, new_n13241, new_n13242, new_n13243, new_n13244,
    new_n13245, new_n13246, new_n13247, new_n13248, new_n13249, new_n13250,
    new_n13251, new_n13252, new_n13253, new_n13254, new_n13255, new_n13256,
    new_n13257, new_n13258, new_n13259, new_n13260, new_n13261, new_n13262,
    new_n13263, new_n13264, new_n13265, new_n13266, new_n13267, new_n13268,
    new_n13269, new_n13270, new_n13271, new_n13272, new_n13273, new_n13274,
    new_n13275, new_n13276, new_n13277, new_n13278, new_n13279, new_n13280,
    new_n13281, new_n13282, new_n13283, new_n13284, new_n13285, new_n13286,
    new_n13287, new_n13288, new_n13289, new_n13290, new_n13291, new_n13292,
    new_n13293, new_n13294, new_n13295, new_n13296, new_n13297, new_n13298,
    new_n13299, new_n13300, new_n13301, new_n13302, new_n13303, new_n13304,
    new_n13305, new_n13306, new_n13307, new_n13308, new_n13309, new_n13310,
    new_n13311, new_n13312, new_n13313, new_n13314, new_n13315, new_n13316,
    new_n13317, new_n13318, new_n13319, new_n13320, new_n13321, new_n13322,
    new_n13323, new_n13324, new_n13325, new_n13326, new_n13327, new_n13328,
    new_n13329, new_n13330, new_n13331, new_n13332, new_n13333, new_n13334,
    new_n13335, new_n13336, new_n13337, new_n13338, new_n13339, new_n13340,
    new_n13341, new_n13342, new_n13343, new_n13344, new_n13345, new_n13346,
    new_n13347, new_n13348, new_n13349, new_n13350, new_n13351, new_n13352,
    new_n13353, new_n13354, new_n13355, new_n13356, new_n13357, new_n13358,
    new_n13359, new_n13360, new_n13361, new_n13362, new_n13363, new_n13364,
    new_n13365, new_n13366, new_n13367, new_n13368, new_n13369, new_n13370,
    new_n13371, new_n13372, new_n13373, new_n13374, new_n13375, new_n13376,
    new_n13377, new_n13378, new_n13379, new_n13380, new_n13381, new_n13382,
    new_n13383, new_n13384, new_n13385, new_n13386, new_n13387, new_n13388,
    new_n13389, new_n13390, new_n13391, new_n13392, new_n13393, new_n13394,
    new_n13395, new_n13396, new_n13397, new_n13398, new_n13399, new_n13400,
    new_n13401, new_n13402, new_n13403, new_n13404, new_n13405, new_n13406,
    new_n13407, new_n13408, new_n13409, new_n13410, new_n13411, new_n13412,
    new_n13413, new_n13414, new_n13415, new_n13416, new_n13417, new_n13418,
    new_n13419, new_n13420, new_n13421, new_n13422, new_n13423, new_n13424,
    new_n13425, new_n13426, new_n13427, new_n13428, new_n13429, new_n13430,
    new_n13431, new_n13432, new_n13433, new_n13434, new_n13435, new_n13436,
    new_n13437, new_n13438, new_n13439, new_n13440, new_n13441, new_n13442,
    new_n13443, new_n13444, new_n13445, new_n13446, new_n13447, new_n13448,
    new_n13449, new_n13450, new_n13451, new_n13452, new_n13453, new_n13454,
    new_n13455, new_n13456, new_n13457, new_n13458, new_n13459, new_n13460,
    new_n13461, new_n13462, new_n13463, new_n13464, new_n13465, new_n13466,
    new_n13467, new_n13468, new_n13469, new_n13470, new_n13471, new_n13472,
    new_n13473, new_n13474, new_n13475, new_n13476, new_n13477, new_n13478,
    new_n13479, new_n13480, new_n13481, new_n13482, new_n13483, new_n13484,
    new_n13485, new_n13486, new_n13487, new_n13488, new_n13489, new_n13490,
    new_n13491, new_n13492, new_n13493, new_n13494, new_n13495, new_n13496,
    new_n13497, new_n13498, new_n13499, new_n13500, new_n13501, new_n13502,
    new_n13503, new_n13504, new_n13505, new_n13506, new_n13507, new_n13508,
    new_n13509, new_n13510, new_n13511, new_n13512, new_n13513, new_n13514,
    new_n13515, new_n13516, new_n13517, new_n13518, new_n13519, new_n13520,
    new_n13521, new_n13522, new_n13523, new_n13524, new_n13525, new_n13526,
    new_n13527, new_n13528, new_n13529, new_n13530, new_n13531, new_n13532,
    new_n13533, new_n13534, new_n13535, new_n13536, new_n13537, new_n13538,
    new_n13539, new_n13540, new_n13541, new_n13542, new_n13543, new_n13544,
    new_n13545, new_n13546, new_n13547, new_n13548, new_n13549, new_n13550,
    new_n13551, new_n13552, new_n13553, new_n13554, new_n13555, new_n13556,
    new_n13557, new_n13558, new_n13559, new_n13560, new_n13561, new_n13562,
    new_n13563, new_n13564, new_n13565, new_n13566, new_n13567, new_n13568,
    new_n13569, new_n13570, new_n13571, new_n13572, new_n13573, new_n13574,
    new_n13575, new_n13576, new_n13577, new_n13578, new_n13579, new_n13580,
    new_n13581, new_n13582, new_n13583, new_n13584, new_n13585, new_n13586,
    new_n13587, new_n13588, new_n13589, new_n13590, new_n13591, new_n13592,
    new_n13593, new_n13594, new_n13595, new_n13596, new_n13597, new_n13598,
    new_n13599, new_n13600, new_n13601, new_n13602, new_n13603, new_n13604,
    new_n13605, new_n13606, new_n13607, new_n13608, new_n13609, new_n13610,
    new_n13611, new_n13612, new_n13613, new_n13614, new_n13615, new_n13616,
    new_n13617, new_n13618, new_n13619, new_n13620, new_n13621, new_n13622,
    new_n13623, new_n13624, new_n13625, new_n13626, new_n13627, new_n13628,
    new_n13629, new_n13630, new_n13631, new_n13632, new_n13633, new_n13634,
    new_n13635, new_n13636, new_n13637, new_n13638, new_n13639, new_n13640,
    new_n13641, new_n13642, new_n13643, new_n13644, new_n13645, new_n13646,
    new_n13647, new_n13648, new_n13649, new_n13650, new_n13651, new_n13652,
    new_n13653, new_n13654, new_n13655, new_n13656, new_n13657, new_n13658,
    new_n13659, new_n13660, new_n13661, new_n13662, new_n13663, new_n13664,
    new_n13665, new_n13666, new_n13667, new_n13668, new_n13669, new_n13670,
    new_n13671, new_n13672, new_n13673, new_n13674, new_n13675, new_n13676,
    new_n13677, new_n13678, new_n13679, new_n13680, new_n13681, new_n13682,
    new_n13683, new_n13684, new_n13685, new_n13686, new_n13687, new_n13688,
    new_n13689, new_n13690, new_n13691, new_n13692, new_n13693, new_n13694,
    new_n13695, new_n13696, new_n13697, new_n13698, new_n13699, new_n13700,
    new_n13701, new_n13702, new_n13703, new_n13704, new_n13705, new_n13706,
    new_n13707, new_n13708, new_n13709, new_n13710, new_n13711, new_n13712,
    new_n13713, new_n13714, new_n13715, new_n13716, new_n13717, new_n13718,
    new_n13719, new_n13720, new_n13721, new_n13722, new_n13723, new_n13724,
    new_n13725, new_n13726, new_n13727, new_n13728, new_n13729, new_n13730,
    new_n13731, new_n13732, new_n13733, new_n13734, new_n13735, new_n13736,
    new_n13737, new_n13738, new_n13739, new_n13740, new_n13741, new_n13742,
    new_n13743, new_n13744, new_n13745, new_n13746, new_n13747, new_n13748,
    new_n13749, new_n13750, new_n13751, new_n13752, new_n13753, new_n13754,
    new_n13755, new_n13756, new_n13757, new_n13758, new_n13759, new_n13760,
    new_n13761, new_n13762, new_n13763, new_n13764, new_n13765, new_n13766,
    new_n13767, new_n13768, new_n13769, new_n13770, new_n13771, new_n13772,
    new_n13773, new_n13774, new_n13775, new_n13776, new_n13777, new_n13778,
    new_n13779, new_n13780, new_n13781, new_n13782, new_n13783, new_n13784,
    new_n13785, new_n13786, new_n13787, new_n13788, new_n13789, new_n13790,
    new_n13791, new_n13792, new_n13793, new_n13794, new_n13795, new_n13796,
    new_n13797, new_n13798, new_n13799, new_n13800, new_n13801, new_n13802,
    new_n13803, new_n13804, new_n13805, new_n13806, new_n13807, new_n13808,
    new_n13809, new_n13810, new_n13811, new_n13812, new_n13813, new_n13814,
    new_n13815, new_n13816, new_n13817, new_n13818, new_n13819, new_n13820,
    new_n13821, new_n13822, new_n13823, new_n13824, new_n13825, new_n13826,
    new_n13827, new_n13828, new_n13829, new_n13830, new_n13831, new_n13832,
    new_n13833, new_n13834, new_n13835, new_n13836, new_n13837, new_n13838,
    new_n13839, new_n13840, new_n13841, new_n13842, new_n13843, new_n13844,
    new_n13845, new_n13846, new_n13847, new_n13848, new_n13849, new_n13850,
    new_n13851, new_n13852, new_n13853, new_n13854, new_n13855, new_n13856,
    new_n13857, new_n13858, new_n13859, new_n13860, new_n13861, new_n13862,
    new_n13863, new_n13864, new_n13865, new_n13866, new_n13867, new_n13868,
    new_n13869, new_n13870, new_n13871, new_n13872, new_n13873, new_n13874,
    new_n13875, new_n13876, new_n13877, new_n13878, new_n13879, new_n13880,
    new_n13881, new_n13882, new_n13883, new_n13884, new_n13885, new_n13886,
    new_n13887, new_n13888, new_n13889, new_n13890, new_n13891, new_n13892,
    new_n13893, new_n13894, new_n13895, new_n13896, new_n13897, new_n13898,
    new_n13899, new_n13900, new_n13901, new_n13902, new_n13903, new_n13904,
    new_n13905, new_n13906, new_n13907, new_n13908, new_n13909, new_n13910,
    new_n13911, new_n13912, new_n13913, new_n13914, new_n13915, new_n13916,
    new_n13917, new_n13918, new_n13919, new_n13920, new_n13921, new_n13922,
    new_n13923, new_n13924, new_n13925, new_n13926, new_n13927, new_n13928,
    new_n13929, new_n13930, new_n13931, new_n13932, new_n13933, new_n13934,
    new_n13935, new_n13936, new_n13937, new_n13938, new_n13939, new_n13940,
    new_n13941, new_n13942, new_n13943, new_n13944, new_n13945, new_n13946,
    new_n13947, new_n13948, new_n13949, new_n13950, new_n13951, new_n13952,
    new_n13953, new_n13954, new_n13955, new_n13956, new_n13957, new_n13958,
    new_n13959, new_n13960, new_n13961, new_n13962, new_n13963, new_n13964,
    new_n13965, new_n13966, new_n13967, new_n13968, new_n13969, new_n13970,
    new_n13971, new_n13972, new_n13973, new_n13974, new_n13975, new_n13976,
    new_n13977, new_n13978, new_n13979, new_n13980, new_n13981, new_n13982,
    new_n13983, new_n13984, new_n13985, new_n13986, new_n13987, new_n13988,
    new_n13989, new_n13990, new_n13991, new_n13992, new_n13993, new_n13994,
    new_n13995, new_n13996, new_n13997, new_n13998, new_n13999, new_n14000,
    new_n14001, new_n14002, new_n14003, new_n14004, new_n14005, new_n14006,
    new_n14007, new_n14008, new_n14009, new_n14010, new_n14011, new_n14012,
    new_n14013, new_n14014, new_n14015, new_n14016, new_n14017, new_n14018,
    new_n14019, new_n14020, new_n14021, new_n14022, new_n14023, new_n14024,
    new_n14025, new_n14026, new_n14027, new_n14028, new_n14029, new_n14030,
    new_n14031, new_n14032, new_n14033, new_n14034, new_n14035, new_n14036,
    new_n14037, new_n14038, new_n14039, new_n14040, new_n14041, new_n14042,
    new_n14043, new_n14044, new_n14045, new_n14046, new_n14047, new_n14048,
    new_n14049, new_n14050, new_n14051, new_n14052, new_n14053, new_n14054,
    new_n14055, new_n14056, new_n14057, new_n14058, new_n14059, new_n14060,
    new_n14061, new_n14062, new_n14063, new_n14064, new_n14065, new_n14066,
    new_n14067, new_n14068, new_n14069, new_n14070, new_n14071, new_n14072,
    new_n14073, new_n14074, new_n14075, new_n14076, new_n14077, new_n14078,
    new_n14079, new_n14080, new_n14081, new_n14082, new_n14083, new_n14084,
    new_n14085, new_n14086, new_n14087, new_n14088, new_n14089, new_n14090,
    new_n14091, new_n14092, new_n14093, new_n14094, new_n14095, new_n14096,
    new_n14097, new_n14098, new_n14099, new_n14100, new_n14101, new_n14102,
    new_n14103, new_n14104, new_n14105, new_n14106, new_n14107, new_n14108,
    new_n14109, new_n14110, new_n14111, new_n14112, new_n14113, new_n14114,
    new_n14115, new_n14116, new_n14117, new_n14118, new_n14119, new_n14120,
    new_n14121, new_n14122, new_n14123, new_n14124, new_n14125, new_n14126,
    new_n14127, new_n14128, new_n14129, new_n14130, new_n14131, new_n14132,
    new_n14133, new_n14134, new_n14135, new_n14136, new_n14137, new_n14138,
    new_n14139, new_n14140, new_n14141, new_n14142, new_n14143, new_n14144,
    new_n14145, new_n14146, new_n14147, new_n14148, new_n14149, new_n14150,
    new_n14151, new_n14152, new_n14153, new_n14154, new_n14155, new_n14156,
    new_n14157, new_n14158, new_n14159, new_n14160, new_n14161, new_n14162,
    new_n14163, new_n14164, new_n14165, new_n14166, new_n14167, new_n14168,
    new_n14169, new_n14170, new_n14171, new_n14172, new_n14173, new_n14174,
    new_n14175, new_n14176, new_n14177, new_n14178, new_n14179, new_n14180,
    new_n14181, new_n14182, new_n14183, new_n14184, new_n14185, new_n14186,
    new_n14187, new_n14188, new_n14189, new_n14190, new_n14191, new_n14192,
    new_n14193, new_n14194, new_n14195, new_n14196, new_n14197, new_n14198,
    new_n14199, new_n14200, new_n14201, new_n14202, new_n14203, new_n14204,
    new_n14205, new_n14206, new_n14207, new_n14208, new_n14209, new_n14210,
    new_n14211, new_n14212, new_n14213, new_n14214, new_n14215, new_n14216,
    new_n14217, new_n14218, new_n14219, new_n14220, new_n14221, new_n14222,
    new_n14223, new_n14224, new_n14225, new_n14226, new_n14227, new_n14228,
    new_n14229, new_n14230, new_n14231, new_n14232, new_n14233, new_n14234,
    new_n14235, new_n14236, new_n14237, new_n14238, new_n14239, new_n14240,
    new_n14241, new_n14242, new_n14243, new_n14244, new_n14245, new_n14246,
    new_n14247, new_n14248, new_n14249, new_n14250, new_n14251, new_n14252,
    new_n14253, new_n14254, new_n14255, new_n14256, new_n14257, new_n14258,
    new_n14259, new_n14260, new_n14261, new_n14262, new_n14263, new_n14264,
    new_n14265, new_n14266, new_n14267, new_n14268, new_n14269, new_n14270,
    new_n14271, new_n14272, new_n14273, new_n14274, new_n14275, new_n14276,
    new_n14277, new_n14278, new_n14279, new_n14280, new_n14281, new_n14282,
    new_n14283, new_n14284, new_n14285, new_n14286, new_n14287, new_n14288,
    new_n14289, new_n14290, new_n14291, new_n14292, new_n14293, new_n14294,
    new_n14295, new_n14296, new_n14297, new_n14298, new_n14299, new_n14300,
    new_n14301, new_n14302, new_n14303, new_n14304, new_n14305, new_n14306,
    new_n14307, new_n14308, new_n14309, new_n14310, new_n14311, new_n14312,
    new_n14313, new_n14314, new_n14315, new_n14316, new_n14317, new_n14318,
    new_n14319, new_n14320, new_n14321, new_n14322, new_n14323, new_n14324,
    new_n14325, new_n14326, new_n14327, new_n14328, new_n14329, new_n14330,
    new_n14331, new_n14332, new_n14333, new_n14334, new_n14335, new_n14336,
    new_n14337, new_n14338, new_n14339, new_n14340, new_n14341, new_n14342,
    new_n14343, new_n14344, new_n14345, new_n14346, new_n14347, new_n14348,
    new_n14349, new_n14350, new_n14351, new_n14352, new_n14353, new_n14354,
    new_n14355, new_n14356, new_n14357, new_n14358, new_n14359, new_n14360,
    new_n14361, new_n14362, new_n14363, new_n14364, new_n14365, new_n14366,
    new_n14367, new_n14368, new_n14369, new_n14370, new_n14371, new_n14372,
    new_n14373, new_n14374, new_n14375, new_n14376, new_n14377, new_n14378,
    new_n14379, new_n14380, new_n14381, new_n14382, new_n14383, new_n14384,
    new_n14385, new_n14386, new_n14387, new_n14388, new_n14389, new_n14390,
    new_n14391, new_n14392, new_n14393, new_n14394, new_n14395, new_n14396,
    new_n14397, new_n14398, new_n14399, new_n14400, new_n14401, new_n14402,
    new_n14403, new_n14404, new_n14405, new_n14406, new_n14407, new_n14408,
    new_n14409, new_n14410, new_n14411, new_n14412, new_n14413, new_n14414,
    new_n14415, new_n14416, new_n14417, new_n14418, new_n14419, new_n14420,
    new_n14421, new_n14422, new_n14423, new_n14424, new_n14425, new_n14426,
    new_n14427, new_n14428, new_n14429, new_n14430, new_n14431, new_n14432,
    new_n14433, new_n14434, new_n14435, new_n14436, new_n14437, new_n14438,
    new_n14439, new_n14440, new_n14441, new_n14442, new_n14443, new_n14444,
    new_n14445, new_n14446, new_n14447, new_n14448, new_n14449, new_n14450,
    new_n14451, new_n14452, new_n14453, new_n14454, new_n14455, new_n14456,
    new_n14457, new_n14458, new_n14459, new_n14460, new_n14461, new_n14462,
    new_n14463, new_n14464, new_n14465, new_n14466, new_n14467, new_n14468,
    new_n14469, new_n14470, new_n14471, new_n14472, new_n14473, new_n14474,
    new_n14475, new_n14476, new_n14477, new_n14478, new_n14479, new_n14480,
    new_n14481, new_n14482, new_n14483, new_n14484, new_n14485, new_n14486,
    new_n14487, new_n14488, new_n14489, new_n14490, new_n14491, new_n14492,
    new_n14493, new_n14494, new_n14495, new_n14496, new_n14497, new_n14498,
    new_n14499, new_n14500, new_n14501, new_n14502, new_n14503, new_n14504,
    new_n14505, new_n14506, new_n14507, new_n14508, new_n14509, new_n14510,
    new_n14511, new_n14512, new_n14513, new_n14514, new_n14515, new_n14516,
    new_n14517, new_n14518, new_n14519, new_n14520, new_n14521, new_n14522,
    new_n14523, new_n14524, new_n14525, new_n14526, new_n14527, new_n14528,
    new_n14529, new_n14530, new_n14531, new_n14532, new_n14533, new_n14534,
    new_n14535, new_n14536, new_n14537, new_n14538, new_n14539, new_n14540,
    new_n14541, new_n14542, new_n14543, new_n14544, new_n14545, new_n14546,
    new_n14547, new_n14548, new_n14549, new_n14550, new_n14551, new_n14552,
    new_n14553, new_n14554, new_n14555, new_n14556, new_n14557, new_n14558,
    new_n14559, new_n14560, new_n14561, new_n14562, new_n14563, new_n14564,
    new_n14565, new_n14566, new_n14567, new_n14568, new_n14569, new_n14570,
    new_n14571, new_n14572, new_n14573, new_n14574, new_n14575, new_n14576,
    new_n14577, new_n14578, new_n14579, new_n14580, new_n14581, new_n14582,
    new_n14583, new_n14584, new_n14585, new_n14586, new_n14587, new_n14588,
    new_n14589, new_n14590, new_n14591, new_n14592, new_n14593, new_n14594,
    new_n14595, new_n14596, new_n14597, new_n14598, new_n14599, new_n14600,
    new_n14601, new_n14602, new_n14603, new_n14604, new_n14605, new_n14606,
    new_n14607, new_n14608, new_n14609, new_n14610, new_n14611, new_n14612,
    new_n14613, new_n14614, new_n14615, new_n14616, new_n14617, new_n14618,
    new_n14619, new_n14620, new_n14621, new_n14622, new_n14623, new_n14624,
    new_n14625, new_n14626, new_n14627, new_n14628, new_n14629, new_n14630,
    new_n14631, new_n14632, new_n14633, new_n14634, new_n14635, new_n14636,
    new_n14637, new_n14638, new_n14639, new_n14640, new_n14641, new_n14642,
    new_n14643, new_n14644, new_n14645, new_n14646, new_n14647, new_n14648,
    new_n14649, new_n14650, new_n14651, new_n14652, new_n14653, new_n14654,
    new_n14655, new_n14656, new_n14657, new_n14658, new_n14659, new_n14660,
    new_n14661, new_n14662, new_n14663, new_n14664, new_n14665, new_n14666,
    new_n14667, new_n14668, new_n14669, new_n14670, new_n14671, new_n14672,
    new_n14673, new_n14674, new_n14675, new_n14676, new_n14677, new_n14678,
    new_n14679, new_n14680, new_n14681, new_n14682, new_n14683, new_n14684,
    new_n14685, new_n14686, new_n14687, new_n14688, new_n14689, new_n14690,
    new_n14691, new_n14692, new_n14693, new_n14694, new_n14695, new_n14696,
    new_n14697, new_n14698, new_n14699, new_n14700, new_n14701, new_n14702,
    new_n14703, new_n14704, new_n14705, new_n14706, new_n14707, new_n14708,
    new_n14709, new_n14710, new_n14711, new_n14712, new_n14713, new_n14714,
    new_n14715, new_n14716, new_n14717, new_n14718, new_n14719, new_n14720,
    new_n14721, new_n14722, new_n14723, new_n14724, new_n14725, new_n14726,
    new_n14727, new_n14728, new_n14729, new_n14730, new_n14731, new_n14732,
    new_n14733, new_n14734, new_n14735, new_n14736, new_n14737, new_n14738,
    new_n14739, new_n14740, new_n14741, new_n14742, new_n14743, new_n14744,
    new_n14745, new_n14746, new_n14747, new_n14748, new_n14749, new_n14750,
    new_n14751, new_n14752, new_n14753, new_n14754, new_n14755, new_n14756,
    new_n14757, new_n14758, new_n14759, new_n14760, new_n14761, new_n14762,
    new_n14763, new_n14764, new_n14765, new_n14766, new_n14767, new_n14768,
    new_n14769, new_n14770, new_n14771, new_n14772, new_n14773, new_n14774,
    new_n14775, new_n14776, new_n14777, new_n14778, new_n14779, new_n14780,
    new_n14781, new_n14782, new_n14783, new_n14784, new_n14785, new_n14786,
    new_n14787, new_n14788, new_n14789, new_n14790, new_n14791, new_n14792,
    new_n14793, new_n14794, new_n14795, new_n14796, new_n14797, new_n14798,
    new_n14799, new_n14800, new_n14801, new_n14802, new_n14803, new_n14804,
    new_n14805, new_n14806, new_n14807, new_n14808, new_n14809, new_n14810,
    new_n14811, new_n14812, new_n14813, new_n14814, new_n14815, new_n14816,
    new_n14817, new_n14818, new_n14819, new_n14820, new_n14821, new_n14822,
    new_n14823, new_n14824, new_n14825, new_n14826, new_n14827, new_n14828,
    new_n14829, new_n14830, new_n14831, new_n14832, new_n14833, new_n14834,
    new_n14835, new_n14836, new_n14837, new_n14838, new_n14839, new_n14840,
    new_n14841, new_n14842, new_n14843, new_n14844, new_n14845, new_n14846,
    new_n14847, new_n14848, new_n14849, new_n14850, new_n14851, new_n14852,
    new_n14853, new_n14854, new_n14855, new_n14856, new_n14857, new_n14858,
    new_n14859, new_n14860, new_n14861, new_n14862, new_n14863, new_n14864,
    new_n14865, new_n14866, new_n14867, new_n14868, new_n14869, new_n14870,
    new_n14871, new_n14872, new_n14873, new_n14874, new_n14875, new_n14876,
    new_n14877, new_n14878, new_n14879, new_n14880, new_n14881, new_n14882,
    new_n14883, new_n14884, new_n14885, new_n14886, new_n14887, new_n14888,
    new_n14889, new_n14890, new_n14891, new_n14892, new_n14893, new_n14894,
    new_n14895, new_n14896, new_n14897, new_n14898, new_n14899, new_n14900,
    new_n14901, new_n14902, new_n14903, new_n14904, new_n14905, new_n14906,
    new_n14907, new_n14908, new_n14909, new_n14910, new_n14911, new_n14912,
    new_n14913, new_n14914, new_n14915, new_n14916, new_n14917, new_n14918,
    new_n14919, new_n14920, new_n14921, new_n14922, new_n14923, new_n14924,
    new_n14925, new_n14926, new_n14927, new_n14928, new_n14929, new_n14930,
    new_n14931, new_n14932, new_n14933, new_n14934, new_n14935, new_n14936,
    new_n14937, new_n14938, new_n14939, new_n14940, new_n14941, new_n14942,
    new_n14943, new_n14944, new_n14945, new_n14946, new_n14947, new_n14948,
    new_n14949, new_n14950, new_n14951, new_n14952, new_n14953, new_n14954,
    new_n14955, new_n14956, new_n14957, new_n14958, new_n14959, new_n14960,
    new_n14961, new_n14962, new_n14963, new_n14964, new_n14965, new_n14966,
    new_n14967, new_n14968, new_n14969, new_n14970, new_n14971, new_n14972,
    new_n14973, new_n14974, new_n14975, new_n14976, new_n14977, new_n14978,
    new_n14979, new_n14980, new_n14981, new_n14982, new_n14983, new_n14984,
    new_n14985, new_n14986, new_n14987, new_n14988, new_n14989, new_n14990,
    new_n14991, new_n14992, new_n14993, new_n14994, new_n14995, new_n14996,
    new_n14997, new_n14998, new_n14999, new_n15000, new_n15001, new_n15002,
    new_n15003, new_n15004, new_n15005, new_n15006, new_n15007, new_n15008,
    new_n15009, new_n15010, new_n15011, new_n15012, new_n15013, new_n15014,
    new_n15015, new_n15016, new_n15017, new_n15018, new_n15019, new_n15020,
    new_n15021, new_n15022, new_n15023, new_n15024, new_n15025, new_n15026,
    new_n15027, new_n15028, new_n15029, new_n15030, new_n15031, new_n15032,
    new_n15033, new_n15034, new_n15035, new_n15036, new_n15037, new_n15038,
    new_n15039, new_n15040, new_n15041, new_n15042, new_n15043, new_n15044,
    new_n15045, new_n15046, new_n15047, new_n15048, new_n15049, new_n15050,
    new_n15051, new_n15052, new_n15053, new_n15054, new_n15055, new_n15056,
    new_n15057, new_n15058, new_n15059, new_n15060, new_n15061, new_n15062,
    new_n15063, new_n15064, new_n15065, new_n15066, new_n15067, new_n15068,
    new_n15069, new_n15070, new_n15071, new_n15072, new_n15073, new_n15074,
    new_n15075, new_n15076, new_n15077, new_n15078, new_n15079, new_n15080,
    new_n15081, new_n15082, new_n15083, new_n15084, new_n15085, new_n15086,
    new_n15087, new_n15088, new_n15089, new_n15090, new_n15091, new_n15092,
    new_n15093, new_n15094, new_n15095, new_n15096, new_n15097, new_n15098,
    new_n15099, new_n15100, new_n15101, new_n15102, new_n15103, new_n15104,
    new_n15105, new_n15106, new_n15107, new_n15108, new_n15109, new_n15110,
    new_n15111, new_n15112, new_n15113, new_n15114, new_n15115, new_n15116,
    new_n15117, new_n15118, new_n15119, new_n15120, new_n15121, new_n15122,
    new_n15123, new_n15124, new_n15125, new_n15126, new_n15127, new_n15128,
    new_n15129, new_n15130, new_n15131, new_n15132, new_n15133, new_n15134,
    new_n15135, new_n15136, new_n15137, new_n15138, new_n15139, new_n15140,
    new_n15141, new_n15142, new_n15143, new_n15144, new_n15145, new_n15146,
    new_n15147, new_n15148, new_n15149, new_n15150, new_n15151, new_n15152,
    new_n15153, new_n15154, new_n15155, new_n15156, new_n15157, new_n15158,
    new_n15159, new_n15160, new_n15161, new_n15162, new_n15163, new_n15164,
    new_n15165, new_n15166, new_n15167, new_n15168, new_n15169, new_n15170,
    new_n15171, new_n15172, new_n15173, new_n15174, new_n15175, new_n15176,
    new_n15177, new_n15178, new_n15179, new_n15180, new_n15181, new_n15182,
    new_n15183, new_n15184, new_n15185, new_n15186, new_n15187, new_n15188,
    new_n15189, new_n15190, new_n15191, new_n15192, new_n15193, new_n15194,
    new_n15195, new_n15196, new_n15197, new_n15198, new_n15199, new_n15200,
    new_n15201, new_n15202, new_n15203, new_n15204, new_n15205, new_n15206,
    new_n15207, new_n15208, new_n15209, new_n15210, new_n15211, new_n15212,
    new_n15213, new_n15214, new_n15215, new_n15216, new_n15217, new_n15218,
    new_n15219, new_n15220, new_n15221, new_n15222, new_n15223, new_n15224,
    new_n15225, new_n15226, new_n15227, new_n15228, new_n15229, new_n15230,
    new_n15231, new_n15232, new_n15233, new_n15234, new_n15235, new_n15236,
    new_n15237, new_n15238, new_n15239, new_n15240, new_n15241, new_n15242,
    new_n15243, new_n15244, new_n15245, new_n15246, new_n15247, new_n15248,
    new_n15249, new_n15250, new_n15251, new_n15252, new_n15253, new_n15254,
    new_n15255, new_n15256, new_n15257, new_n15258, new_n15259, new_n15260,
    new_n15261, new_n15262, new_n15263, new_n15264, new_n15265, new_n15266,
    new_n15267, new_n15268, new_n15269, new_n15270, new_n15271, new_n15272,
    new_n15273, new_n15274, new_n15275, new_n15276, new_n15277, new_n15278,
    new_n15279, new_n15280, new_n15281, new_n15282, new_n15283, new_n15284,
    new_n15285, new_n15286, new_n15287, new_n15288, new_n15289, new_n15290,
    new_n15291, new_n15292, new_n15293, new_n15294, new_n15295, new_n15296,
    new_n15297, new_n15298, new_n15299, new_n15300, new_n15301, new_n15302,
    new_n15303, new_n15304, new_n15305, new_n15306, new_n15307, new_n15308,
    new_n15309, new_n15310, new_n15311, new_n15312, new_n15313, new_n15314,
    new_n15315, new_n15316, new_n15317, new_n15318, new_n15319, new_n15320,
    new_n15321, new_n15322, new_n15323, new_n15324, new_n15325, new_n15326,
    new_n15327, new_n15328, new_n15329, new_n15330, new_n15331, new_n15332,
    new_n15333, new_n15334, new_n15335, new_n15336, new_n15337, new_n15338,
    new_n15339, new_n15340, new_n15341, new_n15342, new_n15343, new_n15344,
    new_n15345, new_n15346, new_n15347, new_n15348, new_n15349, new_n15350,
    new_n15351, new_n15352, new_n15353, new_n15354, new_n15355, new_n15356,
    new_n15357, new_n15358, new_n15359, new_n15360, new_n15361, new_n15362,
    new_n15363, new_n15364, new_n15365, new_n15366, new_n15367, new_n15368,
    new_n15369, new_n15370, new_n15371, new_n15372, new_n15373, new_n15374,
    new_n15375, new_n15376, new_n15377, new_n15378, new_n15379, new_n15380,
    new_n15381, new_n15382, new_n15383, new_n15384, new_n15385, new_n15386,
    new_n15387, new_n15388, new_n15389, new_n15390, new_n15391, new_n15392,
    new_n15393, new_n15394, new_n15395, new_n15396, new_n15397, new_n15398,
    new_n15399, new_n15400, new_n15401, new_n15402, new_n15403, new_n15404,
    new_n15405, new_n15406, new_n15407, new_n15408, new_n15409, new_n15410,
    new_n15411, new_n15412, new_n15413, new_n15414, new_n15415, new_n15416,
    new_n15417, new_n15418, new_n15419, new_n15420, new_n15421, new_n15422,
    new_n15423, new_n15424, new_n15425, new_n15426, new_n15427, new_n15428,
    new_n15429, new_n15430, new_n15431, new_n15432, new_n15433, new_n15434,
    new_n15435, new_n15436, new_n15437, new_n15438, new_n15439, new_n15440,
    new_n15441, new_n15442, new_n15443, new_n15444, new_n15445, new_n15446,
    new_n15447, new_n15448, new_n15449, new_n15450, new_n15451, new_n15452,
    new_n15453, new_n15454, new_n15455, new_n15456, new_n15457, new_n15458,
    new_n15459, new_n15460, new_n15461, new_n15462, new_n15463, new_n15464,
    new_n15465, new_n15466, new_n15467, new_n15468, new_n15469, new_n15470,
    new_n15471, new_n15472, new_n15473, new_n15474, new_n15475, new_n15476,
    new_n15477, new_n15478, new_n15479, new_n15480, new_n15481, new_n15482,
    new_n15483, new_n15484, new_n15485, new_n15486, new_n15487, new_n15488,
    new_n15489, new_n15490, new_n15491, new_n15492, new_n15493, new_n15494,
    new_n15495, new_n15496, new_n15497, new_n15498, new_n15499, new_n15500,
    new_n15501, new_n15502, new_n15503, new_n15504, new_n15505, new_n15506,
    new_n15507, new_n15508, new_n15509, new_n15510, new_n15511, new_n15512,
    new_n15513, new_n15514, new_n15515, new_n15516, new_n15517, new_n15518,
    new_n15519, new_n15520, new_n15521, new_n15522, new_n15523, new_n15524,
    new_n15525, new_n15526, new_n15527, new_n15528, new_n15529, new_n15530,
    new_n15531, new_n15532, new_n15533, new_n15534, new_n15535, new_n15536,
    new_n15537, new_n15538, new_n15539, new_n15540, new_n15541, new_n15542,
    new_n15543, new_n15544, new_n15545, new_n15546, new_n15547, new_n15548,
    new_n15549, new_n15550, new_n15551, new_n15552, new_n15553, new_n15554,
    new_n15555, new_n15556, new_n15557, new_n15558, new_n15559, new_n15560,
    new_n15561, new_n15562, new_n15563, new_n15564, new_n15565, new_n15566,
    new_n15567, new_n15568, new_n15569, new_n15570, new_n15571, new_n15572,
    new_n15573, new_n15574, new_n15575, new_n15576, new_n15577, new_n15578,
    new_n15579, new_n15580, new_n15581, new_n15582, new_n15583, new_n15584,
    new_n15585, new_n15586, new_n15587, new_n15588, new_n15589, new_n15590,
    new_n15591, new_n15592, new_n15593, new_n15594, new_n15595, new_n15596,
    new_n15597, new_n15598, new_n15599, new_n15600, new_n15601, new_n15602,
    new_n15603, new_n15604, new_n15605, new_n15606, new_n15607, new_n15608,
    new_n15609, new_n15610, new_n15611, new_n15612, new_n15613, new_n15614,
    new_n15615, new_n15616, new_n15617, new_n15618, new_n15619, new_n15620,
    new_n15621, new_n15622, new_n15623, new_n15624, new_n15625, new_n15626,
    new_n15627, new_n15628, new_n15629, new_n15630, new_n15631, new_n15632,
    new_n15633, new_n15634, new_n15635, new_n15636, new_n15637, new_n15638,
    new_n15639, new_n15640, new_n15641, new_n15642, new_n15643, new_n15644,
    new_n15645, new_n15646, new_n15647, new_n15648, new_n15649, new_n15650,
    new_n15651, new_n15652, new_n15653, new_n15654, new_n15655, new_n15656,
    new_n15657, new_n15658, new_n15659, new_n15660, new_n15661, new_n15662,
    new_n15663, new_n15664, new_n15665, new_n15666, new_n15667, new_n15668,
    new_n15669, new_n15670, new_n15671, new_n15672, new_n15673, new_n15674,
    new_n15675, new_n15676, new_n15677, new_n15678, new_n15679, new_n15680,
    new_n15681, new_n15682, new_n15683, new_n15684, new_n15685, new_n15686,
    new_n15687, new_n15688, new_n15689, new_n15690, new_n15691, new_n15692,
    new_n15693, new_n15694, new_n15695, new_n15696, new_n15697, new_n15698,
    new_n15699, new_n15700, new_n15701, new_n15702, new_n15703, new_n15704,
    new_n15705, new_n15706, new_n15707, new_n15708, new_n15709, new_n15710,
    new_n15711, new_n15712, new_n15713, new_n15714, new_n15715, new_n15716,
    new_n15717, new_n15718, new_n15719, new_n15720, new_n15721, new_n15722,
    new_n15723, new_n15724, new_n15725, new_n15726, new_n15727, new_n15728,
    new_n15729, new_n15730, new_n15731, new_n15732, new_n15733, new_n15734,
    new_n15735, new_n15736, new_n15737, new_n15738, new_n15739, new_n15740,
    new_n15741, new_n15742, new_n15743, new_n15744, new_n15745, new_n15746,
    new_n15747, new_n15748, new_n15749, new_n15750, new_n15751, new_n15752,
    new_n15753, new_n15754, new_n15755, new_n15756, new_n15757, new_n15758,
    new_n15759, new_n15760, new_n15761, new_n15762, new_n15763, new_n15764,
    new_n15765, new_n15766, new_n15767, new_n15768, new_n15769, new_n15770,
    new_n15771, new_n15772, new_n15773, new_n15774, new_n15775, new_n15776,
    new_n15777, new_n15778, new_n15779, new_n15780, new_n15781, new_n15782,
    new_n15783, new_n15784, new_n15785, new_n15786, new_n15787, new_n15788,
    new_n15789, new_n15790, new_n15791, new_n15792, new_n15793, new_n15794,
    new_n15795, new_n15796, new_n15797, new_n15798, new_n15799, new_n15800,
    new_n15801, new_n15802, new_n15803, new_n15804, new_n15805, new_n15806,
    new_n15807, new_n15808, new_n15809, new_n15810, new_n15811, new_n15812,
    new_n15813, new_n15814, new_n15815, new_n15816, new_n15817, new_n15818,
    new_n15819, new_n15820, new_n15821, new_n15822, new_n15823, new_n15824,
    new_n15825, new_n15826, new_n15827, new_n15828, new_n15829, new_n15830,
    new_n15831, new_n15832, new_n15833, new_n15834, new_n15835, new_n15836,
    new_n15837, new_n15838, new_n15839, new_n15840, new_n15841, new_n15842,
    new_n15843, new_n15844, new_n15845, new_n15846, new_n15847, new_n15848,
    new_n15849, new_n15850, new_n15851, new_n15852, new_n15853, new_n15854,
    new_n15855, new_n15856, new_n15857, new_n15858, new_n15859, new_n15860,
    new_n15861, new_n15862, new_n15863, new_n15864, new_n15865, new_n15866,
    new_n15867, new_n15868, new_n15869, new_n15870, new_n15871, new_n15872,
    new_n15873, new_n15874, new_n15875, new_n15876, new_n15877, new_n15878,
    new_n15879, new_n15880, new_n15881, new_n15882, new_n15883, new_n15884,
    new_n15885, new_n15886, new_n15887, new_n15888, new_n15889, new_n15890,
    new_n15891, new_n15892, new_n15893, new_n15894, new_n15895, new_n15896,
    new_n15897, new_n15898, new_n15899, new_n15900, new_n15901, new_n15902,
    new_n15903, new_n15904, new_n15905, new_n15906, new_n15907, new_n15908,
    new_n15909, new_n15910, new_n15911, new_n15912, new_n15913, new_n15914,
    new_n15915, new_n15916, new_n15917, new_n15918, new_n15919, new_n15920,
    new_n15921, new_n15922, new_n15923, new_n15924, new_n15925, new_n15926,
    new_n15927, new_n15928, new_n15929, new_n15930, new_n15931, new_n15932,
    new_n15933, new_n15934, new_n15935, new_n15936, new_n15937, new_n15938,
    new_n15939, new_n15940, new_n15941, new_n15942, new_n15943, new_n15944,
    new_n15945, new_n15946, new_n15947, new_n15948, new_n15949, new_n15950,
    new_n15951, new_n15952, new_n15953, new_n15954, new_n15955, new_n15956,
    new_n15957, new_n15958, new_n15959, new_n15960, new_n15961, new_n15962,
    new_n15963, new_n15964, new_n15965, new_n15966, new_n15967, new_n15968,
    new_n15969, new_n15970, new_n15971, new_n15972, new_n15973, new_n15974,
    new_n15975, new_n15976, new_n15977, new_n15978, new_n15979, new_n15980,
    new_n15981, new_n15982, new_n15983, new_n15984, new_n15985, new_n15986,
    new_n15987, new_n15988, new_n15989, new_n15990, new_n15991, new_n15992,
    new_n15993, new_n15994, new_n15995, new_n15996, new_n15997, new_n15998,
    new_n15999, new_n16000, new_n16001, new_n16002, new_n16003, new_n16004,
    new_n16005, new_n16006, new_n16007, new_n16008, new_n16009, new_n16010,
    new_n16011, new_n16012, new_n16013, new_n16014, new_n16015, new_n16016,
    new_n16017, new_n16018, new_n16019, new_n16020, new_n16021, new_n16022,
    new_n16023, new_n16024, new_n16025, new_n16026, new_n16027, new_n16028,
    new_n16029, new_n16030, new_n16031, new_n16032, new_n16033, new_n16034,
    new_n16035, new_n16036, new_n16037, new_n16038, new_n16039, new_n16040,
    new_n16041, new_n16042, new_n16043, new_n16044, new_n16045, new_n16046,
    new_n16047, new_n16048, new_n16049, new_n16050, new_n16051, new_n16052,
    new_n16053, new_n16054, new_n16055, new_n16056, new_n16057, new_n16058,
    new_n16059, new_n16060, new_n16061, new_n16062, new_n16063, new_n16064,
    new_n16065, new_n16066, new_n16067, new_n16068, new_n16069, new_n16070,
    new_n16071, new_n16072, new_n16073, new_n16074, new_n16075, new_n16076,
    new_n16077, new_n16078, new_n16079, new_n16080, new_n16081, new_n16082,
    new_n16083, new_n16084, new_n16085, new_n16086, new_n16087, new_n16088,
    new_n16089, new_n16090, new_n16091, new_n16092, new_n16093, new_n16094,
    new_n16095, new_n16096, new_n16097, new_n16098, new_n16099, new_n16100,
    new_n16101, new_n16102, new_n16103, new_n16104, new_n16105, new_n16106,
    new_n16107, new_n16108, new_n16109, new_n16110, new_n16111, new_n16112,
    new_n16113, new_n16114, new_n16115, new_n16116, new_n16117, new_n16118,
    new_n16119, new_n16120, new_n16121, new_n16122, new_n16123, new_n16124,
    new_n16125, new_n16126, new_n16127, new_n16128, new_n16129, new_n16130,
    new_n16131, new_n16132, new_n16133, new_n16134, new_n16135, new_n16136,
    new_n16137, new_n16138, new_n16139, new_n16140, new_n16141, new_n16142,
    new_n16143, new_n16144, new_n16145, new_n16146, new_n16147, new_n16148,
    new_n16149, new_n16150, new_n16151, new_n16152, new_n16153, new_n16154,
    new_n16155, new_n16156, new_n16157, new_n16158, new_n16159, new_n16160,
    new_n16161, new_n16162, new_n16163, new_n16164, new_n16165, new_n16166,
    new_n16167, new_n16168, new_n16169, new_n16170, new_n16171, new_n16172,
    new_n16173, new_n16174, new_n16175, new_n16176, new_n16177, new_n16178,
    new_n16179, new_n16180, new_n16181, new_n16182, new_n16183, new_n16184,
    new_n16185, new_n16186, new_n16187, new_n16188, new_n16189, new_n16190,
    new_n16191, new_n16192, new_n16193, new_n16194, new_n16195, new_n16196,
    new_n16197, new_n16198, new_n16199, new_n16200, new_n16201, new_n16202,
    new_n16203, new_n16204, new_n16205, new_n16206, new_n16207, new_n16208,
    new_n16209, new_n16210, new_n16211, new_n16212, new_n16213, new_n16214,
    new_n16215, new_n16216, new_n16217, new_n16218, new_n16219, new_n16220,
    new_n16221, new_n16222, new_n16223, new_n16224, new_n16225, new_n16226,
    new_n16227, new_n16228, new_n16229, new_n16230, new_n16231, new_n16232,
    new_n16233, new_n16234, new_n16235, new_n16236, new_n16237, new_n16238,
    new_n16239, new_n16240, new_n16241, new_n16242, new_n16243, new_n16244,
    new_n16245, new_n16246, new_n16247, new_n16248, new_n16249, new_n16250,
    new_n16251, new_n16252, new_n16253, new_n16254, new_n16255, new_n16256,
    new_n16257, new_n16258, new_n16259, new_n16260, new_n16261, new_n16262,
    new_n16263, new_n16264, new_n16265, new_n16266, new_n16267, new_n16268,
    new_n16269, new_n16270, new_n16271, new_n16272, new_n16273, new_n16274,
    new_n16275, new_n16276, new_n16277, new_n16278, new_n16279, new_n16280,
    new_n16281, new_n16282, new_n16283, new_n16284, new_n16285, new_n16286,
    new_n16287, new_n16288, new_n16289, new_n16290, new_n16291, new_n16292,
    new_n16293, new_n16294, new_n16295, new_n16296, new_n16297, new_n16298,
    new_n16299, new_n16300, new_n16301, new_n16302, new_n16303, new_n16304,
    new_n16305, new_n16306, new_n16307, new_n16308, new_n16309, new_n16310,
    new_n16311, new_n16312, new_n16313, new_n16314, new_n16315, new_n16316,
    new_n16317, new_n16318, new_n16319, new_n16320, new_n16321, new_n16322,
    new_n16323, new_n16324, new_n16325, new_n16326, new_n16327, new_n16328,
    new_n16329, new_n16330, new_n16331, new_n16332, new_n16333, new_n16334,
    new_n16335, new_n16336, new_n16337, new_n16338, new_n16339, new_n16340,
    new_n16341, new_n16342, new_n16343, new_n16344, new_n16345, new_n16346,
    new_n16347, new_n16348, new_n16349, new_n16350, new_n16351, new_n16352,
    new_n16353, new_n16354, new_n16355, new_n16356, new_n16357, new_n16358,
    new_n16359, new_n16360, new_n16361, new_n16362, new_n16363, new_n16364,
    new_n16365, new_n16366, new_n16367, new_n16368, new_n16369, new_n16370,
    new_n16371, new_n16372, new_n16373, new_n16374, new_n16375, new_n16376,
    new_n16377, new_n16378, new_n16379, new_n16380, new_n16381, new_n16382,
    new_n16383, new_n16384, new_n16385, new_n16386, new_n16387, new_n16388,
    new_n16389, new_n16390, new_n16391, new_n16392, new_n16393, new_n16394,
    new_n16395, new_n16396, new_n16397, new_n16398, new_n16399, new_n16400,
    new_n16401, new_n16402, new_n16403, new_n16404, new_n16405, new_n16406,
    new_n16407, new_n16408, new_n16409, new_n16410, new_n16411, new_n16412,
    new_n16413, new_n16414, new_n16415, new_n16416, new_n16417, new_n16418,
    new_n16419, new_n16420, new_n16421, new_n16422, new_n16423, new_n16424,
    new_n16425, new_n16426, new_n16427, new_n16428, new_n16429, new_n16430,
    new_n16431, new_n16432, new_n16433, new_n16434, new_n16435, new_n16436,
    new_n16437, new_n16438, new_n16439, new_n16440, new_n16441, new_n16442,
    new_n16443, new_n16444, new_n16445, new_n16446, new_n16447, new_n16448,
    new_n16449, new_n16450, new_n16451, new_n16452, new_n16453, new_n16454,
    new_n16455, new_n16456, new_n16457, new_n16458, new_n16459, new_n16460,
    new_n16461, new_n16462, new_n16463, new_n16464, new_n16465, new_n16466,
    new_n16467, new_n16468, new_n16469, new_n16470, new_n16471, new_n16472,
    new_n16473, new_n16474, new_n16475, new_n16476, new_n16477, new_n16478,
    new_n16479, new_n16480, new_n16481, new_n16482, new_n16483, new_n16484,
    new_n16485, new_n16486, new_n16487, new_n16488, new_n16489, new_n16490,
    new_n16491, new_n16492, new_n16493, new_n16494, new_n16495, new_n16496,
    new_n16497, new_n16498, new_n16499, new_n16500, new_n16501, new_n16502,
    new_n16503, new_n16504, new_n16505, new_n16506, new_n16507, new_n16508,
    new_n16509, new_n16510, new_n16511, new_n16512, new_n16513, new_n16514,
    new_n16515, new_n16516, new_n16517, new_n16518, new_n16519, new_n16520,
    new_n16521, new_n16522, new_n16523, new_n16524, new_n16525, new_n16526,
    new_n16527, new_n16528, new_n16529, new_n16530, new_n16531, new_n16532,
    new_n16533, new_n16534, new_n16535, new_n16536, new_n16537, new_n16538,
    new_n16539, new_n16540, new_n16541, new_n16542, new_n16543, new_n16544,
    new_n16545, new_n16546, new_n16547, new_n16548, new_n16549, new_n16550,
    new_n16551, new_n16552, new_n16553, new_n16554, new_n16555, new_n16556,
    new_n16557, new_n16558, new_n16559, new_n16560, new_n16561, new_n16562,
    new_n16563, new_n16564, new_n16565, new_n16566, new_n16567, new_n16568,
    new_n16569, new_n16570, new_n16571, new_n16572, new_n16573, new_n16574,
    new_n16575, new_n16576, new_n16577, new_n16578, new_n16579, new_n16580,
    new_n16581, new_n16582, new_n16583, new_n16584, new_n16585, new_n16586,
    new_n16587, new_n16588, new_n16589, new_n16590, new_n16591, new_n16592,
    new_n16593, new_n16594, new_n16595, new_n16596, new_n16597, new_n16598,
    new_n16599, new_n16600, new_n16601, new_n16602, new_n16603, new_n16604,
    new_n16605, new_n16606, new_n16607, new_n16608, new_n16609, new_n16610,
    new_n16611, new_n16612, new_n16613, new_n16614, new_n16615, new_n16616,
    new_n16617, new_n16618, new_n16619, new_n16620, new_n16621, new_n16622,
    new_n16623, new_n16624, new_n16625, new_n16626, new_n16627, new_n16628,
    new_n16629, new_n16630, new_n16631, new_n16632, new_n16633, new_n16634,
    new_n16635, new_n16636, new_n16637, new_n16638, new_n16639, new_n16640,
    new_n16641, new_n16642, new_n16643, new_n16644, new_n16645, new_n16646,
    new_n16647, new_n16648, new_n16649, new_n16650, new_n16651, new_n16652,
    new_n16653, new_n16654, new_n16655, new_n16656, new_n16657, new_n16658,
    new_n16659, new_n16660, new_n16661, new_n16662, new_n16663, new_n16664,
    new_n16665, new_n16666, new_n16667, new_n16668, new_n16669, new_n16670,
    new_n16671, new_n16672, new_n16673, new_n16674, new_n16675, new_n16676,
    new_n16677, new_n16678, new_n16679, new_n16680, new_n16681, new_n16682,
    new_n16683, new_n16684, new_n16685, new_n16686, new_n16687, new_n16688,
    new_n16689, new_n16690, new_n16691, new_n16692, new_n16693, new_n16694,
    new_n16695, new_n16696, new_n16697, new_n16698, new_n16699, new_n16700,
    new_n16701, new_n16702, new_n16703, new_n16704, new_n16705, new_n16706,
    new_n16707, new_n16708, new_n16709, new_n16710, new_n16711, new_n16712,
    new_n16713, new_n16714, new_n16715, new_n16716, new_n16717, new_n16718,
    new_n16719, new_n16720, new_n16721, new_n16722, new_n16723, new_n16724,
    new_n16725, new_n16726, new_n16727, new_n16728, new_n16729, new_n16730,
    new_n16731, new_n16732, new_n16733, new_n16734, new_n16735, new_n16736,
    new_n16737, new_n16738, new_n16739, new_n16740, new_n16741, new_n16742,
    new_n16743, new_n16744, new_n16745, new_n16746, new_n16747, new_n16748,
    new_n16749, new_n16750, new_n16751, new_n16752, new_n16753, new_n16754,
    new_n16755, new_n16756, new_n16757, new_n16758, new_n16759, new_n16760,
    new_n16761, new_n16762, new_n16763, new_n16764, new_n16765, new_n16766,
    new_n16767, new_n16768, new_n16769, new_n16770, new_n16771, new_n16772,
    new_n16773, new_n16774, new_n16775, new_n16776, new_n16777, new_n16778,
    new_n16779, new_n16780, new_n16781, new_n16782, new_n16783, new_n16784,
    new_n16785, new_n16786, new_n16787, new_n16788, new_n16789, new_n16790,
    new_n16791, new_n16792, new_n16793, new_n16794, new_n16795, new_n16796,
    new_n16797, new_n16798, new_n16799, new_n16800, new_n16801, new_n16802,
    new_n16803, new_n16804, new_n16805, new_n16806, new_n16807, new_n16808,
    new_n16809, new_n16810, new_n16811, new_n16812, new_n16813, new_n16814,
    new_n16815, new_n16816, new_n16817, new_n16818, new_n16819, new_n16820,
    new_n16821, new_n16822, new_n16823, new_n16824, new_n16825, new_n16826,
    new_n16827, new_n16828, new_n16829, new_n16830, new_n16831, new_n16832,
    new_n16833, new_n16834, new_n16835, new_n16836, new_n16837, new_n16838,
    new_n16839, new_n16840, new_n16841, new_n16842, new_n16843, new_n16844,
    new_n16845, new_n16846, new_n16847, new_n16848, new_n16849, new_n16850,
    new_n16851, new_n16852, new_n16853, new_n16854, new_n16855, new_n16856,
    new_n16857, new_n16858, new_n16859, new_n16860, new_n16861, new_n16862,
    new_n16863, new_n16864, new_n16865, new_n16866, new_n16867, new_n16868,
    new_n16869, new_n16870, new_n16871, new_n16872, new_n16873, new_n16874,
    new_n16875, new_n16876, new_n16877, new_n16878, new_n16879, new_n16880,
    new_n16881, new_n16882, new_n16883, new_n16884, new_n16885, new_n16886,
    new_n16887, new_n16888, new_n16889, new_n16890, new_n16891, new_n16892,
    new_n16893, new_n16894, new_n16895, new_n16896, new_n16897, new_n16898,
    new_n16899, new_n16900, new_n16901, new_n16902, new_n16903, new_n16904,
    new_n16905, new_n16906, new_n16907, new_n16908, new_n16909, new_n16910,
    new_n16911, new_n16912, new_n16913, new_n16914, new_n16915, new_n16916,
    new_n16917, new_n16918, new_n16919, new_n16920, new_n16921, new_n16922,
    new_n16923, new_n16924, new_n16925, new_n16926, new_n16927, new_n16928,
    new_n16929, new_n16930, new_n16931, new_n16932, new_n16933, new_n16934,
    new_n16935, new_n16936, new_n16937, new_n16938, new_n16939, new_n16940,
    new_n16941, new_n16942, new_n16943, new_n16944, new_n16945, new_n16946,
    new_n16947, new_n16948, new_n16949, new_n16950, new_n16951, new_n16952,
    new_n16953, new_n16954, new_n16955, new_n16956, new_n16957, new_n16958,
    new_n16959, new_n16960, new_n16961, new_n16962, new_n16963, new_n16964,
    new_n16965, new_n16966, new_n16967, new_n16968, new_n16969, new_n16970,
    new_n16971, new_n16972, new_n16973, new_n16974, new_n16975, new_n16976,
    new_n16977, new_n16978, new_n16979, new_n16980, new_n16981, new_n16982,
    new_n16983, new_n16984, new_n16985, new_n16986, new_n16987, new_n16988,
    new_n16989, new_n16990, new_n16991, new_n16992, new_n16993, new_n16994,
    new_n16995, new_n16996, new_n16997, new_n16998, new_n16999, new_n17000,
    new_n17001, new_n17002, new_n17003, new_n17004, new_n17005, new_n17006,
    new_n17007, new_n17008, new_n17009, new_n17010, new_n17011, new_n17012,
    new_n17013, new_n17014, new_n17015, new_n17016, new_n17017, new_n17018,
    new_n17019, new_n17020, new_n17021, new_n17022, new_n17023, new_n17024,
    new_n17025, new_n17026, new_n17027, new_n17028, new_n17029, new_n17030,
    new_n17031, new_n17032, new_n17033, new_n17034, new_n17035, new_n17036,
    new_n17037, new_n17038, new_n17039, new_n17040, new_n17041, new_n17042,
    new_n17043, new_n17044, new_n17045, new_n17046, new_n17047, new_n17048,
    new_n17049, new_n17050, new_n17051, new_n17052, new_n17053, new_n17054,
    new_n17055, new_n17056, new_n17057, new_n17058, new_n17059, new_n17060,
    new_n17061, new_n17062, new_n17063, new_n17064, new_n17065, new_n17066,
    new_n17067, new_n17068, new_n17069, new_n17070, new_n17071, new_n17072,
    new_n17073, new_n17074, new_n17075, new_n17076, new_n17077, new_n17078,
    new_n17079, new_n17080, new_n17081, new_n17082, new_n17083, new_n17084,
    new_n17085, new_n17086, new_n17087, new_n17088, new_n17089, new_n17090,
    new_n17091, new_n17092, new_n17093, new_n17094, new_n17095, new_n17096,
    new_n17097, new_n17098, new_n17099, new_n17100, new_n17101, new_n17102,
    new_n17103, new_n17104, new_n17105, new_n17106, new_n17107, new_n17108,
    new_n17109, new_n17110, new_n17111, new_n17112, new_n17113, new_n17114,
    new_n17115, new_n17116, new_n17117, new_n17118, new_n17119, new_n17120,
    new_n17121, new_n17122, new_n17123, new_n17124, new_n17125, new_n17126,
    new_n17127, new_n17128, new_n17129, new_n17130, new_n17131, new_n17132,
    new_n17133, new_n17134, new_n17135, new_n17136, new_n17137, new_n17138,
    new_n17139, new_n17140, new_n17141, new_n17142, new_n17143, new_n17144,
    new_n17145, new_n17146, new_n17147, new_n17148, new_n17149, new_n17150,
    new_n17151, new_n17152, new_n17153, new_n17154, new_n17155, new_n17156,
    new_n17157, new_n17158, new_n17159, new_n17160, new_n17161, new_n17162,
    new_n17163, new_n17164, new_n17165, new_n17166, new_n17167, new_n17168,
    new_n17169, new_n17170, new_n17171, new_n17172, new_n17173, new_n17174,
    new_n17175, new_n17176, new_n17177, new_n17178, new_n17179, new_n17180,
    new_n17181, new_n17182, new_n17183, new_n17184, new_n17185, new_n17186,
    new_n17187, new_n17188, new_n17189, new_n17190, new_n17191, new_n17192,
    new_n17193, new_n17194, new_n17195, new_n17196, new_n17197, new_n17198,
    new_n17199, new_n17200, new_n17201, new_n17202, new_n17203, new_n17204,
    new_n17205, new_n17206, new_n17207, new_n17208, new_n17209, new_n17210,
    new_n17211, new_n17212, new_n17213, new_n17214, new_n17215, new_n17216,
    new_n17217, new_n17218, new_n17219, new_n17220, new_n17221, new_n17222,
    new_n17223, new_n17224, new_n17225, new_n17226, new_n17227, new_n17228,
    new_n17229, new_n17230, new_n17231, new_n17232, new_n17233, new_n17234,
    new_n17235, new_n17236, new_n17237, new_n17238, new_n17239, new_n17240,
    new_n17241, new_n17242, new_n17243, new_n17244, new_n17245, new_n17246,
    new_n17247, new_n17248, new_n17249, new_n17250, new_n17251, new_n17252,
    new_n17253, new_n17254, new_n17255, new_n17256, new_n17257, new_n17258,
    new_n17259, new_n17260, new_n17261, new_n17262, new_n17263, new_n17264,
    new_n17265, new_n17266, new_n17267, new_n17268, new_n17269, new_n17270,
    new_n17271, new_n17272, new_n17273, new_n17274, new_n17275, new_n17276,
    new_n17277, new_n17278, new_n17279, new_n17280, new_n17281, new_n17282,
    new_n17283, new_n17284, new_n17285, new_n17286, new_n17287, new_n17288,
    new_n17289, new_n17290, new_n17291, new_n17292, new_n17293, new_n17294,
    new_n17295, new_n17296, new_n17297, new_n17298, new_n17299, new_n17300,
    new_n17301, new_n17302, new_n17303, new_n17304, new_n17305, new_n17306,
    new_n17307, new_n17308, new_n17309, new_n17310, new_n17311, new_n17312,
    new_n17313, new_n17314, new_n17315, new_n17316, new_n17317, new_n17318,
    new_n17319, new_n17320, new_n17321, new_n17322, new_n17323, new_n17324,
    new_n17325, new_n17326, new_n17327, new_n17328, new_n17329, new_n17330,
    new_n17331, new_n17332, new_n17333, new_n17334, new_n17335, new_n17336,
    new_n17337, new_n17338, new_n17339, new_n17340, new_n17341, new_n17342,
    new_n17343, new_n17344, new_n17345, new_n17346, new_n17347, new_n17348,
    new_n17349, new_n17350, new_n17351, new_n17352, new_n17353, new_n17354,
    new_n17355, new_n17356, new_n17357, new_n17358, new_n17359, new_n17360,
    new_n17361, new_n17362, new_n17363, new_n17364, new_n17365, new_n17366,
    new_n17367, new_n17368, new_n17369, new_n17370, new_n17371, new_n17372,
    new_n17373, new_n17374, new_n17375, new_n17376, new_n17377, new_n17378,
    new_n17379, new_n17380, new_n17381, new_n17382, new_n17383, new_n17384,
    new_n17385, new_n17386, new_n17387, new_n17388, new_n17389, new_n17390,
    new_n17391, new_n17392, new_n17393, new_n17394, new_n17395, new_n17396,
    new_n17397, new_n17398, new_n17399, new_n17400, new_n17401, new_n17402,
    new_n17403, new_n17404, new_n17405, new_n17406, new_n17407, new_n17408,
    new_n17409, new_n17410, new_n17411, new_n17412, new_n17413, new_n17414,
    new_n17415, new_n17416, new_n17417, new_n17418, new_n17419, new_n17420,
    new_n17421, new_n17422, new_n17423, new_n17424, new_n17425, new_n17426,
    new_n17427, new_n17428, new_n17429, new_n17430, new_n17431, new_n17432,
    new_n17433, new_n17434, new_n17435, new_n17436, new_n17437, new_n17438,
    new_n17439, new_n17440, new_n17441, new_n17442, new_n17443, new_n17444,
    new_n17445, new_n17446, new_n17447, new_n17448, new_n17449, new_n17450,
    new_n17451, new_n17452, new_n17453, new_n17454, new_n17455, new_n17456,
    new_n17457, new_n17458, new_n17459, new_n17460, new_n17461, new_n17462,
    new_n17463, new_n17464, new_n17465, new_n17466, new_n17467, new_n17468,
    new_n17469, new_n17470, new_n17471, new_n17472, new_n17473, new_n17474,
    new_n17475, new_n17476, new_n17477, new_n17478, new_n17479, new_n17480,
    new_n17481, new_n17482, new_n17483, new_n17484, new_n17485, new_n17486,
    new_n17487, new_n17488, new_n17489, new_n17490, new_n17491, new_n17492,
    new_n17493, new_n17494, new_n17495, new_n17496, new_n17497, new_n17498,
    new_n17499, new_n17500, new_n17501, new_n17502, new_n17503, new_n17504,
    new_n17505, new_n17506, new_n17507, new_n17508, new_n17509, new_n17510,
    new_n17511, new_n17512, new_n17513, new_n17514, new_n17515, new_n17516,
    new_n17517, new_n17518, new_n17519, new_n17520, new_n17521, new_n17522,
    new_n17523, new_n17524, new_n17525, new_n17526, new_n17527, new_n17528,
    new_n17529, new_n17530, new_n17531, new_n17532, new_n17533, new_n17534,
    new_n17535, new_n17536, new_n17537, new_n17538, new_n17539, new_n17540,
    new_n17541, new_n17542, new_n17543, new_n17544, new_n17545, new_n17546,
    new_n17547, new_n17548, new_n17549, new_n17550, new_n17551, new_n17552,
    new_n17553, new_n17554, new_n17555, new_n17556, new_n17557, new_n17558,
    new_n17559, new_n17560, new_n17561, new_n17562, new_n17563, new_n17564,
    new_n17565, new_n17566, new_n17567, new_n17568, new_n17569, new_n17570,
    new_n17571, new_n17572, new_n17573, new_n17574, new_n17575, new_n17576,
    new_n17577, new_n17578, new_n17579, new_n17580, new_n17581, new_n17582,
    new_n17583, new_n17584, new_n17585, new_n17586, new_n17587, new_n17588,
    new_n17589, new_n17590, new_n17591, new_n17592, new_n17593, new_n17594,
    new_n17595, new_n17596, new_n17597, new_n17598, new_n17599, new_n17600,
    new_n17601, new_n17602, new_n17603, new_n17604, new_n17605, new_n17606,
    new_n17607, new_n17608, new_n17609, new_n17610, new_n17611, new_n17612,
    new_n17613, new_n17614, new_n17615, new_n17616, new_n17617, new_n17618,
    new_n17619, new_n17620, new_n17621, new_n17622, new_n17623, new_n17624,
    new_n17625, new_n17626, new_n17627, new_n17628, new_n17629, new_n17630,
    new_n17631, new_n17632, new_n17633, new_n17634, new_n17635, new_n17636,
    new_n17637, new_n17638, new_n17639, new_n17640, new_n17641, new_n17642,
    new_n17643, new_n17644, new_n17645, new_n17646, new_n17647, new_n17648,
    new_n17649, new_n17650, new_n17651, new_n17652, new_n17653, new_n17654,
    new_n17655, new_n17656, new_n17657, new_n17658, new_n17659, new_n17660,
    new_n17661, new_n17662, new_n17663, new_n17664, new_n17665, new_n17666,
    new_n17667, new_n17668, new_n17669, new_n17670, new_n17671, new_n17672,
    new_n17673, new_n17674, new_n17675, new_n17676, new_n17677, new_n17678,
    new_n17679, new_n17680, new_n17681, new_n17682, new_n17683, new_n17684,
    new_n17685, new_n17686, new_n17687, new_n17688, new_n17689, new_n17690,
    new_n17691, new_n17692, new_n17693, new_n17694, new_n17695, new_n17696,
    new_n17697, new_n17698, new_n17699, new_n17700, new_n17701, new_n17702,
    new_n17703, new_n17704, new_n17705, new_n17706, new_n17707, new_n17708,
    new_n17709, new_n17710, new_n17711, new_n17712, new_n17713, new_n17714,
    new_n17715, new_n17716, new_n17717, new_n17718, new_n17719, new_n17720,
    new_n17721, new_n17722, new_n17723, new_n17724, new_n17725, new_n17726,
    new_n17727, new_n17728, new_n17729, new_n17730, new_n17731, new_n17732,
    new_n17733, new_n17734, new_n17735, new_n17736, new_n17737, new_n17738,
    new_n17739, new_n17740, new_n17741, new_n17742, new_n17743, new_n17744,
    new_n17745, new_n17746, new_n17747, new_n17748, new_n17749, new_n17750,
    new_n17751, new_n17752, new_n17753, new_n17754, new_n17755, new_n17756,
    new_n17757, new_n17758, new_n17759, new_n17760, new_n17761, new_n17762,
    new_n17763, new_n17764, new_n17765, new_n17766, new_n17767, new_n17768,
    new_n17769, new_n17770, new_n17771, new_n17772, new_n17773, new_n17774,
    new_n17775, new_n17776, new_n17777, new_n17778, new_n17779, new_n17780,
    new_n17781, new_n17782, new_n17783, new_n17784, new_n17785, new_n17786,
    new_n17787, new_n17788, new_n17789, new_n17790, new_n17791, new_n17792,
    new_n17793, new_n17794, new_n17795, new_n17796, new_n17797, new_n17798,
    new_n17799, new_n17800, new_n17801, new_n17802, new_n17803, new_n17804,
    new_n17805, new_n17806, new_n17807, new_n17808, new_n17809, new_n17810,
    new_n17811, new_n17812, new_n17813, new_n17814, new_n17815, new_n17816,
    new_n17817, new_n17818, new_n17819, new_n17820, new_n17821, new_n17822,
    new_n17823, new_n17824, new_n17825, new_n17826, new_n17827, new_n17828,
    new_n17829, new_n17830, new_n17831, new_n17832, new_n17833, new_n17834,
    new_n17835, new_n17836, new_n17837, new_n17838, new_n17839, new_n17840,
    new_n17841, new_n17842, new_n17843, new_n17844, new_n17845, new_n17846,
    new_n17847, new_n17848, new_n17849, new_n17850, new_n17851, new_n17852,
    new_n17853, new_n17854, new_n17855, new_n17856, new_n17857, new_n17858,
    new_n17859, new_n17860, new_n17861, new_n17862, new_n17863, new_n17864,
    new_n17865, new_n17866, new_n17867, new_n17868, new_n17869, new_n17870,
    new_n17871, new_n17872, new_n17873, new_n17874, new_n17875, new_n17876,
    new_n17877, new_n17878, new_n17879, new_n17880, new_n17881, new_n17882,
    new_n17883, new_n17884, new_n17885, new_n17886, new_n17887, new_n17888,
    new_n17889, new_n17890, new_n17891, new_n17892, new_n17893, new_n17894,
    new_n17895, new_n17896, new_n17897, new_n17898, new_n17899, new_n17900,
    new_n17901, new_n17902, new_n17903, new_n17904, new_n17905, new_n17906,
    new_n17907, new_n17908, new_n17909, new_n17910, new_n17911, new_n17912,
    new_n17913, new_n17914, new_n17915, new_n17916, new_n17917, new_n17918,
    new_n17919, new_n17920, new_n17921, new_n17922, new_n17923, new_n17924,
    new_n17925, new_n17926, new_n17927, new_n17928, new_n17929, new_n17930,
    new_n17931, new_n17932, new_n17933, new_n17934, new_n17935, new_n17936,
    new_n17937, new_n17938, new_n17939, new_n17940, new_n17941, new_n17942,
    new_n17943, new_n17944, new_n17945, new_n17946, new_n17947, new_n17948,
    new_n17949, new_n17950, new_n17951, new_n17952, new_n17953, new_n17954,
    new_n17955, new_n17956, new_n17957, new_n17958, new_n17959, new_n17960,
    new_n17961, new_n17962, new_n17963, new_n17964, new_n17965, new_n17966,
    new_n17967, new_n17968, new_n17969, new_n17970, new_n17971, new_n17972,
    new_n17973, new_n17974, new_n17975, new_n17976, new_n17977, new_n17978,
    new_n17979, new_n17980, new_n17981, new_n17982, new_n17983, new_n17984,
    new_n17985, new_n17986, new_n17987, new_n17988, new_n17989, new_n17990,
    new_n17991, new_n17992, new_n17993, new_n17994, new_n17995, new_n17996,
    new_n17997, new_n17998, new_n17999, new_n18000, new_n18001, new_n18002,
    new_n18003, new_n18004, new_n18005, new_n18006, new_n18007, new_n18008,
    new_n18009, new_n18010, new_n18011, new_n18012, new_n18013, new_n18014,
    new_n18015, new_n18016, new_n18017, new_n18018, new_n18019, new_n18020,
    new_n18021, new_n18022, new_n18023, new_n18024, new_n18025, new_n18026,
    new_n18027, new_n18028, new_n18029, new_n18030, new_n18031, new_n18032,
    new_n18033, new_n18034, new_n18035, new_n18036, new_n18037, new_n18038,
    new_n18039, new_n18040, new_n18041, new_n18042, new_n18043, new_n18044,
    new_n18045, new_n18046, new_n18047, new_n18048, new_n18049, new_n18050,
    new_n18051, new_n18052, new_n18053, new_n18054, new_n18055, new_n18056,
    new_n18057, new_n18058, new_n18059, new_n18060, new_n18061, new_n18062,
    new_n18063, new_n18064, new_n18065, new_n18066, new_n18067, new_n18068,
    new_n18069, new_n18070, new_n18071, new_n18072, new_n18073, new_n18074,
    new_n18075, new_n18076, new_n18077, new_n18078, new_n18079, new_n18080,
    new_n18081, new_n18082, new_n18083, new_n18084, new_n18085, new_n18086,
    new_n18087, new_n18088, new_n18089, new_n18090, new_n18091, new_n18092,
    new_n18093, new_n18094, new_n18095, new_n18096, new_n18097, new_n18098,
    new_n18099, new_n18100, new_n18101, new_n18102, new_n18103, new_n18104,
    new_n18105, new_n18106, new_n18107, new_n18108, new_n18109, new_n18110,
    new_n18111, new_n18112, new_n18113, new_n18114, new_n18115, new_n18116,
    new_n18117, new_n18118, new_n18119, new_n18120, new_n18121, new_n18122,
    new_n18123, new_n18124, new_n18125, new_n18126, new_n18127, new_n18128,
    new_n18129, new_n18130, new_n18131, new_n18132, new_n18133, new_n18134,
    new_n18135, new_n18136, new_n18137, new_n18138, new_n18139, new_n18140,
    new_n18141, new_n18142, new_n18143, new_n18144, new_n18145, new_n18146,
    new_n18147, new_n18148, new_n18149, new_n18150, new_n18151, new_n18152,
    new_n18153, new_n18154, new_n18155, new_n18156, new_n18157, new_n18158,
    new_n18159, new_n18160, new_n18161, new_n18162, new_n18163, new_n18164,
    new_n18165, new_n18166, new_n18167, new_n18168, new_n18169, new_n18170,
    new_n18171, new_n18172, new_n18173, new_n18174, new_n18175, new_n18176,
    new_n18177, new_n18178, new_n18179, new_n18180, new_n18181, new_n18182,
    new_n18183, new_n18184, new_n18185, new_n18186, new_n18187, new_n18188,
    new_n18189, new_n18190, new_n18191, new_n18192, new_n18193, new_n18194,
    new_n18195, new_n18196, new_n18197, new_n18198, new_n18199, new_n18200,
    new_n18201, new_n18202, new_n18203, new_n18204, new_n18205, new_n18206,
    new_n18207, new_n18208, new_n18209, new_n18210, new_n18211, new_n18212,
    new_n18213, new_n18214, new_n18215, new_n18216, new_n18217, new_n18218,
    new_n18219, new_n18220, new_n18221, new_n18222, new_n18223, new_n18224,
    new_n18225, new_n18226, new_n18227, new_n18228, new_n18229, new_n18230,
    new_n18231, new_n18232, new_n18233, new_n18234, new_n18235, new_n18236,
    new_n18237, new_n18238, new_n18239, new_n18240, new_n18241, new_n18242,
    new_n18243, new_n18244, new_n18245, new_n18246, new_n18247, new_n18248,
    new_n18249, new_n18250, new_n18251, new_n18252, new_n18253, new_n18254,
    new_n18255, new_n18256, new_n18257, new_n18258, new_n18259, new_n18260,
    new_n18261, new_n18262, new_n18263, new_n18264, new_n18265, new_n18266,
    new_n18267, new_n18268, new_n18269, new_n18270, new_n18271, new_n18272,
    new_n18273, new_n18274, new_n18275, new_n18276, new_n18277, new_n18278,
    new_n18279, new_n18280, new_n18281, new_n18282, new_n18283, new_n18284,
    new_n18285, new_n18286, new_n18287, new_n18288, new_n18289, new_n18290,
    new_n18291, new_n18292, new_n18293, new_n18294, new_n18295, new_n18296,
    new_n18297, new_n18298, new_n18299, new_n18300, new_n18301, new_n18302,
    new_n18303, new_n18304, new_n18305, new_n18306, new_n18307, new_n18308,
    new_n18309, new_n18310, new_n18311, new_n18312, new_n18313, new_n18314,
    new_n18315, new_n18316, new_n18317, new_n18318, new_n18319, new_n18320,
    new_n18321, new_n18322, new_n18323, new_n18324, new_n18325, new_n18326,
    new_n18327, new_n18328, new_n18329, new_n18330, new_n18331, new_n18332,
    new_n18333, new_n18334, new_n18335, new_n18336, new_n18337, new_n18338,
    new_n18339, new_n18340, new_n18341, new_n18342, new_n18343, new_n18344,
    new_n18345, new_n18346, new_n18347, new_n18348, new_n18349, new_n18350,
    new_n18351, new_n18352, new_n18353, new_n18354, new_n18355, new_n18356,
    new_n18357, new_n18358, new_n18359, new_n18360, new_n18361, new_n18362,
    new_n18363, new_n18364, new_n18365, new_n18366, new_n18367, new_n18368,
    new_n18369, new_n18370, new_n18371, new_n18372, new_n18373, new_n18374,
    new_n18375, new_n18376, new_n18377, new_n18378, new_n18379, new_n18380,
    new_n18381, new_n18382, new_n18383, new_n18384, new_n18385, new_n18386,
    new_n18387, new_n18388, new_n18389, new_n18390, new_n18391, new_n18392,
    new_n18393, new_n18394, new_n18395, new_n18396, new_n18397, new_n18398,
    new_n18399, new_n18400, new_n18401, new_n18402, new_n18403, new_n18404,
    new_n18405, new_n18406, new_n18407, new_n18408, new_n18409, new_n18410,
    new_n18411, new_n18412, new_n18413, new_n18414, new_n18415, new_n18416,
    new_n18417, new_n18418, new_n18419, new_n18420, new_n18421, new_n18422,
    new_n18423, new_n18424, new_n18425, new_n18426, new_n18427, new_n18428,
    new_n18429, new_n18430, new_n18431, new_n18432, new_n18433, new_n18434,
    new_n18435, new_n18436, new_n18437, new_n18438, new_n18439, new_n18440,
    new_n18441, new_n18442, new_n18443, new_n18444, new_n18445, new_n18446,
    new_n18447, new_n18448, new_n18449, new_n18450, new_n18451, new_n18452,
    new_n18453, new_n18454, new_n18455, new_n18456, new_n18457, new_n18458,
    new_n18459, new_n18460, new_n18461, new_n18462, new_n18463, new_n18464,
    new_n18465, new_n18466, new_n18467, new_n18468, new_n18469, new_n18470,
    new_n18471, new_n18472, new_n18473, new_n18474, new_n18475, new_n18476,
    new_n18477, new_n18478, new_n18479, new_n18480, new_n18481, new_n18482,
    new_n18483, new_n18484, new_n18485, new_n18486, new_n18487, new_n18488,
    new_n18489, new_n18490, new_n18491, new_n18492, new_n18493, new_n18494,
    new_n18495, new_n18496, new_n18497, new_n18498, new_n18499, new_n18500,
    new_n18501, new_n18502, new_n18503, new_n18504, new_n18505, new_n18506,
    new_n18507, new_n18508, new_n18509, new_n18510, new_n18511, new_n18512,
    new_n18513, new_n18514, new_n18515, new_n18516, new_n18517, new_n18518,
    new_n18519, new_n18520, new_n18521, new_n18522, new_n18523, new_n18524,
    new_n18525, new_n18526, new_n18527, new_n18528, new_n18529, new_n18530,
    new_n18531, new_n18532, new_n18533, new_n18534, new_n18535, new_n18536,
    new_n18537, new_n18538, new_n18539, new_n18540, new_n18541, new_n18542,
    new_n18543, new_n18544, new_n18545, new_n18546, new_n18547, new_n18548,
    new_n18549, new_n18550, new_n18551, new_n18552, new_n18553, new_n18554,
    new_n18555, new_n18556, new_n18557, new_n18558, new_n18559, new_n18560,
    new_n18561, new_n18562, new_n18563, new_n18564, new_n18565, new_n18566,
    new_n18567, new_n18568, new_n18569, new_n18570, new_n18571, new_n18572,
    new_n18573, new_n18574, new_n18575, new_n18576, new_n18577, new_n18578,
    new_n18579, new_n18580, new_n18581, new_n18582, new_n18583, new_n18584,
    new_n18585, new_n18586, new_n18587, new_n18588, new_n18589, new_n18590,
    new_n18591, new_n18592, new_n18593, new_n18594, new_n18595, new_n18596,
    new_n18597, new_n18598, new_n18599, new_n18600, new_n18601, new_n18602,
    new_n18603, new_n18604, new_n18605, new_n18606, new_n18607, new_n18608,
    new_n18609, new_n18610, new_n18611, new_n18612, new_n18613, new_n18614,
    new_n18615, new_n18616, new_n18617, new_n18618, new_n18619, new_n18620,
    new_n18621, new_n18622, new_n18623, new_n18624, new_n18625, new_n18626,
    new_n18627, new_n18628, new_n18629, new_n18630, new_n18631, new_n18632,
    new_n18633, new_n18634, new_n18635, new_n18636, new_n18637, new_n18638,
    new_n18639, new_n18640, new_n18641, new_n18642, new_n18643, new_n18644,
    new_n18645, new_n18646, new_n18647, new_n18648, new_n18649, new_n18650,
    new_n18651, new_n18652, new_n18653, new_n18654, new_n18655, new_n18656,
    new_n18657, new_n18658, new_n18659, new_n18660, new_n18661, new_n18662,
    new_n18663, new_n18664, new_n18665, new_n18666, new_n18667, new_n18668,
    new_n18669, new_n18670, new_n18671, new_n18672, new_n18673, new_n18674,
    new_n18675, new_n18676, new_n18677, new_n18678, new_n18679, new_n18680,
    new_n18681, new_n18682, new_n18683, new_n18684, new_n18685, new_n18686,
    new_n18687, new_n18688, new_n18689, new_n18690, new_n18691, new_n18692,
    new_n18693, new_n18694, new_n18695, new_n18696, new_n18697, new_n18698,
    new_n18699, new_n18700, new_n18701, new_n18702, new_n18703, new_n18704,
    new_n18705, new_n18706, new_n18707, new_n18708, new_n18709, new_n18710,
    new_n18711, new_n18712, new_n18713, new_n18714, new_n18715, new_n18716,
    new_n18717, new_n18718, new_n18719, new_n18720, new_n18721, new_n18722,
    new_n18723, new_n18724, new_n18725, new_n18726, new_n18727, new_n18728,
    new_n18729, new_n18730, new_n18731, new_n18732, new_n18733, new_n18734,
    new_n18735, new_n18736, new_n18737, new_n18738, new_n18739, new_n18740,
    new_n18741, new_n18742, new_n18743, new_n18744, new_n18745, new_n18746,
    new_n18747, new_n18748, new_n18749, new_n18750, new_n18751, new_n18752,
    new_n18753, new_n18754, new_n18755, new_n18756, new_n18757, new_n18758,
    new_n18759, new_n18760, new_n18761, new_n18762, new_n18763, new_n18764,
    new_n18765, new_n18766, new_n18767, new_n18768, new_n18769, new_n18770,
    new_n18771, new_n18772, new_n18773, new_n18774, new_n18775, new_n18776,
    new_n18777, new_n18778, new_n18779, new_n18780, new_n18781, new_n18782,
    new_n18783, new_n18784, new_n18785, new_n18786, new_n18787, new_n18788,
    new_n18789, new_n18790, new_n18791, new_n18792, new_n18793, new_n18794,
    new_n18795, new_n18796, new_n18797, new_n18798, new_n18799, new_n18800,
    new_n18801, new_n18802, new_n18803, new_n18804, new_n18805, new_n18806,
    new_n18807, new_n18808, new_n18809, new_n18810, new_n18811, new_n18812,
    new_n18813, new_n18814, new_n18815, new_n18816, new_n18817, new_n18818,
    new_n18819, new_n18820, new_n18821, new_n18822, new_n18823, new_n18824,
    new_n18825, new_n18826, new_n18827, new_n18828, new_n18829, new_n18830,
    new_n18831, new_n18832, new_n18833, new_n18834, new_n18835, new_n18836,
    new_n18837, new_n18838, new_n18839, new_n18840, new_n18841, new_n18842,
    new_n18843, new_n18844, new_n18845, new_n18846, new_n18847, new_n18848,
    new_n18849, new_n18850, new_n18851, new_n18852, new_n18853, new_n18854,
    new_n18855, new_n18856, new_n18857, new_n18858, new_n18859, new_n18860,
    new_n18861, new_n18862, new_n18863, new_n18864, new_n18865, new_n18866,
    new_n18867, new_n18868, new_n18869, new_n18870, new_n18871, new_n18872,
    new_n18873, new_n18874, new_n18875, new_n18876, new_n18877, new_n18878,
    new_n18879, new_n18880, new_n18881, new_n18882, new_n18883, new_n18884,
    new_n18885, new_n18886, new_n18887, new_n18888, new_n18889, new_n18890,
    new_n18891, new_n18892, new_n18893, new_n18894, new_n18895, new_n18896,
    new_n18897, new_n18898, new_n18899, new_n18900, new_n18901, new_n18902,
    new_n18903, new_n18904, new_n18905, new_n18906, new_n18907, new_n18908,
    new_n18909, new_n18910, new_n18911, new_n18912, new_n18913, new_n18914,
    new_n18915, new_n18916, new_n18917, new_n18918, new_n18919, new_n18920,
    new_n18921, new_n18922, new_n18923, new_n18924, new_n18925, new_n18926,
    new_n18927, new_n18928, new_n18929, new_n18930, new_n18931, new_n18932,
    new_n18933, new_n18934, new_n18935, new_n18936, new_n18937, new_n18938,
    new_n18939, new_n18940, new_n18941, new_n18942, new_n18943, new_n18944,
    new_n18945, new_n18946, new_n18947, new_n18948, new_n18949, new_n18950,
    new_n18951, new_n18952, new_n18953, new_n18954, new_n18955, new_n18956,
    new_n18957, new_n18958, new_n18959, new_n18960, new_n18961, new_n18962,
    new_n18963, new_n18964, new_n18965, new_n18966, new_n18967, new_n18968,
    new_n18969, new_n18970, new_n18971, new_n18972, new_n18973, new_n18974,
    new_n18975, new_n18976, new_n18977, new_n18978, new_n18979, new_n18980,
    new_n18981, new_n18982, new_n18983, new_n18984, new_n18985, new_n18986,
    new_n18987, new_n18988, new_n18989, new_n18990, new_n18991, new_n18992,
    new_n18993, new_n18994, new_n18995, new_n18996, new_n18997, new_n18998,
    new_n18999, new_n19000, new_n19001, new_n19002, new_n19003, new_n19004,
    new_n19005, new_n19006, new_n19007, new_n19008, new_n19009, new_n19010,
    new_n19011, new_n19012, new_n19013, new_n19014, new_n19015, new_n19016,
    new_n19017, new_n19018, new_n19019, new_n19020, new_n19021, new_n19022,
    new_n19023, new_n19024, new_n19025, new_n19026, new_n19027, new_n19028,
    new_n19029, new_n19030, new_n19031, new_n19032, new_n19033, new_n19034,
    new_n19035, new_n19036, new_n19037, new_n19038, new_n19039, new_n19040,
    new_n19041, new_n19042, new_n19043, new_n19044, new_n19045, new_n19046,
    new_n19047, new_n19048, new_n19049, new_n19050, new_n19051, new_n19052,
    new_n19053, new_n19054, new_n19055, new_n19056, new_n19057, new_n19058,
    new_n19059, new_n19060, new_n19061, new_n19062, new_n19063, new_n19064,
    new_n19065, new_n19066, new_n19067, new_n19068, new_n19069, new_n19070,
    new_n19071, new_n19072, new_n19073, new_n19074, new_n19075, new_n19076,
    new_n19077, new_n19078, new_n19079, new_n19080, new_n19081, new_n19082,
    new_n19083, new_n19084, new_n19085, new_n19086, new_n19087, new_n19088,
    new_n19089, new_n19090, new_n19091, new_n19092, new_n19093, new_n19094,
    new_n19095, new_n19096, new_n19097, new_n19098, new_n19099, new_n19100,
    new_n19101, new_n19102, new_n19103, new_n19104, new_n19105, new_n19106,
    new_n19107, new_n19108, new_n19109, new_n19110, new_n19111, new_n19112,
    new_n19113, new_n19114, new_n19115, new_n19116, new_n19117, new_n19118,
    new_n19119, new_n19120, new_n19121, new_n19122, new_n19123, new_n19124,
    new_n19125, new_n19126, new_n19127, new_n19128, new_n19129, new_n19130,
    new_n19131, new_n19132, new_n19133, new_n19134, new_n19135, new_n19136,
    new_n19137, new_n19138, new_n19139, new_n19140, new_n19141, new_n19142,
    new_n19143, new_n19144, new_n19145, new_n19146, new_n19147, new_n19148,
    new_n19149, new_n19150, new_n19151, new_n19152, new_n19153, new_n19154,
    new_n19155, new_n19156, new_n19157, new_n19158, new_n19159, new_n19160,
    new_n19161, new_n19162, new_n19163, new_n19164, new_n19165, new_n19166,
    new_n19167, new_n19168, new_n19169, new_n19170, new_n19171, new_n19172,
    new_n19173, new_n19174, new_n19175, new_n19176, new_n19177, new_n19178,
    new_n19179, new_n19180, new_n19181, new_n19182, new_n19183, new_n19184,
    new_n19185, new_n19186, new_n19187, new_n19188, new_n19189, new_n19190,
    new_n19191, new_n19192, new_n19193, new_n19194, new_n19195, new_n19196,
    new_n19197, new_n19198, new_n19199, new_n19200, new_n19201, new_n19202,
    new_n19203, new_n19204, new_n19205, new_n19206, new_n19207, new_n19208,
    new_n19209, new_n19210, new_n19211, new_n19212, new_n19213, new_n19214,
    new_n19215, new_n19216, new_n19217, new_n19218, new_n19219, new_n19220,
    new_n19221, new_n19222, new_n19223, new_n19224, new_n19225, new_n19226,
    new_n19227, new_n19228, new_n19229, new_n19230, new_n19231, new_n19232,
    new_n19233, new_n19234, new_n19235, new_n19236, new_n19237, new_n19238,
    new_n19239, new_n19240, new_n19241, new_n19242, new_n19243, new_n19244,
    new_n19245, new_n19246, new_n19247, new_n19248, new_n19249, new_n19250,
    new_n19251, new_n19252, new_n19253, new_n19254, new_n19255, new_n19256,
    new_n19257, new_n19258, new_n19259, new_n19260, new_n19261, new_n19262,
    new_n19263, new_n19264, new_n19265, new_n19266, new_n19267, new_n19268,
    new_n19269, new_n19270, new_n19271, new_n19272, new_n19273, new_n19274,
    new_n19275, new_n19276, new_n19277, new_n19278, new_n19279, new_n19280,
    new_n19281, new_n19282, new_n19283, new_n19284, new_n19285, new_n19286,
    new_n19287, new_n19288, new_n19289, new_n19290, new_n19291, new_n19292,
    new_n19293, new_n19294, new_n19295, new_n19296, new_n19297, new_n19298,
    new_n19299, new_n19300, new_n19301, new_n19302, new_n19303, new_n19304,
    new_n19305, new_n19306, new_n19307, new_n19308, new_n19309, new_n19310,
    new_n19311, new_n19312, new_n19313, new_n19314, new_n19315, new_n19316,
    new_n19317, new_n19318, new_n19319, new_n19320, new_n19321, new_n19322,
    new_n19323, new_n19324, new_n19325, new_n19326, new_n19327, new_n19328,
    new_n19329, new_n19330, new_n19331, new_n19332, new_n19333, new_n19334,
    new_n19335, new_n19336, new_n19337, new_n19338, new_n19339, new_n19340,
    new_n19341, new_n19342, new_n19343, new_n19344, new_n19345, new_n19346,
    new_n19347, new_n19348, new_n19349, new_n19350, new_n19351, new_n19352,
    new_n19353, new_n19354, new_n19355, new_n19356, new_n19357, new_n19358,
    new_n19359, new_n19360, new_n19361, new_n19362, new_n19363, new_n19364,
    new_n19365, new_n19366, new_n19367, new_n19368, new_n19369, new_n19370,
    new_n19371, new_n19372, new_n19373, new_n19374, new_n19375, new_n19376,
    new_n19377, new_n19378, new_n19379, new_n19380, new_n19381, new_n19382,
    new_n19383, new_n19384, new_n19385, new_n19386, new_n19387, new_n19388,
    new_n19389, new_n19390, new_n19391, new_n19392, new_n19393, new_n19394,
    new_n19395, new_n19396, new_n19397, new_n19398, new_n19399, new_n19400,
    new_n19401, new_n19402, new_n19403, new_n19404, new_n19405, new_n19406,
    new_n19407, new_n19408, new_n19409, new_n19410, new_n19411, new_n19412,
    new_n19413, new_n19414, new_n19415, new_n19416, new_n19417, new_n19418,
    new_n19419, new_n19420, new_n19421, new_n19422, new_n19423, new_n19424,
    new_n19425, new_n19426, new_n19427, new_n19428, new_n19429, new_n19430,
    new_n19431, new_n19432, new_n19433, new_n19434, new_n19435, new_n19436,
    new_n19437, new_n19438, new_n19439, new_n19440, new_n19441, new_n19442,
    new_n19443, new_n19444, new_n19445, new_n19446, new_n19447, new_n19448,
    new_n19449, new_n19450, new_n19451, new_n19452, new_n19453, new_n19454,
    new_n19455, new_n19456, new_n19457, new_n19458, new_n19459, new_n19460,
    new_n19461, new_n19462, new_n19463, new_n19464, new_n19465, new_n19466,
    new_n19467, new_n19468, new_n19469, new_n19470, new_n19471, new_n19472,
    new_n19473, new_n19474, new_n19475, new_n19476, new_n19477, new_n19478,
    new_n19479, new_n19480, new_n19481, new_n19482, new_n19483, new_n19484,
    new_n19485, new_n19486, new_n19487, new_n19488, new_n19489, new_n19490,
    new_n19491, new_n19492, new_n19493, new_n19494, new_n19495, new_n19496,
    new_n19497, new_n19498, new_n19499, new_n19500, new_n19501, new_n19502,
    new_n19503, new_n19504, new_n19505, new_n19506, new_n19507, new_n19508,
    new_n19509, new_n19510, new_n19511, new_n19512, new_n19513, new_n19514,
    new_n19515, new_n19516, new_n19517, new_n19518, new_n19519, new_n19520,
    new_n19521, new_n19522, new_n19523, new_n19524, new_n19525, new_n19526,
    new_n19527, new_n19528, new_n19529, new_n19530, new_n19531, new_n19532,
    new_n19533, new_n19534, new_n19535, new_n19536, new_n19537, new_n19538,
    new_n19539, new_n19540, new_n19541, new_n19542, new_n19543, new_n19544,
    new_n19545, new_n19546, new_n19547, new_n19548, new_n19549, new_n19550,
    new_n19551, new_n19552, new_n19553, new_n19554, new_n19555, new_n19556,
    new_n19557, new_n19558, new_n19559, new_n19560, new_n19561, new_n19562,
    new_n19563, new_n19564, new_n19565, new_n19566, new_n19567, new_n19568,
    new_n19569, new_n19570, new_n19571, new_n19572, new_n19573, new_n19574,
    new_n19575, new_n19576, new_n19577, new_n19578, new_n19579, new_n19580,
    new_n19581, new_n19582, new_n19583, new_n19584, new_n19585, new_n19586,
    new_n19587, new_n19588, new_n19589, new_n19590, new_n19591, new_n19592,
    new_n19593, new_n19594, new_n19595, new_n19596, new_n19597, new_n19598,
    new_n19599, new_n19600, new_n19601, new_n19602, new_n19603, new_n19604,
    new_n19605, new_n19606, new_n19607, new_n19608, new_n19609, new_n19610,
    new_n19611, new_n19612, new_n19613, new_n19614, new_n19615, new_n19616,
    new_n19617, new_n19618, new_n19619, new_n19620, new_n19621, new_n19622,
    new_n19623, new_n19624, new_n19625, new_n19626, new_n19627, new_n19628,
    new_n19629, new_n19630, new_n19631, new_n19632, new_n19633, new_n19634,
    new_n19635, new_n19636, new_n19637, new_n19638, new_n19639, new_n19640,
    new_n19641, new_n19642, new_n19643, new_n19644, new_n19645, new_n19646,
    new_n19647, new_n19648, new_n19649, new_n19650, new_n19651, new_n19652,
    new_n19653, new_n19654, new_n19655, new_n19656, new_n19657, new_n19658,
    new_n19659, new_n19660, new_n19661, new_n19662, new_n19663, new_n19664,
    new_n19665, new_n19666, new_n19667, new_n19668, new_n19669, new_n19670,
    new_n19671, new_n19672, new_n19673, new_n19674, new_n19675, new_n19676,
    new_n19677, new_n19678, new_n19679, new_n19680, new_n19681, new_n19682,
    new_n19683, new_n19684, new_n19685, new_n19686, new_n19687, new_n19688,
    new_n19689, new_n19690, new_n19691, new_n19692, new_n19693, new_n19694,
    new_n19695, new_n19696, new_n19697, new_n19698, new_n19699, new_n19700,
    new_n19701, new_n19702, new_n19703, new_n19704, new_n19705, new_n19706,
    new_n19707, new_n19708, new_n19709, new_n19710, new_n19711, new_n19712,
    new_n19713, new_n19714, new_n19715, new_n19716, new_n19717, new_n19718,
    new_n19719, new_n19720, new_n19721, new_n19722, new_n19723, new_n19724,
    new_n19725, new_n19726, new_n19727, new_n19728, new_n19729, new_n19730,
    new_n19731, new_n19732, new_n19733, new_n19734, new_n19735, new_n19736,
    new_n19737, new_n19738, new_n19739, new_n19740, new_n19741, new_n19742,
    new_n19743, new_n19744, new_n19745, new_n19746, new_n19747, new_n19748,
    new_n19749, new_n19750, new_n19751, new_n19752, new_n19753, new_n19754,
    new_n19755, new_n19756, new_n19757, new_n19758, new_n19759, new_n19760,
    new_n19761, new_n19762, new_n19763, new_n19764, new_n19765, new_n19766,
    new_n19767, new_n19768, new_n19769, new_n19770, new_n19771, new_n19772,
    new_n19773, new_n19774, new_n19775, new_n19776, new_n19777, new_n19778,
    new_n19779, new_n19780, new_n19781, new_n19782, new_n19783, new_n19784,
    new_n19785, new_n19786, new_n19787, new_n19788, new_n19789, new_n19790,
    new_n19791, new_n19792, new_n19793, new_n19794, new_n19795, new_n19796,
    new_n19797, new_n19798, new_n19799, new_n19800, new_n19801, new_n19802,
    new_n19803, new_n19804, new_n19805, new_n19806, new_n19807, new_n19808,
    new_n19809, new_n19810, new_n19811, new_n19812, new_n19813, new_n19814,
    new_n19815, new_n19816, new_n19817, new_n19818, new_n19819, new_n19820,
    new_n19821, new_n19822, new_n19823, new_n19824, new_n19825, new_n19826,
    new_n19827, new_n19828, new_n19829, new_n19830, new_n19831, new_n19832,
    new_n19833, new_n19834, new_n19835, new_n19836, new_n19837, new_n19838,
    new_n19839, new_n19840, new_n19841, new_n19842, new_n19843, new_n19844,
    new_n19845, new_n19846, new_n19847, new_n19848, new_n19849, new_n19850,
    new_n19851, new_n19852, new_n19853, new_n19854, new_n19855, new_n19856,
    new_n19857, new_n19858, new_n19859, new_n19860, new_n19861, new_n19862,
    new_n19863, new_n19864, new_n19865, new_n19866, new_n19867, new_n19868,
    new_n19869, new_n19870, new_n19871, new_n19872, new_n19873, new_n19874,
    new_n19875, new_n19876, new_n19877, new_n19878, new_n19879, new_n19880,
    new_n19881, new_n19882, new_n19883, new_n19884, new_n19885, new_n19886,
    new_n19887, new_n19888, new_n19889, new_n19890, new_n19891, new_n19892,
    new_n19893, new_n19894, new_n19895, new_n19896, new_n19897, new_n19898,
    new_n19899, new_n19900, new_n19901, new_n19902, new_n19903, new_n19904,
    new_n19905, new_n19906, new_n19907, new_n19908, new_n19909, new_n19910,
    new_n19911, new_n19912, new_n19913, new_n19914, new_n19915, new_n19916,
    new_n19917, new_n19918, new_n19919, new_n19920, new_n19921, new_n19922,
    new_n19923, new_n19924, new_n19925, new_n19926, new_n19927, new_n19928,
    new_n19929, new_n19930, new_n19931, new_n19932, new_n19933, new_n19934,
    new_n19935, new_n19936, new_n19937, new_n19938, new_n19939, new_n19940,
    new_n19941, new_n19942, new_n19943, new_n19944, new_n19945, new_n19946,
    new_n19947, new_n19948, new_n19949, new_n19950, new_n19951, new_n19952,
    new_n19953, new_n19954, new_n19955, new_n19956, new_n19957, new_n19958,
    new_n19959, new_n19960, new_n19961, new_n19962, new_n19963, new_n19964,
    new_n19965, new_n19966, new_n19967, new_n19968, new_n19969, new_n19970,
    new_n19971, new_n19972, new_n19973, new_n19974, new_n19975, new_n19976,
    new_n19977, new_n19978, new_n19979, new_n19980, new_n19981, new_n19982,
    new_n19983, new_n19984, new_n19985, new_n19986, new_n19987, new_n19988,
    new_n19989, new_n19990, new_n19991, new_n19992, new_n19993, new_n19994,
    new_n19995, new_n19996, new_n19997, new_n19998, new_n19999, new_n20000,
    new_n20001, new_n20002, new_n20003, new_n20004, new_n20005, new_n20006,
    new_n20007, new_n20008, new_n20009, new_n20010, new_n20011, new_n20012,
    new_n20013, new_n20014, new_n20015, new_n20016, new_n20017, new_n20018,
    new_n20019, new_n20020, new_n20021, new_n20022, new_n20023, new_n20024,
    new_n20025, new_n20026, new_n20027, new_n20028, new_n20029, new_n20030,
    new_n20031, new_n20032, new_n20033, new_n20034, new_n20035, new_n20036,
    new_n20037, new_n20038, new_n20039, new_n20040, new_n20041, new_n20042,
    new_n20043, new_n20044, new_n20045, new_n20046, new_n20047, new_n20048,
    new_n20049, new_n20050, new_n20051, new_n20052, new_n20053, new_n20054,
    new_n20055, new_n20056, new_n20057, new_n20058, new_n20059, new_n20060,
    new_n20061, new_n20062, new_n20063, new_n20064, new_n20065, new_n20066,
    new_n20067, new_n20068, new_n20069, new_n20070, new_n20071, new_n20072,
    new_n20073, new_n20074, new_n20075, new_n20076, new_n20077, new_n20078,
    new_n20079, new_n20080, new_n20081, new_n20082, new_n20083, new_n20084,
    new_n20085, new_n20086, new_n20087, new_n20088, new_n20089, new_n20090,
    new_n20091, new_n20092, new_n20093, new_n20094, new_n20095, new_n20096,
    new_n20097, new_n20098, new_n20099, new_n20100, new_n20101, new_n20102,
    new_n20103, new_n20104, new_n20105, new_n20106, new_n20107, new_n20108,
    new_n20109, new_n20110, new_n20111, new_n20112, new_n20113, new_n20114,
    new_n20115, new_n20116, new_n20117, new_n20118, new_n20119, new_n20120,
    new_n20121, new_n20122, new_n20123, new_n20124, new_n20125, new_n20126,
    new_n20127, new_n20128, new_n20129, new_n20130, new_n20131, new_n20132,
    new_n20133, new_n20134, new_n20135, new_n20136, new_n20137, new_n20138,
    new_n20139, new_n20140, new_n20141, new_n20142, new_n20143, new_n20144,
    new_n20145, new_n20146, new_n20147, new_n20148, new_n20149, new_n20150,
    new_n20151, new_n20152, new_n20153, new_n20154, new_n20155, new_n20156,
    new_n20157, new_n20158, new_n20159, new_n20160, new_n20161, new_n20162,
    new_n20163, new_n20164, new_n20165, new_n20166, new_n20167, new_n20168,
    new_n20169, new_n20170, new_n20171, new_n20172, new_n20173, new_n20174,
    new_n20175, new_n20176, new_n20177, new_n20178, new_n20179, new_n20180,
    new_n20181, new_n20182, new_n20183, new_n20184, new_n20185, new_n20186,
    new_n20187, new_n20188, new_n20189, new_n20190, new_n20191, new_n20192,
    new_n20193, new_n20194, new_n20195, new_n20196, new_n20197, new_n20198,
    new_n20199, new_n20200, new_n20201, new_n20202, new_n20203, new_n20204,
    new_n20205, new_n20206, new_n20207, new_n20208, new_n20209, new_n20210,
    new_n20211, new_n20212, new_n20213, new_n20214, new_n20215, new_n20216,
    new_n20217, new_n20218, new_n20219, new_n20220, new_n20221, new_n20222,
    new_n20223, new_n20224, new_n20225, new_n20226, new_n20227, new_n20228,
    new_n20229, new_n20230, new_n20231, new_n20232, new_n20233, new_n20234,
    new_n20235, new_n20236, new_n20237, new_n20238, new_n20239, new_n20240,
    new_n20241, new_n20242, new_n20243, new_n20244, new_n20245, new_n20246,
    new_n20247, new_n20248, new_n20249, new_n20250, new_n20251, new_n20252,
    new_n20253, new_n20254, new_n20255, new_n20256, new_n20257, new_n20258,
    new_n20259, new_n20260, new_n20261, new_n20262, new_n20263, new_n20264,
    new_n20265, new_n20266, new_n20267, new_n20268, new_n20269, new_n20270,
    new_n20271, new_n20272, new_n20273, new_n20274, new_n20275, new_n20276,
    new_n20277, new_n20278, new_n20279, new_n20280, new_n20281, new_n20282,
    new_n20283, new_n20284, new_n20285, new_n20286, new_n20287, new_n20288,
    new_n20289, new_n20290, new_n20291, new_n20292, new_n20293, new_n20294,
    new_n20295, new_n20296, new_n20297, new_n20298, new_n20299, new_n20300,
    new_n20301, new_n20302, new_n20303, new_n20304, new_n20305, new_n20306,
    new_n20307, new_n20308, new_n20309, new_n20310, new_n20311, new_n20312,
    new_n20313, new_n20314, new_n20315, new_n20316, new_n20317, new_n20318,
    new_n20319, new_n20320, new_n20321, new_n20322, new_n20323, new_n20324,
    new_n20325, new_n20326, new_n20327, new_n20328, new_n20329, new_n20330,
    new_n20331, new_n20332, new_n20333, new_n20334, new_n20335, new_n20336,
    new_n20337, new_n20338, new_n20339, new_n20340, new_n20341, new_n20342,
    new_n20343, new_n20344, new_n20345, new_n20346, new_n20347, new_n20348,
    new_n20349, new_n20350, new_n20351, new_n20352, new_n20353, new_n20354,
    new_n20355, new_n20356, new_n20357, new_n20358, new_n20359, new_n20360,
    new_n20361, new_n20362, new_n20363, new_n20364, new_n20365, new_n20366,
    new_n20367, new_n20368, new_n20369, new_n20370, new_n20371, new_n20372,
    new_n20373, new_n20374, new_n20375, new_n20376, new_n20377, new_n20378,
    new_n20379, new_n20380, new_n20381, new_n20382, new_n20383, new_n20384,
    new_n20385, new_n20386, new_n20387, new_n20388, new_n20389, new_n20390,
    new_n20391, new_n20392, new_n20393, new_n20394, new_n20395, new_n20396,
    new_n20397, new_n20398, new_n20399, new_n20400, new_n20401, new_n20402,
    new_n20403, new_n20404, new_n20405, new_n20406, new_n20407, new_n20408,
    new_n20409, new_n20410, new_n20411, new_n20412, new_n20413, new_n20414,
    new_n20415, new_n20416, new_n20417, new_n20418, new_n20419, new_n20420,
    new_n20421, new_n20422, new_n20423, new_n20424, new_n20425, new_n20426,
    new_n20427, new_n20428, new_n20429, new_n20430, new_n20431, new_n20432,
    new_n20433, new_n20434, new_n20435, new_n20436, new_n20437, new_n20438,
    new_n20439, new_n20440, new_n20441, new_n20442, new_n20443, new_n20444,
    new_n20445, new_n20446, new_n20447, new_n20448, new_n20449, new_n20450,
    new_n20451, new_n20452, new_n20453, new_n20454, new_n20455, new_n20456,
    new_n20457, new_n20458, new_n20459, new_n20460, new_n20461, new_n20462,
    new_n20463, new_n20464, new_n20465, new_n20466, new_n20467, new_n20468,
    new_n20469, new_n20470, new_n20471, new_n20472, new_n20473, new_n20474,
    new_n20475, new_n20476, new_n20477, new_n20478, new_n20479, new_n20480,
    new_n20481, new_n20482, new_n20483, new_n20484, new_n20485, new_n20486,
    new_n20487, new_n20488, new_n20489, new_n20490, new_n20491, new_n20492,
    new_n20493, new_n20494, new_n20495, new_n20496, new_n20497, new_n20498,
    new_n20499, new_n20500, new_n20501, new_n20502, new_n20503, new_n20504,
    new_n20505, new_n20506, new_n20507, new_n20508, new_n20509, new_n20510,
    new_n20511, new_n20512, new_n20513, new_n20514, new_n20515, new_n20516,
    new_n20517, new_n20518, new_n20519, new_n20520, new_n20521, new_n20522,
    new_n20523, new_n20524, new_n20525, new_n20526, new_n20527, new_n20528,
    new_n20529, new_n20530, new_n20531, new_n20532, new_n20533, new_n20534,
    new_n20535, new_n20536, new_n20537, new_n20538, new_n20539, new_n20540,
    new_n20541, new_n20542, new_n20543, new_n20544, new_n20545, new_n20546,
    new_n20547, new_n20548, new_n20549, new_n20550, new_n20551, new_n20552,
    new_n20553, new_n20554, new_n20555, new_n20556, new_n20557, new_n20558,
    new_n20559, new_n20560, new_n20561, new_n20562, new_n20563, new_n20564,
    new_n20565, new_n20566, new_n20567, new_n20568, new_n20569, new_n20570,
    new_n20571, new_n20572, new_n20573, new_n20574, new_n20575, new_n20576,
    new_n20577, new_n20578, new_n20579, new_n20580, new_n20581, new_n20582,
    new_n20583, new_n20584, new_n20585, new_n20586, new_n20587, new_n20588,
    new_n20589, new_n20590, new_n20591, new_n20592, new_n20593, new_n20594,
    new_n20595, new_n20596, new_n20597, new_n20598, new_n20599, new_n20600,
    new_n20601, new_n20602, new_n20603, new_n20604, new_n20605, new_n20606,
    new_n20607, new_n20608, new_n20609, new_n20610, new_n20611, new_n20612,
    new_n20613, new_n20614, new_n20615, new_n20616, new_n20617, new_n20618,
    new_n20619, new_n20620, new_n20621, new_n20622, new_n20623, new_n20624,
    new_n20625, new_n20626, new_n20627, new_n20628, new_n20629, new_n20630,
    new_n20631, new_n20632, new_n20633, new_n20634, new_n20635, new_n20636,
    new_n20637, new_n20638, new_n20639, new_n20640, new_n20641, new_n20642,
    new_n20643, new_n20644, new_n20645, new_n20646, new_n20647, new_n20648,
    new_n20649, new_n20650, new_n20651, new_n20652, new_n20653, new_n20654,
    new_n20655, new_n20656, new_n20657, new_n20658, new_n20659, new_n20660,
    new_n20661, new_n20662, new_n20663, new_n20664, new_n20665, new_n20666,
    new_n20667, new_n20668, new_n20669, new_n20670, new_n20671, new_n20672,
    new_n20673, new_n20674, new_n20675, new_n20676, new_n20677, new_n20678,
    new_n20679, new_n20680, new_n20681, new_n20682, new_n20683, new_n20684,
    new_n20685, new_n20686, new_n20687, new_n20688, new_n20689, new_n20690,
    new_n20691, new_n20692, new_n20693, new_n20694, new_n20695, new_n20696,
    new_n20697, new_n20698, new_n20699, new_n20700, new_n20701, new_n20702,
    new_n20703, new_n20704, new_n20705, new_n20706, new_n20707, new_n20708,
    new_n20709, new_n20710, new_n20711, new_n20712, new_n20713, new_n20714,
    new_n20715, new_n20716, new_n20717, new_n20718, new_n20719, new_n20720,
    new_n20721, new_n20722, new_n20723, new_n20724, new_n20725, new_n20726,
    new_n20727, new_n20728, new_n20729, new_n20730, new_n20731, new_n20732,
    new_n20733, new_n20734, new_n20735, new_n20736, new_n20737, new_n20738,
    new_n20739, new_n20740, new_n20741, new_n20742, new_n20743, new_n20744,
    new_n20745, new_n20746, new_n20747, new_n20748, new_n20749, new_n20750,
    new_n20751, new_n20752, new_n20753, new_n20754, new_n20755, new_n20756,
    new_n20757, new_n20758, new_n20759, new_n20760, new_n20761, new_n20762,
    new_n20763, new_n20764, new_n20765, new_n20766, new_n20767, new_n20768,
    new_n20769, new_n20770, new_n20771, new_n20772, new_n20773, new_n20774,
    new_n20775, new_n20776, new_n20777, new_n20778, new_n20779, new_n20780,
    new_n20781, new_n20782, new_n20783, new_n20784, new_n20785, new_n20786,
    new_n20787, new_n20788, new_n20789, new_n20790, new_n20791, new_n20792,
    new_n20793, new_n20794, new_n20795, new_n20796, new_n20797, new_n20798,
    new_n20799, new_n20800, new_n20801, new_n20802, new_n20803, new_n20804,
    new_n20805, new_n20806, new_n20807, new_n20808, new_n20809, new_n20810,
    new_n20811, new_n20812, new_n20813, new_n20814, new_n20815, new_n20816,
    new_n20817, new_n20818, new_n20819, new_n20820, new_n20821, new_n20822,
    new_n20823, new_n20824, new_n20825, new_n20826, new_n20827, new_n20828,
    new_n20829, new_n20830, new_n20831, new_n20832, new_n20833, new_n20834,
    new_n20835, new_n20836, new_n20837, new_n20838, new_n20839, new_n20840,
    new_n20841, new_n20842, new_n20843, new_n20844, new_n20845, new_n20846,
    new_n20847, new_n20848, new_n20849, new_n20850, new_n20851, new_n20852,
    new_n20853, new_n20854, new_n20855, new_n20856, new_n20857, new_n20858,
    new_n20859, new_n20860, new_n20861, new_n20862, new_n20863, new_n20864,
    new_n20865, new_n20866, new_n20867, new_n20868, new_n20869, new_n20870,
    new_n20871, new_n20872, new_n20873, new_n20874, new_n20875, new_n20876,
    new_n20877, new_n20878, new_n20879, new_n20880, new_n20881, new_n20882,
    new_n20883, new_n20884, new_n20885, new_n20886, new_n20887, new_n20888,
    new_n20889, new_n20890, new_n20891, new_n20892, new_n20893, new_n20894,
    new_n20895, new_n20896, new_n20897, new_n20898, new_n20899, new_n20900,
    new_n20901, new_n20902, new_n20903, new_n20904, new_n20905, new_n20906,
    new_n20907, new_n20908, new_n20909, new_n20910, new_n20911, new_n20912,
    new_n20913, new_n20914, new_n20915, new_n20916, new_n20917, new_n20918,
    new_n20919, new_n20920, new_n20921, new_n20922, new_n20923, new_n20924,
    new_n20925, new_n20926, new_n20927, new_n20928, new_n20929, new_n20930,
    new_n20931, new_n20932, new_n20933, new_n20934, new_n20935, new_n20936,
    new_n20937, new_n20938, new_n20939, new_n20940, new_n20941, new_n20942,
    new_n20943, new_n20944, new_n20945, new_n20946, new_n20947, new_n20948,
    new_n20949, new_n20950, new_n20951, new_n20952, new_n20953, new_n20954,
    new_n20955, new_n20956, new_n20957, new_n20958, new_n20959, new_n20960,
    new_n20961, new_n20962, new_n20963, new_n20964, new_n20965, new_n20966,
    new_n20967, new_n20968, new_n20969, new_n20970, new_n20971, new_n20972,
    new_n20973, new_n20974, new_n20975, new_n20976, new_n20977, new_n20978,
    new_n20979, new_n20980, new_n20981, new_n20982, new_n20983, new_n20984,
    new_n20985, new_n20986, new_n20987, new_n20988, new_n20989, new_n20990,
    new_n20991, new_n20992, new_n20993, new_n20994, new_n20995, new_n20996,
    new_n20997, new_n20998, new_n20999, new_n21000, new_n21001, new_n21002,
    new_n21003, new_n21004, new_n21005, new_n21006, new_n21007, new_n21008,
    new_n21009, new_n21010, new_n21011, new_n21012, new_n21013, new_n21014,
    new_n21015, new_n21016, new_n21017, new_n21018, new_n21019, new_n21020,
    new_n21021, new_n21022, new_n21023, new_n21024, new_n21025, new_n21026,
    new_n21027, new_n21028, new_n21029, new_n21030, new_n21031, new_n21032,
    new_n21033, new_n21034, new_n21035, new_n21036, new_n21037, new_n21038,
    new_n21039, new_n21040, new_n21041, new_n21042, new_n21043, new_n21044,
    new_n21045, new_n21046, new_n21047, new_n21048, new_n21049, new_n21050,
    new_n21051, new_n21052, new_n21053, new_n21054, new_n21055, new_n21056,
    new_n21057, new_n21058, new_n21059, new_n21060, new_n21061, new_n21062,
    new_n21063, new_n21064, new_n21065, new_n21066, new_n21067, new_n21068,
    new_n21069, new_n21070, new_n21071, new_n21072, new_n21073, new_n21074,
    new_n21075, new_n21076, new_n21077, new_n21078, new_n21079, new_n21080,
    new_n21081, new_n21082, new_n21083, new_n21084, new_n21085, new_n21086,
    new_n21087, new_n21088, new_n21089, new_n21090, new_n21091, new_n21092,
    new_n21093, new_n21094, new_n21095, new_n21096, new_n21097, new_n21098,
    new_n21099, new_n21100, new_n21101, new_n21102, new_n21103, new_n21104,
    new_n21105, new_n21106, new_n21107, new_n21108, new_n21109, new_n21110,
    new_n21111, new_n21112, new_n21113, new_n21114, new_n21115, new_n21116,
    new_n21117, new_n21118, new_n21119, new_n21120, new_n21121, new_n21122,
    new_n21123, new_n21124, new_n21125, new_n21126, new_n21127, new_n21128,
    new_n21129, new_n21130, new_n21131, new_n21132, new_n21133, new_n21134,
    new_n21135, new_n21136, new_n21137, new_n21138, new_n21139, new_n21140,
    new_n21141, new_n21142, new_n21143, new_n21144, new_n21145, new_n21146,
    new_n21147, new_n21148, new_n21149, new_n21150, new_n21151, new_n21152,
    new_n21153, new_n21154, new_n21155, new_n21156, new_n21157, new_n21158,
    new_n21159, new_n21160, new_n21161, new_n21162, new_n21163, new_n21164,
    new_n21165, new_n21166, new_n21167, new_n21168, new_n21169, new_n21170,
    new_n21171, new_n21172, new_n21173, new_n21174, new_n21175, new_n21176,
    new_n21177, new_n21178, new_n21179, new_n21180, new_n21181, new_n21182,
    new_n21183, new_n21184, new_n21185, new_n21186, new_n21187, new_n21188,
    new_n21189, new_n21190, new_n21191, new_n21192, new_n21193, new_n21194,
    new_n21195, new_n21196, new_n21197, new_n21198, new_n21199, new_n21200,
    new_n21201, new_n21202, new_n21203, new_n21204, new_n21205, new_n21206,
    new_n21207, new_n21208, new_n21209, new_n21210, new_n21211, new_n21212,
    new_n21213, new_n21214, new_n21215, new_n21216, new_n21217, new_n21218,
    new_n21219, new_n21220, new_n21221, new_n21222, new_n21223, new_n21224,
    new_n21225, new_n21226, new_n21227, new_n21228, new_n21229, new_n21230,
    new_n21231, new_n21232, new_n21233, new_n21234, new_n21235, new_n21236,
    new_n21237, new_n21238, new_n21239, new_n21240, new_n21241, new_n21242,
    new_n21243, new_n21244, new_n21245, new_n21246, new_n21247, new_n21248,
    new_n21249, new_n21250, new_n21251, new_n21252, new_n21253, new_n21254,
    new_n21255, new_n21256, new_n21257, new_n21258, new_n21259, new_n21260,
    new_n21261, new_n21262, new_n21263, new_n21264, new_n21265, new_n21266,
    new_n21267, new_n21268, new_n21269, new_n21270, new_n21271, new_n21272,
    new_n21273, new_n21274, new_n21275, new_n21276, new_n21277, new_n21278,
    new_n21279, new_n21280, new_n21281, new_n21282, new_n21283, new_n21284,
    new_n21285, new_n21286, new_n21287, new_n21288, new_n21289, new_n21290,
    new_n21291, new_n21292, new_n21293, new_n21294, new_n21295, new_n21296,
    new_n21297, new_n21298, new_n21299, new_n21300, new_n21301, new_n21302,
    new_n21303, new_n21304, new_n21305, new_n21306, new_n21307, new_n21308,
    new_n21309, new_n21310, new_n21311, new_n21312, new_n21313, new_n21314,
    new_n21315, new_n21316, new_n21317, new_n21318, new_n21319, new_n21320,
    new_n21321, new_n21322, new_n21323, new_n21324, new_n21325, new_n21326,
    new_n21327, new_n21328, new_n21329, new_n21330, new_n21331, new_n21332,
    new_n21333, new_n21334, new_n21335, new_n21336, new_n21337, new_n21338,
    new_n21339, new_n21340, new_n21341, new_n21342, new_n21343, new_n21344,
    new_n21345, new_n21346, new_n21347, new_n21348, new_n21349, new_n21350,
    new_n21351, new_n21352, new_n21353, new_n21354, new_n21355, new_n21356,
    new_n21357, new_n21358, new_n21359, new_n21360, new_n21361, new_n21362,
    new_n21363, new_n21364, new_n21365, new_n21366, new_n21367, new_n21368,
    new_n21369, new_n21370, new_n21371, new_n21372, new_n21373, new_n21374,
    new_n21375, new_n21376, new_n21377, new_n21378, new_n21379, new_n21380,
    new_n21381, new_n21382, new_n21383, new_n21384, new_n21385, new_n21386,
    new_n21387, new_n21388, new_n21389, new_n21390, new_n21391, new_n21392,
    new_n21393, new_n21394, new_n21395, new_n21396, new_n21397, new_n21398,
    new_n21399, new_n21400, new_n21401, new_n21402, new_n21403, new_n21404,
    new_n21405, new_n21406, new_n21407, new_n21408, new_n21409, new_n21410,
    new_n21411, new_n21412, new_n21413, new_n21414, new_n21415, new_n21416,
    new_n21417, new_n21418, new_n21419, new_n21420, new_n21421, new_n21422,
    new_n21423, new_n21424, new_n21425, new_n21426, new_n21427, new_n21428,
    new_n21429, new_n21430, new_n21431, new_n21432, new_n21433, new_n21434,
    new_n21435, new_n21436, new_n21437, new_n21438, new_n21439, new_n21440,
    new_n21441, new_n21442, new_n21443, new_n21444, new_n21445, new_n21446,
    new_n21447, new_n21448, new_n21449, new_n21450, new_n21451, new_n21452,
    new_n21453, new_n21454, new_n21455, new_n21456, new_n21457, new_n21458,
    new_n21459, new_n21460, new_n21461, new_n21462, new_n21463, new_n21464,
    new_n21465, new_n21466, new_n21467, new_n21468, new_n21469, new_n21470,
    new_n21471, new_n21472, new_n21473, new_n21474, new_n21475, new_n21476,
    new_n21477, new_n21478, new_n21479, new_n21480, new_n21481, new_n21482,
    new_n21483, new_n21484, new_n21485, new_n21486, new_n21487, new_n21488,
    new_n21489, new_n21490, new_n21491, new_n21492, new_n21493, new_n21494,
    new_n21495, new_n21496, new_n21497, new_n21498, new_n21499, new_n21500,
    new_n21501, new_n21502, new_n21503, new_n21504, new_n21505, new_n21506,
    new_n21507, new_n21508, new_n21509, new_n21510, new_n21511, new_n21512,
    new_n21513, new_n21514, new_n21515, new_n21516, new_n21517, new_n21518,
    new_n21519, new_n21520, new_n21521, new_n21522, new_n21523, new_n21524,
    new_n21525, new_n21526, new_n21527, new_n21528, new_n21529, new_n21530,
    new_n21531, new_n21532, new_n21533, new_n21534, new_n21535, new_n21536,
    new_n21537, new_n21538, new_n21539, new_n21540, new_n21541, new_n21542,
    new_n21543, new_n21544, new_n21545, new_n21546, new_n21547, new_n21548,
    new_n21549, new_n21550, new_n21551, new_n21552, new_n21553, new_n21554,
    new_n21555, new_n21556, new_n21557, new_n21558, new_n21559, new_n21560,
    new_n21561, new_n21562, new_n21563, new_n21564, new_n21565, new_n21566,
    new_n21567, new_n21568, new_n21569, new_n21570, new_n21571, new_n21572,
    new_n21573, new_n21574, new_n21575, new_n21576, new_n21577, new_n21578,
    new_n21579, new_n21580, new_n21581, new_n21582, new_n21583, new_n21584,
    new_n21585, new_n21586, new_n21587, new_n21588, new_n21589, new_n21590,
    new_n21591, new_n21592, new_n21593, new_n21594, new_n21595, new_n21596,
    new_n21597, new_n21598, new_n21599, new_n21600, new_n21601, new_n21602,
    new_n21603, new_n21604, new_n21605, new_n21606, new_n21607, new_n21608,
    new_n21609, new_n21610, new_n21611, new_n21612, new_n21613, new_n21614,
    new_n21615, new_n21616, new_n21617, new_n21618, new_n21619, new_n21620,
    new_n21621, new_n21622, new_n21623, new_n21624, new_n21625, new_n21626,
    new_n21627, new_n21628, new_n21629, new_n21630, new_n21631, new_n21632,
    new_n21633, new_n21634, new_n21635, new_n21636, new_n21637, new_n21638,
    new_n21639, new_n21640, new_n21641, new_n21642, new_n21643, new_n21644,
    new_n21645, new_n21646, new_n21647, new_n21648, new_n21649, new_n21650,
    new_n21651, new_n21652, new_n21653, new_n21654, new_n21655, new_n21656,
    new_n21657, new_n21658, new_n21659, new_n21660, new_n21661, new_n21662,
    new_n21663, new_n21664, new_n21665, new_n21666, new_n21667, new_n21668,
    new_n21669, new_n21670, new_n21671, new_n21672, new_n21673, new_n21674,
    new_n21675, new_n21676, new_n21677, new_n21678, new_n21679, new_n21680,
    new_n21681, new_n21682, new_n21683, new_n21684, new_n21685, new_n21686,
    new_n21687, new_n21688, new_n21689, new_n21690, new_n21691, new_n21692,
    new_n21693, new_n21694, new_n21695, new_n21696, new_n21697, new_n21698,
    new_n21699, new_n21700, new_n21701, new_n21702, new_n21703, new_n21704,
    new_n21705, new_n21706, new_n21707, new_n21708, new_n21709, new_n21710,
    new_n21711, new_n21712, new_n21713, new_n21714, new_n21715, new_n21716,
    new_n21717, new_n21718, new_n21719, new_n21720, new_n21721, new_n21722,
    new_n21723, new_n21724, new_n21725, new_n21726, new_n21727, new_n21728,
    new_n21729, new_n21730, new_n21731, new_n21732, new_n21733, new_n21734,
    new_n21735, new_n21736, new_n21737, new_n21738, new_n21739, new_n21740,
    new_n21741, new_n21742, new_n21743, new_n21744, new_n21745, new_n21746,
    new_n21747, new_n21748, new_n21749, new_n21750, new_n21751, new_n21752,
    new_n21753, new_n21754, new_n21755, new_n21756, new_n21757, new_n21758,
    new_n21759, new_n21760, new_n21761, new_n21762, new_n21763, new_n21764,
    new_n21765, new_n21766, new_n21767, new_n21768, new_n21769, new_n21770,
    new_n21771, new_n21772, new_n21773, new_n21774, new_n21775, new_n21776,
    new_n21777, new_n21778, new_n21779, new_n21780, new_n21781, new_n21782,
    new_n21783, new_n21784, new_n21785, new_n21786, new_n21787, new_n21788,
    new_n21789, new_n21790, new_n21791, new_n21792, new_n21793, new_n21794,
    new_n21795, new_n21796, new_n21797, new_n21798, new_n21799, new_n21800,
    new_n21801, new_n21802, new_n21803, new_n21804, new_n21805, new_n21806,
    new_n21807, new_n21808, new_n21809, new_n21810, new_n21811, new_n21812,
    new_n21813, new_n21814, new_n21815, new_n21816, new_n21817, new_n21818,
    new_n21819, new_n21820, new_n21821, new_n21822, new_n21823, new_n21824,
    new_n21825, new_n21826, new_n21827, new_n21828, new_n21829, new_n21830,
    new_n21831, new_n21832, new_n21833, new_n21834, new_n21835, new_n21836,
    new_n21837, new_n21838, new_n21839, new_n21840, new_n21841, new_n21842,
    new_n21843, new_n21844, new_n21845, new_n21846, new_n21847, new_n21848,
    new_n21849, new_n21850, new_n21851, new_n21852, new_n21853, new_n21854,
    new_n21855, new_n21856, new_n21857, new_n21858, new_n21859, new_n21860,
    new_n21861, new_n21862, new_n21863, new_n21864, new_n21865, new_n21866,
    new_n21867, new_n21868, new_n21869, new_n21870, new_n21871, new_n21872,
    new_n21873, new_n21874, new_n21875, new_n21876, new_n21877, new_n21878,
    new_n21879, new_n21880, new_n21881, new_n21882, new_n21883, new_n21884,
    new_n21885, new_n21886, new_n21887, new_n21888, new_n21889, new_n21890,
    new_n21891, new_n21892, new_n21893, new_n21894, new_n21895, new_n21896,
    new_n21897, new_n21898, new_n21899, new_n21900, new_n21901, new_n21902,
    new_n21903, new_n21904, new_n21905, new_n21906, new_n21907, new_n21908,
    new_n21909, new_n21910, new_n21911, new_n21912, new_n21913, new_n21914,
    new_n21915, new_n21916, new_n21917, new_n21918, new_n21919, new_n21920,
    new_n21921, new_n21922, new_n21923, new_n21924, new_n21925, new_n21926,
    new_n21927, new_n21928, new_n21929, new_n21930, new_n21931, new_n21932,
    new_n21933, new_n21934, new_n21935, new_n21936, new_n21937, new_n21938,
    new_n21939, new_n21940, new_n21941, new_n21942, new_n21943, new_n21944,
    new_n21945, new_n21946, new_n21947, new_n21948, new_n21949, new_n21950,
    new_n21951, new_n21952, new_n21953, new_n21954, new_n21955, new_n21956,
    new_n21957, new_n21958, new_n21959, new_n21960, new_n21961, new_n21962,
    new_n21963, new_n21964, new_n21965, new_n21966, new_n21967, new_n21968,
    new_n21969, new_n21970, new_n21971, new_n21972, new_n21973, new_n21974,
    new_n21975, new_n21976, new_n21977, new_n21978, new_n21979, new_n21980,
    new_n21981, new_n21982, new_n21983, new_n21984, new_n21985, new_n21986,
    new_n21987, new_n21988, new_n21989, new_n21990, new_n21991, new_n21992,
    new_n21993, new_n21994, new_n21995, new_n21996, new_n21997, new_n21998,
    new_n21999, new_n22000, new_n22001, new_n22002, new_n22003, new_n22004,
    new_n22005, new_n22006, new_n22007, new_n22008, new_n22009, new_n22010,
    new_n22011, new_n22012, new_n22013, new_n22014, new_n22015, new_n22016,
    new_n22017, new_n22018, new_n22019, new_n22020, new_n22021, new_n22022,
    new_n22023, new_n22024, new_n22025, new_n22026, new_n22027, new_n22028,
    new_n22029, new_n22030, new_n22031, new_n22032, new_n22033, new_n22034,
    new_n22035, new_n22036, new_n22037, new_n22038, new_n22039, new_n22040,
    new_n22041, new_n22042, new_n22043, new_n22044, new_n22045, new_n22046,
    new_n22047, new_n22048, new_n22049, new_n22050, new_n22051, new_n22052,
    new_n22053, new_n22054, new_n22055, new_n22056, new_n22057, new_n22058,
    new_n22059, new_n22060, new_n22061, new_n22062, new_n22063, new_n22064,
    new_n22065, new_n22066, new_n22067, new_n22068, new_n22069, new_n22070,
    new_n22071, new_n22072, new_n22073, new_n22074, new_n22075, new_n22076,
    new_n22077, new_n22078, new_n22079, new_n22080, new_n22081, new_n22082,
    new_n22083, new_n22084, new_n22085, new_n22086, new_n22087, new_n22088,
    new_n22089, new_n22090, new_n22091, new_n22092, new_n22093, new_n22094,
    new_n22095, new_n22096, new_n22097, new_n22098, new_n22099, new_n22100,
    new_n22101, new_n22102, new_n22103, new_n22104, new_n22105, new_n22106,
    new_n22107, new_n22108, new_n22109, new_n22110, new_n22111, new_n22112,
    new_n22113, new_n22114, new_n22115, new_n22116, new_n22117, new_n22118,
    new_n22119, new_n22120, new_n22121, new_n22122, new_n22123, new_n22124,
    new_n22125, new_n22126, new_n22127, new_n22128, new_n22129, new_n22130,
    new_n22131, new_n22132, new_n22133, new_n22134, new_n22135, new_n22136,
    new_n22137, new_n22138, new_n22139, new_n22140, new_n22141, new_n22142,
    new_n22143, new_n22144, new_n22145, new_n22146, new_n22147, new_n22148,
    new_n22149, new_n22150, new_n22151, new_n22152, new_n22153, new_n22154,
    new_n22155, new_n22156, new_n22157, new_n22158, new_n22159, new_n22160,
    new_n22161, new_n22162, new_n22163, new_n22164, new_n22165, new_n22166,
    new_n22167, new_n22168, new_n22169, new_n22170, new_n22171, new_n22172,
    new_n22173, new_n22174, new_n22175, new_n22176, new_n22177, new_n22178,
    new_n22179, new_n22180, new_n22181, new_n22182, new_n22183, new_n22184,
    new_n22185, new_n22186, new_n22187, new_n22188, new_n22189, new_n22190,
    new_n22191, new_n22192, new_n22193, new_n22194, new_n22195, new_n22196,
    new_n22197, new_n22198, new_n22199, new_n22200, new_n22201, new_n22202,
    new_n22203, new_n22204, new_n22205, new_n22206, new_n22207, new_n22208,
    new_n22209, new_n22210, new_n22211, new_n22212, new_n22213, new_n22214,
    new_n22215, new_n22216, new_n22217, new_n22218, new_n22219, new_n22220,
    new_n22221, new_n22222, new_n22223, new_n22224, new_n22225, new_n22226,
    new_n22227, new_n22228, new_n22229, new_n22230, new_n22231, new_n22232,
    new_n22233, new_n22234, new_n22235, new_n22236, new_n22237, new_n22238,
    new_n22239, new_n22240, new_n22241, new_n22242, new_n22243, new_n22244,
    new_n22245, new_n22246, new_n22247, new_n22248, new_n22249, new_n22250,
    new_n22251, new_n22252, new_n22253, new_n22254, new_n22255, new_n22256,
    new_n22257, new_n22258, new_n22259, new_n22260, new_n22261, new_n22262,
    new_n22263, new_n22264, new_n22265, new_n22266, new_n22267, new_n22268,
    new_n22269, new_n22270, new_n22271, new_n22272, new_n22273, new_n22274,
    new_n22275, new_n22276, new_n22277, new_n22278, new_n22279, new_n22280,
    new_n22281, new_n22282, new_n22283, new_n22284, new_n22285, new_n22286,
    new_n22287, new_n22288, new_n22289, new_n22290, new_n22291, new_n22292,
    new_n22293, new_n22294, new_n22295, new_n22296, new_n22297, new_n22298,
    new_n22299, new_n22300, new_n22301, new_n22302, new_n22303, new_n22304,
    new_n22305, new_n22306, new_n22307, new_n22308, new_n22309, new_n22310,
    new_n22311, new_n22312, new_n22313, new_n22314, new_n22315, new_n22316,
    new_n22317, new_n22318, new_n22319, new_n22320, new_n22321, new_n22322,
    new_n22323, new_n22324, new_n22325, new_n22326, new_n22327, new_n22328,
    new_n22329, new_n22330, new_n22331, new_n22332, new_n22333, new_n22334,
    new_n22335, new_n22336, new_n22337, new_n22338, new_n22339, new_n22340,
    new_n22341, new_n22342, new_n22343, new_n22344, new_n22345, new_n22346,
    new_n22347, new_n22348, new_n22349, new_n22350, new_n22351, new_n22352,
    new_n22353, new_n22354, new_n22355, new_n22356, new_n22357, new_n22358,
    new_n22359, new_n22360, new_n22361, new_n22362, new_n22363, new_n22364,
    new_n22365, new_n22366, new_n22367, new_n22368, new_n22369, new_n22370,
    new_n22371, new_n22372, new_n22373, new_n22374, new_n22375, new_n22376,
    new_n22377, new_n22378, new_n22379, new_n22380, new_n22381, new_n22382,
    new_n22383, new_n22384, new_n22385, new_n22386, new_n22387, new_n22388,
    new_n22389, new_n22390, new_n22391, new_n22392, new_n22393, new_n22394,
    new_n22395, new_n22396, new_n22397, new_n22398, new_n22399, new_n22400,
    new_n22401, new_n22402, new_n22403, new_n22404, new_n22405, new_n22406,
    new_n22407, new_n22408, new_n22409, new_n22410, new_n22411, new_n22412,
    new_n22413, new_n22414, new_n22415, new_n22416, new_n22417, new_n22418,
    new_n22419, new_n22420, new_n22421, new_n22422, new_n22423, new_n22424,
    new_n22425, new_n22426, new_n22427, new_n22428, new_n22429, new_n22430,
    new_n22431, new_n22432, new_n22433, new_n22434, new_n22435, new_n22436,
    new_n22437, new_n22438, new_n22439, new_n22440, new_n22441, new_n22442,
    new_n22443, new_n22444, new_n22445, new_n22446, new_n22447, new_n22448,
    new_n22449, new_n22450, new_n22451, new_n22452, new_n22453, new_n22454,
    new_n22455, new_n22456, new_n22457, new_n22458, new_n22459, new_n22460,
    new_n22461, new_n22462, new_n22463, new_n22464, new_n22465, new_n22466,
    new_n22467, new_n22468, new_n22469, new_n22470, new_n22471, new_n22472,
    new_n22473, new_n22474, new_n22475, new_n22476, new_n22477, new_n22478,
    new_n22479, new_n22480, new_n22481, new_n22482, new_n22483, new_n22484,
    new_n22485, new_n22486, new_n22487, new_n22488, new_n22489, new_n22490,
    new_n22491, new_n22492, new_n22493, new_n22494, new_n22495, new_n22496,
    new_n22497, new_n22498, new_n22499, new_n22500, new_n22501, new_n22502,
    new_n22503, new_n22504, new_n22505, new_n22506, new_n22507, new_n22508,
    new_n22509, new_n22510, new_n22511, new_n22512, new_n22513, new_n22514,
    new_n22515, new_n22516, new_n22517, new_n22518, new_n22519, new_n22520,
    new_n22521, new_n22522, new_n22523, new_n22524, new_n22525, new_n22526,
    new_n22527, new_n22528, new_n22529, new_n22530, new_n22531, new_n22532,
    new_n22533, new_n22534, new_n22535, new_n22536, new_n22537, new_n22538,
    new_n22539, new_n22540, new_n22541, new_n22542, new_n22543, new_n22544,
    new_n22545, new_n22546, new_n22547, new_n22548, new_n22549, new_n22550,
    new_n22551, new_n22552, new_n22553, new_n22554, new_n22555, new_n22556,
    new_n22557, new_n22558, new_n22559, new_n22560, new_n22561, new_n22562,
    new_n22563, new_n22564, new_n22565, new_n22566, new_n22567, new_n22568,
    new_n22569, new_n22570, new_n22571, new_n22572, new_n22573, new_n22574,
    new_n22575, new_n22576, new_n22577, new_n22578, new_n22579, new_n22580,
    new_n22581, new_n22582, new_n22583, new_n22584, new_n22585, new_n22586,
    new_n22587, new_n22588, new_n22589, new_n22590, new_n22591, new_n22592,
    new_n22593, new_n22594, new_n22595, new_n22596, new_n22597, new_n22598,
    new_n22599, new_n22600, new_n22601, new_n22602, new_n22603, new_n22604,
    new_n22605, new_n22606, new_n22607, new_n22608, new_n22609, new_n22610,
    new_n22611, new_n22612, new_n22613, new_n22614, new_n22615, new_n22616,
    new_n22617, new_n22618, new_n22619, new_n22620, new_n22621, new_n22622,
    new_n22623, new_n22624, new_n22625, new_n22626, new_n22627, new_n22628,
    new_n22629, new_n22630, new_n22631, new_n22632, new_n22633, new_n22634,
    new_n22635, new_n22636, new_n22637, new_n22638, new_n22639, new_n22640,
    new_n22641, new_n22642, new_n22643, new_n22644, new_n22645, new_n22646,
    new_n22647, new_n22648, new_n22649, new_n22650, new_n22651, new_n22652,
    new_n22653, new_n22654, new_n22655, new_n22656, new_n22657, new_n22658,
    new_n22659, new_n22660, new_n22661, new_n22662, new_n22663, new_n22664,
    new_n22665, new_n22666, new_n22667, new_n22668, new_n22669, new_n22670,
    new_n22671, new_n22672, new_n22673, new_n22674, new_n22675, new_n22676,
    new_n22677, new_n22678, new_n22679, new_n22680, new_n22681, new_n22682,
    new_n22683, new_n22684, new_n22685, new_n22686, new_n22687, new_n22688,
    new_n22689, new_n22690, new_n22691, new_n22692, new_n22693, new_n22694,
    new_n22695, new_n22696, new_n22697, new_n22698, new_n22699, new_n22700,
    new_n22701, new_n22702, new_n22703, new_n22704, new_n22705, new_n22706,
    new_n22707, new_n22708, new_n22709, new_n22710, new_n22711, new_n22712,
    new_n22713, new_n22714, new_n22715, new_n22716, new_n22717, new_n22718,
    new_n22719, new_n22720, new_n22721, new_n22722, new_n22723, new_n22724,
    new_n22725, new_n22726, new_n22727, new_n22728, new_n22729, new_n22730,
    new_n22731, new_n22732, new_n22733, new_n22734, new_n22735, new_n22736,
    new_n22737, new_n22738, new_n22739, new_n22740, new_n22741, new_n22742,
    new_n22743, new_n22744, new_n22745, new_n22746, new_n22747, new_n22748,
    new_n22749, new_n22750, new_n22751, new_n22752, new_n22753, new_n22754,
    new_n22755, new_n22756, new_n22757, new_n22758, new_n22759, new_n22760,
    new_n22761, new_n22762, new_n22763, new_n22764, new_n22765, new_n22766,
    new_n22767, new_n22768, new_n22769, new_n22770, new_n22771, new_n22772,
    new_n22773, new_n22774, new_n22775, new_n22776, new_n22777, new_n22778,
    new_n22779, new_n22780, new_n22781, new_n22782, new_n22783, new_n22784,
    new_n22785, new_n22786, new_n22787, new_n22788, new_n22789, new_n22790,
    new_n22791, new_n22792, new_n22793, new_n22794, new_n22795, new_n22796,
    new_n22797, new_n22798, new_n22799, new_n22800, new_n22801, new_n22802,
    new_n22803, new_n22804, new_n22805, new_n22806, new_n22807, new_n22808,
    new_n22809, new_n22810, new_n22811, new_n22812, new_n22813, new_n22814,
    new_n22815, new_n22816, new_n22817, new_n22818, new_n22819, new_n22820,
    new_n22821, new_n22822, new_n22823, new_n22824, new_n22825, new_n22826,
    new_n22827, new_n22828, new_n22829, new_n22830, new_n22831, new_n22832,
    new_n22833, new_n22834, new_n22835, new_n22836, new_n22837, new_n22838,
    new_n22839, new_n22840, new_n22841, new_n22842, new_n22843, new_n22844,
    new_n22845, new_n22846, new_n22847, new_n22848, new_n22849, new_n22850,
    new_n22851, new_n22852, new_n22853, new_n22854, new_n22855, new_n22856,
    new_n22857, new_n22858, new_n22859, new_n22860, new_n22861, new_n22862,
    new_n22863, new_n22864, new_n22865, new_n22866, new_n22867, new_n22868,
    new_n22869, new_n22870, new_n22871, new_n22872, new_n22873, new_n22874,
    new_n22875, new_n22876, new_n22877, new_n22878, new_n22879, new_n22880,
    new_n22881, new_n22882, new_n22883, new_n22884, new_n22885, new_n22886,
    new_n22887, new_n22888, new_n22889, new_n22890, new_n22891, new_n22892,
    new_n22893, new_n22894, new_n22895, new_n22896, new_n22897, new_n22898,
    new_n22899, new_n22900, new_n22901, new_n22902, new_n22903, new_n22904,
    new_n22905, new_n22906, new_n22907, new_n22908, new_n22909, new_n22910,
    new_n22911, new_n22912, new_n22913, new_n22914, new_n22915, new_n22916,
    new_n22917, new_n22918, new_n22919, new_n22920, new_n22921, new_n22922,
    new_n22923, new_n22924, new_n22925, new_n22926, new_n22927, new_n22928,
    new_n22929, new_n22930, new_n22931, new_n22932, new_n22933, new_n22934,
    new_n22935, new_n22936, new_n22937, new_n22938, new_n22939, new_n22940,
    new_n22941, new_n22942, new_n22943, new_n22944, new_n22945, new_n22946,
    new_n22947, new_n22948, new_n22949, new_n22950, new_n22951, new_n22952,
    new_n22953, new_n22954, new_n22955, new_n22956, new_n22957, new_n22958,
    new_n22959, new_n22960, new_n22961, new_n22962, new_n22963, new_n22964,
    new_n22965, new_n22966, new_n22967, new_n22968, new_n22969, new_n22970,
    new_n22971, new_n22972, new_n22973, new_n22974, new_n22975, new_n22976,
    new_n22977, new_n22978, new_n22979, new_n22980, new_n22981, new_n22982,
    new_n22983, new_n22984, new_n22985, new_n22986, new_n22987, new_n22988,
    new_n22989, new_n22990, new_n22991, new_n22992, new_n22993, new_n22994,
    new_n22995, new_n22996, new_n22997, new_n22998, new_n22999, new_n23000,
    new_n23001, new_n23002, new_n23003, new_n23004, new_n23005, new_n23006,
    new_n23007, new_n23008, new_n23009, new_n23010, new_n23011, new_n23012,
    new_n23013, new_n23014, new_n23015, new_n23016, new_n23017, new_n23018,
    new_n23019, new_n23020, new_n23021, new_n23022, new_n23023, new_n23024,
    new_n23025, new_n23026, new_n23027, new_n23028, new_n23029, new_n23030,
    new_n23031, new_n23032, new_n23033, new_n23034, new_n23035, new_n23036,
    new_n23037, new_n23038, new_n23039, new_n23040, new_n23041, new_n23042,
    new_n23043, new_n23044, new_n23045, new_n23046, new_n23047, new_n23048,
    new_n23049, new_n23050, new_n23051, new_n23052, new_n23053, new_n23054,
    new_n23055, new_n23056, new_n23057, new_n23058, new_n23059, new_n23060,
    new_n23061, new_n23062, new_n23063, new_n23064, new_n23065, new_n23066,
    new_n23067, new_n23068, new_n23069, new_n23070, new_n23071, new_n23072,
    new_n23073, new_n23074, new_n23075, new_n23076, new_n23077, new_n23078,
    new_n23079, new_n23080, new_n23081, new_n23082, new_n23083, new_n23084,
    new_n23085, new_n23086, new_n23087, new_n23088, new_n23089, new_n23090,
    new_n23091, new_n23092, new_n23093, new_n23094, new_n23095, new_n23096,
    new_n23097, new_n23098, new_n23099, new_n23100, new_n23101, new_n23102,
    new_n23103, new_n23104, new_n23105, new_n23106, new_n23107, new_n23108,
    new_n23109, new_n23110, new_n23111, new_n23112, new_n23113, new_n23114,
    new_n23115, new_n23116, new_n23117, new_n23118, new_n23119, new_n23120,
    new_n23121, new_n23122, new_n23123, new_n23124, new_n23125, new_n23126,
    new_n23127, new_n23128, new_n23129, new_n23130, new_n23131, new_n23132,
    new_n23133, new_n23134, new_n23135, new_n23136, new_n23137, new_n23138,
    new_n23139, new_n23140, new_n23141, new_n23142, new_n23143, new_n23144,
    new_n23145, new_n23146, new_n23147, new_n23148, new_n23149, new_n23150,
    new_n23151, new_n23152, new_n23153, new_n23154, new_n23155, new_n23156,
    new_n23157, new_n23158, new_n23159, new_n23160, new_n23161, new_n23162,
    new_n23163, new_n23164, new_n23165, new_n23166, new_n23167, new_n23168,
    new_n23169, new_n23170, new_n23171, new_n23172, new_n23173, new_n23174,
    new_n23175, new_n23176, new_n23177, new_n23178, new_n23179, new_n23180,
    new_n23181, new_n23182, new_n23183, new_n23184, new_n23185, new_n23186,
    new_n23187, new_n23188, new_n23189, new_n23190, new_n23191, new_n23192,
    new_n23193, new_n23194, new_n23195, new_n23196, new_n23197, new_n23198,
    new_n23199, new_n23200, new_n23201, new_n23202, new_n23203, new_n23204,
    new_n23205, new_n23206, new_n23207, new_n23208, new_n23209, new_n23210,
    new_n23211, new_n23212, new_n23213, new_n23214, new_n23215, new_n23216,
    new_n23217, new_n23218, new_n23219, new_n23220, new_n23221, new_n23222,
    new_n23223, new_n23224, new_n23225, new_n23226, new_n23227, new_n23228,
    new_n23229, new_n23230, new_n23231, new_n23232, new_n23233, new_n23234,
    new_n23235, new_n23236, new_n23237, new_n23238, new_n23239, new_n23240,
    new_n23241, new_n23242, new_n23243, new_n23244, new_n23245, new_n23246,
    new_n23247, new_n23248, new_n23249, new_n23250, new_n23251, new_n23252,
    new_n23253, new_n23254, new_n23255, new_n23256, new_n23257, new_n23258,
    new_n23259, new_n23260, new_n23261, new_n23262, new_n23263, new_n23264,
    new_n23265, new_n23266, new_n23267, new_n23268, new_n23269, new_n23270,
    new_n23271, new_n23272, new_n23273, new_n23274, new_n23275, new_n23276,
    new_n23277, new_n23278, new_n23279, new_n23280, new_n23281, new_n23282,
    new_n23283, new_n23284, new_n23285, new_n23286, new_n23287, new_n23288,
    new_n23289, new_n23290, new_n23291, new_n23292, new_n23293, new_n23294,
    new_n23295, new_n23296, new_n23297, new_n23298, new_n23299, new_n23300,
    new_n23301, new_n23302, new_n23303, new_n23304, new_n23305, new_n23306,
    new_n23307, new_n23308, new_n23309, new_n23310, new_n23311, new_n23312,
    new_n23313, new_n23314, new_n23315, new_n23316, new_n23317, new_n23318,
    new_n23319, new_n23320, new_n23321, new_n23322, new_n23323, new_n23324,
    new_n23325, new_n23326, new_n23327, new_n23328, new_n23329, new_n23330,
    new_n23331, new_n23332, new_n23333, new_n23334, new_n23335, new_n23336,
    new_n23337, new_n23338, new_n23339, new_n23340, new_n23341, new_n23342,
    new_n23343, new_n23344, new_n23345, new_n23346, new_n23347, new_n23348,
    new_n23349, new_n23350, new_n23351, new_n23352, new_n23353, new_n23354,
    new_n23355, new_n23356, new_n23357, new_n23358, new_n23359, new_n23360,
    new_n23361, new_n23362, new_n23363, new_n23364, new_n23365, new_n23366,
    new_n23367, new_n23368, new_n23369, new_n23370, new_n23371, new_n23372,
    new_n23373, new_n23374, new_n23375, new_n23376, new_n23377, new_n23378,
    new_n23379, new_n23380, new_n23381, new_n23382, new_n23383, new_n23384,
    new_n23385, new_n23386, new_n23387, new_n23388, new_n23389, new_n23390,
    new_n23391, new_n23392, new_n23393, new_n23394, new_n23395, new_n23396,
    new_n23397, new_n23398, new_n23399, new_n23400, new_n23401, new_n23402,
    new_n23403, new_n23404, new_n23405, new_n23406, new_n23407, new_n23408,
    new_n23409, new_n23410, new_n23411, new_n23412, new_n23413, new_n23414,
    new_n23415, new_n23416, new_n23417, new_n23418, new_n23419, new_n23420,
    new_n23421, new_n23422, new_n23423, new_n23424, new_n23425, new_n23426,
    new_n23427, new_n23428, new_n23429, new_n23430, new_n23431, new_n23432,
    new_n23433, new_n23434, new_n23435, new_n23436, new_n23437, new_n23438,
    new_n23439, new_n23440, new_n23441, new_n23442, new_n23443, new_n23444,
    new_n23445, new_n23446, new_n23447, new_n23448, new_n23449, new_n23450,
    new_n23451, new_n23452, new_n23453, new_n23454, new_n23455, new_n23456,
    new_n23457, new_n23458, new_n23459, new_n23460, new_n23461, new_n23462,
    new_n23463, new_n23464, new_n23465, new_n23466, new_n23467, new_n23468,
    new_n23469, new_n23470, new_n23471, new_n23472, new_n23473, new_n23474,
    new_n23475, new_n23476, new_n23477, new_n23478, new_n23479, new_n23480,
    new_n23481, new_n23482, new_n23483, new_n23484, new_n23485, new_n23486,
    new_n23487, new_n23488, new_n23489, new_n23490, new_n23491, new_n23492,
    new_n23493, new_n23494, new_n23495, new_n23496, new_n23497, new_n23498,
    new_n23499, new_n23500, new_n23501, new_n23502, new_n23503, new_n23504,
    new_n23505, new_n23506, new_n23507, new_n23508, new_n23509, new_n23510,
    new_n23511, new_n23512, new_n23513, new_n23514, new_n23515, new_n23516,
    new_n23517, new_n23518, new_n23519, new_n23520, new_n23521, new_n23522,
    new_n23523, new_n23524, new_n23525, new_n23526, new_n23527, new_n23528,
    new_n23529, new_n23530, new_n23531, new_n23532, new_n23533, new_n23534,
    new_n23535, new_n23536, new_n23537, new_n23538, new_n23539, new_n23540,
    new_n23541, new_n23542, new_n23543, new_n23544, new_n23545, new_n23546,
    new_n23547, new_n23548, new_n23549, new_n23550, new_n23551, new_n23552,
    new_n23553, new_n23554, new_n23555, new_n23556, new_n23557, new_n23558,
    new_n23559, new_n23560, new_n23561, new_n23562, new_n23563, new_n23564,
    new_n23565, new_n23566, new_n23567, new_n23568, new_n23569, new_n23570,
    new_n23571, new_n23572, new_n23573, new_n23574, new_n23575, new_n23576,
    new_n23577, new_n23578, new_n23579, new_n23580, new_n23581, new_n23582,
    new_n23583, new_n23584, new_n23585, new_n23586, new_n23587, new_n23588,
    new_n23589, new_n23590, new_n23591, new_n23592, new_n23593, new_n23594,
    new_n23595, new_n23596, new_n23597, new_n23598, new_n23599, new_n23600,
    new_n23601, new_n23602, new_n23603, new_n23604, new_n23605, new_n23606,
    new_n23607, new_n23608, new_n23609, new_n23610, new_n23611, new_n23612,
    new_n23613, new_n23614, new_n23615, new_n23616, new_n23617, new_n23618,
    new_n23619, new_n23620, new_n23621, new_n23622, new_n23623, new_n23624,
    new_n23625, new_n23626, new_n23627, new_n23628, new_n23629, new_n23630,
    new_n23631, new_n23632, new_n23633, new_n23634, new_n23635, new_n23636,
    new_n23637, new_n23638, new_n23639, new_n23640, new_n23641, new_n23642,
    new_n23643, new_n23644, new_n23645, new_n23646, new_n23647, new_n23648,
    new_n23649, new_n23650, new_n23651, new_n23652, new_n23653, new_n23654,
    new_n23655, new_n23656, new_n23657, new_n23658, new_n23659, new_n23660,
    new_n23661, new_n23662, new_n23663, new_n23664, new_n23665, new_n23666,
    new_n23667, new_n23668, new_n23669, new_n23670, new_n23671, new_n23672,
    new_n23673, new_n23674, new_n23675, new_n23676, new_n23677, new_n23678,
    new_n23679, new_n23680, new_n23681, new_n23682, new_n23683, new_n23684,
    new_n23685, new_n23686, new_n23687, new_n23688, new_n23689, new_n23690,
    new_n23691, new_n23692, new_n23693, new_n23694, new_n23695, new_n23696,
    new_n23697, new_n23698, new_n23699, new_n23700, new_n23701, new_n23702,
    new_n23703, new_n23704, new_n23705, new_n23706, new_n23707, new_n23708,
    new_n23709, new_n23710, new_n23711, new_n23712, new_n23713, new_n23714,
    new_n23715, new_n23716, new_n23717, new_n23718, new_n23719, new_n23720,
    new_n23721, new_n23722, new_n23723, new_n23724, new_n23725, new_n23726,
    new_n23727, new_n23728, new_n23729, new_n23730, new_n23731, new_n23732,
    new_n23733, new_n23734, new_n23735, new_n23736, new_n23737, new_n23738,
    new_n23739, new_n23740, new_n23741, new_n23742, new_n23743, new_n23744,
    new_n23745, new_n23746, new_n23747, new_n23748, new_n23749, new_n23750,
    new_n23751, new_n23752, new_n23753, new_n23754, new_n23755, new_n23756,
    new_n23757, new_n23758, new_n23759, new_n23760, new_n23761, new_n23762,
    new_n23763, new_n23764, new_n23765, new_n23766, new_n23767, new_n23768,
    new_n23769, new_n23770, new_n23771, new_n23772, new_n23773, new_n23774,
    new_n23775, new_n23776, new_n23777, new_n23778, new_n23779, new_n23780,
    new_n23781, new_n23782, new_n23783, new_n23784, new_n23785, new_n23786,
    new_n23787, new_n23788, new_n23789, new_n23790, new_n23791, new_n23792,
    new_n23793, new_n23794, new_n23795, new_n23796, new_n23797, new_n23798,
    new_n23799, new_n23800, new_n23801, new_n23802, new_n23803, new_n23804,
    new_n23805, new_n23806, new_n23807, new_n23808, new_n23809, new_n23810,
    new_n23811, new_n23812, new_n23813, new_n23814, new_n23815, new_n23816,
    new_n23817, new_n23818, new_n23819, new_n23820, new_n23821, new_n23822,
    new_n23823, new_n23824, new_n23825, new_n23826, new_n23827, new_n23828,
    new_n23829, new_n23830, new_n23831, new_n23832, new_n23833, new_n23834,
    new_n23835, new_n23836, new_n23837, new_n23838, new_n23839, new_n23840,
    new_n23841, new_n23842, new_n23843, new_n23844, new_n23845, new_n23846,
    new_n23847, new_n23848, new_n23849, new_n23850, new_n23851, new_n23852,
    new_n23853, new_n23854, new_n23855, new_n23856, new_n23857, new_n23858,
    new_n23859, new_n23860, new_n23861, new_n23862, new_n23863, new_n23864,
    new_n23865, new_n23866, new_n23867, new_n23868, new_n23869, new_n23870,
    new_n23871, new_n23872, new_n23873, new_n23874, new_n23875, new_n23876,
    new_n23877, new_n23878, new_n23879, new_n23880, new_n23881, new_n23882,
    new_n23883, new_n23884, new_n23885, new_n23886, new_n23887, new_n23888,
    new_n23889, new_n23890, new_n23891, new_n23892, new_n23893, new_n23894,
    new_n23895, new_n23896, new_n23897, new_n23898, new_n23899, new_n23900,
    new_n23901, new_n23902, new_n23903, new_n23904, new_n23905, new_n23906,
    new_n23907, new_n23908, new_n23909, new_n23910, new_n23911, new_n23912,
    new_n23913, new_n23914, new_n23915, new_n23916, new_n23917, new_n23918,
    new_n23919, new_n23920, new_n23921, new_n23922, new_n23923, new_n23924,
    new_n23925, new_n23926, new_n23927, new_n23928, new_n23929, new_n23930,
    new_n23931, new_n23932, new_n23933, new_n23934, new_n23935, new_n23936,
    new_n23937, new_n23938, new_n23939, new_n23940, new_n23941, new_n23942,
    new_n23943, new_n23944, new_n23945, new_n23946, new_n23947, new_n23948,
    new_n23949, new_n23950, new_n23951, new_n23952, new_n23953, new_n23954,
    new_n23955, new_n23956, new_n23957, new_n23958, new_n23959, new_n23960,
    new_n23961, new_n23962, new_n23963, new_n23964, new_n23965, new_n23966,
    new_n23967, new_n23968, new_n23969, new_n23970, new_n23971, new_n23972,
    new_n23973, new_n23974, new_n23975, new_n23976, new_n23977, new_n23978,
    new_n23979, new_n23980, new_n23981, new_n23982, new_n23983, new_n23984,
    new_n23985, new_n23986, new_n23987, new_n23988, new_n23989, new_n23990,
    new_n23991, new_n23992, new_n23993, new_n23994, new_n23995, new_n23996,
    new_n23997, new_n23998, new_n23999, new_n24000, new_n24001, new_n24002,
    new_n24003, new_n24004, new_n24005, new_n24006, new_n24007, new_n24008,
    new_n24009, new_n24010, new_n24011, new_n24012, new_n24013, new_n24014,
    new_n24015, new_n24016, new_n24017, new_n24018, new_n24019, new_n24020,
    new_n24021, new_n24022, new_n24023, new_n24024, new_n24025, new_n24026,
    new_n24027, new_n24028, new_n24029, new_n24030, new_n24031, new_n24032,
    new_n24033, new_n24034, new_n24035, new_n24036, new_n24037, new_n24038,
    new_n24039, new_n24040, new_n24041, new_n24042, new_n24043, new_n24044,
    new_n24045, new_n24046, new_n24047, new_n24048, new_n24049, new_n24050,
    new_n24051, new_n24052, new_n24053, new_n24054, new_n24055, new_n24056,
    new_n24057, new_n24058, new_n24059, new_n24060, new_n24061, new_n24062,
    new_n24063, new_n24064, new_n24065, new_n24066, new_n24067, new_n24068,
    new_n24069, new_n24070, new_n24071, new_n24072, new_n24073, new_n24074,
    new_n24075, new_n24076, new_n24077, new_n24078, new_n24079, new_n24080,
    new_n24081, new_n24082, new_n24083, new_n24084, new_n24085, new_n24086,
    new_n24087, new_n24088, new_n24089, new_n24090, new_n24091, new_n24092,
    new_n24093, new_n24094, new_n24095, new_n24096, new_n24097, new_n24098,
    new_n24099, new_n24100, new_n24101, new_n24102, new_n24103, new_n24104,
    new_n24105, new_n24106, new_n24107, new_n24108, new_n24109, new_n24110,
    new_n24111, new_n24112, new_n24113, new_n24114, new_n24115, new_n24116,
    new_n24117, new_n24118, new_n24119, new_n24120, new_n24121, new_n24122,
    new_n24123, new_n24124, new_n24125, new_n24126, new_n24127, new_n24128,
    new_n24129, new_n24130, new_n24131, new_n24132, new_n24133, new_n24134,
    new_n24135, new_n24136, new_n24137, new_n24138, new_n24139, new_n24140,
    new_n24141, new_n24142, new_n24143, new_n24144, new_n24145, new_n24146,
    new_n24147, new_n24148, new_n24149, new_n24150, new_n24151, new_n24152,
    new_n24153, new_n24154, new_n24155, new_n24156, new_n24157, new_n24158,
    new_n24159, new_n24160, new_n24161, new_n24162, new_n24163, new_n24164,
    new_n24165, new_n24166, new_n24167, new_n24168, new_n24169, new_n24170,
    new_n24171, new_n24172, new_n24173, new_n24174, new_n24175, new_n24176,
    new_n24177, new_n24178, new_n24179, new_n24180, new_n24181, new_n24182,
    new_n24183, new_n24184, new_n24185, new_n24186, new_n24187, new_n24188,
    new_n24189, new_n24190, new_n24191, new_n24192, new_n24193, new_n24194,
    new_n24195, new_n24196, new_n24197, new_n24198, new_n24199, new_n24200,
    new_n24201, new_n24202, new_n24203, new_n24204, new_n24205, new_n24206,
    new_n24207, new_n24208, new_n24209, new_n24210, new_n24211, new_n24212,
    new_n24213, new_n24214, new_n24215, new_n24216, new_n24217, new_n24218,
    new_n24219, new_n24220, new_n24221, new_n24222, new_n24223, new_n24224,
    new_n24225, new_n24226, new_n24227, new_n24228, new_n24229, new_n24230,
    new_n24231, new_n24232, new_n24233, new_n24234, new_n24235, new_n24236,
    new_n24237, new_n24238, new_n24239, new_n24240, new_n24241, new_n24242,
    new_n24243, new_n24244, new_n24245, new_n24246, new_n24247, new_n24248,
    new_n24249, new_n24250, new_n24251, new_n24252, new_n24253, new_n24254,
    new_n24255, new_n24256, new_n24257, new_n24258, new_n24259, new_n24260,
    new_n24261, new_n24262, new_n24263, new_n24264, new_n24265, new_n24266,
    new_n24267, new_n24268, new_n24269, new_n24270, new_n24271, new_n24272,
    new_n24273, new_n24274, new_n24275, new_n24276, new_n24277, new_n24278,
    new_n24279, new_n24280, new_n24281, new_n24282, new_n24283, new_n24284,
    new_n24285, new_n24286, new_n24287, new_n24288, new_n24289, new_n24290,
    new_n24291, new_n24292, new_n24293, new_n24294, new_n24295, new_n24296,
    new_n24297, new_n24298, new_n24299, new_n24300, new_n24301, new_n24302,
    new_n24303, new_n24304, new_n24305, new_n24306, new_n24307, new_n24308,
    new_n24309, new_n24310, new_n24311, new_n24312, new_n24313, new_n24314,
    new_n24315, new_n24316, new_n24317, new_n24318, new_n24319, new_n24320,
    new_n24321, new_n24322, new_n24323, new_n24324, new_n24325, new_n24326,
    new_n24327, new_n24328, new_n24329, new_n24330, new_n24331, new_n24332,
    new_n24333, new_n24334, new_n24335, new_n24336, new_n24337, new_n24338,
    new_n24339, new_n24340, new_n24341, new_n24342, new_n24343, new_n24344,
    new_n24345, new_n24346, new_n24347, new_n24348, new_n24349, new_n24350,
    new_n24351, new_n24352, new_n24353, new_n24354, new_n24355, new_n24356,
    new_n24357, new_n24358, new_n24359, new_n24360, new_n24361, new_n24362,
    new_n24363, new_n24364, new_n24365, new_n24366, new_n24367, new_n24368,
    new_n24369, new_n24370, new_n24371, new_n24372, new_n24373, new_n24374,
    new_n24375, new_n24376, new_n24377, new_n24378, new_n24379, new_n24380,
    new_n24381, new_n24382, new_n24383, new_n24384, new_n24385, new_n24386,
    new_n24387, new_n24388, new_n24389, new_n24390, new_n24391, new_n24392,
    new_n24393, new_n24394, new_n24395, new_n24396, new_n24397, new_n24398,
    new_n24399, new_n24400, new_n24401, new_n24402, new_n24403, new_n24404,
    new_n24405, new_n24406, new_n24407, new_n24408, new_n24409, new_n24410,
    new_n24411, new_n24412, new_n24413, new_n24414, new_n24415, new_n24416,
    new_n24417, new_n24418, new_n24419, new_n24420, new_n24421, new_n24422,
    new_n24423, new_n24424, new_n24425, new_n24426, new_n24427, new_n24428,
    new_n24429, new_n24430, new_n24431, new_n24432, new_n24433, new_n24434,
    new_n24435, new_n24436, new_n24437, new_n24438, new_n24439, new_n24440,
    new_n24441, new_n24442, new_n24443, new_n24444, new_n24445, new_n24446,
    new_n24447, new_n24448, new_n24449, new_n24450, new_n24451, new_n24452,
    new_n24453, new_n24454, new_n24455, new_n24456, new_n24457, new_n24458,
    new_n24459, new_n24460, new_n24461, new_n24462, new_n24463, new_n24464,
    new_n24465, new_n24466, new_n24467, new_n24468, new_n24469, new_n24470,
    new_n24471, new_n24472, new_n24473, new_n24474, new_n24475, new_n24476,
    new_n24477, new_n24478, new_n24479, new_n24480, new_n24481, new_n24482,
    new_n24483, new_n24484, new_n24485, new_n24486, new_n24487, new_n24488,
    new_n24489, new_n24490, new_n24491, new_n24492, new_n24493, new_n24494,
    new_n24495, new_n24496, new_n24497, new_n24498, new_n24499, new_n24500,
    new_n24501, new_n24502, new_n24503, new_n24504, new_n24505, new_n24506,
    new_n24507, new_n24508, new_n24509, new_n24510, new_n24511, new_n24512,
    new_n24513, new_n24514, new_n24515, new_n24516, new_n24517, new_n24518,
    new_n24519, new_n24520, new_n24521, new_n24522, new_n24523, new_n24524,
    new_n24525, new_n24526, new_n24527, new_n24528, new_n24529, new_n24530,
    new_n24531, new_n24532, new_n24533, new_n24534, new_n24535, new_n24536,
    new_n24537, new_n24538, new_n24539, new_n24540, new_n24541, new_n24542,
    new_n24543, new_n24544, new_n24545, new_n24546, new_n24547, new_n24548,
    new_n24549, new_n24550, new_n24551, new_n24552, new_n24553, new_n24554,
    new_n24555, new_n24556, new_n24557, new_n24558, new_n24559, new_n24560,
    new_n24561, new_n24562, new_n24563, new_n24564, new_n24565, new_n24566,
    new_n24567, new_n24568, new_n24569, new_n24570, new_n24571, new_n24572,
    new_n24573, new_n24574, new_n24575, new_n24576, new_n24577, new_n24578,
    new_n24579, new_n24580, new_n24581, new_n24582, new_n24583, new_n24584,
    new_n24585, new_n24586, new_n24587, new_n24588, new_n24589, new_n24590,
    new_n24591, new_n24592, new_n24593, new_n24594, new_n24595, new_n24596,
    new_n24597, new_n24598, new_n24599, new_n24600, new_n24601, new_n24602,
    new_n24603, new_n24604, new_n24605, new_n24606, new_n24607, new_n24608,
    new_n24609, new_n24610, new_n24611, new_n24612, new_n24613, new_n24614,
    new_n24615, new_n24616, new_n24617, new_n24618, new_n24619, new_n24620,
    new_n24621, new_n24622, new_n24623, new_n24624, new_n24625, new_n24626,
    new_n24627, new_n24628, new_n24629, new_n24630, new_n24631, new_n24632,
    new_n24633, new_n24634, new_n24635, new_n24636, new_n24637, new_n24638,
    new_n24639, new_n24640, new_n24641, new_n24642, new_n24643, new_n24644,
    new_n24645, new_n24646, new_n24647, new_n24648, new_n24649, new_n24650,
    new_n24651, new_n24652, new_n24653, new_n24654, new_n24655, new_n24656,
    new_n24657, new_n24658, new_n24659, new_n24660, new_n24661, new_n24662,
    new_n24663, new_n24664, new_n24665, new_n24666, new_n24667, new_n24668,
    new_n24669, new_n24670, new_n24671, new_n24672, new_n24673, new_n24674,
    new_n24675, new_n24676, new_n24677, new_n24678, new_n24679, new_n24680,
    new_n24681, new_n24682, new_n24683, new_n24684, new_n24685, new_n24686,
    new_n24687, new_n24688, new_n24689, new_n24690, new_n24691, new_n24692,
    new_n24693, new_n24694, new_n24695, new_n24696, new_n24697, new_n24698,
    new_n24699, new_n24700, new_n24701, new_n24702, new_n24703, new_n24704,
    new_n24705, new_n24706, new_n24707, new_n24708, new_n24709, new_n24710,
    new_n24711, new_n24712, new_n24713, new_n24714, new_n24715, new_n24716,
    new_n24717, new_n24718, new_n24719, new_n24720, new_n24721, new_n24722,
    new_n24723, new_n24724, new_n24725, new_n24726, new_n24727, new_n24728,
    new_n24729, new_n24730, new_n24731, new_n24732, new_n24733, new_n24734,
    new_n24735, new_n24736, new_n24737, new_n24738, new_n24739, new_n24740,
    new_n24741, new_n24742, new_n24743, new_n24744, new_n24745, new_n24746,
    new_n24747, new_n24748, new_n24749, new_n24750, new_n24751, new_n24752,
    new_n24753, new_n24754, new_n24755, new_n24756, new_n24757, new_n24758,
    new_n24759, new_n24760, new_n24761, new_n24762, new_n24763, new_n24764,
    new_n24765, new_n24766, new_n24767, new_n24768, new_n24769, new_n24770,
    new_n24771, new_n24772, new_n24773, new_n24774, new_n24775, new_n24776,
    new_n24777, new_n24778, new_n24779, new_n24780, new_n24781, new_n24782,
    new_n24783, new_n24784, new_n24785, new_n24786, new_n24787, new_n24788,
    new_n24789, new_n24790, new_n24791, new_n24792, new_n24793, new_n24794,
    new_n24795, new_n24796, new_n24797, new_n24798, new_n24799, new_n24800,
    new_n24801, new_n24802, new_n24803, new_n24804, new_n24805, new_n24806,
    new_n24807, new_n24808, new_n24809, new_n24810, new_n24811, new_n24812,
    new_n24813, new_n24814, new_n24815, new_n24816, new_n24817, new_n24818,
    new_n24819, new_n24820, new_n24821, new_n24822, new_n24823, new_n24824,
    new_n24825, new_n24826, new_n24827, new_n24828, new_n24829, new_n24830,
    new_n24831, new_n24832, new_n24833, new_n24834, new_n24835, new_n24836,
    new_n24837, new_n24838, new_n24839, new_n24840, new_n24841, new_n24842,
    new_n24843, new_n24844, new_n24845, new_n24846, new_n24847, new_n24848,
    new_n24849, new_n24850, new_n24851, new_n24852, new_n24853, new_n24854,
    new_n24855, new_n24856, new_n24857, new_n24858, new_n24859, new_n24860,
    new_n24861, new_n24862, new_n24863, new_n24864, new_n24865, new_n24866,
    new_n24867, new_n24868, new_n24869, new_n24870, new_n24871, new_n24872,
    new_n24873, new_n24874, new_n24875, new_n24876, new_n24877, new_n24878,
    new_n24879, new_n24880, new_n24881, new_n24882, new_n24883, new_n24884,
    new_n24885, new_n24886, new_n24887, new_n24888, new_n24889, new_n24890,
    new_n24891, new_n24892, new_n24893, new_n24894, new_n24895, new_n24896,
    new_n24897, new_n24898, new_n24899, new_n24900, new_n24901, new_n24902,
    new_n24903, new_n24904, new_n24905, new_n24906, new_n24907, new_n24908,
    new_n24909, new_n24910, new_n24911, new_n24912, new_n24913, new_n24914,
    new_n24915, new_n24916, new_n24917, new_n24918, new_n24919, new_n24920,
    new_n24921, new_n24922, new_n24923, new_n24924, new_n24925, new_n24926,
    new_n24927, new_n24928, new_n24929, new_n24930, new_n24931, new_n24932,
    new_n24933, new_n24934, new_n24935, new_n24936, new_n24937, new_n24938,
    new_n24939, new_n24940, new_n24941, new_n24942, new_n24943, new_n24944,
    new_n24945, new_n24946, new_n24947, new_n24948, new_n24949, new_n24950,
    new_n24951, new_n24952, new_n24953, new_n24954, new_n24955, new_n24956,
    new_n24957, new_n24958, new_n24959, new_n24960, new_n24961, new_n24962,
    new_n24963, new_n24964, new_n24965, new_n24966, new_n24967, new_n24968,
    new_n24969, new_n24970, new_n24971, new_n24972, new_n24973, new_n24974,
    new_n24975, new_n24976, new_n24977, new_n24978, new_n24979, new_n24980,
    new_n24981, new_n24982, new_n24983, new_n24984, new_n24985, new_n24986,
    new_n24987, new_n24988, new_n24989, new_n24990, new_n24991, new_n24992,
    new_n24993, new_n24994, new_n24995, new_n24996, new_n24997, new_n24998,
    new_n24999, new_n25000, new_n25001, new_n25002, new_n25003, new_n25004,
    new_n25005, new_n25006, new_n25007, new_n25008, new_n25009, new_n25010,
    new_n25011, new_n25012, new_n25013, new_n25014, new_n25015, new_n25016,
    new_n25017, new_n25018, new_n25019, new_n25020, new_n25021, new_n25022,
    new_n25023, new_n25024, new_n25025, new_n25026, new_n25027, new_n25028,
    new_n25029, new_n25030, new_n25031, new_n25032, new_n25033, new_n25034,
    new_n25035, new_n25036, new_n25037, new_n25038, new_n25039, new_n25040,
    new_n25041, new_n25042, new_n25043, new_n25044, new_n25045, new_n25046,
    new_n25047, new_n25048, new_n25049, new_n25050, new_n25051, new_n25052,
    new_n25053, new_n25054, new_n25055, new_n25056, new_n25057, new_n25058,
    new_n25059, new_n25060, new_n25061, new_n25062, new_n25063, new_n25064,
    new_n25065, new_n25066, new_n25067, new_n25068, new_n25069, new_n25070,
    new_n25071, new_n25072, new_n25073, new_n25074, new_n25075, new_n25076,
    new_n25077, new_n25078, new_n25079, new_n25080, new_n25081, new_n25082,
    new_n25083, new_n25084, new_n25085, new_n25086, new_n25087, new_n25088,
    new_n25089, new_n25090, new_n25091, new_n25092, new_n25093, new_n25094,
    new_n25095, new_n25096, new_n25097, new_n25098, new_n25099, new_n25100,
    new_n25101, new_n25102, new_n25103, new_n25104, new_n25105, new_n25106,
    new_n25107, new_n25108, new_n25109, new_n25110, new_n25111, new_n25112,
    new_n25113, new_n25114, new_n25115, new_n25116, new_n25117, new_n25118,
    new_n25119, new_n25120, new_n25121, new_n25122, new_n25123, new_n25124,
    new_n25125, new_n25126, new_n25127, new_n25128, new_n25129, new_n25130,
    new_n25131, new_n25132, new_n25133, new_n25134, new_n25135, new_n25136,
    new_n25137, new_n25138, new_n25139, new_n25140, new_n25141, new_n25142,
    new_n25143, new_n25144, new_n25145, new_n25146, new_n25147, new_n25148,
    new_n25149, new_n25150, new_n25151, new_n25152, new_n25153, new_n25154,
    new_n25155, new_n25156, new_n25157, new_n25158, new_n25159, new_n25160,
    new_n25161, new_n25162, new_n25163, new_n25164, new_n25165, new_n25166,
    new_n25167, new_n25168, new_n25169, new_n25170, new_n25171, new_n25172,
    new_n25173, new_n25174, new_n25175, new_n25176, new_n25177, new_n25178,
    new_n25179, new_n25180, new_n25181, new_n25182, new_n25183, new_n25184,
    new_n25185, new_n25186, new_n25187, new_n25188, new_n25189, new_n25190,
    new_n25191, new_n25192, new_n25193, new_n25194, new_n25195, new_n25196,
    new_n25197, new_n25198, new_n25199, new_n25200, new_n25201, new_n25202,
    new_n25203, new_n25204, new_n25205, new_n25206, new_n25207, new_n25208,
    new_n25209, new_n25210, new_n25211, new_n25212, new_n25213, new_n25214,
    new_n25215, new_n25216, new_n25217, new_n25218, new_n25219, new_n25220,
    new_n25221, new_n25222, new_n25223, new_n25224, new_n25225, new_n25226,
    new_n25227, new_n25228, new_n25229, new_n25230, new_n25231, new_n25232,
    new_n25233, new_n25234, new_n25235, new_n25236, new_n25237, new_n25238,
    new_n25239, new_n25240, new_n25241, new_n25242, new_n25243, new_n25244,
    new_n25245, new_n25246, new_n25247, new_n25248, new_n25249, new_n25250,
    new_n25251, new_n25252, new_n25253, new_n25254, new_n25255, new_n25256,
    new_n25257, new_n25258, new_n25259, new_n25260, new_n25261, new_n25262,
    new_n25263, new_n25264, new_n25265, new_n25266, new_n25267, new_n25268,
    new_n25269, new_n25270, new_n25271, new_n25272, new_n25273, new_n25274,
    new_n25275, new_n25276, new_n25277, new_n25278, new_n25279, new_n25280,
    new_n25281, new_n25282, new_n25283, new_n25284, new_n25285, new_n25286,
    new_n25287, new_n25288, new_n25289, new_n25290, new_n25291, new_n25292,
    new_n25293, new_n25294, new_n25295, new_n25296, new_n25297, new_n25298,
    new_n25299, new_n25300, new_n25301, new_n25302, new_n25303, new_n25304,
    new_n25305, new_n25306, new_n25307, new_n25308, new_n25309, new_n25310,
    new_n25311, new_n25312, new_n25313, new_n25314, new_n25315, new_n25316,
    new_n25317, new_n25318, new_n25319, new_n25320, new_n25321, new_n25322,
    new_n25323, new_n25324, new_n25325, new_n25326, new_n25327, new_n25328,
    new_n25329, new_n25330, new_n25331, new_n25332, new_n25333, new_n25334,
    new_n25335, new_n25336, new_n25337, new_n25338, new_n25339, new_n25340,
    new_n25341, new_n25342, new_n25343, new_n25344, new_n25345, new_n25346,
    new_n25347, new_n25348, new_n25349, new_n25350, new_n25351, new_n25352,
    new_n25353, new_n25354, new_n25355, new_n25356, new_n25357, new_n25358,
    new_n25359, new_n25360, new_n25361, new_n25362, new_n25363, new_n25364,
    new_n25365, new_n25366, new_n25367, new_n25368, new_n25369, new_n25370,
    new_n25371, new_n25372, new_n25373, new_n25374, new_n25375, new_n25376,
    new_n25377, new_n25378, new_n25379, new_n25380, new_n25381, new_n25382,
    new_n25383, new_n25384, new_n25385, new_n25386, new_n25387, new_n25388,
    new_n25389, new_n25390, new_n25391, new_n25392, new_n25393, new_n25394,
    new_n25395, new_n25396, new_n25397, new_n25398, new_n25399, new_n25400,
    new_n25401, new_n25402, new_n25403, new_n25404, new_n25405, new_n25406,
    new_n25407, new_n25408, new_n25409, new_n25410, new_n25411, new_n25412,
    new_n25413, new_n25414, new_n25415, new_n25416, new_n25417, new_n25418,
    new_n25419, new_n25420, new_n25421, new_n25422, new_n25423, new_n25424,
    new_n25425, new_n25426, new_n25427, new_n25428, new_n25429, new_n25430,
    new_n25431, new_n25432, new_n25433, new_n25434, new_n25435, new_n25436,
    new_n25437, new_n25438, new_n25439, new_n25440, new_n25441, new_n25442,
    new_n25443, new_n25444, new_n25445, new_n25446, new_n25447, new_n25448,
    new_n25449, new_n25450, new_n25451, new_n25452, new_n25453, new_n25454,
    new_n25455, new_n25456, new_n25457, new_n25458, new_n25459, new_n25460,
    new_n25461, new_n25462, new_n25463, new_n25464, new_n25465, new_n25466,
    new_n25467, new_n25468, new_n25469, new_n25470, new_n25471, new_n25472,
    new_n25473, new_n25474, new_n25475, new_n25476, new_n25477, new_n25478,
    new_n25479, new_n25480, new_n25481, new_n25482, new_n25483, new_n25484,
    new_n25485, new_n25486, new_n25487, new_n25488, new_n25489, new_n25490,
    new_n25491, new_n25492, new_n25493, new_n25494, new_n25495, new_n25496,
    new_n25497, new_n25498, new_n25499, new_n25500, new_n25501, new_n25502,
    new_n25503, new_n25504, new_n25505, new_n25506, new_n25507, new_n25508,
    new_n25509, new_n25510, new_n25511, new_n25512, new_n25513, new_n25514,
    new_n25515, new_n25516, new_n25517, new_n25518, new_n25519, new_n25520,
    new_n25521, new_n25522, new_n25523, new_n25524, new_n25525, new_n25526,
    new_n25527, new_n25528, new_n25529, new_n25530, new_n25531, new_n25532,
    new_n25533, new_n25534, new_n25535, new_n25536, new_n25537, new_n25538,
    new_n25539, new_n25540, new_n25541, new_n25542, new_n25543, new_n25544,
    new_n25545, new_n25546, new_n25547, new_n25548, new_n25549, new_n25550,
    new_n25551, new_n25552, new_n25553, new_n25554, new_n25555, new_n25556,
    new_n25557, new_n25558, new_n25559, new_n25560, new_n25561, new_n25562,
    new_n25563, new_n25564, new_n25565, new_n25566, new_n25567, new_n25568,
    new_n25569, new_n25570, new_n25571, new_n25572, new_n25573, new_n25574,
    new_n25575, new_n25576, new_n25577, new_n25578, new_n25579, new_n25580,
    new_n25581, new_n25582, new_n25583, new_n25584, new_n25585, new_n25586,
    new_n25587, new_n25588, new_n25589, new_n25590, new_n25591, new_n25592,
    new_n25593, new_n25594, new_n25595, new_n25596, new_n25597, new_n25598,
    new_n25599, new_n25600, new_n25601, new_n25602, new_n25603, new_n25604,
    new_n25605, new_n25606, new_n25607, new_n25608, new_n25609, new_n25610,
    new_n25611, new_n25612, new_n25613, new_n25614, new_n25615, new_n25616,
    new_n25617, new_n25618, new_n25619, new_n25620, new_n25621, new_n25622,
    new_n25623, new_n25624, new_n25625, new_n25626, new_n25627, new_n25628,
    new_n25629, new_n25630, new_n25631, new_n25632, new_n25633, new_n25634,
    new_n25635, new_n25636, new_n25637, new_n25638, new_n25639, new_n25640,
    new_n25641, new_n25642, new_n25643, new_n25644, new_n25645, new_n25646,
    new_n25647, new_n25648, new_n25649, new_n25650, new_n25651, new_n25652,
    new_n25653, new_n25654, new_n25655, new_n25656, new_n25657, new_n25658,
    new_n25659, new_n25660, new_n25661, new_n25662, new_n25663, new_n25664,
    new_n25665, new_n25666, new_n25667, new_n25668, new_n25669, new_n25670,
    new_n25671, new_n25672, new_n25673, new_n25674, new_n25675, new_n25676,
    new_n25677, new_n25678, new_n25679, new_n25680, new_n25681, new_n25682,
    new_n25683, new_n25684, new_n25685, new_n25686, new_n25687, new_n25688,
    new_n25689, new_n25690, new_n25691, new_n25692, new_n25693, new_n25694,
    new_n25695, new_n25696, new_n25697, new_n25698, new_n25699, new_n25700,
    new_n25701, new_n25702, new_n25703, new_n25704, new_n25705, new_n25706,
    new_n25707, new_n25708, new_n25709, new_n25710, new_n25711, new_n25712,
    new_n25713, new_n25714, new_n25715, new_n25716, new_n25717, new_n25718,
    new_n25719, new_n25720, new_n25721, new_n25722, new_n25723, new_n25724,
    new_n25725, new_n25726, new_n25727, new_n25728, new_n25729, new_n25730,
    new_n25731, new_n25732, new_n25733, new_n25734, new_n25735, new_n25736,
    new_n25737, new_n25738, new_n25739, new_n25740, new_n25741, new_n25742,
    new_n25743, new_n25744, new_n25745, new_n25746, new_n25747, new_n25748,
    new_n25749, new_n25750, new_n25751, new_n25752, new_n25753, new_n25754,
    new_n25755, new_n25756, new_n25757, new_n25758, new_n25759, new_n25760,
    new_n25761, new_n25762, new_n25763, new_n25764, new_n25765, new_n25766,
    new_n25767, new_n25768, new_n25769, new_n25770, new_n25771, new_n25772,
    new_n25773, new_n25774, new_n25775, new_n25776, new_n25777, new_n25778,
    new_n25779, new_n25780, new_n25781, new_n25782, new_n25783, new_n25784,
    new_n25785, new_n25786, new_n25787, new_n25788, new_n25789, new_n25790,
    new_n25791, new_n25792, new_n25793, new_n25794, new_n25795, new_n25796,
    new_n25797, new_n25798, new_n25799, new_n25800, new_n25801, new_n25802,
    new_n25803, new_n25804, new_n25805, new_n25806, new_n25807, new_n25808,
    new_n25809, new_n25810, new_n25811, new_n25812, new_n25813, new_n25814,
    new_n25815, new_n25816, new_n25817, new_n25818, new_n25819, new_n25820,
    new_n25821, new_n25822, new_n25823, new_n25824, new_n25825, new_n25826,
    new_n25827, new_n25828, new_n25829, new_n25830, new_n25831, new_n25832,
    new_n25833, new_n25834, new_n25835, new_n25836, new_n25837, new_n25838,
    new_n25839, new_n25840, new_n25841, new_n25842, new_n25843, new_n25844,
    new_n25845, new_n25846, new_n25847, new_n25848, new_n25849, new_n25850,
    new_n25851, new_n25852, new_n25853, new_n25854, new_n25855, new_n25856,
    new_n25857, new_n25858, new_n25859, new_n25860, new_n25861, new_n25862,
    new_n25863, new_n25864, new_n25865, new_n25866, new_n25867, new_n25868,
    new_n25869, new_n25870, new_n25871, new_n25872, new_n25873, new_n25874,
    new_n25875, new_n25876, new_n25877, new_n25878, new_n25879, new_n25880,
    new_n25881, new_n25882, new_n25883, new_n25884, new_n25885, new_n25886,
    new_n25887, new_n25888, new_n25889, new_n25890, new_n25891, new_n25892,
    new_n25893, new_n25894, new_n25895, new_n25896, new_n25897, new_n25898,
    new_n25899, new_n25900, new_n25901, new_n25902, new_n25903, new_n25904,
    new_n25905, new_n25906, new_n25907, new_n25908, new_n25909, new_n25910,
    new_n25911, new_n25912, new_n25913, new_n25914, new_n25915, new_n25916,
    new_n25917, new_n25918, new_n25919, new_n25920, new_n25921, new_n25922,
    new_n25923, new_n25924, new_n25925, new_n25926, new_n25927, new_n25928,
    new_n25929, new_n25930, new_n25931, new_n25932, new_n25933, new_n25934,
    new_n25935, new_n25936, new_n25937, new_n25938, new_n25939, new_n25940,
    new_n25941, new_n25942, new_n25943, new_n25944, new_n25945, new_n25946,
    new_n25947, new_n25948, new_n25949, new_n25950, new_n25951, new_n25952,
    new_n25953, new_n25954, new_n25955, new_n25956, new_n25957, new_n25958,
    new_n25959, new_n25960, new_n25961, new_n25962, new_n25963, new_n25964,
    new_n25965, new_n25966, new_n25967, new_n25968, new_n25969, new_n25970,
    new_n25971, new_n25972, new_n25973, new_n25974, new_n25975, new_n25976,
    new_n25977, new_n25978, new_n25979, new_n25980, new_n25981, new_n25982,
    new_n25983, new_n25984, new_n25985, new_n25986, new_n25987, new_n25988,
    new_n25989, new_n25990, new_n25991, new_n25992, new_n25993, new_n25994,
    new_n25995, new_n25996, new_n25997, new_n25998, new_n25999, new_n26000,
    new_n26001, new_n26002, new_n26003, new_n26004, new_n26005, new_n26006,
    new_n26007, new_n26008, new_n26009, new_n26010, new_n26011, new_n26012,
    new_n26013, new_n26014, new_n26015, new_n26016, new_n26017, new_n26018,
    new_n26019, new_n26020, new_n26021, new_n26022, new_n26023, new_n26024,
    new_n26025, new_n26026, new_n26027, new_n26028, new_n26029, new_n26030,
    new_n26031, new_n26032, new_n26033, new_n26034, new_n26035, new_n26036,
    new_n26037, new_n26038, new_n26039, new_n26040, new_n26041, new_n26042,
    new_n26043, new_n26044, new_n26045, new_n26046, new_n26047, new_n26048,
    new_n26049, new_n26050, new_n26051, new_n26052, new_n26053, new_n26054,
    new_n26055, new_n26056, new_n26057, new_n26058, new_n26059, new_n26060,
    new_n26061, new_n26062, new_n26063, new_n26064, new_n26065, new_n26066,
    new_n26067, new_n26068, new_n26069, new_n26070, new_n26071, new_n26072,
    new_n26073, new_n26074, new_n26075, new_n26076, new_n26077, new_n26078,
    new_n26079, new_n26080, new_n26081, new_n26082, new_n26083, new_n26084,
    new_n26085, new_n26086, new_n26087, new_n26088, new_n26089, new_n26090,
    new_n26091, new_n26092, new_n26093, new_n26094, new_n26095, new_n26096,
    new_n26097, new_n26098, new_n26099, new_n26100, new_n26101, new_n26102,
    new_n26103, new_n26104, new_n26105, new_n26106, new_n26107, new_n26108,
    new_n26109, new_n26110, new_n26111, new_n26112, new_n26113, new_n26114,
    new_n26115, new_n26116, new_n26117, new_n26118, new_n26119, new_n26120,
    new_n26121, new_n26122, new_n26123, new_n26124, new_n26125, new_n26126,
    new_n26127, new_n26128, new_n26129, new_n26130, new_n26131, new_n26132,
    new_n26133, new_n26134, new_n26135, new_n26136, new_n26137, new_n26138,
    new_n26139, new_n26140, new_n26141, new_n26142, new_n26143, new_n26144,
    new_n26145, new_n26146, new_n26147, new_n26148, new_n26149, new_n26150,
    new_n26151, new_n26152, new_n26153, new_n26154, new_n26155, new_n26156,
    new_n26157, new_n26158, new_n26159, new_n26160, new_n26161, new_n26162,
    new_n26163, new_n26164, new_n26165, new_n26166, new_n26167, new_n26168,
    new_n26169, new_n26170, new_n26171, new_n26172, new_n26173, new_n26174,
    new_n26175, new_n26176, new_n26177, new_n26178, new_n26179, new_n26180,
    new_n26181, new_n26182, new_n26183, new_n26184, new_n26185, new_n26186,
    new_n26187, new_n26188, new_n26189, new_n26190, new_n26191, new_n26192,
    new_n26193, new_n26194, new_n26195, new_n26196, new_n26197, new_n26198,
    new_n26199, new_n26200, new_n26201, new_n26202, new_n26203, new_n26204,
    new_n26205, new_n26206, new_n26207, new_n26208, new_n26209, new_n26210,
    new_n26211, new_n26212, new_n26213, new_n26214, new_n26215, new_n26216,
    new_n26217, new_n26218, new_n26219, new_n26220, new_n26221, new_n26222,
    new_n26223, new_n26224, new_n26225, new_n26226, new_n26227, new_n26228,
    new_n26229, new_n26230, new_n26231, new_n26232, new_n26233, new_n26234,
    new_n26235, new_n26236, new_n26237, new_n26238, new_n26239, new_n26240,
    new_n26241, new_n26242, new_n26243, new_n26244, new_n26245, new_n26246,
    new_n26247, new_n26248, new_n26249, new_n26250, new_n26251, new_n26252,
    new_n26253, new_n26254, new_n26255, new_n26256, new_n26257, new_n26258,
    new_n26259, new_n26260, new_n26261, new_n26262, new_n26263, new_n26264,
    new_n26265, new_n26266, new_n26267, new_n26268, new_n26269, new_n26270,
    new_n26271, new_n26272, new_n26273, new_n26274, new_n26275, new_n26276,
    new_n26277, new_n26278, new_n26279, new_n26280, new_n26281, new_n26282,
    new_n26283, new_n26284, new_n26285, new_n26286, new_n26287, new_n26288,
    new_n26289, new_n26290, new_n26291, new_n26292, new_n26293, new_n26294,
    new_n26295, new_n26296, new_n26297, new_n26298, new_n26299, new_n26300,
    new_n26301, new_n26302, new_n26303, new_n26304, new_n26305, new_n26306,
    new_n26307, new_n26308, new_n26309, new_n26310, new_n26311, new_n26312,
    new_n26313, new_n26314, new_n26315, new_n26316, new_n26317, new_n26318,
    new_n26319, new_n26320, new_n26321, new_n26322, new_n26323, new_n26324,
    new_n26325, new_n26326, new_n26327, new_n26328, new_n26329, new_n26330,
    new_n26331, new_n26332, new_n26333, new_n26334, new_n26335, new_n26336,
    new_n26337, new_n26338, new_n26339, new_n26340, new_n26341, new_n26342,
    new_n26343, new_n26344, new_n26345, new_n26346, new_n26347, new_n26348,
    new_n26349, new_n26350, new_n26351, new_n26352, new_n26353, new_n26354,
    new_n26355, new_n26356, new_n26357, new_n26358, new_n26359, new_n26360,
    new_n26361, new_n26362, new_n26363, new_n26364, new_n26365, new_n26366,
    new_n26367, new_n26368, new_n26369, new_n26370, new_n26371, new_n26372,
    new_n26373, new_n26374, new_n26375, new_n26376, new_n26377, new_n26378,
    new_n26379, new_n26380, new_n26381, new_n26382, new_n26383, new_n26384,
    new_n26385, new_n26386, new_n26387, new_n26388, new_n26389, new_n26390,
    new_n26391, new_n26392, new_n26393, new_n26394, new_n26395, new_n26396,
    new_n26397, new_n26398, new_n26399, new_n26400, new_n26401, new_n26402,
    new_n26403, new_n26404, new_n26405, new_n26406, new_n26407, new_n26408,
    new_n26409, new_n26410, new_n26411, new_n26412, new_n26413, new_n26414,
    new_n26415, new_n26416, new_n26417, new_n26418, new_n26419, new_n26420,
    new_n26421, new_n26422, new_n26423, new_n26424, new_n26425, new_n26426,
    new_n26427, new_n26428, new_n26429, new_n26430, new_n26431, new_n26432,
    new_n26433, new_n26434, new_n26435, new_n26436, new_n26437, new_n26438,
    new_n26439, new_n26440, new_n26441, new_n26442, new_n26443, new_n26444,
    new_n26445, new_n26446, new_n26447, new_n26448, new_n26449, new_n26450,
    new_n26451, new_n26452, new_n26453, new_n26454, new_n26455, new_n26456,
    new_n26457, new_n26458, new_n26459, new_n26460, new_n26461, new_n26462,
    new_n26463, new_n26464, new_n26465, new_n26466, new_n26467, new_n26468,
    new_n26469, new_n26470, new_n26471, new_n26472, new_n26473, new_n26474,
    new_n26475, new_n26476, new_n26477, new_n26478, new_n26479, new_n26480,
    new_n26481, new_n26482, new_n26483, new_n26484, new_n26485, new_n26486,
    new_n26487, new_n26488, new_n26489, new_n26490, new_n26491, new_n26492,
    new_n26493, new_n26494, new_n26495, new_n26496, new_n26497, new_n26498,
    new_n26499, new_n26500, new_n26501, new_n26502, new_n26503, new_n26504,
    new_n26505, new_n26506, new_n26507, new_n26508, new_n26509, new_n26510,
    new_n26511, new_n26512, new_n26513, new_n26514, new_n26515, new_n26516,
    new_n26517, new_n26518, new_n26519, new_n26520, new_n26521, new_n26522,
    new_n26523, new_n26524, new_n26525, new_n26526, new_n26527, new_n26528,
    new_n26529, new_n26530, new_n26531, new_n26532, new_n26533, new_n26534,
    new_n26535, new_n26536, new_n26537, new_n26538, new_n26539, new_n26540,
    new_n26541, new_n26542, new_n26543, new_n26544, new_n26545, new_n26546,
    new_n26547, new_n26548, new_n26549, new_n26550, new_n26551, new_n26552,
    new_n26553, new_n26554, new_n26555, new_n26556, new_n26557, new_n26558,
    new_n26559, new_n26560, new_n26561, new_n26562, new_n26563, new_n26564,
    new_n26565, new_n26566, new_n26567, new_n26568, new_n26569, new_n26570,
    new_n26571, new_n26572, new_n26573, new_n26574, new_n26575, new_n26576,
    new_n26577, new_n26578, new_n26579, new_n26580, new_n26581, new_n26582,
    new_n26583, new_n26584, new_n26585, new_n26586, new_n26587, new_n26588,
    new_n26589, new_n26590, new_n26591, new_n26592, new_n26593, new_n26594,
    new_n26595, new_n26596, new_n26597, new_n26598, new_n26599, new_n26600,
    new_n26601, new_n26602, new_n26603, new_n26604, new_n26605, new_n26606,
    new_n26607, new_n26608, new_n26609, new_n26610, new_n26611, new_n26612,
    new_n26613, new_n26614, new_n26615, new_n26616, new_n26617, new_n26618,
    new_n26619, new_n26620, new_n26621, new_n26622, new_n26623, new_n26624,
    new_n26625, new_n26626, new_n26627, new_n26628, new_n26629, new_n26630,
    new_n26631, new_n26632, new_n26633, new_n26634, new_n26635, new_n26636,
    new_n26637, new_n26638, new_n26639, new_n26640, new_n26641, new_n26642,
    new_n26643, new_n26644, new_n26645, new_n26646, new_n26647, new_n26648,
    new_n26649, new_n26650, new_n26651, new_n26652, new_n26653, new_n26654,
    new_n26655, new_n26656, new_n26657, new_n26658, new_n26659, new_n26660,
    new_n26661, new_n26662, new_n26663, new_n26664, new_n26665, new_n26666,
    new_n26667, new_n26668, new_n26669, new_n26670, new_n26671, new_n26672,
    new_n26673, new_n26674, new_n26675, new_n26676, new_n26677, new_n26678,
    new_n26679, new_n26680, new_n26681, new_n26682, new_n26683, new_n26684,
    new_n26685, new_n26686, new_n26687, new_n26688, new_n26689, new_n26690,
    new_n26691, new_n26692, new_n26693, new_n26694, new_n26695, new_n26696,
    new_n26697, new_n26698, new_n26699, new_n26700, new_n26701, new_n26702,
    new_n26703, new_n26704, new_n26705, new_n26706, new_n26707, new_n26708,
    new_n26709, new_n26710, new_n26711, new_n26712, new_n26713, new_n26714,
    new_n26715, new_n26716, new_n26717, new_n26718, new_n26719, new_n26720,
    new_n26721, new_n26722, new_n26723, new_n26724, new_n26725, new_n26726,
    new_n26727, new_n26728, new_n26729, new_n26730, new_n26731, new_n26732,
    new_n26733, new_n26734, new_n26735, new_n26736, new_n26737, new_n26738,
    new_n26739, new_n26740, new_n26741, new_n26742, new_n26743, new_n26744,
    new_n26745, new_n26746, new_n26747, new_n26748, new_n26749, new_n26750,
    new_n26751, new_n26752, new_n26753, new_n26754, new_n26755, new_n26756,
    new_n26757, new_n26758, new_n26759, new_n26760, new_n26761, new_n26762,
    new_n26763, new_n26764, new_n26765, new_n26766, new_n26767, new_n26768,
    new_n26769, new_n26770, new_n26771, new_n26772, new_n26773, new_n26774,
    new_n26775, new_n26776, new_n26777, new_n26778, new_n26779, new_n26780,
    new_n26781, new_n26782, new_n26783, new_n26784, new_n26785, new_n26786,
    new_n26787, new_n26788, new_n26789, new_n26790, new_n26791, new_n26792,
    new_n26793, new_n26794, new_n26795, new_n26796, new_n26797, new_n26798,
    new_n26799, new_n26800, new_n26801, new_n26802, new_n26803, new_n26804,
    new_n26805, new_n26806, new_n26807, new_n26808, new_n26809, new_n26810,
    new_n26811, new_n26812, new_n26813, new_n26814, new_n26815, new_n26816,
    new_n26817, new_n26818, new_n26819, new_n26820, new_n26821, new_n26822,
    new_n26823, new_n26824, new_n26825, new_n26826, new_n26827, new_n26828,
    new_n26829, new_n26830, new_n26831, new_n26832, new_n26833, new_n26834,
    new_n26835, new_n26836, new_n26837, new_n26838, new_n26839, new_n26840,
    new_n26841, new_n26842, new_n26843, new_n26844, new_n26845, new_n26846,
    new_n26847, new_n26848, new_n26849, new_n26850, new_n26851, new_n26852,
    new_n26853, new_n26854, new_n26855, new_n26856, new_n26857, new_n26858,
    new_n26859, new_n26860, new_n26861, new_n26862, new_n26863, new_n26864,
    new_n26865, new_n26866, new_n26867, new_n26868, new_n26869, new_n26870,
    new_n26871, new_n26872, new_n26873, new_n26874, new_n26875, new_n26876,
    new_n26877, new_n26878, new_n26879, new_n26880, new_n26881, new_n26882,
    new_n26883, new_n26884, new_n26885, new_n26886, new_n26887, new_n26888,
    new_n26889, new_n26890, new_n26891, new_n26892, new_n26893, new_n26894,
    new_n26895, new_n26896, new_n26897, new_n26898, new_n26899, new_n26900,
    new_n26901, new_n26902, new_n26903, new_n26904, new_n26905, new_n26906,
    new_n26907, new_n26908, new_n26909, new_n26910, new_n26911, new_n26912,
    new_n26913, new_n26914, new_n26915, new_n26916, new_n26917, new_n26918,
    new_n26919, new_n26920, new_n26921, new_n26922, new_n26923, new_n26924,
    new_n26925, new_n26926, new_n26927, new_n26928, new_n26929, new_n26930,
    new_n26931, new_n26932, new_n26933, new_n26934, new_n26935, new_n26936,
    new_n26937, new_n26938, new_n26939, new_n26940, new_n26941, new_n26942,
    new_n26943, new_n26944, new_n26945, new_n26946, new_n26947, new_n26948,
    new_n26949, new_n26950, new_n26951, new_n26952, new_n26953, new_n26954,
    new_n26955, new_n26956, new_n26957, new_n26958, new_n26959, new_n26960,
    new_n26961, new_n26962, new_n26963, new_n26964, new_n26965, new_n26966,
    new_n26967, new_n26968, new_n26969, new_n26970, new_n26971, new_n26972,
    new_n26973, new_n26974, new_n26975, new_n26976, new_n26977, new_n26978,
    new_n26979, new_n26980, new_n26981, new_n26982, new_n26983, new_n26984,
    new_n26985, new_n26986, new_n26987, new_n26988, new_n26989, new_n26990,
    new_n26991, new_n26992, new_n26993, new_n26994, new_n26995, new_n26996,
    new_n26997, new_n26998, new_n26999, new_n27000, new_n27001, new_n27002,
    new_n27003, new_n27004, new_n27005, new_n27006, new_n27007, new_n27008,
    new_n27009, new_n27010, new_n27011, new_n27012, new_n27013, new_n27014,
    new_n27015, new_n27016, new_n27017, new_n27018, new_n27019, new_n27020,
    new_n27021, new_n27022, new_n27023, new_n27024, new_n27025, new_n27026,
    new_n27027, new_n27028, new_n27029, new_n27030, new_n27031, new_n27032,
    new_n27033, new_n27034, new_n27035, new_n27036, new_n27037, new_n27038,
    new_n27039, new_n27040, new_n27041, new_n27042, new_n27043, new_n27044,
    new_n27045, new_n27046, new_n27047, new_n27048, new_n27049, new_n27050,
    new_n27051, new_n27052, new_n27053, new_n27054, new_n27055, new_n27056,
    new_n27057, new_n27058, new_n27059, new_n27060, new_n27061, new_n27062,
    new_n27063, new_n27064, new_n27065, new_n27066, new_n27067, new_n27068,
    new_n27069, new_n27070, new_n27071, new_n27072, new_n27073, new_n27074,
    new_n27075, new_n27076, new_n27077, new_n27078, new_n27079, new_n27080,
    new_n27081, new_n27082, new_n27083, new_n27084, new_n27085, new_n27086,
    new_n27087, new_n27088, new_n27089, new_n27090, new_n27091, new_n27092,
    new_n27093, new_n27094, new_n27095, new_n27096, new_n27097, new_n27098,
    new_n27099, new_n27100, new_n27101, new_n27102, new_n27103, new_n27104,
    new_n27105, new_n27106, new_n27107, new_n27108, new_n27109, new_n27110,
    new_n27111, new_n27112, new_n27113, new_n27114, new_n27115, new_n27116,
    new_n27117, new_n27118, new_n27119, new_n27120, new_n27121, new_n27122,
    new_n27123, new_n27124, new_n27125, new_n27126, new_n27127, new_n27128,
    new_n27129, new_n27130, new_n27131, new_n27132, new_n27133, new_n27134,
    new_n27135, new_n27136, new_n27137, new_n27138, new_n27139, new_n27140,
    new_n27141, new_n27142, new_n27143, new_n27144, new_n27145, new_n27146,
    new_n27147, new_n27148, new_n27149, new_n27150, new_n27151, new_n27152,
    new_n27153, new_n27154, new_n27155, new_n27156, new_n27157, new_n27158,
    new_n27159, new_n27160, new_n27161, new_n27162, new_n27163, new_n27164,
    new_n27165, new_n27166, new_n27167, new_n27168, new_n27169, new_n27170,
    new_n27171, new_n27172, new_n27173, new_n27174, new_n27175, new_n27176,
    new_n27177, new_n27178, new_n27179, new_n27180, new_n27181, new_n27182,
    new_n27183, new_n27184, new_n27185, new_n27186, new_n27187, new_n27188,
    new_n27189, new_n27190, new_n27191, new_n27192, new_n27193, new_n27194,
    new_n27195, new_n27196, new_n27197, new_n27198, new_n27199, new_n27200,
    new_n27201, new_n27202, new_n27203, new_n27204, new_n27205, new_n27206,
    new_n27207, new_n27208, new_n27209, new_n27210, new_n27211, new_n27212,
    new_n27213, new_n27214, new_n27215, new_n27216, new_n27217, new_n27218,
    new_n27219, new_n27220, new_n27221, new_n27222, new_n27223, new_n27224,
    new_n27225, new_n27226, new_n27227, new_n27228, new_n27229, new_n27230,
    new_n27231, new_n27232, new_n27233, new_n27234, new_n27235, new_n27236,
    new_n27237, new_n27238, new_n27239, new_n27240, new_n27241, new_n27242,
    new_n27243, new_n27244, new_n27245, new_n27246, new_n27247, new_n27248,
    new_n27249, new_n27250, new_n27251, new_n27252, new_n27253, new_n27254,
    new_n27255, new_n27256, new_n27257, new_n27258, new_n27259, new_n27260,
    new_n27261, new_n27262, new_n27263, new_n27264, new_n27265, new_n27266,
    new_n27267, new_n27268, new_n27269, new_n27270, new_n27271, new_n27272,
    new_n27273, new_n27274, new_n27275, new_n27276, new_n27277, new_n27278,
    new_n27279, new_n27280, new_n27281, new_n27282, new_n27283, new_n27284,
    new_n27285, new_n27286, new_n27287, new_n27288, new_n27289, new_n27290,
    new_n27291, new_n27292, new_n27293, new_n27294, new_n27295, new_n27296,
    new_n27297, new_n27298, new_n27299, new_n27300, new_n27301, new_n27302,
    new_n27303, new_n27304, new_n27305, new_n27306, new_n27307, new_n27308,
    new_n27309, new_n27310, new_n27311, new_n27312, new_n27313, new_n27314,
    new_n27315, new_n27316, new_n27317, new_n27318, new_n27319, new_n27320,
    new_n27321, new_n27322, new_n27323, new_n27324, new_n27325, new_n27326,
    new_n27327, new_n27328, new_n27329, new_n27330, new_n27331, new_n27332,
    new_n27333, new_n27334, new_n27335, new_n27336, new_n27337, new_n27338,
    new_n27339, new_n27340, new_n27341, new_n27342, new_n27343, new_n27344,
    new_n27345, new_n27346, new_n27347, new_n27348, new_n27349, new_n27350,
    new_n27351, new_n27352, new_n27353, new_n27354, new_n27355, new_n27356,
    new_n27357, new_n27358, new_n27359, new_n27360, new_n27361, new_n27362,
    new_n27363, new_n27364, new_n27365, new_n27366, new_n27367, new_n27368,
    new_n27369, new_n27370, new_n27371, new_n27372, new_n27373, new_n27374,
    new_n27375, new_n27376, new_n27377, new_n27378, new_n27379, new_n27380,
    new_n27381, new_n27382, new_n27383, new_n27384, new_n27385, new_n27386,
    new_n27387, new_n27388, new_n27389, new_n27390, new_n27391, new_n27392,
    new_n27393, new_n27394, new_n27395, new_n27396, new_n27397, new_n27398,
    new_n27399, new_n27400, new_n27401, new_n27402, new_n27403, new_n27404,
    new_n27405, new_n27406, new_n27407, new_n27408, new_n27409, new_n27410,
    new_n27411, new_n27412, new_n27413, new_n27414, new_n27415, new_n27416,
    new_n27417, new_n27418, new_n27419, new_n27420, new_n27421, new_n27422,
    new_n27423, new_n27424, new_n27425, new_n27426, new_n27427, new_n27428,
    new_n27429, new_n27430, new_n27431, new_n27432, new_n27433, new_n27434,
    new_n27435, new_n27436, new_n27437, new_n27438, new_n27439, new_n27440,
    new_n27441, new_n27442, new_n27443, new_n27444, new_n27445, new_n27446,
    new_n27447, new_n27448, new_n27449, new_n27450, new_n27451, new_n27452,
    new_n27453, new_n27454, new_n27455, new_n27456, new_n27457, new_n27458,
    new_n27459, new_n27460, new_n27461, new_n27462, new_n27463, new_n27464,
    new_n27465, new_n27466, new_n27467, new_n27468, new_n27469, new_n27470,
    new_n27471, new_n27472, new_n27473, new_n27474, new_n27475, new_n27476,
    new_n27477, new_n27478, new_n27479, new_n27480, new_n27481, new_n27482,
    new_n27483, new_n27484, new_n27485, new_n27486, new_n27487, new_n27488,
    new_n27489, new_n27490, new_n27491, new_n27492, new_n27493, new_n27494,
    new_n27495, new_n27496, new_n27497, new_n27498, new_n27499, new_n27500,
    new_n27501, new_n27502, new_n27503, new_n27504, new_n27505, new_n27506,
    new_n27507, new_n27508, new_n27509, new_n27510, new_n27511, new_n27512,
    new_n27513, new_n27514, new_n27515, new_n27516, new_n27517, new_n27518,
    new_n27519, new_n27520, new_n27521, new_n27522, new_n27523, new_n27524,
    new_n27525, new_n27526, new_n27527, new_n27528, new_n27529, new_n27530,
    new_n27531, new_n27532, new_n27533, new_n27534, new_n27535, new_n27536,
    new_n27537, new_n27538, new_n27539, new_n27540, new_n27541, new_n27542,
    new_n27543, new_n27544, new_n27545, new_n27546, new_n27547, new_n27548,
    new_n27549, new_n27550, new_n27551, new_n27552, new_n27553, new_n27554,
    new_n27555, new_n27556, new_n27557, new_n27558, new_n27559, new_n27560,
    new_n27561, new_n27562, new_n27563, new_n27564, new_n27565, new_n27566,
    new_n27567, new_n27568, new_n27569, new_n27570, new_n27571, new_n27572,
    new_n27573, new_n27574, new_n27575, new_n27576, new_n27577, new_n27578,
    new_n27579, new_n27580, new_n27581, new_n27582, new_n27583, new_n27584,
    new_n27585, new_n27586, new_n27587, new_n27588, new_n27589, new_n27590,
    new_n27591, new_n27592, new_n27593, new_n27594, new_n27595, new_n27596,
    new_n27597, new_n27598, new_n27599, new_n27600, new_n27601, new_n27602,
    new_n27603, new_n27604, new_n27605, new_n27606, new_n27607, new_n27608,
    new_n27609, new_n27610, new_n27611, new_n27612, new_n27613, new_n27614,
    new_n27615, new_n27616, new_n27617, new_n27618, new_n27619, new_n27620,
    new_n27621, new_n27622, new_n27623, new_n27624, new_n27625, new_n27626,
    new_n27627, new_n27628, new_n27629, new_n27630, new_n27631, new_n27632,
    new_n27633, new_n27634, new_n27635, new_n27636, new_n27637, new_n27638,
    new_n27639, new_n27640, new_n27641, new_n27642, new_n27643, new_n27644,
    new_n27645, new_n27646, new_n27647, new_n27648, new_n27649, new_n27650,
    new_n27651, new_n27652, new_n27653, new_n27654, new_n27655, new_n27656,
    new_n27657, new_n27658, new_n27659, new_n27660, new_n27661, new_n27662,
    new_n27663, new_n27664, new_n27665, new_n27666, new_n27667, new_n27668,
    new_n27669, new_n27670, new_n27671, new_n27672, new_n27673, new_n27674,
    new_n27675, new_n27676, new_n27677, new_n27678, new_n27679, new_n27680,
    new_n27681, new_n27682, new_n27683, new_n27684, new_n27685, new_n27686,
    new_n27687, new_n27688, new_n27689, new_n27690, new_n27691, new_n27692,
    new_n27693, new_n27694, new_n27695, new_n27696, new_n27697, new_n27698,
    new_n27699, new_n27700, new_n27701, new_n27702, new_n27703, new_n27704,
    new_n27705, new_n27706, new_n27707, new_n27708, new_n27709, new_n27710,
    new_n27711, new_n27712, new_n27713, new_n27714, new_n27715, new_n27716,
    new_n27717, new_n27718, new_n27719, new_n27720, new_n27721, new_n27722,
    new_n27723, new_n27724, new_n27725, new_n27726, new_n27727, new_n27728,
    new_n27729, new_n27730, new_n27731, new_n27732, new_n27733, new_n27734,
    new_n27735, new_n27736, new_n27737, new_n27738, new_n27739, new_n27740,
    new_n27741, new_n27742, new_n27743, new_n27744, new_n27745, new_n27746,
    new_n27747, new_n27748, new_n27749, new_n27750, new_n27751, new_n27752,
    new_n27753, new_n27754, new_n27755, new_n27756, new_n27757, new_n27758,
    new_n27759, new_n27760, new_n27761, new_n27762, new_n27763, new_n27764,
    new_n27765, new_n27766, new_n27767, new_n27768, new_n27769, new_n27770,
    new_n27771, new_n27772, new_n27773, new_n27774, new_n27775, new_n27776,
    new_n27777, new_n27778, new_n27779, new_n27780, new_n27781, new_n27782,
    new_n27783, new_n27784, new_n27785, new_n27786, new_n27787, new_n27788,
    new_n27789, new_n27790, new_n27791, new_n27792, new_n27793, new_n27794,
    new_n27795, new_n27796, new_n27797, new_n27798, new_n27799, new_n27800,
    new_n27801, new_n27802, new_n27803, new_n27804, new_n27805, new_n27806,
    new_n27807, new_n27808, new_n27809, new_n27810, new_n27811, new_n27812,
    new_n27813, new_n27814, new_n27815, new_n27816, new_n27817, new_n27818,
    new_n27819, new_n27820, new_n27821, new_n27822, new_n27823, new_n27824,
    new_n27825, new_n27826, new_n27827, new_n27828, new_n27829, new_n27830,
    new_n27831, new_n27832, new_n27833, new_n27834, new_n27835, new_n27836,
    new_n27837, new_n27838, new_n27839, new_n27840, new_n27841, new_n27842,
    new_n27843, new_n27844, new_n27845, new_n27846, new_n27847, new_n27848,
    new_n27849, new_n27850, new_n27851, new_n27852, new_n27853, new_n27854,
    new_n27855, new_n27856, new_n27857, new_n27858, new_n27859, new_n27860,
    new_n27861, new_n27862, new_n27863, new_n27864, new_n27865, new_n27866,
    new_n27867, new_n27868, new_n27869, new_n27870, new_n27871, new_n27872,
    new_n27873, new_n27874, new_n27875, new_n27876, new_n27877, new_n27878,
    new_n27879, new_n27880, new_n27881, new_n27882, new_n27883, new_n27884,
    new_n27885, new_n27886, new_n27887, new_n27888, new_n27889, new_n27890,
    new_n27891, new_n27892, new_n27893, new_n27894, new_n27895, new_n27896,
    new_n27897, new_n27898, new_n27899, new_n27900, new_n27901, new_n27902,
    new_n27903, new_n27904, new_n27905, new_n27906, new_n27907, new_n27908,
    new_n27909, new_n27910, new_n27911, new_n27912, new_n27913, new_n27914,
    new_n27915, new_n27916, new_n27917, new_n27918, new_n27919, new_n27920,
    new_n27921, new_n27922, new_n27923, new_n27924, new_n27925, new_n27926,
    new_n27927, new_n27928, new_n27929, new_n27930, new_n27931, new_n27932,
    new_n27933, new_n27934, new_n27935, new_n27936, new_n27937, new_n27938,
    new_n27939, new_n27940, new_n27941, new_n27942, new_n27943, new_n27944,
    new_n27945, new_n27946, new_n27947, new_n27948, new_n27949, new_n27950,
    new_n27951, new_n27952, new_n27953, new_n27954, new_n27955, new_n27956,
    new_n27957, new_n27958, new_n27959, new_n27960, new_n27961, new_n27962,
    new_n27963, new_n27964, new_n27965, new_n27966, new_n27967, new_n27968,
    new_n27969, new_n27970, new_n27971, new_n27972, new_n27973, new_n27974,
    new_n27975, new_n27976, new_n27977, new_n27978, new_n27979, new_n27980,
    new_n27981, new_n27982, new_n27983, new_n27984, new_n27985, new_n27986,
    new_n27987, new_n27988, new_n27989, new_n27990, new_n27991, new_n27992,
    new_n27993, new_n27994, new_n27995, new_n27996, new_n27997, new_n27998,
    new_n27999, new_n28000, new_n28001, new_n28002, new_n28003, new_n28004,
    new_n28005, new_n28006, new_n28007, new_n28008, new_n28009, new_n28010,
    new_n28011, new_n28012, new_n28013, new_n28014, new_n28015, new_n28016,
    new_n28017, new_n28018, new_n28019, new_n28020, new_n28021, new_n28022,
    new_n28023, new_n28024, new_n28025, new_n28026, new_n28027, new_n28028,
    new_n28029, new_n28030, new_n28031, new_n28032, new_n28033, new_n28034,
    new_n28035, new_n28036, new_n28037, new_n28038, new_n28039, new_n28040,
    new_n28041, new_n28042, new_n28043, new_n28044, new_n28045, new_n28046,
    new_n28047, new_n28048, new_n28049, new_n28050, new_n28051, new_n28052,
    new_n28053, new_n28054, new_n28055, new_n28056, new_n28057, new_n28058,
    new_n28059, new_n28060, new_n28061, new_n28062, new_n28063, new_n28064,
    new_n28065, new_n28066, new_n28067, new_n28068, new_n28069, new_n28070,
    new_n28071, new_n28072, new_n28073, new_n28074, new_n28075, new_n28076,
    new_n28077, new_n28078, new_n28079, new_n28080, new_n28081, new_n28082,
    new_n28083, new_n28084, new_n28085, new_n28086, new_n28087, new_n28088,
    new_n28089, new_n28090, new_n28091, new_n28092, new_n28093, new_n28094,
    new_n28095, new_n28096, new_n28097, new_n28098, new_n28099, new_n28100,
    new_n28101, new_n28102, new_n28103, new_n28104, new_n28105, new_n28106,
    new_n28107, new_n28108, new_n28109, new_n28110, new_n28111, new_n28112,
    new_n28113, new_n28114, new_n28115, new_n28116, new_n28117, new_n28118,
    new_n28119, new_n28120, new_n28121, new_n28122, new_n28123, new_n28124,
    new_n28125, new_n28126, new_n28127, new_n28128, new_n28129, new_n28130,
    new_n28131, new_n28132, new_n28133, new_n28134, new_n28135, new_n28136,
    new_n28137, new_n28138, new_n28139, new_n28140, new_n28141, new_n28142,
    new_n28143, new_n28144, new_n28145, new_n28146, new_n28147, new_n28148,
    new_n28149, new_n28150, new_n28151, new_n28152, new_n28153, new_n28154,
    new_n28155, new_n28156, new_n28157, new_n28158, new_n28159, new_n28160,
    new_n28161, new_n28162, new_n28163, new_n28164, new_n28165, new_n28166,
    new_n28167, new_n28168, new_n28169, new_n28170, new_n28171, new_n28172,
    new_n28173, new_n28174, new_n28175, new_n28176, new_n28177, new_n28178,
    new_n28179, new_n28180, new_n28181, new_n28182, new_n28183, new_n28184,
    new_n28185, new_n28186, new_n28187, new_n28188, new_n28189, new_n28190,
    new_n28191, new_n28192, new_n28193, new_n28194, new_n28195, new_n28196,
    new_n28197, new_n28198, new_n28199, new_n28200, new_n28201, new_n28202,
    new_n28203, new_n28204, new_n28205, new_n28206, new_n28207, new_n28208,
    new_n28209, new_n28210, new_n28211, new_n28212, new_n28213, new_n28214,
    new_n28215, new_n28216, new_n28217, new_n28218, new_n28219, new_n28220,
    new_n28221, new_n28222, new_n28223, new_n28224, new_n28225, new_n28226,
    new_n28227, new_n28228, new_n28229, new_n28230, new_n28231, new_n28232,
    new_n28233, new_n28234, new_n28235, new_n28236, new_n28237, new_n28238,
    new_n28239, new_n28240, new_n28241, new_n28242, new_n28243, new_n28244,
    new_n28245, new_n28246, new_n28247, new_n28248, new_n28249, new_n28250,
    new_n28251, new_n28252, new_n28253, new_n28254, new_n28255, new_n28256,
    new_n28257, new_n28258, new_n28259, new_n28260, new_n28261, new_n28262,
    new_n28263, new_n28264, new_n28265, new_n28266, new_n28267, new_n28268,
    new_n28269, new_n28270, new_n28271, new_n28272, new_n28273, new_n28274,
    new_n28275, new_n28276, new_n28277, new_n28278, new_n28279, new_n28280,
    new_n28281, new_n28282, new_n28283, new_n28284, new_n28285, new_n28286,
    new_n28287, new_n28288, new_n28289, new_n28290, new_n28291, new_n28292,
    new_n28293, new_n28294, new_n28295, new_n28296, new_n28297, new_n28298,
    new_n28299, new_n28300, new_n28301, new_n28302, new_n28303, new_n28304,
    new_n28305, new_n28306, new_n28307, new_n28308, new_n28309, new_n28310,
    new_n28311, new_n28312, new_n28313, new_n28314, new_n28315, new_n28316,
    new_n28317, new_n28318, new_n28319, new_n28320, new_n28321, new_n28322,
    new_n28323, new_n28324, new_n28325, new_n28326, new_n28327, new_n28328,
    new_n28329, new_n28330, new_n28331, new_n28332, new_n28333, new_n28334,
    new_n28335, new_n28336, new_n28337, new_n28338, new_n28339, new_n28340,
    new_n28341, new_n28342, new_n28343, new_n28344, new_n28345, new_n28346,
    new_n28347, new_n28348, new_n28349, new_n28350, new_n28351, new_n28352,
    new_n28353, new_n28354, new_n28355, new_n28356, new_n28357, new_n28358,
    new_n28359, new_n28360, new_n28361, new_n28362, new_n28363, new_n28364,
    new_n28365, new_n28366, new_n28367, new_n28368, new_n28369, new_n28370,
    new_n28371, new_n28372, new_n28373, new_n28374, new_n28375, new_n28376,
    new_n28377, new_n28378, new_n28379, new_n28380, new_n28381, new_n28382,
    new_n28383, new_n28384, new_n28385, new_n28386, new_n28387, new_n28388,
    new_n28389, new_n28390, new_n28391, new_n28392, new_n28393, new_n28394,
    new_n28395, new_n28396, new_n28397, new_n28398, new_n28399, new_n28400,
    new_n28401, new_n28402, new_n28403, new_n28404, new_n28405, new_n28406,
    new_n28407, new_n28408, new_n28409, new_n28410, new_n28411, new_n28412,
    new_n28413, new_n28414, new_n28415, new_n28416, new_n28417, new_n28418,
    new_n28419, new_n28420, new_n28421, new_n28422, new_n28423, new_n28424,
    new_n28425, new_n28426, new_n28427, new_n28428, new_n28429, new_n28430,
    new_n28431, new_n28432, new_n28433, new_n28434, new_n28435, new_n28436,
    new_n28437, new_n28438, new_n28439, new_n28440, new_n28441, new_n28442,
    new_n28443, new_n28444, new_n28445, new_n28446, new_n28447, new_n28448,
    new_n28449, new_n28450, new_n28451, new_n28452, new_n28453, new_n28454,
    new_n28455, new_n28456, new_n28457, new_n28458, new_n28459, new_n28460,
    new_n28461, new_n28462, new_n28463, new_n28464, new_n28465, new_n28466,
    new_n28467, new_n28468, new_n28469, new_n28470, new_n28471, new_n28472,
    new_n28473, new_n28474, new_n28475, new_n28476, new_n28477, new_n28478,
    new_n28479, new_n28480, new_n28481, new_n28482, new_n28483, new_n28484,
    new_n28485, new_n28486, new_n28487, new_n28488, new_n28489, new_n28490,
    new_n28491, new_n28492, new_n28493, new_n28494, new_n28495, new_n28496,
    new_n28497, new_n28498, new_n28499, new_n28500, new_n28501, new_n28502,
    new_n28503, new_n28504, new_n28505, new_n28506, new_n28507, new_n28508,
    new_n28509, new_n28510, new_n28511, new_n28512, new_n28513, new_n28514,
    new_n28515, new_n28516, new_n28517, new_n28518, new_n28519, new_n28520,
    new_n28521, new_n28522, new_n28523, new_n28524, new_n28525, new_n28526,
    new_n28527, new_n28528, new_n28529, new_n28530, new_n28531, new_n28532,
    new_n28533, new_n28534, new_n28535, new_n28536, new_n28537, new_n28538,
    new_n28539, new_n28540, new_n28541, new_n28542, new_n28543, new_n28544,
    new_n28545, new_n28546, new_n28547, new_n28548, new_n28549, new_n28550,
    new_n28551, new_n28552, new_n28553, new_n28554, new_n28555, new_n28556,
    new_n28557, new_n28558, new_n28559, new_n28560, new_n28561, new_n28562,
    new_n28563, new_n28564, new_n28565, new_n28566, new_n28567, new_n28568,
    new_n28569, new_n28570, new_n28571, new_n28572, new_n28573, new_n28574,
    new_n28575, new_n28576, new_n28577, new_n28578, new_n28579, new_n28580,
    new_n28581, new_n28582, new_n28583, new_n28584, new_n28585, new_n28586,
    new_n28587, new_n28588, new_n28589, new_n28590, new_n28591, new_n28592,
    new_n28593, new_n28594, new_n28595, new_n28596, new_n28597, new_n28598,
    new_n28599, new_n28600, new_n28601, new_n28602, new_n28603, new_n28604,
    new_n28605, new_n28606, new_n28607, new_n28608, new_n28609, new_n28610,
    new_n28611, new_n28612, new_n28613, new_n28614, new_n28615, new_n28616,
    new_n28617, new_n28618, new_n28619, new_n28620, new_n28621, new_n28622,
    new_n28623, new_n28624, new_n28625, new_n28626, new_n28627, new_n28628,
    new_n28629, new_n28630, new_n28631, new_n28632, new_n28633, new_n28634,
    new_n28635, new_n28636, new_n28637, new_n28638, new_n28639, new_n28640,
    new_n28641, new_n28642, new_n28643, new_n28644, new_n28645, new_n28646,
    new_n28647, new_n28648, new_n28649, new_n28650, new_n28651, new_n28652,
    new_n28653, new_n28654, new_n28655, new_n28656, new_n28657, new_n28658,
    new_n28659, new_n28660, new_n28661, new_n28662, new_n28663, new_n28664,
    new_n28665, new_n28666, new_n28667, new_n28668, new_n28669, new_n28670,
    new_n28671, new_n28672, new_n28673, new_n28674, new_n28675, new_n28676,
    new_n28677, new_n28678, new_n28679, new_n28680, new_n28681, new_n28682,
    new_n28683, new_n28684, new_n28685, new_n28686, new_n28687, new_n28688,
    new_n28689, new_n28690, new_n28691, new_n28692, new_n28693, new_n28694,
    new_n28695, new_n28696, new_n28697, new_n28698, new_n28699, new_n28700,
    new_n28701, new_n28702, new_n28703, new_n28704, new_n28705, new_n28706,
    new_n28707, new_n28708, new_n28709, new_n28710, new_n28711, new_n28712,
    new_n28713, new_n28714, new_n28715, new_n28716, new_n28717, new_n28718,
    new_n28719, new_n28720, new_n28721, new_n28722, new_n28723, new_n28724,
    new_n28725, new_n28726, new_n28727, new_n28728, new_n28729, new_n28730,
    new_n28731, new_n28732, new_n28733, new_n28734, new_n28735, new_n28736,
    new_n28737, new_n28738, new_n28739, new_n28740, new_n28741, new_n28742,
    new_n28743, new_n28744, new_n28745, new_n28746, new_n28747, new_n28748,
    new_n28749, new_n28750, new_n28751, new_n28752, new_n28753, new_n28754,
    new_n28755, new_n28756, new_n28757, new_n28758, new_n28759, new_n28760,
    new_n28761, new_n28762, new_n28763, new_n28764, new_n28765, new_n28766,
    new_n28767, new_n28768, new_n28769, new_n28770, new_n28771, new_n28772,
    new_n28773, new_n28774, new_n28775, new_n28776, new_n28777, new_n28778,
    new_n28779, new_n28780, new_n28781, new_n28782, new_n28783, new_n28784,
    new_n28785, new_n28786, new_n28787, new_n28788, new_n28789, new_n28790,
    new_n28791, new_n28792, new_n28793, new_n28794, new_n28795, new_n28796,
    new_n28797, new_n28798, new_n28799, new_n28800, new_n28801, new_n28802,
    new_n28803, new_n28804, new_n28805, new_n28806, new_n28807, new_n28808,
    new_n28809, new_n28810, new_n28811, new_n28812, new_n28813, new_n28814,
    new_n28815, new_n28816, new_n28817, new_n28818, new_n28819, new_n28820,
    new_n28821, new_n28822, new_n28823, new_n28824, new_n28825, new_n28826,
    new_n28827, new_n28828, new_n28829, new_n28830, new_n28831, new_n28832,
    new_n28833, new_n28834, new_n28835, new_n28836, new_n28837, new_n28838,
    new_n28839, new_n28840, new_n28841, new_n28842, new_n28843, new_n28844,
    new_n28845, new_n28846, new_n28847, new_n28848, new_n28849, new_n28850,
    new_n28851, new_n28852, new_n28853, new_n28854, new_n28855, new_n28856,
    new_n28857, new_n28858, new_n28859, new_n28860, new_n28861, new_n28862,
    new_n28863, new_n28864, new_n28865, new_n28866, new_n28867, new_n28868,
    new_n28869, new_n28870, new_n28871, new_n28872, new_n28873, new_n28874,
    new_n28875, new_n28876, new_n28877, new_n28878, new_n28879, new_n28880,
    new_n28881, new_n28882, new_n28883, new_n28884, new_n28885, new_n28886,
    new_n28887, new_n28888, new_n28889, new_n28890, new_n28891, new_n28892,
    new_n28893, new_n28894, new_n28895, new_n28896, new_n28897, new_n28898,
    new_n28899, new_n28900, new_n28901, new_n28902, new_n28903, new_n28904,
    new_n28905, new_n28906, new_n28907, new_n28908, new_n28909, new_n28910,
    new_n28911, new_n28912, new_n28913, new_n28914, new_n28915, new_n28916,
    new_n28917, new_n28918, new_n28919, new_n28920, new_n28921, new_n28922,
    new_n28923, new_n28924, new_n28925, new_n28926, new_n28927, new_n28928,
    new_n28929, new_n28930, new_n28931, new_n28932, new_n28933, new_n28934,
    new_n28935, new_n28936, new_n28937, new_n28938, new_n28939, new_n28940,
    new_n28941, new_n28942, new_n28943, new_n28944, new_n28945, new_n28946,
    new_n28947, new_n28948, new_n28949, new_n28950, new_n28951, new_n28952,
    new_n28953, new_n28954, new_n28955, new_n28956, new_n28957, new_n28958,
    new_n28959, new_n28960, new_n28961, new_n28962, new_n28963, new_n28964,
    new_n28965, new_n28966, new_n28967, new_n28968, new_n28969, new_n28970,
    new_n28971, new_n28972, new_n28973, new_n28974, new_n28975, new_n28976,
    new_n28977, new_n28978, new_n28979, new_n28980, new_n28981, new_n28982,
    new_n28983, new_n28984, new_n28985, new_n28986, new_n28987, new_n28988,
    new_n28989, new_n28990, new_n28991, new_n28992, new_n28993, new_n28994,
    new_n28995, new_n28996, new_n28997, new_n28998, new_n28999, new_n29000,
    new_n29001, new_n29002, new_n29003, new_n29004, new_n29005, new_n29006,
    new_n29007, new_n29008, new_n29009, new_n29010, new_n29011, new_n29012,
    new_n29013, new_n29014, new_n29015, new_n29016, new_n29017, new_n29018,
    new_n29019, new_n29020, new_n29021, new_n29022, new_n29023, new_n29024,
    new_n29025, new_n29026, new_n29027, new_n29028, new_n29029, new_n29030,
    new_n29031, new_n29032, new_n29033, new_n29034, new_n29035, new_n29036,
    new_n29037, new_n29038, new_n29039, new_n29040, new_n29041, new_n29042,
    new_n29043, new_n29044, new_n29045, new_n29046, new_n29047, new_n29048,
    new_n29049, new_n29050, new_n29051, new_n29052, new_n29053, new_n29054,
    new_n29055, new_n29056, new_n29057, new_n29058, new_n29059, new_n29060,
    new_n29061, new_n29062, new_n29063, new_n29064, new_n29065, new_n29066,
    new_n29067, new_n29068, new_n29069, new_n29070, new_n29071, new_n29072,
    new_n29073, new_n29074, new_n29075, new_n29076, new_n29077, new_n29078,
    new_n29079, new_n29080, new_n29081, new_n29082, new_n29083, new_n29084,
    new_n29085, new_n29086, new_n29087, new_n29088, new_n29089, new_n29090,
    new_n29091, new_n29092, new_n29093, new_n29094, new_n29095, new_n29096,
    new_n29097, new_n29098, new_n29099, new_n29100, new_n29101, new_n29102,
    new_n29103, new_n29104, new_n29105, new_n29106, new_n29107, new_n29108,
    new_n29109, new_n29110, new_n29111, new_n29112, new_n29113, new_n29114,
    new_n29115, new_n29116, new_n29117, new_n29118, new_n29119, new_n29120,
    new_n29121, new_n29122, new_n29123, new_n29124, new_n29125, new_n29126,
    new_n29127, new_n29128, new_n29129, new_n29130, new_n29131, new_n29132,
    new_n29133, new_n29134, new_n29135, new_n29136, new_n29137, new_n29138,
    new_n29139, new_n29140, new_n29141, new_n29142, new_n29143, new_n29144,
    new_n29145, new_n29146, new_n29147, new_n29148, new_n29149, new_n29150,
    new_n29151, new_n29152, new_n29153, new_n29154, new_n29155, new_n29156,
    new_n29157, new_n29158, new_n29159, new_n29160, new_n29161, new_n29162,
    new_n29163, new_n29164, new_n29165, new_n29166, new_n29167, new_n29168,
    new_n29169, new_n29170, new_n29171, new_n29172, new_n29173, new_n29174,
    new_n29175, new_n29176, new_n29177, new_n29178, new_n29179, new_n29180,
    new_n29181, new_n29182, new_n29183, new_n29184, new_n29185, new_n29186,
    new_n29187, new_n29188, new_n29189, new_n29190, new_n29191, new_n29192,
    new_n29193, new_n29194, new_n29195, new_n29196, new_n29197, new_n29198,
    new_n29199, new_n29200, new_n29201, new_n29202, new_n29203, new_n29204,
    new_n29205, new_n29206, new_n29207, new_n29208, new_n29209, new_n29210,
    new_n29211, new_n29212, new_n29213, new_n29214, new_n29215, new_n29216,
    new_n29217, new_n29218, new_n29219, new_n29220, new_n29221, new_n29222,
    new_n29223, new_n29224, new_n29225, new_n29226, new_n29227, new_n29228,
    new_n29229, new_n29230, new_n29231, new_n29232, new_n29233, new_n29234,
    new_n29235, new_n29236, new_n29237, new_n29238, new_n29239, new_n29240,
    new_n29241, new_n29242, new_n29243, new_n29244, new_n29245, new_n29246,
    new_n29247, new_n29248, new_n29249, new_n29250, new_n29251, new_n29252,
    new_n29253, new_n29254, new_n29255, new_n29256, new_n29257, new_n29258,
    new_n29259, new_n29260, new_n29261, new_n29262, new_n29263, new_n29264,
    new_n29265, new_n29266, new_n29267, new_n29268, new_n29269, new_n29270,
    new_n29271, new_n29272, new_n29273, new_n29274, new_n29275, new_n29276,
    new_n29277, new_n29278, new_n29279, new_n29280, new_n29281, new_n29282,
    new_n29283, new_n29284, new_n29285, new_n29286, new_n29287, new_n29288,
    new_n29289, new_n29290, new_n29291, new_n29292, new_n29293, new_n29294,
    new_n29295, new_n29296, new_n29297, new_n29298, new_n29299, new_n29300,
    new_n29301, new_n29302, new_n29303, new_n29304, new_n29305, new_n29306,
    new_n29307, new_n29308, new_n29309, new_n29310, new_n29311, new_n29312,
    new_n29313, new_n29314, new_n29315, new_n29316, new_n29317, new_n29318,
    new_n29319, new_n29320, new_n29321, new_n29322, new_n29323, new_n29324,
    new_n29325, new_n29326, new_n29327, new_n29328, new_n29329, new_n29330,
    new_n29331, new_n29332, new_n29333, new_n29334, new_n29335, new_n29336,
    new_n29337, new_n29338, new_n29339, new_n29340, new_n29341, new_n29342,
    new_n29343, new_n29344, new_n29345, new_n29346, new_n29347, new_n29348,
    new_n29349, new_n29350, new_n29351, new_n29352, new_n29353, new_n29354,
    new_n29355, new_n29356, new_n29357, new_n29358, new_n29359, new_n29360,
    new_n29361, new_n29362, new_n29363, new_n29364, new_n29365, new_n29366,
    new_n29367, new_n29368, new_n29369, new_n29370, new_n29371, new_n29372,
    new_n29373, new_n29374, new_n29375, new_n29376, new_n29377, new_n29378,
    new_n29379, new_n29380, new_n29381, new_n29382, new_n29383, new_n29384,
    new_n29385, new_n29386, new_n29387, new_n29388, new_n29389, new_n29390,
    new_n29391, new_n29392, new_n29393, new_n29394, new_n29395, new_n29396,
    new_n29397, new_n29398, new_n29399, new_n29400, new_n29401, new_n29402,
    new_n29403, new_n29404, new_n29405, new_n29406, new_n29407, new_n29408,
    new_n29409, new_n29410, new_n29411, new_n29412, new_n29413, new_n29414,
    new_n29415, new_n29416, new_n29417, new_n29418, new_n29419, new_n29420,
    new_n29421, new_n29422, new_n29423, new_n29424, new_n29425, new_n29426,
    new_n29427, new_n29428, new_n29429, new_n29430, new_n29431, new_n29432,
    new_n29433, new_n29434, new_n29435, new_n29436, new_n29437, new_n29438,
    new_n29439, new_n29440, new_n29441, new_n29442, new_n29443, new_n29444,
    new_n29445, new_n29446, new_n29447, new_n29448, new_n29449, new_n29450,
    new_n29451, new_n29452, new_n29453, new_n29454, new_n29455, new_n29456,
    new_n29457, new_n29458, new_n29459, new_n29460, new_n29461, new_n29462,
    new_n29463, new_n29464, new_n29465, new_n29466, new_n29467, new_n29468,
    new_n29469, new_n29470, new_n29471, new_n29472, new_n29473, new_n29474,
    new_n29475, new_n29476, new_n29477, new_n29478, new_n29479, new_n29480,
    new_n29481, new_n29482, new_n29483, new_n29484, new_n29485, new_n29486,
    new_n29487, new_n29488, new_n29489, new_n29490, new_n29491, new_n29492,
    new_n29493, new_n29494, new_n29495, new_n29496, new_n29497, new_n29498,
    new_n29499, new_n29500, new_n29501, new_n29502, new_n29503, new_n29504,
    new_n29505, new_n29506, new_n29507, new_n29508, new_n29509, new_n29510,
    new_n29511, new_n29512, new_n29513, new_n29514, new_n29515, new_n29516,
    new_n29517, new_n29518, new_n29519, new_n29520, new_n29521, new_n29522,
    new_n29523, new_n29524, new_n29525, new_n29526, new_n29527, new_n29528,
    new_n29529, new_n29530, new_n29531, new_n29532, new_n29533, new_n29534,
    new_n29535, new_n29536, new_n29537, new_n29538, new_n29539, new_n29540,
    new_n29541, new_n29542, new_n29543, new_n29544, new_n29545, new_n29546,
    new_n29547, new_n29548, new_n29549, new_n29550, new_n29551, new_n29552,
    new_n29553, new_n29554, new_n29555, new_n29556, new_n29557, new_n29558,
    new_n29559, new_n29560, new_n29561, new_n29562, new_n29563, new_n29564,
    new_n29565, new_n29566, new_n29567, new_n29568, new_n29569, new_n29570,
    new_n29571, new_n29572, new_n29573, new_n29574, new_n29575, new_n29576,
    new_n29577, new_n29578, new_n29579, new_n29580, new_n29581, new_n29582,
    new_n29583, new_n29584, new_n29585, new_n29586, new_n29587, new_n29588,
    new_n29589, new_n29590, new_n29591, new_n29592, new_n29593, new_n29594,
    new_n29595, new_n29596, new_n29597, new_n29598, new_n29599, new_n29600,
    new_n29601, new_n29602, new_n29603, new_n29604, new_n29605, new_n29606,
    new_n29607, new_n29608, new_n29609, new_n29610, new_n29611, new_n29612,
    new_n29613, new_n29614, new_n29615, new_n29616, new_n29617, new_n29618,
    new_n29619, new_n29620, new_n29621, new_n29622, new_n29623, new_n29624,
    new_n29625, new_n29626, new_n29627, new_n29628, new_n29629, new_n29630,
    new_n29631, new_n29632, new_n29633, new_n29634, new_n29635, new_n29636,
    new_n29637, new_n29638, new_n29639, new_n29640, new_n29641, new_n29642,
    new_n29643, new_n29644, new_n29645, new_n29646, new_n29647, new_n29648,
    new_n29649, new_n29650, new_n29651, new_n29652, new_n29653, new_n29654,
    new_n29655, new_n29656, new_n29657, new_n29658, new_n29659, new_n29660,
    new_n29661, new_n29662, new_n29663, new_n29664, new_n29665, new_n29666,
    new_n29667, new_n29668, new_n29669, new_n29670, new_n29671, new_n29672,
    new_n29673, new_n29674, new_n29675, new_n29676, new_n29677, new_n29678,
    new_n29679, new_n29680, new_n29681, new_n29682, new_n29683, new_n29684,
    new_n29685, new_n29686, new_n29687, new_n29688, new_n29689, new_n29690,
    new_n29691, new_n29692, new_n29693, new_n29694, new_n29695, new_n29696,
    new_n29697, new_n29698, new_n29699, new_n29700, new_n29701, new_n29702,
    new_n29703, new_n29704, new_n29705, new_n29706, new_n29707, new_n29708,
    new_n29709, new_n29710, new_n29711, new_n29712, new_n29713, new_n29714,
    new_n29715, new_n29716, new_n29717, new_n29718, new_n29719, new_n29720,
    new_n29721, new_n29722, new_n29723, new_n29724, new_n29725, new_n29726,
    new_n29727, new_n29728, new_n29729, new_n29730, new_n29731, new_n29732,
    new_n29733, new_n29734, new_n29735, new_n29736, new_n29737, new_n29738,
    new_n29739, new_n29740, new_n29741, new_n29742, new_n29743, new_n29744,
    new_n29745, new_n29746, new_n29747, new_n29748, new_n29749, new_n29750,
    new_n29751, new_n29752, new_n29753, new_n29754, new_n29755, new_n29756,
    new_n29757, new_n29758, new_n29759, new_n29760, new_n29761, new_n29762,
    new_n29763, new_n29764, new_n29765, new_n29766, new_n29767, new_n29768,
    new_n29769, new_n29770, new_n29771, new_n29772, new_n29773, new_n29774,
    new_n29775, new_n29776, new_n29777, new_n29778, new_n29779, new_n29780,
    new_n29781, new_n29782, new_n29783, new_n29784, new_n29785, new_n29786,
    new_n29787, new_n29788, new_n29789, new_n29790, new_n29791, new_n29792,
    new_n29793, new_n29794, new_n29795, new_n29796, new_n29797, new_n29798,
    new_n29799, new_n29800, new_n29801, new_n29802, new_n29803, new_n29804,
    new_n29805, new_n29806, new_n29807, new_n29808, new_n29809, new_n29810,
    new_n29811, new_n29812, new_n29813, new_n29814, new_n29815, new_n29816,
    new_n29817, new_n29818, new_n29819, new_n29820, new_n29821, new_n29822,
    new_n29823, new_n29824, new_n29825, new_n29826, new_n29827, new_n29828,
    new_n29829, new_n29830, new_n29831, new_n29832, new_n29833, new_n29834,
    new_n29835, new_n29836, new_n29837, new_n29838, new_n29839, new_n29840,
    new_n29841, new_n29842, new_n29843, new_n29844, new_n29845, new_n29846,
    new_n29847, new_n29848, new_n29849, new_n29850, new_n29851, new_n29852,
    new_n29853, new_n29854, new_n29855, new_n29856, new_n29857, new_n29858,
    new_n29859, new_n29860, new_n29861, new_n29862, new_n29863, new_n29864,
    new_n29865, new_n29866, new_n29867, new_n29868, new_n29869, new_n29870,
    new_n29871, new_n29872, new_n29873, new_n29874, new_n29875, new_n29876,
    new_n29877, new_n29878, new_n29879, new_n29880, new_n29881, new_n29882,
    new_n29883, new_n29884, new_n29885, new_n29886, new_n29887, new_n29888,
    new_n29889, new_n29890, new_n29891, new_n29892, new_n29893, new_n29894,
    new_n29895, new_n29896, new_n29897, new_n29898, new_n29899, new_n29900,
    new_n29901, new_n29902, new_n29903, new_n29904, new_n29905, new_n29906,
    new_n29907, new_n29908, new_n29909, new_n29910, new_n29911, new_n29912,
    new_n29913, new_n29914, new_n29915, new_n29916, new_n29917, new_n29918,
    new_n29919, new_n29920, new_n29921, new_n29922, new_n29923, new_n29924,
    new_n29925, new_n29926, new_n29927, new_n29928, new_n29929, new_n29930,
    new_n29931, new_n29932, new_n29933, new_n29934, new_n29935, new_n29936,
    new_n29937, new_n29938, new_n29939, new_n29940, new_n29941, new_n29942,
    new_n29943, new_n29944, new_n29945, new_n29946, new_n29947, new_n29948,
    new_n29949, new_n29950, new_n29951, new_n29952, new_n29953, new_n29954,
    new_n29955, new_n29956, new_n29957, new_n29958, new_n29959, new_n29960,
    new_n29961, new_n29962, new_n29963, new_n29964, new_n29965, new_n29966,
    new_n29967, new_n29968, new_n29969, new_n29970, new_n29971, new_n29972,
    new_n29973, new_n29974, new_n29975, new_n29976, new_n29977, new_n29978,
    new_n29979, new_n29980, new_n29981, new_n29982, new_n29983, new_n29984,
    new_n29985, new_n29986, new_n29987, new_n29988, new_n29989, new_n29990,
    new_n29991, new_n29992, new_n29993, new_n29994, new_n29995, new_n29996,
    new_n29997, new_n29998, new_n29999, new_n30000, new_n30001, new_n30002,
    new_n30003, new_n30004, new_n30005, new_n30006, new_n30007, new_n30008,
    new_n30009, new_n30010, new_n30011, new_n30012, new_n30013, new_n30014,
    new_n30015, new_n30016, new_n30017, new_n30018, new_n30019, new_n30020,
    new_n30021, new_n30022, new_n30023, new_n30024, new_n30025, new_n30026,
    new_n30027, new_n30028, new_n30029, new_n30030, new_n30031, new_n30032,
    new_n30033, new_n30034, new_n30035, new_n30036, new_n30037, new_n30038,
    new_n30039, new_n30040, new_n30041, new_n30042, new_n30043, new_n30044,
    new_n30045, new_n30046, new_n30047, new_n30048, new_n30049, new_n30050,
    new_n30051, new_n30052, new_n30053, new_n30054, new_n30055, new_n30056,
    new_n30057, new_n30058, new_n30059, new_n30060, new_n30061, new_n30062,
    new_n30063, new_n30064, new_n30065, new_n30066, new_n30067, new_n30068,
    new_n30069, new_n30070, new_n30071, new_n30072, new_n30073, new_n30074,
    new_n30075, new_n30076, new_n30077, new_n30078, new_n30079, new_n30080,
    new_n30081, new_n30082, new_n30083, new_n30084, new_n30085, new_n30086,
    new_n30087, new_n30088, new_n30089, new_n30090, new_n30091, new_n30092,
    new_n30093, new_n30094, new_n30095, new_n30096, new_n30097, new_n30098,
    new_n30099, new_n30100, new_n30101, new_n30102, new_n30103, new_n30104,
    new_n30105, new_n30106, new_n30107, new_n30108, new_n30109, new_n30110,
    new_n30111, new_n30112, new_n30113, new_n30114, new_n30115, new_n30116,
    new_n30117, new_n30118, new_n30119, new_n30120, new_n30121, new_n30122,
    new_n30123, new_n30124, new_n30125, new_n30126, new_n30127, new_n30128,
    new_n30129, new_n30130, new_n30131, new_n30132, new_n30133, new_n30134,
    new_n30135, new_n30136, new_n30137, new_n30138, new_n30139, new_n30140,
    new_n30141, new_n30142, new_n30143, new_n30144, new_n30145, new_n30146,
    new_n30147, new_n30148, new_n30149, new_n30150, new_n30151, new_n30152,
    new_n30153, new_n30154, new_n30155, new_n30156, new_n30157, new_n30158,
    new_n30159, new_n30160, new_n30161, new_n30162, new_n30163, new_n30164,
    new_n30165, new_n30166, new_n30167, new_n30168, new_n30169, new_n30170,
    new_n30171, new_n30172, new_n30173, new_n30174, new_n30175, new_n30176,
    new_n30177, new_n30178, new_n30179, new_n30180, new_n30181, new_n30182,
    new_n30183, new_n30184, new_n30185, new_n30186, new_n30187, new_n30188,
    new_n30189, new_n30190, new_n30191, new_n30192, new_n30193, new_n30194,
    new_n30195, new_n30196, new_n30197, new_n30198, new_n30199, new_n30200,
    new_n30201, new_n30202, new_n30203, new_n30204, new_n30205, new_n30206,
    new_n30207, new_n30208, new_n30209, new_n30210, new_n30211, new_n30212,
    new_n30213, new_n30214, new_n30215, new_n30216, new_n30217, new_n30218,
    new_n30219, new_n30220, new_n30221, new_n30222, new_n30223, new_n30224,
    new_n30225, new_n30226, new_n30227, new_n30228, new_n30229, new_n30230,
    new_n30231, new_n30232, new_n30233, new_n30234, new_n30235, new_n30236,
    new_n30237, new_n30238, new_n30239, new_n30240, new_n30241, new_n30242,
    new_n30243, new_n30244, new_n30245, new_n30246, new_n30247, new_n30248,
    new_n30249, new_n30250, new_n30251, new_n30252, new_n30253, new_n30254,
    new_n30255, new_n30256, new_n30257, new_n30258, new_n30259, new_n30260,
    new_n30261, new_n30262, new_n30263, new_n30264, new_n30265, new_n30266,
    new_n30267, new_n30268, new_n30269, new_n30270, new_n30271, new_n30272,
    new_n30273, new_n30274, new_n30275, new_n30276, new_n30277, new_n30278,
    new_n30279, new_n30280, new_n30281, new_n30282, new_n30283, new_n30284,
    new_n30285, new_n30286, new_n30287, new_n30288, new_n30289, new_n30290,
    new_n30291, new_n30292, new_n30293, new_n30294, new_n30295, new_n30296,
    new_n30297, new_n30298, new_n30299, new_n30300, new_n30301, new_n30302,
    new_n30303, new_n30304, new_n30305, new_n30306, new_n30307, new_n30308,
    new_n30309, new_n30310, new_n30311, new_n30312, new_n30313, new_n30314,
    new_n30315, new_n30316, new_n30317, new_n30318, new_n30319, new_n30320,
    new_n30321, new_n30322, new_n30323, new_n30324, new_n30325, new_n30326,
    new_n30327, new_n30328, new_n30329, new_n30330, new_n30331, new_n30332,
    new_n30333, new_n30334, new_n30335, new_n30336, new_n30337, new_n30338,
    new_n30339, new_n30340, new_n30341, new_n30342, new_n30343, new_n30344,
    new_n30345, new_n30346, new_n30347, new_n30348, new_n30349, new_n30350,
    new_n30351, new_n30352, new_n30353, new_n30354, new_n30355, new_n30356,
    new_n30357, new_n30358, new_n30359, new_n30360, new_n30361, new_n30362,
    new_n30363, new_n30364, new_n30365, new_n30366, new_n30367, new_n30368,
    new_n30369, new_n30370, new_n30371, new_n30372, new_n30373, new_n30374,
    new_n30375, new_n30376, new_n30377, new_n30378, new_n30379, new_n30380,
    new_n30381, new_n30382, new_n30383, new_n30384, new_n30385, new_n30386,
    new_n30387, new_n30388, new_n30389, new_n30390, new_n30391, new_n30392,
    new_n30393, new_n30394, new_n30395, new_n30396, new_n30397, new_n30398,
    new_n30399, new_n30400, new_n30401, new_n30402, new_n30403, new_n30404,
    new_n30405, new_n30406, new_n30407, new_n30408, new_n30409, new_n30410,
    new_n30411, new_n30412, new_n30413, new_n30414, new_n30415, new_n30416,
    new_n30417, new_n30418, new_n30419, new_n30420, new_n30421, new_n30422,
    new_n30423, new_n30424, new_n30425, new_n30426, new_n30427, new_n30428,
    new_n30429, new_n30430, new_n30431, new_n30432, new_n30433, new_n30434,
    new_n30435, new_n30436, new_n30437, new_n30438, new_n30439, new_n30440,
    new_n30441, new_n30442, new_n30443, new_n30444, new_n30445, new_n30446,
    new_n30447, new_n30448, new_n30449, new_n30450, new_n30451, new_n30452,
    new_n30453, new_n30454, new_n30455, new_n30456, new_n30457, new_n30458,
    new_n30459, new_n30460, new_n30461, new_n30462, new_n30463, new_n30464,
    new_n30465, new_n30466, new_n30467, new_n30468, new_n30469, new_n30470,
    new_n30471, new_n30472, new_n30473, new_n30474, new_n30475, new_n30476,
    new_n30477, new_n30478, new_n30479, new_n30480, new_n30481, new_n30482,
    new_n30483, new_n30484, new_n30485, new_n30486, new_n30487, new_n30488,
    new_n30489, new_n30490, new_n30491, new_n30492, new_n30493, new_n30494,
    new_n30495, new_n30496, new_n30497, new_n30498, new_n30499, new_n30500,
    new_n30501, new_n30502, new_n30503, new_n30504, new_n30505, new_n30506,
    new_n30507, new_n30508, new_n30509, new_n30510, new_n30511, new_n30512,
    new_n30513, new_n30514, new_n30515, new_n30516, new_n30517, new_n30518,
    new_n30519, new_n30520, new_n30521, new_n30522, new_n30523, new_n30524,
    new_n30525, new_n30526, new_n30527, new_n30528, new_n30529, new_n30530,
    new_n30531, new_n30532, new_n30533, new_n30534, new_n30535, new_n30536,
    new_n30537, new_n30538, new_n30539, new_n30540, new_n30541, new_n30542,
    new_n30543, new_n30544, new_n30545, new_n30546, new_n30547, new_n30548,
    new_n30549, new_n30550, new_n30551, new_n30552, new_n30553, new_n30554,
    new_n30555, new_n30556, new_n30557, new_n30558, new_n30559, new_n30560,
    new_n30561, new_n30562, new_n30563, new_n30564, new_n30565, new_n30566,
    new_n30567, new_n30568, new_n30569, new_n30570, new_n30571, new_n30572,
    new_n30573, new_n30574, new_n30575, new_n30576, new_n30577, new_n30578,
    new_n30579, new_n30580, new_n30581, new_n30582, new_n30583, new_n30584,
    new_n30585, new_n30586, new_n30587, new_n30588, new_n30589, new_n30590,
    new_n30591, new_n30592, new_n30593, new_n30594, new_n30595, new_n30596,
    new_n30597, new_n30598, new_n30599, new_n30600, new_n30601, new_n30602,
    new_n30603, new_n30604, new_n30605, new_n30606, new_n30607, new_n30608,
    new_n30609, new_n30610, new_n30611, new_n30612, new_n30613, new_n30614,
    new_n30615, new_n30616, new_n30617, new_n30618, new_n30619, new_n30620,
    new_n30621, new_n30622, new_n30623, new_n30624, new_n30625, new_n30626,
    new_n30627, new_n30628, new_n30629, new_n30630, new_n30631, new_n30632,
    new_n30633, new_n30634, new_n30635, new_n30636, new_n30637, new_n30638,
    new_n30639, new_n30640, new_n30641, new_n30642, new_n30643, new_n30644,
    new_n30645, new_n30646, new_n30647, new_n30648, new_n30649, new_n30650,
    new_n30651, new_n30652, new_n30653, new_n30654, new_n30655, new_n30656,
    new_n30657, new_n30658, new_n30659, new_n30660, new_n30661, new_n30662,
    new_n30663, new_n30664, new_n30665, new_n30666, new_n30667, new_n30668,
    new_n30669, new_n30670, new_n30671, new_n30672, new_n30673, new_n30674,
    new_n30675, new_n30676, new_n30677, new_n30678, new_n30679, new_n30680,
    new_n30681, new_n30682, new_n30683, new_n30684, new_n30685, new_n30686,
    new_n30687, new_n30688, new_n30689, new_n30690, new_n30691, new_n30692,
    new_n30693, new_n30694, new_n30695, new_n30696, new_n30697, new_n30698,
    new_n30699, new_n30700, new_n30701, new_n30702, new_n30703, new_n30704,
    new_n30705, new_n30706, new_n30707, new_n30708, new_n30709, new_n30710,
    new_n30711, new_n30712, new_n30713, new_n30714, new_n30715, new_n30716,
    new_n30717, new_n30718, new_n30719, new_n30720, new_n30721, new_n30722,
    new_n30723, new_n30724, new_n30725, new_n30726, new_n30727, new_n30728,
    new_n30729, new_n30730, new_n30731, new_n30732, new_n30733, new_n30734,
    new_n30735, new_n30736, new_n30737, new_n30738, new_n30739, new_n30740,
    new_n30741, new_n30742, new_n30743, new_n30744, new_n30745, new_n30746,
    new_n30747, new_n30748, new_n30749, new_n30750, new_n30751, new_n30752,
    new_n30753, new_n30754, new_n30755, new_n30756, new_n30757, new_n30758,
    new_n30759, new_n30760, new_n30761, new_n30762, new_n30763, new_n30764,
    new_n30765, new_n30766, new_n30767, new_n30768, new_n30769, new_n30770,
    new_n30771, new_n30772, new_n30773, new_n30774, new_n30775, new_n30776,
    new_n30777, new_n30778, new_n30779, new_n30780, new_n30781, new_n30782,
    new_n30783, new_n30784, new_n30785, new_n30786, new_n30787, new_n30788,
    new_n30789, new_n30790, new_n30791, new_n30792, new_n30793, new_n30794,
    new_n30795, new_n30796, new_n30797, new_n30798, new_n30799, new_n30800,
    new_n30801, new_n30802, new_n30803, new_n30804, new_n30805, new_n30806,
    new_n30807, new_n30808, new_n30809, new_n30810, new_n30811, new_n30812,
    new_n30813, new_n30814, new_n30815, new_n30816, new_n30817, new_n30818,
    new_n30819, new_n30820, new_n30821, new_n30822, new_n30823, new_n30824,
    new_n30825, new_n30826, new_n30827, new_n30828, new_n30829, new_n30830,
    new_n30831, new_n30832, new_n30833, new_n30834, new_n30835, new_n30836,
    new_n30837, new_n30838, new_n30839, new_n30840, new_n30841, new_n30842,
    new_n30843, new_n30844, new_n30845, new_n30846, new_n30847, new_n30848,
    new_n30849, new_n30850, new_n30851, new_n30852, new_n30853, new_n30854,
    new_n30855, new_n30856, new_n30857, new_n30858, new_n30859, new_n30860,
    new_n30861, new_n30862, new_n30863, new_n30864, new_n30865, new_n30866,
    new_n30867, new_n30868, new_n30869, new_n30870, new_n30871, new_n30872,
    new_n30873, new_n30874, new_n30875, new_n30876, new_n30877, new_n30878,
    new_n30879, new_n30880, new_n30881, new_n30882, new_n30883, new_n30884,
    new_n30885, new_n30886, new_n30887, new_n30888, new_n30889, new_n30890,
    new_n30891, new_n30892, new_n30893, new_n30894, new_n30895, new_n30896,
    new_n30897, new_n30898, new_n30899, new_n30900, new_n30901, new_n30902,
    new_n30903, new_n30904, new_n30905, new_n30906, new_n30907, new_n30908,
    new_n30909, new_n30910, new_n30911, new_n30912, new_n30913, new_n30914,
    new_n30915, new_n30916, new_n30917, new_n30918, new_n30919, new_n30920,
    new_n30921, new_n30922, new_n30923, new_n30924, new_n30925, new_n30926,
    new_n30927, new_n30928, new_n30929, new_n30930, new_n30931, new_n30932,
    new_n30933, new_n30934, new_n30935, new_n30936, new_n30937, new_n30938,
    new_n30939, new_n30940, new_n30941, new_n30942, new_n30943, new_n30944,
    new_n30945, new_n30946, new_n30947, new_n30948, new_n30949, new_n30950,
    new_n30951, new_n30952, new_n30953, new_n30954, new_n30955, new_n30956,
    new_n30957, new_n30958, new_n30959, new_n30960, new_n30961, new_n30962,
    new_n30963, new_n30964, new_n30965, new_n30966, new_n30967, new_n30968,
    new_n30969, new_n30970, new_n30971, new_n30972, new_n30973, new_n30974,
    new_n30975, new_n30976, new_n30977, new_n30978, new_n30979, new_n30980,
    new_n30981, new_n30982, new_n30983, new_n30984, new_n30985, new_n30986,
    new_n30987, new_n30988, new_n30989, new_n30990, new_n30991, new_n30992,
    new_n30993, new_n30994, new_n30995, new_n30996, new_n30997, new_n30998,
    new_n30999, new_n31000, new_n31001, new_n31002, new_n31003, new_n31004,
    new_n31005, new_n31006, new_n31007, new_n31008, new_n31009, new_n31010,
    new_n31011, new_n31012, new_n31013, new_n31014, new_n31015, new_n31016,
    new_n31017, new_n31018, new_n31019, new_n31020, new_n31021, new_n31022,
    new_n31023, new_n31024, new_n31025, new_n31026, new_n31027, new_n31028,
    new_n31029, new_n31030, new_n31031, new_n31032, new_n31033, new_n31034,
    new_n31035, new_n31036, new_n31037, new_n31038, new_n31039, new_n31040,
    new_n31041, new_n31042, new_n31043, new_n31044, new_n31045, new_n31046,
    new_n31047, new_n31048, new_n31049, new_n31050, new_n31051, new_n31052,
    new_n31053, new_n31054, new_n31055, new_n31056, new_n31057, new_n31058,
    new_n31059, new_n31060, new_n31061, new_n31062, new_n31063, new_n31064,
    new_n31065, new_n31066, new_n31067, new_n31068, new_n31069, new_n31070,
    new_n31071, new_n31072, new_n31073, new_n31074, new_n31075, new_n31076,
    new_n31077, new_n31078, new_n31079, new_n31080, new_n31081, new_n31082,
    new_n31083, new_n31084, new_n31085, new_n31086, new_n31087, new_n31088,
    new_n31089, new_n31090, new_n31091, new_n31092, new_n31093, new_n31094,
    new_n31095, new_n31096, new_n31097, new_n31098, new_n31099, new_n31100,
    new_n31101, new_n31102, new_n31103, new_n31104, new_n31105, new_n31106,
    new_n31107, new_n31108, new_n31109, new_n31110, new_n31111, new_n31112,
    new_n31113, new_n31114, new_n31115, new_n31116, new_n31117, new_n31118,
    new_n31119, new_n31120, new_n31121, new_n31122, new_n31123, new_n31124,
    new_n31125, new_n31126, new_n31127, new_n31128, new_n31129, new_n31130,
    new_n31131, new_n31132, new_n31133, new_n31134, new_n31135, new_n31136,
    new_n31137, new_n31138, new_n31139, new_n31140, new_n31141, new_n31142,
    new_n31143, new_n31144, new_n31145, new_n31146, new_n31147, new_n31148,
    new_n31149, new_n31150, new_n31151, new_n31152, new_n31153, new_n31154,
    new_n31155, new_n31156, new_n31157, new_n31158, new_n31159, new_n31160,
    new_n31161, new_n31162, new_n31163, new_n31164, new_n31165, new_n31166,
    new_n31167, new_n31168, new_n31169, new_n31170, new_n31171, new_n31172,
    new_n31173, new_n31174, new_n31175, new_n31176, new_n31177, new_n31178,
    new_n31179, new_n31180, new_n31181, new_n31182, new_n31183, new_n31184,
    new_n31185, new_n31186, new_n31187, new_n31188, new_n31189, new_n31190,
    new_n31191, new_n31192, new_n31193, new_n31194, new_n31195, new_n31196,
    new_n31197, new_n31198, new_n31199, new_n31200, new_n31201, new_n31202,
    new_n31203, new_n31204, new_n31205, new_n31206, new_n31207, new_n31208,
    new_n31209, new_n31210, new_n31211, new_n31212, new_n31213, new_n31214,
    new_n31215, new_n31216, new_n31217, new_n31218, new_n31219, new_n31220,
    new_n31221, new_n31222, new_n31223, new_n31224, new_n31225, new_n31226,
    new_n31227, new_n31228, new_n31229, new_n31230, new_n31231, new_n31232,
    new_n31233, new_n31234, new_n31235, new_n31236, new_n31237, new_n31238,
    new_n31239, new_n31240, new_n31241, new_n31242, new_n31243, new_n31244,
    new_n31245, new_n31246, new_n31247, new_n31248, new_n31249, new_n31250,
    new_n31251, new_n31252, new_n31253, new_n31254, new_n31255, new_n31256,
    new_n31257, new_n31258, new_n31259, new_n31260, new_n31261, new_n31262,
    new_n31263, new_n31264, new_n31265, new_n31266, new_n31267, new_n31268,
    new_n31269, new_n31270, new_n31271, new_n31272, new_n31273, new_n31274,
    new_n31275, new_n31276, new_n31277, new_n31278, new_n31279, new_n31280,
    new_n31281, new_n31282, new_n31283, new_n31284, new_n31285, new_n31286,
    new_n31287, new_n31288, new_n31289, new_n31290, new_n31291, new_n31292,
    new_n31293, new_n31294, new_n31295, new_n31296, new_n31297, new_n31298,
    new_n31299, new_n31300, new_n31301, new_n31302, new_n31303, new_n31304,
    new_n31305, new_n31306, new_n31307, new_n31308, new_n31309, new_n31310,
    new_n31311, new_n31312, new_n31313, new_n31314, new_n31315, new_n31316,
    new_n31317, new_n31318, new_n31319, new_n31320, new_n31321, new_n31322,
    new_n31323, new_n31324, new_n31325, new_n31326, new_n31327, new_n31328,
    new_n31329, new_n31330, new_n31331, new_n31332, new_n31333, new_n31334,
    new_n31335, new_n31336, new_n31337, new_n31338, new_n31339, new_n31340,
    new_n31341, new_n31342, new_n31343, new_n31344, new_n31345, new_n31346,
    new_n31347, new_n31348, new_n31349, new_n31350, new_n31351, new_n31352,
    new_n31353, new_n31354, new_n31355, new_n31356, new_n31357, new_n31358,
    new_n31359, new_n31360, new_n31361, new_n31362, new_n31363, new_n31364,
    new_n31365, new_n31366, new_n31367, new_n31368, new_n31369, new_n31370,
    new_n31371, new_n31372, new_n31373, new_n31374, new_n31375, new_n31376,
    new_n31377, new_n31378, new_n31379, new_n31380, new_n31381, new_n31382,
    new_n31383, new_n31384, new_n31385, new_n31386, new_n31387, new_n31388,
    new_n31389, new_n31390, new_n31391, new_n31392, new_n31393, new_n31394,
    new_n31395, new_n31396, new_n31397, new_n31398, new_n31399, new_n31400,
    new_n31401, new_n31402, new_n31403, new_n31404, new_n31405, new_n31406,
    new_n31407, new_n31408, new_n31409, new_n31410, new_n31411, new_n31412,
    new_n31413, new_n31414, new_n31415, new_n31416, new_n31417, new_n31418,
    new_n31419, new_n31420, new_n31421, new_n31422, new_n31423, new_n31424,
    new_n31425, new_n31426, new_n31427, new_n31428, new_n31429, new_n31430,
    new_n31431, new_n31432, new_n31433, new_n31434, new_n31435, new_n31436,
    new_n31437, new_n31438, new_n31439, new_n31440, new_n31441, new_n31442,
    new_n31443, new_n31444, new_n31445, new_n31446, new_n31447, new_n31448,
    new_n31449, new_n31450, new_n31451, new_n31452, new_n31453, new_n31454,
    new_n31455, new_n31456, new_n31457, new_n31458, new_n31459, new_n31460,
    new_n31461, new_n31462, new_n31463, new_n31464, new_n31465, new_n31466,
    new_n31467, new_n31468, new_n31469, new_n31470, new_n31471, new_n31472,
    new_n31473, new_n31474, new_n31475, new_n31476, new_n31477, new_n31478,
    new_n31479, new_n31480, new_n31481, new_n31482, new_n31483, new_n31484,
    new_n31485, new_n31486, new_n31487, new_n31488, new_n31489, new_n31490,
    new_n31491, new_n31492, new_n31493, new_n31494, new_n31495, new_n31496,
    new_n31497, new_n31498, new_n31499, new_n31500, new_n31501, new_n31502,
    new_n31503, new_n31504, new_n31505, new_n31506, new_n31507, new_n31508,
    new_n31509, new_n31510, new_n31511, new_n31512, new_n31513, new_n31514,
    new_n31515, new_n31516, new_n31517, new_n31518, new_n31519, new_n31520,
    new_n31521, new_n31522, new_n31523, new_n31524, new_n31525, new_n31526,
    new_n31527, new_n31528, new_n31529, new_n31530, new_n31531, new_n31532,
    new_n31533, new_n31534, new_n31535, new_n31536, new_n31537, new_n31538,
    new_n31539, new_n31540, new_n31541, new_n31542, new_n31543, new_n31544,
    new_n31545, new_n31546, new_n31547, new_n31548, new_n31549, new_n31550,
    new_n31551, new_n31552, new_n31553, new_n31554, new_n31555, new_n31556,
    new_n31557, new_n31558, new_n31559, new_n31560, new_n31561, new_n31562,
    new_n31563, new_n31564, new_n31565, new_n31566, new_n31567, new_n31568,
    new_n31569, new_n31570, new_n31571, new_n31572, new_n31573, new_n31574,
    new_n31575, new_n31576, new_n31577, new_n31578, new_n31579, new_n31580,
    new_n31581, new_n31582, new_n31583, new_n31584, new_n31585, new_n31586,
    new_n31587, new_n31588, new_n31589, new_n31590, new_n31591, new_n31592,
    new_n31593, new_n31594, new_n31595, new_n31596, new_n31597, new_n31598,
    new_n31599, new_n31600, new_n31601, new_n31602, new_n31603, new_n31604,
    new_n31605, new_n31606, new_n31607, new_n31608, new_n31609, new_n31610,
    new_n31611, new_n31612, new_n31613, new_n31614, new_n31615, new_n31616,
    new_n31617, new_n31618, new_n31619, new_n31620, new_n31621, new_n31622,
    new_n31623, new_n31624, new_n31625, new_n31626, new_n31627, new_n31628,
    new_n31629, new_n31630, new_n31631, new_n31632, new_n31633, new_n31634,
    new_n31635, new_n31636, new_n31637, new_n31638, new_n31639, new_n31640,
    new_n31641, new_n31642, new_n31643, new_n31644, new_n31645, new_n31646,
    new_n31647, new_n31648, new_n31649, new_n31650, new_n31651, new_n31652,
    new_n31653, new_n31654, new_n31655, new_n31656, new_n31657, new_n31658,
    new_n31659, new_n31660, new_n31661, new_n31662, new_n31663, new_n31664,
    new_n31665, new_n31666, new_n31667, new_n31668, new_n31669, new_n31670,
    new_n31671, new_n31672, new_n31673, new_n31674, new_n31675, new_n31676,
    new_n31677, new_n31678, new_n31679, new_n31680, new_n31681, new_n31682,
    new_n31683, new_n31684, new_n31685, new_n31686, new_n31687, new_n31688,
    new_n31689, new_n31690, new_n31691, new_n31692, new_n31693, new_n31694,
    new_n31695, new_n31696, new_n31697, new_n31698, new_n31699, new_n31700,
    new_n31701, new_n31702, new_n31703, new_n31704, new_n31705, new_n31706,
    new_n31707, new_n31708, new_n31709, new_n31710, new_n31711, new_n31712,
    new_n31713, new_n31714, new_n31715, new_n31716, new_n31717, new_n31718,
    new_n31719, new_n31720, new_n31721, new_n31722, new_n31723, new_n31724,
    new_n31725, new_n31726, new_n31727, new_n31728, new_n31729, new_n31730,
    new_n31731, new_n31732, new_n31733, new_n31734, new_n31735, new_n31736,
    new_n31737, new_n31738, new_n31739, new_n31740, new_n31741, new_n31742,
    new_n31743, new_n31744, new_n31745, new_n31746, new_n31747, new_n31748,
    new_n31749, new_n31750, new_n31751, new_n31752, new_n31753, new_n31754,
    new_n31755, new_n31756, new_n31757, new_n31758, new_n31759, new_n31760,
    new_n31761, new_n31762, new_n31763, new_n31764, new_n31765, new_n31766,
    new_n31767, new_n31768, new_n31769, new_n31770, new_n31771, new_n31772,
    new_n31773, new_n31774, new_n31775, new_n31776, new_n31777, new_n31778,
    new_n31779, new_n31780, new_n31781, new_n31782, new_n31783, new_n31784,
    new_n31785, new_n31786, new_n31787, new_n31788, new_n31789, new_n31790,
    new_n31791, new_n31792, new_n31793, new_n31794, new_n31795, new_n31796,
    new_n31797, new_n31798, new_n31799, new_n31800, new_n31801, new_n31802,
    new_n31803, new_n31804, new_n31805, new_n31806, new_n31807, new_n31808,
    new_n31809, new_n31810, new_n31811, new_n31812, new_n31813, new_n31814,
    new_n31815, new_n31816, new_n31817, new_n31818, new_n31819, new_n31820,
    new_n31821, new_n31822, new_n31823, new_n31824, new_n31825, new_n31826,
    new_n31827, new_n31828, new_n31829, new_n31830, new_n31831, new_n31832,
    new_n31833, new_n31834, new_n31835, new_n31836, new_n31837, new_n31838,
    new_n31839, new_n31840, new_n31841, new_n31842, new_n31843, new_n31844,
    new_n31845, new_n31846, new_n31847, new_n31848, new_n31849, new_n31850,
    new_n31851, new_n31852, new_n31853, new_n31854, new_n31855, new_n31856,
    new_n31857, new_n31858, new_n31859, new_n31860, new_n31861, new_n31862,
    new_n31863, new_n31864, new_n31865, new_n31866, new_n31867, new_n31868,
    new_n31869, new_n31870, new_n31871, new_n31872, new_n31873, new_n31874,
    new_n31875, new_n31876, new_n31877, new_n31878, new_n31879, new_n31880,
    new_n31881, new_n31882, new_n31883, new_n31884, new_n31885, new_n31886,
    new_n31887, new_n31888, new_n31889, new_n31890, new_n31891, new_n31892,
    new_n31893, new_n31894, new_n31895, new_n31896, new_n31897, new_n31898,
    new_n31899, new_n31900, new_n31901, new_n31902, new_n31903, new_n31904,
    new_n31905, new_n31906, new_n31907, new_n31908, new_n31909, new_n31910,
    new_n31911, new_n31912, new_n31913, new_n31914, new_n31915, new_n31916,
    new_n31917, new_n31918, new_n31919, new_n31920, new_n31921, new_n31922,
    new_n31923, new_n31924, new_n31925, new_n31926, new_n31927, new_n31928,
    new_n31929, new_n31930, new_n31931, new_n31932, new_n31933, new_n31934,
    new_n31935, new_n31936, new_n31937, new_n31938, new_n31939, new_n31940,
    new_n31941, new_n31942, new_n31943, new_n31944, new_n31945, new_n31946,
    new_n31947, new_n31948, new_n31949, new_n31950, new_n31951, new_n31952,
    new_n31953, new_n31954, new_n31955, new_n31956, new_n31957, new_n31958,
    new_n31959, new_n31960, new_n31961, new_n31962, new_n31963, new_n31964,
    new_n31965, new_n31966, new_n31967, new_n31968, new_n31969, new_n31970,
    new_n31971, new_n31972, new_n31973, new_n31974, new_n31975, new_n31976,
    new_n31977, new_n31978, new_n31979, new_n31980, new_n31981, new_n31982,
    new_n31983, new_n31984, new_n31985, new_n31986, new_n31987, new_n31988,
    new_n31989, new_n31990, new_n31991, new_n31992, new_n31993, new_n31994,
    new_n31995, new_n31996, new_n31997, new_n31998, new_n31999, new_n32000,
    new_n32001, new_n32002, new_n32003, new_n32004, new_n32005, new_n32006,
    new_n32007, new_n32008, new_n32009, new_n32010, new_n32011, new_n32012,
    new_n32013, new_n32014, new_n32015, new_n32016, new_n32017, new_n32018,
    new_n32019, new_n32020, new_n32021, new_n32022, new_n32023, new_n32024,
    new_n32025, new_n32026, new_n32027, new_n32028, new_n32029, new_n32030,
    new_n32031, new_n32032, new_n32033, new_n32034, new_n32035, new_n32036,
    new_n32037, new_n32038, new_n32039, new_n32040, new_n32041, new_n32042,
    new_n32043, new_n32044, new_n32045, new_n32046, new_n32047, new_n32048,
    new_n32049, new_n32050, new_n32051, new_n32052, new_n32053, new_n32054,
    new_n32055, new_n32056, new_n32057, new_n32058, new_n32059, new_n32060,
    new_n32061, new_n32062, new_n32063, new_n32064, new_n32065, new_n32066,
    new_n32067, new_n32068, new_n32069, new_n32070, new_n32071, new_n32072,
    new_n32073, new_n32074, new_n32075, new_n32076, new_n32077, new_n32078,
    new_n32079, new_n32080, new_n32081, new_n32082, new_n32083, new_n32084,
    new_n32085, new_n32086, new_n32087, new_n32088, new_n32089, new_n32090,
    new_n32091, new_n32092, new_n32093, new_n32094, new_n32095, new_n32096,
    new_n32097, new_n32098, new_n32099, new_n32100, new_n32101, new_n32102,
    new_n32103, new_n32104, new_n32105, new_n32106, new_n32107, new_n32108,
    new_n32109, new_n32110, new_n32111, new_n32112, new_n32113, new_n32114,
    new_n32115, new_n32116, new_n32117, new_n32118, new_n32119, new_n32120,
    new_n32121, new_n32122, new_n32123, new_n32124, new_n32125, new_n32126,
    new_n32127, new_n32128, new_n32129, new_n32130, new_n32131, new_n32132,
    new_n32133, new_n32134, new_n32135, new_n32136, new_n32137, new_n32138,
    new_n32139, new_n32140, new_n32141, new_n32142, new_n32143, new_n32144,
    new_n32145, new_n32146, new_n32147, new_n32148, new_n32149, new_n32150,
    new_n32151, new_n32152, new_n32153, new_n32154, new_n32155, new_n32156,
    new_n32157, new_n32158, new_n32159, new_n32160, new_n32161, new_n32162,
    new_n32163, new_n32164, new_n32165, new_n32166, new_n32167, new_n32168,
    new_n32169, new_n32170, new_n32171, new_n32172, new_n32173, new_n32174,
    new_n32175, new_n32176, new_n32177, new_n32178, new_n32179, new_n32180,
    new_n32181, new_n32182, new_n32183, new_n32184, new_n32185, new_n32186,
    new_n32187, new_n32188, new_n32189, new_n32190, new_n32191, new_n32192,
    new_n32193, new_n32194, new_n32195, new_n32196, new_n32197, new_n32198,
    new_n32199, new_n32200, new_n32201, new_n32202, new_n32203, new_n32204,
    new_n32205, new_n32206, new_n32207, new_n32208, new_n32209, new_n32210,
    new_n32211, new_n32212, new_n32213, new_n32214, new_n32215, new_n32216,
    new_n32217, new_n32218, new_n32219, new_n32220, new_n32221, new_n32222,
    new_n32223, new_n32224, new_n32225, new_n32226, new_n32227, new_n32228,
    new_n32229, new_n32230, new_n32231, new_n32232, new_n32233, new_n32234,
    new_n32235, new_n32236, new_n32237, new_n32238, new_n32239, new_n32240,
    new_n32241, new_n32242, new_n32243, new_n32244, new_n32245, new_n32246,
    new_n32247, new_n32248, new_n32249, new_n32250, new_n32251, new_n32252,
    new_n32253, new_n32254, new_n32255, new_n32256, new_n32257, new_n32258,
    new_n32259, new_n32260, new_n32261, new_n32262, new_n32263, new_n32264,
    new_n32265, new_n32266, new_n32267, new_n32268, new_n32269, new_n32270,
    new_n32271, new_n32272, new_n32273, new_n32274, new_n32275, new_n32276,
    new_n32277, new_n32278, new_n32279, new_n32280, new_n32281, new_n32282,
    new_n32283, new_n32284, new_n32285, new_n32286, new_n32287, new_n32288,
    new_n32289, new_n32290, new_n32291, new_n32292, new_n32293, new_n32294,
    new_n32295, new_n32296, new_n32297, new_n32298, new_n32299, new_n32300,
    new_n32301, new_n32302, new_n32303, new_n32304, new_n32305, new_n32306,
    new_n32307, new_n32308, new_n32309, new_n32310, new_n32311, new_n32312,
    new_n32313, new_n32314, new_n32315, new_n32316, new_n32317, new_n32318,
    new_n32319, new_n32320, new_n32321, new_n32322, new_n32323, new_n32324,
    new_n32325, new_n32326, new_n32327, new_n32328, new_n32329, new_n32330,
    new_n32331, new_n32332, new_n32333, new_n32334, new_n32335, new_n32336,
    new_n32337, new_n32338, new_n32339, new_n32340, new_n32341, new_n32342,
    new_n32343, new_n32344, new_n32345, new_n32346, new_n32347, new_n32348,
    new_n32349, new_n32350, new_n32351, new_n32352, new_n32353, new_n32354,
    new_n32355, new_n32356, new_n32357, new_n32358, new_n32359, new_n32360,
    new_n32361, new_n32362, new_n32363, new_n32364, new_n32365, new_n32366,
    new_n32367, new_n32368, new_n32369, new_n32370, new_n32371, new_n32372,
    new_n32373, new_n32374, new_n32375, new_n32376, new_n32377, new_n32378,
    new_n32379, new_n32380, new_n32381, new_n32382, new_n32383, new_n32384,
    new_n32385, new_n32386, new_n32387, new_n32388, new_n32389, new_n32390,
    new_n32391, new_n32392, new_n32393, new_n32394, new_n32395, new_n32396,
    new_n32397, new_n32398, new_n32399, new_n32400, new_n32401, new_n32402,
    new_n32403, new_n32404, new_n32405, new_n32406, new_n32407, new_n32408,
    new_n32409, new_n32410, new_n32411, new_n32412, new_n32413, new_n32414,
    new_n32415, new_n32416, new_n32417, new_n32418, new_n32419, new_n32420,
    new_n32421, new_n32422, new_n32423, new_n32424, new_n32425, new_n32426,
    new_n32427, new_n32428, new_n32429, new_n32430, new_n32431, new_n32432,
    new_n32433, new_n32434, new_n32435, new_n32436, new_n32437, new_n32438,
    new_n32439, new_n32440, new_n32441, new_n32442, new_n32443, new_n32444,
    new_n32445, new_n32446, new_n32447, new_n32448, new_n32449, new_n32450,
    new_n32451, new_n32452, new_n32453, new_n32454, new_n32455, new_n32456,
    new_n32457, new_n32458, new_n32459, new_n32460, new_n32461, new_n32462,
    new_n32463, new_n32464, new_n32465, new_n32466, new_n32467, new_n32468,
    new_n32469, new_n32470, new_n32471, new_n32472, new_n32473, new_n32474,
    new_n32475, new_n32476, new_n32477, new_n32478, new_n32479, new_n32480,
    new_n32481, new_n32482, new_n32483, new_n32484, new_n32485, new_n32486,
    new_n32487, new_n32488, new_n32489, new_n32490, new_n32491, new_n32492,
    new_n32493, new_n32494, new_n32495, new_n32496, new_n32497, new_n32498,
    new_n32499, new_n32500, new_n32501, new_n32502, new_n32503, new_n32504,
    new_n32505, new_n32506, new_n32507, new_n32508, new_n32509, new_n32510,
    new_n32511, new_n32512, new_n32513, new_n32514, new_n32515, new_n32516,
    new_n32517, new_n32518, new_n32519, new_n32520, new_n32521, new_n32522,
    new_n32523, new_n32524, new_n32525, new_n32526, new_n32527, new_n32528,
    new_n32529, new_n32530, new_n32531, new_n32532, new_n32533, new_n32534,
    new_n32535, new_n32536, new_n32537, new_n32538, new_n32539, new_n32540,
    new_n32541, new_n32542, new_n32543, new_n32544, new_n32545, new_n32546,
    new_n32547, new_n32548, new_n32549, new_n32550, new_n32551, new_n32552,
    new_n32553, new_n32554, new_n32555, new_n32556, new_n32557, new_n32558,
    new_n32559, new_n32560, new_n32561, new_n32562, new_n32563, new_n32564,
    new_n32565, new_n32566, new_n32567, new_n32568, new_n32569, new_n32570,
    new_n32571, new_n32572, new_n32573, new_n32574, new_n32575, new_n32576,
    new_n32577, new_n32578, new_n32579, new_n32580, new_n32581, new_n32582,
    new_n32583, new_n32584, new_n32585, new_n32586, new_n32587, new_n32588,
    new_n32589, new_n32590, new_n32591, new_n32592, new_n32593, new_n32594,
    new_n32595, new_n32596, new_n32597, new_n32598, new_n32599, new_n32600,
    new_n32601, new_n32602, new_n32603, new_n32604, new_n32605, new_n32606,
    new_n32607, new_n32608, new_n32609, new_n32610, new_n32611, new_n32612,
    new_n32613, new_n32614, new_n32615, new_n32616, new_n32617, new_n32618,
    new_n32619, new_n32620, new_n32621, new_n32622, new_n32623, new_n32624,
    new_n32625, new_n32626, new_n32627, new_n32628, new_n32629, new_n32630,
    new_n32631, new_n32632, new_n32633, new_n32634, new_n32635, new_n32636,
    new_n32637, new_n32638, new_n32639, new_n32640, new_n32641, new_n32642,
    new_n32643, new_n32644, new_n32645, new_n32646, new_n32647, new_n32648,
    new_n32649, new_n32650, new_n32651, new_n32652, new_n32653, new_n32654,
    new_n32655, new_n32656, new_n32657, new_n32658, new_n32659, new_n32660,
    new_n32661, new_n32662, new_n32663, new_n32664, new_n32665, new_n32666,
    new_n32667, new_n32668, new_n32669, new_n32670, new_n32671, new_n32672,
    new_n32673, new_n32674, new_n32675, new_n32676, new_n32677, new_n32678,
    new_n32679, new_n32680, new_n32681, new_n32682, new_n32683, new_n32684,
    new_n32685, new_n32686, new_n32687, new_n32688, new_n32689, new_n32690,
    new_n32691, new_n32692, new_n32693, new_n32694, new_n32695, new_n32696,
    new_n32697, new_n32698, new_n32699, new_n32700, new_n32701, new_n32702,
    new_n32703, new_n32704, new_n32705, new_n32706, new_n32707, new_n32708,
    new_n32709, new_n32710, new_n32711, new_n32712, new_n32713, new_n32714,
    new_n32715, new_n32716, new_n32717, new_n32718, new_n32719, new_n32720,
    new_n32721, new_n32722, new_n32723, new_n32724, new_n32725, new_n32726,
    new_n32727, new_n32728, new_n32729, new_n32730, new_n32731, new_n32732,
    new_n32733, new_n32734, new_n32735, new_n32736, new_n32737, new_n32738,
    new_n32739, new_n32740, new_n32741, new_n32742, new_n32743, new_n32744,
    new_n32745, new_n32746, new_n32747, new_n32748, new_n32749, new_n32750,
    new_n32751, new_n32752, new_n32753, new_n32754, new_n32755, new_n32756,
    new_n32757, new_n32758, new_n32759, new_n32760, new_n32761, new_n32762,
    new_n32763, new_n32764, new_n32765, new_n32766, new_n32767, new_n32768,
    new_n32769, new_n32770, new_n32771, new_n32772, new_n32773, new_n32774,
    new_n32775, new_n32776, new_n32777, new_n32778, new_n32779, new_n32780,
    new_n32781, new_n32782, new_n32783, new_n32784, new_n32785, new_n32786,
    new_n32787, new_n32788, new_n32789, new_n32790, new_n32791, new_n32792,
    new_n32793, new_n32794, new_n32795, new_n32796, new_n32797, new_n32798,
    new_n32799, new_n32800, new_n32801, new_n32802, new_n32803, new_n32804,
    new_n32805, new_n32806, new_n32807, new_n32808, new_n32809, new_n32810,
    new_n32811, new_n32812, new_n32813, new_n32814, new_n32815, new_n32816,
    new_n32817, new_n32818, new_n32819, new_n32820, new_n32821, new_n32822,
    new_n32823, new_n32824, new_n32825, new_n32826, new_n32827, new_n32828,
    new_n32829, new_n32830, new_n32831, new_n32832, new_n32833, new_n32834,
    new_n32835, new_n32836, new_n32837, new_n32838, new_n32839, new_n32840,
    new_n32841, new_n32842, new_n32843, new_n32844, new_n32845, new_n32846,
    new_n32847, new_n32848, new_n32849, new_n32850, new_n32851, new_n32852,
    new_n32853, new_n32854, new_n32855, new_n32856, new_n32857, new_n32858,
    new_n32859, new_n32860, new_n32861, new_n32862, new_n32863, new_n32864,
    new_n32865, new_n32866, new_n32867, new_n32868, new_n32869, new_n32870,
    new_n32871, new_n32872, new_n32873, new_n32874, new_n32875, new_n32876,
    new_n32877, new_n32878, new_n32879, new_n32880, new_n32881, new_n32882,
    new_n32883, new_n32884, new_n32885, new_n32886, new_n32887, new_n32888,
    new_n32889, new_n32890, new_n32891, new_n32892, new_n32893, new_n32894,
    new_n32895, new_n32896, new_n32897, new_n32898, new_n32899, new_n32900,
    new_n32901, new_n32902, new_n32903, new_n32904, new_n32905, new_n32906,
    new_n32907, new_n32908, new_n32909, new_n32910, new_n32911, new_n32912,
    new_n32913, new_n32914, new_n32915, new_n32916, new_n32917, new_n32918,
    new_n32919, new_n32920, new_n32921, new_n32922, new_n32923, new_n32924,
    new_n32925, new_n32926, new_n32927, new_n32928, new_n32929, new_n32930,
    new_n32931, new_n32932, new_n32933, new_n32934, new_n32935, new_n32936,
    new_n32937, new_n32938, new_n32939, new_n32940, new_n32941, new_n32942,
    new_n32943, new_n32944, new_n32945, new_n32946, new_n32947, new_n32948,
    new_n32949, new_n32950, new_n32951, new_n32952, new_n32953, new_n32954,
    new_n32955, new_n32956, new_n32957, new_n32958, new_n32959, new_n32960,
    new_n32961, new_n32962, new_n32963, new_n32964, new_n32965, new_n32966,
    new_n32967, new_n32968, new_n32969, new_n32970, new_n32971, new_n32972,
    new_n32973, new_n32974, new_n32975, new_n32976, new_n32977, new_n32978,
    new_n32979, new_n32980, new_n32981, new_n32982, new_n32983, new_n32984,
    new_n32985, new_n32986, new_n32987, new_n32988, new_n32989, new_n32990,
    new_n32991, new_n32992, new_n32993, new_n32994, new_n32995, new_n32996,
    new_n32997, new_n32998, new_n32999, new_n33000, new_n33001, new_n33002,
    new_n33003, new_n33004, new_n33005, new_n33006, new_n33007, new_n33008,
    new_n33009, new_n33010, new_n33011, new_n33012, new_n33013, new_n33014,
    new_n33015, new_n33016, new_n33017, new_n33018, new_n33019, new_n33020,
    new_n33021, new_n33022, new_n33023, new_n33024, new_n33025, new_n33026,
    new_n33027, new_n33028, new_n33029, new_n33030, new_n33031, new_n33032,
    new_n33033, new_n33034, new_n33035, new_n33036, new_n33037, new_n33038,
    new_n33039, new_n33040, new_n33041, new_n33042, new_n33043, new_n33044,
    new_n33045, new_n33046, new_n33047, new_n33048, new_n33049, new_n33050,
    new_n33051, new_n33052, new_n33053, new_n33054, new_n33055, new_n33056,
    new_n33057, new_n33058, new_n33059, new_n33060, new_n33061, new_n33062,
    new_n33063, new_n33064, new_n33065, new_n33066, new_n33067, new_n33068,
    new_n33069, new_n33070, new_n33071, new_n33072, new_n33073, new_n33074,
    new_n33075, new_n33076, new_n33077, new_n33078, new_n33079, new_n33080,
    new_n33081, new_n33082, new_n33083, new_n33084, new_n33085, new_n33086,
    new_n33087, new_n33088, new_n33089, new_n33090, new_n33091, new_n33092,
    new_n33093, new_n33094, new_n33095, new_n33096, new_n33097, new_n33098,
    new_n33099, new_n33100, new_n33101, new_n33102, new_n33103, new_n33104,
    new_n33105, new_n33106, new_n33107, new_n33108, new_n33109, new_n33110,
    new_n33111, new_n33112, new_n33113, new_n33114, new_n33115, new_n33116,
    new_n33117, new_n33118, new_n33119, new_n33120, new_n33121, new_n33122,
    new_n33123, new_n33124, new_n33125, new_n33126, new_n33127, new_n33128,
    new_n33129, new_n33130, new_n33131, new_n33132, new_n33133, new_n33134,
    new_n33135, new_n33136, new_n33137, new_n33138, new_n33139, new_n33140,
    new_n33141, new_n33142, new_n33143, new_n33144, new_n33145, new_n33146,
    new_n33147, new_n33148, new_n33149, new_n33150, new_n33151, new_n33152,
    new_n33153, new_n33154, new_n33155, new_n33156, new_n33157, new_n33158,
    new_n33159, new_n33160, new_n33161, new_n33162, new_n33163, new_n33164,
    new_n33165, new_n33166, new_n33167, new_n33168, new_n33169, new_n33170,
    new_n33171, new_n33172, new_n33173, new_n33174, new_n33175, new_n33176,
    new_n33177, new_n33178, new_n33179, new_n33180, new_n33181, new_n33182,
    new_n33183, new_n33184, new_n33185, new_n33186, new_n33187, new_n33188,
    new_n33189, new_n33190, new_n33191, new_n33192, new_n33193, new_n33194,
    new_n33195, new_n33196, new_n33197, new_n33198, new_n33199, new_n33200,
    new_n33201, new_n33202, new_n33203, new_n33204, new_n33205, new_n33206,
    new_n33207, new_n33208, new_n33209, new_n33210, new_n33211, new_n33212,
    new_n33213, new_n33214, new_n33215, new_n33216, new_n33217, new_n33218,
    new_n33219, new_n33220, new_n33221, new_n33222, new_n33223, new_n33224,
    new_n33225, new_n33226, new_n33227, new_n33228, new_n33229, new_n33230,
    new_n33231, new_n33232, new_n33233, new_n33234, new_n33235, new_n33236,
    new_n33237, new_n33238, new_n33239, new_n33240, new_n33241, new_n33242,
    new_n33243, new_n33244, new_n33245, new_n33246, new_n33247, new_n33248,
    new_n33249, new_n33250, new_n33251, new_n33252, new_n33253, new_n33254,
    new_n33255, new_n33256, new_n33257, new_n33258, new_n33259, new_n33260,
    new_n33261, new_n33262, new_n33263, new_n33264, new_n33265, new_n33266,
    new_n33267, new_n33268, new_n33269, new_n33270, new_n33271, new_n33272,
    new_n33273, new_n33274, new_n33275, new_n33276, new_n33277, new_n33278,
    new_n33279, new_n33280, new_n33281, new_n33282, new_n33283, new_n33284,
    new_n33285, new_n33286, new_n33287, new_n33288, new_n33289, new_n33290,
    new_n33291, new_n33292, new_n33293, new_n33294, new_n33295, new_n33296,
    new_n33297, new_n33298, new_n33299, new_n33300, new_n33301, new_n33302,
    new_n33303, new_n33304, new_n33305, new_n33306, new_n33307, new_n33308,
    new_n33309, new_n33310, new_n33311, new_n33312, new_n33313, new_n33314,
    new_n33315, new_n33316, new_n33317, new_n33318, new_n33319, new_n33320,
    new_n33321, new_n33322, new_n33323, new_n33324, new_n33325, new_n33326,
    new_n33327, new_n33328, new_n33329, new_n33330, new_n33331, new_n33332,
    new_n33333, new_n33334, new_n33335, new_n33336, new_n33337, new_n33338,
    new_n33339, new_n33340, new_n33341, new_n33342, new_n33343, new_n33344,
    new_n33345, new_n33346, new_n33347, new_n33348, new_n33349, new_n33350,
    new_n33351, new_n33352, new_n33353, new_n33354, new_n33355, new_n33356,
    new_n33357, new_n33358, new_n33359, new_n33360, new_n33361, new_n33362,
    new_n33363, new_n33364, new_n33365, new_n33366, new_n33367, new_n33368,
    new_n33369, new_n33370, new_n33371, new_n33372, new_n33373, new_n33374,
    new_n33375, new_n33376, new_n33377, new_n33378, new_n33379, new_n33380,
    new_n33381, new_n33382, new_n33383, new_n33384, new_n33385, new_n33386,
    new_n33387, new_n33388, new_n33389, new_n33390, new_n33391, new_n33392,
    new_n33393, new_n33394, new_n33395, new_n33396, new_n33397, new_n33398,
    new_n33399, new_n33400, new_n33401, new_n33402, new_n33403, new_n33404,
    new_n33405, new_n33406, new_n33407, new_n33408, new_n33409, new_n33410,
    new_n33411, new_n33412, new_n33413, new_n33414, new_n33415, new_n33416,
    new_n33417, new_n33418, new_n33419, new_n33420, new_n33421, new_n33422,
    new_n33423, new_n33424, new_n33425, new_n33426, new_n33427, new_n33428,
    new_n33429, new_n33430, new_n33431, new_n33432, new_n33433, new_n33434,
    new_n33435, new_n33436, new_n33437, new_n33438, new_n33439, new_n33440,
    new_n33441, new_n33442, new_n33443, new_n33444, new_n33445, new_n33446,
    new_n33447, new_n33448, new_n33449, new_n33450, new_n33451, new_n33452,
    new_n33453, new_n33454, new_n33455, new_n33456, new_n33457, new_n33458,
    new_n33459, new_n33460, new_n33461, new_n33462, new_n33463, new_n33464,
    new_n33465, new_n33466, new_n33467, new_n33468, new_n33469, new_n33470,
    new_n33471, new_n33472, new_n33473, new_n33474, new_n33475, new_n33476,
    new_n33477, new_n33478, new_n33479, new_n33480, new_n33481, new_n33482,
    new_n33483, new_n33484, new_n33485, new_n33486, new_n33487, new_n33488,
    new_n33489, new_n33490, new_n33491, new_n33492, new_n33493, new_n33494,
    new_n33495, new_n33496, new_n33497, new_n33498, new_n33499, new_n33500,
    new_n33501, new_n33502, new_n33503, new_n33504, new_n33505, new_n33506,
    new_n33507, new_n33508, new_n33509, new_n33510, new_n33511, new_n33512,
    new_n33513, new_n33514, new_n33515, new_n33516, new_n33517, new_n33518,
    new_n33519, new_n33520, new_n33521, new_n33522, new_n33523, new_n33524,
    new_n33525, new_n33526, new_n33527, new_n33528, new_n33529, new_n33530,
    new_n33531, new_n33532, new_n33533, new_n33534, new_n33535, new_n33536,
    new_n33537, new_n33538, new_n33539, new_n33540, new_n33541, new_n33542,
    new_n33543, new_n33544, new_n33545, new_n33546, new_n33547, new_n33548,
    new_n33549, new_n33550, new_n33551, new_n33552, new_n33553, new_n33554,
    new_n33555, new_n33556, new_n33557, new_n33558, new_n33559, new_n33560,
    new_n33561, new_n33562, new_n33563, new_n33564, new_n33565, new_n33566,
    new_n33567, new_n33568, new_n33569, new_n33570, new_n33571, new_n33572,
    new_n33573, new_n33574, new_n33575, new_n33576, new_n33577, new_n33578,
    new_n33579, new_n33580, new_n33581, new_n33582, new_n33583, new_n33584,
    new_n33585, new_n33586, new_n33587, new_n33588, new_n33589, new_n33590,
    new_n33591, new_n33592, new_n33593, new_n33594, new_n33595, new_n33596,
    new_n33597, new_n33598, new_n33599, new_n33600, new_n33601, new_n33602,
    new_n33603, new_n33604, new_n33605, new_n33606, new_n33607, new_n33608,
    new_n33609, new_n33610, new_n33611, new_n33612, new_n33613, new_n33614,
    new_n33615, new_n33616, new_n33617, new_n33618, new_n33619, new_n33620,
    new_n33621, new_n33622, new_n33623, new_n33624, new_n33625, new_n33626,
    new_n33627, new_n33628, new_n33629, new_n33630, new_n33631, new_n33632,
    new_n33633, new_n33634, new_n33635, new_n33636, new_n33637, new_n33638,
    new_n33639, new_n33640, new_n33641, new_n33642, new_n33643, new_n33644,
    new_n33645, new_n33646, new_n33647, new_n33648, new_n33649, new_n33650,
    new_n33651, new_n33652, new_n33653, new_n33654, new_n33655, new_n33656,
    new_n33657, new_n33658, new_n33659, new_n33660, new_n33661, new_n33662,
    new_n33663, new_n33664, new_n33665, new_n33666, new_n33667, new_n33668,
    new_n33669, new_n33670, new_n33671, new_n33672, new_n33673, new_n33674,
    new_n33675, new_n33676, new_n33677, new_n33678, new_n33679, new_n33680,
    new_n33681, new_n33682, new_n33683, new_n33684, new_n33685, new_n33686,
    new_n33687, new_n33688, new_n33689, new_n33690, new_n33691, new_n33692,
    new_n33693, new_n33694, new_n33695, new_n33696, new_n33697, new_n33698,
    new_n33699, new_n33700, new_n33701, new_n33702, new_n33703, new_n33704,
    new_n33705, new_n33706, new_n33707, new_n33708, new_n33709, new_n33710,
    new_n33711, new_n33712, new_n33713, new_n33714, new_n33715, new_n33716,
    new_n33717, new_n33718, new_n33719, new_n33720, new_n33721, new_n33722,
    new_n33723, new_n33724, new_n33725, new_n33726, new_n33727, new_n33728,
    new_n33729, new_n33730, new_n33731, new_n33732, new_n33733, new_n33734,
    new_n33735, new_n33736, new_n33737, new_n33738, new_n33739, new_n33740,
    new_n33741, new_n33742, new_n33743, new_n33744, new_n33745, new_n33746,
    new_n33747, new_n33748, new_n33749, new_n33750, new_n33751, new_n33752,
    new_n33753, new_n33754, new_n33755, new_n33756, new_n33757, new_n33758,
    new_n33759, new_n33760, new_n33761, new_n33762, new_n33763, new_n33764,
    new_n33765, new_n33766, new_n33767, new_n33768, new_n33769, new_n33770,
    new_n33771, new_n33772, new_n33773, new_n33774, new_n33775, new_n33776,
    new_n33777, new_n33778, new_n33779, new_n33780, new_n33781, new_n33782,
    new_n33783, new_n33784, new_n33785, new_n33786, new_n33787, new_n33788,
    new_n33789, new_n33790, new_n33791, new_n33792, new_n33793, new_n33794,
    new_n33795, new_n33796, new_n33797, new_n33798, new_n33799, new_n33800,
    new_n33801, new_n33802, new_n33803, new_n33804, new_n33805, new_n33806,
    new_n33807, new_n33808, new_n33809, new_n33810, new_n33811, new_n33812,
    new_n33813, new_n33814, new_n33815, new_n33816, new_n33817, new_n33818,
    new_n33819, new_n33820, new_n33821, new_n33822, new_n33823, new_n33824,
    new_n33825, new_n33826, new_n33827, new_n33828, new_n33829, new_n33830,
    new_n33831, new_n33832, new_n33833, new_n33834, new_n33835, new_n33836,
    new_n33837, new_n33838, new_n33839, new_n33840, new_n33841, new_n33842,
    new_n33843, new_n33844, new_n33845, new_n33846, new_n33847, new_n33848,
    new_n33849, new_n33850, new_n33851, new_n33852, new_n33853, new_n33854,
    new_n33855, new_n33856, new_n33857, new_n33858, new_n33859, new_n33860,
    new_n33861, new_n33862, new_n33863, new_n33864, new_n33865, new_n33866,
    new_n33867, new_n33868, new_n33869, new_n33870, new_n33871, new_n33872,
    new_n33873, new_n33874, new_n33875, new_n33876, new_n33877, new_n33878,
    new_n33879, new_n33880, new_n33881, new_n33882, new_n33883, new_n33884,
    new_n33885, new_n33886, new_n33887, new_n33888, new_n33889, new_n33890,
    new_n33891, new_n33892, new_n33893, new_n33894, new_n33895, new_n33896,
    new_n33897, new_n33898, new_n33899, new_n33900, new_n33901, new_n33902,
    new_n33903, new_n33904, new_n33905, new_n33906, new_n33907, new_n33908,
    new_n33909, new_n33910, new_n33911, new_n33912, new_n33913, new_n33914,
    new_n33915, new_n33916, new_n33917, new_n33918, new_n33919, new_n33920,
    new_n33921, new_n33922, new_n33923, new_n33924, new_n33925, new_n33926,
    new_n33927, new_n33928, new_n33929, new_n33930, new_n33931, new_n33932,
    new_n33933, new_n33934, new_n33935, new_n33936, new_n33937, new_n33938,
    new_n33939, new_n33940, new_n33941, new_n33942, new_n33943, new_n33944,
    new_n33945, new_n33946, new_n33947, new_n33948, new_n33949, new_n33950,
    new_n33951, new_n33952, new_n33953, new_n33954, new_n33955, new_n33956,
    new_n33957, new_n33958, new_n33959, new_n33960, new_n33961, new_n33962,
    new_n33963, new_n33964, new_n33965, new_n33966, new_n33967, new_n33968,
    new_n33969, new_n33970, new_n33971, new_n33972, new_n33973, new_n33974,
    new_n33975, new_n33976, new_n33977, new_n33978, new_n33979, new_n33980,
    new_n33981, new_n33982, new_n33983, new_n33984, new_n33985, new_n33986,
    new_n33987, new_n33988, new_n33989, new_n33990, new_n33991, new_n33992,
    new_n33993, new_n33994, new_n33995, new_n33996, new_n33997, new_n33998,
    new_n33999, new_n34000, new_n34001, new_n34002, new_n34003, new_n34004,
    new_n34005, new_n34006, new_n34007, new_n34008, new_n34009, new_n34010,
    new_n34011, new_n34012, new_n34013, new_n34014, new_n34015, new_n34016,
    new_n34017, new_n34018, new_n34019, new_n34020, new_n34021, new_n34022,
    new_n34023, new_n34024, new_n34025, new_n34026, new_n34027, new_n34028,
    new_n34029, new_n34030, new_n34031, new_n34032, new_n34033, new_n34034,
    new_n34035, new_n34036, new_n34037, new_n34038, new_n34039, new_n34040,
    new_n34041, new_n34042, new_n34043, new_n34044, new_n34045, new_n34046,
    new_n34047, new_n34048, new_n34049, new_n34050, new_n34051, new_n34052,
    new_n34053, new_n34054, new_n34055, new_n34056, new_n34057, new_n34058,
    new_n34059, new_n34060, new_n34061, new_n34062, new_n34063, new_n34064,
    new_n34065, new_n34066, new_n34067, new_n34068, new_n34069, new_n34070,
    new_n34071, new_n34072, new_n34073, new_n34074, new_n34075, new_n34076,
    new_n34077, new_n34078, new_n34079, new_n34080, new_n34081, new_n34082,
    new_n34083, new_n34084, new_n34085, new_n34086, new_n34087, new_n34088,
    new_n34089, new_n34090, new_n34091, new_n34092, new_n34093, new_n34094,
    new_n34095, new_n34096, new_n34097, new_n34098, new_n34099, new_n34100,
    new_n34101, new_n34102, new_n34103, new_n34104, new_n34105, new_n34106,
    new_n34107, new_n34108, new_n34109, new_n34110, new_n34111, new_n34112,
    new_n34113, new_n34114, new_n34115, new_n34116, new_n34117, new_n34118,
    new_n34119, new_n34120, new_n34121, new_n34122, new_n34123, new_n34124,
    new_n34125, new_n34126, new_n34127, new_n34128, new_n34129, new_n34130,
    new_n34131, new_n34132, new_n34133, new_n34134, new_n34135, new_n34136,
    new_n34137, new_n34138, new_n34139, new_n34140, new_n34141, new_n34142,
    new_n34143, new_n34144, new_n34145, new_n34146, new_n34147, new_n34148,
    new_n34149, new_n34150, new_n34151, new_n34152, new_n34153, new_n34154,
    new_n34155, new_n34156, new_n34157, new_n34158, new_n34159, new_n34160,
    new_n34161, new_n34162, new_n34163, new_n34164, new_n34165, new_n34166,
    new_n34167, new_n34168, new_n34169, new_n34170, new_n34171, new_n34172,
    new_n34173, new_n34174, new_n34175, new_n34176, new_n34177, new_n34178,
    new_n34179, new_n34180, new_n34181, new_n34182, new_n34183, new_n34184,
    new_n34185, new_n34186, new_n34187, new_n34188, new_n34189, new_n34190,
    new_n34191, new_n34192, new_n34193, new_n34194, new_n34195, new_n34196,
    new_n34197, new_n34198, new_n34199, new_n34200, new_n34201, new_n34202,
    new_n34203, new_n34204, new_n34205, new_n34206, new_n34207, new_n34208,
    new_n34209, new_n34210, new_n34211, new_n34212, new_n34213, new_n34214,
    new_n34215, new_n34216, new_n34217, new_n34218, new_n34219, new_n34220,
    new_n34221, new_n34222, new_n34223, new_n34224, new_n34225, new_n34226,
    new_n34227, new_n34228, new_n34229, new_n34230, new_n34231, new_n34232,
    new_n34233, new_n34234, new_n34235, new_n34236, new_n34237, new_n34238,
    new_n34239, new_n34240, new_n34241, new_n34242, new_n34243, new_n34244,
    new_n34245, new_n34246, new_n34247, new_n34248, new_n34249, new_n34250,
    new_n34251, new_n34252, new_n34253, new_n34254, new_n34255, new_n34256,
    new_n34257, new_n34258, new_n34259, new_n34260, new_n34261, new_n34262,
    new_n34263, new_n34264, new_n34265, new_n34266, new_n34267, new_n34268,
    new_n34269, new_n34270, new_n34271, new_n34272, new_n34273, new_n34274,
    new_n34275, new_n34276, new_n34277, new_n34278, new_n34279, new_n34280,
    new_n34281, new_n34282, new_n34283, new_n34284, new_n34285, new_n34286,
    new_n34287, new_n34288, new_n34289, new_n34290, new_n34291, new_n34292,
    new_n34293, new_n34294, new_n34295, new_n34296, new_n34297, new_n34298,
    new_n34299, new_n34300, new_n34301, new_n34302, new_n34303, new_n34304,
    new_n34305, new_n34306, new_n34307, new_n34308, new_n34309, new_n34310,
    new_n34311, new_n34312, new_n34313, new_n34314, new_n34315, new_n34316,
    new_n34317, new_n34318, new_n34319, new_n34320, new_n34321, new_n34322,
    new_n34323, new_n34324, new_n34325, new_n34326, new_n34327, new_n34328,
    new_n34329, new_n34330, new_n34331, new_n34332, new_n34333, new_n34334,
    new_n34335, new_n34336, new_n34337, new_n34338, new_n34339, new_n34340,
    new_n34341, new_n34342, new_n34343, new_n34344, new_n34345, new_n34346,
    new_n34347, new_n34348, new_n34349, new_n34350, new_n34351, new_n34352,
    new_n34353, new_n34354, new_n34355, new_n34356, new_n34357, new_n34358,
    new_n34359, new_n34360, new_n34361, new_n34362, new_n34363, new_n34364,
    new_n34365, new_n34366, new_n34367, new_n34368, new_n34369, new_n34370,
    new_n34371, new_n34372, new_n34373, new_n34374, new_n34375, new_n34376,
    new_n34377, new_n34378, new_n34379, new_n34380, new_n34381, new_n34382,
    new_n34383, new_n34384, new_n34385, new_n34386, new_n34387, new_n34388,
    new_n34389, new_n34390, new_n34391, new_n34392, new_n34393, new_n34394,
    new_n34395, new_n34396, new_n34397, new_n34398, new_n34399, new_n34400,
    new_n34401, new_n34402, new_n34403, new_n34404, new_n34405, new_n34406,
    new_n34407, new_n34408, new_n34409, new_n34410, new_n34411, new_n34412,
    new_n34413, new_n34414, new_n34415, new_n34416, new_n34417, new_n34418,
    new_n34419, new_n34420, new_n34421, new_n34422, new_n34423, new_n34424,
    new_n34425, new_n34426, new_n34427, new_n34428, new_n34429, new_n34430,
    new_n34431, new_n34432, new_n34433, new_n34434, new_n34435, new_n34436,
    new_n34437, new_n34438, new_n34439, new_n34440, new_n34441, new_n34442,
    new_n34443, new_n34444, new_n34445, new_n34446, new_n34447, new_n34448,
    new_n34449, new_n34450, new_n34451, new_n34452, new_n34453, new_n34454,
    new_n34455, new_n34456, new_n34457, new_n34458, new_n34459, new_n34460,
    new_n34461, new_n34462, new_n34463, new_n34464, new_n34465, new_n34466,
    new_n34467, new_n34468, new_n34469, new_n34470, new_n34471, new_n34472,
    new_n34473, new_n34474, new_n34475, new_n34476, new_n34477, new_n34478,
    new_n34479, new_n34480, new_n34481, new_n34482, new_n34483, new_n34484,
    new_n34485, new_n34486, new_n34487, new_n34488, new_n34489, new_n34490,
    new_n34491, new_n34492, new_n34493, new_n34494, new_n34495, new_n34496,
    new_n34497, new_n34498, new_n34499, new_n34500, new_n34501, new_n34502,
    new_n34503, new_n34504, new_n34505, new_n34506, new_n34507, new_n34508,
    new_n34509, new_n34510, new_n34511, new_n34512, new_n34513, new_n34514,
    new_n34515, new_n34516, new_n34517, new_n34518, new_n34519, new_n34520,
    new_n34521, new_n34522, new_n34523, new_n34524, new_n34525, new_n34526,
    new_n34527, new_n34528, new_n34529, new_n34530, new_n34531, new_n34532,
    new_n34533, new_n34534, new_n34535, new_n34536, new_n34537, new_n34538,
    new_n34539, new_n34540, new_n34541, new_n34542, new_n34543, new_n34544,
    new_n34545, new_n34546, new_n34547, new_n34548, new_n34549, new_n34550,
    new_n34551, new_n34552, new_n34553, new_n34554, new_n34555, new_n34556,
    new_n34557, new_n34558, new_n34559, new_n34560, new_n34561, new_n34562,
    new_n34563, new_n34564, new_n34565, new_n34566, new_n34567, new_n34568,
    new_n34569, new_n34570, new_n34571, new_n34572, new_n34573, new_n34574,
    new_n34575, new_n34576, new_n34577, new_n34578, new_n34579, new_n34580,
    new_n34581, new_n34582, new_n34583, new_n34584, new_n34585, new_n34586,
    new_n34587, new_n34588, new_n34589, new_n34590, new_n34591, new_n34592,
    new_n34593, new_n34594, new_n34595, new_n34596, new_n34597, new_n34598,
    new_n34599, new_n34600, new_n34601, new_n34602, new_n34603, new_n34604,
    new_n34605, new_n34606, new_n34607, new_n34608, new_n34609, new_n34610,
    new_n34611, new_n34612, new_n34613, new_n34614, new_n34615, new_n34616,
    new_n34617, new_n34618, new_n34619, new_n34620, new_n34621, new_n34622,
    new_n34623, new_n34624, new_n34625, new_n34626, new_n34627, new_n34628,
    new_n34629, new_n34630, new_n34631, new_n34632, new_n34633, new_n34634,
    new_n34635, new_n34636, new_n34637, new_n34638, new_n34639, new_n34640,
    new_n34641, new_n34642, new_n34643, new_n34644, new_n34645, new_n34646,
    new_n34647, new_n34648, new_n34649, new_n34650, new_n34651, new_n34652,
    new_n34653, new_n34654, new_n34655, new_n34656, new_n34657, new_n34658,
    new_n34659, new_n34660, new_n34661, new_n34662, new_n34663, new_n34664,
    new_n34665, new_n34666, new_n34667, new_n34668, new_n34669, new_n34670,
    new_n34671, new_n34672, new_n34673, new_n34674, new_n34675, new_n34676,
    new_n34677, new_n34678, new_n34679, new_n34680, new_n34681, new_n34682,
    new_n34683, new_n34684, new_n34685, new_n34686, new_n34687, new_n34688,
    new_n34689, new_n34690, new_n34691, new_n34692, new_n34693, new_n34694,
    new_n34695, new_n34696, new_n34697, new_n34698, new_n34699, new_n34700,
    new_n34701, new_n34702, new_n34703, new_n34704, new_n34705, new_n34706,
    new_n34707, new_n34708, new_n34709, new_n34710, new_n34711, new_n34712,
    new_n34713, new_n34714, new_n34715, new_n34716, new_n34717, new_n34718,
    new_n34719, new_n34720, new_n34721, new_n34722, new_n34723, new_n34724,
    new_n34725, new_n34726, new_n34727, new_n34728, new_n34729, new_n34730,
    new_n34731, new_n34732, new_n34733, new_n34734, new_n34735, new_n34736,
    new_n34737, new_n34738, new_n34739, new_n34740, new_n34741, new_n34742,
    new_n34743, new_n34744, new_n34745, new_n34746, new_n34747, new_n34748,
    new_n34749, new_n34750, new_n34751, new_n34752, new_n34753, new_n34754,
    new_n34755, new_n34756, new_n34757, new_n34758, new_n34759, new_n34760,
    new_n34761, new_n34762, new_n34763, new_n34764, new_n34765, new_n34766,
    new_n34767, new_n34768, new_n34769, new_n34770, new_n34771, new_n34772,
    new_n34773, new_n34774, new_n34775, new_n34776, new_n34777, new_n34778,
    new_n34779, new_n34780, new_n34781, new_n34782, new_n34783, new_n34784,
    new_n34785, new_n34786, new_n34787, new_n34788, new_n34789, new_n34790,
    new_n34791, new_n34792, new_n34793, new_n34794, new_n34795, new_n34796,
    new_n34797, new_n34798, new_n34799, new_n34800, new_n34801, new_n34802,
    new_n34803, new_n34804, new_n34805, new_n34806, new_n34807, new_n34808,
    new_n34809, new_n34810, new_n34811, new_n34812, new_n34813, new_n34814,
    new_n34815, new_n34816, new_n34817, new_n34818, new_n34819, new_n34820,
    new_n34821, new_n34822, new_n34823, new_n34824, new_n34825, new_n34826,
    new_n34827, new_n34828, new_n34829, new_n34830, new_n34831, new_n34832,
    new_n34833, new_n34834, new_n34835, new_n34836, new_n34837, new_n34838,
    new_n34839, new_n34840, new_n34841, new_n34842, new_n34843, new_n34844,
    new_n34845, new_n34846, new_n34847, new_n34848, new_n34849, new_n34850,
    new_n34851, new_n34852, new_n34853, new_n34854, new_n34855, new_n34856,
    new_n34857, new_n34858, new_n34859, new_n34860, new_n34861, new_n34862,
    new_n34863, new_n34864, new_n34865, new_n34866, new_n34867, new_n34868,
    new_n34869, new_n34870, new_n34871, new_n34872, new_n34873, new_n34874,
    new_n34875, new_n34876, new_n34877, new_n34878, new_n34879, new_n34880,
    new_n34881, new_n34882, new_n34883, new_n34884, new_n34885, new_n34886,
    new_n34887, new_n34888, new_n34889, new_n34890, new_n34891, new_n34892,
    new_n34893, new_n34894, new_n34895, new_n34896, new_n34897, new_n34898,
    new_n34899, new_n34900, new_n34901, new_n34902, new_n34903, new_n34904,
    new_n34905, new_n34906, new_n34907, new_n34908, new_n34909, new_n34910,
    new_n34911, new_n34912, new_n34913, new_n34914, new_n34915, new_n34916,
    new_n34917, new_n34918, new_n34919, new_n34920, new_n34921, new_n34922,
    new_n34923, new_n34924, new_n34925, new_n34926, new_n34927, new_n34928,
    new_n34929, new_n34930, new_n34931, new_n34932, new_n34933, new_n34934,
    new_n34935, new_n34936, new_n34937, new_n34938, new_n34939, new_n34940,
    new_n34941, new_n34942, new_n34943, new_n34944, new_n34945, new_n34946,
    new_n34947, new_n34948, new_n34949, new_n34950, new_n34951, new_n34952,
    new_n34953, new_n34954, new_n34955, new_n34956, new_n34957, new_n34958,
    new_n34959, new_n34960, new_n34961, new_n34962, new_n34963, new_n34964,
    new_n34965, new_n34966, new_n34967, new_n34968, new_n34969, new_n34970,
    new_n34971, new_n34972, new_n34973, new_n34974, new_n34975, new_n34976,
    new_n34977, new_n34978, new_n34979, new_n34980, new_n34981, new_n34982,
    new_n34983, new_n34984, new_n34985, new_n34986, new_n34987, new_n34988,
    new_n34989, new_n34990, new_n34991, new_n34992, new_n34993, new_n34994,
    new_n34995, new_n34996, new_n34997, new_n34998, new_n34999, new_n35000,
    new_n35001, new_n35002, new_n35003, new_n35004, new_n35005, new_n35006,
    new_n35007, new_n35008, new_n35009, new_n35010, new_n35011, new_n35012,
    new_n35013, new_n35014, new_n35015, new_n35016, new_n35017, new_n35018,
    new_n35019, new_n35020, new_n35021, new_n35022, new_n35023, new_n35024,
    new_n35025, new_n35026, new_n35027, new_n35028, new_n35029, new_n35030,
    new_n35031, new_n35032, new_n35033, new_n35034, new_n35035, new_n35036,
    new_n35037, new_n35038, new_n35039, new_n35040, new_n35041, new_n35042,
    new_n35043, new_n35044, new_n35045, new_n35046, new_n35047, new_n35048,
    new_n35049, new_n35050, new_n35051, new_n35052, new_n35053, new_n35054,
    new_n35055, new_n35056, new_n35057, new_n35058, new_n35059, new_n35060,
    new_n35061, new_n35062, new_n35063, new_n35064, new_n35065, new_n35066,
    new_n35067, new_n35068, new_n35069, new_n35070, new_n35071, new_n35072,
    new_n35073, new_n35074, new_n35075, new_n35076, new_n35077, new_n35078,
    new_n35079, new_n35080, new_n35081, new_n35082, new_n35083, new_n35084,
    new_n35085, new_n35086, new_n35087, new_n35088, new_n35089, new_n35090,
    new_n35091, new_n35092, new_n35093, new_n35094, new_n35095, new_n35096,
    new_n35097, new_n35098, new_n35099, new_n35100, new_n35101, new_n35102,
    new_n35103, new_n35104, new_n35105, new_n35106, new_n35107, new_n35108,
    new_n35109, new_n35110, new_n35111, new_n35112, new_n35113, new_n35114,
    new_n35115, new_n35116, new_n35117, new_n35118, new_n35119, new_n35120,
    new_n35121, new_n35122, new_n35123, new_n35124, new_n35125, new_n35126,
    new_n35127, new_n35128, new_n35129, new_n35130, new_n35131, new_n35132,
    new_n35133, new_n35134, new_n35135, new_n35136, new_n35137, new_n35138,
    new_n35139, new_n35140, new_n35141, new_n35142, new_n35143, new_n35144,
    new_n35145, new_n35146, new_n35147, new_n35148, new_n35149, new_n35150,
    new_n35151, new_n35152, new_n35153, new_n35154, new_n35155, new_n35156,
    new_n35157, new_n35158, new_n35159, new_n35160, new_n35161, new_n35162,
    new_n35163, new_n35164, new_n35165, new_n35166, new_n35167, new_n35168,
    new_n35169, new_n35170, new_n35171, new_n35172, new_n35173, new_n35174,
    new_n35175, new_n35176, new_n35177, new_n35178, new_n35179, new_n35180,
    new_n35181, new_n35182, new_n35183, new_n35184, new_n35185, new_n35186,
    new_n35187, new_n35188, new_n35189, new_n35190, new_n35191, new_n35192,
    new_n35193, new_n35194, new_n35195, new_n35196, new_n35197, new_n35198,
    new_n35199, new_n35200, new_n35201, new_n35202, new_n35203, new_n35204,
    new_n35205, new_n35206, new_n35207, new_n35208, new_n35209, new_n35210,
    new_n35211, new_n35212, new_n35213, new_n35214, new_n35215, new_n35216,
    new_n35217, new_n35218, new_n35219, new_n35220, new_n35221, new_n35222,
    new_n35223, new_n35224, new_n35225, new_n35226, new_n35227, new_n35228,
    new_n35229, new_n35230, new_n35231, new_n35232, new_n35233, new_n35234,
    new_n35235, new_n35236, new_n35237, new_n35238, new_n35239, new_n35240,
    new_n35241, new_n35242, new_n35243, new_n35244, new_n35245, new_n35246,
    new_n35247, new_n35248, new_n35249, new_n35250, new_n35251, new_n35252,
    new_n35253, new_n35254, new_n35255, new_n35256, new_n35257, new_n35258,
    new_n35259, new_n35260, new_n35261, new_n35262, new_n35263, new_n35264,
    new_n35265, new_n35266, new_n35267, new_n35268, new_n35269, new_n35270,
    new_n35271, new_n35272, new_n35273, new_n35274, new_n35275, new_n35276,
    new_n35277, new_n35278, new_n35279, new_n35280, new_n35281, new_n35282,
    new_n35283, new_n35284, new_n35285, new_n35286, new_n35287, new_n35288,
    new_n35289, new_n35290, new_n35291, new_n35292, new_n35293, new_n35294,
    new_n35295, new_n35296, new_n35297, new_n35298, new_n35299, new_n35300,
    new_n35301, new_n35302, new_n35303, new_n35304, new_n35305, new_n35306,
    new_n35307, new_n35308, new_n35309, new_n35310, new_n35311, new_n35312,
    new_n35313, new_n35314, new_n35315, new_n35316, new_n35317, new_n35318,
    new_n35319, new_n35320, new_n35321, new_n35322, new_n35323, new_n35324,
    new_n35325, new_n35326, new_n35327, new_n35328, new_n35329, new_n35330,
    new_n35331, new_n35332, new_n35333, new_n35334, new_n35335, new_n35336,
    new_n35337, new_n35338, new_n35339, new_n35340, new_n35341, new_n35342,
    new_n35343, new_n35344, new_n35345, new_n35346, new_n35347, new_n35348,
    new_n35349, new_n35350, new_n35351, new_n35352, new_n35353, new_n35354,
    new_n35355, new_n35356, new_n35357, new_n35358, new_n35359, new_n35360,
    new_n35361, new_n35362, new_n35363, new_n35364, new_n35365, new_n35366,
    new_n35367, new_n35368, new_n35369, new_n35370, new_n35371, new_n35372,
    new_n35373, new_n35374, new_n35375, new_n35376, new_n35377, new_n35378,
    new_n35379, new_n35380, new_n35381, new_n35382, new_n35383, new_n35384,
    new_n35385, new_n35386, new_n35387, new_n35388, new_n35389, new_n35390,
    new_n35391, new_n35392, new_n35393, new_n35394, new_n35395, new_n35396,
    new_n35397, new_n35398, new_n35399, new_n35400, new_n35401, new_n35402,
    new_n35403, new_n35404, new_n35405, new_n35406, new_n35407, new_n35408,
    new_n35409, new_n35410, new_n35411, new_n35412, new_n35413, new_n35414,
    new_n35415, new_n35416, new_n35417, new_n35418, new_n35419, new_n35420,
    new_n35421, new_n35422, new_n35423, new_n35424, new_n35425, new_n35426,
    new_n35427, new_n35428, new_n35429, new_n35430, new_n35431, new_n35432,
    new_n35433, new_n35434, new_n35435, new_n35436, new_n35437, new_n35438,
    new_n35439, new_n35440, new_n35441, new_n35442, new_n35443, new_n35444,
    new_n35445, new_n35446, new_n35447, new_n35448, new_n35449, new_n35450,
    new_n35451, new_n35452, new_n35453, new_n35454, new_n35455, new_n35456,
    new_n35457, new_n35458, new_n35459, new_n35460, new_n35461, new_n35462,
    new_n35463, new_n35464, new_n35465, new_n35466, new_n35467, new_n35468,
    new_n35469, new_n35470, new_n35471, new_n35472, new_n35473, new_n35474,
    new_n35475, new_n35476, new_n35477, new_n35478, new_n35479, new_n35480,
    new_n35481, new_n35482, new_n35483, new_n35484, new_n35485, new_n35486,
    new_n35487, new_n35488, new_n35489, new_n35490, new_n35491, new_n35492,
    new_n35493, new_n35494, new_n35495, new_n35496, new_n35497, new_n35498,
    new_n35499, new_n35500, new_n35501, new_n35502, new_n35503, new_n35504,
    new_n35505, new_n35506, new_n35507, new_n35508, new_n35509, new_n35510,
    new_n35511, new_n35512, new_n35513, new_n35514, new_n35515, new_n35516,
    new_n35517, new_n35518, new_n35519, new_n35520, new_n35521, new_n35522,
    new_n35523, new_n35524, new_n35525, new_n35526, new_n35527, new_n35528,
    new_n35529, new_n35530, new_n35531, new_n35532, new_n35533, new_n35534,
    new_n35535, new_n35536, new_n35537, new_n35538, new_n35539, new_n35540,
    new_n35541, new_n35542, new_n35543, new_n35544, new_n35545, new_n35546,
    new_n35547, new_n35548, new_n35549, new_n35550, new_n35551, new_n35552,
    new_n35553, new_n35554, new_n35555, new_n35556, new_n35557, new_n35558,
    new_n35559, new_n35560, new_n35561, new_n35562, new_n35563, new_n35564,
    new_n35565, new_n35566, new_n35567, new_n35568, new_n35569, new_n35570,
    new_n35571, new_n35572, new_n35573, new_n35574, new_n35575, new_n35576,
    new_n35577, new_n35578, new_n35579, new_n35580, new_n35581, new_n35582,
    new_n35583, new_n35584, new_n35585, new_n35586, new_n35587, new_n35588,
    new_n35589, new_n35590, new_n35591, new_n35592, new_n35593, new_n35594,
    new_n35595, new_n35596, new_n35597, new_n35598, new_n35599, new_n35600,
    new_n35601, new_n35602, new_n35603, new_n35604, new_n35605, new_n35606,
    new_n35607, new_n35608, new_n35609, new_n35610, new_n35611, new_n35612,
    new_n35613, new_n35614, new_n35615, new_n35616, new_n35617, new_n35618,
    new_n35619, new_n35620, new_n35621, new_n35622, new_n35623, new_n35624,
    new_n35625, new_n35626, new_n35627, new_n35628, new_n35629, new_n35630,
    new_n35631, new_n35632, new_n35633, new_n35634, new_n35635, new_n35636,
    new_n35637, new_n35638, new_n35639, new_n35640, new_n35641, new_n35642,
    new_n35643, new_n35644, new_n35645, new_n35646, new_n35647, new_n35648,
    new_n35649, new_n35650, new_n35651, new_n35652, new_n35653, new_n35654,
    new_n35655, new_n35656, new_n35657, new_n35658, new_n35659, new_n35660,
    new_n35661, new_n35662, new_n35663, new_n35664, new_n35665, new_n35666,
    new_n35667, new_n35668, new_n35669, new_n35670, new_n35671, new_n35672,
    new_n35673, new_n35674, new_n35675, new_n35676, new_n35677, new_n35678,
    new_n35679, new_n35680, new_n35681, new_n35682, new_n35683, new_n35684,
    new_n35685, new_n35686, new_n35687, new_n35688, new_n35689, new_n35690,
    new_n35691, new_n35692, new_n35693, new_n35694, new_n35695, new_n35696,
    new_n35697, new_n35698, new_n35699, new_n35700, new_n35701, new_n35702,
    new_n35703, new_n35704, new_n35705, new_n35706, new_n35707, new_n35708,
    new_n35709, new_n35710, new_n35711, new_n35712, new_n35713, new_n35714,
    new_n35715, new_n35716, new_n35717, new_n35718, new_n35719, new_n35720,
    new_n35721, new_n35722, new_n35723, new_n35724, new_n35725, new_n35726,
    new_n35727, new_n35728, new_n35729, new_n35730, new_n35731, new_n35732,
    new_n35733, new_n35734, new_n35735, new_n35736, new_n35737, new_n35738,
    new_n35739, new_n35740, new_n35741, new_n35742, new_n35743, new_n35744,
    new_n35745, new_n35746, new_n35747, new_n35748, new_n35749, new_n35750,
    new_n35751, new_n35752, new_n35753, new_n35754, new_n35755, new_n35756,
    new_n35757, new_n35758, new_n35759, new_n35760, new_n35761, new_n35762,
    new_n35763, new_n35764, new_n35765, new_n35766, new_n35767, new_n35768,
    new_n35769, new_n35770, new_n35771, new_n35772, new_n35773, new_n35774,
    new_n35775, new_n35776, new_n35777, new_n35778, new_n35779, new_n35780,
    new_n35781, new_n35782, new_n35783, new_n35784, new_n35785, new_n35786,
    new_n35787, new_n35788, new_n35789, new_n35790, new_n35791, new_n35792,
    new_n35793, new_n35794, new_n35795, new_n35796, new_n35797, new_n35798,
    new_n35799, new_n35800, new_n35801, new_n35802, new_n35803, new_n35804,
    new_n35805, new_n35806, new_n35807, new_n35808, new_n35809, new_n35810,
    new_n35811, new_n35812, new_n35813, new_n35814, new_n35815, new_n35816,
    new_n35817, new_n35818, new_n35819, new_n35820, new_n35821, new_n35822,
    new_n35823, new_n35824, new_n35825, new_n35826, new_n35827, new_n35828,
    new_n35829, new_n35830, new_n35831, new_n35832, new_n35833, new_n35834,
    new_n35835, new_n35836, new_n35837, new_n35838, new_n35839, new_n35840,
    new_n35841, new_n35842, new_n35843, new_n35844, new_n35845, new_n35846,
    new_n35847, new_n35848, new_n35849, new_n35850, new_n35851, new_n35852,
    new_n35853, new_n35854, new_n35855, new_n35856, new_n35857, new_n35858,
    new_n35859, new_n35860, new_n35861, new_n35862, new_n35863, new_n35864,
    new_n35865, new_n35866, new_n35867, new_n35868, new_n35869, new_n35870,
    new_n35871, new_n35872, new_n35873, new_n35874, new_n35875, new_n35876,
    new_n35877, new_n35878, new_n35879, new_n35880, new_n35881, new_n35882,
    new_n35883, new_n35884, new_n35885, new_n35886, new_n35887, new_n35888,
    new_n35889, new_n35890, new_n35891, new_n35892, new_n35893, new_n35894,
    new_n35895, new_n35896, new_n35897, new_n35898, new_n35899, new_n35900,
    new_n35901, new_n35902, new_n35903, new_n35904, new_n35905, new_n35906,
    new_n35907, new_n35908, new_n35909, new_n35910, new_n35911, new_n35912,
    new_n35913, new_n35914, new_n35915, new_n35916, new_n35917, new_n35918,
    new_n35919, new_n35920, new_n35921, new_n35922, new_n35923, new_n35924,
    new_n35925, new_n35926, new_n35927, new_n35928, new_n35929, new_n35930,
    new_n35931, new_n35932, new_n35933, new_n35934, new_n35935, new_n35936,
    new_n35937, new_n35938, new_n35939, new_n35940, new_n35941, new_n35942,
    new_n35943, new_n35944, new_n35945, new_n35946, new_n35947, new_n35948,
    new_n35949, new_n35950, new_n35951, new_n35952, new_n35953, new_n35954,
    new_n35955, new_n35956, new_n35957, new_n35958, new_n35959, new_n35960,
    new_n35961, new_n35962, new_n35963, new_n35964, new_n35965, new_n35966,
    new_n35967, new_n35968, new_n35969, new_n35970, new_n35971, new_n35972,
    new_n35973, new_n35974, new_n35975, new_n35976, new_n35977, new_n35978,
    new_n35979, new_n35980, new_n35981, new_n35982, new_n35983, new_n35984,
    new_n35985, new_n35986, new_n35987, new_n35988, new_n35989, new_n35990,
    new_n35991, new_n35992, new_n35993, new_n35994, new_n35995, new_n35996,
    new_n35997, new_n35998, new_n35999, new_n36000, new_n36001, new_n36002,
    new_n36003, new_n36004, new_n36005, new_n36006, new_n36007, new_n36008,
    new_n36009, new_n36010, new_n36011, new_n36012, new_n36013, new_n36014,
    new_n36015, new_n36016, new_n36017, new_n36018, new_n36019, new_n36020,
    new_n36021, new_n36022, new_n36023, new_n36024, new_n36025, new_n36026,
    new_n36027, new_n36028, new_n36029, new_n36030, new_n36031, new_n36032,
    new_n36033, new_n36034, new_n36035, new_n36036, new_n36037, new_n36038,
    new_n36039, new_n36040, new_n36041, new_n36042, new_n36043, new_n36044,
    new_n36045, new_n36046, new_n36047, new_n36048, new_n36049, new_n36050,
    new_n36051, new_n36052, new_n36053, new_n36054, new_n36055, new_n36056,
    new_n36057, new_n36058, new_n36059, new_n36060, new_n36061, new_n36062,
    new_n36063, new_n36064, new_n36065, new_n36066, new_n36067, new_n36068,
    new_n36069, new_n36070, new_n36071, new_n36072, new_n36073, new_n36074,
    new_n36075, new_n36076, new_n36077, new_n36078, new_n36079, new_n36080,
    new_n36081, new_n36082, new_n36083, new_n36084, new_n36085, new_n36086,
    new_n36087, new_n36088, new_n36089, new_n36090, new_n36091, new_n36092,
    new_n36093, new_n36094, new_n36095, new_n36096, new_n36097, new_n36098,
    new_n36099, new_n36100, new_n36101, new_n36102, new_n36103, new_n36104,
    new_n36105, new_n36106, new_n36107, new_n36108, new_n36109, new_n36110,
    new_n36111, new_n36112, new_n36113, new_n36114, new_n36115, new_n36116,
    new_n36117, new_n36118, new_n36119, new_n36120, new_n36121, new_n36122,
    new_n36123, new_n36124, new_n36125, new_n36126, new_n36127, new_n36128,
    new_n36129, new_n36130, new_n36131, new_n36132, new_n36133, new_n36134,
    new_n36135, new_n36136, new_n36137, new_n36138, new_n36139, new_n36140,
    new_n36141, new_n36142, new_n36143, new_n36144, new_n36145, new_n36146,
    new_n36147, new_n36148, new_n36149, new_n36150, new_n36151, new_n36152,
    new_n36153, new_n36154, new_n36155, new_n36156, new_n36157, new_n36158,
    new_n36159, new_n36160, new_n36161, new_n36162, new_n36163, new_n36164,
    new_n36165, new_n36166, new_n36167, new_n36168, new_n36169, new_n36170,
    new_n36171, new_n36172, new_n36173, new_n36174, new_n36175, new_n36176,
    new_n36177, new_n36178, new_n36179, new_n36180, new_n36181, new_n36182,
    new_n36183, new_n36184, new_n36185, new_n36186, new_n36187, new_n36188,
    new_n36189, new_n36190, new_n36191, new_n36192, new_n36193, new_n36194,
    new_n36195, new_n36196, new_n36197, new_n36198, new_n36199, new_n36200,
    new_n36201, new_n36202, new_n36203, new_n36204, new_n36205, new_n36206,
    new_n36207, new_n36208, new_n36209, new_n36210, new_n36211, new_n36212,
    new_n36213, new_n36214, new_n36215, new_n36216, new_n36217, new_n36218,
    new_n36219, new_n36220, new_n36221, new_n36222, new_n36223, new_n36224,
    new_n36225, new_n36226, new_n36227, new_n36228, new_n36229, new_n36230,
    new_n36231, new_n36232, new_n36233, new_n36234, new_n36235, new_n36236,
    new_n36237, new_n36238, new_n36239, new_n36240, new_n36241, new_n36242,
    new_n36243, new_n36244, new_n36245, new_n36246, new_n36247, new_n36248,
    new_n36249, new_n36250, new_n36251, new_n36252, new_n36253, new_n36254,
    new_n36255, new_n36256, new_n36257, new_n36258, new_n36259, new_n36260,
    new_n36261, new_n36262, new_n36263, new_n36264, new_n36265, new_n36266,
    new_n36267, new_n36268, new_n36269, new_n36270, new_n36271, new_n36272,
    new_n36273, new_n36274, new_n36275, new_n36276, new_n36277, new_n36278,
    new_n36279, new_n36280, new_n36281, new_n36282, new_n36283, new_n36284,
    new_n36285, new_n36286, new_n36287, new_n36288, new_n36289, new_n36290,
    new_n36291, new_n36292, new_n36293, new_n36294, new_n36295, new_n36296,
    new_n36297, new_n36298, new_n36299, new_n36300, new_n36301, new_n36302,
    new_n36303, new_n36304, new_n36305, new_n36306, new_n36307, new_n36308,
    new_n36309, new_n36310, new_n36311, new_n36312, new_n36313, new_n36314,
    new_n36315, new_n36316, new_n36317, new_n36318, new_n36319, new_n36320,
    new_n36321, new_n36322, new_n36323, new_n36324, new_n36325;
  assign new_n257 = n28 ^ n27;
  assign new_n258 = n30 ^ n25;
  assign new_n259 = new_n258 ^ new_n257;
  assign new_n260 = n31 ^ n27;
  assign new_n261 = n27 ^ n26;
  assign new_n262 = new_n261 ^ n32;
  assign new_n263 = new_n262 ^ n31;
  assign new_n264 = new_n263 ^ new_n258;
  assign new_n265 = n28 ^ n25;
  assign new_n266 = n31 ^ n29;
  assign new_n267 = new_n266 ^ new_n265;
  assign new_n268 = new_n267 ^ n32;
  assign new_n269 = new_n264 & new_n268;
  assign new_n270 = ~n31 & ~new_n262;
  assign new_n271 = new_n270 ^ n31;
  assign new_n272 = new_n271 ^ new_n269;
  assign new_n273 = n27 ^ n25;
  assign new_n274 = ~new_n261 & n32;
  assign new_n275 = ~n32 & n28;
  assign new_n276 = new_n275 ^ new_n274;
  assign new_n277 = new_n276 ^ n28;
  assign new_n278 = new_n277 ^ new_n269;
  assign new_n279 = n30 ^ n28;
  assign new_n280 = new_n259 & new_n279;
  assign new_n281 = new_n267 ^ new_n261;
  assign new_n282 = new_n258 & new_n281;
  assign new_n283 = new_n282 ^ new_n280;
  assign new_n284 = new_n283 ^ new_n278;
  assign new_n285 = new_n284 ^ new_n273;
  assign new_n286 = n30 ^ n29;
  assign new_n287 = new_n286 ^ n31;
  assign new_n288 = new_n287 ^ n27;
  assign new_n289 = n31 ^ n25;
  assign new_n290 = new_n288 & new_n289;
  assign new_n291 = new_n290 ^ new_n271;
  assign new_n292 = new_n291 ^ new_n258;
  assign new_n293 = new_n287 ^ n26;
  assign new_n294 = new_n265 & new_n293;
  assign new_n295 = new_n294 ^ new_n280;
  assign new_n296 = n29 ^ n27;
  assign new_n297 = new_n296 ^ new_n295;
  assign new_n298 = new_n297 ^ new_n292;
  assign new_n299 = n31 ^ n28;
  assign new_n300 = new_n299 ^ new_n258;
  assign new_n301 = new_n267 & new_n300;
  assign new_n302 = new_n301 ^ n26;
  assign new_n303 = new_n302 ^ new_n267;
  assign new_n304 = new_n294 ^ new_n269;
  assign new_n305 = new_n280 ^ n30;
  assign new_n306 = new_n305 ^ new_n304;
  assign new_n307 = new_n306 ^ new_n303;
  assign new_n308 = ~new_n298 & new_n307;
  assign new_n309 = new_n294 ^ new_n282;
  assign new_n310 = new_n309 ^ new_n288;
  assign new_n311 = new_n293 ^ n32;
  assign new_n312 = new_n262 ^ n25;
  assign new_n313 = new_n311 & new_n312;
  assign new_n314 = new_n313 ^ new_n290;
  assign new_n315 = new_n314 ^ n25;
  assign new_n316 = new_n315 ^ new_n310;
  assign new_n317 = new_n316 ^ new_n308;
  assign new_n318 = new_n285 & new_n317;
  assign new_n319 = new_n302 ^ new_n276;
  assign new_n320 = new_n319 ^ new_n318;
  assign new_n321 = new_n320 ^ new_n310;
  assign new_n322 = new_n319 ^ new_n308;
  assign new_n323 = new_n322 ^ new_n310;
  assign new_n324 = new_n313 ^ new_n270;
  assign new_n325 = new_n324 ^ new_n283;
  assign new_n326 = ~new_n325 & new_n323;
  assign new_n327 = new_n326 ^ new_n308;
  assign new_n328 = new_n316 & new_n327;
  assign new_n329 = new_n328 ^ new_n317;
  assign new_n330 = new_n321 & new_n329;
  assign new_n331 = new_n330 ^ new_n328;
  assign new_n332 = new_n331 ^ new_n272;
  assign new_n333 = new_n332 ^ new_n260;
  assign new_n334 = new_n333 ^ n28;
  assign new_n335 = new_n318 ^ new_n290;
  assign new_n336 = new_n335 ^ new_n302;
  assign new_n337 = new_n336 ^ new_n334;
  assign new_n338 = ~new_n337 & new_n259;
  assign new_n339 = new_n330 ^ new_n285;
  assign new_n340 = new_n262 & new_n339;
  assign new_n341 = new_n328 ^ new_n326;
  assign new_n342 = new_n341 ^ new_n325;
  assign new_n343 = ~new_n342 & new_n264;
  assign new_n344 = ~new_n337 & new_n279;
  assign new_n345 = new_n326 ^ new_n318;
  assign new_n346 = new_n319 ^ new_n315;
  assign new_n347 = new_n346 ^ new_n345;
  assign new_n348 = new_n265 & new_n347;
  assign new_n349 = new_n348 ^ new_n344;
  assign new_n350 = new_n349 ^ new_n343;
  assign new_n351 = new_n350 ^ new_n340;
  assign new_n352 = new_n330 ^ new_n318;
  assign new_n353 = new_n352 ^ new_n307;
  assign new_n354 = new_n288 & new_n353;
  assign new_n355 = new_n354 ^ new_n351;
  assign new_n356 = new_n355 ^ new_n338;
  assign new_n357 = new_n293 & new_n347;
  assign new_n358 = new_n328 ^ new_n298;
  assign new_n359 = ~new_n358 & new_n300;
  assign new_n360 = new_n359 ^ new_n357;
  assign new_n361 = new_n360 ^ new_n356;
  assign new_n362 = new_n361 ^ n65;
  assign new_n363 = new_n362 ^ n97;
  assign new_n364 = new_n363 ^ n33;
  assign new_n365 = new_n364 ^ n1;
  assign new_n366 = ~new_n342 & new_n268;
  assign new_n367 = ~new_n358 & new_n267;
  assign new_n368 = new_n367 ^ new_n366;
  assign new_n369 = new_n368 ^ new_n359;
  assign new_n370 = new_n369 ^ new_n355;
  assign new_n371 = new_n370 ^ n68;
  assign new_n372 = new_n371 ^ n100;
  assign new_n373 = new_n372 ^ n36;
  assign new_n374 = new_n373 ^ n4;
  assign new_n375 = new_n374 ^ new_n365;
  assign new_n376 = new_n326 ^ n25;
  assign new_n377 = new_n313 ^ new_n277;
  assign new_n378 = new_n377 ^ new_n333;
  assign new_n379 = new_n378 ^ new_n376;
  assign new_n380 = ~new_n379 & new_n281;
  assign new_n381 = new_n289 & new_n353;
  assign new_n382 = new_n381 ^ new_n380;
  assign new_n383 = new_n311 & new_n321;
  assign new_n384 = new_n263 & new_n339;
  assign new_n385 = new_n384 ^ new_n383;
  assign new_n386 = new_n385 ^ new_n349;
  assign new_n387 = new_n340 ^ new_n338;
  assign new_n388 = new_n387 ^ new_n386;
  assign new_n389 = new_n388 ^ new_n382;
  assign new_n390 = new_n389 ^ n103;
  assign new_n391 = new_n390 ^ n71;
  assign new_n392 = new_n391 ^ n39;
  assign new_n393 = new_n392 ^ n7;
  assign new_n394 = new_n383 ^ new_n359;
  assign new_n395 = new_n326 ^ new_n316;
  assign new_n396 = n32 & new_n395;
  assign new_n397 = new_n396 ^ new_n366;
  assign new_n398 = new_n397 ^ new_n351;
  assign new_n399 = new_n398 ^ new_n394;
  assign new_n400 = new_n399 ^ n69;
  assign new_n401 = new_n400 ^ n101;
  assign new_n402 = new_n401 ^ n37;
  assign new_n403 = new_n402 ^ n5;
  assign new_n404 = new_n403 ^ new_n393;
  assign new_n405 = new_n404 ^ new_n375;
  assign new_n406 = new_n396 ^ new_n367;
  assign new_n407 = new_n406 ^ new_n381;
  assign new_n408 = new_n407 ^ new_n354;
  assign new_n409 = new_n408 ^ new_n386;
  assign new_n410 = new_n409 ^ n104;
  assign new_n411 = new_n410 ^ n72;
  assign new_n412 = new_n411 ^ n40;
  assign new_n413 = new_n412 ^ n8;
  assign new_n414 = new_n413 ^ new_n405;
  assign new_n415 = new_n262 ^ n28;
  assign new_n416 = new_n395 & new_n415;
  assign new_n417 = new_n416 ^ new_n356;
  assign new_n418 = new_n312 & new_n321;
  assign new_n419 = new_n418 ^ new_n380;
  assign new_n420 = new_n419 ^ new_n407;
  assign new_n421 = new_n420 ^ new_n417;
  assign new_n422 = new_n421 ^ n70;
  assign new_n423 = new_n422 ^ n102;
  assign new_n424 = new_n423 ^ n38;
  assign new_n425 = new_n424 ^ n6;
  assign new_n426 = new_n425 ^ new_n404;
  assign new_n427 = new_n357 ^ new_n338;
  assign new_n428 = new_n369 ^ new_n350;
  assign new_n429 = new_n428 ^ new_n427;
  assign new_n430 = new_n429 ^ n98;
  assign new_n431 = new_n430 ^ n66;
  assign new_n432 = new_n431 ^ n34;
  assign new_n433 = new_n432 ^ n2;
  assign new_n434 = new_n433 ^ new_n426;
  assign new_n435 = new_n375 & new_n434;
  assign new_n436 = new_n425 ^ new_n365;
  assign new_n437 = new_n357 ^ new_n348;
  assign new_n438 = ~new_n379 & new_n258;
  assign new_n439 = new_n438 ^ new_n420;
  assign new_n440 = new_n439 ^ new_n437;
  assign new_n441 = new_n440 ^ n99;
  assign new_n442 = new_n441 ^ n67;
  assign new_n443 = new_n442 ^ n35;
  assign new_n444 = new_n443 ^ n3;
  assign new_n445 = new_n444 ^ new_n433;
  assign new_n446 = new_n445 ^ new_n405;
  assign new_n447 = ~new_n446 & new_n436;
  assign new_n448 = new_n447 ^ new_n435;
  assign new_n449 = new_n444 ^ new_n426;
  assign new_n450 = new_n449 ^ new_n448;
  assign new_n451 = new_n393 ^ new_n365;
  assign new_n452 = ~new_n451 & new_n449;
  assign new_n453 = new_n434 ^ new_n413;
  assign new_n454 = new_n445 ^ new_n413;
  assign new_n455 = new_n454 ^ new_n365;
  assign new_n456 = ~new_n453 & ~new_n455;
  assign new_n457 = new_n456 ^ new_n452;
  assign new_n458 = new_n457 ^ new_n365;
  assign new_n459 = new_n458 ^ new_n450;
  assign new_n460 = new_n393 & new_n454;
  assign new_n461 = new_n460 ^ new_n393;
  assign new_n462 = new_n461 ^ new_n452;
  assign new_n463 = new_n462 ^ new_n436;
  assign new_n464 = new_n444 ^ new_n374;
  assign new_n465 = new_n464 ^ new_n436;
  assign new_n466 = new_n425 ^ new_n374;
  assign new_n467 = ~new_n465 & new_n466;
  assign new_n468 = new_n467 ^ new_n435;
  assign new_n469 = new_n444 ^ new_n403;
  assign new_n470 = new_n469 ^ new_n468;
  assign new_n471 = new_n470 ^ new_n463;
  assign new_n472 = new_n393 ^ new_n374;
  assign new_n473 = new_n472 ^ new_n436;
  assign new_n474 = ~new_n405 & ~new_n473;
  assign new_n475 = new_n474 ^ new_n433;
  assign new_n476 = new_n475 ^ new_n405;
  assign new_n477 = new_n454 ^ new_n393;
  assign new_n478 = new_n477 ^ new_n436;
  assign new_n479 = new_n414 & new_n478;
  assign new_n480 = new_n479 ^ new_n425;
  assign new_n481 = new_n480 ^ new_n468;
  assign new_n482 = new_n481 ^ new_n476;
  assign new_n483 = ~new_n471 & new_n482;
  assign new_n484 = new_n454 ^ new_n374;
  assign new_n485 = ~new_n413 & ~new_n484;
  assign new_n486 = new_n485 ^ new_n374;
  assign new_n487 = new_n486 ^ new_n475;
  assign new_n488 = new_n487 ^ new_n483;
  assign new_n489 = new_n488 ^ new_n450;
  assign new_n490 = new_n460 ^ new_n456;
  assign new_n491 = new_n467 ^ new_n447;
  assign new_n492 = new_n491 ^ new_n490;
  assign new_n493 = ~new_n489 & ~new_n492;
  assign new_n494 = new_n493 ^ new_n483;
  assign new_n495 = ~new_n494 & new_n459;
  assign new_n496 = new_n495 ^ new_n459;
  assign new_n497 = new_n496 ^ new_n493;
  assign new_n498 = new_n497 ^ new_n492;
  assign new_n499 = ~new_n498 & new_n414;
  assign new_n500 = new_n496 ^ new_n471;
  assign new_n501 = ~new_n405 & ~new_n500;
  assign new_n502 = new_n501 ^ new_n499;
  assign new_n503 = ~new_n473 & ~new_n500;
  assign new_n504 = new_n503 ^ new_n502;
  assign new_n505 = ~new_n498 & new_n478;
  assign new_n506 = new_n444 ^ new_n365;
  assign new_n507 = new_n485 ^ new_n479;
  assign new_n508 = new_n507 ^ new_n491;
  assign new_n509 = new_n508 ^ new_n506;
  assign new_n510 = new_n483 ^ new_n459;
  assign new_n511 = ~new_n509 & new_n510;
  assign new_n512 = new_n511 ^ new_n493;
  assign new_n513 = new_n487 ^ new_n458;
  assign new_n514 = new_n513 ^ new_n512;
  assign new_n515 = ~new_n514 & new_n375;
  assign new_n516 = new_n444 ^ new_n393;
  assign new_n517 = new_n479 ^ new_n461;
  assign new_n518 = new_n511 ^ new_n487;
  assign new_n519 = new_n518 ^ new_n450;
  assign new_n520 = new_n495 ^ new_n483;
  assign new_n521 = ~new_n519 & new_n520;
  assign new_n522 = new_n521 ^ new_n496;
  assign new_n523 = new_n522 ^ new_n517;
  assign new_n524 = new_n523 ^ new_n516;
  assign new_n525 = new_n524 ^ new_n374;
  assign new_n526 = new_n511 ^ new_n452;
  assign new_n527 = new_n526 ^ new_n475;
  assign new_n528 = new_n527 ^ new_n525;
  assign new_n529 = ~new_n528 & new_n466;
  assign new_n530 = new_n529 ^ new_n515;
  assign new_n531 = new_n530 ^ new_n505;
  assign new_n532 = new_n521 ^ new_n509;
  assign new_n533 = ~new_n454 & ~new_n532;
  assign new_n534 = new_n533 ^ new_n531;
  assign new_n535 = new_n521 ^ new_n511;
  assign new_n536 = new_n535 ^ new_n482;
  assign new_n537 = new_n449 & new_n536;
  assign new_n538 = new_n537 ^ new_n534;
  assign new_n539 = new_n538 ^ new_n504;
  assign new_n540 = new_n539 ^ n76;
  assign new_n541 = new_n540 ^ n12;
  assign new_n542 = ~new_n514 & new_n434;
  assign new_n543 = new_n542 ^ new_n515;
  assign new_n544 = new_n493 ^ new_n365;
  assign new_n545 = new_n485 ^ new_n456;
  assign new_n546 = new_n545 ^ new_n524;
  assign new_n547 = new_n546 ^ new_n544;
  assign new_n548 = new_n436 & new_n547;
  assign new_n549 = ~new_n455 & ~new_n519;
  assign new_n550 = ~new_n446 & new_n547;
  assign new_n551 = new_n550 ^ new_n549;
  assign new_n552 = new_n493 ^ new_n459;
  assign new_n553 = ~new_n413 & new_n552;
  assign new_n554 = new_n553 ^ new_n501;
  assign new_n555 = ~new_n451 & new_n536;
  assign new_n556 = new_n555 ^ new_n554;
  assign new_n557 = new_n556 ^ new_n551;
  assign new_n558 = new_n557 ^ new_n548;
  assign new_n559 = new_n558 ^ new_n543;
  assign new_n560 = new_n559 ^ n75;
  assign new_n561 = new_n560 ^ n11;
  assign new_n562 = ~new_n465 & ~new_n528;
  assign new_n563 = new_n562 ^ new_n542;
  assign new_n564 = new_n531 ^ new_n504;
  assign new_n565 = new_n564 ^ new_n563;
  assign new_n566 = new_n565 ^ n74;
  assign new_n567 = new_n566 ^ n10;
  assign new_n568 = new_n567 ^ new_n561;
  assign new_n569 = new_n556 ^ new_n537;
  assign new_n570 = ~new_n532 & new_n477;
  assign new_n571 = ~new_n453 & ~new_n519;
  assign new_n572 = new_n571 ^ new_n570;
  assign new_n573 = new_n572 ^ new_n530;
  assign new_n574 = new_n573 ^ new_n569;
  assign new_n575 = new_n574 ^ n80;
  assign new_n576 = new_n575 ^ n16;
  assign new_n577 = new_n576 ^ new_n568;
  assign new_n578 = new_n577 ^ new_n541;
  assign new_n579 = ~new_n576 & ~new_n578;
  assign new_n580 = new_n579 ^ new_n541;
  assign new_n581 = new_n562 ^ new_n538;
  assign new_n582 = new_n542 ^ new_n503;
  assign new_n583 = new_n582 ^ new_n581;
  assign new_n584 = new_n583 ^ n73;
  assign new_n585 = new_n584 ^ n9;
  assign new_n586 = new_n585 ^ new_n541;
  assign new_n587 = new_n555 ^ new_n550;
  assign new_n588 = new_n562 ^ new_n533;
  assign new_n589 = new_n588 ^ new_n573;
  assign new_n590 = new_n589 ^ new_n587;
  assign new_n591 = new_n590 ^ n79;
  assign new_n592 = new_n591 ^ n15;
  assign new_n593 = new_n571 ^ new_n503;
  assign new_n594 = new_n553 ^ new_n499;
  assign new_n595 = new_n594 ^ new_n534;
  assign new_n596 = new_n595 ^ new_n593;
  assign new_n597 = new_n596 ^ n77;
  assign new_n598 = new_n597 ^ n13;
  assign new_n599 = new_n598 ^ new_n592;
  assign new_n600 = new_n599 ^ new_n586;
  assign new_n601 = new_n592 ^ new_n541;
  assign new_n602 = ~new_n484 & new_n552;
  assign new_n603 = new_n602 ^ new_n581;
  assign new_n604 = new_n603 ^ new_n557;
  assign new_n605 = new_n604 ^ n78;
  assign new_n606 = new_n605 ^ n14;
  assign new_n607 = new_n606 ^ new_n585;
  assign new_n608 = new_n607 ^ new_n601;
  assign new_n609 = ~new_n600 & ~new_n608;
  assign new_n610 = new_n609 ^ new_n567;
  assign new_n611 = new_n610 ^ new_n580;
  assign new_n612 = new_n577 & new_n592;
  assign new_n613 = new_n612 ^ new_n592;
  assign new_n614 = new_n606 ^ new_n599;
  assign new_n615 = new_n614 ^ new_n561;
  assign new_n616 = new_n592 ^ new_n585;
  assign new_n617 = ~new_n616 & new_n615;
  assign new_n618 = new_n617 ^ new_n613;
  assign new_n619 = new_n618 ^ new_n607;
  assign new_n620 = new_n561 ^ new_n541;
  assign new_n621 = new_n620 ^ new_n607;
  assign new_n622 = new_n606 ^ new_n541;
  assign new_n623 = ~new_n621 & new_n622;
  assign new_n624 = new_n614 ^ new_n567;
  assign new_n625 = new_n586 & new_n624;
  assign new_n626 = new_n625 ^ new_n623;
  assign new_n627 = new_n598 ^ new_n561;
  assign new_n628 = new_n627 ^ new_n626;
  assign new_n629 = new_n628 ^ new_n619;
  assign new_n630 = new_n610 ^ new_n600;
  assign new_n631 = new_n600 ^ new_n576;
  assign new_n632 = new_n592 ^ new_n577;
  assign new_n633 = new_n632 ^ new_n607;
  assign new_n634 = new_n631 & new_n633;
  assign new_n635 = new_n634 ^ new_n606;
  assign new_n636 = new_n635 ^ new_n626;
  assign new_n637 = new_n636 ^ new_n630;
  assign new_n638 = ~new_n629 & new_n637;
  assign new_n639 = new_n638 ^ new_n611;
  assign new_n640 = new_n600 ^ new_n568;
  assign new_n641 = ~new_n640 & new_n607;
  assign new_n642 = new_n641 ^ new_n625;
  assign new_n643 = new_n642 ^ new_n615;
  assign new_n644 = new_n643 ^ new_n639;
  assign new_n645 = new_n641 ^ new_n623;
  assign new_n646 = new_n585 ^ new_n577;
  assign new_n647 = new_n624 ^ new_n576;
  assign new_n648 = ~new_n646 & ~new_n647;
  assign new_n649 = new_n648 ^ new_n612;
  assign new_n650 = new_n649 ^ new_n645;
  assign new_n651 = ~new_n644 & ~new_n650;
  assign new_n652 = new_n648 ^ new_n617;
  assign new_n653 = new_n652 ^ new_n585;
  assign new_n654 = new_n653 ^ new_n643;
  assign new_n655 = new_n654 ^ new_n651;
  assign new_n656 = ~new_n578 & new_n655;
  assign new_n657 = new_n592 ^ new_n561;
  assign new_n658 = new_n634 ^ new_n613;
  assign new_n659 = new_n651 ^ new_n638;
  assign new_n660 = ~new_n654 & ~new_n659;
  assign new_n661 = new_n660 ^ new_n651;
  assign new_n662 = new_n654 ^ new_n638;
  assign new_n663 = new_n585 ^ new_n561;
  assign new_n664 = new_n634 ^ new_n579;
  assign new_n665 = new_n664 ^ new_n645;
  assign new_n666 = new_n665 ^ new_n663;
  assign new_n667 = ~new_n666 & new_n662;
  assign new_n668 = new_n667 ^ new_n611;
  assign new_n669 = new_n668 ^ new_n643;
  assign new_n670 = ~new_n661 & ~new_n669;
  assign new_n671 = new_n662 ^ new_n661;
  assign new_n672 = new_n671 ^ new_n670;
  assign new_n673 = new_n672 ^ new_n658;
  assign new_n674 = new_n673 ^ new_n657;
  assign new_n675 = new_n674 ^ new_n541;
  assign new_n676 = new_n667 ^ new_n617;
  assign new_n677 = new_n676 ^ new_n610;
  assign new_n678 = new_n677 ^ new_n675;
  assign new_n679 = ~new_n621 & new_n678;
  assign new_n680 = new_n670 ^ new_n666;
  assign new_n681 = ~new_n577 & ~new_n680;
  assign new_n682 = new_n622 & new_n678;
  assign new_n683 = new_n667 ^ new_n651;
  assign new_n684 = new_n653 ^ new_n611;
  assign new_n685 = new_n684 ^ new_n683;
  assign new_n686 = ~new_n685 & new_n586;
  assign new_n687 = new_n686 ^ new_n682;
  assign new_n688 = new_n671 ^ new_n651;
  assign new_n689 = new_n688 ^ new_n650;
  assign new_n690 = new_n633 & new_n689;
  assign new_n691 = new_n690 ^ new_n687;
  assign new_n692 = new_n691 ^ new_n681;
  assign new_n693 = new_n670 ^ new_n667;
  assign new_n694 = new_n693 ^ new_n637;
  assign new_n695 = new_n615 & new_n694;
  assign new_n696 = new_n695 ^ new_n692;
  assign new_n697 = new_n696 ^ new_n679;
  assign new_n698 = new_n697 ^ new_n656;
  assign new_n699 = ~new_n646 & ~new_n669;
  assign new_n700 = new_n651 ^ new_n585;
  assign new_n701 = new_n648 ^ new_n579;
  assign new_n702 = new_n701 ^ new_n674;
  assign new_n703 = new_n702 ^ new_n700;
  assign new_n704 = ~new_n640 & ~new_n703;
  assign new_n705 = new_n704 ^ new_n699;
  assign new_n706 = ~new_n576 & new_n655;
  assign new_n707 = new_n671 ^ new_n629;
  assign new_n708 = ~new_n600 & new_n707;
  assign new_n709 = new_n708 ^ new_n706;
  assign new_n710 = ~new_n616 & new_n694;
  assign new_n711 = new_n710 ^ new_n709;
  assign new_n712 = new_n711 ^ new_n705;
  assign new_n713 = new_n712 ^ new_n698;
  assign new_n714 = new_n713 ^ n54;
  assign new_n715 = n4 ^ n3;
  assign new_n716 = n6 ^ n1;
  assign new_n717 = new_n716 ^ new_n715;
  assign new_n718 = n7 ^ n3;
  assign new_n719 = n3 ^ n2;
  assign new_n720 = new_n719 ^ n8;
  assign new_n721 = new_n720 ^ n7;
  assign new_n722 = new_n721 ^ new_n716;
  assign new_n723 = n7 ^ n5;
  assign new_n724 = n4 ^ n1;
  assign new_n725 = new_n724 ^ new_n723;
  assign new_n726 = new_n725 ^ n8;
  assign new_n727 = new_n722 & new_n726;
  assign new_n728 = ~n7 & ~new_n720;
  assign new_n729 = new_n728 ^ n7;
  assign new_n730 = new_n729 ^ new_n727;
  assign new_n731 = n6 ^ n5;
  assign new_n732 = new_n731 ^ n7;
  assign new_n733 = new_n732 ^ n3;
  assign new_n734 = n7 ^ n1;
  assign new_n735 = new_n733 & new_n734;
  assign new_n736 = new_n735 ^ new_n729;
  assign new_n737 = new_n736 ^ new_n716;
  assign new_n738 = n6 ^ n4;
  assign new_n739 = new_n717 & new_n738;
  assign new_n740 = new_n732 ^ n2;
  assign new_n741 = new_n724 & new_n740;
  assign new_n742 = new_n741 ^ new_n739;
  assign new_n743 = n5 ^ n3;
  assign new_n744 = new_n743 ^ new_n742;
  assign new_n745 = new_n744 ^ new_n737;
  assign new_n746 = n7 ^ n4;
  assign new_n747 = new_n746 ^ new_n716;
  assign new_n748 = new_n725 & new_n747;
  assign new_n749 = new_n748 ^ n2;
  assign new_n750 = new_n749 ^ new_n725;
  assign new_n751 = new_n741 ^ new_n727;
  assign new_n752 = new_n739 ^ n6;
  assign new_n753 = new_n752 ^ new_n751;
  assign new_n754 = new_n753 ^ new_n750;
  assign new_n755 = ~new_n745 & new_n754;
  assign new_n756 = new_n725 ^ new_n719;
  assign new_n757 = new_n716 & new_n756;
  assign new_n758 = new_n757 ^ new_n741;
  assign new_n759 = new_n758 ^ new_n733;
  assign new_n760 = new_n720 ^ n1;
  assign new_n761 = new_n740 ^ n8;
  assign new_n762 = new_n760 & new_n761;
  assign new_n763 = new_n762 ^ new_n735;
  assign new_n764 = new_n763 ^ n1;
  assign new_n765 = new_n764 ^ new_n759;
  assign new_n766 = new_n765 ^ new_n755;
  assign new_n767 = ~new_n719 & n8;
  assign new_n768 = ~n8 & n4;
  assign new_n769 = new_n768 ^ new_n767;
  assign new_n770 = new_n769 ^ new_n749;
  assign new_n771 = new_n770 ^ new_n755;
  assign new_n772 = new_n771 ^ new_n759;
  assign new_n773 = new_n757 ^ new_n739;
  assign new_n774 = new_n762 ^ new_n728;
  assign new_n775 = new_n774 ^ new_n773;
  assign new_n776 = ~new_n775 & new_n772;
  assign new_n777 = new_n776 ^ new_n755;
  assign new_n778 = ~new_n765 & ~new_n777;
  assign new_n779 = new_n778 ^ new_n776;
  assign new_n780 = new_n779 ^ new_n766;
  assign new_n781 = n3 ^ n1;
  assign new_n782 = new_n769 ^ n4;
  assign new_n783 = new_n782 ^ new_n727;
  assign new_n784 = new_n783 ^ new_n773;
  assign new_n785 = new_n784 ^ new_n781;
  assign new_n786 = new_n766 & new_n785;
  assign new_n787 = new_n786 ^ new_n770;
  assign new_n788 = new_n787 ^ new_n759;
  assign new_n789 = ~new_n779 & new_n788;
  assign new_n790 = new_n789 ^ new_n780;
  assign new_n791 = new_n790 ^ new_n730;
  assign new_n792 = new_n791 ^ new_n718;
  assign new_n793 = new_n792 ^ n4;
  assign new_n794 = new_n786 ^ new_n735;
  assign new_n795 = new_n794 ^ new_n749;
  assign new_n796 = new_n795 ^ new_n793;
  assign new_n797 = new_n717 & new_n796;
  assign new_n798 = new_n786 ^ new_n776;
  assign new_n799 = new_n770 ^ new_n764;
  assign new_n800 = new_n799 ^ new_n798;
  assign new_n801 = new_n740 & new_n800;
  assign new_n802 = new_n801 ^ new_n797;
  assign new_n803 = new_n780 ^ new_n776;
  assign new_n804 = new_n803 ^ new_n775;
  assign new_n805 = new_n722 & new_n804;
  assign new_n806 = new_n738 & new_n796;
  assign new_n807 = new_n724 & new_n800;
  assign new_n808 = new_n807 ^ new_n806;
  assign new_n809 = new_n808 ^ new_n805;
  assign new_n810 = new_n780 ^ new_n745;
  assign new_n811 = new_n747 & new_n810;
  assign new_n812 = new_n726 & new_n804;
  assign new_n813 = new_n725 & new_n810;
  assign new_n814 = new_n813 ^ new_n812;
  assign new_n815 = new_n814 ^ new_n811;
  assign new_n816 = new_n815 ^ new_n809;
  assign new_n817 = new_n816 ^ new_n802;
  assign new_n818 = new_n817 ^ n106;
  assign new_n819 = new_n818 ^ n74;
  assign new_n820 = new_n819 ^ n42;
  assign new_n821 = new_n820 ^ n10;
  assign new_n822 = new_n807 ^ new_n801;
  assign new_n823 = new_n776 ^ n1;
  assign new_n824 = new_n782 ^ new_n762;
  assign new_n825 = new_n824 ^ new_n792;
  assign new_n826 = new_n825 ^ new_n823;
  assign new_n827 = new_n756 & new_n826;
  assign new_n828 = new_n760 & new_n788;
  assign new_n829 = new_n828 ^ new_n827;
  assign new_n830 = new_n789 ^ new_n786;
  assign new_n831 = new_n830 ^ new_n754;
  assign new_n832 = new_n734 & new_n831;
  assign new_n833 = new_n776 ^ new_n765;
  assign new_n834 = n8 & new_n833;
  assign new_n835 = new_n834 ^ new_n813;
  assign new_n836 = new_n835 ^ new_n832;
  assign new_n837 = new_n836 ^ new_n829;
  assign new_n838 = new_n716 & new_n826;
  assign new_n839 = new_n838 ^ new_n837;
  assign new_n840 = new_n839 ^ new_n822;
  assign new_n841 = new_n840 ^ n107;
  assign new_n842 = new_n841 ^ n75;
  assign new_n843 = new_n842 ^ n43;
  assign new_n844 = new_n843 ^ n11;
  assign new_n845 = new_n844 ^ new_n821;
  assign new_n846 = new_n761 & new_n788;
  assign new_n847 = new_n789 ^ new_n785;
  assign new_n848 = new_n721 & new_n847;
  assign new_n849 = new_n848 ^ new_n846;
  assign new_n850 = new_n849 ^ new_n808;
  assign new_n851 = new_n733 & new_n831;
  assign new_n852 = new_n851 ^ new_n836;
  assign new_n853 = new_n852 ^ new_n850;
  assign new_n854 = new_n853 ^ n112;
  assign new_n855 = new_n854 ^ n80;
  assign new_n856 = new_n855 ^ n48;
  assign new_n857 = new_n856 ^ n16;
  assign new_n858 = new_n857 ^ new_n845;
  assign new_n859 = new_n720 & new_n847;
  assign new_n860 = new_n859 ^ new_n809;
  assign new_n861 = new_n860 ^ new_n851;
  assign new_n862 = new_n861 ^ new_n815;
  assign new_n863 = new_n862 ^ n76;
  assign new_n864 = new_n863 ^ n108;
  assign new_n865 = new_n864 ^ n44;
  assign new_n866 = new_n865 ^ n12;
  assign new_n867 = new_n866 ^ new_n858;
  assign new_n868 = ~new_n857 & ~new_n867;
  assign new_n869 = new_n868 ^ new_n866;
  assign new_n870 = new_n811 ^ new_n801;
  assign new_n871 = new_n861 ^ new_n797;
  assign new_n872 = new_n871 ^ new_n870;
  assign new_n873 = new_n872 ^ n73;
  assign new_n874 = new_n873 ^ n105;
  assign new_n875 = new_n874 ^ n41;
  assign new_n876 = new_n875 ^ n9;
  assign new_n877 = new_n876 ^ new_n866;
  assign new_n878 = new_n846 ^ new_n811;
  assign new_n879 = new_n834 ^ new_n812;
  assign new_n880 = new_n879 ^ new_n860;
  assign new_n881 = new_n880 ^ new_n878;
  assign new_n882 = new_n881 ^ n77;
  assign new_n883 = new_n882 ^ n109;
  assign new_n884 = new_n883 ^ n45;
  assign new_n885 = new_n884 ^ n13;
  assign new_n886 = new_n832 ^ new_n827;
  assign new_n887 = new_n859 ^ new_n797;
  assign new_n888 = new_n887 ^ new_n850;
  assign new_n889 = new_n888 ^ new_n886;
  assign new_n890 = new_n889 ^ n111;
  assign new_n891 = new_n890 ^ n79;
  assign new_n892 = new_n891 ^ n47;
  assign new_n893 = new_n892 ^ n15;
  assign new_n894 = new_n893 ^ new_n885;
  assign new_n895 = new_n894 ^ new_n877;
  assign new_n896 = new_n893 ^ new_n866;
  assign new_n897 = new_n720 ^ n4;
  assign new_n898 = new_n833 & new_n897;
  assign new_n899 = new_n898 ^ new_n871;
  assign new_n900 = new_n899 ^ new_n837;
  assign new_n901 = new_n900 ^ n78;
  assign new_n902 = new_n901 ^ n110;
  assign new_n903 = new_n902 ^ n46;
  assign new_n904 = new_n903 ^ n14;
  assign new_n905 = new_n904 ^ new_n876;
  assign new_n906 = new_n905 ^ new_n896;
  assign new_n907 = ~new_n895 & ~new_n906;
  assign new_n908 = new_n907 ^ new_n821;
  assign new_n909 = new_n908 ^ new_n869;
  assign new_n910 = new_n858 & new_n893;
  assign new_n911 = new_n910 ^ new_n893;
  assign new_n912 = new_n893 ^ new_n876;
  assign new_n913 = new_n904 ^ new_n894;
  assign new_n914 = new_n913 ^ new_n844;
  assign new_n915 = ~new_n912 & new_n914;
  assign new_n916 = new_n915 ^ new_n911;
  assign new_n917 = new_n916 ^ new_n905;
  assign new_n918 = new_n866 ^ new_n844;
  assign new_n919 = new_n918 ^ new_n905;
  assign new_n920 = new_n904 ^ new_n866;
  assign new_n921 = ~new_n919 & new_n920;
  assign new_n922 = new_n913 ^ new_n821;
  assign new_n923 = new_n877 & new_n922;
  assign new_n924 = new_n923 ^ new_n921;
  assign new_n925 = new_n885 ^ new_n844;
  assign new_n926 = new_n925 ^ new_n924;
  assign new_n927 = new_n926 ^ new_n917;
  assign new_n928 = new_n908 ^ new_n895;
  assign new_n929 = new_n895 ^ new_n857;
  assign new_n930 = new_n893 ^ new_n858;
  assign new_n931 = new_n930 ^ new_n905;
  assign new_n932 = new_n929 & new_n931;
  assign new_n933 = new_n932 ^ new_n904;
  assign new_n934 = new_n933 ^ new_n924;
  assign new_n935 = new_n934 ^ new_n928;
  assign new_n936 = ~new_n927 & new_n935;
  assign new_n937 = new_n936 ^ new_n909;
  assign new_n938 = new_n895 ^ new_n845;
  assign new_n939 = ~new_n938 & new_n905;
  assign new_n940 = new_n939 ^ new_n923;
  assign new_n941 = new_n940 ^ new_n914;
  assign new_n942 = new_n941 ^ new_n937;
  assign new_n943 = new_n876 ^ new_n858;
  assign new_n944 = new_n922 ^ new_n857;
  assign new_n945 = ~new_n943 & ~new_n944;
  assign new_n946 = new_n945 ^ new_n910;
  assign new_n947 = new_n939 ^ new_n921;
  assign new_n948 = new_n947 ^ new_n946;
  assign new_n949 = ~new_n942 & ~new_n948;
  assign new_n950 = new_n945 ^ new_n915;
  assign new_n951 = new_n950 ^ new_n876;
  assign new_n952 = new_n951 ^ new_n941;
  assign new_n953 = new_n952 ^ new_n949;
  assign new_n954 = ~new_n867 & new_n953;
  assign new_n955 = new_n952 ^ new_n936;
  assign new_n956 = new_n949 ^ new_n936;
  assign new_n957 = ~new_n952 & ~new_n956;
  assign new_n958 = new_n957 ^ new_n949;
  assign new_n959 = new_n958 ^ new_n955;
  assign new_n960 = new_n959 ^ new_n949;
  assign new_n961 = new_n960 ^ new_n948;
  assign new_n962 = new_n931 & new_n961;
  assign new_n963 = new_n876 ^ new_n844;
  assign new_n964 = new_n932 ^ new_n868;
  assign new_n965 = new_n964 ^ new_n947;
  assign new_n966 = new_n965 ^ new_n963;
  assign new_n967 = ~new_n966 & new_n955;
  assign new_n968 = new_n967 ^ new_n949;
  assign new_n969 = new_n951 ^ new_n909;
  assign new_n970 = new_n969 ^ new_n968;
  assign new_n971 = ~new_n970 & new_n877;
  assign new_n972 = new_n893 ^ new_n844;
  assign new_n973 = new_n932 ^ new_n911;
  assign new_n974 = new_n967 ^ new_n909;
  assign new_n975 = new_n974 ^ new_n941;
  assign new_n976 = ~new_n958 & ~new_n975;
  assign new_n977 = new_n976 ^ new_n959;
  assign new_n978 = new_n977 ^ new_n973;
  assign new_n979 = new_n978 ^ new_n972;
  assign new_n980 = new_n979 ^ new_n866;
  assign new_n981 = new_n967 ^ new_n915;
  assign new_n982 = new_n981 ^ new_n908;
  assign new_n983 = new_n982 ^ new_n980;
  assign new_n984 = new_n920 & new_n983;
  assign new_n985 = new_n984 ^ new_n971;
  assign new_n986 = new_n985 ^ new_n962;
  assign new_n987 = new_n976 ^ new_n966;
  assign new_n988 = ~new_n858 & ~new_n987;
  assign new_n989 = new_n988 ^ new_n986;
  assign new_n990 = new_n976 ^ new_n967;
  assign new_n991 = new_n990 ^ new_n935;
  assign new_n992 = new_n914 & new_n991;
  assign new_n993 = new_n992 ^ new_n989;
  assign new_n994 = ~new_n919 & new_n983;
  assign new_n995 = new_n994 ^ new_n993;
  assign new_n996 = new_n995 ^ new_n954;
  assign new_n997 = ~new_n943 & ~new_n975;
  assign new_n998 = new_n949 ^ new_n876;
  assign new_n999 = new_n945 ^ new_n868;
  assign new_n1000 = new_n999 ^ new_n979;
  assign new_n1001 = new_n1000 ^ new_n998;
  assign new_n1002 = ~new_n938 & ~new_n1001;
  assign new_n1003 = new_n1002 ^ new_n997;
  assign new_n1004 = ~new_n857 & new_n953;
  assign new_n1005 = new_n959 ^ new_n927;
  assign new_n1006 = ~new_n895 & new_n1005;
  assign new_n1007 = new_n1006 ^ new_n1004;
  assign new_n1008 = ~new_n912 & new_n991;
  assign new_n1009 = new_n1008 ^ new_n1007;
  assign new_n1010 = new_n1009 ^ new_n1003;
  assign new_n1011 = new_n1010 ^ new_n996;
  assign new_n1012 = new_n1011 ^ n86;
  assign new_n1013 = new_n1012 ^ new_n714;
  assign new_n1014 = n14 ^ n13;
  assign new_n1015 = new_n1014 ^ n15;
  assign new_n1016 = new_n1015 ^ n10;
  assign new_n1017 = n11 ^ n9;
  assign new_n1018 = n11 ^ n10;
  assign new_n1019 = ~new_n1018 & n16;
  assign new_n1020 = ~n16 & n12;
  assign new_n1021 = new_n1020 ^ new_n1019;
  assign new_n1022 = new_n1021 ^ n12;
  assign new_n1023 = n12 ^ n9;
  assign new_n1024 = n15 ^ n13;
  assign new_n1025 = new_n1024 ^ new_n1023;
  assign new_n1026 = new_n1025 ^ n16;
  assign new_n1027 = new_n1018 ^ n16;
  assign new_n1028 = new_n1027 ^ n15;
  assign new_n1029 = n14 ^ n9;
  assign new_n1030 = new_n1029 ^ new_n1028;
  assign new_n1031 = new_n1026 & new_n1030;
  assign new_n1032 = new_n1031 ^ new_n1022;
  assign new_n1033 = n12 ^ n11;
  assign new_n1034 = new_n1033 ^ new_n1029;
  assign new_n1035 = n14 ^ n12;
  assign new_n1036 = new_n1034 & new_n1035;
  assign new_n1037 = new_n1025 ^ new_n1018;
  assign new_n1038 = new_n1029 & new_n1037;
  assign new_n1039 = new_n1038 ^ new_n1036;
  assign new_n1040 = new_n1039 ^ new_n1032;
  assign new_n1041 = new_n1040 ^ new_n1017;
  assign new_n1042 = ~n15 & ~new_n1027;
  assign new_n1043 = new_n1042 ^ n15;
  assign new_n1044 = new_n1015 ^ n11;
  assign new_n1045 = n15 ^ n9;
  assign new_n1046 = new_n1044 & new_n1045;
  assign new_n1047 = new_n1046 ^ new_n1043;
  assign new_n1048 = new_n1047 ^ new_n1029;
  assign new_n1049 = new_n1016 & new_n1023;
  assign new_n1050 = new_n1049 ^ new_n1036;
  assign new_n1051 = n13 ^ n11;
  assign new_n1052 = new_n1051 ^ new_n1050;
  assign new_n1053 = new_n1052 ^ new_n1048;
  assign new_n1054 = n15 ^ n12;
  assign new_n1055 = new_n1054 ^ new_n1029;
  assign new_n1056 = new_n1025 & new_n1055;
  assign new_n1057 = new_n1056 ^ n10;
  assign new_n1058 = new_n1057 ^ new_n1025;
  assign new_n1059 = new_n1049 ^ new_n1031;
  assign new_n1060 = new_n1036 ^ n14;
  assign new_n1061 = new_n1060 ^ new_n1059;
  assign new_n1062 = new_n1061 ^ new_n1058;
  assign new_n1063 = ~new_n1053 & new_n1062;
  assign new_n1064 = new_n1049 ^ new_n1038;
  assign new_n1065 = new_n1064 ^ new_n1044;
  assign new_n1066 = new_n1016 ^ n16;
  assign new_n1067 = new_n1027 ^ n9;
  assign new_n1068 = new_n1066 & new_n1067;
  assign new_n1069 = new_n1068 ^ new_n1046;
  assign new_n1070 = new_n1069 ^ n9;
  assign new_n1071 = new_n1070 ^ new_n1065;
  assign new_n1072 = new_n1071 ^ new_n1063;
  assign new_n1073 = new_n1041 & new_n1072;
  assign new_n1074 = new_n1057 ^ new_n1021;
  assign new_n1075 = new_n1074 ^ new_n1063;
  assign new_n1076 = new_n1075 ^ new_n1065;
  assign new_n1077 = new_n1068 ^ new_n1042;
  assign new_n1078 = new_n1077 ^ new_n1039;
  assign new_n1079 = ~new_n1078 & new_n1076;
  assign new_n1080 = new_n1079 ^ new_n1073;
  assign new_n1081 = new_n1074 ^ new_n1070;
  assign new_n1082 = new_n1081 ^ new_n1080;
  assign new_n1083 = new_n1016 & new_n1082;
  assign new_n1084 = n15 ^ n11;
  assign new_n1085 = new_n1043 ^ new_n1031;
  assign new_n1086 = new_n1074 ^ new_n1073;
  assign new_n1087 = new_n1086 ^ new_n1065;
  assign new_n1088 = new_n1079 ^ new_n1063;
  assign new_n1089 = new_n1071 & new_n1088;
  assign new_n1090 = new_n1089 ^ new_n1072;
  assign new_n1091 = new_n1087 & new_n1090;
  assign new_n1092 = new_n1091 ^ new_n1089;
  assign new_n1093 = new_n1092 ^ new_n1085;
  assign new_n1094 = new_n1093 ^ new_n1084;
  assign new_n1095 = new_n1094 ^ n12;
  assign new_n1096 = new_n1073 ^ new_n1046;
  assign new_n1097 = new_n1096 ^ new_n1057;
  assign new_n1098 = new_n1097 ^ new_n1095;
  assign new_n1099 = ~new_n1098 & new_n1034;
  assign new_n1100 = new_n1099 ^ new_n1083;
  assign new_n1101 = new_n1089 ^ new_n1079;
  assign new_n1102 = new_n1101 ^ new_n1078;
  assign new_n1103 = ~new_n1102 & new_n1030;
  assign new_n1104 = ~new_n1098 & new_n1035;
  assign new_n1105 = new_n1023 & new_n1082;
  assign new_n1106 = new_n1105 ^ new_n1104;
  assign new_n1107 = new_n1106 ^ new_n1103;
  assign new_n1108 = new_n1089 ^ new_n1053;
  assign new_n1109 = ~new_n1108 & new_n1055;
  assign new_n1110 = ~new_n1102 & new_n1026;
  assign new_n1111 = ~new_n1108 & new_n1025;
  assign new_n1112 = new_n1111 ^ new_n1110;
  assign new_n1113 = new_n1112 ^ new_n1109;
  assign new_n1114 = new_n1113 ^ new_n1107;
  assign new_n1115 = new_n1114 ^ new_n1100;
  assign new_n1116 = new_n1115 ^ n114;
  assign new_n1117 = new_n1116 ^ n82;
  assign new_n1118 = new_n1117 ^ n50;
  assign new_n1119 = new_n1118 ^ n18;
  assign new_n1120 = new_n1105 ^ new_n1083;
  assign new_n1121 = new_n1079 ^ n9;
  assign new_n1122 = new_n1068 ^ new_n1022;
  assign new_n1123 = new_n1122 ^ new_n1094;
  assign new_n1124 = new_n1123 ^ new_n1121;
  assign new_n1125 = ~new_n1124 & new_n1029;
  assign new_n1126 = ~new_n1124 & new_n1037;
  assign new_n1127 = new_n1067 & new_n1087;
  assign new_n1128 = new_n1127 ^ new_n1126;
  assign new_n1129 = new_n1091 ^ new_n1073;
  assign new_n1130 = new_n1129 ^ new_n1062;
  assign new_n1131 = new_n1045 & new_n1130;
  assign new_n1132 = new_n1079 ^ new_n1071;
  assign new_n1133 = n16 & new_n1132;
  assign new_n1134 = new_n1133 ^ new_n1111;
  assign new_n1135 = new_n1134 ^ new_n1131;
  assign new_n1136 = new_n1135 ^ new_n1128;
  assign new_n1137 = new_n1136 ^ new_n1125;
  assign new_n1138 = new_n1137 ^ new_n1120;
  assign new_n1139 = new_n1138 ^ n83;
  assign new_n1140 = new_n1139 ^ n115;
  assign new_n1141 = new_n1140 ^ n51;
  assign new_n1142 = new_n1141 ^ n19;
  assign new_n1143 = new_n1142 ^ new_n1119;
  assign new_n1144 = new_n1044 & new_n1130;
  assign new_n1145 = new_n1144 ^ new_n1135;
  assign new_n1146 = new_n1066 & new_n1087;
  assign new_n1147 = new_n1091 ^ new_n1041;
  assign new_n1148 = new_n1028 & new_n1147;
  assign new_n1149 = new_n1148 ^ new_n1146;
  assign new_n1150 = new_n1149 ^ new_n1106;
  assign new_n1151 = new_n1150 ^ new_n1145;
  assign new_n1152 = new_n1151 ^ n120;
  assign new_n1153 = new_n1152 ^ n88;
  assign new_n1154 = new_n1153 ^ n56;
  assign new_n1155 = new_n1154 ^ n24;
  assign new_n1156 = new_n1155 ^ new_n1143;
  assign new_n1157 = new_n1027 & new_n1147;
  assign new_n1158 = new_n1157 ^ new_n1107;
  assign new_n1159 = new_n1158 ^ new_n1144;
  assign new_n1160 = new_n1159 ^ new_n1113;
  assign new_n1161 = new_n1160 ^ n84;
  assign new_n1162 = new_n1161 ^ n116;
  assign new_n1163 = new_n1162 ^ n52;
  assign new_n1164 = new_n1163 ^ n20;
  assign new_n1165 = new_n1164 ^ new_n1156;
  assign new_n1166 = ~new_n1155 & ~new_n1165;
  assign new_n1167 = new_n1166 ^ new_n1164;
  assign new_n1168 = new_n1146 ^ new_n1109;
  assign new_n1169 = new_n1133 ^ new_n1110;
  assign new_n1170 = new_n1169 ^ new_n1158;
  assign new_n1171 = new_n1170 ^ new_n1168;
  assign new_n1172 = new_n1171 ^ n85;
  assign new_n1173 = new_n1172 ^ n117;
  assign new_n1174 = new_n1173 ^ n53;
  assign new_n1175 = new_n1174 ^ n21;
  assign new_n1176 = new_n1131 ^ new_n1126;
  assign new_n1177 = new_n1157 ^ new_n1099;
  assign new_n1178 = new_n1177 ^ new_n1150;
  assign new_n1179 = new_n1178 ^ new_n1176;
  assign new_n1180 = new_n1179 ^ n119;
  assign new_n1181 = new_n1180 ^ n87;
  assign new_n1182 = new_n1181 ^ n55;
  assign new_n1183 = new_n1182 ^ n23;
  assign new_n1184 = new_n1183 ^ new_n1175;
  assign new_n1185 = new_n1109 ^ new_n1083;
  assign new_n1186 = new_n1159 ^ new_n1099;
  assign new_n1187 = new_n1186 ^ new_n1185;
  assign new_n1188 = new_n1187 ^ n81;
  assign new_n1189 = new_n1188 ^ n113;
  assign new_n1190 = new_n1189 ^ n49;
  assign new_n1191 = new_n1190 ^ n17;
  assign new_n1192 = new_n1191 ^ new_n1164;
  assign new_n1193 = new_n1192 ^ new_n1184;
  assign new_n1194 = new_n1183 ^ new_n1164;
  assign new_n1195 = new_n1027 ^ n12;
  assign new_n1196 = new_n1132 & new_n1195;
  assign new_n1197 = new_n1196 ^ new_n1186;
  assign new_n1198 = new_n1197 ^ new_n1136;
  assign new_n1199 = new_n1198 ^ n86;
  assign new_n1200 = new_n1199 ^ n118;
  assign new_n1201 = new_n1200 ^ n54;
  assign new_n1202 = new_n1201 ^ n22;
  assign new_n1203 = new_n1202 ^ new_n1191;
  assign new_n1204 = new_n1203 ^ new_n1194;
  assign new_n1205 = ~new_n1193 & ~new_n1204;
  assign new_n1206 = new_n1205 ^ new_n1119;
  assign new_n1207 = new_n1206 ^ new_n1167;
  assign new_n1208 = new_n1191 ^ new_n1142;
  assign new_n1209 = new_n1202 ^ new_n1164;
  assign new_n1210 = new_n1164 ^ new_n1142;
  assign new_n1211 = new_n1210 ^ new_n1203;
  assign new_n1212 = ~new_n1211 & new_n1209;
  assign new_n1213 = new_n1193 ^ new_n1143;
  assign new_n1214 = ~new_n1213 & new_n1203;
  assign new_n1215 = new_n1214 ^ new_n1212;
  assign new_n1216 = new_n1193 ^ new_n1155;
  assign new_n1217 = new_n1183 ^ new_n1156;
  assign new_n1218 = new_n1217 ^ new_n1203;
  assign new_n1219 = new_n1216 & new_n1218;
  assign new_n1220 = new_n1219 ^ new_n1166;
  assign new_n1221 = new_n1220 ^ new_n1215;
  assign new_n1222 = new_n1221 ^ new_n1208;
  assign new_n1223 = new_n1156 & new_n1183;
  assign new_n1224 = new_n1223 ^ new_n1183;
  assign new_n1225 = new_n1202 ^ new_n1184;
  assign new_n1226 = new_n1225 ^ new_n1142;
  assign new_n1227 = new_n1191 ^ new_n1183;
  assign new_n1228 = ~new_n1227 & new_n1226;
  assign new_n1229 = new_n1228 ^ new_n1224;
  assign new_n1230 = new_n1229 ^ new_n1203;
  assign new_n1231 = new_n1225 ^ new_n1119;
  assign new_n1232 = new_n1192 & new_n1231;
  assign new_n1233 = new_n1232 ^ new_n1212;
  assign new_n1234 = new_n1175 ^ new_n1142;
  assign new_n1235 = new_n1234 ^ new_n1233;
  assign new_n1236 = new_n1235 ^ new_n1230;
  assign new_n1237 = new_n1206 ^ new_n1193;
  assign new_n1238 = new_n1219 ^ new_n1202;
  assign new_n1239 = new_n1238 ^ new_n1233;
  assign new_n1240 = new_n1239 ^ new_n1237;
  assign new_n1241 = ~new_n1236 & new_n1240;
  assign new_n1242 = new_n1232 ^ new_n1214;
  assign new_n1243 = new_n1242 ^ new_n1226;
  assign new_n1244 = new_n1191 ^ new_n1156;
  assign new_n1245 = new_n1231 ^ new_n1155;
  assign new_n1246 = ~new_n1244 & ~new_n1245;
  assign new_n1247 = new_n1246 ^ new_n1228;
  assign new_n1248 = new_n1247 ^ new_n1191;
  assign new_n1249 = new_n1248 ^ new_n1243;
  assign new_n1250 = new_n1249 ^ new_n1241;
  assign new_n1251 = ~new_n1222 & new_n1250;
  assign new_n1252 = new_n1251 ^ new_n1207;
  assign new_n1253 = new_n1252 ^ new_n1243;
  assign new_n1254 = new_n1241 ^ new_n1207;
  assign new_n1255 = new_n1254 ^ new_n1243;
  assign new_n1256 = new_n1246 ^ new_n1223;
  assign new_n1257 = new_n1256 ^ new_n1215;
  assign new_n1258 = ~new_n1255 & ~new_n1257;
  assign new_n1259 = new_n1258 ^ new_n1241;
  assign new_n1260 = new_n1249 & new_n1259;
  assign new_n1261 = new_n1260 ^ new_n1250;
  assign new_n1262 = ~new_n1253 & new_n1261;
  assign new_n1263 = new_n1262 ^ new_n1222;
  assign new_n1264 = ~new_n1156 & ~new_n1263;
  assign new_n1265 = new_n1260 ^ new_n1258;
  assign new_n1266 = new_n1265 ^ new_n1257;
  assign new_n1267 = ~new_n1266 & new_n1218;
  assign new_n1268 = new_n1258 ^ new_n1251;
  assign new_n1269 = new_n1248 ^ new_n1207;
  assign new_n1270 = new_n1269 ^ new_n1268;
  assign new_n1271 = ~new_n1270 & new_n1192;
  assign new_n1272 = new_n1183 ^ new_n1142;
  assign new_n1273 = new_n1224 ^ new_n1219;
  assign new_n1274 = new_n1262 ^ new_n1260;
  assign new_n1275 = new_n1274 ^ new_n1273;
  assign new_n1276 = new_n1275 ^ new_n1272;
  assign new_n1277 = new_n1276 ^ new_n1164;
  assign new_n1278 = new_n1251 ^ new_n1228;
  assign new_n1279 = new_n1278 ^ new_n1206;
  assign new_n1280 = new_n1279 ^ new_n1277;
  assign new_n1281 = ~new_n1280 & new_n1209;
  assign new_n1282 = new_n1281 ^ new_n1271;
  assign new_n1283 = new_n1282 ^ new_n1267;
  assign new_n1284 = new_n1283 ^ new_n1264;
  assign new_n1285 = new_n1262 ^ new_n1251;
  assign new_n1286 = new_n1285 ^ new_n1240;
  assign new_n1287 = new_n1226 & new_n1286;
  assign new_n1288 = new_n1287 ^ new_n1284;
  assign new_n1289 = new_n1260 ^ new_n1236;
  assign new_n1290 = ~new_n1193 & ~new_n1289;
  assign new_n1291 = ~new_n1266 & new_n1216;
  assign new_n1292 = new_n1291 ^ new_n1290;
  assign new_n1293 = ~new_n1204 & ~new_n1289;
  assign new_n1294 = new_n1293 ^ new_n1292;
  assign new_n1295 = new_n1294 ^ new_n1288;
  assign new_n1296 = n19 ^ n18;
  assign new_n1297 = new_n1296 ^ n24;
  assign new_n1298 = n19 ^ n17;
  assign new_n1299 = ~new_n1296 & n24;
  assign new_n1300 = ~n24 & n20;
  assign new_n1301 = new_n1300 ^ new_n1299;
  assign new_n1302 = new_n1301 ^ n20;
  assign new_n1303 = n20 ^ n17;
  assign new_n1304 = n23 ^ n21;
  assign new_n1305 = new_n1304 ^ new_n1303;
  assign new_n1306 = new_n1305 ^ n24;
  assign new_n1307 = new_n1297 ^ n23;
  assign new_n1308 = n22 ^ n17;
  assign new_n1309 = new_n1308 ^ new_n1307;
  assign new_n1310 = new_n1306 & new_n1309;
  assign new_n1311 = new_n1310 ^ new_n1302;
  assign new_n1312 = n20 ^ n19;
  assign new_n1313 = new_n1312 ^ new_n1308;
  assign new_n1314 = n22 ^ n20;
  assign new_n1315 = new_n1313 & new_n1314;
  assign new_n1316 = new_n1305 ^ new_n1296;
  assign new_n1317 = new_n1308 & new_n1316;
  assign new_n1318 = new_n1317 ^ new_n1315;
  assign new_n1319 = new_n1318 ^ new_n1311;
  assign new_n1320 = new_n1319 ^ new_n1298;
  assign new_n1321 = ~n23 & ~new_n1297;
  assign new_n1322 = new_n1321 ^ n23;
  assign new_n1323 = n22 ^ n21;
  assign new_n1324 = new_n1323 ^ n23;
  assign new_n1325 = new_n1324 ^ n19;
  assign new_n1326 = n23 ^ n17;
  assign new_n1327 = new_n1325 & new_n1326;
  assign new_n1328 = new_n1327 ^ new_n1322;
  assign new_n1329 = new_n1328 ^ new_n1308;
  assign new_n1330 = new_n1324 ^ n18;
  assign new_n1331 = new_n1303 & new_n1330;
  assign new_n1332 = new_n1331 ^ new_n1315;
  assign new_n1333 = n21 ^ n19;
  assign new_n1334 = new_n1333 ^ new_n1332;
  assign new_n1335 = new_n1334 ^ new_n1329;
  assign new_n1336 = n23 ^ n20;
  assign new_n1337 = new_n1336 ^ new_n1308;
  assign new_n1338 = new_n1305 & new_n1337;
  assign new_n1339 = new_n1338 ^ n18;
  assign new_n1340 = new_n1339 ^ new_n1305;
  assign new_n1341 = new_n1331 ^ new_n1310;
  assign new_n1342 = new_n1315 ^ n22;
  assign new_n1343 = new_n1342 ^ new_n1341;
  assign new_n1344 = new_n1343 ^ new_n1340;
  assign new_n1345 = ~new_n1335 & new_n1344;
  assign new_n1346 = new_n1330 ^ n24;
  assign new_n1347 = new_n1297 ^ n17;
  assign new_n1348 = new_n1346 & new_n1347;
  assign new_n1349 = new_n1348 ^ new_n1327;
  assign new_n1350 = new_n1349 ^ n17;
  assign new_n1351 = new_n1331 ^ new_n1317;
  assign new_n1352 = new_n1351 ^ new_n1325;
  assign new_n1353 = new_n1352 ^ new_n1350;
  assign new_n1354 = new_n1353 ^ new_n1345;
  assign new_n1355 = new_n1320 & new_n1354;
  assign new_n1356 = new_n1339 ^ new_n1301;
  assign new_n1357 = new_n1356 ^ new_n1355;
  assign new_n1358 = new_n1357 ^ new_n1352;
  assign new_n1359 = new_n1356 ^ new_n1345;
  assign new_n1360 = new_n1359 ^ new_n1352;
  assign new_n1361 = new_n1348 ^ new_n1321;
  assign new_n1362 = new_n1361 ^ new_n1318;
  assign new_n1363 = ~new_n1362 & new_n1360;
  assign new_n1364 = new_n1363 ^ new_n1345;
  assign new_n1365 = new_n1353 & new_n1364;
  assign new_n1366 = new_n1365 ^ new_n1354;
  assign new_n1367 = new_n1358 & new_n1366;
  assign new_n1368 = new_n1367 ^ new_n1320;
  assign new_n1369 = new_n1297 & new_n1368;
  assign new_n1370 = n23 ^ n19;
  assign new_n1371 = new_n1322 ^ new_n1310;
  assign new_n1372 = new_n1367 ^ new_n1365;
  assign new_n1373 = new_n1372 ^ new_n1371;
  assign new_n1374 = new_n1373 ^ new_n1370;
  assign new_n1375 = new_n1374 ^ n20;
  assign new_n1376 = new_n1355 ^ new_n1327;
  assign new_n1377 = new_n1376 ^ new_n1339;
  assign new_n1378 = new_n1377 ^ new_n1375;
  assign new_n1379 = ~new_n1378 & new_n1314;
  assign new_n1380 = new_n1363 ^ new_n1355;
  assign new_n1381 = new_n1356 ^ new_n1350;
  assign new_n1382 = new_n1381 ^ new_n1380;
  assign new_n1383 = new_n1303 & new_n1382;
  assign new_n1384 = new_n1383 ^ new_n1379;
  assign new_n1385 = new_n1365 ^ new_n1363;
  assign new_n1386 = new_n1385 ^ new_n1362;
  assign new_n1387 = ~new_n1386 & new_n1309;
  assign new_n1388 = new_n1387 ^ new_n1384;
  assign new_n1389 = new_n1388 ^ new_n1369;
  assign new_n1390 = new_n1367 ^ new_n1355;
  assign new_n1391 = new_n1390 ^ new_n1344;
  assign new_n1392 = new_n1325 & new_n1391;
  assign new_n1393 = new_n1392 ^ new_n1389;
  assign new_n1394 = new_n1365 ^ new_n1335;
  assign new_n1395 = ~new_n1394 & new_n1337;
  assign new_n1396 = ~new_n1386 & new_n1306;
  assign new_n1397 = ~new_n1394 & new_n1305;
  assign new_n1398 = new_n1397 ^ new_n1396;
  assign new_n1399 = new_n1398 ^ new_n1395;
  assign new_n1400 = new_n1399 ^ new_n1393;
  assign new_n1401 = new_n1400 ^ new_n1295;
  assign new_n1402 = new_n1401 ^ n124;
  assign new_n1403 = new_n1402 ^ n60;
  assign new_n1404 = n210 ^ n82;
  assign new_n1405 = n214 ^ n86;
  assign new_n1406 = n215 ^ n87;
  assign new_n1407 = n213 ^ n85;
  assign new_n1408 = new_n1407 ^ new_n1406;
  assign new_n1409 = new_n1408 ^ new_n1405;
  assign new_n1410 = new_n1409 ^ new_n1404;
  assign new_n1411 = n216 ^ n88;
  assign new_n1412 = new_n1411 ^ new_n1410;
  assign new_n1413 = n211 ^ n83;
  assign new_n1414 = n209 ^ n81;
  assign new_n1415 = new_n1414 ^ new_n1413;
  assign new_n1416 = new_n1413 ^ new_n1404;
  assign new_n1417 = ~new_n1416 & new_n1411;
  assign new_n1418 = n212 ^ n84;
  assign new_n1419 = ~new_n1411 & new_n1418;
  assign new_n1420 = new_n1419 ^ new_n1417;
  assign new_n1421 = new_n1420 ^ new_n1418;
  assign new_n1422 = new_n1418 ^ new_n1414;
  assign new_n1423 = new_n1422 ^ new_n1408;
  assign new_n1424 = new_n1423 ^ new_n1411;
  assign new_n1425 = new_n1416 ^ new_n1411;
  assign new_n1426 = new_n1425 ^ new_n1406;
  assign new_n1427 = new_n1414 ^ new_n1405;
  assign new_n1428 = new_n1427 ^ new_n1426;
  assign new_n1429 = new_n1424 & new_n1428;
  assign new_n1430 = new_n1429 ^ new_n1421;
  assign new_n1431 = new_n1418 ^ new_n1413;
  assign new_n1432 = new_n1431 ^ new_n1427;
  assign new_n1433 = new_n1418 ^ new_n1405;
  assign new_n1434 = new_n1432 & new_n1433;
  assign new_n1435 = new_n1423 ^ new_n1416;
  assign new_n1436 = new_n1427 & new_n1435;
  assign new_n1437 = new_n1436 ^ new_n1434;
  assign new_n1438 = new_n1437 ^ new_n1430;
  assign new_n1439 = new_n1438 ^ new_n1415;
  assign new_n1440 = ~new_n1406 & ~new_n1425;
  assign new_n1441 = new_n1440 ^ new_n1406;
  assign new_n1442 = new_n1413 ^ new_n1409;
  assign new_n1443 = new_n1414 ^ new_n1406;
  assign new_n1444 = new_n1442 & new_n1443;
  assign new_n1445 = new_n1444 ^ new_n1441;
  assign new_n1446 = new_n1445 ^ new_n1427;
  assign new_n1447 = new_n1410 & new_n1422;
  assign new_n1448 = new_n1447 ^ new_n1434;
  assign new_n1449 = new_n1413 ^ new_n1407;
  assign new_n1450 = new_n1449 ^ new_n1448;
  assign new_n1451 = new_n1450 ^ new_n1446;
  assign new_n1452 = new_n1418 ^ new_n1406;
  assign new_n1453 = new_n1452 ^ new_n1427;
  assign new_n1454 = new_n1423 & new_n1453;
  assign new_n1455 = new_n1454 ^ new_n1404;
  assign new_n1456 = new_n1455 ^ new_n1423;
  assign new_n1457 = new_n1429 ^ new_n1405;
  assign new_n1458 = new_n1457 ^ new_n1448;
  assign new_n1459 = new_n1458 ^ new_n1456;
  assign new_n1460 = ~new_n1451 & new_n1459;
  assign new_n1461 = new_n1447 ^ new_n1436;
  assign new_n1462 = new_n1461 ^ new_n1442;
  assign new_n1463 = new_n1425 ^ new_n1414;
  assign new_n1464 = new_n1412 & new_n1463;
  assign new_n1465 = new_n1464 ^ new_n1444;
  assign new_n1466 = new_n1465 ^ new_n1414;
  assign new_n1467 = new_n1466 ^ new_n1462;
  assign new_n1468 = new_n1467 ^ new_n1460;
  assign new_n1469 = new_n1439 & new_n1468;
  assign new_n1470 = new_n1455 ^ new_n1420;
  assign new_n1471 = new_n1470 ^ new_n1469;
  assign new_n1472 = new_n1471 ^ new_n1462;
  assign new_n1473 = new_n1412 & new_n1472;
  assign new_n1474 = new_n1470 ^ new_n1460;
  assign new_n1475 = new_n1474 ^ new_n1462;
  assign new_n1476 = new_n1464 ^ new_n1440;
  assign new_n1477 = new_n1476 ^ new_n1437;
  assign new_n1478 = ~new_n1477 & new_n1475;
  assign new_n1479 = new_n1478 ^ new_n1460;
  assign new_n1480 = ~new_n1479 & new_n1467;
  assign new_n1481 = new_n1480 ^ new_n1467;
  assign new_n1482 = new_n1481 ^ new_n1451;
  assign new_n1483 = ~new_n1482 & new_n1453;
  assign new_n1484 = new_n1483 ^ new_n1473;
  assign new_n1485 = new_n1478 ^ new_n1467;
  assign new_n1486 = new_n1411 & new_n1485;
  assign new_n1487 = new_n1481 ^ new_n1478;
  assign new_n1488 = new_n1487 ^ new_n1477;
  assign new_n1489 = ~new_n1488 & new_n1424;
  assign new_n1490 = new_n1489 ^ new_n1486;
  assign new_n1491 = new_n1480 ^ new_n1460;
  assign new_n1492 = new_n1472 & new_n1491;
  assign new_n1493 = new_n1492 ^ new_n1439;
  assign new_n1494 = new_n1425 & new_n1493;
  assign new_n1495 = ~new_n1488 & new_n1428;
  assign new_n1496 = new_n1413 ^ new_n1406;
  assign new_n1497 = new_n1441 ^ new_n1429;
  assign new_n1498 = new_n1492 ^ new_n1481;
  assign new_n1499 = new_n1498 ^ new_n1497;
  assign new_n1500 = new_n1499 ^ new_n1496;
  assign new_n1501 = new_n1500 ^ new_n1418;
  assign new_n1502 = new_n1469 ^ new_n1444;
  assign new_n1503 = new_n1502 ^ new_n1455;
  assign new_n1504 = new_n1503 ^ new_n1501;
  assign new_n1505 = ~new_n1504 & new_n1433;
  assign new_n1506 = new_n1478 ^ new_n1469;
  assign new_n1507 = new_n1470 ^ new_n1466;
  assign new_n1508 = new_n1507 ^ new_n1506;
  assign new_n1509 = new_n1422 & new_n1508;
  assign new_n1510 = new_n1509 ^ new_n1505;
  assign new_n1511 = new_n1510 ^ new_n1495;
  assign new_n1512 = new_n1511 ^ new_n1494;
  assign new_n1513 = new_n1512 ^ new_n1490;
  assign new_n1514 = new_n1513 ^ new_n1484;
  assign new_n1515 = new_n1514 ^ n109;
  assign new_n1516 = new_n1515 ^ new_n881;
  assign new_n1517 = n135 ^ n7;
  assign new_n1518 = n136 ^ n8;
  assign new_n1519 = n131 ^ n3;
  assign new_n1520 = n130 ^ n2;
  assign new_n1521 = new_n1520 ^ new_n1519;
  assign new_n1522 = new_n1521 ^ new_n1518;
  assign new_n1523 = ~new_n1517 & ~new_n1522;
  assign new_n1524 = new_n1523 ^ new_n1517;
  assign new_n1525 = n129 ^ n1;
  assign new_n1526 = new_n1525 ^ new_n1517;
  assign new_n1527 = n133 ^ n5;
  assign new_n1528 = new_n1527 ^ new_n1517;
  assign new_n1529 = n134 ^ n6;
  assign new_n1530 = new_n1529 ^ new_n1528;
  assign new_n1531 = new_n1530 ^ new_n1519;
  assign new_n1532 = new_n1526 & new_n1531;
  assign new_n1533 = new_n1532 ^ new_n1524;
  assign new_n1534 = new_n1529 ^ new_n1525;
  assign new_n1535 = new_n1534 ^ new_n1533;
  assign new_n1536 = new_n1530 ^ new_n1520;
  assign new_n1537 = n132 ^ n4;
  assign new_n1538 = new_n1537 ^ new_n1525;
  assign new_n1539 = new_n1536 & new_n1538;
  assign new_n1540 = new_n1537 ^ new_n1519;
  assign new_n1541 = new_n1540 ^ new_n1534;
  assign new_n1542 = new_n1537 ^ new_n1529;
  assign new_n1543 = new_n1541 & new_n1542;
  assign new_n1544 = new_n1543 ^ new_n1539;
  assign new_n1545 = new_n1527 ^ new_n1519;
  assign new_n1546 = new_n1545 ^ new_n1544;
  assign new_n1547 = new_n1546 ^ new_n1535;
  assign new_n1548 = new_n1538 ^ new_n1528;
  assign new_n1549 = new_n1537 ^ new_n1517;
  assign new_n1550 = new_n1549 ^ new_n1534;
  assign new_n1551 = new_n1548 & new_n1550;
  assign new_n1552 = new_n1551 ^ new_n1520;
  assign new_n1553 = new_n1552 ^ new_n1548;
  assign new_n1554 = new_n1548 ^ new_n1518;
  assign new_n1555 = new_n1522 ^ new_n1517;
  assign new_n1556 = new_n1555 ^ new_n1534;
  assign new_n1557 = new_n1554 & new_n1556;
  assign new_n1558 = new_n1557 ^ new_n1529;
  assign new_n1559 = new_n1558 ^ new_n1544;
  assign new_n1560 = new_n1559 ^ new_n1553;
  assign new_n1561 = ~new_n1547 & new_n1560;
  assign new_n1562 = ~new_n1521 & new_n1518;
  assign new_n1563 = ~new_n1518 & new_n1537;
  assign new_n1564 = new_n1563 ^ new_n1562;
  assign new_n1565 = new_n1564 ^ new_n1552;
  assign new_n1566 = new_n1565 ^ new_n1561;
  assign new_n1567 = new_n1548 ^ new_n1521;
  assign new_n1568 = new_n1534 & new_n1567;
  assign new_n1569 = new_n1568 ^ new_n1539;
  assign new_n1570 = new_n1569 ^ new_n1531;
  assign new_n1571 = new_n1570 ^ new_n1566;
  assign new_n1572 = new_n1525 ^ new_n1522;
  assign new_n1573 = new_n1536 ^ new_n1518;
  assign new_n1574 = new_n1572 & new_n1573;
  assign new_n1575 = new_n1574 ^ new_n1523;
  assign new_n1576 = new_n1568 ^ new_n1543;
  assign new_n1577 = new_n1576 ^ new_n1575;
  assign new_n1578 = ~new_n1577 & new_n1571;
  assign new_n1579 = new_n1574 ^ new_n1532;
  assign new_n1580 = new_n1579 ^ new_n1525;
  assign new_n1581 = new_n1580 ^ new_n1570;
  assign new_n1582 = new_n1581 ^ new_n1578;
  assign new_n1583 = new_n1537 ^ new_n1522;
  assign new_n1584 = new_n1582 & new_n1583;
  assign new_n1585 = new_n1519 ^ new_n1517;
  assign new_n1586 = new_n1557 ^ new_n1524;
  assign new_n1587 = new_n1525 ^ new_n1519;
  assign new_n1588 = new_n1564 ^ new_n1537;
  assign new_n1589 = new_n1588 ^ new_n1557;
  assign new_n1590 = new_n1589 ^ new_n1576;
  assign new_n1591 = new_n1590 ^ new_n1587;
  assign new_n1592 = new_n1581 ^ new_n1561;
  assign new_n1593 = new_n1591 & new_n1592;
  assign new_n1594 = new_n1593 ^ new_n1565;
  assign new_n1595 = new_n1594 ^ new_n1570;
  assign new_n1596 = new_n1578 ^ new_n1561;
  assign new_n1597 = new_n1581 & new_n1596;
  assign new_n1598 = new_n1597 ^ new_n1592;
  assign new_n1599 = new_n1595 & new_n1598;
  assign new_n1600 = new_n1599 ^ new_n1597;
  assign new_n1601 = new_n1600 ^ new_n1586;
  assign new_n1602 = new_n1601 ^ new_n1585;
  assign new_n1603 = new_n1602 ^ new_n1537;
  assign new_n1604 = new_n1593 ^ new_n1532;
  assign new_n1605 = new_n1604 ^ new_n1552;
  assign new_n1606 = new_n1605 ^ new_n1603;
  assign new_n1607 = ~new_n1606 & new_n1541;
  assign new_n1608 = new_n1597 ^ new_n1578;
  assign new_n1609 = new_n1608 ^ new_n1577;
  assign new_n1610 = ~new_n1609 & new_n1556;
  assign new_n1611 = ~new_n1606 & new_n1542;
  assign new_n1612 = new_n1593 ^ new_n1578;
  assign new_n1613 = new_n1580 ^ new_n1565;
  assign new_n1614 = new_n1613 ^ new_n1612;
  assign new_n1615 = new_n1538 & new_n1614;
  assign new_n1616 = new_n1615 ^ new_n1611;
  assign new_n1617 = new_n1616 ^ new_n1610;
  assign new_n1618 = new_n1599 ^ new_n1591;
  assign new_n1619 = new_n1522 & new_n1618;
  assign new_n1620 = new_n1619 ^ new_n1617;
  assign new_n1621 = new_n1599 ^ new_n1593;
  assign new_n1622 = new_n1621 ^ new_n1560;
  assign new_n1623 = new_n1531 & new_n1622;
  assign new_n1624 = new_n1623 ^ new_n1620;
  assign new_n1625 = new_n1624 ^ new_n1607;
  assign new_n1626 = new_n1625 ^ new_n1584;
  assign new_n1627 = new_n1572 & new_n1595;
  assign new_n1628 = new_n1578 ^ new_n1525;
  assign new_n1629 = new_n1588 ^ new_n1574;
  assign new_n1630 = new_n1629 ^ new_n1602;
  assign new_n1631 = new_n1630 ^ new_n1628;
  assign new_n1632 = ~new_n1631 & new_n1567;
  assign new_n1633 = new_n1632 ^ new_n1627;
  assign new_n1634 = new_n1597 ^ new_n1547;
  assign new_n1635 = ~new_n1634 & new_n1548;
  assign new_n1636 = new_n1518 & new_n1582;
  assign new_n1637 = new_n1636 ^ new_n1635;
  assign new_n1638 = new_n1526 & new_n1622;
  assign new_n1639 = new_n1638 ^ new_n1637;
  assign new_n1640 = new_n1639 ^ new_n1633;
  assign new_n1641 = new_n1640 ^ new_n1626;
  assign new_n1642 = n170 ^ n42;
  assign new_n1643 = n171 ^ n43;
  assign new_n1644 = new_n1643 ^ new_n1642;
  assign new_n1645 = n176 ^ n48;
  assign new_n1646 = new_n1645 ^ new_n1644;
  assign new_n1647 = n172 ^ n44;
  assign new_n1648 = new_n1647 ^ new_n1646;
  assign new_n1649 = new_n1645 & new_n1648;
  assign new_n1650 = new_n1649 ^ new_n1647;
  assign new_n1651 = n169 ^ n41;
  assign new_n1652 = new_n1651 ^ new_n1647;
  assign new_n1653 = n175 ^ n47;
  assign new_n1654 = n173 ^ n45;
  assign new_n1655 = new_n1654 ^ new_n1653;
  assign new_n1656 = new_n1655 ^ new_n1652;
  assign new_n1657 = new_n1653 ^ new_n1647;
  assign new_n1658 = n174 ^ n46;
  assign new_n1659 = new_n1658 ^ new_n1651;
  assign new_n1660 = new_n1659 ^ new_n1657;
  assign new_n1661 = new_n1656 & new_n1660;
  assign new_n1662 = new_n1661 ^ new_n1642;
  assign new_n1663 = new_n1662 ^ new_n1650;
  assign new_n1664 = new_n1653 ^ new_n1651;
  assign new_n1665 = new_n1658 ^ new_n1655;
  assign new_n1666 = new_n1665 ^ new_n1643;
  assign new_n1667 = new_n1664 & new_n1666;
  assign new_n1668 = ~new_n1646 & ~new_n1653;
  assign new_n1669 = new_n1668 ^ new_n1653;
  assign new_n1670 = new_n1669 ^ new_n1667;
  assign new_n1671 = new_n1670 ^ new_n1659;
  assign new_n1672 = new_n1665 ^ new_n1642;
  assign new_n1673 = new_n1652 & new_n1672;
  assign new_n1674 = new_n1647 ^ new_n1643;
  assign new_n1675 = new_n1674 ^ new_n1659;
  assign new_n1676 = new_n1658 ^ new_n1647;
  assign new_n1677 = new_n1675 & new_n1676;
  assign new_n1678 = new_n1677 ^ new_n1673;
  assign new_n1679 = new_n1654 ^ new_n1643;
  assign new_n1680 = new_n1679 ^ new_n1678;
  assign new_n1681 = new_n1680 ^ new_n1671;
  assign new_n1682 = new_n1662 ^ new_n1656;
  assign new_n1683 = new_n1656 ^ new_n1645;
  assign new_n1684 = new_n1653 ^ new_n1646;
  assign new_n1685 = new_n1684 ^ new_n1659;
  assign new_n1686 = new_n1683 & new_n1685;
  assign new_n1687 = new_n1686 ^ new_n1658;
  assign new_n1688 = new_n1687 ^ new_n1678;
  assign new_n1689 = new_n1688 ^ new_n1682;
  assign new_n1690 = ~new_n1681 & new_n1689;
  assign new_n1691 = new_n1690 ^ new_n1663;
  assign new_n1692 = new_n1656 ^ new_n1644;
  assign new_n1693 = new_n1659 & new_n1692;
  assign new_n1694 = new_n1693 ^ new_n1673;
  assign new_n1695 = new_n1694 ^ new_n1666;
  assign new_n1696 = new_n1695 ^ new_n1691;
  assign new_n1697 = new_n1693 ^ new_n1677;
  assign new_n1698 = new_n1651 ^ new_n1646;
  assign new_n1699 = new_n1672 ^ new_n1645;
  assign new_n1700 = new_n1698 & new_n1699;
  assign new_n1701 = new_n1700 ^ new_n1668;
  assign new_n1702 = new_n1701 ^ new_n1697;
  assign new_n1703 = ~new_n1702 & new_n1696;
  assign new_n1704 = new_n1700 ^ new_n1667;
  assign new_n1705 = new_n1704 ^ new_n1651;
  assign new_n1706 = new_n1705 ^ new_n1695;
  assign new_n1707 = new_n1706 ^ new_n1703;
  assign new_n1708 = new_n1648 & new_n1707;
  assign new_n1709 = new_n1653 ^ new_n1643;
  assign new_n1710 = new_n1686 ^ new_n1669;
  assign new_n1711 = new_n1703 ^ new_n1690;
  assign new_n1712 = ~new_n1706 & ~new_n1711;
  assign new_n1713 = new_n1712 ^ new_n1703;
  assign new_n1714 = new_n1706 ^ new_n1690;
  assign new_n1715 = new_n1651 ^ new_n1643;
  assign new_n1716 = new_n1686 ^ new_n1649;
  assign new_n1717 = new_n1716 ^ new_n1697;
  assign new_n1718 = new_n1717 ^ new_n1715;
  assign new_n1719 = new_n1714 & new_n1718;
  assign new_n1720 = new_n1719 ^ new_n1663;
  assign new_n1721 = new_n1720 ^ new_n1695;
  assign new_n1722 = ~new_n1713 & new_n1721;
  assign new_n1723 = new_n1714 ^ new_n1713;
  assign new_n1724 = new_n1723 ^ new_n1722;
  assign new_n1725 = new_n1724 ^ new_n1710;
  assign new_n1726 = new_n1725 ^ new_n1709;
  assign new_n1727 = new_n1726 ^ new_n1647;
  assign new_n1728 = new_n1719 ^ new_n1667;
  assign new_n1729 = new_n1728 ^ new_n1662;
  assign new_n1730 = new_n1729 ^ new_n1727;
  assign new_n1731 = new_n1675 & new_n1730;
  assign new_n1732 = new_n1722 ^ new_n1718;
  assign new_n1733 = new_n1646 & new_n1732;
  assign new_n1734 = new_n1676 & new_n1730;
  assign new_n1735 = new_n1719 ^ new_n1703;
  assign new_n1736 = new_n1705 ^ new_n1663;
  assign new_n1737 = new_n1736 ^ new_n1735;
  assign new_n1738 = new_n1652 & new_n1737;
  assign new_n1739 = new_n1738 ^ new_n1734;
  assign new_n1740 = new_n1723 ^ new_n1703;
  assign new_n1741 = new_n1740 ^ new_n1702;
  assign new_n1742 = new_n1685 & new_n1741;
  assign new_n1743 = new_n1742 ^ new_n1739;
  assign new_n1744 = new_n1743 ^ new_n1733;
  assign new_n1745 = new_n1722 ^ new_n1719;
  assign new_n1746 = new_n1745 ^ new_n1689;
  assign new_n1747 = new_n1666 & new_n1746;
  assign new_n1748 = new_n1747 ^ new_n1744;
  assign new_n1749 = new_n1748 ^ new_n1731;
  assign new_n1750 = new_n1749 ^ new_n1708;
  assign new_n1751 = new_n1664 & new_n1746;
  assign new_n1752 = new_n1645 & new_n1707;
  assign new_n1753 = new_n1723 ^ new_n1681;
  assign new_n1754 = new_n1656 & new_n1753;
  assign new_n1755 = new_n1754 ^ new_n1752;
  assign new_n1756 = new_n1755 ^ new_n1751;
  assign new_n1757 = new_n1703 ^ new_n1651;
  assign new_n1758 = new_n1700 ^ new_n1649;
  assign new_n1759 = new_n1758 ^ new_n1726;
  assign new_n1760 = new_n1759 ^ new_n1757;
  assign new_n1761 = new_n1692 & new_n1760;
  assign new_n1762 = new_n1698 & new_n1721;
  assign new_n1763 = new_n1762 ^ new_n1761;
  assign new_n1764 = new_n1763 ^ new_n1756;
  assign new_n1765 = new_n1764 ^ new_n1750;
  assign new_n1766 = new_n1765 ^ new_n1641;
  assign new_n1767 = new_n1672 & new_n1737;
  assign new_n1768 = new_n1660 & new_n1753;
  assign new_n1769 = new_n1768 ^ new_n1767;
  assign new_n1770 = new_n1769 ^ new_n1749;
  assign new_n1771 = ~new_n1634 & new_n1550;
  assign new_n1772 = new_n1536 & new_n1614;
  assign new_n1773 = new_n1772 ^ new_n1771;
  assign new_n1774 = new_n1773 ^ new_n1625;
  assign new_n1775 = new_n1774 ^ new_n1770;
  assign new_n1776 = new_n1775 ^ new_n1766;
  assign new_n1777 = n250 ^ n122;
  assign new_n1778 = n254 ^ n126;
  assign new_n1779 = n255 ^ n127;
  assign new_n1780 = n253 ^ n125;
  assign new_n1781 = new_n1780 ^ new_n1779;
  assign new_n1782 = new_n1781 ^ new_n1778;
  assign new_n1783 = new_n1782 ^ new_n1777;
  assign new_n1784 = n256 ^ n128;
  assign new_n1785 = new_n1784 ^ new_n1783;
  assign new_n1786 = n251 ^ n123;
  assign new_n1787 = new_n1786 ^ new_n1777;
  assign new_n1788 = new_n1787 ^ new_n1784;
  assign new_n1789 = ~new_n1779 & new_n1788;
  assign new_n1790 = new_n1786 ^ new_n1782;
  assign new_n1791 = n249 ^ n121;
  assign new_n1792 = new_n1791 ^ new_n1779;
  assign new_n1793 = new_n1790 & new_n1792;
  assign new_n1794 = new_n1793 ^ new_n1789;
  assign new_n1795 = new_n1791 ^ new_n1778;
  assign new_n1796 = new_n1795 ^ new_n1794;
  assign new_n1797 = n252 ^ n124;
  assign new_n1798 = new_n1797 ^ new_n1786;
  assign new_n1799 = new_n1798 ^ new_n1795;
  assign new_n1800 = new_n1797 ^ new_n1778;
  assign new_n1801 = new_n1799 & new_n1800;
  assign new_n1802 = new_n1797 ^ new_n1791;
  assign new_n1803 = new_n1783 & new_n1802;
  assign new_n1804 = new_n1803 ^ new_n1801;
  assign new_n1805 = new_n1786 ^ new_n1780;
  assign new_n1806 = new_n1805 ^ new_n1804;
  assign new_n1807 = new_n1806 ^ new_n1796;
  assign new_n1808 = new_n1802 ^ new_n1781;
  assign new_n1809 = new_n1797 ^ new_n1779;
  assign new_n1810 = new_n1809 ^ new_n1795;
  assign new_n1811 = new_n1808 & new_n1810;
  assign new_n1812 = new_n1811 ^ new_n1777;
  assign new_n1813 = new_n1812 ^ new_n1808;
  assign new_n1814 = new_n1808 ^ new_n1784;
  assign new_n1815 = new_n1788 ^ new_n1779;
  assign new_n1816 = new_n1815 ^ new_n1795;
  assign new_n1817 = new_n1814 & new_n1816;
  assign new_n1818 = new_n1817 ^ new_n1778;
  assign new_n1819 = new_n1818 ^ new_n1804;
  assign new_n1820 = new_n1819 ^ new_n1813;
  assign new_n1821 = new_n1807 & new_n1820;
  assign new_n1822 = new_n1808 ^ new_n1787;
  assign new_n1823 = new_n1795 & new_n1822;
  assign new_n1824 = new_n1823 ^ new_n1803;
  assign new_n1825 = new_n1824 ^ new_n1790;
  assign new_n1826 = new_n1791 ^ new_n1788;
  assign new_n1827 = new_n1785 & new_n1826;
  assign new_n1828 = new_n1827 ^ new_n1793;
  assign new_n1829 = new_n1828 ^ new_n1791;
  assign new_n1830 = new_n1829 ^ new_n1825;
  assign new_n1831 = new_n1830 ^ new_n1821;
  assign new_n1832 = new_n1791 ^ new_n1786;
  assign new_n1833 = ~new_n1787 & new_n1784;
  assign new_n1834 = ~new_n1784 & new_n1797;
  assign new_n1835 = new_n1834 ^ new_n1833;
  assign new_n1836 = new_n1835 ^ new_n1797;
  assign new_n1837 = new_n1836 ^ new_n1817;
  assign new_n1838 = new_n1823 ^ new_n1801;
  assign new_n1839 = new_n1838 ^ new_n1837;
  assign new_n1840 = new_n1839 ^ new_n1832;
  assign new_n1841 = new_n1831 & new_n1840;
  assign new_n1842 = new_n1835 ^ new_n1812;
  assign new_n1843 = new_n1842 ^ new_n1841;
  assign new_n1844 = new_n1843 ^ new_n1825;
  assign new_n1845 = new_n1785 & new_n1844;
  assign new_n1846 = new_n1789 ^ new_n1779;
  assign new_n1847 = new_n1846 ^ new_n1827;
  assign new_n1848 = new_n1847 ^ new_n1838;
  assign new_n1849 = new_n1842 ^ new_n1821;
  assign new_n1850 = new_n1849 ^ new_n1825;
  assign new_n1851 = new_n1848 & new_n1850;
  assign new_n1852 = new_n1851 ^ new_n1821;
  assign new_n1853 = ~new_n1830 & ~new_n1852;
  assign new_n1854 = new_n1853 ^ new_n1851;
  assign new_n1855 = new_n1854 ^ new_n1831;
  assign new_n1856 = new_n1855 ^ new_n1807;
  assign new_n1857 = ~new_n1856 & new_n1810;
  assign new_n1858 = new_n1857 ^ new_n1845;
  assign new_n1859 = new_n1851 ^ new_n1830;
  assign new_n1860 = new_n1784 & new_n1859;
  assign new_n1861 = new_n1855 ^ new_n1851;
  assign new_n1862 = new_n1861 ^ new_n1848;
  assign new_n1863 = ~new_n1862 & new_n1814;
  assign new_n1864 = new_n1863 ^ new_n1860;
  assign new_n1865 = ~new_n1854 & new_n1844;
  assign new_n1866 = new_n1865 ^ new_n1840;
  assign new_n1867 = new_n1788 & new_n1866;
  assign new_n1868 = ~new_n1862 & new_n1816;
  assign new_n1869 = new_n1786 ^ new_n1779;
  assign new_n1870 = new_n1817 ^ new_n1789;
  assign new_n1871 = new_n1865 ^ new_n1855;
  assign new_n1872 = new_n1871 ^ new_n1870;
  assign new_n1873 = new_n1872 ^ new_n1869;
  assign new_n1874 = new_n1873 ^ new_n1797;
  assign new_n1875 = new_n1841 ^ new_n1793;
  assign new_n1876 = new_n1875 ^ new_n1812;
  assign new_n1877 = new_n1876 ^ new_n1874;
  assign new_n1878 = ~new_n1877 & new_n1800;
  assign new_n1879 = new_n1851 ^ new_n1841;
  assign new_n1880 = new_n1842 ^ new_n1829;
  assign new_n1881 = new_n1880 ^ new_n1879;
  assign new_n1882 = new_n1802 & new_n1881;
  assign new_n1883 = new_n1882 ^ new_n1878;
  assign new_n1884 = new_n1883 ^ new_n1868;
  assign new_n1885 = new_n1884 ^ new_n1867;
  assign new_n1886 = new_n1885 ^ new_n1864;
  assign new_n1887 = new_n1886 ^ new_n1858;
  assign new_n1888 = new_n1573 & new_n1595;
  assign new_n1889 = new_n1888 ^ new_n1771;
  assign new_n1890 = ~new_n1609 & new_n1554;
  assign new_n1891 = new_n1890 ^ new_n1636;
  assign new_n1892 = new_n1891 ^ new_n1620;
  assign new_n1893 = new_n1892 ^ new_n1889;
  assign new_n1894 = new_n1893 ^ new_n1887;
  assign new_n1895 = new_n1894 ^ new_n1776;
  assign new_n1896 = new_n1895 ^ new_n1516;
  assign new_n1897 = new_n1478 ^ new_n1414;
  assign new_n1898 = new_n1464 ^ new_n1421;
  assign new_n1899 = new_n1898 ^ new_n1500;
  assign new_n1900 = new_n1899 ^ new_n1897;
  assign new_n1901 = ~new_n1900 & new_n1435;
  assign new_n1902 = new_n1492 ^ new_n1469;
  assign new_n1903 = new_n1902 ^ new_n1459;
  assign new_n1904 = new_n1443 & new_n1903;
  assign new_n1905 = new_n1904 ^ new_n1901;
  assign new_n1906 = ~new_n1504 & new_n1432;
  assign new_n1907 = new_n1906 ^ new_n1494;
  assign new_n1908 = new_n1426 & new_n1493;
  assign new_n1909 = new_n1908 ^ new_n1473;
  assign new_n1910 = new_n1909 ^ new_n1510;
  assign new_n1911 = new_n1910 ^ new_n1907;
  assign new_n1912 = new_n1911 ^ new_n1905;
  assign new_n1913 = new_n1638 ^ new_n1632;
  assign new_n1914 = new_n1619 ^ new_n1607;
  assign new_n1915 = new_n1555 & new_n1618;
  assign new_n1916 = new_n1915 ^ new_n1888;
  assign new_n1917 = new_n1916 ^ new_n1616;
  assign new_n1918 = new_n1917 ^ new_n1914;
  assign new_n1919 = new_n1918 ^ new_n1913;
  assign new_n1920 = new_n1919 ^ new_n1912;
  assign new_n1921 = new_n1756 ^ new_n1747;
  assign new_n1922 = new_n1684 & new_n1732;
  assign new_n1923 = new_n1699 & new_n1721;
  assign new_n1924 = new_n1923 ^ new_n1922;
  assign new_n1925 = new_n1924 ^ new_n1739;
  assign new_n1926 = new_n1925 ^ new_n1921;
  assign new_n1927 = new_n1639 ^ new_n1623;
  assign new_n1928 = new_n1927 ^ new_n1917;
  assign new_n1929 = new_n1928 ^ new_n1926;
  assign new_n1930 = new_n1929 ^ new_n1775;
  assign new_n1931 = new_n1930 ^ new_n1920;
  assign new_n1932 = new_n1851 ^ new_n1791;
  assign new_n1933 = new_n1836 ^ new_n1827;
  assign new_n1934 = new_n1933 ^ new_n1873;
  assign new_n1935 = new_n1934 ^ new_n1932;
  assign new_n1936 = ~new_n1935 & new_n1822;
  assign new_n1937 = new_n1865 ^ new_n1841;
  assign new_n1938 = new_n1937 ^ new_n1820;
  assign new_n1939 = new_n1792 & new_n1938;
  assign new_n1940 = new_n1939 ^ new_n1936;
  assign new_n1941 = ~new_n1877 & new_n1799;
  assign new_n1942 = new_n1941 ^ new_n1867;
  assign new_n1943 = new_n1815 & new_n1866;
  assign new_n1944 = new_n1943 ^ new_n1845;
  assign new_n1945 = new_n1944 ^ new_n1883;
  assign new_n1946 = new_n1945 ^ new_n1942;
  assign new_n1947 = new_n1946 ^ new_n1940;
  assign new_n1948 = new_n1947 ^ new_n890;
  assign new_n1949 = new_n1948 ^ new_n1931;
  assign new_n1950 = new_n1949 ^ new_n1896;
  assign new_n1951 = new_n1923 ^ new_n1768;
  assign new_n1952 = new_n1683 & new_n1741;
  assign new_n1953 = new_n1952 ^ new_n1752;
  assign new_n1954 = new_n1953 ^ new_n1744;
  assign new_n1955 = new_n1954 ^ new_n1951;
  assign new_n1956 = new_n1955 ^ new_n1893;
  assign new_n1957 = new_n1956 ^ new_n1775;
  assign new_n1958 = new_n1890 ^ new_n1635;
  assign new_n1959 = new_n1958 ^ new_n1771;
  assign new_n1960 = new_n1959 ^ new_n1624;
  assign new_n1961 = new_n1790 & new_n1938;
  assign new_n1962 = new_n1961 ^ new_n1885;
  assign new_n1963 = ~new_n1856 & new_n1808;
  assign new_n1964 = new_n1963 ^ new_n1863;
  assign new_n1965 = new_n1964 ^ new_n1857;
  assign new_n1966 = new_n1965 ^ new_n1962;
  assign new_n1967 = new_n1966 ^ new_n1960;
  assign new_n1968 = new_n1967 ^ new_n1957;
  assign new_n1969 = new_n1442 & new_n1903;
  assign new_n1970 = new_n1969 ^ new_n1512;
  assign new_n1971 = ~new_n1482 & new_n1423;
  assign new_n1972 = new_n1971 ^ new_n1489;
  assign new_n1973 = new_n1972 ^ new_n1483;
  assign new_n1974 = new_n1973 ^ new_n1970;
  assign new_n1975 = new_n1974 ^ n108;
  assign new_n1976 = new_n1975 ^ new_n862;
  assign new_n1977 = new_n1976 ^ new_n1968;
  assign new_n1978 = new_n1767 ^ new_n1731;
  assign new_n1979 = new_n1952 ^ new_n1754;
  assign new_n1980 = new_n1979 ^ new_n1768;
  assign new_n1981 = new_n1980 ^ new_n1743;
  assign new_n1982 = new_n1981 ^ new_n1978;
  assign new_n1983 = new_n1772 ^ new_n1607;
  assign new_n1984 = new_n1959 ^ new_n1617;
  assign new_n1985 = new_n1984 ^ new_n1983;
  assign new_n1986 = new_n1985 ^ new_n1982;
  assign new_n1987 = new_n1962 ^ new_n1941;
  assign new_n1988 = new_n1783 & new_n1881;
  assign new_n1989 = new_n1988 ^ new_n1857;
  assign new_n1990 = new_n1989 ^ new_n1987;
  assign new_n1991 = new_n1990 ^ new_n1774;
  assign new_n1992 = new_n1991 ^ new_n1986;
  assign new_n1993 = new_n1970 ^ new_n1906;
  assign new_n1994 = new_n1410 & new_n1508;
  assign new_n1995 = new_n1994 ^ new_n1483;
  assign new_n1996 = new_n1995 ^ new_n1993;
  assign new_n1997 = new_n1996 ^ n105;
  assign new_n1998 = new_n1997 ^ new_n872;
  assign new_n1999 = new_n1998 ^ new_n1992;
  assign new_n2000 = new_n1999 ^ new_n1977;
  assign new_n2001 = new_n2000 ^ new_n1950;
  assign new_n2002 = new_n1761 ^ new_n1751;
  assign new_n2003 = new_n1733 ^ new_n1731;
  assign new_n2004 = new_n2003 ^ new_n1925;
  assign new_n2005 = new_n2004 ^ new_n2002;
  assign new_n2006 = new_n2005 ^ new_n1919;
  assign new_n2007 = new_n1797 ^ new_n1788;
  assign new_n2008 = new_n1859 & new_n2007;
  assign new_n2009 = new_n2008 ^ new_n1987;
  assign new_n2010 = new_n1826 & new_n1844;
  assign new_n2011 = new_n2010 ^ new_n1936;
  assign new_n2012 = new_n1963 ^ new_n1860;
  assign new_n2013 = new_n2012 ^ new_n1939;
  assign new_n2014 = new_n2013 ^ new_n2011;
  assign new_n2015 = new_n2014 ^ new_n2009;
  assign new_n2016 = new_n2015 ^ new_n1641;
  assign new_n2017 = new_n2016 ^ new_n2006;
  assign new_n2018 = new_n1425 ^ new_n1418;
  assign new_n2019 = new_n1485 & new_n2018;
  assign new_n2020 = new_n2019 ^ new_n1993;
  assign new_n2021 = new_n1463 & new_n1472;
  assign new_n2022 = new_n2021 ^ new_n1901;
  assign new_n2023 = new_n1971 ^ new_n1486;
  assign new_n2024 = new_n2023 ^ new_n1904;
  assign new_n2025 = new_n2024 ^ new_n2022;
  assign new_n2026 = new_n2025 ^ new_n2020;
  assign new_n2027 = new_n2026 ^ n110;
  assign new_n2028 = new_n2027 ^ new_n900;
  assign new_n2029 = new_n2028 ^ new_n2017;
  assign new_n2030 = new_n2029 ^ new_n1950;
  assign new_n2031 = new_n1994 ^ new_n1906;
  assign new_n2032 = new_n1973 ^ new_n1511;
  assign new_n2033 = new_n2032 ^ new_n2031;
  assign new_n2034 = new_n2033 ^ new_n818;
  assign new_n2035 = new_n1772 ^ new_n1615;
  assign new_n2036 = ~new_n1631 & new_n1534;
  assign new_n2037 = new_n2036 ^ new_n1640;
  assign new_n2038 = new_n2037 ^ new_n2035;
  assign new_n2039 = new_n1767 ^ new_n1738;
  assign new_n2040 = new_n1659 & new_n1760;
  assign new_n2041 = new_n2040 ^ new_n1764;
  assign new_n2042 = new_n2041 ^ new_n2039;
  assign new_n2043 = new_n2042 ^ new_n2038;
  assign new_n2044 = new_n1988 ^ new_n1941;
  assign new_n2045 = new_n1965 ^ new_n1884;
  assign new_n2046 = new_n2045 ^ new_n2044;
  assign new_n2047 = new_n2046 ^ new_n1985;
  assign new_n2048 = new_n2047 ^ new_n2043;
  assign new_n2049 = new_n2048 ^ new_n2034;
  assign new_n2050 = new_n2049 ^ new_n2030;
  assign new_n2051 = new_n2000 & new_n2050;
  assign new_n2052 = new_n2029 ^ new_n1999;
  assign new_n2053 = new_n1994 ^ new_n1509;
  assign new_n2054 = ~new_n1900 & new_n1427;
  assign new_n2055 = new_n2054 ^ new_n2025;
  assign new_n2056 = new_n2055 ^ new_n2053;
  assign new_n2057 = new_n2056 ^ new_n841;
  assign new_n2058 = new_n1980 ^ new_n1748;
  assign new_n2059 = new_n2058 ^ new_n1960;
  assign new_n2060 = new_n1988 ^ new_n1882;
  assign new_n2061 = ~new_n1935 & new_n1795;
  assign new_n2062 = new_n2061 ^ new_n2014;
  assign new_n2063 = new_n2062 ^ new_n2060;
  assign new_n2064 = new_n2063 ^ new_n2038;
  assign new_n2065 = new_n2064 ^ new_n2059;
  assign new_n2066 = new_n2065 ^ new_n2057;
  assign new_n2067 = new_n2066 ^ new_n2049;
  assign new_n2068 = new_n2067 ^ new_n2001;
  assign new_n2069 = new_n2052 & new_n2068;
  assign new_n2070 = new_n2069 ^ new_n2051;
  assign new_n2071 = new_n2066 ^ new_n2030;
  assign new_n2072 = new_n2071 ^ new_n2070;
  assign new_n2073 = new_n1999 ^ new_n1949;
  assign new_n2074 = new_n2071 & new_n2073;
  assign new_n2075 = new_n2013 ^ new_n1961;
  assign new_n2076 = new_n2075 ^ new_n1945;
  assign new_n2077 = new_n2076 ^ new_n854;
  assign new_n2078 = new_n2024 ^ new_n1969;
  assign new_n2079 = new_n2078 ^ new_n1910;
  assign new_n2080 = new_n2079 ^ new_n1928;
  assign new_n2081 = new_n2080 ^ new_n1775;
  assign new_n2082 = new_n2081 ^ new_n2077;
  assign new_n2083 = new_n2082 ^ new_n2067;
  assign new_n2084 = new_n2083 ^ new_n1999;
  assign new_n2085 = new_n2082 ^ new_n2050;
  assign new_n2086 = new_n2084 & new_n2085;
  assign new_n2087 = new_n2086 ^ new_n2074;
  assign new_n2088 = new_n2087 ^ new_n1999;
  assign new_n2089 = new_n2088 ^ new_n2072;
  assign new_n2090 = new_n2083 ^ new_n1977;
  assign new_n2091 = new_n2082 & new_n2090;
  assign new_n2092 = new_n2091 ^ new_n1977;
  assign new_n2093 = new_n1977 ^ new_n1949;
  assign new_n2094 = new_n2093 ^ new_n2052;
  assign new_n2095 = new_n2001 & new_n2094;
  assign new_n2096 = new_n2095 ^ new_n2049;
  assign new_n2097 = new_n2096 ^ new_n2092;
  assign new_n2098 = ~new_n1949 & ~new_n2083;
  assign new_n2099 = new_n2098 ^ new_n1949;
  assign new_n2100 = new_n2099 ^ new_n2074;
  assign new_n2101 = new_n2100 ^ new_n2052;
  assign new_n2102 = new_n2029 ^ new_n1977;
  assign new_n2103 = new_n2066 ^ new_n1977;
  assign new_n2104 = new_n2103 ^ new_n2052;
  assign new_n2105 = new_n2102 & new_n2104;
  assign new_n2106 = new_n2105 ^ new_n2051;
  assign new_n2107 = new_n2066 ^ new_n1896;
  assign new_n2108 = new_n2107 ^ new_n2106;
  assign new_n2109 = new_n2108 ^ new_n2101;
  assign new_n2110 = new_n2096 ^ new_n2001;
  assign new_n2111 = new_n2082 ^ new_n2001;
  assign new_n2112 = new_n2083 ^ new_n1949;
  assign new_n2113 = new_n2112 ^ new_n2052;
  assign new_n2114 = new_n2111 & new_n2113;
  assign new_n2115 = new_n2114 ^ new_n2106;
  assign new_n2116 = new_n2115 ^ new_n2029;
  assign new_n2117 = new_n2116 ^ new_n2110;
  assign new_n2118 = ~new_n2109 & new_n2117;
  assign new_n2119 = new_n2118 ^ new_n2097;
  assign new_n2120 = new_n2119 ^ new_n2072;
  assign new_n2121 = new_n2098 ^ new_n2086;
  assign new_n2122 = new_n2105 ^ new_n2069;
  assign new_n2123 = new_n2122 ^ new_n2121;
  assign new_n2124 = ~new_n2123 & new_n2120;
  assign new_n2125 = new_n2124 ^ new_n2118;
  assign new_n2126 = new_n2089 & new_n2125;
  assign new_n2127 = new_n2126 ^ new_n2109;
  assign new_n2128 = ~new_n2127 & new_n2001;
  assign new_n2129 = new_n2126 ^ new_n2124;
  assign new_n2130 = new_n2129 ^ new_n2123;
  assign new_n2131 = ~new_n2130 & new_n2111;
  assign new_n2132 = new_n2131 ^ new_n2128;
  assign new_n2133 = ~new_n2127 & new_n2094;
  assign new_n2134 = new_n2133 ^ new_n2132;
  assign new_n2135 = new_n2066 ^ new_n1999;
  assign new_n2136 = new_n2114 ^ new_n2091;
  assign new_n2137 = new_n2136 ^ new_n2122;
  assign new_n2138 = new_n2137 ^ new_n2135;
  assign new_n2139 = new_n2118 ^ new_n2089;
  assign new_n2140 = new_n2138 & new_n2139;
  assign new_n2141 = new_n2140 ^ new_n2097;
  assign new_n2142 = new_n2141 ^ new_n2072;
  assign new_n2143 = new_n2139 ^ new_n2126;
  assign new_n2144 = new_n2142 & new_n2143;
  assign new_n2145 = new_n2144 ^ new_n2140;
  assign new_n2146 = new_n2145 ^ new_n2117;
  assign new_n2147 = new_n2071 & new_n2146;
  assign new_n2148 = ~new_n2130 & new_n2113;
  assign new_n2149 = new_n2140 ^ new_n2124;
  assign new_n2150 = new_n2097 ^ new_n2088;
  assign new_n2151 = new_n2150 ^ new_n2149;
  assign new_n2152 = new_n2000 & new_n2151;
  assign new_n2153 = new_n2066 ^ new_n1949;
  assign new_n2154 = new_n2114 ^ new_n2099;
  assign new_n2155 = new_n2144 ^ new_n2126;
  assign new_n2156 = new_n2155 ^ new_n2154;
  assign new_n2157 = new_n2156 ^ new_n2153;
  assign new_n2158 = new_n2157 ^ new_n1977;
  assign new_n2159 = new_n2140 ^ new_n2074;
  assign new_n2160 = new_n2159 ^ new_n2096;
  assign new_n2161 = new_n2160 ^ new_n2158;
  assign new_n2162 = ~new_n2161 & new_n2102;
  assign new_n2163 = new_n2162 ^ new_n2152;
  assign new_n2164 = new_n2163 ^ new_n2148;
  assign new_n2165 = new_n2144 ^ new_n2138;
  assign new_n2166 = new_n2083 & new_n2165;
  assign new_n2167 = new_n2166 ^ new_n2164;
  assign new_n2168 = new_n2167 ^ new_n2147;
  assign new_n2169 = new_n2168 ^ new_n2134;
  assign new_n2170 = n139 ^ n11;
  assign new_n2171 = n138 ^ n10;
  assign new_n2172 = new_n2171 ^ new_n2170;
  assign new_n2173 = n143 ^ n15;
  assign new_n2174 = n141 ^ n13;
  assign new_n2175 = new_n2174 ^ new_n2173;
  assign new_n2176 = n137 ^ n9;
  assign new_n2177 = n140 ^ n12;
  assign new_n2178 = new_n2177 ^ new_n2176;
  assign new_n2179 = new_n2178 ^ new_n2175;
  assign new_n2180 = new_n2179 ^ new_n2172;
  assign new_n2181 = n144 ^ n16;
  assign new_n2182 = new_n2181 ^ new_n2172;
  assign new_n2183 = ~new_n2173 & ~new_n2182;
  assign new_n2184 = new_n2183 ^ new_n2173;
  assign new_n2185 = new_n2176 ^ new_n2173;
  assign new_n2186 = n142 ^ n14;
  assign new_n2187 = new_n2186 ^ new_n2175;
  assign new_n2188 = new_n2187 ^ new_n2170;
  assign new_n2189 = new_n2185 & new_n2188;
  assign new_n2190 = new_n2189 ^ new_n2184;
  assign new_n2191 = new_n2186 ^ new_n2176;
  assign new_n2192 = new_n2191 ^ new_n2190;
  assign new_n2193 = new_n2177 ^ new_n2170;
  assign new_n2194 = new_n2193 ^ new_n2191;
  assign new_n2195 = new_n2186 ^ new_n2177;
  assign new_n2196 = new_n2194 & new_n2195;
  assign new_n2197 = new_n2187 ^ new_n2171;
  assign new_n2198 = new_n2178 & new_n2197;
  assign new_n2199 = new_n2198 ^ new_n2196;
  assign new_n2200 = new_n2174 ^ new_n2170;
  assign new_n2201 = new_n2200 ^ new_n2199;
  assign new_n2202 = new_n2201 ^ new_n2192;
  assign new_n2203 = new_n2177 ^ new_n2173;
  assign new_n2204 = new_n2203 ^ new_n2191;
  assign new_n2205 = new_n2179 & new_n2204;
  assign new_n2206 = new_n2205 ^ new_n2171;
  assign new_n2207 = new_n2206 ^ new_n2179;
  assign new_n2208 = new_n2181 ^ new_n2179;
  assign new_n2209 = new_n2182 ^ new_n2173;
  assign new_n2210 = new_n2209 ^ new_n2191;
  assign new_n2211 = new_n2208 & new_n2210;
  assign new_n2212 = new_n2211 ^ new_n2186;
  assign new_n2213 = new_n2212 ^ new_n2199;
  assign new_n2214 = new_n2213 ^ new_n2207;
  assign new_n2215 = ~new_n2202 & new_n2214;
  assign new_n2216 = ~new_n2172 & new_n2181;
  assign new_n2217 = ~new_n2181 & new_n2177;
  assign new_n2218 = new_n2217 ^ new_n2216;
  assign new_n2219 = new_n2218 ^ new_n2206;
  assign new_n2220 = new_n2219 ^ new_n2215;
  assign new_n2221 = new_n2180 & new_n2191;
  assign new_n2222 = new_n2221 ^ new_n2198;
  assign new_n2223 = new_n2222 ^ new_n2188;
  assign new_n2224 = new_n2223 ^ new_n2220;
  assign new_n2225 = new_n2221 ^ new_n2196;
  assign new_n2226 = new_n2182 ^ new_n2176;
  assign new_n2227 = new_n2197 ^ new_n2181;
  assign new_n2228 = new_n2226 & new_n2227;
  assign new_n2229 = new_n2228 ^ new_n2183;
  assign new_n2230 = new_n2229 ^ new_n2225;
  assign new_n2231 = ~new_n2230 & new_n2224;
  assign new_n2232 = new_n2231 ^ new_n2176;
  assign new_n2233 = new_n2218 ^ new_n2177;
  assign new_n2234 = new_n2233 ^ new_n2228;
  assign new_n2235 = new_n2173 ^ new_n2170;
  assign new_n2236 = new_n2211 ^ new_n2184;
  assign new_n2237 = new_n2176 ^ new_n2170;
  assign new_n2238 = new_n2233 ^ new_n2211;
  assign new_n2239 = new_n2238 ^ new_n2225;
  assign new_n2240 = new_n2239 ^ new_n2237;
  assign new_n2241 = new_n2228 ^ new_n2189;
  assign new_n2242 = new_n2241 ^ new_n2176;
  assign new_n2243 = new_n2242 ^ new_n2223;
  assign new_n2244 = new_n2243 ^ new_n2215;
  assign new_n2245 = new_n2240 & new_n2244;
  assign new_n2246 = new_n2245 ^ new_n2219;
  assign new_n2247 = new_n2246 ^ new_n2223;
  assign new_n2248 = new_n2231 ^ new_n2215;
  assign new_n2249 = ~new_n2248 & new_n2243;
  assign new_n2250 = new_n2249 ^ new_n2215;
  assign new_n2251 = new_n2247 & new_n2250;
  assign new_n2252 = new_n2249 ^ new_n2243;
  assign new_n2253 = new_n2252 ^ new_n2251;
  assign new_n2254 = new_n2253 ^ new_n2236;
  assign new_n2255 = new_n2254 ^ new_n2235;
  assign new_n2256 = new_n2255 ^ new_n2234;
  assign new_n2257 = new_n2256 ^ new_n2232;
  assign new_n2258 = ~new_n2257 & new_n2180;
  assign new_n2259 = new_n2251 ^ new_n2245;
  assign new_n2260 = new_n2259 ^ new_n2214;
  assign new_n2261 = new_n2185 & new_n2260;
  assign new_n2262 = new_n2261 ^ new_n2258;
  assign new_n2263 = new_n2251 ^ new_n2240;
  assign new_n2264 = new_n2182 & new_n2263;
  assign new_n2265 = new_n2255 ^ new_n2177;
  assign new_n2266 = new_n2245 ^ new_n2189;
  assign new_n2267 = new_n2266 ^ new_n2206;
  assign new_n2268 = new_n2267 ^ new_n2265;
  assign new_n2269 = ~new_n2268 & new_n2194;
  assign new_n2270 = new_n2269 ^ new_n2264;
  assign new_n2271 = new_n2209 & new_n2263;
  assign new_n2272 = new_n2227 & new_n2247;
  assign new_n2273 = new_n2272 ^ new_n2271;
  assign new_n2274 = ~new_n2268 & new_n2195;
  assign new_n2275 = new_n2245 ^ new_n2231;
  assign new_n2276 = new_n2242 ^ new_n2219;
  assign new_n2277 = new_n2276 ^ new_n2275;
  assign new_n2278 = new_n2178 & new_n2277;
  assign new_n2279 = new_n2278 ^ new_n2274;
  assign new_n2280 = new_n2279 ^ new_n2273;
  assign new_n2281 = new_n2280 ^ new_n2270;
  assign new_n2282 = new_n2281 ^ new_n2262;
  assign new_n2283 = n178 ^ n50;
  assign new_n2284 = n179 ^ n51;
  assign new_n2285 = new_n2284 ^ new_n2283;
  assign new_n2286 = n183 ^ n55;
  assign new_n2287 = n181 ^ n53;
  assign new_n2288 = new_n2287 ^ new_n2286;
  assign new_n2289 = n177 ^ n49;
  assign new_n2290 = n180 ^ n52;
  assign new_n2291 = new_n2290 ^ new_n2289;
  assign new_n2292 = new_n2291 ^ new_n2288;
  assign new_n2293 = new_n2292 ^ new_n2285;
  assign new_n2294 = n184 ^ n56;
  assign new_n2295 = new_n2294 ^ new_n2285;
  assign new_n2296 = ~new_n2286 & ~new_n2295;
  assign new_n2297 = new_n2296 ^ new_n2286;
  assign new_n2298 = n182 ^ n54;
  assign new_n2299 = new_n2298 ^ new_n2288;
  assign new_n2300 = new_n2299 ^ new_n2284;
  assign new_n2301 = new_n2289 ^ new_n2286;
  assign new_n2302 = new_n2300 & new_n2301;
  assign new_n2303 = new_n2302 ^ new_n2297;
  assign new_n2304 = new_n2298 ^ new_n2289;
  assign new_n2305 = new_n2304 ^ new_n2303;
  assign new_n2306 = new_n2298 ^ new_n2290;
  assign new_n2307 = new_n2290 ^ new_n2284;
  assign new_n2308 = new_n2307 ^ new_n2304;
  assign new_n2309 = new_n2306 & new_n2308;
  assign new_n2310 = new_n2299 ^ new_n2283;
  assign new_n2311 = new_n2291 & new_n2310;
  assign new_n2312 = new_n2311 ^ new_n2309;
  assign new_n2313 = new_n2287 ^ new_n2284;
  assign new_n2314 = new_n2313 ^ new_n2312;
  assign new_n2315 = new_n2314 ^ new_n2305;
  assign new_n2316 = new_n2290 ^ new_n2286;
  assign new_n2317 = new_n2316 ^ new_n2304;
  assign new_n2318 = new_n2292 & new_n2317;
  assign new_n2319 = new_n2318 ^ new_n2283;
  assign new_n2320 = new_n2319 ^ new_n2292;
  assign new_n2321 = new_n2294 ^ new_n2292;
  assign new_n2322 = new_n2295 ^ new_n2286;
  assign new_n2323 = new_n2322 ^ new_n2304;
  assign new_n2324 = new_n2321 & new_n2323;
  assign new_n2325 = new_n2324 ^ new_n2298;
  assign new_n2326 = new_n2325 ^ new_n2312;
  assign new_n2327 = new_n2326 ^ new_n2320;
  assign new_n2328 = ~new_n2315 & new_n2327;
  assign new_n2329 = ~new_n2285 & new_n2294;
  assign new_n2330 = ~new_n2294 & new_n2290;
  assign new_n2331 = new_n2330 ^ new_n2329;
  assign new_n2332 = new_n2331 ^ new_n2319;
  assign new_n2333 = new_n2332 ^ new_n2328;
  assign new_n2334 = new_n2293 & new_n2304;
  assign new_n2335 = new_n2334 ^ new_n2311;
  assign new_n2336 = new_n2335 ^ new_n2300;
  assign new_n2337 = new_n2336 ^ new_n2333;
  assign new_n2338 = new_n2295 ^ new_n2289;
  assign new_n2339 = new_n2310 ^ new_n2294;
  assign new_n2340 = new_n2338 & new_n2339;
  assign new_n2341 = new_n2340 ^ new_n2296;
  assign new_n2342 = new_n2334 ^ new_n2309;
  assign new_n2343 = new_n2342 ^ new_n2341;
  assign new_n2344 = ~new_n2343 & new_n2337;
  assign new_n2345 = new_n2344 ^ new_n2289;
  assign new_n2346 = new_n2331 ^ new_n2290;
  assign new_n2347 = new_n2346 ^ new_n2340;
  assign new_n2348 = new_n2286 ^ new_n2284;
  assign new_n2349 = new_n2324 ^ new_n2297;
  assign new_n2350 = new_n2289 ^ new_n2284;
  assign new_n2351 = new_n2346 ^ new_n2324;
  assign new_n2352 = new_n2351 ^ new_n2342;
  assign new_n2353 = new_n2352 ^ new_n2350;
  assign new_n2354 = new_n2340 ^ new_n2302;
  assign new_n2355 = new_n2354 ^ new_n2289;
  assign new_n2356 = new_n2355 ^ new_n2336;
  assign new_n2357 = new_n2356 ^ new_n2328;
  assign new_n2358 = new_n2353 & new_n2357;
  assign new_n2359 = new_n2358 ^ new_n2332;
  assign new_n2360 = new_n2359 ^ new_n2336;
  assign new_n2361 = new_n2344 ^ new_n2328;
  assign new_n2362 = ~new_n2361 & new_n2356;
  assign new_n2363 = new_n2362 ^ new_n2328;
  assign new_n2364 = new_n2360 & new_n2363;
  assign new_n2365 = new_n2362 ^ new_n2356;
  assign new_n2366 = new_n2365 ^ new_n2364;
  assign new_n2367 = new_n2366 ^ new_n2349;
  assign new_n2368 = new_n2367 ^ new_n2348;
  assign new_n2369 = new_n2368 ^ new_n2347;
  assign new_n2370 = new_n2369 ^ new_n2345;
  assign new_n2371 = ~new_n2370 & new_n2293;
  assign new_n2372 = new_n2364 ^ new_n2358;
  assign new_n2373 = new_n2372 ^ new_n2327;
  assign new_n2374 = new_n2301 & new_n2373;
  assign new_n2375 = new_n2374 ^ new_n2371;
  assign new_n2376 = new_n2364 ^ new_n2353;
  assign new_n2377 = new_n2295 & new_n2376;
  assign new_n2378 = new_n2368 ^ new_n2290;
  assign new_n2379 = new_n2358 ^ new_n2302;
  assign new_n2380 = new_n2379 ^ new_n2319;
  assign new_n2381 = new_n2380 ^ new_n2378;
  assign new_n2382 = ~new_n2381 & new_n2308;
  assign new_n2383 = new_n2382 ^ new_n2377;
  assign new_n2384 = new_n2339 & new_n2360;
  assign new_n2385 = new_n2322 & new_n2376;
  assign new_n2386 = new_n2385 ^ new_n2384;
  assign new_n2387 = ~new_n2381 & new_n2306;
  assign new_n2388 = new_n2358 ^ new_n2344;
  assign new_n2389 = new_n2355 ^ new_n2332;
  assign new_n2390 = new_n2389 ^ new_n2388;
  assign new_n2391 = new_n2291 & new_n2390;
  assign new_n2392 = new_n2391 ^ new_n2387;
  assign new_n2393 = new_n2392 ^ new_n2386;
  assign new_n2394 = new_n2393 ^ new_n2383;
  assign new_n2395 = new_n2394 ^ new_n2375;
  assign new_n2396 = new_n2395 ^ new_n2282;
  assign new_n2397 = n226 ^ n98;
  assign new_n2398 = n227 ^ n99;
  assign new_n2399 = new_n2398 ^ new_n2397;
  assign new_n2400 = n232 ^ n104;
  assign new_n2401 = new_n2400 ^ new_n2399;
  assign new_n2402 = n230 ^ n102;
  assign new_n2403 = n225 ^ n97;
  assign new_n2404 = new_n2403 ^ new_n2402;
  assign new_n2405 = n228 ^ n100;
  assign new_n2406 = new_n2405 ^ new_n2403;
  assign new_n2407 = n231 ^ n103;
  assign new_n2408 = n229 ^ n101;
  assign new_n2409 = new_n2408 ^ new_n2407;
  assign new_n2410 = new_n2409 ^ new_n2406;
  assign new_n2411 = new_n2410 ^ new_n2399;
  assign new_n2412 = new_n2404 & new_n2411;
  assign new_n2413 = new_n2409 ^ new_n2402;
  assign new_n2414 = new_n2413 ^ new_n2397;
  assign new_n2415 = new_n2406 & new_n2414;
  assign new_n2416 = new_n2415 ^ new_n2412;
  assign new_n2417 = new_n2413 ^ new_n2398;
  assign new_n2418 = new_n2417 ^ new_n2416;
  assign new_n2419 = new_n2403 ^ new_n2401;
  assign new_n2420 = new_n2414 ^ new_n2400;
  assign new_n2421 = new_n2419 & new_n2420;
  assign new_n2422 = new_n2407 ^ new_n2403;
  assign new_n2423 = new_n2417 & new_n2422;
  assign new_n2424 = new_n2423 ^ new_n2421;
  assign new_n2425 = new_n2424 ^ new_n2403;
  assign new_n2426 = new_n2425 ^ new_n2418;
  assign new_n2427 = new_n2405 ^ new_n2401;
  assign new_n2428 = new_n2400 & new_n2427;
  assign new_n2429 = new_n2428 ^ new_n2405;
  assign new_n2430 = new_n2407 ^ new_n2405;
  assign new_n2431 = new_n2430 ^ new_n2404;
  assign new_n2432 = new_n2410 & new_n2431;
  assign new_n2433 = new_n2432 ^ new_n2397;
  assign new_n2434 = new_n2433 ^ new_n2429;
  assign new_n2435 = ~new_n2401 & ~new_n2407;
  assign new_n2436 = new_n2435 ^ new_n2407;
  assign new_n2437 = new_n2436 ^ new_n2423;
  assign new_n2438 = new_n2437 ^ new_n2404;
  assign new_n2439 = new_n2405 ^ new_n2398;
  assign new_n2440 = new_n2439 ^ new_n2404;
  assign new_n2441 = new_n2405 ^ new_n2402;
  assign new_n2442 = new_n2440 & new_n2441;
  assign new_n2443 = new_n2442 ^ new_n2415;
  assign new_n2444 = new_n2408 ^ new_n2398;
  assign new_n2445 = new_n2444 ^ new_n2443;
  assign new_n2446 = new_n2445 ^ new_n2438;
  assign new_n2447 = new_n2433 ^ new_n2410;
  assign new_n2448 = new_n2410 ^ new_n2400;
  assign new_n2449 = new_n2407 ^ new_n2401;
  assign new_n2450 = new_n2449 ^ new_n2404;
  assign new_n2451 = new_n2448 & new_n2450;
  assign new_n2452 = new_n2451 ^ new_n2402;
  assign new_n2453 = new_n2452 ^ new_n2443;
  assign new_n2454 = new_n2453 ^ new_n2447;
  assign new_n2455 = ~new_n2446 & new_n2454;
  assign new_n2456 = new_n2455 ^ new_n2434;
  assign new_n2457 = new_n2456 ^ new_n2418;
  assign new_n2458 = new_n2442 ^ new_n2412;
  assign new_n2459 = new_n2435 ^ new_n2421;
  assign new_n2460 = new_n2459 ^ new_n2458;
  assign new_n2461 = ~new_n2460 & new_n2457;
  assign new_n2462 = new_n2461 ^ new_n2455;
  assign new_n2463 = ~new_n2426 & ~new_n2462;
  assign new_n2464 = new_n2463 ^ new_n2461;
  assign new_n2465 = new_n2455 ^ new_n2426;
  assign new_n2466 = new_n2403 ^ new_n2398;
  assign new_n2467 = new_n2451 ^ new_n2428;
  assign new_n2468 = new_n2467 ^ new_n2458;
  assign new_n2469 = new_n2468 ^ new_n2466;
  assign new_n2470 = new_n2465 & new_n2469;
  assign new_n2471 = new_n2470 ^ new_n2434;
  assign new_n2472 = new_n2471 ^ new_n2418;
  assign new_n2473 = ~new_n2464 & new_n2472;
  assign new_n2474 = new_n2473 ^ new_n2469;
  assign new_n2475 = new_n2401 & new_n2474;
  assign new_n2476 = new_n2407 ^ new_n2398;
  assign new_n2477 = new_n2451 ^ new_n2436;
  assign new_n2478 = new_n2465 ^ new_n2464;
  assign new_n2479 = new_n2478 ^ new_n2473;
  assign new_n2480 = new_n2479 ^ new_n2477;
  assign new_n2481 = new_n2480 ^ new_n2476;
  assign new_n2482 = new_n2481 ^ new_n2405;
  assign new_n2483 = new_n2470 ^ new_n2423;
  assign new_n2484 = new_n2483 ^ new_n2433;
  assign new_n2485 = new_n2484 ^ new_n2482;
  assign new_n2486 = new_n2441 & new_n2485;
  assign new_n2487 = new_n2470 ^ new_n2461;
  assign new_n2488 = new_n2434 ^ new_n2425;
  assign new_n2489 = new_n2488 ^ new_n2487;
  assign new_n2490 = new_n2406 & new_n2489;
  assign new_n2491 = new_n2490 ^ new_n2486;
  assign new_n2492 = new_n2478 ^ new_n2461;
  assign new_n2493 = new_n2492 ^ new_n2460;
  assign new_n2494 = new_n2450 & new_n2493;
  assign new_n2495 = new_n2494 ^ new_n2491;
  assign new_n2496 = new_n2495 ^ new_n2475;
  assign new_n2497 = new_n2473 ^ new_n2470;
  assign new_n2498 = new_n2497 ^ new_n2454;
  assign new_n2499 = new_n2417 & new_n2498;
  assign new_n2500 = new_n2499 ^ new_n2496;
  assign new_n2501 = new_n2440 & new_n2485;
  assign new_n2502 = new_n2501 ^ new_n2500;
  assign new_n2503 = new_n2414 & new_n2489;
  assign new_n2504 = new_n2478 ^ new_n2446;
  assign new_n2505 = new_n2431 & new_n2504;
  assign new_n2506 = new_n2505 ^ new_n2503;
  assign new_n2507 = new_n2506 ^ new_n2502;
  assign new_n2508 = n220 ^ n92;
  assign new_n2509 = n219 ^ n91;
  assign new_n2510 = new_n2509 ^ new_n2508;
  assign new_n2511 = n217 ^ n89;
  assign new_n2512 = n222 ^ n94;
  assign new_n2513 = new_n2512 ^ new_n2511;
  assign new_n2514 = new_n2513 ^ new_n2510;
  assign new_n2515 = n223 ^ n95;
  assign new_n2516 = new_n2515 ^ new_n2509;
  assign new_n2517 = new_n2511 ^ new_n2508;
  assign new_n2518 = n221 ^ n93;
  assign new_n2519 = new_n2518 ^ new_n2515;
  assign new_n2520 = new_n2519 ^ new_n2517;
  assign new_n2521 = n224 ^ n96;
  assign new_n2522 = new_n2521 ^ new_n2520;
  assign new_n2523 = n218 ^ n90;
  assign new_n2524 = new_n2523 ^ new_n2509;
  assign new_n2525 = new_n2524 ^ new_n2521;
  assign new_n2526 = new_n2525 ^ new_n2515;
  assign new_n2527 = new_n2526 ^ new_n2513;
  assign new_n2528 = new_n2522 & new_n2527;
  assign new_n2529 = ~new_n2515 & ~new_n2525;
  assign new_n2530 = new_n2529 ^ new_n2515;
  assign new_n2531 = new_n2530 ^ new_n2528;
  assign new_n2532 = new_n2519 ^ new_n2512;
  assign new_n2533 = new_n2532 ^ new_n2523;
  assign new_n2534 = new_n2517 & new_n2533;
  assign new_n2535 = new_n2524 ^ new_n2520;
  assign new_n2536 = new_n2513 & new_n2535;
  assign new_n2537 = new_n2536 ^ new_n2534;
  assign new_n2538 = new_n2532 ^ new_n2509;
  assign new_n2539 = new_n2538 ^ new_n2537;
  assign new_n2540 = new_n2515 ^ new_n2511;
  assign new_n2541 = new_n2538 & new_n2540;
  assign new_n2542 = new_n2525 ^ new_n2511;
  assign new_n2543 = new_n2533 ^ new_n2521;
  assign new_n2544 = new_n2542 & new_n2543;
  assign new_n2545 = new_n2544 ^ new_n2541;
  assign new_n2546 = new_n2545 ^ new_n2511;
  assign new_n2547 = new_n2546 ^ new_n2539;
  assign new_n2548 = new_n2525 ^ new_n2508;
  assign new_n2549 = new_n2521 & new_n2548;
  assign new_n2550 = new_n2549 ^ new_n2508;
  assign new_n2551 = new_n2515 ^ new_n2508;
  assign new_n2552 = new_n2551 ^ new_n2513;
  assign new_n2553 = new_n2520 & new_n2552;
  assign new_n2554 = new_n2553 ^ new_n2523;
  assign new_n2555 = new_n2554 ^ new_n2550;
  assign new_n2556 = new_n2541 ^ new_n2530;
  assign new_n2557 = new_n2556 ^ new_n2513;
  assign new_n2558 = new_n2512 ^ new_n2508;
  assign new_n2559 = new_n2514 & new_n2558;
  assign new_n2560 = new_n2559 ^ new_n2534;
  assign new_n2561 = new_n2518 ^ new_n2509;
  assign new_n2562 = new_n2561 ^ new_n2560;
  assign new_n2563 = new_n2562 ^ new_n2557;
  assign new_n2564 = new_n2554 ^ new_n2520;
  assign new_n2565 = new_n2528 ^ new_n2512;
  assign new_n2566 = new_n2565 ^ new_n2560;
  assign new_n2567 = new_n2566 ^ new_n2564;
  assign new_n2568 = ~new_n2563 & new_n2567;
  assign new_n2569 = new_n2568 ^ new_n2555;
  assign new_n2570 = new_n2569 ^ new_n2539;
  assign new_n2571 = new_n2559 ^ new_n2536;
  assign new_n2572 = new_n2544 ^ new_n2529;
  assign new_n2573 = new_n2572 ^ new_n2571;
  assign new_n2574 = ~new_n2573 & new_n2570;
  assign new_n2575 = new_n2574 ^ new_n2568;
  assign new_n2576 = ~new_n2547 & ~new_n2575;
  assign new_n2577 = new_n2576 ^ new_n2574;
  assign new_n2578 = new_n2568 ^ new_n2547;
  assign new_n2579 = new_n2511 ^ new_n2509;
  assign new_n2580 = new_n2549 ^ new_n2528;
  assign new_n2581 = new_n2580 ^ new_n2571;
  assign new_n2582 = new_n2581 ^ new_n2579;
  assign new_n2583 = new_n2578 & new_n2582;
  assign new_n2584 = new_n2583 ^ new_n2555;
  assign new_n2585 = new_n2584 ^ new_n2539;
  assign new_n2586 = ~new_n2577 & new_n2585;
  assign new_n2587 = new_n2578 ^ new_n2577;
  assign new_n2588 = new_n2587 ^ new_n2586;
  assign new_n2589 = new_n2588 ^ new_n2531;
  assign new_n2590 = new_n2589 ^ new_n2516;
  assign new_n2591 = new_n2590 ^ new_n2508;
  assign new_n2592 = new_n2583 ^ new_n2541;
  assign new_n2593 = new_n2592 ^ new_n2554;
  assign new_n2594 = new_n2593 ^ new_n2591;
  assign new_n2595 = new_n2514 & new_n2594;
  assign new_n2596 = new_n2586 ^ new_n2583;
  assign new_n2597 = new_n2596 ^ new_n2567;
  assign new_n2598 = new_n2538 & new_n2597;
  assign new_n2599 = new_n2558 & new_n2594;
  assign new_n2600 = new_n2583 ^ new_n2574;
  assign new_n2601 = new_n2555 ^ new_n2546;
  assign new_n2602 = new_n2601 ^ new_n2600;
  assign new_n2603 = new_n2517 & new_n2602;
  assign new_n2604 = new_n2603 ^ new_n2599;
  assign new_n2605 = new_n2587 ^ new_n2574;
  assign new_n2606 = new_n2605 ^ new_n2573;
  assign new_n2607 = new_n2527 & new_n2606;
  assign new_n2608 = new_n2607 ^ new_n2604;
  assign new_n2609 = new_n2586 ^ new_n2582;
  assign new_n2610 = new_n2525 & new_n2609;
  assign new_n2611 = new_n2610 ^ new_n2608;
  assign new_n2612 = new_n2611 ^ new_n2598;
  assign new_n2613 = new_n2612 ^ new_n2595;
  assign new_n2614 = new_n2587 ^ new_n2563;
  assign new_n2615 = new_n2552 & new_n2614;
  assign new_n2616 = new_n2533 & new_n2602;
  assign new_n2617 = new_n2616 ^ new_n2615;
  assign new_n2618 = new_n2617 ^ new_n2613;
  assign new_n2619 = new_n2618 ^ new_n2507;
  assign new_n2620 = new_n2449 & new_n2474;
  assign new_n2621 = new_n2420 & new_n2472;
  assign new_n2622 = new_n2621 ^ new_n2620;
  assign new_n2623 = new_n2622 ^ new_n2491;
  assign new_n2624 = new_n2422 & new_n2498;
  assign new_n2625 = new_n2461 ^ new_n2426;
  assign new_n2626 = new_n2400 & new_n2625;
  assign new_n2627 = new_n2410 & new_n2504;
  assign new_n2628 = new_n2627 ^ new_n2626;
  assign new_n2629 = new_n2628 ^ new_n2624;
  assign new_n2630 = new_n2629 ^ new_n2499;
  assign new_n2631 = new_n2630 ^ new_n2623;
  assign new_n2632 = new_n2631 ^ new_n2619;
  assign new_n2633 = new_n2632 ^ new_n2396;
  assign new_n2634 = new_n2574 ^ new_n2511;
  assign new_n2635 = new_n2549 ^ new_n2544;
  assign new_n2636 = new_n2635 ^ new_n2590;
  assign new_n2637 = new_n2636 ^ new_n2634;
  assign new_n2638 = new_n2535 & new_n2637;
  assign new_n2639 = new_n2540 & new_n2597;
  assign new_n2640 = new_n2639 ^ new_n2638;
  assign new_n2641 = new_n2610 ^ new_n2595;
  assign new_n2642 = new_n2526 & new_n2609;
  assign new_n2643 = new_n2543 & new_n2585;
  assign new_n2644 = new_n2643 ^ new_n2642;
  assign new_n2645 = new_n2644 ^ new_n2604;
  assign new_n2646 = new_n2645 ^ new_n2641;
  assign new_n2647 = new_n2646 ^ new_n2640;
  assign new_n2648 = new_n2647 ^ new_n391;
  assign new_n2649 = new_n2574 ^ new_n2547;
  assign new_n2650 = new_n2521 & new_n2649;
  assign new_n2651 = new_n2520 & new_n2614;
  assign new_n2652 = new_n2651 ^ new_n2650;
  assign new_n2653 = new_n2652 ^ new_n2639;
  assign new_n2654 = new_n2653 ^ new_n2598;
  assign new_n2655 = new_n2654 ^ new_n2645;
  assign new_n2656 = new_n2655 ^ new_n2648;
  assign new_n2657 = new_n2656 ^ new_n2633;
  assign new_n2658 = new_n2427 & new_n2625;
  assign new_n2659 = new_n2658 ^ new_n2502;
  assign new_n2660 = new_n2461 ^ new_n2403;
  assign new_n2661 = new_n2428 ^ new_n2421;
  assign new_n2662 = new_n2661 ^ new_n2481;
  assign new_n2663 = new_n2662 ^ new_n2660;
  assign new_n2664 = new_n2411 & new_n2663;
  assign new_n2665 = new_n2419 & new_n2472;
  assign new_n2666 = new_n2665 ^ new_n2664;
  assign new_n2667 = new_n2666 ^ new_n2629;
  assign new_n2668 = new_n2667 ^ new_n2659;
  assign new_n2669 = new_n2643 ^ new_n2615;
  assign new_n2670 = new_n2522 & new_n2606;
  assign new_n2671 = new_n2670 ^ new_n2650;
  assign new_n2672 = new_n2671 ^ new_n2611;
  assign new_n2673 = new_n2672 ^ new_n2669;
  assign new_n2674 = new_n2673 ^ new_n2668;
  assign new_n2675 = new_n2548 & new_n2649;
  assign new_n2676 = new_n2675 ^ new_n2613;
  assign new_n2677 = new_n2542 & new_n2585;
  assign new_n2678 = new_n2677 ^ new_n2638;
  assign new_n2679 = new_n2678 ^ new_n2653;
  assign new_n2680 = new_n2679 ^ new_n2676;
  assign new_n2681 = new_n2680 ^ new_n2674;
  assign new_n2682 = new_n2252 ^ new_n2202;
  assign new_n2683 = ~new_n2682 & new_n2204;
  assign new_n2684 = new_n2683 ^ new_n2272;
  assign new_n2685 = new_n2243 ^ new_n2231;
  assign new_n2686 = new_n2181 & new_n2685;
  assign new_n2687 = new_n2252 ^ new_n2231;
  assign new_n2688 = new_n2687 ^ new_n2230;
  assign new_n2689 = ~new_n2688 & new_n2208;
  assign new_n2690 = new_n2689 ^ new_n2686;
  assign new_n2691 = ~new_n2688 & new_n2210;
  assign new_n2692 = new_n2691 ^ new_n2279;
  assign new_n2693 = new_n2692 ^ new_n2264;
  assign new_n2694 = new_n2693 ^ new_n2690;
  assign new_n2695 = new_n2694 ^ new_n2684;
  assign new_n2696 = new_n2365 ^ new_n2315;
  assign new_n2697 = ~new_n2696 & new_n2317;
  assign new_n2698 = new_n2697 ^ new_n2384;
  assign new_n2699 = new_n2356 ^ new_n2344;
  assign new_n2700 = new_n2294 & new_n2699;
  assign new_n2701 = new_n2365 ^ new_n2344;
  assign new_n2702 = new_n2701 ^ new_n2343;
  assign new_n2703 = ~new_n2702 & new_n2321;
  assign new_n2704 = new_n2703 ^ new_n2700;
  assign new_n2705 = ~new_n2702 & new_n2323;
  assign new_n2706 = new_n2705 ^ new_n2392;
  assign new_n2707 = new_n2706 ^ new_n2377;
  assign new_n2708 = new_n2707 ^ new_n2704;
  assign new_n2709 = new_n2708 ^ new_n2698;
  assign new_n2710 = new_n2709 ^ new_n2695;
  assign new_n2711 = new_n2619 ^ new_n401;
  assign new_n2712 = new_n2711 ^ new_n2710;
  assign new_n2713 = new_n2712 ^ new_n2681;
  assign new_n2714 = new_n2713 ^ new_n2657;
  assign new_n2715 = new_n2188 & new_n2260;
  assign new_n2716 = new_n2715 ^ new_n2693;
  assign new_n2717 = ~new_n2682 & new_n2179;
  assign new_n2718 = new_n2717 ^ new_n2689;
  assign new_n2719 = new_n2718 ^ new_n2683;
  assign new_n2720 = new_n2719 ^ new_n2716;
  assign new_n2721 = new_n2300 & new_n2373;
  assign new_n2722 = new_n2721 ^ new_n2707;
  assign new_n2723 = ~new_n2696 & new_n2292;
  assign new_n2724 = new_n2723 ^ new_n2703;
  assign new_n2725 = new_n2724 ^ new_n2697;
  assign new_n2726 = new_n2725 ^ new_n2722;
  assign new_n2727 = new_n2726 ^ new_n2720;
  assign new_n2728 = new_n2727 ^ new_n372;
  assign new_n2729 = new_n2728 ^ new_n2619;
  assign new_n2730 = new_n2621 ^ new_n2505;
  assign new_n2731 = new_n2448 & new_n2493;
  assign new_n2732 = new_n2731 ^ new_n2626;
  assign new_n2733 = new_n2732 ^ new_n2496;
  assign new_n2734 = new_n2733 ^ new_n2730;
  assign new_n2735 = new_n2670 ^ new_n2651;
  assign new_n2736 = new_n2735 ^ new_n2615;
  assign new_n2737 = new_n2736 ^ new_n2612;
  assign new_n2738 = new_n2737 ^ new_n2734;
  assign new_n2739 = new_n2738 ^ new_n2673;
  assign new_n2740 = new_n2739 ^ new_n2729;
  assign new_n2741 = new_n2716 ^ new_n2269;
  assign new_n2742 = new_n2197 & new_n2277;
  assign new_n2743 = new_n2742 ^ new_n2683;
  assign new_n2744 = new_n2743 ^ new_n2741;
  assign new_n2745 = new_n2722 ^ new_n2382;
  assign new_n2746 = new_n2310 & new_n2390;
  assign new_n2747 = new_n2746 ^ new_n2697;
  assign new_n2748 = new_n2747 ^ new_n2745;
  assign new_n2749 = new_n2748 ^ new_n2744;
  assign new_n2750 = new_n2503 ^ new_n2501;
  assign new_n2751 = new_n2731 ^ new_n2627;
  assign new_n2752 = new_n2751 ^ new_n2505;
  assign new_n2753 = new_n2752 ^ new_n2495;
  assign new_n2754 = new_n2753 ^ new_n2750;
  assign new_n2755 = new_n2754 ^ new_n2749;
  assign new_n2756 = new_n2618 ^ new_n363;
  assign new_n2757 = new_n2616 ^ new_n2595;
  assign new_n2758 = new_n2736 ^ new_n2608;
  assign new_n2759 = new_n2758 ^ new_n2757;
  assign new_n2760 = new_n2759 ^ new_n2756;
  assign new_n2761 = new_n2760 ^ new_n2755;
  assign new_n2762 = new_n2761 ^ new_n2740;
  assign new_n2763 = new_n2762 ^ new_n2714;
  assign new_n2764 = new_n2182 ^ new_n2177;
  assign new_n2765 = new_n2685 & new_n2764;
  assign new_n2766 = new_n2765 ^ new_n2741;
  assign new_n2767 = new_n2226 & new_n2247;
  assign new_n2768 = new_n2767 ^ new_n2258;
  assign new_n2769 = new_n2717 ^ new_n2686;
  assign new_n2770 = new_n2769 ^ new_n2261;
  assign new_n2771 = new_n2770 ^ new_n2768;
  assign new_n2772 = new_n2771 ^ new_n2766;
  assign new_n2773 = new_n2295 ^ new_n2290;
  assign new_n2774 = new_n2699 & new_n2773;
  assign new_n2775 = new_n2774 ^ new_n2745;
  assign new_n2776 = new_n2338 & new_n2360;
  assign new_n2777 = new_n2776 ^ new_n2371;
  assign new_n2778 = new_n2723 ^ new_n2700;
  assign new_n2779 = new_n2778 ^ new_n2374;
  assign new_n2780 = new_n2779 ^ new_n2777;
  assign new_n2781 = new_n2780 ^ new_n2775;
  assign new_n2782 = new_n2781 ^ new_n2772;
  assign new_n2783 = new_n2664 ^ new_n2624;
  assign new_n2784 = new_n2501 ^ new_n2475;
  assign new_n2785 = new_n2784 ^ new_n2623;
  assign new_n2786 = new_n2785 ^ new_n2783;
  assign new_n2787 = new_n2786 ^ new_n2782;
  assign new_n2788 = new_n2680 ^ new_n423;
  assign new_n2789 = new_n2788 ^ new_n2647;
  assign new_n2790 = new_n2789 ^ new_n2787;
  assign new_n2791 = new_n2790 ^ new_n2714;
  assign new_n2792 = new_n2742 ^ new_n2269;
  assign new_n2793 = new_n2719 ^ new_n2692;
  assign new_n2794 = new_n2793 ^ new_n2792;
  assign new_n2795 = new_n2746 ^ new_n2382;
  assign new_n2796 = new_n2725 ^ new_n2706;
  assign new_n2797 = new_n2796 ^ new_n2795;
  assign new_n2798 = new_n2797 ^ new_n2794;
  assign new_n2799 = new_n2503 ^ new_n2490;
  assign new_n2800 = new_n2404 & new_n2663;
  assign new_n2801 = new_n2800 ^ new_n2667;
  assign new_n2802 = new_n2801 ^ new_n2799;
  assign new_n2803 = new_n2802 ^ new_n2798;
  assign new_n2804 = new_n2759 ^ new_n431;
  assign new_n2805 = new_n2616 ^ new_n2603;
  assign new_n2806 = new_n2513 & new_n2637;
  assign new_n2807 = new_n2806 ^ new_n2679;
  assign new_n2808 = new_n2807 ^ new_n2805;
  assign new_n2809 = new_n2808 ^ new_n2804;
  assign new_n2810 = new_n2809 ^ new_n2803;
  assign new_n2811 = new_n2810 ^ new_n2791;
  assign new_n2812 = new_n2762 & new_n2811;
  assign new_n2813 = new_n2790 ^ new_n2761;
  assign new_n2814 = new_n2742 ^ new_n2278;
  assign new_n2815 = ~new_n2257 & new_n2191;
  assign new_n2816 = new_n2815 ^ new_n2771;
  assign new_n2817 = new_n2816 ^ new_n2814;
  assign new_n2818 = new_n2746 ^ new_n2391;
  assign new_n2819 = ~new_n2370 & new_n2304;
  assign new_n2820 = new_n2819 ^ new_n2780;
  assign new_n2821 = new_n2820 ^ new_n2818;
  assign new_n2822 = new_n2821 ^ new_n2817;
  assign new_n2823 = new_n2822 ^ new_n2808;
  assign new_n2824 = new_n2752 ^ new_n2500;
  assign new_n2825 = new_n2824 ^ new_n2737;
  assign new_n2826 = new_n2825 ^ new_n442;
  assign new_n2827 = new_n2826 ^ new_n2823;
  assign new_n2828 = new_n2827 ^ new_n2810;
  assign new_n2829 = new_n2828 ^ new_n2763;
  assign new_n2830 = new_n2813 & new_n2829;
  assign new_n2831 = new_n2830 ^ new_n2812;
  assign new_n2832 = new_n2827 ^ new_n2791;
  assign new_n2833 = new_n2832 ^ new_n2831;
  assign new_n2834 = new_n2761 ^ new_n2657;
  assign new_n2835 = new_n2832 & new_n2834;
  assign new_n2836 = new_n2655 ^ new_n411;
  assign new_n2837 = new_n2779 ^ new_n2721;
  assign new_n2838 = new_n2837 ^ new_n2393;
  assign new_n2839 = new_n2770 ^ new_n2715;
  assign new_n2840 = new_n2839 ^ new_n2280;
  assign new_n2841 = new_n2840 ^ new_n2838;
  assign new_n2842 = new_n2841 ^ new_n2619;
  assign new_n2843 = new_n2842 ^ new_n2836;
  assign new_n2844 = new_n2843 ^ new_n2828;
  assign new_n2845 = new_n2844 ^ new_n2761;
  assign new_n2846 = new_n2843 ^ new_n2811;
  assign new_n2847 = new_n2845 & new_n2846;
  assign new_n2848 = new_n2847 ^ new_n2835;
  assign new_n2849 = new_n2848 ^ new_n2761;
  assign new_n2850 = new_n2849 ^ new_n2833;
  assign new_n2851 = new_n2844 ^ new_n2740;
  assign new_n2852 = new_n2843 & new_n2851;
  assign new_n2853 = new_n2852 ^ new_n2740;
  assign new_n2854 = new_n2790 ^ new_n2740;
  assign new_n2855 = new_n2854 ^ new_n2834;
  assign new_n2856 = new_n2763 & new_n2855;
  assign new_n2857 = new_n2856 ^ new_n2810;
  assign new_n2858 = new_n2857 ^ new_n2853;
  assign new_n2859 = ~new_n2657 & ~new_n2844;
  assign new_n2860 = new_n2859 ^ new_n2657;
  assign new_n2861 = new_n2860 ^ new_n2835;
  assign new_n2862 = new_n2861 ^ new_n2813;
  assign new_n2863 = new_n2827 ^ new_n2740;
  assign new_n2864 = new_n2863 ^ new_n2813;
  assign new_n2865 = new_n2854 & new_n2864;
  assign new_n2866 = new_n2865 ^ new_n2812;
  assign new_n2867 = new_n2827 ^ new_n2713;
  assign new_n2868 = new_n2867 ^ new_n2866;
  assign new_n2869 = new_n2868 ^ new_n2862;
  assign new_n2870 = new_n2857 ^ new_n2763;
  assign new_n2871 = new_n2843 ^ new_n2763;
  assign new_n2872 = new_n2844 ^ new_n2657;
  assign new_n2873 = new_n2872 ^ new_n2813;
  assign new_n2874 = new_n2871 & new_n2873;
  assign new_n2875 = new_n2874 ^ new_n2866;
  assign new_n2876 = new_n2875 ^ new_n2790;
  assign new_n2877 = new_n2876 ^ new_n2870;
  assign new_n2878 = ~new_n2869 & new_n2877;
  assign new_n2879 = new_n2878 ^ new_n2858;
  assign new_n2880 = new_n2879 ^ new_n2833;
  assign new_n2881 = new_n2859 ^ new_n2847;
  assign new_n2882 = new_n2865 ^ new_n2830;
  assign new_n2883 = new_n2882 ^ new_n2881;
  assign new_n2884 = ~new_n2883 & new_n2880;
  assign new_n2885 = new_n2884 ^ new_n2878;
  assign new_n2886 = new_n2850 & new_n2885;
  assign new_n2887 = new_n2886 ^ new_n2869;
  assign new_n2888 = ~new_n2887 & new_n2763;
  assign new_n2889 = new_n2886 ^ new_n2884;
  assign new_n2890 = new_n2889 ^ new_n2883;
  assign new_n2891 = ~new_n2890 & new_n2871;
  assign new_n2892 = new_n2891 ^ new_n2888;
  assign new_n2893 = ~new_n2887 & new_n2855;
  assign new_n2894 = new_n2893 ^ new_n2892;
  assign new_n2895 = new_n2827 ^ new_n2761;
  assign new_n2896 = new_n2874 ^ new_n2852;
  assign new_n2897 = new_n2896 ^ new_n2882;
  assign new_n2898 = new_n2897 ^ new_n2895;
  assign new_n2899 = new_n2878 ^ new_n2850;
  assign new_n2900 = new_n2898 & new_n2899;
  assign new_n2901 = new_n2900 ^ new_n2858;
  assign new_n2902 = new_n2901 ^ new_n2833;
  assign new_n2903 = new_n2899 ^ new_n2886;
  assign new_n2904 = new_n2902 & new_n2903;
  assign new_n2905 = new_n2904 ^ new_n2900;
  assign new_n2906 = new_n2905 ^ new_n2877;
  assign new_n2907 = new_n2832 & new_n2906;
  assign new_n2908 = ~new_n2890 & new_n2873;
  assign new_n2909 = new_n2900 ^ new_n2884;
  assign new_n2910 = new_n2858 ^ new_n2849;
  assign new_n2911 = new_n2910 ^ new_n2909;
  assign new_n2912 = new_n2762 & new_n2911;
  assign new_n2913 = new_n2827 ^ new_n2657;
  assign new_n2914 = new_n2874 ^ new_n2860;
  assign new_n2915 = new_n2904 ^ new_n2886;
  assign new_n2916 = new_n2915 ^ new_n2914;
  assign new_n2917 = new_n2916 ^ new_n2913;
  assign new_n2918 = new_n2917 ^ new_n2740;
  assign new_n2919 = new_n2900 ^ new_n2835;
  assign new_n2920 = new_n2919 ^ new_n2857;
  assign new_n2921 = new_n2920 ^ new_n2918;
  assign new_n2922 = ~new_n2921 & new_n2854;
  assign new_n2923 = new_n2922 ^ new_n2912;
  assign new_n2924 = new_n2923 ^ new_n2908;
  assign new_n2925 = new_n2904 ^ new_n2898;
  assign new_n2926 = new_n2844 & new_n2925;
  assign new_n2927 = new_n2926 ^ new_n2924;
  assign new_n2928 = new_n2927 ^ new_n2907;
  assign new_n2929 = new_n2928 ^ new_n2894;
  assign new_n2930 = new_n2929 ^ new_n2169;
  assign new_n2931 = new_n2930 ^ new_n1403;
  assign new_n2932 = n239 ^ n111;
  assign new_n2933 = n233 ^ n105;
  assign new_n2934 = new_n2933 ^ new_n2932;
  assign new_n2935 = n235 ^ n107;
  assign new_n2936 = new_n2935 ^ new_n2933;
  assign new_n2937 = n236 ^ n108;
  assign new_n2938 = new_n2937 ^ new_n2933;
  assign new_n2939 = n237 ^ n109;
  assign new_n2940 = new_n2939 ^ new_n2932;
  assign new_n2941 = new_n2940 ^ new_n2938;
  assign new_n2942 = n240 ^ n112;
  assign new_n2943 = new_n2942 ^ new_n2941;
  assign new_n2944 = n234 ^ n106;
  assign new_n2945 = new_n2944 ^ new_n2935;
  assign new_n2946 = new_n2945 ^ new_n2942;
  assign new_n2947 = new_n2946 ^ new_n2932;
  assign new_n2948 = n238 ^ n110;
  assign new_n2949 = new_n2948 ^ new_n2933;
  assign new_n2950 = new_n2949 ^ new_n2947;
  assign new_n2951 = new_n2943 & new_n2950;
  assign new_n2952 = new_n2946 ^ new_n2937;
  assign new_n2953 = new_n2942 & new_n2952;
  assign new_n2954 = new_n2953 ^ new_n2951;
  assign new_n2955 = new_n2937 ^ new_n2935;
  assign new_n2956 = new_n2955 ^ new_n2949;
  assign new_n2957 = new_n2948 ^ new_n2937;
  assign new_n2958 = new_n2956 & new_n2957;
  assign new_n2959 = new_n2945 ^ new_n2941;
  assign new_n2960 = new_n2949 & new_n2959;
  assign new_n2961 = new_n2960 ^ new_n2958;
  assign new_n2962 = new_n2961 ^ new_n2954;
  assign new_n2963 = new_n2962 ^ new_n2936;
  assign new_n2964 = ~new_n2932 & ~new_n2946;
  assign new_n2965 = new_n2964 ^ new_n2932;
  assign new_n2966 = new_n2948 ^ new_n2940;
  assign new_n2967 = new_n2966 ^ new_n2935;
  assign new_n2968 = new_n2934 & new_n2967;
  assign new_n2969 = new_n2968 ^ new_n2965;
  assign new_n2970 = new_n2969 ^ new_n2949;
  assign new_n2971 = new_n2966 ^ new_n2944;
  assign new_n2972 = new_n2938 & new_n2971;
  assign new_n2973 = new_n2972 ^ new_n2958;
  assign new_n2974 = new_n2939 ^ new_n2935;
  assign new_n2975 = new_n2974 ^ new_n2973;
  assign new_n2976 = new_n2975 ^ new_n2970;
  assign new_n2977 = new_n2937 ^ new_n2932;
  assign new_n2978 = new_n2977 ^ new_n2949;
  assign new_n2979 = new_n2941 & new_n2978;
  assign new_n2980 = new_n2979 ^ new_n2944;
  assign new_n2981 = new_n2980 ^ new_n2941;
  assign new_n2982 = new_n2951 ^ new_n2948;
  assign new_n2983 = new_n2982 ^ new_n2973;
  assign new_n2984 = new_n2983 ^ new_n2981;
  assign new_n2985 = ~new_n2976 & new_n2984;
  assign new_n2986 = new_n2972 ^ new_n2960;
  assign new_n2987 = new_n2986 ^ new_n2967;
  assign new_n2988 = new_n2971 ^ new_n2942;
  assign new_n2989 = new_n2946 ^ new_n2933;
  assign new_n2990 = new_n2988 & new_n2989;
  assign new_n2991 = new_n2990 ^ new_n2968;
  assign new_n2992 = new_n2991 ^ new_n2933;
  assign new_n2993 = new_n2992 ^ new_n2987;
  assign new_n2994 = new_n2993 ^ new_n2985;
  assign new_n2995 = new_n2963 & new_n2994;
  assign new_n2996 = new_n2953 ^ new_n2937;
  assign new_n2997 = new_n2996 ^ new_n2980;
  assign new_n2998 = new_n2997 ^ new_n2995;
  assign new_n2999 = new_n2998 ^ new_n2987;
  assign new_n3000 = new_n2997 ^ new_n2985;
  assign new_n3001 = new_n3000 ^ new_n2987;
  assign new_n3002 = new_n2990 ^ new_n2964;
  assign new_n3003 = new_n3002 ^ new_n2961;
  assign new_n3004 = ~new_n3003 & new_n3001;
  assign new_n3005 = new_n3004 ^ new_n2985;
  assign new_n3006 = new_n2993 & new_n3005;
  assign new_n3007 = new_n3006 ^ new_n2994;
  assign new_n3008 = new_n2999 & new_n3007;
  assign new_n3009 = new_n3008 ^ new_n2995;
  assign new_n3010 = new_n3009 ^ new_n2984;
  assign new_n3011 = new_n2934 & new_n3010;
  assign new_n3012 = new_n3004 ^ new_n2933;
  assign new_n3013 = new_n2935 ^ new_n2932;
  assign new_n3014 = new_n2965 ^ new_n2951;
  assign new_n3015 = new_n3008 ^ new_n3006;
  assign new_n3016 = new_n3015 ^ new_n3014;
  assign new_n3017 = new_n3016 ^ new_n3013;
  assign new_n3018 = new_n2990 ^ new_n2953;
  assign new_n3019 = new_n3018 ^ new_n3017;
  assign new_n3020 = new_n3019 ^ new_n3012;
  assign new_n3021 = ~new_n3020 & new_n2959;
  assign new_n3022 = new_n3021 ^ new_n3011;
  assign new_n3023 = new_n3008 ^ new_n2963;
  assign new_n3024 = new_n2946 & new_n3023;
  assign new_n3025 = new_n3017 ^ new_n2937;
  assign new_n3026 = new_n2995 ^ new_n2968;
  assign new_n3027 = new_n3026 ^ new_n2980;
  assign new_n3028 = new_n3027 ^ new_n3025;
  assign new_n3029 = ~new_n3028 & new_n2956;
  assign new_n3030 = new_n3029 ^ new_n3024;
  assign new_n3031 = new_n2988 & new_n2999;
  assign new_n3032 = new_n2947 & new_n3023;
  assign new_n3033 = new_n3032 ^ new_n3031;
  assign new_n3034 = ~new_n3028 & new_n2957;
  assign new_n3035 = new_n3004 ^ new_n2995;
  assign new_n3036 = new_n2997 ^ new_n2992;
  assign new_n3037 = new_n3036 ^ new_n3035;
  assign new_n3038 = new_n2938 & new_n3037;
  assign new_n3039 = new_n3038 ^ new_n3034;
  assign new_n3040 = new_n3039 ^ new_n3033;
  assign new_n3041 = new_n3040 ^ new_n3030;
  assign new_n3042 = new_n3041 ^ new_n3022;
  assign new_n3043 = n199 ^ n71;
  assign new_n3044 = n193 ^ n65;
  assign new_n3045 = new_n3044 ^ new_n3043;
  assign new_n3046 = n195 ^ n67;
  assign new_n3047 = new_n3046 ^ new_n3044;
  assign new_n3048 = n200 ^ n72;
  assign new_n3049 = n197 ^ n69;
  assign new_n3050 = new_n3049 ^ new_n3043;
  assign new_n3051 = n196 ^ n68;
  assign new_n3052 = new_n3051 ^ new_n3044;
  assign new_n3053 = new_n3052 ^ new_n3050;
  assign new_n3054 = new_n3053 ^ new_n3048;
  assign new_n3055 = n194 ^ n66;
  assign new_n3056 = new_n3055 ^ new_n3046;
  assign new_n3057 = new_n3056 ^ new_n3048;
  assign new_n3058 = new_n3057 ^ new_n3043;
  assign new_n3059 = n198 ^ n70;
  assign new_n3060 = new_n3059 ^ new_n3044;
  assign new_n3061 = new_n3060 ^ new_n3058;
  assign new_n3062 = new_n3054 & new_n3061;
  assign new_n3063 = new_n3057 ^ new_n3051;
  assign new_n3064 = new_n3048 & new_n3063;
  assign new_n3065 = new_n3064 ^ new_n3062;
  assign new_n3066 = new_n3051 ^ new_n3046;
  assign new_n3067 = new_n3066 ^ new_n3060;
  assign new_n3068 = new_n3059 ^ new_n3051;
  assign new_n3069 = new_n3067 & new_n3068;
  assign new_n3070 = new_n3056 ^ new_n3053;
  assign new_n3071 = new_n3060 & new_n3070;
  assign new_n3072 = new_n3071 ^ new_n3069;
  assign new_n3073 = new_n3072 ^ new_n3065;
  assign new_n3074 = new_n3073 ^ new_n3047;
  assign new_n3075 = ~new_n3043 & ~new_n3057;
  assign new_n3076 = new_n3075 ^ new_n3043;
  assign new_n3077 = new_n3059 ^ new_n3050;
  assign new_n3078 = new_n3077 ^ new_n3046;
  assign new_n3079 = new_n3045 & new_n3078;
  assign new_n3080 = new_n3079 ^ new_n3076;
  assign new_n3081 = new_n3080 ^ new_n3060;
  assign new_n3082 = new_n3077 ^ new_n3055;
  assign new_n3083 = new_n3052 & new_n3082;
  assign new_n3084 = new_n3083 ^ new_n3069;
  assign new_n3085 = new_n3049 ^ new_n3046;
  assign new_n3086 = new_n3085 ^ new_n3084;
  assign new_n3087 = new_n3086 ^ new_n3081;
  assign new_n3088 = new_n3051 ^ new_n3043;
  assign new_n3089 = new_n3088 ^ new_n3060;
  assign new_n3090 = new_n3053 & new_n3089;
  assign new_n3091 = new_n3090 ^ new_n3055;
  assign new_n3092 = new_n3091 ^ new_n3053;
  assign new_n3093 = new_n3062 ^ new_n3059;
  assign new_n3094 = new_n3093 ^ new_n3084;
  assign new_n3095 = new_n3094 ^ new_n3092;
  assign new_n3096 = ~new_n3087 & new_n3095;
  assign new_n3097 = new_n3083 ^ new_n3071;
  assign new_n3098 = new_n3097 ^ new_n3078;
  assign new_n3099 = new_n3082 ^ new_n3048;
  assign new_n3100 = new_n3057 ^ new_n3044;
  assign new_n3101 = new_n3099 & new_n3100;
  assign new_n3102 = new_n3101 ^ new_n3079;
  assign new_n3103 = new_n3102 ^ new_n3044;
  assign new_n3104 = new_n3103 ^ new_n3098;
  assign new_n3105 = new_n3104 ^ new_n3096;
  assign new_n3106 = new_n3074 & new_n3105;
  assign new_n3107 = new_n3064 ^ new_n3051;
  assign new_n3108 = new_n3107 ^ new_n3091;
  assign new_n3109 = new_n3108 ^ new_n3106;
  assign new_n3110 = new_n3109 ^ new_n3098;
  assign new_n3111 = new_n3108 ^ new_n3096;
  assign new_n3112 = new_n3111 ^ new_n3098;
  assign new_n3113 = new_n3101 ^ new_n3075;
  assign new_n3114 = new_n3113 ^ new_n3072;
  assign new_n3115 = ~new_n3114 & new_n3112;
  assign new_n3116 = new_n3115 ^ new_n3096;
  assign new_n3117 = new_n3104 & new_n3116;
  assign new_n3118 = new_n3117 ^ new_n3105;
  assign new_n3119 = new_n3110 & new_n3118;
  assign new_n3120 = new_n3119 ^ new_n3106;
  assign new_n3121 = new_n3120 ^ new_n3095;
  assign new_n3122 = new_n3045 & new_n3121;
  assign new_n3123 = new_n3115 ^ new_n3044;
  assign new_n3124 = new_n3101 ^ new_n3064;
  assign new_n3125 = new_n3046 ^ new_n3043;
  assign new_n3126 = new_n3076 ^ new_n3062;
  assign new_n3127 = new_n3119 ^ new_n3117;
  assign new_n3128 = new_n3127 ^ new_n3126;
  assign new_n3129 = new_n3128 ^ new_n3125;
  assign new_n3130 = new_n3129 ^ new_n3124;
  assign new_n3131 = new_n3130 ^ new_n3123;
  assign new_n3132 = ~new_n3131 & new_n3070;
  assign new_n3133 = new_n3132 ^ new_n3122;
  assign new_n3134 = new_n3119 ^ new_n3074;
  assign new_n3135 = new_n3057 & new_n3134;
  assign new_n3136 = new_n3129 ^ new_n3051;
  assign new_n3137 = new_n3106 ^ new_n3079;
  assign new_n3138 = new_n3137 ^ new_n3091;
  assign new_n3139 = new_n3138 ^ new_n3136;
  assign new_n3140 = ~new_n3139 & new_n3067;
  assign new_n3141 = new_n3140 ^ new_n3135;
  assign new_n3142 = new_n3099 & new_n3110;
  assign new_n3143 = new_n3058 & new_n3134;
  assign new_n3144 = new_n3143 ^ new_n3142;
  assign new_n3145 = ~new_n3139 & new_n3068;
  assign new_n3146 = new_n3115 ^ new_n3106;
  assign new_n3147 = new_n3108 ^ new_n3103;
  assign new_n3148 = new_n3147 ^ new_n3146;
  assign new_n3149 = new_n3052 & new_n3148;
  assign new_n3150 = new_n3149 ^ new_n3145;
  assign new_n3151 = new_n3150 ^ new_n3144;
  assign new_n3152 = new_n3151 ^ new_n3141;
  assign new_n3153 = new_n3152 ^ new_n3133;
  assign new_n3154 = new_n3153 ^ new_n3042;
  assign new_n3155 = n151 ^ n23;
  assign new_n3156 = n149 ^ n21;
  assign new_n3157 = new_n3156 ^ new_n3155;
  assign new_n3158 = n150 ^ n22;
  assign new_n3159 = new_n3158 ^ new_n3157;
  assign new_n3160 = n147 ^ n19;
  assign new_n3161 = new_n3160 ^ new_n3159;
  assign new_n3162 = n146 ^ n18;
  assign new_n3163 = new_n3162 ^ new_n3159;
  assign new_n3164 = n148 ^ n20;
  assign new_n3165 = n145 ^ n17;
  assign new_n3166 = new_n3165 ^ new_n3164;
  assign new_n3167 = new_n3163 & new_n3166;
  assign new_n3168 = new_n3165 ^ new_n3158;
  assign new_n3169 = new_n3166 ^ new_n3157;
  assign new_n3170 = new_n3162 ^ new_n3160;
  assign new_n3171 = new_n3170 ^ new_n3169;
  assign new_n3172 = new_n3168 & new_n3171;
  assign new_n3173 = new_n3172 ^ new_n3167;
  assign new_n3174 = new_n3173 ^ new_n3161;
  assign new_n3175 = new_n3165 ^ new_n3155;
  assign new_n3176 = new_n3161 & new_n3175;
  assign new_n3177 = n152 ^ n24;
  assign new_n3178 = new_n3177 ^ new_n3170;
  assign new_n3179 = new_n3178 ^ new_n3165;
  assign new_n3180 = new_n3177 ^ new_n3163;
  assign new_n3181 = new_n3179 & new_n3180;
  assign new_n3182 = new_n3181 ^ new_n3176;
  assign new_n3183 = new_n3182 ^ new_n3165;
  assign new_n3184 = new_n3183 ^ new_n3174;
  assign new_n3185 = new_n3164 ^ new_n3155;
  assign new_n3186 = new_n3185 ^ new_n3168;
  assign new_n3187 = new_n3169 & new_n3186;
  assign new_n3188 = new_n3187 ^ new_n3162;
  assign new_n3189 = ~new_n3170 & new_n3177;
  assign new_n3190 = ~new_n3177 & new_n3164;
  assign new_n3191 = new_n3190 ^ new_n3189;
  assign new_n3192 = new_n3191 ^ new_n3188;
  assign new_n3193 = ~new_n3155 & ~new_n3178;
  assign new_n3194 = new_n3193 ^ new_n3155;
  assign new_n3195 = new_n3194 ^ new_n3176;
  assign new_n3196 = new_n3195 ^ new_n3168;
  assign new_n3197 = new_n3164 ^ new_n3160;
  assign new_n3198 = new_n3197 ^ new_n3168;
  assign new_n3199 = new_n3164 ^ new_n3158;
  assign new_n3200 = new_n3198 & new_n3199;
  assign new_n3201 = new_n3200 ^ new_n3167;
  assign new_n3202 = new_n3160 ^ new_n3156;
  assign new_n3203 = new_n3202 ^ new_n3201;
  assign new_n3204 = new_n3203 ^ new_n3196;
  assign new_n3205 = new_n3188 ^ new_n3169;
  assign new_n3206 = new_n3177 ^ new_n3169;
  assign new_n3207 = new_n3178 ^ new_n3155;
  assign new_n3208 = new_n3207 ^ new_n3168;
  assign new_n3209 = new_n3206 & new_n3208;
  assign new_n3210 = new_n3209 ^ new_n3158;
  assign new_n3211 = new_n3210 ^ new_n3201;
  assign new_n3212 = new_n3211 ^ new_n3205;
  assign new_n3213 = ~new_n3204 & new_n3212;
  assign new_n3214 = new_n3213 ^ new_n3192;
  assign new_n3215 = new_n3214 ^ new_n3174;
  assign new_n3216 = new_n3193 ^ new_n3181;
  assign new_n3217 = new_n3200 ^ new_n3172;
  assign new_n3218 = new_n3217 ^ new_n3216;
  assign new_n3219 = ~new_n3218 & new_n3215;
  assign new_n3220 = new_n3219 ^ new_n3213;
  assign new_n3221 = ~new_n3184 & ~new_n3220;
  assign new_n3222 = new_n3221 ^ new_n3219;
  assign new_n3223 = new_n3213 ^ new_n3184;
  assign new_n3224 = new_n3165 ^ new_n3160;
  assign new_n3225 = new_n3191 ^ new_n3164;
  assign new_n3226 = new_n3225 ^ new_n3209;
  assign new_n3227 = new_n3226 ^ new_n3217;
  assign new_n3228 = new_n3227 ^ new_n3224;
  assign new_n3229 = new_n3223 & new_n3228;
  assign new_n3230 = new_n3229 ^ new_n3192;
  assign new_n3231 = new_n3230 ^ new_n3174;
  assign new_n3232 = ~new_n3222 & new_n3231;
  assign new_n3233 = new_n3232 ^ new_n3229;
  assign new_n3234 = new_n3233 ^ new_n3212;
  assign new_n3235 = new_n3161 & new_n3234;
  assign new_n3236 = new_n3175 & new_n3234;
  assign new_n3237 = new_n3219 ^ new_n3184;
  assign new_n3238 = new_n3177 & new_n3237;
  assign new_n3239 = new_n3223 ^ new_n3222;
  assign new_n3240 = new_n3239 ^ new_n3204;
  assign new_n3241 = new_n3169 & new_n3240;
  assign new_n3242 = new_n3241 ^ new_n3238;
  assign new_n3243 = new_n3242 ^ new_n3236;
  assign new_n3244 = new_n3243 ^ new_n3235;
  assign new_n3245 = new_n3232 ^ new_n3228;
  assign new_n3246 = new_n3207 & new_n3245;
  assign new_n3247 = new_n3180 & new_n3231;
  assign new_n3248 = new_n3247 ^ new_n3246;
  assign new_n3249 = new_n3160 ^ new_n3155;
  assign new_n3250 = new_n3209 ^ new_n3194;
  assign new_n3251 = new_n3239 ^ new_n3232;
  assign new_n3252 = new_n3251 ^ new_n3250;
  assign new_n3253 = new_n3252 ^ new_n3249;
  assign new_n3254 = new_n3253 ^ new_n3164;
  assign new_n3255 = new_n3229 ^ new_n3176;
  assign new_n3256 = new_n3255 ^ new_n3188;
  assign new_n3257 = new_n3256 ^ new_n3254;
  assign new_n3258 = new_n3199 & new_n3257;
  assign new_n3259 = new_n3229 ^ new_n3219;
  assign new_n3260 = new_n3192 ^ new_n3183;
  assign new_n3261 = new_n3260 ^ new_n3259;
  assign new_n3262 = new_n3166 & new_n3261;
  assign new_n3263 = new_n3262 ^ new_n3258;
  assign new_n3264 = new_n3263 ^ new_n3248;
  assign new_n3265 = new_n3264 ^ new_n3244;
  assign new_n3266 = new_n3265 ^ new_n3154;
  assign new_n3267 = n190 ^ n62;
  assign new_n3268 = n191 ^ n63;
  assign new_n3269 = n189 ^ n61;
  assign new_n3270 = new_n3269 ^ new_n3268;
  assign new_n3271 = new_n3270 ^ new_n3267;
  assign new_n3272 = n186 ^ n58;
  assign new_n3273 = new_n3272 ^ new_n3271;
  assign new_n3274 = n187 ^ n59;
  assign new_n3275 = new_n3274 ^ new_n3272;
  assign new_n3276 = n192 ^ n64;
  assign new_n3277 = new_n3276 ^ new_n3275;
  assign new_n3278 = ~new_n3268 & ~new_n3277;
  assign new_n3279 = new_n3278 ^ new_n3268;
  assign new_n3280 = new_n3274 ^ new_n3271;
  assign new_n3281 = n185 ^ n57;
  assign new_n3282 = new_n3281 ^ new_n3268;
  assign new_n3283 = new_n3280 & new_n3282;
  assign new_n3284 = new_n3283 ^ new_n3279;
  assign new_n3285 = new_n3281 ^ new_n3267;
  assign new_n3286 = new_n3285 ^ new_n3284;
  assign new_n3287 = n188 ^ n60;
  assign new_n3288 = new_n3287 ^ new_n3274;
  assign new_n3289 = new_n3288 ^ new_n3285;
  assign new_n3290 = new_n3287 ^ new_n3267;
  assign new_n3291 = new_n3289 & new_n3290;
  assign new_n3292 = new_n3287 ^ new_n3281;
  assign new_n3293 = new_n3273 & new_n3292;
  assign new_n3294 = new_n3293 ^ new_n3291;
  assign new_n3295 = new_n3274 ^ new_n3269;
  assign new_n3296 = new_n3295 ^ new_n3294;
  assign new_n3297 = new_n3296 ^ new_n3286;
  assign new_n3298 = new_n3292 ^ new_n3270;
  assign new_n3299 = new_n3287 ^ new_n3268;
  assign new_n3300 = new_n3299 ^ new_n3285;
  assign new_n3301 = new_n3298 & new_n3300;
  assign new_n3302 = new_n3301 ^ new_n3272;
  assign new_n3303 = new_n3302 ^ new_n3298;
  assign new_n3304 = new_n3298 ^ new_n3276;
  assign new_n3305 = new_n3277 ^ new_n3268;
  assign new_n3306 = new_n3305 ^ new_n3285;
  assign new_n3307 = new_n3304 & new_n3306;
  assign new_n3308 = new_n3307 ^ new_n3267;
  assign new_n3309 = new_n3308 ^ new_n3294;
  assign new_n3310 = new_n3309 ^ new_n3303;
  assign new_n3311 = ~new_n3297 & new_n3310;
  assign new_n3312 = new_n3298 ^ new_n3275;
  assign new_n3313 = new_n3285 & new_n3312;
  assign new_n3314 = new_n3313 ^ new_n3293;
  assign new_n3315 = new_n3314 ^ new_n3280;
  assign new_n3316 = new_n3281 ^ new_n3277;
  assign new_n3317 = new_n3276 ^ new_n3273;
  assign new_n3318 = new_n3316 & new_n3317;
  assign new_n3319 = new_n3318 ^ new_n3283;
  assign new_n3320 = new_n3319 ^ new_n3281;
  assign new_n3321 = new_n3320 ^ new_n3315;
  assign new_n3322 = new_n3321 ^ new_n3311;
  assign new_n3323 = new_n3281 ^ new_n3274;
  assign new_n3324 = new_n3287 ^ new_n3277;
  assign new_n3325 = new_n3276 & new_n3324;
  assign new_n3326 = new_n3325 ^ new_n3307;
  assign new_n3327 = new_n3313 ^ new_n3291;
  assign new_n3328 = new_n3327 ^ new_n3326;
  assign new_n3329 = new_n3328 ^ new_n3323;
  assign new_n3330 = new_n3322 & new_n3329;
  assign new_n3331 = new_n3325 ^ new_n3287;
  assign new_n3332 = new_n3331 ^ new_n3302;
  assign new_n3333 = new_n3332 ^ new_n3311;
  assign new_n3334 = new_n3333 ^ new_n3315;
  assign new_n3335 = new_n3318 ^ new_n3278;
  assign new_n3336 = new_n3335 ^ new_n3327;
  assign new_n3337 = ~new_n3336 & new_n3334;
  assign new_n3338 = new_n3337 ^ new_n3330;
  assign new_n3339 = new_n3332 ^ new_n3320;
  assign new_n3340 = new_n3339 ^ new_n3338;
  assign new_n3341 = new_n3273 & new_n3340;
  assign new_n3342 = new_n3337 ^ new_n3311;
  assign new_n3343 = new_n3321 & new_n3342;
  assign new_n3344 = new_n3343 ^ new_n3297;
  assign new_n3345 = ~new_n3344 & new_n3300;
  assign new_n3346 = new_n3345 ^ new_n3341;
  assign new_n3347 = new_n3332 ^ new_n3330;
  assign new_n3348 = new_n3347 ^ new_n3315;
  assign new_n3349 = new_n3343 ^ new_n3322;
  assign new_n3350 = new_n3348 & new_n3349;
  assign new_n3351 = new_n3350 ^ new_n3329;
  assign new_n3352 = new_n3277 & new_n3351;
  assign new_n3353 = new_n3343 ^ new_n3337;
  assign new_n3354 = new_n3353 ^ new_n3336;
  assign new_n3355 = ~new_n3354 & new_n3306;
  assign new_n3356 = new_n3274 ^ new_n3268;
  assign new_n3357 = new_n3307 ^ new_n3279;
  assign new_n3358 = new_n3350 ^ new_n3343;
  assign new_n3359 = new_n3358 ^ new_n3357;
  assign new_n3360 = new_n3359 ^ new_n3356;
  assign new_n3361 = new_n3360 ^ new_n3287;
  assign new_n3362 = new_n3330 ^ new_n3283;
  assign new_n3363 = new_n3362 ^ new_n3302;
  assign new_n3364 = new_n3363 ^ new_n3361;
  assign new_n3365 = ~new_n3364 & new_n3290;
  assign new_n3366 = new_n3292 & new_n3340;
  assign new_n3367 = new_n3366 ^ new_n3365;
  assign new_n3368 = new_n3367 ^ new_n3355;
  assign new_n3369 = new_n3368 ^ new_n3352;
  assign new_n3370 = new_n3350 ^ new_n3330;
  assign new_n3371 = new_n3370 ^ new_n3310;
  assign new_n3372 = new_n3280 & new_n3371;
  assign new_n3373 = new_n3372 ^ new_n3369;
  assign new_n3374 = ~new_n3364 & new_n3289;
  assign new_n3375 = new_n3374 ^ new_n3373;
  assign new_n3376 = new_n3375 ^ new_n3346;
  assign new_n3377 = new_n3198 & new_n3257;
  assign new_n3378 = new_n3239 ^ new_n3219;
  assign new_n3379 = new_n3378 ^ new_n3218;
  assign new_n3380 = new_n3208 & new_n3379;
  assign new_n3381 = new_n3380 ^ new_n3263;
  assign new_n3382 = new_n3178 & new_n3245;
  assign new_n3383 = new_n3382 ^ new_n3381;
  assign new_n3384 = new_n3383 ^ new_n3235;
  assign new_n3385 = new_n3384 ^ new_n3377;
  assign new_n3386 = new_n3186 & new_n3240;
  assign new_n3387 = new_n3163 & new_n3261;
  assign new_n3388 = new_n3387 ^ new_n3386;
  assign new_n3389 = new_n3388 ^ new_n3385;
  assign new_n3390 = new_n3389 ^ new_n3376;
  assign new_n3391 = new_n3390 ^ new_n3266;
  assign new_n3392 = new_n3337 ^ new_n3321;
  assign new_n3393 = new_n3276 & new_n3392;
  assign new_n3394 = ~new_n3344 & new_n3298;
  assign new_n3395 = new_n3394 ^ new_n3393;
  assign new_n3396 = new_n3282 & new_n3371;
  assign new_n3397 = new_n3396 ^ new_n3395;
  assign new_n3398 = new_n3397 ^ new_n3372;
  assign new_n3399 = new_n3305 & new_n3351;
  assign new_n3400 = new_n3317 & new_n3348;
  assign new_n3401 = new_n3400 ^ new_n3399;
  assign new_n3402 = new_n3401 ^ new_n3367;
  assign new_n3403 = new_n3402 ^ new_n3398;
  assign new_n3404 = new_n1326 & new_n1391;
  assign new_n3405 = new_n1363 ^ n17;
  assign new_n3406 = new_n1348 ^ new_n1302;
  assign new_n3407 = new_n3406 ^ new_n1374;
  assign new_n3408 = new_n3407 ^ new_n3405;
  assign new_n3409 = ~new_n3408 & new_n1316;
  assign new_n3410 = new_n3409 ^ new_n3404;
  assign new_n3411 = ~new_n1378 & new_n1313;
  assign new_n3412 = new_n3411 ^ new_n1369;
  assign new_n3413 = new_n1346 & new_n1358;
  assign new_n3414 = new_n1307 & new_n1368;
  assign new_n3415 = new_n3414 ^ new_n3413;
  assign new_n3416 = new_n3415 ^ new_n1384;
  assign new_n3417 = new_n3416 ^ new_n3412;
  assign new_n3418 = new_n3417 ^ new_n3410;
  assign new_n3419 = new_n3418 ^ n127;
  assign new_n3420 = new_n3419 ^ n95;
  assign new_n3421 = new_n3420 ^ n63;
  assign new_n3422 = new_n3421 ^ new_n3403;
  assign new_n3423 = new_n3219 ^ new_n3165;
  assign new_n3424 = new_n3225 ^ new_n3181;
  assign new_n3425 = new_n3424 ^ new_n3253;
  assign new_n3426 = new_n3425 ^ new_n3423;
  assign new_n3427 = new_n3171 & new_n3426;
  assign new_n3428 = new_n3427 ^ new_n3236;
  assign new_n3429 = new_n3382 ^ new_n3377;
  assign new_n3430 = new_n3429 ^ new_n3264;
  assign new_n3431 = new_n3430 ^ new_n3428;
  assign new_n3432 = new_n3431 ^ new_n3422;
  assign new_n3433 = new_n3432 ^ new_n3391;
  assign new_n3434 = new_n3082 & new_n3148;
  assign new_n3435 = new_n3117 ^ new_n3087;
  assign new_n3436 = ~new_n3435 & new_n3089;
  assign new_n3437 = new_n3436 ^ new_n3434;
  assign new_n3438 = new_n3117 ^ new_n3115;
  assign new_n3439 = new_n3438 ^ new_n3114;
  assign new_n3440 = ~new_n3439 & new_n3061;
  assign new_n3441 = new_n3440 ^ new_n3150;
  assign new_n3442 = new_n3441 ^ new_n3135;
  assign new_n3443 = new_n3078 & new_n3121;
  assign new_n3444 = new_n3443 ^ new_n3442;
  assign new_n3445 = new_n3444 ^ new_n3140;
  assign new_n3446 = new_n3445 ^ new_n3437;
  assign new_n3447 = new_n3006 ^ new_n3004;
  assign new_n3448 = new_n3447 ^ new_n3003;
  assign new_n3449 = ~new_n3448 & new_n2950;
  assign new_n3450 = new_n3449 ^ new_n3039;
  assign new_n3451 = new_n3450 ^ new_n3024;
  assign new_n3452 = new_n2967 & new_n3010;
  assign new_n3453 = new_n3452 ^ new_n3451;
  assign new_n3454 = new_n3453 ^ new_n3029;
  assign new_n3455 = new_n3006 ^ new_n2976;
  assign new_n3456 = ~new_n3455 & new_n2978;
  assign new_n3457 = new_n2971 & new_n3037;
  assign new_n3458 = new_n3457 ^ new_n3456;
  assign new_n3459 = new_n3458 ^ new_n3454;
  assign new_n3460 = new_n3459 ^ new_n3446;
  assign new_n3461 = new_n3387 ^ new_n3377;
  assign new_n3462 = new_n3206 & new_n3379;
  assign new_n3463 = new_n3462 ^ new_n3241;
  assign new_n3464 = new_n3463 ^ new_n3386;
  assign new_n3465 = new_n3464 ^ new_n3381;
  assign new_n3466 = new_n3465 ^ new_n3461;
  assign new_n3467 = new_n3466 ^ new_n3460;
  assign new_n3468 = new_n3411 ^ new_n1393;
  assign new_n3469 = new_n1330 & new_n1382;
  assign new_n3470 = new_n3469 ^ new_n1395;
  assign new_n3471 = new_n3470 ^ new_n3468;
  assign new_n3472 = new_n3471 ^ n89;
  assign new_n3473 = new_n3472 ^ n121;
  assign new_n3474 = new_n3473 ^ n57;
  assign new_n3475 = new_n3474 ^ new_n3389;
  assign new_n3476 = new_n3374 ^ new_n3341;
  assign new_n3477 = ~new_n3354 & new_n3304;
  assign new_n3478 = new_n3477 ^ new_n3394;
  assign new_n3479 = new_n3478 ^ new_n3345;
  assign new_n3480 = new_n3479 ^ new_n3368;
  assign new_n3481 = new_n3480 ^ new_n3476;
  assign new_n3482 = new_n3481 ^ new_n3475;
  assign new_n3483 = new_n3482 ^ new_n3467;
  assign new_n3484 = new_n3483 ^ new_n3433;
  assign new_n3485 = new_n3115 ^ new_n3104;
  assign new_n3486 = new_n3063 & new_n3485;
  assign new_n3487 = new_n3486 ^ new_n3445;
  assign new_n3488 = new_n3048 & new_n3485;
  assign new_n3489 = ~new_n3435 & new_n3053;
  assign new_n3490 = new_n3489 ^ new_n3488;
  assign new_n3491 = new_n3490 ^ new_n3122;
  assign new_n3492 = new_n3100 & new_n3110;
  assign new_n3493 = new_n3492 ^ new_n3132;
  assign new_n3494 = new_n3493 ^ new_n3491;
  assign new_n3495 = new_n3494 ^ new_n3487;
  assign new_n3496 = new_n3004 ^ new_n2993;
  assign new_n3497 = new_n2952 & new_n3496;
  assign new_n3498 = new_n3497 ^ new_n3454;
  assign new_n3499 = new_n2942 & new_n3496;
  assign new_n3500 = ~new_n3455 & new_n2941;
  assign new_n3501 = new_n3500 ^ new_n3499;
  assign new_n3502 = new_n3501 ^ new_n3011;
  assign new_n3503 = new_n2989 & new_n2999;
  assign new_n3504 = new_n3503 ^ new_n3021;
  assign new_n3505 = new_n3504 ^ new_n3502;
  assign new_n3506 = new_n3505 ^ new_n3498;
  assign new_n3507 = new_n3506 ^ new_n3495;
  assign new_n3508 = new_n3507 ^ new_n3431;
  assign new_n3509 = new_n3178 ^ new_n3164;
  assign new_n3510 = new_n3237 & new_n3509;
  assign new_n3511 = new_n3510 ^ new_n3385;
  assign new_n3512 = new_n3179 & new_n3231;
  assign new_n3513 = new_n3512 ^ new_n3427;
  assign new_n3514 = new_n3513 ^ new_n3243;
  assign new_n3515 = new_n3514 ^ new_n3511;
  assign new_n3516 = new_n1363 ^ new_n1353;
  assign new_n3517 = new_n1297 ^ n20;
  assign new_n3518 = new_n3516 & new_n3517;
  assign new_n3519 = new_n3518 ^ new_n3468;
  assign new_n3520 = n24 & new_n3516;
  assign new_n3521 = new_n3520 ^ new_n1397;
  assign new_n3522 = new_n3521 ^ new_n3404;
  assign new_n3523 = new_n1347 & new_n1358;
  assign new_n3524 = new_n3523 ^ new_n3409;
  assign new_n3525 = new_n3524 ^ new_n3522;
  assign new_n3526 = new_n3525 ^ new_n3519;
  assign new_n3527 = new_n3526 ^ n94;
  assign new_n3528 = new_n3527 ^ n126;
  assign new_n3529 = new_n3528 ^ n62;
  assign new_n3530 = new_n3529 ^ new_n3515;
  assign new_n3531 = new_n3337 ^ new_n3281;
  assign new_n3532 = new_n3325 ^ new_n3318;
  assign new_n3533 = new_n3532 ^ new_n3360;
  assign new_n3534 = new_n3533 ^ new_n3531;
  assign new_n3535 = ~new_n3534 & new_n3312;
  assign new_n3536 = new_n3535 ^ new_n3396;
  assign new_n3537 = new_n3374 ^ new_n3352;
  assign new_n3538 = new_n3537 ^ new_n3402;
  assign new_n3539 = new_n3538 ^ new_n3536;
  assign new_n3540 = new_n3539 ^ new_n3530;
  assign new_n3541 = new_n3540 ^ new_n3508;
  assign new_n3542 = ~new_n3439 & new_n3054;
  assign new_n3543 = new_n3542 ^ new_n3489;
  assign new_n3544 = new_n3543 ^ new_n3436;
  assign new_n3545 = new_n3544 ^ new_n3444;
  assign new_n3546 = ~new_n3448 & new_n2943;
  assign new_n3547 = new_n3546 ^ new_n3500;
  assign new_n3548 = new_n3547 ^ new_n3456;
  assign new_n3549 = new_n3548 ^ new_n3453;
  assign new_n3550 = new_n3549 ^ new_n3545;
  assign new_n3551 = new_n1400 ^ n92;
  assign new_n3552 = new_n3551 ^ n124;
  assign new_n3553 = new_n3552 ^ n60;
  assign new_n3554 = new_n3553 ^ new_n3550;
  assign new_n3555 = new_n3554 ^ new_n3390;
  assign new_n3556 = new_n3386 ^ new_n3247;
  assign new_n3557 = new_n3462 ^ new_n3238;
  assign new_n3558 = new_n3557 ^ new_n3383;
  assign new_n3559 = new_n3558 ^ new_n3556;
  assign new_n3560 = new_n3464 ^ new_n3384;
  assign new_n3561 = new_n3560 ^ new_n3559;
  assign new_n3562 = new_n3400 ^ new_n3345;
  assign new_n3563 = new_n3477 ^ new_n3393;
  assign new_n3564 = new_n3563 ^ new_n3369;
  assign new_n3565 = new_n3564 ^ new_n3562;
  assign new_n3566 = new_n3565 ^ new_n3561;
  assign new_n3567 = new_n3566 ^ new_n3555;
  assign new_n3568 = new_n3567 ^ new_n3541;
  assign new_n3569 = new_n3568 ^ new_n3484;
  assign new_n3570 = new_n3567 ^ new_n3483;
  assign new_n3571 = new_n3559 ^ new_n3515;
  assign new_n3572 = new_n3324 & new_n3392;
  assign new_n3573 = new_n3572 ^ new_n3375;
  assign new_n3574 = new_n3316 & new_n3348;
  assign new_n3575 = new_n3574 ^ new_n3535;
  assign new_n3576 = new_n3575 ^ new_n3397;
  assign new_n3577 = new_n3576 ^ new_n3573;
  assign new_n3578 = new_n3577 ^ new_n3571;
  assign new_n3579 = new_n3436 ^ new_n3142;
  assign new_n3580 = new_n3542 ^ new_n3488;
  assign new_n3581 = new_n3580 ^ new_n3442;
  assign new_n3582 = new_n3581 ^ new_n3579;
  assign new_n3583 = new_n3456 ^ new_n3031;
  assign new_n3584 = new_n3546 ^ new_n3499;
  assign new_n3585 = new_n3584 ^ new_n3451;
  assign new_n3586 = new_n3585 ^ new_n3583;
  assign new_n3587 = new_n3586 ^ new_n3582;
  assign new_n3588 = new_n3413 ^ new_n1395;
  assign new_n3589 = new_n3520 ^ new_n1396;
  assign new_n3590 = new_n3589 ^ new_n1389;
  assign new_n3591 = new_n3590 ^ new_n3588;
  assign new_n3592 = new_n3591 ^ n93;
  assign new_n3593 = new_n3592 ^ n125;
  assign new_n3594 = new_n3593 ^ n61;
  assign new_n3595 = new_n3594 ^ new_n3587;
  assign new_n3596 = new_n3595 ^ new_n3390;
  assign new_n3597 = new_n3596 ^ new_n3578;
  assign new_n3598 = new_n3597 ^ new_n3433;
  assign new_n3599 = new_n3598 ^ new_n3541;
  assign new_n3600 = new_n3434 ^ new_n3140;
  assign new_n3601 = new_n3544 ^ new_n3441;
  assign new_n3602 = new_n3601 ^ new_n3600;
  assign new_n3603 = new_n3457 ^ new_n3029;
  assign new_n3604 = new_n3548 ^ new_n3450;
  assign new_n3605 = new_n3604 ^ new_n3603;
  assign new_n3606 = new_n3605 ^ new_n3602;
  assign new_n3607 = new_n3387 ^ new_n3262;
  assign new_n3608 = new_n3168 & new_n3426;
  assign new_n3609 = new_n3608 ^ new_n3514;
  assign new_n3610 = new_n3609 ^ new_n3607;
  assign new_n3611 = new_n3610 ^ new_n3606;
  assign new_n3612 = new_n3366 ^ new_n3341;
  assign new_n3613 = ~new_n3534 & new_n3285;
  assign new_n3614 = new_n3613 ^ new_n3576;
  assign new_n3615 = new_n3614 ^ new_n3612;
  assign new_n3616 = new_n3469 ^ new_n3411;
  assign new_n3617 = new_n1399 ^ new_n1388;
  assign new_n3618 = new_n3617 ^ new_n3616;
  assign new_n3619 = new_n3618 ^ n122;
  assign new_n3620 = new_n3619 ^ n90;
  assign new_n3621 = new_n3620 ^ n58;
  assign new_n3622 = new_n3621 ^ new_n3615;
  assign new_n3623 = new_n3622 ^ new_n3466;
  assign new_n3624 = new_n3623 ^ new_n3611;
  assign new_n3625 = new_n3624 ^ new_n3599;
  assign new_n3626 = new_n3570 & new_n3625;
  assign new_n3627 = new_n3541 ^ new_n3483;
  assign new_n3628 = new_n3434 ^ new_n3149;
  assign new_n3629 = ~new_n3131 & new_n3060;
  assign new_n3630 = new_n3629 ^ new_n3494;
  assign new_n3631 = new_n3630 ^ new_n3628;
  assign new_n3632 = new_n3457 ^ new_n3038;
  assign new_n3633 = ~new_n3020 & new_n2949;
  assign new_n3634 = new_n3633 ^ new_n3505;
  assign new_n3635 = new_n3634 ^ new_n3632;
  assign new_n3636 = new_n3635 ^ new_n3631;
  assign new_n3637 = new_n3636 ^ new_n3610;
  assign new_n3638 = new_n3479 ^ new_n3373;
  assign new_n3639 = new_n3638 ^ new_n3560;
  assign new_n3640 = new_n3469 ^ new_n1383;
  assign new_n3641 = ~new_n3408 & new_n1308;
  assign new_n3642 = new_n3641 ^ new_n3525;
  assign new_n3643 = new_n3642 ^ new_n3640;
  assign new_n3644 = new_n3643 ^ n91;
  assign new_n3645 = new_n3644 ^ n123;
  assign new_n3646 = new_n3645 ^ n59;
  assign new_n3647 = new_n3646 ^ new_n3639;
  assign new_n3648 = new_n3647 ^ new_n3637;
  assign new_n3649 = new_n3648 ^ new_n3624;
  assign new_n3650 = new_n3598 ^ new_n3570;
  assign new_n3651 = new_n3650 ^ new_n3649;
  assign new_n3652 = new_n3627 & new_n3651;
  assign new_n3653 = new_n3652 ^ new_n3626;
  assign new_n3654 = new_n3648 ^ new_n3599;
  assign new_n3655 = new_n3654 ^ new_n3653;
  assign new_n3656 = new_n3484 & new_n3654;
  assign new_n3657 = new_n3522 ^ new_n1392;
  assign new_n3658 = new_n3657 ^ new_n3416;
  assign new_n3659 = new_n3658 ^ n128;
  assign new_n3660 = new_n3659 ^ n96;
  assign new_n3661 = new_n3660 ^ n64;
  assign new_n3662 = new_n3661 ^ new_n3265;
  assign new_n3663 = new_n3502 ^ new_n3452;
  assign new_n3664 = new_n3663 ^ new_n3040;
  assign new_n3665 = new_n3491 ^ new_n3443;
  assign new_n3666 = new_n3665 ^ new_n3151;
  assign new_n3667 = new_n3666 ^ new_n3664;
  assign new_n3668 = new_n3667 ^ new_n3390;
  assign new_n3669 = new_n3668 ^ new_n3662;
  assign new_n3670 = new_n3669 ^ new_n3649;
  assign new_n3671 = new_n3670 ^ new_n3483;
  assign new_n3672 = new_n3669 ^ new_n3625;
  assign new_n3673 = ~new_n3671 & ~new_n3672;
  assign new_n3674 = new_n3673 ^ new_n3656;
  assign new_n3675 = new_n3674 ^ new_n3483;
  assign new_n3676 = new_n3675 ^ new_n3655;
  assign new_n3677 = new_n3569 & new_n3650;
  assign new_n3678 = new_n3677 ^ new_n3624;
  assign new_n3679 = ~new_n3649 & ~new_n3669;
  assign new_n3680 = new_n3567 & new_n3669;
  assign new_n3681 = new_n3680 ^ new_n3679;
  assign new_n3682 = new_n3681 ^ new_n3678;
  assign new_n3683 = ~new_n3433 & new_n3670;
  assign new_n3684 = new_n3683 ^ new_n3433;
  assign new_n3685 = new_n3684 ^ new_n3656;
  assign new_n3686 = new_n3685 ^ new_n3627;
  assign new_n3687 = new_n3648 ^ new_n3567;
  assign new_n3688 = new_n3687 ^ new_n3627;
  assign new_n3689 = new_n3568 & new_n3688;
  assign new_n3690 = new_n3689 ^ new_n3626;
  assign new_n3691 = new_n3648 ^ new_n3597;
  assign new_n3692 = new_n3691 ^ new_n3690;
  assign new_n3693 = new_n3692 ^ new_n3686;
  assign new_n3694 = new_n3678 ^ new_n3650;
  assign new_n3695 = new_n3669 ^ new_n3650;
  assign new_n3696 = new_n3670 ^ new_n3433;
  assign new_n3697 = new_n3696 ^ new_n3627;
  assign new_n3698 = ~new_n3695 & ~new_n3697;
  assign new_n3699 = new_n3698 ^ new_n3626;
  assign new_n3700 = new_n3689 ^ new_n3541;
  assign new_n3701 = new_n3700 ^ new_n3699;
  assign new_n3702 = new_n3701 ^ new_n3694;
  assign new_n3703 = ~new_n3693 & new_n3702;
  assign new_n3704 = new_n3703 ^ new_n3682;
  assign new_n3705 = new_n3704 ^ new_n3655;
  assign new_n3706 = new_n3683 ^ new_n3673;
  assign new_n3707 = new_n3689 ^ new_n3652;
  assign new_n3708 = new_n3707 ^ new_n3706;
  assign new_n3709 = ~new_n3708 & new_n3705;
  assign new_n3710 = new_n3709 ^ new_n3703;
  assign new_n3711 = new_n3676 & new_n3710;
  assign new_n3712 = new_n3711 ^ new_n3693;
  assign new_n3713 = ~new_n3712 & new_n3569;
  assign new_n3714 = new_n3648 ^ new_n3483;
  assign new_n3715 = new_n3681 ^ new_n3567;
  assign new_n3716 = new_n3715 ^ new_n3698;
  assign new_n3717 = new_n3716 ^ new_n3707;
  assign new_n3718 = new_n3717 ^ new_n3714;
  assign new_n3719 = new_n3703 ^ new_n3676;
  assign new_n3720 = new_n3718 & new_n3719;
  assign new_n3721 = new_n3720 ^ new_n3709;
  assign new_n3722 = new_n3682 ^ new_n3675;
  assign new_n3723 = new_n3722 ^ new_n3721;
  assign new_n3724 = new_n3625 & new_n3723;
  assign new_n3725 = new_n3724 ^ new_n3713;
  assign new_n3726 = new_n3720 ^ new_n3682;
  assign new_n3727 = new_n3726 ^ new_n3655;
  assign new_n3728 = new_n3719 ^ new_n3711;
  assign new_n3729 = new_n3727 & new_n3728;
  assign new_n3730 = new_n3729 ^ new_n3720;
  assign new_n3731 = new_n3730 ^ new_n3702;
  assign new_n3732 = new_n3654 & new_n3731;
  assign new_n3733 = new_n3729 ^ new_n3718;
  assign new_n3734 = ~new_n3670 & new_n3733;
  assign new_n3735 = new_n3711 ^ new_n3709;
  assign new_n3736 = new_n3735 ^ new_n3708;
  assign new_n3737 = ~new_n3697 & ~new_n3736;
  assign new_n3738 = new_n3570 & new_n3723;
  assign new_n3739 = new_n3648 ^ new_n3433;
  assign new_n3740 = new_n3698 ^ new_n3684;
  assign new_n3741 = new_n3729 ^ new_n3711;
  assign new_n3742 = new_n3741 ^ new_n3740;
  assign new_n3743 = new_n3742 ^ new_n3739;
  assign new_n3744 = new_n3743 ^ new_n3567;
  assign new_n3745 = new_n3720 ^ new_n3656;
  assign new_n3746 = new_n3745 ^ new_n3678;
  assign new_n3747 = new_n3746 ^ new_n3744;
  assign new_n3748 = ~new_n3747 & new_n3568;
  assign new_n3749 = new_n3748 ^ new_n3738;
  assign new_n3750 = new_n3749 ^ new_n3737;
  assign new_n3751 = new_n3750 ^ new_n3734;
  assign new_n3752 = new_n3751 ^ new_n3732;
  assign new_n3753 = ~new_n3747 & new_n3688;
  assign new_n3754 = new_n3753 ^ new_n3752;
  assign new_n3755 = new_n3754 ^ new_n3725;
  assign new_n3756 = n203 ^ n75;
  assign new_n3757 = n202 ^ n74;
  assign new_n3758 = new_n3757 ^ new_n3756;
  assign new_n3759 = n208 ^ n80;
  assign new_n3760 = new_n3759 ^ new_n3758;
  assign new_n3761 = n204 ^ n76;
  assign new_n3762 = new_n3761 ^ new_n3760;
  assign new_n3763 = new_n3759 & new_n3762;
  assign new_n3764 = new_n3763 ^ new_n3761;
  assign new_n3765 = n207 ^ n79;
  assign new_n3766 = n205 ^ n77;
  assign new_n3767 = new_n3766 ^ new_n3765;
  assign new_n3768 = n201 ^ n73;
  assign new_n3769 = new_n3768 ^ new_n3761;
  assign new_n3770 = new_n3769 ^ new_n3767;
  assign new_n3771 = new_n3765 ^ new_n3761;
  assign new_n3772 = n206 ^ n78;
  assign new_n3773 = new_n3772 ^ new_n3768;
  assign new_n3774 = new_n3773 ^ new_n3771;
  assign new_n3775 = new_n3770 & new_n3774;
  assign new_n3776 = new_n3775 ^ new_n3757;
  assign new_n3777 = new_n3776 ^ new_n3764;
  assign new_n3778 = ~new_n3760 & ~new_n3765;
  assign new_n3779 = new_n3778 ^ new_n3765;
  assign new_n3780 = new_n3772 ^ new_n3767;
  assign new_n3781 = new_n3780 ^ new_n3756;
  assign new_n3782 = new_n3768 ^ new_n3765;
  assign new_n3783 = new_n3781 & new_n3782;
  assign new_n3784 = new_n3783 ^ new_n3779;
  assign new_n3785 = new_n3784 ^ new_n3773;
  assign new_n3786 = new_n3761 ^ new_n3756;
  assign new_n3787 = new_n3786 ^ new_n3773;
  assign new_n3788 = new_n3772 ^ new_n3761;
  assign new_n3789 = new_n3787 & new_n3788;
  assign new_n3790 = new_n3780 ^ new_n3757;
  assign new_n3791 = new_n3769 & new_n3790;
  assign new_n3792 = new_n3791 ^ new_n3789;
  assign new_n3793 = new_n3766 ^ new_n3756;
  assign new_n3794 = new_n3793 ^ new_n3792;
  assign new_n3795 = new_n3794 ^ new_n3785;
  assign new_n3796 = new_n3776 ^ new_n3770;
  assign new_n3797 = new_n3770 ^ new_n3759;
  assign new_n3798 = new_n3765 ^ new_n3760;
  assign new_n3799 = new_n3798 ^ new_n3773;
  assign new_n3800 = new_n3797 & new_n3799;
  assign new_n3801 = new_n3800 ^ new_n3772;
  assign new_n3802 = new_n3801 ^ new_n3792;
  assign new_n3803 = new_n3802 ^ new_n3796;
  assign new_n3804 = ~new_n3795 & new_n3803;
  assign new_n3805 = new_n3804 ^ new_n3777;
  assign new_n3806 = new_n3770 ^ new_n3758;
  assign new_n3807 = new_n3773 & new_n3806;
  assign new_n3808 = new_n3807 ^ new_n3791;
  assign new_n3809 = new_n3808 ^ new_n3781;
  assign new_n3810 = new_n3809 ^ new_n3805;
  assign new_n3811 = new_n3807 ^ new_n3789;
  assign new_n3812 = new_n3790 ^ new_n3759;
  assign new_n3813 = new_n3768 ^ new_n3760;
  assign new_n3814 = new_n3812 & new_n3813;
  assign new_n3815 = new_n3814 ^ new_n3778;
  assign new_n3816 = new_n3815 ^ new_n3811;
  assign new_n3817 = ~new_n3816 & new_n3810;
  assign new_n3818 = new_n3814 ^ new_n3783;
  assign new_n3819 = new_n3818 ^ new_n3768;
  assign new_n3820 = new_n3819 ^ new_n3809;
  assign new_n3821 = new_n3820 ^ new_n3817;
  assign new_n3822 = new_n3762 & new_n3821;
  assign new_n3823 = new_n3765 ^ new_n3756;
  assign new_n3824 = new_n3800 ^ new_n3779;
  assign new_n3825 = new_n3817 ^ new_n3804;
  assign new_n3826 = ~new_n3820 & ~new_n3825;
  assign new_n3827 = new_n3826 ^ new_n3817;
  assign new_n3828 = new_n3820 ^ new_n3804;
  assign new_n3829 = new_n3768 ^ new_n3756;
  assign new_n3830 = new_n3800 ^ new_n3763;
  assign new_n3831 = new_n3830 ^ new_n3811;
  assign new_n3832 = new_n3831 ^ new_n3829;
  assign new_n3833 = new_n3828 & new_n3832;
  assign new_n3834 = new_n3833 ^ new_n3777;
  assign new_n3835 = new_n3834 ^ new_n3809;
  assign new_n3836 = ~new_n3827 & new_n3835;
  assign new_n3837 = new_n3828 ^ new_n3827;
  assign new_n3838 = new_n3837 ^ new_n3836;
  assign new_n3839 = new_n3838 ^ new_n3824;
  assign new_n3840 = new_n3839 ^ new_n3823;
  assign new_n3841 = new_n3840 ^ new_n3761;
  assign new_n3842 = new_n3833 ^ new_n3783;
  assign new_n3843 = new_n3842 ^ new_n3776;
  assign new_n3844 = new_n3843 ^ new_n3841;
  assign new_n3845 = new_n3787 & new_n3844;
  assign new_n3846 = new_n3836 ^ new_n3833;
  assign new_n3847 = new_n3846 ^ new_n3803;
  assign new_n3848 = new_n3781 & new_n3847;
  assign new_n3849 = new_n3837 ^ new_n3817;
  assign new_n3850 = new_n3849 ^ new_n3816;
  assign new_n3851 = new_n3799 & new_n3850;
  assign new_n3852 = new_n3833 ^ new_n3817;
  assign new_n3853 = new_n3819 ^ new_n3777;
  assign new_n3854 = new_n3853 ^ new_n3852;
  assign new_n3855 = new_n3769 & new_n3854;
  assign new_n3856 = new_n3788 & new_n3844;
  assign new_n3857 = new_n3856 ^ new_n3855;
  assign new_n3858 = new_n3857 ^ new_n3851;
  assign new_n3859 = new_n3836 ^ new_n3832;
  assign new_n3860 = new_n3760 & new_n3859;
  assign new_n3861 = new_n3860 ^ new_n3858;
  assign new_n3862 = new_n3861 ^ new_n3848;
  assign new_n3863 = new_n3862 ^ new_n3845;
  assign new_n3864 = new_n3863 ^ new_n3822;
  assign new_n3865 = new_n3759 & new_n3821;
  assign new_n3866 = new_n3837 ^ new_n3795;
  assign new_n3867 = new_n3770 & new_n3866;
  assign new_n3868 = new_n3867 ^ new_n3865;
  assign new_n3869 = new_n3782 & new_n3847;
  assign new_n3870 = new_n3869 ^ new_n3868;
  assign new_n3871 = new_n3813 & new_n3835;
  assign new_n3872 = new_n3817 ^ new_n3768;
  assign new_n3873 = new_n3814 ^ new_n3763;
  assign new_n3874 = new_n3873 ^ new_n3840;
  assign new_n3875 = new_n3874 ^ new_n3872;
  assign new_n3876 = new_n3806 & new_n3875;
  assign new_n3877 = new_n3876 ^ new_n3871;
  assign new_n3878 = new_n3877 ^ new_n3870;
  assign new_n3879 = new_n3878 ^ new_n3864;
  assign new_n3880 = new_n3812 & new_n3835;
  assign new_n3881 = new_n3774 & new_n3866;
  assign new_n3882 = new_n3881 ^ new_n3880;
  assign new_n3883 = new_n3797 & new_n3850;
  assign new_n3884 = new_n3883 ^ new_n3865;
  assign new_n3885 = new_n3884 ^ new_n3861;
  assign new_n3886 = new_n3885 ^ new_n3882;
  assign new_n3887 = new_n3886 ^ new_n3879;
  assign new_n3888 = n244 ^ n116;
  assign new_n3889 = n243 ^ n115;
  assign new_n3890 = n242 ^ n114;
  assign new_n3891 = new_n3890 ^ new_n3889;
  assign new_n3892 = n248 ^ n120;
  assign new_n3893 = new_n3892 ^ new_n3891;
  assign new_n3894 = new_n3893 ^ new_n3888;
  assign new_n3895 = n247 ^ n119;
  assign new_n3896 = ~new_n3893 & ~new_n3895;
  assign new_n3897 = new_n3896 ^ new_n3895;
  assign new_n3898 = n245 ^ n117;
  assign new_n3899 = new_n3898 ^ new_n3895;
  assign new_n3900 = n246 ^ n118;
  assign new_n3901 = new_n3900 ^ new_n3899;
  assign new_n3902 = new_n3901 ^ new_n3889;
  assign new_n3903 = n241 ^ n113;
  assign new_n3904 = new_n3903 ^ new_n3895;
  assign new_n3905 = new_n3902 & new_n3904;
  assign new_n3906 = new_n3905 ^ new_n3897;
  assign new_n3907 = new_n3903 ^ new_n3900;
  assign new_n3908 = new_n3907 ^ new_n3906;
  assign new_n3909 = new_n3889 ^ new_n3888;
  assign new_n3910 = new_n3909 ^ new_n3907;
  assign new_n3911 = new_n3900 ^ new_n3888;
  assign new_n3912 = new_n3910 & new_n3911;
  assign new_n3913 = new_n3901 ^ new_n3890;
  assign new_n3914 = new_n3903 ^ new_n3888;
  assign new_n3915 = new_n3913 & new_n3914;
  assign new_n3916 = new_n3915 ^ new_n3912;
  assign new_n3917 = new_n3898 ^ new_n3889;
  assign new_n3918 = new_n3917 ^ new_n3916;
  assign new_n3919 = new_n3918 ^ new_n3908;
  assign new_n3920 = new_n3914 ^ new_n3899;
  assign new_n3921 = new_n3895 ^ new_n3888;
  assign new_n3922 = new_n3921 ^ new_n3907;
  assign new_n3923 = new_n3920 & new_n3922;
  assign new_n3924 = new_n3923 ^ new_n3890;
  assign new_n3925 = new_n3924 ^ new_n3920;
  assign new_n3926 = new_n3920 ^ new_n3892;
  assign new_n3927 = new_n3895 ^ new_n3893;
  assign new_n3928 = new_n3927 ^ new_n3907;
  assign new_n3929 = new_n3926 & new_n3928;
  assign new_n3930 = new_n3929 ^ new_n3900;
  assign new_n3931 = new_n3930 ^ new_n3916;
  assign new_n3932 = new_n3931 ^ new_n3925;
  assign new_n3933 = ~new_n3919 & new_n3932;
  assign new_n3934 = new_n3892 & new_n3894;
  assign new_n3935 = new_n3934 ^ new_n3888;
  assign new_n3936 = new_n3935 ^ new_n3924;
  assign new_n3937 = new_n3936 ^ new_n3933;
  assign new_n3938 = new_n3920 ^ new_n3891;
  assign new_n3939 = new_n3907 & new_n3938;
  assign new_n3940 = new_n3939 ^ new_n3915;
  assign new_n3941 = new_n3940 ^ new_n3902;
  assign new_n3942 = new_n3941 ^ new_n3937;
  assign new_n3943 = new_n3913 ^ new_n3892;
  assign new_n3944 = new_n3903 ^ new_n3893;
  assign new_n3945 = new_n3943 & new_n3944;
  assign new_n3946 = new_n3945 ^ new_n3896;
  assign new_n3947 = new_n3939 ^ new_n3912;
  assign new_n3948 = new_n3947 ^ new_n3946;
  assign new_n3949 = ~new_n3948 & new_n3942;
  assign new_n3950 = new_n3945 ^ new_n3905;
  assign new_n3951 = new_n3950 ^ new_n3903;
  assign new_n3952 = new_n3951 ^ new_n3941;
  assign new_n3953 = new_n3952 ^ new_n3949;
  assign new_n3954 = new_n3894 & new_n3953;
  assign new_n3955 = new_n3903 ^ new_n3889;
  assign new_n3956 = new_n3934 ^ new_n3929;
  assign new_n3957 = new_n3956 ^ new_n3947;
  assign new_n3958 = new_n3957 ^ new_n3955;
  assign new_n3959 = new_n3952 ^ new_n3933;
  assign new_n3960 = new_n3958 & new_n3959;
  assign new_n3961 = new_n3960 ^ new_n3936;
  assign new_n3962 = new_n3961 ^ new_n3941;
  assign new_n3963 = new_n3949 ^ new_n3933;
  assign new_n3964 = ~new_n3963 & new_n3952;
  assign new_n3965 = new_n3964 ^ new_n3933;
  assign new_n3966 = new_n3962 & new_n3965;
  assign new_n3967 = new_n3966 ^ new_n3958;
  assign new_n3968 = new_n3893 & new_n3967;
  assign new_n3969 = new_n3964 ^ new_n3952;
  assign new_n3970 = new_n3969 ^ new_n3949;
  assign new_n3971 = new_n3970 ^ new_n3948;
  assign new_n3972 = ~new_n3971 & new_n3928;
  assign new_n3973 = new_n3895 ^ new_n3889;
  assign new_n3974 = new_n3929 ^ new_n3897;
  assign new_n3975 = new_n3969 ^ new_n3966;
  assign new_n3976 = new_n3975 ^ new_n3974;
  assign new_n3977 = new_n3976 ^ new_n3973;
  assign new_n3978 = new_n3977 ^ new_n3888;
  assign new_n3979 = new_n3960 ^ new_n3905;
  assign new_n3980 = new_n3979 ^ new_n3924;
  assign new_n3981 = new_n3980 ^ new_n3978;
  assign new_n3982 = ~new_n3981 & new_n3911;
  assign new_n3983 = new_n3960 ^ new_n3949;
  assign new_n3984 = new_n3951 ^ new_n3936;
  assign new_n3985 = new_n3984 ^ new_n3983;
  assign new_n3986 = new_n3914 & new_n3985;
  assign new_n3987 = new_n3986 ^ new_n3982;
  assign new_n3988 = new_n3987 ^ new_n3972;
  assign new_n3989 = new_n3988 ^ new_n3968;
  assign new_n3990 = new_n3966 ^ new_n3960;
  assign new_n3991 = new_n3990 ^ new_n3932;
  assign new_n3992 = new_n3902 & new_n3991;
  assign new_n3993 = new_n3992 ^ new_n3989;
  assign new_n3994 = ~new_n3981 & new_n3910;
  assign new_n3995 = new_n3994 ^ new_n3993;
  assign new_n3996 = new_n3995 ^ new_n3954;
  assign new_n3997 = new_n3944 & new_n3962;
  assign new_n3998 = new_n3949 ^ new_n3903;
  assign new_n3999 = new_n3945 ^ new_n3934;
  assign new_n4000 = new_n3999 ^ new_n3977;
  assign new_n4001 = new_n4000 ^ new_n3998;
  assign new_n4002 = ~new_n4001 & new_n3938;
  assign new_n4003 = new_n4002 ^ new_n3997;
  assign new_n4004 = new_n3969 ^ new_n3919;
  assign new_n4005 = ~new_n4004 & new_n3920;
  assign new_n4006 = new_n3892 & new_n3953;
  assign new_n4007 = new_n4006 ^ new_n4005;
  assign new_n4008 = new_n3904 & new_n3991;
  assign new_n4009 = new_n4008 ^ new_n4007;
  assign new_n4010 = new_n4009 ^ new_n4003;
  assign new_n4011 = new_n4010 ^ new_n3996;
  assign new_n4012 = new_n4011 ^ new_n3887;
  assign new_n4013 = ~new_n4004 & new_n3922;
  assign new_n4014 = new_n3913 & new_n3985;
  assign new_n4015 = new_n4014 ^ new_n4013;
  assign new_n4016 = new_n4015 ^ new_n3995;
  assign new_n4017 = new_n3790 & new_n3854;
  assign new_n4018 = new_n4017 ^ new_n3881;
  assign new_n4019 = new_n4018 ^ new_n3863;
  assign new_n4020 = new_n4019 ^ new_n4016;
  assign new_n4021 = new_n4020 ^ new_n1175;
  assign new_n4022 = n159 ^ n31;
  assign new_n4023 = n157 ^ n29;
  assign new_n4024 = new_n4023 ^ new_n4022;
  assign new_n4025 = n158 ^ n30;
  assign new_n4026 = new_n4025 ^ new_n4024;
  assign new_n4027 = n154 ^ n26;
  assign new_n4028 = new_n4027 ^ new_n4026;
  assign new_n4029 = n160 ^ n32;
  assign new_n4030 = new_n4029 ^ new_n4028;
  assign new_n4031 = n155 ^ n27;
  assign new_n4032 = n153 ^ n25;
  assign new_n4033 = new_n4032 ^ new_n4031;
  assign new_n4034 = n156 ^ n28;
  assign new_n4035 = new_n4034 ^ new_n4032;
  assign new_n4036 = new_n4035 ^ new_n4024;
  assign new_n4037 = new_n4036 ^ new_n4029;
  assign new_n4038 = new_n4031 ^ new_n4027;
  assign new_n4039 = new_n4038 ^ new_n4029;
  assign new_n4040 = new_n4039 ^ new_n4022;
  assign new_n4041 = new_n4032 ^ new_n4025;
  assign new_n4042 = new_n4041 ^ new_n4040;
  assign new_n4043 = new_n4037 & new_n4042;
  assign new_n4044 = new_n4039 ^ new_n4034;
  assign new_n4045 = new_n4029 & new_n4044;
  assign new_n4046 = new_n4045 ^ new_n4043;
  assign new_n4047 = new_n4034 ^ new_n4025;
  assign new_n4048 = new_n4034 ^ new_n4031;
  assign new_n4049 = new_n4048 ^ new_n4041;
  assign new_n4050 = new_n4047 & new_n4049;
  assign new_n4051 = new_n4038 ^ new_n4036;
  assign new_n4052 = new_n4041 & new_n4051;
  assign new_n4053 = new_n4052 ^ new_n4050;
  assign new_n4054 = new_n4053 ^ new_n4046;
  assign new_n4055 = new_n4054 ^ new_n4033;
  assign new_n4056 = ~new_n4022 & ~new_n4039;
  assign new_n4057 = new_n4056 ^ new_n4022;
  assign new_n4058 = new_n4032 ^ new_n4022;
  assign new_n4059 = new_n4031 ^ new_n4026;
  assign new_n4060 = new_n4058 & new_n4059;
  assign new_n4061 = new_n4060 ^ new_n4057;
  assign new_n4062 = new_n4061 ^ new_n4041;
  assign new_n4063 = new_n4028 & new_n4035;
  assign new_n4064 = new_n4063 ^ new_n4050;
  assign new_n4065 = new_n4031 ^ new_n4023;
  assign new_n4066 = new_n4065 ^ new_n4064;
  assign new_n4067 = new_n4066 ^ new_n4062;
  assign new_n4068 = new_n4058 ^ new_n4047;
  assign new_n4069 = new_n4036 & new_n4068;
  assign new_n4070 = new_n4069 ^ new_n4027;
  assign new_n4071 = new_n4070 ^ new_n4036;
  assign new_n4072 = new_n4043 ^ new_n4025;
  assign new_n4073 = new_n4072 ^ new_n4064;
  assign new_n4074 = new_n4073 ^ new_n4071;
  assign new_n4075 = ~new_n4067 & new_n4074;
  assign new_n4076 = new_n4063 ^ new_n4052;
  assign new_n4077 = new_n4076 ^ new_n4059;
  assign new_n4078 = new_n4039 ^ new_n4032;
  assign new_n4079 = new_n4030 & new_n4078;
  assign new_n4080 = new_n4079 ^ new_n4060;
  assign new_n4081 = new_n4080 ^ new_n4032;
  assign new_n4082 = new_n4081 ^ new_n4077;
  assign new_n4083 = new_n4082 ^ new_n4075;
  assign new_n4084 = new_n4055 & new_n4083;
  assign new_n4085 = new_n4045 ^ new_n4034;
  assign new_n4086 = new_n4085 ^ new_n4070;
  assign new_n4087 = new_n4086 ^ new_n4084;
  assign new_n4088 = new_n4087 ^ new_n4077;
  assign new_n4089 = new_n4030 & new_n4088;
  assign new_n4090 = new_n4086 ^ new_n4075;
  assign new_n4091 = new_n4090 ^ new_n4077;
  assign new_n4092 = new_n4079 ^ new_n4056;
  assign new_n4093 = new_n4092 ^ new_n4053;
  assign new_n4094 = ~new_n4093 & new_n4091;
  assign new_n4095 = new_n4094 ^ new_n4075;
  assign new_n4096 = ~new_n4095 & new_n4082;
  assign new_n4097 = new_n4096 ^ new_n4082;
  assign new_n4098 = new_n4097 ^ new_n4067;
  assign new_n4099 = ~new_n4098 & new_n4068;
  assign new_n4100 = new_n4099 ^ new_n4089;
  assign new_n4101 = new_n4097 ^ new_n4094;
  assign new_n4102 = new_n4101 ^ new_n4093;
  assign new_n4103 = ~new_n4102 & new_n4037;
  assign new_n4104 = new_n4094 ^ new_n4082;
  assign new_n4105 = new_n4029 & new_n4104;
  assign new_n4106 = new_n4105 ^ new_n4103;
  assign new_n4107 = new_n4096 ^ new_n4075;
  assign new_n4108 = new_n4088 & new_n4107;
  assign new_n4109 = new_n4108 ^ new_n4055;
  assign new_n4110 = new_n4039 & new_n4109;
  assign new_n4111 = ~new_n4102 & new_n4042;
  assign new_n4112 = new_n4031 ^ new_n4022;
  assign new_n4113 = new_n4057 ^ new_n4043;
  assign new_n4114 = new_n4108 ^ new_n4097;
  assign new_n4115 = new_n4114 ^ new_n4113;
  assign new_n4116 = new_n4115 ^ new_n4112;
  assign new_n4117 = new_n4116 ^ new_n4034;
  assign new_n4118 = new_n4084 ^ new_n4060;
  assign new_n4119 = new_n4118 ^ new_n4070;
  assign new_n4120 = new_n4119 ^ new_n4117;
  assign new_n4121 = ~new_n4120 & new_n4047;
  assign new_n4122 = new_n4094 ^ new_n4084;
  assign new_n4123 = new_n4086 ^ new_n4081;
  assign new_n4124 = new_n4123 ^ new_n4122;
  assign new_n4125 = new_n4035 & new_n4124;
  assign new_n4126 = new_n4125 ^ new_n4121;
  assign new_n4127 = new_n4126 ^ new_n4111;
  assign new_n4128 = new_n4127 ^ new_n4110;
  assign new_n4129 = new_n4128 ^ new_n4106;
  assign new_n4130 = new_n4129 ^ new_n4100;
  assign new_n4131 = n168 ^ n40;
  assign new_n4132 = n162 ^ n34;
  assign new_n4133 = n167 ^ n39;
  assign new_n4134 = n165 ^ n37;
  assign new_n4135 = new_n4134 ^ new_n4133;
  assign new_n4136 = n166 ^ n38;
  assign new_n4137 = new_n4136 ^ new_n4135;
  assign new_n4138 = new_n4137 ^ new_n4132;
  assign new_n4139 = new_n4138 ^ new_n4131;
  assign new_n4140 = n163 ^ n35;
  assign new_n4141 = n161 ^ n33;
  assign new_n4142 = new_n4141 ^ new_n4140;
  assign new_n4143 = n164 ^ n36;
  assign new_n4144 = new_n4143 ^ new_n4141;
  assign new_n4145 = new_n4144 ^ new_n4135;
  assign new_n4146 = new_n4145 ^ new_n4131;
  assign new_n4147 = new_n4140 ^ new_n4132;
  assign new_n4148 = new_n4147 ^ new_n4131;
  assign new_n4149 = new_n4148 ^ new_n4133;
  assign new_n4150 = new_n4141 ^ new_n4136;
  assign new_n4151 = new_n4150 ^ new_n4149;
  assign new_n4152 = new_n4146 & new_n4151;
  assign new_n4153 = new_n4148 ^ new_n4143;
  assign new_n4154 = new_n4131 & new_n4153;
  assign new_n4155 = new_n4154 ^ new_n4152;
  assign new_n4156 = new_n4143 ^ new_n4140;
  assign new_n4157 = new_n4156 ^ new_n4150;
  assign new_n4158 = new_n4143 ^ new_n4136;
  assign new_n4159 = new_n4157 & new_n4158;
  assign new_n4160 = new_n4147 ^ new_n4145;
  assign new_n4161 = new_n4150 & new_n4160;
  assign new_n4162 = new_n4161 ^ new_n4159;
  assign new_n4163 = new_n4162 ^ new_n4155;
  assign new_n4164 = new_n4163 ^ new_n4142;
  assign new_n4165 = ~new_n4133 & ~new_n4148;
  assign new_n4166 = new_n4165 ^ new_n4133;
  assign new_n4167 = new_n4140 ^ new_n4137;
  assign new_n4168 = new_n4141 ^ new_n4133;
  assign new_n4169 = new_n4167 & new_n4168;
  assign new_n4170 = new_n4169 ^ new_n4166;
  assign new_n4171 = new_n4170 ^ new_n4150;
  assign new_n4172 = new_n4138 & new_n4144;
  assign new_n4173 = new_n4172 ^ new_n4159;
  assign new_n4174 = new_n4140 ^ new_n4134;
  assign new_n4175 = new_n4174 ^ new_n4173;
  assign new_n4176 = new_n4175 ^ new_n4171;
  assign new_n4177 = new_n4143 ^ new_n4133;
  assign new_n4178 = new_n4177 ^ new_n4150;
  assign new_n4179 = new_n4145 & new_n4178;
  assign new_n4180 = new_n4179 ^ new_n4132;
  assign new_n4181 = new_n4180 ^ new_n4145;
  assign new_n4182 = new_n4152 ^ new_n4136;
  assign new_n4183 = new_n4182 ^ new_n4173;
  assign new_n4184 = new_n4183 ^ new_n4181;
  assign new_n4185 = ~new_n4176 & new_n4184;
  assign new_n4186 = new_n4172 ^ new_n4161;
  assign new_n4187 = new_n4186 ^ new_n4167;
  assign new_n4188 = new_n4148 ^ new_n4141;
  assign new_n4189 = new_n4139 & new_n4188;
  assign new_n4190 = new_n4189 ^ new_n4169;
  assign new_n4191 = new_n4190 ^ new_n4141;
  assign new_n4192 = new_n4191 ^ new_n4187;
  assign new_n4193 = new_n4192 ^ new_n4185;
  assign new_n4194 = new_n4164 & new_n4193;
  assign new_n4195 = new_n4154 ^ new_n4143;
  assign new_n4196 = new_n4195 ^ new_n4180;
  assign new_n4197 = new_n4196 ^ new_n4194;
  assign new_n4198 = new_n4197 ^ new_n4187;
  assign new_n4199 = new_n4139 & new_n4198;
  assign new_n4200 = new_n4196 ^ new_n4185;
  assign new_n4201 = new_n4200 ^ new_n4187;
  assign new_n4202 = new_n4189 ^ new_n4165;
  assign new_n4203 = new_n4202 ^ new_n4162;
  assign new_n4204 = ~new_n4203 & new_n4201;
  assign new_n4205 = new_n4204 ^ new_n4185;
  assign new_n4206 = ~new_n4205 & new_n4192;
  assign new_n4207 = new_n4206 ^ new_n4192;
  assign new_n4208 = new_n4207 ^ new_n4176;
  assign new_n4209 = ~new_n4208 & new_n4178;
  assign new_n4210 = new_n4209 ^ new_n4199;
  assign new_n4211 = new_n4207 ^ new_n4204;
  assign new_n4212 = new_n4211 ^ new_n4203;
  assign new_n4213 = ~new_n4212 & new_n4146;
  assign new_n4214 = new_n4204 ^ new_n4192;
  assign new_n4215 = new_n4131 & new_n4214;
  assign new_n4216 = new_n4215 ^ new_n4213;
  assign new_n4217 = ~new_n4212 & new_n4151;
  assign new_n4218 = new_n4140 ^ new_n4133;
  assign new_n4219 = new_n4166 ^ new_n4152;
  assign new_n4220 = new_n4206 ^ new_n4185;
  assign new_n4221 = new_n4198 & new_n4220;
  assign new_n4222 = new_n4221 ^ new_n4207;
  assign new_n4223 = new_n4222 ^ new_n4219;
  assign new_n4224 = new_n4223 ^ new_n4218;
  assign new_n4225 = new_n4224 ^ new_n4143;
  assign new_n4226 = new_n4194 ^ new_n4169;
  assign new_n4227 = new_n4226 ^ new_n4180;
  assign new_n4228 = new_n4227 ^ new_n4225;
  assign new_n4229 = ~new_n4228 & new_n4158;
  assign new_n4230 = new_n4204 ^ new_n4194;
  assign new_n4231 = new_n4196 ^ new_n4191;
  assign new_n4232 = new_n4231 ^ new_n4230;
  assign new_n4233 = new_n4144 & new_n4232;
  assign new_n4234 = new_n4233 ^ new_n4229;
  assign new_n4235 = new_n4234 ^ new_n4217;
  assign new_n4236 = new_n4221 ^ new_n4164;
  assign new_n4237 = new_n4148 & new_n4236;
  assign new_n4238 = new_n4237 ^ new_n4235;
  assign new_n4239 = new_n4238 ^ new_n4216;
  assign new_n4240 = new_n4239 ^ new_n4210;
  assign new_n4241 = new_n4240 ^ new_n4130;
  assign new_n4242 = new_n4241 ^ new_n4021;
  assign new_n4243 = new_n4242 ^ new_n4012;
  assign new_n4244 = new_n4009 ^ new_n3992;
  assign new_n4245 = new_n3927 & new_n3967;
  assign new_n4246 = new_n3943 & new_n3962;
  assign new_n4247 = new_n4246 ^ new_n4245;
  assign new_n4248 = new_n4247 ^ new_n3987;
  assign new_n4249 = new_n4248 ^ new_n4244;
  assign new_n4250 = new_n4249 ^ new_n4020;
  assign new_n4251 = new_n4221 ^ new_n4194;
  assign new_n4252 = new_n4251 ^ new_n4184;
  assign new_n4253 = new_n4168 & new_n4252;
  assign new_n4254 = new_n4204 ^ new_n4141;
  assign new_n4255 = new_n4189 ^ new_n4154;
  assign new_n4256 = new_n4255 ^ new_n4224;
  assign new_n4257 = new_n4256 ^ new_n4254;
  assign new_n4258 = ~new_n4257 & new_n4160;
  assign new_n4259 = new_n4258 ^ new_n4253;
  assign new_n4260 = ~new_n4228 & new_n4157;
  assign new_n4261 = new_n4260 ^ new_n4237;
  assign new_n4262 = new_n4149 & new_n4236;
  assign new_n4263 = new_n4262 ^ new_n4199;
  assign new_n4264 = new_n4263 ^ new_n4234;
  assign new_n4265 = new_n4264 ^ new_n4261;
  assign new_n4266 = new_n4265 ^ new_n4259;
  assign new_n4267 = new_n4094 ^ new_n4032;
  assign new_n4268 = new_n4079 ^ new_n4045;
  assign new_n4269 = new_n4268 ^ new_n4116;
  assign new_n4270 = new_n4269 ^ new_n4267;
  assign new_n4271 = ~new_n4270 & new_n4051;
  assign new_n4272 = new_n4108 ^ new_n4084;
  assign new_n4273 = new_n4272 ^ new_n4074;
  assign new_n4274 = new_n4058 & new_n4273;
  assign new_n4275 = new_n4274 ^ new_n4271;
  assign new_n4276 = ~new_n4120 & new_n4049;
  assign new_n4277 = new_n4276 ^ new_n4110;
  assign new_n4278 = new_n4040 & new_n4109;
  assign new_n4279 = new_n4278 ^ new_n4089;
  assign new_n4280 = new_n4279 ^ new_n4126;
  assign new_n4281 = new_n4280 ^ new_n4277;
  assign new_n4282 = new_n4281 ^ new_n4275;
  assign new_n4283 = new_n4282 ^ new_n4266;
  assign new_n4284 = new_n4283 ^ new_n4250;
  assign new_n4285 = new_n3876 ^ new_n3869;
  assign new_n4286 = new_n3860 ^ new_n3845;
  assign new_n4287 = new_n3798 & new_n3859;
  assign new_n4288 = new_n4287 ^ new_n3880;
  assign new_n4289 = new_n4288 ^ new_n3857;
  assign new_n4290 = new_n4289 ^ new_n4286;
  assign new_n4291 = new_n4290 ^ new_n4285;
  assign new_n4292 = new_n4291 ^ new_n1183;
  assign new_n4293 = new_n3870 ^ new_n3848;
  assign new_n4294 = new_n4293 ^ new_n4289;
  assign new_n4295 = new_n4294 ^ new_n4292;
  assign new_n4296 = new_n4295 ^ new_n4284;
  assign new_n4297 = new_n4296 ^ new_n4243;
  assign new_n4298 = new_n4044 & new_n4104;
  assign new_n4299 = new_n4059 & new_n4273;
  assign new_n4300 = new_n4299 ^ new_n4128;
  assign new_n4301 = new_n4300 ^ new_n4276;
  assign new_n4302 = new_n4301 ^ new_n4298;
  assign new_n4303 = new_n4078 & new_n4088;
  assign new_n4304 = new_n4303 ^ new_n4271;
  assign new_n4305 = ~new_n4098 & new_n4036;
  assign new_n4306 = new_n4305 ^ new_n4105;
  assign new_n4307 = new_n4306 ^ new_n4274;
  assign new_n4308 = new_n4307 ^ new_n4304;
  assign new_n4309 = new_n4308 ^ new_n4302;
  assign new_n4310 = new_n4153 & new_n4214;
  assign new_n4311 = new_n4167 & new_n4252;
  assign new_n4312 = new_n4311 ^ new_n4238;
  assign new_n4313 = new_n4312 ^ new_n4260;
  assign new_n4314 = new_n4313 ^ new_n4310;
  assign new_n4315 = ~new_n4208 & new_n4145;
  assign new_n4316 = new_n4315 ^ new_n4215;
  assign new_n4317 = new_n4316 ^ new_n4253;
  assign new_n4318 = new_n4188 & new_n4198;
  assign new_n4319 = new_n4318 ^ new_n4258;
  assign new_n4320 = new_n4319 ^ new_n4317;
  assign new_n4321 = new_n4320 ^ new_n4314;
  assign new_n4322 = new_n4321 ^ new_n4309;
  assign new_n4323 = new_n4008 ^ new_n4002;
  assign new_n4324 = new_n3994 ^ new_n3968;
  assign new_n4325 = new_n4324 ^ new_n4248;
  assign new_n4326 = new_n4325 ^ new_n4323;
  assign new_n4327 = new_n4326 ^ new_n4322;
  assign new_n4328 = new_n3879 ^ new_n1202;
  assign new_n4329 = new_n4328 ^ new_n4291;
  assign new_n4330 = new_n4329 ^ new_n4327;
  assign new_n4331 = new_n4330 ^ new_n4297;
  assign new_n4332 = new_n4028 & new_n4124;
  assign new_n4333 = new_n4332 ^ new_n4276;
  assign new_n4334 = new_n4305 ^ new_n4103;
  assign new_n4335 = new_n4334 ^ new_n4099;
  assign new_n4336 = new_n4335 ^ new_n4127;
  assign new_n4337 = new_n4336 ^ new_n4333;
  assign new_n4338 = new_n4337 ^ new_n1119;
  assign new_n4339 = new_n4017 ^ new_n3855;
  assign new_n4340 = new_n3773 & new_n3875;
  assign new_n4341 = new_n4340 ^ new_n3878;
  assign new_n4342 = new_n4341 ^ new_n4339;
  assign new_n4343 = new_n4014 ^ new_n3986;
  assign new_n4344 = ~new_n4001 & new_n3907;
  assign new_n4345 = new_n4344 ^ new_n4010;
  assign new_n4346 = new_n4345 ^ new_n4343;
  assign new_n4347 = new_n4346 ^ new_n4342;
  assign new_n4348 = new_n4017 ^ new_n3845;
  assign new_n4349 = new_n3883 ^ new_n3867;
  assign new_n4350 = new_n4349 ^ new_n3881;
  assign new_n4351 = new_n4350 ^ new_n3858;
  assign new_n4352 = new_n4351 ^ new_n4348;
  assign new_n4353 = new_n4138 & new_n4232;
  assign new_n4354 = new_n4353 ^ new_n4260;
  assign new_n4355 = new_n4315 ^ new_n4213;
  assign new_n4356 = new_n4355 ^ new_n4209;
  assign new_n4357 = new_n4356 ^ new_n4235;
  assign new_n4358 = new_n4357 ^ new_n4354;
  assign new_n4359 = new_n4358 ^ new_n4352;
  assign new_n4360 = new_n4359 ^ new_n4347;
  assign new_n4361 = new_n4360 ^ new_n4338;
  assign new_n4362 = new_n4361 ^ new_n4331;
  assign new_n4363 = new_n4332 ^ new_n4099;
  assign new_n4364 = new_n4363 ^ new_n4301;
  assign new_n4365 = new_n4364 ^ new_n1191;
  assign new_n4366 = new_n4014 ^ new_n3994;
  assign new_n4367 = ~new_n3971 & new_n3926;
  assign new_n4368 = new_n4367 ^ new_n4005;
  assign new_n4369 = new_n4368 ^ new_n4013;
  assign new_n4370 = new_n4369 ^ new_n3988;
  assign new_n4371 = new_n4370 ^ new_n4366;
  assign new_n4372 = new_n4371 ^ new_n4352;
  assign new_n4373 = new_n4353 ^ new_n4209;
  assign new_n4374 = new_n4373 ^ new_n4313;
  assign new_n4375 = new_n4374 ^ new_n4019;
  assign new_n4376 = new_n4375 ^ new_n4372;
  assign new_n4377 = new_n4376 ^ new_n4365;
  assign new_n4378 = new_n4020 ^ new_n1164;
  assign new_n4379 = new_n4350 ^ new_n3862;
  assign new_n4380 = new_n4356 ^ new_n4312;
  assign new_n4381 = new_n4380 ^ new_n4379;
  assign new_n4382 = new_n4381 ^ new_n4378;
  assign new_n4383 = new_n4246 ^ new_n4013;
  assign new_n4384 = new_n4367 ^ new_n4006;
  assign new_n4385 = new_n4384 ^ new_n3989;
  assign new_n4386 = new_n4385 ^ new_n4383;
  assign new_n4387 = new_n4386 ^ new_n3886;
  assign new_n4388 = new_n4335 ^ new_n4300;
  assign new_n4389 = new_n4388 ^ new_n4387;
  assign new_n4390 = new_n4389 ^ new_n4382;
  assign new_n4391 = new_n4390 ^ new_n4377;
  assign new_n4392 = new_n4391 ^ new_n4297;
  assign new_n4393 = new_n4377 ^ new_n4296;
  assign new_n4394 = new_n4390 ^ new_n4330;
  assign new_n4395 = new_n4394 ^ new_n4393;
  assign new_n4396 = new_n4392 & new_n4395;
  assign new_n4397 = new_n4396 ^ new_n4361;
  assign new_n4398 = new_n4294 ^ new_n1155;
  assign new_n4399 = new_n4317 ^ new_n4311;
  assign new_n4400 = new_n4399 ^ new_n4264;
  assign new_n4401 = new_n4307 ^ new_n4299;
  assign new_n4402 = new_n4401 ^ new_n4280;
  assign new_n4403 = new_n4402 ^ new_n4400;
  assign new_n4404 = new_n4403 ^ new_n4020;
  assign new_n4405 = new_n4404 ^ new_n4398;
  assign new_n4406 = new_n4332 ^ new_n4125;
  assign new_n4407 = ~new_n4270 & new_n4041;
  assign new_n4408 = new_n4407 ^ new_n4308;
  assign new_n4409 = new_n4408 ^ new_n4406;
  assign new_n4410 = new_n4409 ^ new_n1142;
  assign new_n4411 = new_n4369 ^ new_n3993;
  assign new_n4412 = new_n4411 ^ new_n4379;
  assign new_n4413 = new_n4353 ^ new_n4233;
  assign new_n4414 = ~new_n4257 & new_n4150;
  assign new_n4415 = new_n4414 ^ new_n4320;
  assign new_n4416 = new_n4415 ^ new_n4413;
  assign new_n4417 = new_n4416 ^ new_n4342;
  assign new_n4418 = new_n4417 ^ new_n4412;
  assign new_n4419 = new_n4418 ^ new_n4410;
  assign new_n4420 = new_n4419 ^ new_n4361;
  assign new_n4421 = ~new_n4420 & new_n4405;
  assign new_n4422 = ~new_n4405 & new_n4390;
  assign new_n4423 = new_n4422 ^ new_n4421;
  assign new_n4424 = new_n4423 ^ new_n4397;
  assign new_n4425 = new_n4420 ^ new_n4405;
  assign new_n4426 = ~new_n4296 & ~new_n4425;
  assign new_n4427 = new_n4426 ^ new_n4296;
  assign new_n4428 = new_n4419 ^ new_n4331;
  assign new_n4429 = new_n4393 & new_n4428;
  assign new_n4430 = new_n4429 ^ new_n4427;
  assign new_n4431 = new_n4377 ^ new_n4330;
  assign new_n4432 = new_n4431 ^ new_n4430;
  assign new_n4433 = new_n4362 & new_n4391;
  assign new_n4434 = new_n4419 ^ new_n4390;
  assign new_n4435 = new_n4434 ^ new_n4431;
  assign new_n4436 = new_n4394 & new_n4435;
  assign new_n4437 = new_n4436 ^ new_n4433;
  assign new_n4438 = new_n4419 ^ new_n4243;
  assign new_n4439 = new_n4438 ^ new_n4437;
  assign new_n4440 = new_n4439 ^ new_n4432;
  assign new_n4441 = new_n4397 ^ new_n4392;
  assign new_n4442 = new_n4425 ^ new_n4296;
  assign new_n4443 = new_n4442 ^ new_n4431;
  assign new_n4444 = new_n4405 ^ new_n4392;
  assign new_n4445 = new_n4443 & new_n4444;
  assign new_n4446 = new_n4445 ^ new_n4433;
  assign new_n4447 = new_n4436 ^ new_n4330;
  assign new_n4448 = new_n4447 ^ new_n4446;
  assign new_n4449 = new_n4448 ^ new_n4441;
  assign new_n4450 = ~new_n4440 & new_n4449;
  assign new_n4451 = new_n4450 ^ new_n4424;
  assign new_n4452 = new_n4420 ^ new_n4392;
  assign new_n4453 = new_n4431 & new_n4452;
  assign new_n4454 = new_n4453 ^ new_n4433;
  assign new_n4455 = new_n4454 ^ new_n4428;
  assign new_n4456 = new_n4455 ^ new_n4451;
  assign new_n4457 = new_n4425 ^ new_n4377;
  assign new_n4458 = new_n4405 ^ new_n4362;
  assign new_n4459 = new_n4457 & new_n4458;
  assign new_n4460 = new_n4459 ^ new_n4426;
  assign new_n4461 = new_n4453 ^ new_n4436;
  assign new_n4462 = new_n4461 ^ new_n4460;
  assign new_n4463 = ~new_n4462 & new_n4456;
  assign new_n4464 = new_n4419 ^ new_n4377;
  assign new_n4465 = new_n4423 ^ new_n4390;
  assign new_n4466 = new_n4465 ^ new_n4445;
  assign new_n4467 = new_n4466 ^ new_n4461;
  assign new_n4468 = new_n4467 ^ new_n4464;
  assign new_n4469 = new_n4459 ^ new_n4429;
  assign new_n4470 = new_n4469 ^ new_n4377;
  assign new_n4471 = new_n4470 ^ new_n4455;
  assign new_n4472 = new_n4471 ^ new_n4450;
  assign new_n4473 = new_n4468 & new_n4472;
  assign new_n4474 = new_n4473 ^ new_n4463;
  assign new_n4475 = new_n4470 ^ new_n4424;
  assign new_n4476 = new_n4475 ^ new_n4474;
  assign new_n4477 = new_n4362 & new_n4476;
  assign new_n4478 = new_n4463 ^ new_n4450;
  assign new_n4479 = new_n4471 & new_n4478;
  assign new_n4480 = new_n4479 ^ new_n4440;
  assign new_n4481 = ~new_n4480 & new_n4395;
  assign new_n4482 = new_n4481 ^ new_n4477;
  assign new_n4483 = new_n4479 ^ new_n4463;
  assign new_n4484 = new_n4483 ^ new_n4462;
  assign new_n4485 = ~new_n4484 & new_n4443;
  assign new_n4486 = new_n4391 & new_n4476;
  assign new_n4487 = new_n4419 ^ new_n4296;
  assign new_n4488 = new_n4445 ^ new_n4427;
  assign new_n4489 = new_n4473 ^ new_n4424;
  assign new_n4490 = new_n4489 ^ new_n4455;
  assign new_n4491 = new_n4479 ^ new_n4472;
  assign new_n4492 = new_n4490 & new_n4491;
  assign new_n4493 = new_n4492 ^ new_n4479;
  assign new_n4494 = new_n4493 ^ new_n4488;
  assign new_n4495 = new_n4494 ^ new_n4487;
  assign new_n4496 = new_n4495 ^ new_n4390;
  assign new_n4497 = new_n4473 ^ new_n4429;
  assign new_n4498 = new_n4497 ^ new_n4397;
  assign new_n4499 = new_n4498 ^ new_n4496;
  assign new_n4500 = ~new_n4499 & new_n4394;
  assign new_n4501 = new_n4500 ^ new_n4486;
  assign new_n4502 = new_n4501 ^ new_n4485;
  assign new_n4503 = new_n4492 ^ new_n4468;
  assign new_n4504 = new_n4425 & new_n4503;
  assign new_n4505 = new_n4504 ^ new_n4502;
  assign new_n4506 = new_n4492 ^ new_n4473;
  assign new_n4507 = new_n4506 ^ new_n4449;
  assign new_n4508 = new_n4428 & new_n4507;
  assign new_n4509 = new_n4508 ^ new_n4505;
  assign new_n4510 = ~new_n4499 & new_n4435;
  assign new_n4511 = new_n4510 ^ new_n4509;
  assign new_n4512 = new_n4511 ^ new_n4482;
  assign new_n4513 = new_n4512 ^ new_n3755;
  assign new_n4514 = new_n4513 ^ new_n2931;
  assign new_n4515 = ~new_n4484 & new_n4444;
  assign new_n4516 = ~new_n4480 & new_n4392;
  assign new_n4517 = new_n4516 ^ new_n4515;
  assign new_n4518 = new_n4517 ^ new_n4481;
  assign new_n4519 = new_n4518 ^ new_n4509;
  assign new_n4520 = new_n4458 & new_n4490;
  assign new_n4521 = new_n4520 ^ new_n4481;
  assign new_n4522 = new_n4471 ^ new_n4463;
  assign new_n4523 = new_n4405 & new_n4522;
  assign new_n4524 = new_n4523 ^ new_n4515;
  assign new_n4525 = new_n4524 ^ new_n4505;
  assign new_n4526 = new_n4525 ^ new_n4521;
  assign new_n4527 = new_n4526 ^ new_n4519;
  assign new_n4528 = ~new_n3672 & new_n3727;
  assign new_n4529 = new_n4528 ^ new_n3713;
  assign new_n4530 = ~new_n3695 & ~new_n3736;
  assign new_n4531 = new_n3709 ^ new_n3676;
  assign new_n4532 = ~new_n3669 & new_n4531;
  assign new_n4533 = new_n4532 ^ new_n4530;
  assign new_n4534 = new_n4533 ^ new_n3751;
  assign new_n4535 = new_n4534 ^ new_n4529;
  assign new_n4536 = new_n4535 ^ new_n4527;
  assign new_n4537 = new_n4536 ^ new_n4514;
  assign new_n4538 = new_n2050 & new_n2151;
  assign new_n4539 = new_n4538 ^ new_n2152;
  assign new_n4540 = new_n2124 ^ new_n1999;
  assign new_n4541 = new_n2091 ^ new_n2086;
  assign new_n4542 = new_n4541 ^ new_n2157;
  assign new_n4543 = new_n4542 ^ new_n4540;
  assign new_n4544 = ~new_n4543 & new_n2052;
  assign new_n4545 = new_n2084 & new_n2142;
  assign new_n4546 = ~new_n4543 & new_n2068;
  assign new_n4547 = new_n4546 ^ new_n4545;
  assign new_n4548 = new_n2124 ^ new_n2089;
  assign new_n4549 = new_n2082 & new_n4548;
  assign new_n4550 = new_n4549 ^ new_n2128;
  assign new_n4551 = new_n2073 & new_n2146;
  assign new_n4552 = new_n4551 ^ new_n4550;
  assign new_n4553 = new_n4552 ^ new_n4547;
  assign new_n4554 = new_n4553 ^ new_n4544;
  assign new_n4555 = new_n4554 ^ new_n4539;
  assign new_n4556 = new_n2811 & new_n2911;
  assign new_n4557 = new_n4556 ^ new_n2912;
  assign new_n4558 = new_n2884 ^ new_n2761;
  assign new_n4559 = new_n2852 ^ new_n2847;
  assign new_n4560 = new_n4559 ^ new_n2917;
  assign new_n4561 = new_n4560 ^ new_n4558;
  assign new_n4562 = ~new_n4561 & new_n2813;
  assign new_n4563 = new_n2845 & new_n2902;
  assign new_n4564 = ~new_n4561 & new_n2829;
  assign new_n4565 = new_n4564 ^ new_n4563;
  assign new_n4566 = new_n2884 ^ new_n2850;
  assign new_n4567 = new_n2843 & new_n4566;
  assign new_n4568 = new_n4567 ^ new_n2888;
  assign new_n4569 = new_n2834 & new_n2906;
  assign new_n4570 = new_n4569 ^ new_n4568;
  assign new_n4571 = new_n4570 ^ new_n4565;
  assign new_n4572 = new_n4571 ^ new_n4562;
  assign new_n4573 = new_n4572 ^ new_n4557;
  assign new_n4574 = new_n4573 ^ new_n4555;
  assign new_n4575 = new_n4486 ^ new_n4477;
  assign new_n4576 = new_n4463 ^ new_n4377;
  assign new_n4577 = new_n4465 ^ new_n4459;
  assign new_n4578 = new_n4577 ^ new_n4495;
  assign new_n4579 = new_n4578 ^ new_n4576;
  assign new_n4580 = ~new_n4579 & new_n4431;
  assign new_n4581 = new_n4393 & new_n4507;
  assign new_n4582 = new_n4523 ^ new_n4516;
  assign new_n4583 = new_n4582 ^ new_n4581;
  assign new_n4584 = ~new_n4579 & new_n4452;
  assign new_n4585 = new_n4457 & new_n4490;
  assign new_n4586 = new_n4585 ^ new_n4584;
  assign new_n4587 = new_n4586 ^ new_n4583;
  assign new_n4588 = new_n4587 ^ new_n4580;
  assign new_n4589 = new_n4588 ^ new_n4575;
  assign new_n4590 = new_n4589 ^ new_n4574;
  assign new_n4591 = ~new_n3712 & new_n3650;
  assign new_n4592 = new_n4591 ^ new_n4530;
  assign new_n4593 = new_n4592 ^ new_n3713;
  assign new_n4594 = new_n4593 ^ new_n3752;
  assign new_n4595 = new_n4594 ^ new_n4519;
  assign new_n4596 = ~new_n1270 & new_n1231;
  assign new_n4597 = new_n4596 ^ new_n1271;
  assign new_n4598 = ~new_n1244 & ~new_n1253;
  assign new_n4599 = new_n1258 ^ new_n1191;
  assign new_n4600 = new_n1246 ^ new_n1166;
  assign new_n4601 = new_n4600 ^ new_n1276;
  assign new_n4602 = new_n4601 ^ new_n4599;
  assign new_n4603 = ~new_n1213 & new_n4602;
  assign new_n4604 = new_n4603 ^ new_n4598;
  assign new_n4605 = new_n1258 ^ new_n1249;
  assign new_n4606 = ~new_n1155 & new_n4605;
  assign new_n4607 = new_n4606 ^ new_n1290;
  assign new_n4608 = ~new_n1227 & new_n1286;
  assign new_n4609 = new_n4608 ^ new_n4607;
  assign new_n4610 = new_n4609 ^ new_n4604;
  assign new_n4611 = new_n1203 & new_n4602;
  assign new_n4612 = new_n4611 ^ new_n4610;
  assign new_n4613 = new_n4612 ^ new_n4597;
  assign new_n4614 = new_n4613 ^ new_n3643;
  assign new_n4615 = new_n4614 ^ n123;
  assign new_n4616 = new_n4615 ^ n59;
  assign new_n4617 = new_n4616 ^ new_n4595;
  assign new_n4618 = new_n4617 ^ new_n4590;
  assign new_n4619 = ~new_n2921 & new_n2864;
  assign new_n4620 = new_n4619 ^ new_n4556;
  assign new_n4621 = new_n2924 ^ new_n2894;
  assign new_n4622 = new_n4621 ^ new_n4620;
  assign new_n4623 = ~new_n2161 & new_n2104;
  assign new_n4624 = new_n4623 ^ new_n4538;
  assign new_n4625 = new_n2164 ^ new_n2134;
  assign new_n4626 = new_n4625 ^ new_n4624;
  assign new_n4627 = new_n4626 ^ new_n4622;
  assign new_n4628 = new_n4627 ^ new_n4589;
  assign new_n4629 = ~new_n1211 & ~new_n1280;
  assign new_n4630 = new_n4629 ^ new_n4596;
  assign new_n4631 = new_n1294 ^ new_n1283;
  assign new_n4632 = new_n4631 ^ new_n4630;
  assign new_n4633 = new_n4632 ^ new_n3619;
  assign new_n4634 = new_n4633 ^ n58;
  assign new_n4635 = new_n3738 ^ new_n3724;
  assign new_n4636 = new_n3709 ^ new_n3483;
  assign new_n4637 = new_n3715 ^ new_n3673;
  assign new_n4638 = new_n4637 ^ new_n3743;
  assign new_n4639 = new_n4638 ^ new_n4636;
  assign new_n4640 = ~new_n4639 & new_n3627;
  assign new_n4641 = new_n4591 ^ new_n4532;
  assign new_n4642 = new_n3484 & new_n3731;
  assign new_n4643 = new_n4642 ^ new_n4641;
  assign new_n4644 = ~new_n3671 & new_n3727;
  assign new_n4645 = ~new_n4639 & new_n3651;
  assign new_n4646 = new_n4645 ^ new_n4644;
  assign new_n4647 = new_n4646 ^ new_n4643;
  assign new_n4648 = new_n4647 ^ new_n4640;
  assign new_n4649 = new_n4648 ^ new_n4635;
  assign new_n4650 = new_n4649 ^ new_n4634;
  assign new_n4651 = new_n4510 ^ new_n4477;
  assign new_n4652 = new_n4518 ^ new_n4502;
  assign new_n4653 = new_n4652 ^ new_n4651;
  assign new_n4654 = new_n4653 ^ new_n4650;
  assign new_n4655 = new_n4654 ^ new_n4628;
  assign new_n4656 = new_n4655 ^ new_n4618;
  assign new_n4657 = new_n4609 ^ new_n1287;
  assign new_n4658 = ~new_n1263 & new_n1217;
  assign new_n4659 = ~new_n1245 & ~new_n1253;
  assign new_n4660 = new_n4659 ^ new_n4658;
  assign new_n4661 = new_n4660 ^ new_n1282;
  assign new_n4662 = new_n4661 ^ new_n4657;
  assign new_n4663 = new_n4662 ^ new_n3659;
  assign new_n4664 = new_n4663 ^ n64;
  assign new_n4665 = new_n4583 ^ new_n4508;
  assign new_n4666 = new_n4442 & new_n4503;
  assign new_n4667 = new_n4666 ^ new_n4520;
  assign new_n4668 = new_n4667 ^ new_n4501;
  assign new_n4669 = new_n4668 ^ new_n4665;
  assign new_n4670 = new_n4669 ^ new_n4664;
  assign new_n4671 = new_n4570 ^ new_n2907;
  assign new_n4672 = new_n2872 & new_n2925;
  assign new_n4673 = new_n2846 & new_n2902;
  assign new_n4674 = new_n4673 ^ new_n4672;
  assign new_n4675 = new_n4674 ^ new_n2923;
  assign new_n4676 = new_n4675 ^ new_n4671;
  assign new_n4677 = new_n4552 ^ new_n2147;
  assign new_n4678 = new_n2112 & new_n2165;
  assign new_n4679 = new_n2085 & new_n2142;
  assign new_n4680 = new_n4679 ^ new_n4678;
  assign new_n4681 = new_n4680 ^ new_n2163;
  assign new_n4682 = new_n4681 ^ new_n4677;
  assign new_n4683 = new_n4682 ^ new_n4676;
  assign new_n4684 = new_n4683 ^ new_n4513;
  assign new_n4685 = new_n4684 ^ new_n4670;
  assign new_n4686 = new_n4685 ^ new_n4656;
  assign new_n4687 = new_n4686 ^ new_n4537;
  assign new_n4688 = new_n4569 ^ new_n4564;
  assign new_n4689 = new_n4619 ^ new_n2926;
  assign new_n4690 = new_n4689 ^ new_n4675;
  assign new_n4691 = new_n4690 ^ new_n4688;
  assign new_n4692 = new_n4551 ^ new_n4546;
  assign new_n4693 = new_n4623 ^ new_n2166;
  assign new_n4694 = new_n4693 ^ new_n4681;
  assign new_n4695 = new_n4694 ^ new_n4692;
  assign new_n4696 = new_n4695 ^ new_n4691;
  assign new_n4697 = new_n4696 ^ new_n4669;
  assign new_n4698 = new_n4697 ^ new_n4513;
  assign new_n4699 = new_n4608 ^ new_n4603;
  assign new_n4700 = new_n4629 ^ new_n1264;
  assign new_n4701 = new_n4700 ^ new_n4661;
  assign new_n4702 = new_n4701 ^ new_n4699;
  assign new_n4703 = new_n4702 ^ new_n3419;
  assign new_n4704 = new_n4703 ^ n63;
  assign new_n4705 = new_n4643 ^ new_n3732;
  assign new_n4706 = ~new_n3696 & new_n3733;
  assign new_n4707 = new_n4706 ^ new_n4528;
  assign new_n4708 = new_n4707 ^ new_n3749;
  assign new_n4709 = new_n4708 ^ new_n4705;
  assign new_n4710 = new_n4709 ^ new_n4704;
  assign new_n4711 = new_n4584 ^ new_n4581;
  assign new_n4712 = new_n4510 ^ new_n4504;
  assign new_n4713 = new_n4712 ^ new_n4668;
  assign new_n4714 = new_n4713 ^ new_n4711;
  assign new_n4715 = new_n4714 ^ new_n4710;
  assign new_n4716 = new_n4715 ^ new_n4698;
  assign new_n4717 = ~new_n4686 & ~new_n4716;
  assign new_n4718 = new_n4717 ^ new_n4716;
  assign new_n4719 = new_n4556 ^ new_n2893;
  assign new_n4720 = new_n4619 ^ new_n2928;
  assign new_n4721 = new_n4720 ^ new_n4719;
  assign new_n4722 = new_n4538 ^ new_n2133;
  assign new_n4723 = new_n4623 ^ new_n2168;
  assign new_n4724 = new_n4723 ^ new_n4722;
  assign new_n4725 = new_n4724 ^ new_n4721;
  assign new_n4726 = new_n4725 ^ new_n4653;
  assign new_n4727 = new_n4596 ^ new_n1293;
  assign new_n4728 = new_n4629 ^ new_n1288;
  assign new_n4729 = new_n4728 ^ new_n4727;
  assign new_n4730 = new_n4729 ^ new_n3471;
  assign new_n4731 = new_n4730 ^ n121;
  assign new_n4732 = new_n4731 ^ n57;
  assign new_n4733 = new_n4732 ^ new_n4512;
  assign new_n4734 = new_n3753 ^ new_n3724;
  assign new_n4735 = new_n4593 ^ new_n3750;
  assign new_n4736 = new_n4735 ^ new_n4734;
  assign new_n4737 = new_n4736 ^ new_n4733;
  assign new_n4738 = new_n4737 ^ new_n4726;
  assign new_n4739 = new_n4738 ^ new_n4716;
  assign new_n4740 = new_n2090 & new_n4548;
  assign new_n4741 = new_n4740 ^ new_n4723;
  assign new_n4742 = new_n4741 ^ new_n4553;
  assign new_n4743 = new_n2851 & new_n4566;
  assign new_n4744 = new_n4743 ^ new_n4720;
  assign new_n4745 = new_n4744 ^ new_n4571;
  assign new_n4746 = new_n4745 ^ new_n4742;
  assign new_n4747 = new_n4746 ^ new_n4714;
  assign new_n4748 = ~new_n1165 & new_n4605;
  assign new_n4749 = new_n4748 ^ new_n4728;
  assign new_n4750 = new_n4749 ^ new_n4610;
  assign new_n4751 = new_n4750 ^ new_n3526;
  assign new_n4752 = new_n4751 ^ n126;
  assign new_n4753 = new_n4752 ^ n62;
  assign new_n4754 = new_n4425 ^ new_n4390;
  assign new_n4755 = new_n4522 & new_n4754;
  assign new_n4756 = new_n4755 ^ new_n4511;
  assign new_n4757 = new_n4756 ^ new_n4587;
  assign new_n4758 = new_n4757 ^ new_n4753;
  assign new_n4759 = new_n4645 ^ new_n4642;
  assign new_n4760 = new_n3753 ^ new_n3734;
  assign new_n4761 = new_n4760 ^ new_n4708;
  assign new_n4762 = new_n4761 ^ new_n4759;
  assign new_n4763 = new_n4762 ^ new_n4758;
  assign new_n4764 = new_n4763 ^ new_n4747;
  assign new_n4765 = new_n4757 ^ new_n4526;
  assign new_n4766 = new_n3670 ^ new_n3567;
  assign new_n4767 = ~new_n4766 & new_n4531;
  assign new_n4768 = new_n4767 ^ new_n3754;
  assign new_n4769 = new_n4768 ^ new_n4647;
  assign new_n4770 = new_n4769 ^ new_n4765;
  assign new_n4771 = new_n4659 ^ new_n1293;
  assign new_n4772 = new_n4606 ^ new_n1291;
  assign new_n4773 = new_n4772 ^ new_n1284;
  assign new_n4774 = new_n4773 ^ new_n4771;
  assign new_n4775 = new_n4774 ^ new_n3591;
  assign new_n4776 = new_n4775 ^ n125;
  assign new_n4777 = new_n4776 ^ n61;
  assign new_n4778 = new_n4673 ^ new_n2893;
  assign new_n4779 = new_n4567 ^ new_n2891;
  assign new_n4780 = new_n4779 ^ new_n2927;
  assign new_n4781 = new_n4780 ^ new_n4778;
  assign new_n4782 = new_n4679 ^ new_n2133;
  assign new_n4783 = new_n4549 ^ new_n2131;
  assign new_n4784 = new_n4783 ^ new_n2167;
  assign new_n4785 = new_n4784 ^ new_n4782;
  assign new_n4786 = new_n4785 ^ new_n4781;
  assign new_n4787 = new_n4786 ^ new_n4777;
  assign new_n4788 = new_n4787 ^ new_n4513;
  assign new_n4789 = new_n4788 ^ new_n4770;
  assign new_n4790 = new_n4789 ^ new_n4716;
  assign new_n4791 = new_n4790 ^ new_n4764;
  assign new_n4792 = new_n4791 ^ new_n4618;
  assign new_n4793 = ~new_n4792 & new_n4739;
  assign new_n4794 = new_n4793 ^ new_n4718;
  assign new_n4795 = new_n4764 ^ new_n4738;
  assign new_n4796 = new_n4795 ^ new_n4794;
  assign new_n4797 = new_n4791 ^ new_n4655;
  assign new_n4798 = new_n4738 ^ new_n4537;
  assign new_n4799 = ~new_n4797 & new_n4798;
  assign new_n4800 = new_n4618 ^ new_n4537;
  assign new_n4801 = new_n4800 ^ new_n4795;
  assign new_n4802 = new_n4764 ^ new_n4537;
  assign new_n4803 = ~new_n4801 & new_n4802;
  assign new_n4804 = new_n4803 ^ new_n4799;
  assign new_n4805 = new_n4789 ^ new_n4618;
  assign new_n4806 = new_n4805 ^ new_n4804;
  assign new_n4807 = new_n4806 ^ new_n4796;
  assign new_n4808 = new_n4798 ^ new_n4790;
  assign new_n4809 = new_n4716 ^ new_n4537;
  assign new_n4810 = new_n4809 ^ new_n4795;
  assign new_n4811 = new_n4808 & new_n4810;
  assign new_n4812 = new_n4811 ^ new_n4655;
  assign new_n4813 = new_n4812 ^ new_n4808;
  assign new_n4814 = new_n4808 ^ new_n4685;
  assign new_n4815 = new_n4716 ^ new_n4686;
  assign new_n4816 = new_n4815 ^ new_n4795;
  assign new_n4817 = new_n4814 & new_n4816;
  assign new_n4818 = new_n4817 ^ new_n4804;
  assign new_n4819 = new_n4818 ^ new_n4764;
  assign new_n4820 = new_n4819 ^ new_n4813;
  assign new_n4821 = ~new_n4820 & new_n4807;
  assign new_n4822 = new_n4685 & new_n4687;
  assign new_n4823 = new_n4822 ^ new_n4537;
  assign new_n4824 = new_n4823 ^ new_n4812;
  assign new_n4825 = new_n4824 ^ new_n4821;
  assign new_n4826 = new_n4808 ^ new_n4656;
  assign new_n4827 = new_n4795 & new_n4826;
  assign new_n4828 = new_n4827 ^ new_n4799;
  assign new_n4829 = new_n4828 ^ new_n4792;
  assign new_n4830 = new_n4829 ^ new_n4825;
  assign new_n4831 = new_n4738 ^ new_n4686;
  assign new_n4832 = new_n4797 ^ new_n4685;
  assign new_n4833 = ~new_n4832 & new_n4831;
  assign new_n4834 = new_n4833 ^ new_n4717;
  assign new_n4835 = new_n4827 ^ new_n4803;
  assign new_n4836 = new_n4835 ^ new_n4834;
  assign new_n4837 = ~new_n4836 & new_n4830;
  assign new_n4838 = new_n4833 ^ new_n4793;
  assign new_n4839 = new_n4838 ^ new_n4738;
  assign new_n4840 = new_n4839 ^ new_n4829;
  assign new_n4841 = new_n4840 ^ new_n4837;
  assign new_n4842 = ~new_n4841 & new_n4687;
  assign new_n4843 = new_n4716 ^ new_n4618;
  assign new_n4844 = new_n4817 ^ new_n4718;
  assign new_n4845 = new_n4738 ^ new_n4618;
  assign new_n4846 = new_n4822 ^ new_n4817;
  assign new_n4847 = new_n4846 ^ new_n4835;
  assign new_n4848 = new_n4847 ^ new_n4845;
  assign new_n4849 = new_n4840 ^ new_n4821;
  assign new_n4850 = ~new_n4848 & ~new_n4849;
  assign new_n4851 = new_n4850 ^ new_n4824;
  assign new_n4852 = new_n4851 ^ new_n4829;
  assign new_n4853 = new_n4837 ^ new_n4821;
  assign new_n4854 = ~new_n4840 & ~new_n4853;
  assign new_n4855 = new_n4854 ^ new_n4821;
  assign new_n4856 = new_n4852 & new_n4855;
  assign new_n4857 = new_n4854 ^ new_n4840;
  assign new_n4858 = new_n4857 ^ new_n4856;
  assign new_n4859 = new_n4858 ^ new_n4844;
  assign new_n4860 = new_n4859 ^ new_n4843;
  assign new_n4861 = new_n4860 ^ new_n4537;
  assign new_n4862 = new_n4850 ^ new_n4793;
  assign new_n4863 = new_n4862 ^ new_n4812;
  assign new_n4864 = new_n4863 ^ new_n4861;
  assign new_n4865 = ~new_n4801 & new_n4864;
  assign new_n4866 = new_n4856 ^ new_n4848;
  assign new_n4867 = ~new_n4866 & new_n4686;
  assign new_n4868 = new_n4802 & new_n4864;
  assign new_n4869 = new_n4850 ^ new_n4837;
  assign new_n4870 = new_n4839 ^ new_n4824;
  assign new_n4871 = new_n4870 ^ new_n4869;
  assign new_n4872 = ~new_n4871 & new_n4798;
  assign new_n4873 = new_n4872 ^ new_n4868;
  assign new_n4874 = new_n4857 ^ new_n4837;
  assign new_n4875 = new_n4874 ^ new_n4836;
  assign new_n4876 = new_n4816 & new_n4875;
  assign new_n4877 = new_n4876 ^ new_n4873;
  assign new_n4878 = new_n4877 ^ new_n4867;
  assign new_n4879 = new_n4856 ^ new_n4850;
  assign new_n4880 = new_n4879 ^ new_n4820;
  assign new_n4881 = ~new_n4792 & ~new_n4880;
  assign new_n4882 = new_n4881 ^ new_n4878;
  assign new_n4883 = new_n4882 ^ new_n4865;
  assign new_n4884 = new_n4883 ^ new_n4842;
  assign new_n4885 = new_n4831 & new_n4852;
  assign new_n4886 = new_n4837 ^ new_n4738;
  assign new_n4887 = new_n4833 ^ new_n4822;
  assign new_n4888 = new_n4887 ^ new_n4860;
  assign new_n4889 = new_n4888 ^ new_n4886;
  assign new_n4890 = ~new_n4889 & new_n4826;
  assign new_n4891 = new_n4890 ^ new_n4885;
  assign new_n4892 = new_n4857 ^ new_n4807;
  assign new_n4893 = ~new_n4892 & new_n4808;
  assign new_n4894 = ~new_n4841 & new_n4685;
  assign new_n4895 = new_n4894 ^ new_n4893;
  assign new_n4896 = ~new_n4880 & new_n4739;
  assign new_n4897 = new_n4896 ^ new_n4895;
  assign new_n4898 = new_n4897 ^ new_n4891;
  assign new_n4899 = new_n4898 ^ new_n4884;
  assign new_n4900 = new_n4899 ^ new_n1013;
  assign new_n4901 = new_n818 ^ new_n565;
  assign new_n4902 = new_n2759 ^ new_n1117;
  assign new_n4903 = new_n2794 ^ new_n2754;
  assign new_n4904 = new_n4903 ^ new_n2822;
  assign new_n4905 = new_n4904 ^ new_n4902;
  assign new_n4906 = new_n2680 ^ new_n1200;
  assign new_n4907 = new_n2772 ^ new_n2668;
  assign new_n4908 = new_n4907 ^ new_n2396;
  assign new_n4909 = new_n4908 ^ new_n4906;
  assign new_n4910 = new_n2786 ^ new_n2282;
  assign new_n4911 = new_n4910 ^ new_n2841;
  assign new_n4912 = new_n2647 ^ new_n1181;
  assign new_n4913 = new_n4912 ^ new_n2749;
  assign new_n4914 = new_n4913 ^ new_n4911;
  assign new_n4915 = new_n2673 ^ new_n1173;
  assign new_n4916 = new_n4915 ^ new_n2749;
  assign new_n4917 = new_n2734 ^ new_n2695;
  assign new_n4918 = new_n4917 ^ new_n2782;
  assign new_n4919 = new_n4918 ^ new_n4916;
  assign new_n4920 = new_n4919 ^ new_n4914;
  assign new_n4921 = new_n4920 ^ new_n4909;
  assign new_n4922 = new_n4921 ^ new_n4905;
  assign new_n4923 = new_n2808 ^ new_n1140;
  assign new_n4924 = new_n2817 ^ new_n2802;
  assign new_n4925 = new_n4924 ^ new_n2727;
  assign new_n4926 = new_n4925 ^ new_n4923;
  assign new_n4927 = new_n2618 ^ new_n1189;
  assign new_n4928 = new_n2744 ^ new_n2507;
  assign new_n4929 = new_n4928 ^ new_n2798;
  assign new_n4930 = new_n4929 ^ new_n4927;
  assign new_n4931 = new_n4930 ^ new_n4926;
  assign new_n4932 = new_n2655 ^ new_n1153;
  assign new_n4933 = new_n2840 ^ new_n2631;
  assign new_n4934 = new_n4933 ^ new_n2749;
  assign new_n4935 = new_n4934 ^ new_n4932;
  assign new_n4936 = new_n2824 ^ new_n2720;
  assign new_n4937 = new_n4936 ^ new_n2710;
  assign new_n4938 = new_n2737 ^ new_n1162;
  assign new_n4939 = new_n4938 ^ new_n2749;
  assign new_n4940 = new_n4939 ^ new_n4937;
  assign new_n4941 = new_n4940 ^ new_n4930;
  assign new_n4942 = new_n4941 ^ new_n4920;
  assign new_n4943 = new_n4942 ^ new_n4935;
  assign new_n4944 = new_n4926 ^ new_n4905;
  assign new_n4945 = new_n4944 ^ new_n4935;
  assign new_n4946 = new_n4945 ^ new_n4914;
  assign new_n4947 = new_n4930 ^ new_n4909;
  assign new_n4948 = new_n4947 ^ new_n4946;
  assign new_n4949 = new_n4943 & new_n4948;
  assign new_n4950 = new_n4945 ^ new_n4940;
  assign new_n4951 = new_n4935 & new_n4950;
  assign new_n4952 = new_n4951 ^ new_n4949;
  assign new_n4953 = new_n4940 ^ new_n4926;
  assign new_n4954 = new_n4953 ^ new_n4947;
  assign new_n4955 = new_n4940 ^ new_n4909;
  assign new_n4956 = new_n4954 & new_n4955;
  assign new_n4957 = new_n4944 ^ new_n4942;
  assign new_n4958 = new_n4947 & new_n4957;
  assign new_n4959 = new_n4958 ^ new_n4956;
  assign new_n4960 = new_n4959 ^ new_n4952;
  assign new_n4961 = new_n4960 ^ new_n4931;
  assign new_n4962 = ~new_n4914 & ~new_n4945;
  assign new_n4963 = new_n4962 ^ new_n4914;
  assign new_n4964 = new_n4926 ^ new_n4921;
  assign new_n4965 = new_n4930 ^ new_n4914;
  assign new_n4966 = new_n4964 & new_n4965;
  assign new_n4967 = new_n4966 ^ new_n4963;
  assign new_n4968 = new_n4967 ^ new_n4947;
  assign new_n4969 = new_n4922 & new_n4941;
  assign new_n4970 = new_n4969 ^ new_n4956;
  assign new_n4971 = new_n4926 ^ new_n4919;
  assign new_n4972 = new_n4971 ^ new_n4970;
  assign new_n4973 = new_n4972 ^ new_n4968;
  assign new_n4974 = new_n4940 ^ new_n4914;
  assign new_n4975 = new_n4974 ^ new_n4947;
  assign new_n4976 = new_n4942 & new_n4975;
  assign new_n4977 = new_n4976 ^ new_n4905;
  assign new_n4978 = new_n4977 ^ new_n4942;
  assign new_n4979 = new_n4969 ^ new_n4949;
  assign new_n4980 = new_n4956 ^ new_n4909;
  assign new_n4981 = new_n4980 ^ new_n4979;
  assign new_n4982 = new_n4981 ^ new_n4978;
  assign new_n4983 = ~new_n4973 & new_n4982;
  assign new_n4984 = new_n4945 ^ new_n4930;
  assign new_n4985 = new_n4935 ^ new_n4922;
  assign new_n4986 = new_n4984 & new_n4985;
  assign new_n4987 = new_n4986 ^ new_n4966;
  assign new_n4988 = new_n4987 ^ new_n4930;
  assign new_n4989 = new_n4969 ^ new_n4958;
  assign new_n4990 = new_n4989 ^ new_n4964;
  assign new_n4991 = new_n4990 ^ new_n4988;
  assign new_n4992 = new_n4991 ^ new_n4983;
  assign new_n4993 = new_n4961 & new_n4992;
  assign new_n4994 = new_n4951 ^ new_n4940;
  assign new_n4995 = new_n4994 ^ new_n4977;
  assign new_n4996 = new_n4995 ^ new_n4983;
  assign new_n4997 = new_n4996 ^ new_n4990;
  assign new_n4998 = new_n4986 ^ new_n4962;
  assign new_n4999 = new_n4998 ^ new_n4959;
  assign new_n5000 = ~new_n4999 & new_n4997;
  assign new_n5001 = new_n5000 ^ new_n4993;
  assign new_n5002 = new_n4995 ^ new_n4988;
  assign new_n5003 = new_n5002 ^ new_n5001;
  assign new_n5004 = new_n4922 & new_n5003;
  assign new_n5005 = new_n4926 ^ new_n4914;
  assign new_n5006 = new_n4963 ^ new_n4949;
  assign new_n5007 = new_n4995 ^ new_n4993;
  assign new_n5008 = new_n5007 ^ new_n4990;
  assign new_n5009 = new_n5000 ^ new_n4983;
  assign new_n5010 = ~new_n5009 & new_n4991;
  assign new_n5011 = new_n5010 ^ new_n4983;
  assign new_n5012 = new_n5008 & new_n5011;
  assign new_n5013 = new_n5010 ^ new_n4991;
  assign new_n5014 = new_n5013 ^ new_n5012;
  assign new_n5015 = new_n5014 ^ new_n5006;
  assign new_n5016 = new_n5015 ^ new_n5005;
  assign new_n5017 = new_n5016 ^ new_n4940;
  assign new_n5018 = new_n4993 ^ new_n4966;
  assign new_n5019 = new_n5018 ^ new_n4977;
  assign new_n5020 = new_n5019 ^ new_n5017;
  assign new_n5021 = ~new_n5020 & new_n4954;
  assign new_n5022 = new_n5021 ^ new_n5004;
  assign new_n5023 = new_n5013 ^ new_n5000;
  assign new_n5024 = new_n5023 ^ new_n4999;
  assign new_n5025 = ~new_n5024 & new_n4943;
  assign new_n5026 = new_n5013 ^ new_n4973;
  assign new_n5027 = ~new_n5026 & new_n4942;
  assign new_n5028 = new_n5027 ^ new_n5025;
  assign new_n5029 = ~new_n5026 & new_n4975;
  assign new_n5030 = new_n5029 ^ new_n5028;
  assign new_n5031 = ~new_n5024 & new_n4948;
  assign new_n5032 = new_n4941 & new_n5003;
  assign new_n5033 = ~new_n5020 & new_n4955;
  assign new_n5034 = new_n5033 ^ new_n5032;
  assign new_n5035 = new_n5034 ^ new_n5031;
  assign new_n5036 = new_n5035 ^ new_n5030;
  assign new_n5037 = new_n5036 ^ new_n5022;
  assign new_n5038 = new_n5037 ^ new_n4901;
  assign new_n5039 = new_n3606 ^ new_n875;
  assign new_n5040 = new_n3446 ^ new_n3376;
  assign new_n5041 = new_n5040 ^ new_n3389;
  assign new_n5042 = new_n5041 ^ new_n5039;
  assign new_n5043 = new_n3460 ^ new_n865;
  assign new_n5044 = new_n5043 ^ new_n3587;
  assign new_n5045 = new_n3638 ^ new_n3545;
  assign new_n5046 = new_n5045 ^ new_n3560;
  assign new_n5047 = new_n5046 ^ new_n5044;
  assign new_n5048 = new_n5047 ^ new_n5042;
  assign new_n5049 = new_n3515 ^ new_n3495;
  assign new_n5050 = new_n5049 ^ new_n3577;
  assign new_n5051 = new_n3154 ^ new_n903;
  assign new_n5052 = new_n5051 ^ new_n5050;
  assign new_n5053 = new_n5052 ^ new_n5042;
  assign new_n5054 = new_n3582 ^ new_n3559;
  assign new_n5055 = new_n5054 ^ new_n3565;
  assign new_n5056 = new_n3460 ^ new_n884;
  assign new_n5057 = new_n5056 ^ new_n3507;
  assign new_n5058 = new_n5057 ^ new_n5055;
  assign new_n5059 = new_n3460 ^ new_n3431;
  assign new_n5060 = new_n5059 ^ new_n3667;
  assign new_n5061 = new_n3539 ^ new_n892;
  assign new_n5062 = new_n5061 ^ new_n3153;
  assign new_n5063 = new_n5062 ^ new_n5060;
  assign new_n5064 = new_n5063 ^ new_n5058;
  assign new_n5065 = new_n5064 ^ new_n5048;
  assign new_n5066 = new_n3636 ^ new_n3466;
  assign new_n5067 = new_n3481 ^ new_n820;
  assign new_n5068 = new_n5067 ^ new_n3602;
  assign new_n5069 = new_n5068 ^ new_n5066;
  assign new_n5070 = new_n3610 ^ new_n3550;
  assign new_n5071 = new_n3615 ^ new_n843;
  assign new_n5072 = new_n5071 ^ new_n3631;
  assign new_n5073 = new_n5072 ^ new_n5070;
  assign new_n5074 = new_n5073 ^ new_n5069;
  assign new_n5075 = new_n5074 ^ new_n5065;
  assign new_n5076 = new_n5053 & new_n5075;
  assign new_n5077 = new_n5064 ^ new_n5052;
  assign new_n5078 = new_n5077 ^ new_n5069;
  assign new_n5079 = new_n5048 & new_n5078;
  assign new_n5080 = new_n5079 ^ new_n5076;
  assign new_n5081 = new_n5077 ^ new_n5073;
  assign new_n5082 = new_n5081 ^ new_n5080;
  assign new_n5083 = new_n3460 ^ new_n3265;
  assign new_n5084 = new_n3403 ^ new_n856;
  assign new_n5085 = new_n5084 ^ new_n3666;
  assign new_n5086 = new_n5085 ^ new_n5083;
  assign new_n5087 = new_n5086 ^ new_n5074;
  assign new_n5088 = new_n5087 ^ new_n5042;
  assign new_n5089 = new_n5086 ^ new_n5078;
  assign new_n5090 = new_n5088 & new_n5089;
  assign new_n5091 = new_n5063 ^ new_n5042;
  assign new_n5092 = new_n5081 & new_n5091;
  assign new_n5093 = new_n5092 ^ new_n5090;
  assign new_n5094 = new_n5093 ^ new_n5042;
  assign new_n5095 = new_n5094 ^ new_n5082;
  assign new_n5096 = ~new_n5063 & ~new_n5087;
  assign new_n5097 = new_n5096 ^ new_n5063;
  assign new_n5098 = new_n5097 ^ new_n5092;
  assign new_n5099 = new_n5098 ^ new_n5053;
  assign new_n5100 = new_n5052 ^ new_n5047;
  assign new_n5101 = new_n5073 ^ new_n5047;
  assign new_n5102 = new_n5101 ^ new_n5053;
  assign new_n5103 = new_n5100 & new_n5102;
  assign new_n5104 = new_n5103 ^ new_n5079;
  assign new_n5105 = new_n5073 ^ new_n5058;
  assign new_n5106 = new_n5105 ^ new_n5104;
  assign new_n5107 = new_n5106 ^ new_n5099;
  assign new_n5108 = new_n5100 ^ new_n5091;
  assign new_n5109 = new_n5065 & new_n5108;
  assign new_n5110 = new_n5109 ^ new_n5069;
  assign new_n5111 = new_n5110 ^ new_n5065;
  assign new_n5112 = new_n5087 ^ new_n5063;
  assign new_n5113 = new_n5112 ^ new_n5053;
  assign new_n5114 = new_n5086 ^ new_n5065;
  assign new_n5115 = new_n5113 & new_n5114;
  assign new_n5116 = new_n5115 ^ new_n5104;
  assign new_n5117 = new_n5116 ^ new_n5052;
  assign new_n5118 = new_n5117 ^ new_n5111;
  assign new_n5119 = ~new_n5107 & new_n5118;
  assign new_n5120 = new_n5119 ^ new_n5095;
  assign new_n5121 = new_n5073 ^ new_n5042;
  assign new_n5122 = new_n5087 ^ new_n5047;
  assign new_n5123 = new_n5086 & new_n5122;
  assign new_n5124 = new_n5123 ^ new_n5115;
  assign new_n5125 = new_n5103 ^ new_n5076;
  assign new_n5126 = new_n5125 ^ new_n5124;
  assign new_n5127 = new_n5126 ^ new_n5121;
  assign new_n5128 = new_n5120 & new_n5127;
  assign new_n5129 = new_n5123 ^ new_n5047;
  assign new_n5130 = new_n5129 ^ new_n5110;
  assign new_n5131 = new_n5130 ^ new_n5119;
  assign new_n5132 = new_n5131 ^ new_n5082;
  assign new_n5133 = new_n5096 ^ new_n5090;
  assign new_n5134 = new_n5133 ^ new_n5125;
  assign new_n5135 = ~new_n5134 & new_n5132;
  assign new_n5136 = new_n5135 ^ new_n5128;
  assign new_n5137 = new_n5130 ^ new_n5094;
  assign new_n5138 = new_n5137 ^ new_n5136;
  assign new_n5139 = new_n5048 & new_n5138;
  assign new_n5140 = new_n5078 & new_n5138;
  assign new_n5141 = new_n5140 ^ new_n5139;
  assign new_n5142 = new_n5135 ^ new_n5042;
  assign new_n5143 = new_n5123 ^ new_n5090;
  assign new_n5144 = new_n5073 ^ new_n5063;
  assign new_n5145 = new_n5115 ^ new_n5097;
  assign new_n5146 = new_n5135 ^ new_n5119;
  assign new_n5147 = ~new_n5095 & ~new_n5146;
  assign new_n5148 = new_n5147 ^ new_n5135;
  assign new_n5149 = new_n5130 ^ new_n5128;
  assign new_n5150 = new_n5149 ^ new_n5082;
  assign new_n5151 = ~new_n5148 & new_n5150;
  assign new_n5152 = new_n5148 ^ new_n5120;
  assign new_n5153 = new_n5152 ^ new_n5151;
  assign new_n5154 = new_n5153 ^ new_n5145;
  assign new_n5155 = new_n5154 ^ new_n5144;
  assign new_n5156 = new_n5155 ^ new_n5143;
  assign new_n5157 = new_n5156 ^ new_n5142;
  assign new_n5158 = new_n5053 & new_n5157;
  assign new_n5159 = new_n5152 ^ new_n5107;
  assign new_n5160 = new_n5065 & new_n5159;
  assign new_n5161 = new_n5135 ^ new_n5095;
  assign new_n5162 = new_n5086 & new_n5161;
  assign new_n5163 = new_n5162 ^ new_n5160;
  assign new_n5164 = new_n5151 ^ new_n5128;
  assign new_n5165 = new_n5164 ^ new_n5118;
  assign new_n5166 = new_n5091 & new_n5165;
  assign new_n5167 = new_n5166 ^ new_n5163;
  assign new_n5168 = new_n5075 & new_n5157;
  assign new_n5169 = new_n5088 & new_n5150;
  assign new_n5170 = new_n5169 ^ new_n5168;
  assign new_n5171 = new_n5170 ^ new_n5167;
  assign new_n5172 = new_n5171 ^ new_n5158;
  assign new_n5173 = new_n5172 ^ new_n5141;
  assign new_n5174 = new_n4283 ^ new_n425;
  assign new_n5175 = new_n4309 ^ new_n3879;
  assign new_n5176 = new_n5175 ^ new_n4011;
  assign new_n5177 = new_n5176 ^ new_n5174;
  assign new_n5178 = new_n4374 ^ new_n4364;
  assign new_n5179 = new_n5178 ^ new_n4282;
  assign new_n5180 = new_n5179 ^ new_n4403;
  assign new_n5181 = new_n4291 ^ new_n393;
  assign new_n5182 = new_n5181 ^ new_n4326;
  assign new_n5183 = new_n5182 ^ new_n5180;
  assign new_n5184 = new_n5178 ^ new_n403;
  assign new_n5185 = new_n5184 ^ new_n4322;
  assign new_n5186 = new_n4387 ^ new_n4130;
  assign new_n5187 = new_n5186 ^ new_n5185;
  assign new_n5188 = new_n5187 ^ new_n5183;
  assign new_n5189 = new_n5188 ^ new_n5177;
  assign new_n5190 = new_n4416 ^ new_n4372;
  assign new_n5191 = new_n4337 ^ new_n433;
  assign new_n5192 = new_n5191 ^ new_n4409;
  assign new_n5193 = new_n5192 ^ new_n5190;
  assign new_n5194 = new_n5193 ^ new_n5189;
  assign new_n5195 = new_n4358 ^ new_n4020;
  assign new_n5196 = new_n4364 ^ new_n365;
  assign new_n5197 = new_n5196 ^ new_n4337;
  assign new_n5198 = new_n5197 ^ new_n5195;
  assign new_n5199 = new_n4409 ^ new_n4347;
  assign new_n5200 = new_n4388 ^ new_n4380;
  assign new_n5201 = new_n5200 ^ new_n444;
  assign new_n5202 = new_n5201 ^ new_n5199;
  assign new_n5203 = new_n5202 ^ new_n5198;
  assign new_n5204 = new_n5202 ^ new_n5193;
  assign new_n5205 = new_n5178 ^ new_n4402;
  assign new_n5206 = new_n4294 ^ new_n413;
  assign new_n5207 = new_n5206 ^ new_n4249;
  assign new_n5208 = new_n5207 ^ new_n5205;
  assign new_n5209 = new_n5208 ^ new_n5204;
  assign new_n5210 = new_n5209 ^ new_n5183;
  assign new_n5211 = new_n5198 ^ new_n5177;
  assign new_n5212 = new_n5211 ^ new_n5210;
  assign new_n5213 = new_n5178 ^ new_n4412;
  assign new_n5214 = new_n4388 ^ new_n374;
  assign new_n5215 = new_n5214 ^ new_n4241;
  assign new_n5216 = new_n5215 ^ new_n5213;
  assign new_n5217 = new_n5216 ^ new_n5198;
  assign new_n5218 = new_n5217 ^ new_n5188;
  assign new_n5219 = new_n5218 ^ new_n5208;
  assign new_n5220 = new_n5212 & new_n5219;
  assign new_n5221 = new_n5216 ^ new_n5209;
  assign new_n5222 = new_n5208 & new_n5221;
  assign new_n5223 = new_n5222 ^ new_n5220;
  assign new_n5224 = new_n5218 ^ new_n5204;
  assign new_n5225 = new_n5211 & new_n5224;
  assign new_n5226 = new_n5216 ^ new_n5202;
  assign new_n5227 = new_n5226 ^ new_n5211;
  assign new_n5228 = new_n5216 ^ new_n5177;
  assign new_n5229 = new_n5227 & new_n5228;
  assign new_n5230 = new_n5229 ^ new_n5225;
  assign new_n5231 = new_n5230 ^ new_n5223;
  assign new_n5232 = new_n5231 ^ new_n5203;
  assign new_n5233 = new_n5208 ^ new_n5194;
  assign new_n5234 = new_n5209 ^ new_n5198;
  assign new_n5235 = new_n5233 & new_n5234;
  assign new_n5236 = new_n5202 ^ new_n5189;
  assign new_n5237 = new_n5198 ^ new_n5183;
  assign new_n5238 = new_n5236 & new_n5237;
  assign new_n5239 = new_n5238 ^ new_n5235;
  assign new_n5240 = new_n5239 ^ new_n5198;
  assign new_n5241 = new_n5194 & new_n5217;
  assign new_n5242 = new_n5241 ^ new_n5225;
  assign new_n5243 = new_n5242 ^ new_n5236;
  assign new_n5244 = new_n5243 ^ new_n5240;
  assign new_n5245 = ~new_n5183 & ~new_n5209;
  assign new_n5246 = new_n5245 ^ new_n5183;
  assign new_n5247 = new_n5246 ^ new_n5238;
  assign new_n5248 = new_n5247 ^ new_n5211;
  assign new_n5249 = new_n5241 ^ new_n5229;
  assign new_n5250 = new_n5202 ^ new_n5187;
  assign new_n5251 = new_n5250 ^ new_n5249;
  assign new_n5252 = new_n5251 ^ new_n5248;
  assign new_n5253 = new_n5216 ^ new_n5183;
  assign new_n5254 = new_n5253 ^ new_n5211;
  assign new_n5255 = new_n5218 & new_n5254;
  assign new_n5256 = new_n5255 ^ new_n5193;
  assign new_n5257 = new_n5256 ^ new_n5218;
  assign new_n5258 = new_n5249 ^ new_n5220;
  assign new_n5259 = new_n5258 ^ new_n5177;
  assign new_n5260 = new_n5259 ^ new_n5257;
  assign new_n5261 = ~new_n5252 & new_n5260;
  assign new_n5262 = new_n5261 ^ new_n5244;
  assign new_n5263 = new_n5232 & new_n5262;
  assign new_n5264 = new_n5222 ^ new_n5216;
  assign new_n5265 = new_n5264 ^ new_n5256;
  assign new_n5266 = new_n5265 ^ new_n5261;
  assign new_n5267 = new_n5266 ^ new_n5243;
  assign new_n5268 = new_n5245 ^ new_n5235;
  assign new_n5269 = new_n5268 ^ new_n5230;
  assign new_n5270 = ~new_n5269 & new_n5267;
  assign new_n5271 = new_n5270 ^ new_n5263;
  assign new_n5272 = new_n5265 ^ new_n5240;
  assign new_n5273 = new_n5272 ^ new_n5271;
  assign new_n5274 = new_n5194 & new_n5273;
  assign new_n5275 = new_n5217 & new_n5273;
  assign new_n5276 = new_n5275 ^ new_n5274;
  assign new_n5277 = new_n5270 ^ new_n5198;
  assign new_n5278 = new_n5235 ^ new_n5222;
  assign new_n5279 = new_n5202 ^ new_n5183;
  assign new_n5280 = new_n5246 ^ new_n5220;
  assign new_n5281 = new_n5265 ^ new_n5263;
  assign new_n5282 = new_n5281 ^ new_n5243;
  assign new_n5283 = new_n5270 ^ new_n5261;
  assign new_n5284 = ~new_n5283 & new_n5244;
  assign new_n5285 = new_n5284 ^ new_n5261;
  assign new_n5286 = new_n5282 & new_n5285;
  assign new_n5287 = new_n5284 ^ new_n5244;
  assign new_n5288 = new_n5287 ^ new_n5286;
  assign new_n5289 = new_n5288 ^ new_n5280;
  assign new_n5290 = new_n5289 ^ new_n5279;
  assign new_n5291 = new_n5290 ^ new_n5278;
  assign new_n5292 = new_n5291 ^ new_n5277;
  assign new_n5293 = ~new_n5292 & new_n5211;
  assign new_n5294 = ~new_n5292 & new_n5224;
  assign new_n5295 = new_n5234 & new_n5282;
  assign new_n5296 = new_n5295 ^ new_n5294;
  assign new_n5297 = new_n5286 ^ new_n5263;
  assign new_n5298 = new_n5297 ^ new_n5260;
  assign new_n5299 = new_n5237 & new_n5298;
  assign new_n5300 = new_n5287 ^ new_n5252;
  assign new_n5301 = ~new_n5300 & new_n5218;
  assign new_n5302 = new_n5270 ^ new_n5244;
  assign new_n5303 = new_n5208 & new_n5302;
  assign new_n5304 = new_n5303 ^ new_n5301;
  assign new_n5305 = new_n5304 ^ new_n5299;
  assign new_n5306 = new_n5305 ^ new_n5296;
  assign new_n5307 = new_n5306 ^ new_n5293;
  assign new_n5308 = new_n5307 ^ new_n5276;
  assign new_n5309 = new_n5308 ^ new_n5173;
  assign new_n5310 = new_n3619 ^ new_n2033;
  assign new_n5311 = new_n2063 ^ new_n2056;
  assign new_n5312 = new_n5311 ^ new_n1986;
  assign new_n5313 = new_n5312 ^ new_n5310;
  assign new_n5314 = new_n1947 ^ new_n1912;
  assign new_n5315 = new_n5314 ^ new_n1766;
  assign new_n5316 = new_n2026 ^ n126;
  assign new_n5317 = new_n5316 ^ new_n3526;
  assign new_n5318 = new_n5317 ^ new_n5315;
  assign new_n5319 = new_n2015 ^ new_n1514;
  assign new_n5320 = new_n2026 ^ n125;
  assign new_n5321 = new_n5320 ^ new_n5319;
  assign new_n5322 = new_n1996 ^ new_n1990;
  assign new_n5323 = new_n5322 ^ new_n3591;
  assign new_n5324 = new_n5323 ^ new_n1956;
  assign new_n5325 = new_n5324 ^ new_n5321;
  assign new_n5326 = new_n5325 ^ new_n5318;
  assign new_n5327 = new_n5322 ^ new_n2076;
  assign new_n5328 = new_n5327 ^ new_n1920;
  assign new_n5329 = new_n2079 ^ new_n2005;
  assign new_n5330 = new_n5329 ^ new_n3419;
  assign new_n5331 = new_n5330 ^ new_n5328;
  assign new_n5332 = new_n5331 ^ new_n5326;
  assign new_n5333 = new_n5332 ^ new_n5313;
  assign new_n5334 = new_n1974 ^ new_n1966;
  assign new_n5335 = new_n5334 ^ n123;
  assign new_n5336 = new_n3643 ^ new_n2056;
  assign new_n5337 = new_n5336 ^ new_n2043;
  assign new_n5338 = new_n5337 ^ new_n5335;
  assign new_n5339 = new_n2046 ^ new_n2033;
  assign new_n5340 = new_n5339 ^ new_n1775;
  assign new_n5341 = new_n1996 ^ n121;
  assign new_n5342 = new_n5341 ^ new_n3471;
  assign new_n5343 = new_n5342 ^ new_n5340;
  assign new_n5344 = new_n5343 ^ new_n5338;
  assign new_n5345 = new_n3659 ^ new_n1926;
  assign new_n5346 = new_n5322 ^ new_n2080;
  assign new_n5347 = new_n5346 ^ new_n5345;
  assign new_n5348 = new_n5331 ^ new_n5325;
  assign new_n5349 = new_n2059 ^ new_n1400;
  assign new_n5350 = new_n5349 ^ new_n5322;
  assign new_n5351 = new_n1974 ^ new_n1887;
  assign new_n5352 = new_n1514 ^ n124;
  assign new_n5353 = new_n5352 ^ new_n5351;
  assign new_n5354 = new_n5353 ^ new_n5350;
  assign new_n5355 = new_n5354 ^ new_n5343;
  assign new_n5356 = new_n5355 ^ new_n5348;
  assign new_n5357 = new_n5356 ^ new_n5347;
  assign new_n5358 = new_n5338 ^ new_n5313;
  assign new_n5359 = new_n5358 ^ new_n5347;
  assign new_n5360 = new_n5359 ^ new_n5331;
  assign new_n5361 = new_n5343 ^ new_n5318;
  assign new_n5362 = new_n5361 ^ new_n5360;
  assign new_n5363 = ~new_n5357 & ~new_n5362;
  assign new_n5364 = new_n5359 ^ new_n5354;
  assign new_n5365 = ~new_n5347 & ~new_n5364;
  assign new_n5366 = new_n5365 ^ new_n5363;
  assign new_n5367 = new_n5354 ^ new_n5338;
  assign new_n5368 = new_n5367 ^ new_n5361;
  assign new_n5369 = new_n5354 ^ new_n5318;
  assign new_n5370 = new_n5368 & new_n5369;
  assign new_n5371 = new_n5358 ^ new_n5356;
  assign new_n5372 = new_n5361 & new_n5371;
  assign new_n5373 = new_n5372 ^ new_n5370;
  assign new_n5374 = new_n5373 ^ new_n5366;
  assign new_n5375 = new_n5374 ^ new_n5344;
  assign new_n5376 = ~new_n5331 & new_n5359;
  assign new_n5377 = new_n5376 ^ new_n5331;
  assign new_n5378 = new_n5338 ^ new_n5332;
  assign new_n5379 = new_n5343 ^ new_n5331;
  assign new_n5380 = new_n5378 & new_n5379;
  assign new_n5381 = new_n5380 ^ new_n5377;
  assign new_n5382 = new_n5381 ^ new_n5361;
  assign new_n5383 = new_n5333 & new_n5355;
  assign new_n5384 = new_n5383 ^ new_n5370;
  assign new_n5385 = new_n5338 ^ new_n5325;
  assign new_n5386 = new_n5385 ^ new_n5384;
  assign new_n5387 = new_n5386 ^ new_n5382;
  assign new_n5388 = new_n5354 ^ new_n5331;
  assign new_n5389 = new_n5388 ^ new_n5361;
  assign new_n5390 = new_n5356 & new_n5389;
  assign new_n5391 = new_n5390 ^ new_n5313;
  assign new_n5392 = new_n5391 ^ new_n5356;
  assign new_n5393 = new_n5383 ^ new_n5363;
  assign new_n5394 = new_n5370 ^ new_n5318;
  assign new_n5395 = new_n5394 ^ new_n5393;
  assign new_n5396 = new_n5395 ^ new_n5392;
  assign new_n5397 = ~new_n5387 & new_n5396;
  assign new_n5398 = new_n5383 ^ new_n5372;
  assign new_n5399 = new_n5398 ^ new_n5378;
  assign new_n5400 = new_n5347 ^ new_n5333;
  assign new_n5401 = new_n5359 ^ new_n5343;
  assign new_n5402 = ~new_n5400 & ~new_n5401;
  assign new_n5403 = new_n5402 ^ new_n5380;
  assign new_n5404 = new_n5403 ^ new_n5343;
  assign new_n5405 = new_n5404 ^ new_n5399;
  assign new_n5406 = new_n5405 ^ new_n5397;
  assign new_n5407 = new_n5375 & new_n5406;
  assign new_n5408 = new_n5365 ^ new_n5354;
  assign new_n5409 = new_n5408 ^ new_n5391;
  assign new_n5410 = new_n5409 ^ new_n5397;
  assign new_n5411 = new_n5410 ^ new_n5399;
  assign new_n5412 = new_n5402 ^ new_n5376;
  assign new_n5413 = new_n5412 ^ new_n5373;
  assign new_n5414 = ~new_n5413 & new_n5411;
  assign new_n5415 = new_n5414 ^ new_n5407;
  assign new_n5416 = new_n5409 ^ new_n5404;
  assign new_n5417 = new_n5416 ^ new_n5415;
  assign new_n5418 = new_n5333 & new_n5417;
  assign new_n5419 = new_n5338 ^ new_n5331;
  assign new_n5420 = new_n5377 ^ new_n5363;
  assign new_n5421 = new_n5409 ^ new_n5407;
  assign new_n5422 = new_n5421 ^ new_n5399;
  assign new_n5423 = new_n5414 ^ new_n5397;
  assign new_n5424 = ~new_n5423 & new_n5405;
  assign new_n5425 = new_n5424 ^ new_n5397;
  assign new_n5426 = new_n5422 & new_n5425;
  assign new_n5427 = new_n5424 ^ new_n5405;
  assign new_n5428 = new_n5427 ^ new_n5426;
  assign new_n5429 = new_n5428 ^ new_n5420;
  assign new_n5430 = new_n5429 ^ new_n5419;
  assign new_n5431 = new_n5430 ^ new_n5354;
  assign new_n5432 = new_n5407 ^ new_n5380;
  assign new_n5433 = new_n5432 ^ new_n5391;
  assign new_n5434 = new_n5433 ^ new_n5431;
  assign new_n5435 = ~new_n5434 & new_n5368;
  assign new_n5436 = new_n5435 ^ new_n5418;
  assign new_n5437 = new_n5427 ^ new_n5414;
  assign new_n5438 = new_n5437 ^ new_n5413;
  assign new_n5439 = ~new_n5357 & ~new_n5438;
  assign new_n5440 = new_n5427 ^ new_n5387;
  assign new_n5441 = ~new_n5440 & new_n5356;
  assign new_n5442 = new_n5441 ^ new_n5439;
  assign new_n5443 = ~new_n5440 & new_n5389;
  assign new_n5444 = new_n5443 ^ new_n5442;
  assign new_n5445 = ~new_n5362 & ~new_n5438;
  assign new_n5446 = new_n5355 & new_n5417;
  assign new_n5447 = ~new_n5434 & new_n5369;
  assign new_n5448 = new_n5447 ^ new_n5446;
  assign new_n5449 = new_n5448 ^ new_n5445;
  assign new_n5450 = new_n5449 ^ new_n5444;
  assign new_n5451 = new_n5450 ^ new_n5436;
  assign new_n5452 = new_n5290 ^ new_n5216;
  assign new_n5453 = new_n5263 ^ new_n5238;
  assign new_n5454 = new_n5453 ^ new_n5256;
  assign new_n5455 = new_n5454 ^ new_n5452;
  assign new_n5456 = ~new_n5455 & new_n5227;
  assign new_n5457 = new_n5456 ^ new_n5274;
  assign new_n5458 = new_n5287 ^ new_n5270;
  assign new_n5459 = new_n5458 ^ new_n5269;
  assign new_n5460 = ~new_n5459 & new_n5219;
  assign new_n5461 = new_n5460 ^ new_n5301;
  assign new_n5462 = ~new_n5300 & new_n5254;
  assign new_n5463 = new_n5462 ^ new_n5461;
  assign new_n5464 = ~new_n5459 & new_n5212;
  assign new_n5465 = ~new_n5455 & new_n5228;
  assign new_n5466 = new_n5465 ^ new_n5275;
  assign new_n5467 = new_n5466 ^ new_n5464;
  assign new_n5468 = new_n5467 ^ new_n5463;
  assign new_n5469 = new_n5468 ^ new_n5457;
  assign new_n5470 = new_n5469 ^ new_n5451;
  assign new_n5471 = new_n5470 ^ new_n5309;
  assign new_n5472 = new_n5471 ^ new_n5038;
  assign new_n5473 = new_n841 ^ new_n559;
  assign new_n5474 = new_n5032 ^ new_n5004;
  assign new_n5475 = new_n4984 & new_n5008;
  assign new_n5476 = new_n5000 ^ new_n4930;
  assign new_n5477 = new_n4986 ^ new_n4951;
  assign new_n5478 = new_n5477 ^ new_n5016;
  assign new_n5479 = new_n5478 ^ new_n5476;
  assign new_n5480 = ~new_n5479 & new_n4957;
  assign new_n5481 = new_n5480 ^ new_n5475;
  assign new_n5482 = new_n5012 ^ new_n4993;
  assign new_n5483 = new_n5482 ^ new_n4982;
  assign new_n5484 = new_n4965 & new_n5483;
  assign new_n5485 = new_n5000 ^ new_n4991;
  assign new_n5486 = new_n4935 & new_n5485;
  assign new_n5487 = new_n5486 ^ new_n5027;
  assign new_n5488 = new_n5487 ^ new_n5484;
  assign new_n5489 = new_n5488 ^ new_n5481;
  assign new_n5490 = ~new_n5479 & new_n4947;
  assign new_n5491 = new_n5490 ^ new_n5489;
  assign new_n5492 = new_n5491 ^ new_n5474;
  assign new_n5493 = new_n5492 ^ new_n5473;
  assign new_n5494 = new_n5152 ^ new_n5135;
  assign new_n5495 = new_n5494 ^ new_n5134;
  assign new_n5496 = new_n5114 & new_n5495;
  assign new_n5497 = new_n5496 ^ new_n5160;
  assign new_n5498 = new_n5108 & new_n5159;
  assign new_n5499 = new_n5498 ^ new_n5497;
  assign new_n5500 = new_n5113 & new_n5495;
  assign new_n5501 = new_n5155 ^ new_n5047;
  assign new_n5502 = new_n5128 ^ new_n5092;
  assign new_n5503 = new_n5502 ^ new_n5110;
  assign new_n5504 = new_n5503 ^ new_n5501;
  assign new_n5505 = new_n5100 & new_n5504;
  assign new_n5506 = new_n5505 ^ new_n5139;
  assign new_n5507 = new_n5506 ^ new_n5500;
  assign new_n5508 = new_n5151 ^ new_n5127;
  assign new_n5509 = new_n5087 & new_n5508;
  assign new_n5510 = new_n5509 ^ new_n5507;
  assign new_n5511 = new_n5081 & new_n5165;
  assign new_n5512 = new_n5511 ^ new_n5510;
  assign new_n5513 = new_n5512 ^ new_n5499;
  assign new_n5514 = new_n5286 ^ new_n5232;
  assign new_n5515 = new_n5209 & new_n5514;
  assign new_n5516 = new_n5515 ^ new_n5467;
  assign new_n5517 = new_n5236 & new_n5298;
  assign new_n5518 = new_n5517 ^ new_n5516;
  assign new_n5519 = new_n5518 ^ new_n5463;
  assign new_n5520 = new_n5519 ^ new_n5513;
  assign new_n5521 = new_n5446 ^ new_n5418;
  assign new_n5522 = ~new_n5401 & new_n5422;
  assign new_n5523 = new_n5414 ^ new_n5343;
  assign new_n5524 = new_n5402 ^ new_n5365;
  assign new_n5525 = new_n5524 ^ new_n5430;
  assign new_n5526 = new_n5525 ^ new_n5523;
  assign new_n5527 = ~new_n5526 & new_n5371;
  assign new_n5528 = new_n5527 ^ new_n5522;
  assign new_n5529 = new_n5426 ^ new_n5407;
  assign new_n5530 = new_n5529 ^ new_n5396;
  assign new_n5531 = new_n5379 & new_n5530;
  assign new_n5532 = new_n5414 ^ new_n5405;
  assign new_n5533 = ~new_n5347 & new_n5532;
  assign new_n5534 = new_n5533 ^ new_n5441;
  assign new_n5535 = new_n5534 ^ new_n5531;
  assign new_n5536 = new_n5535 ^ new_n5528;
  assign new_n5537 = ~new_n5526 & new_n5361;
  assign new_n5538 = new_n5537 ^ new_n5536;
  assign new_n5539 = new_n5538 ^ new_n5521;
  assign new_n5540 = new_n5539 ^ new_n5308;
  assign new_n5541 = new_n5540 ^ new_n5520;
  assign new_n5542 = new_n5541 ^ new_n5493;
  assign new_n5543 = new_n5542 ^ new_n5472;
  assign new_n5544 = new_n854 ^ new_n574;
  assign new_n5545 = ~new_n5400 & new_n5422;
  assign new_n5546 = new_n5426 ^ new_n5375;
  assign new_n5547 = ~new_n5360 & new_n5546;
  assign new_n5548 = new_n5547 ^ new_n5545;
  assign new_n5549 = new_n5548 ^ new_n5448;
  assign new_n5550 = new_n5378 & new_n5530;
  assign new_n5551 = new_n5550 ^ new_n5535;
  assign new_n5552 = new_n5551 ^ new_n5549;
  assign new_n5553 = new_n5552 ^ new_n5544;
  assign new_n5554 = new_n5518 ^ new_n5456;
  assign new_n5555 = new_n5462 ^ new_n5274;
  assign new_n5556 = new_n5555 ^ new_n5554;
  assign new_n5557 = new_n5102 & new_n5504;
  assign new_n5558 = new_n5557 ^ new_n5512;
  assign new_n5559 = new_n5498 ^ new_n5140;
  assign new_n5560 = new_n5559 ^ new_n5558;
  assign new_n5561 = new_n5560 ^ new_n5556;
  assign new_n5562 = new_n5210 & new_n5514;
  assign new_n5563 = new_n5233 & new_n5282;
  assign new_n5564 = new_n5563 ^ new_n5562;
  assign new_n5565 = new_n5564 ^ new_n5466;
  assign new_n5566 = new_n5517 ^ new_n5305;
  assign new_n5567 = new_n5566 ^ new_n5565;
  assign new_n5568 = new_n5012 ^ new_n4961;
  assign new_n5569 = new_n4946 & new_n5568;
  assign new_n5570 = new_n4985 & new_n5008;
  assign new_n5571 = new_n5570 ^ new_n5569;
  assign new_n5572 = new_n5571 ^ new_n5034;
  assign new_n5573 = new_n4964 & new_n5483;
  assign new_n5574 = new_n5573 ^ new_n5488;
  assign new_n5575 = new_n5574 ^ new_n5572;
  assign new_n5576 = new_n5575 ^ new_n5567;
  assign new_n5577 = new_n5576 ^ new_n5561;
  assign new_n5578 = new_n5577 ^ new_n5553;
  assign new_n5579 = new_n5578 ^ new_n5543;
  assign new_n5580 = new_n5089 & new_n5150;
  assign new_n5581 = new_n5580 ^ new_n5498;
  assign new_n5582 = new_n5496 ^ new_n5162;
  assign new_n5583 = new_n5582 ^ new_n5510;
  assign new_n5584 = new_n5583 ^ new_n5581;
  assign new_n5585 = new_n5563 ^ new_n5462;
  assign new_n5586 = new_n5460 ^ new_n5303;
  assign new_n5587 = new_n5586 ^ new_n5516;
  assign new_n5588 = new_n5587 ^ new_n5585;
  assign new_n5589 = new_n5588 ^ new_n5584;
  assign new_n5590 = ~new_n5359 & new_n5546;
  assign new_n5591 = new_n5590 ^ new_n5449;
  assign new_n5592 = new_n5591 ^ new_n5550;
  assign new_n5593 = new_n5592 ^ new_n5444;
  assign new_n5594 = new_n5593 ^ new_n5519;
  assign new_n5595 = new_n5594 ^ new_n5589;
  assign new_n5596 = new_n862 ^ new_n539;
  assign new_n5597 = new_n5596 ^ n108;
  assign new_n5598 = new_n4945 & new_n5568;
  assign new_n5599 = new_n5598 ^ new_n5035;
  assign new_n5600 = new_n5599 ^ new_n5573;
  assign new_n5601 = new_n5600 ^ new_n5030;
  assign new_n5602 = new_n5601 ^ new_n5597;
  assign new_n5603 = new_n5602 ^ new_n5561;
  assign new_n5604 = new_n5603 ^ new_n5595;
  assign new_n5605 = new_n5604 ^ new_n5579;
  assign new_n5606 = ~new_n5578 & ~new_n5605;
  assign new_n5607 = new_n5606 ^ new_n5604;
  assign new_n5608 = new_n872 ^ new_n583;
  assign new_n5609 = new_n5608 ^ n105;
  assign new_n5610 = new_n5029 ^ new_n5004;
  assign new_n5611 = new_n5600 ^ new_n5021;
  assign new_n5612 = new_n5611 ^ new_n5610;
  assign new_n5613 = new_n5612 ^ new_n5609;
  assign new_n5614 = new_n5557 ^ new_n5140;
  assign new_n5615 = new_n5507 ^ new_n5499;
  assign new_n5616 = new_n5615 ^ new_n5614;
  assign new_n5617 = new_n5616 ^ new_n5469;
  assign new_n5618 = new_n5443 ^ new_n5418;
  assign new_n5619 = new_n5592 ^ new_n5435;
  assign new_n5620 = new_n5619 ^ new_n5618;
  assign new_n5621 = new_n5620 ^ new_n5556;
  assign new_n5622 = new_n5621 ^ new_n5617;
  assign new_n5623 = new_n5622 ^ new_n5613;
  assign new_n5624 = new_n5623 ^ new_n5604;
  assign new_n5625 = new_n5299 ^ new_n5294;
  assign new_n5626 = new_n5515 ^ new_n5456;
  assign new_n5627 = new_n5626 ^ new_n5565;
  assign new_n5628 = new_n5627 ^ new_n5625;
  assign new_n5629 = new_n5484 ^ new_n5480;
  assign new_n5630 = new_n5598 ^ new_n5021;
  assign new_n5631 = new_n5630 ^ new_n5572;
  assign new_n5632 = new_n5631 ^ new_n5629;
  assign new_n5633 = new_n5632 ^ new_n5628;
  assign new_n5634 = new_n5633 ^ new_n5561;
  assign new_n5635 = new_n5112 & new_n5508;
  assign new_n5636 = new_n5635 ^ new_n5580;
  assign new_n5637 = new_n5636 ^ new_n5506;
  assign new_n5638 = new_n5511 ^ new_n5167;
  assign new_n5639 = new_n5638 ^ new_n5637;
  assign new_n5640 = new_n5639 ^ new_n5567;
  assign new_n5641 = new_n890 ^ new_n590;
  assign new_n5642 = new_n5531 ^ new_n5527;
  assign new_n5643 = new_n5590 ^ new_n5435;
  assign new_n5644 = new_n5643 ^ new_n5549;
  assign new_n5645 = new_n5644 ^ new_n5642;
  assign new_n5646 = new_n5645 ^ new_n5641;
  assign new_n5647 = new_n5646 ^ new_n5640;
  assign new_n5648 = new_n5647 ^ new_n5634;
  assign new_n5649 = new_n881 ^ new_n596;
  assign new_n5650 = new_n5649 ^ n109;
  assign new_n5651 = new_n5570 ^ new_n5029;
  assign new_n5652 = new_n5486 ^ new_n5025;
  assign new_n5653 = new_n5652 ^ new_n5599;
  assign new_n5654 = new_n5653 ^ new_n5651;
  assign new_n5655 = new_n5654 ^ new_n5650;
  assign new_n5656 = new_n5655 ^ new_n5561;
  assign new_n5657 = new_n5221 & new_n5302;
  assign new_n5658 = new_n5657 ^ new_n5554;
  assign new_n5659 = new_n5658 ^ new_n5306;
  assign new_n5660 = new_n5122 & new_n5161;
  assign new_n5661 = new_n5660 ^ new_n5558;
  assign new_n5662 = new_n5661 ^ new_n5171;
  assign new_n5663 = new_n5662 ^ new_n5659;
  assign new_n5664 = new_n5545 ^ new_n5443;
  assign new_n5665 = new_n5533 ^ new_n5439;
  assign new_n5666 = new_n5665 ^ new_n5591;
  assign new_n5667 = new_n5666 ^ new_n5664;
  assign new_n5668 = new_n5667 ^ new_n5588;
  assign new_n5669 = new_n5668 ^ new_n5663;
  assign new_n5670 = new_n5669 ^ new_n5656;
  assign new_n5671 = new_n5670 ^ new_n5648;
  assign new_n5672 = new_n5671 ^ new_n5624;
  assign new_n5673 = new_n5648 ^ new_n5604;
  assign new_n5674 = new_n5168 ^ new_n5166;
  assign new_n5675 = new_n5557 ^ new_n5509;
  assign new_n5676 = new_n5675 ^ new_n5637;
  assign new_n5677 = new_n5676 ^ new_n5674;
  assign new_n5678 = ~new_n5364 & new_n5532;
  assign new_n5679 = new_n5678 ^ new_n5619;
  assign new_n5680 = new_n5679 ^ new_n5536;
  assign new_n5681 = new_n5680 ^ new_n5659;
  assign new_n5682 = new_n5681 ^ new_n5677;
  assign new_n5683 = new_n900 ^ new_n604;
  assign new_n5684 = new_n5683 ^ n110;
  assign new_n5685 = new_n4950 & new_n5485;
  assign new_n5686 = new_n5685 ^ new_n5611;
  assign new_n5687 = new_n5686 ^ new_n5489;
  assign new_n5688 = new_n5687 ^ new_n5684;
  assign new_n5689 = new_n5688 ^ new_n5628;
  assign new_n5690 = new_n5689 ^ new_n5682;
  assign new_n5691 = new_n5690 ^ new_n5623;
  assign new_n5692 = new_n5691 ^ new_n5673;
  assign new_n5693 = ~new_n5672 & ~new_n5692;
  assign new_n5694 = new_n5693 ^ new_n5472;
  assign new_n5695 = new_n5694 ^ new_n5607;
  assign new_n5696 = new_n5648 ^ new_n5623;
  assign new_n5697 = new_n5690 ^ new_n5671;
  assign new_n5698 = new_n5697 ^ new_n5542;
  assign new_n5699 = ~new_n5696 & new_n5698;
  assign new_n5700 = new_n5579 & new_n5648;
  assign new_n5701 = new_n5700 ^ new_n5648;
  assign new_n5702 = new_n5701 ^ new_n5699;
  assign new_n5703 = new_n5702 ^ new_n5691;
  assign new_n5704 = new_n5697 ^ new_n5472;
  assign new_n5705 = new_n5624 & new_n5704;
  assign new_n5706 = new_n5604 ^ new_n5542;
  assign new_n5707 = new_n5706 ^ new_n5691;
  assign new_n5708 = new_n5690 ^ new_n5604;
  assign new_n5709 = ~new_n5707 & new_n5708;
  assign new_n5710 = new_n5709 ^ new_n5705;
  assign new_n5711 = new_n5670 ^ new_n5542;
  assign new_n5712 = new_n5711 ^ new_n5710;
  assign new_n5713 = new_n5712 ^ new_n5703;
  assign new_n5714 = new_n5694 ^ new_n5672;
  assign new_n5715 = new_n5672 ^ new_n5578;
  assign new_n5716 = new_n5648 ^ new_n5579;
  assign new_n5717 = new_n5716 ^ new_n5691;
  assign new_n5718 = new_n5715 & new_n5717;
  assign new_n5719 = new_n5718 ^ new_n5710;
  assign new_n5720 = new_n5719 ^ new_n5690;
  assign new_n5721 = new_n5720 ^ new_n5714;
  assign new_n5722 = ~new_n5713 & new_n5721;
  assign new_n5723 = new_n5722 ^ new_n5695;
  assign new_n5724 = new_n5672 ^ new_n5543;
  assign new_n5725 = ~new_n5724 & new_n5691;
  assign new_n5726 = new_n5725 ^ new_n5705;
  assign new_n5727 = new_n5726 ^ new_n5698;
  assign new_n5728 = new_n5727 ^ new_n5723;
  assign new_n5729 = new_n5725 ^ new_n5709;
  assign new_n5730 = new_n5623 ^ new_n5579;
  assign new_n5731 = new_n5704 ^ new_n5578;
  assign new_n5732 = ~new_n5730 & ~new_n5731;
  assign new_n5733 = new_n5732 ^ new_n5700;
  assign new_n5734 = new_n5733 ^ new_n5729;
  assign new_n5735 = ~new_n5728 & ~new_n5734;
  assign new_n5736 = new_n5732 ^ new_n5699;
  assign new_n5737 = new_n5736 ^ new_n5623;
  assign new_n5738 = new_n5737 ^ new_n5727;
  assign new_n5739 = new_n5738 ^ new_n5735;
  assign new_n5740 = ~new_n5605 & new_n5739;
  assign new_n5741 = new_n5735 ^ new_n5722;
  assign new_n5742 = ~new_n5738 & ~new_n5741;
  assign new_n5743 = new_n5742 ^ new_n5735;
  assign new_n5744 = new_n5738 ^ new_n5722;
  assign new_n5745 = new_n5623 ^ new_n5542;
  assign new_n5746 = new_n5718 ^ new_n5606;
  assign new_n5747 = new_n5746 ^ new_n5729;
  assign new_n5748 = new_n5747 ^ new_n5745;
  assign new_n5749 = ~new_n5748 & new_n5744;
  assign new_n5750 = new_n5749 ^ new_n5695;
  assign new_n5751 = new_n5750 ^ new_n5727;
  assign new_n5752 = ~new_n5743 & ~new_n5751;
  assign new_n5753 = new_n5752 ^ new_n5749;
  assign new_n5754 = new_n5753 ^ new_n5721;
  assign new_n5755 = new_n5698 & new_n5754;
  assign new_n5756 = new_n5752 ^ new_n5748;
  assign new_n5757 = ~new_n5579 & ~new_n5756;
  assign new_n5758 = new_n5749 ^ new_n5735;
  assign new_n5759 = new_n5737 ^ new_n5695;
  assign new_n5760 = new_n5759 ^ new_n5758;
  assign new_n5761 = ~new_n5760 & new_n5624;
  assign new_n5762 = new_n5648 ^ new_n5542;
  assign new_n5763 = new_n5718 ^ new_n5701;
  assign new_n5764 = new_n5744 ^ new_n5743;
  assign new_n5765 = new_n5764 ^ new_n5752;
  assign new_n5766 = new_n5765 ^ new_n5763;
  assign new_n5767 = new_n5766 ^ new_n5762;
  assign new_n5768 = new_n5767 ^ new_n5604;
  assign new_n5769 = new_n5749 ^ new_n5699;
  assign new_n5770 = new_n5769 ^ new_n5694;
  assign new_n5771 = new_n5770 ^ new_n5768;
  assign new_n5772 = new_n5708 & new_n5771;
  assign new_n5773 = new_n5772 ^ new_n5761;
  assign new_n5774 = new_n5764 ^ new_n5735;
  assign new_n5775 = new_n5774 ^ new_n5734;
  assign new_n5776 = new_n5717 & new_n5775;
  assign new_n5777 = new_n5776 ^ new_n5773;
  assign new_n5778 = new_n5777 ^ new_n5757;
  assign new_n5779 = new_n5778 ^ new_n5755;
  assign new_n5780 = ~new_n5707 & new_n5771;
  assign new_n5781 = new_n5780 ^ new_n5779;
  assign new_n5782 = new_n5781 ^ new_n5740;
  assign new_n5783 = ~new_n5730 & ~new_n5751;
  assign new_n5784 = new_n5735 ^ new_n5623;
  assign new_n5785 = new_n5732 ^ new_n5606;
  assign new_n5786 = new_n5785 ^ new_n5767;
  assign new_n5787 = new_n5786 ^ new_n5784;
  assign new_n5788 = ~new_n5724 & ~new_n5787;
  assign new_n5789 = new_n5788 ^ new_n5783;
  assign new_n5790 = new_n5764 ^ new_n5713;
  assign new_n5791 = ~new_n5672 & new_n5790;
  assign new_n5792 = ~new_n5578 & new_n5739;
  assign new_n5793 = new_n5792 ^ new_n5791;
  assign new_n5794 = ~new_n5696 & new_n5754;
  assign new_n5795 = new_n5794 ^ new_n5793;
  assign new_n5796 = new_n5795 ^ new_n5789;
  assign new_n5797 = new_n5796 ^ new_n5782;
  assign new_n5798 = new_n4359 ^ new_n876;
  assign new_n5799 = new_n4364 ^ new_n4016;
  assign new_n5800 = new_n5799 ^ new_n4374;
  assign new_n5801 = new_n5800 ^ new_n5798;
  assign new_n5802 = new_n4240 ^ new_n3886;
  assign new_n5803 = new_n5802 ^ new_n866;
  assign new_n5804 = new_n5803 ^ new_n4375;
  assign new_n5805 = new_n5200 ^ new_n4411;
  assign new_n5806 = new_n5805 ^ new_n5804;
  assign new_n5807 = new_n5806 ^ new_n5801;
  assign new_n5808 = new_n4321 ^ new_n3879;
  assign new_n5809 = new_n4386 ^ new_n885;
  assign new_n5810 = new_n5809 ^ new_n5808;
  assign new_n5811 = new_n4375 ^ new_n4241;
  assign new_n5812 = new_n5811 ^ new_n5810;
  assign new_n5813 = new_n4375 ^ new_n4283;
  assign new_n5814 = new_n4400 ^ new_n4294;
  assign new_n5815 = new_n4326 ^ new_n893;
  assign new_n5816 = new_n5815 ^ new_n5814;
  assign new_n5817 = new_n5816 ^ new_n5813;
  assign new_n5818 = new_n5817 ^ new_n5812;
  assign new_n5819 = new_n5818 ^ new_n5807;
  assign new_n5820 = new_n4249 ^ new_n857;
  assign new_n5821 = new_n4403 ^ new_n4375;
  assign new_n5822 = new_n5821 ^ new_n5820;
  assign new_n5823 = new_n5822 ^ new_n5819;
  assign new_n5824 = new_n4011 ^ new_n904;
  assign new_n5825 = new_n4291 ^ new_n4266;
  assign new_n5826 = new_n5825 ^ new_n4322;
  assign new_n5827 = new_n5826 ^ new_n5824;
  assign new_n5828 = new_n5827 ^ new_n5818;
  assign new_n5829 = new_n4417 ^ new_n4358;
  assign new_n5830 = new_n4371 ^ new_n821;
  assign new_n5831 = new_n5830 ^ new_n4337;
  assign new_n5832 = new_n5831 ^ new_n5829;
  assign new_n5833 = new_n5832 ^ new_n5828;
  assign new_n5834 = new_n5807 & new_n5833;
  assign new_n5835 = new_n5827 ^ new_n5801;
  assign new_n5836 = new_n4416 ^ new_n4381;
  assign new_n5837 = new_n4346 ^ new_n844;
  assign new_n5838 = new_n5837 ^ new_n4409;
  assign new_n5839 = new_n5838 ^ new_n5836;
  assign new_n5840 = new_n5839 ^ new_n5832;
  assign new_n5841 = new_n5840 ^ new_n5819;
  assign new_n5842 = new_n5835 & new_n5841;
  assign new_n5843 = new_n5842 ^ new_n5834;
  assign new_n5844 = new_n5839 ^ new_n5828;
  assign new_n5845 = new_n5844 ^ new_n5843;
  assign new_n5846 = new_n5817 ^ new_n5801;
  assign new_n5847 = new_n5844 & new_n5846;
  assign new_n5848 = new_n5833 ^ new_n5822;
  assign new_n5849 = new_n5840 ^ new_n5822;
  assign new_n5850 = new_n5849 ^ new_n5801;
  assign new_n5851 = new_n5848 & new_n5850;
  assign new_n5852 = new_n5851 ^ new_n5847;
  assign new_n5853 = new_n5852 ^ new_n5801;
  assign new_n5854 = new_n5853 ^ new_n5845;
  assign new_n5855 = new_n5849 ^ new_n5806;
  assign new_n5856 = new_n5822 & new_n5855;
  assign new_n5857 = new_n5856 ^ new_n5806;
  assign new_n5858 = new_n5817 ^ new_n5806;
  assign new_n5859 = new_n5858 ^ new_n5835;
  assign new_n5860 = new_n5819 & new_n5859;
  assign new_n5861 = new_n5860 ^ new_n5832;
  assign new_n5862 = new_n5861 ^ new_n5857;
  assign new_n5863 = ~new_n5817 & ~new_n5849;
  assign new_n5864 = new_n5863 ^ new_n5817;
  assign new_n5865 = new_n5864 ^ new_n5847;
  assign new_n5866 = new_n5865 ^ new_n5835;
  assign new_n5867 = new_n5839 ^ new_n5806;
  assign new_n5868 = new_n5867 ^ new_n5835;
  assign new_n5869 = new_n5827 ^ new_n5806;
  assign new_n5870 = new_n5868 & new_n5869;
  assign new_n5871 = new_n5870 ^ new_n5834;
  assign new_n5872 = new_n5839 ^ new_n5812;
  assign new_n5873 = new_n5872 ^ new_n5871;
  assign new_n5874 = new_n5873 ^ new_n5866;
  assign new_n5875 = new_n5861 ^ new_n5819;
  assign new_n5876 = new_n5849 ^ new_n5817;
  assign new_n5877 = new_n5876 ^ new_n5835;
  assign new_n5878 = new_n5823 & new_n5877;
  assign new_n5879 = new_n5878 ^ new_n5834;
  assign new_n5880 = new_n5870 ^ new_n5827;
  assign new_n5881 = new_n5880 ^ new_n5879;
  assign new_n5882 = new_n5881 ^ new_n5875;
  assign new_n5883 = ~new_n5874 & new_n5882;
  assign new_n5884 = new_n5883 ^ new_n5862;
  assign new_n5885 = new_n5884 ^ new_n5845;
  assign new_n5886 = new_n5863 ^ new_n5851;
  assign new_n5887 = new_n5870 ^ new_n5842;
  assign new_n5888 = new_n5887 ^ new_n5886;
  assign new_n5889 = ~new_n5888 & new_n5885;
  assign new_n5890 = new_n5889 ^ new_n5883;
  assign new_n5891 = new_n5854 & new_n5890;
  assign new_n5892 = new_n5891 ^ new_n5889;
  assign new_n5893 = new_n5892 ^ new_n5888;
  assign new_n5894 = ~new_n5893 & new_n5823;
  assign new_n5895 = new_n5891 ^ new_n5874;
  assign new_n5896 = ~new_n5895 & new_n5819;
  assign new_n5897 = new_n5896 ^ new_n5894;
  assign new_n5898 = ~new_n5895 & new_n5859;
  assign new_n5899 = new_n5898 ^ new_n5897;
  assign new_n5900 = new_n5839 ^ new_n5801;
  assign new_n5901 = new_n5878 ^ new_n5856;
  assign new_n5902 = new_n5901 ^ new_n5887;
  assign new_n5903 = new_n5902 ^ new_n5900;
  assign new_n5904 = new_n5883 ^ new_n5854;
  assign new_n5905 = new_n5903 & new_n5904;
  assign new_n5906 = new_n5905 ^ new_n5862;
  assign new_n5907 = new_n5906 ^ new_n5845;
  assign new_n5908 = new_n5904 ^ new_n5891;
  assign new_n5909 = new_n5907 & new_n5908;
  assign new_n5910 = new_n5909 ^ new_n5905;
  assign new_n5911 = new_n5910 ^ new_n5882;
  assign new_n5912 = new_n5844 & new_n5911;
  assign new_n5913 = ~new_n5893 & new_n5877;
  assign new_n5914 = new_n5905 ^ new_n5889;
  assign new_n5915 = new_n5862 ^ new_n5853;
  assign new_n5916 = new_n5915 ^ new_n5914;
  assign new_n5917 = new_n5807 & new_n5916;
  assign new_n5918 = new_n5839 ^ new_n5817;
  assign new_n5919 = new_n5878 ^ new_n5864;
  assign new_n5920 = new_n5909 ^ new_n5891;
  assign new_n5921 = new_n5920 ^ new_n5919;
  assign new_n5922 = new_n5921 ^ new_n5918;
  assign new_n5923 = new_n5922 ^ new_n5806;
  assign new_n5924 = new_n5905 ^ new_n5847;
  assign new_n5925 = new_n5924 ^ new_n5861;
  assign new_n5926 = new_n5925 ^ new_n5923;
  assign new_n5927 = ~new_n5926 & new_n5869;
  assign new_n5928 = new_n5927 ^ new_n5917;
  assign new_n5929 = new_n5928 ^ new_n5913;
  assign new_n5930 = new_n5909 ^ new_n5903;
  assign new_n5931 = new_n5849 & new_n5930;
  assign new_n5932 = new_n5931 ^ new_n5929;
  assign new_n5933 = new_n5932 ^ new_n5912;
  assign new_n5934 = new_n5933 ^ new_n5899;
  assign new_n5935 = new_n3376 ^ new_n1190;
  assign new_n5936 = new_n3605 ^ new_n3466;
  assign new_n5937 = new_n5936 ^ new_n3460;
  assign new_n5938 = new_n5937 ^ new_n5935;
  assign new_n5939 = new_n3586 ^ new_n3559;
  assign new_n5940 = new_n5939 ^ new_n3550;
  assign new_n5941 = new_n3638 ^ new_n1163;
  assign new_n5942 = new_n3459 ^ new_n3389;
  assign new_n5943 = new_n5942 ^ new_n5941;
  assign new_n5944 = new_n5943 ^ new_n5940;
  assign new_n5945 = new_n5944 ^ new_n5938;
  assign new_n5946 = new_n3565 ^ new_n1174;
  assign new_n5947 = new_n5946 ^ new_n5942;
  assign new_n5948 = new_n3515 ^ new_n3506;
  assign new_n5949 = new_n5948 ^ new_n3587;
  assign new_n5950 = new_n5949 ^ new_n5947;
  assign new_n5951 = new_n3664 ^ new_n3265;
  assign new_n5952 = new_n5951 ^ new_n3154;
  assign new_n5953 = new_n3539 ^ new_n1182;
  assign new_n5954 = new_n5953 ^ new_n5942;
  assign new_n5955 = new_n5954 ^ new_n5952;
  assign new_n5956 = new_n5955 ^ new_n5950;
  assign new_n5957 = new_n5956 ^ new_n5945;
  assign new_n5958 = new_n3403 ^ new_n1154;
  assign new_n5959 = new_n5942 ^ new_n3667;
  assign new_n5960 = new_n5959 ^ new_n5958;
  assign new_n5961 = new_n5960 ^ new_n5957;
  assign new_n5962 = new_n3577 ^ new_n1201;
  assign new_n5963 = new_n3431 ^ new_n3042;
  assign new_n5964 = new_n5963 ^ new_n3507;
  assign new_n5965 = new_n5964 ^ new_n5962;
  assign new_n5966 = new_n5965 ^ new_n5956;
  assign new_n5967 = new_n3481 ^ new_n1118;
  assign new_n5968 = new_n3635 ^ new_n3610;
  assign new_n5969 = new_n5968 ^ new_n3606;
  assign new_n5970 = new_n5969 ^ new_n5967;
  assign new_n5971 = new_n5970 ^ new_n5966;
  assign new_n5972 = new_n5971 ^ new_n5960;
  assign new_n5973 = new_n3615 ^ new_n1141;
  assign new_n5974 = new_n3560 ^ new_n3549;
  assign new_n5975 = new_n5974 ^ new_n3636;
  assign new_n5976 = new_n5975 ^ new_n5973;
  assign new_n5977 = new_n5976 ^ new_n5970;
  assign new_n5978 = new_n5977 ^ new_n5960;
  assign new_n5979 = new_n5978 ^ new_n5938;
  assign new_n5980 = new_n5972 & new_n5979;
  assign new_n5981 = new_n5976 ^ new_n5966;
  assign new_n5982 = new_n5955 ^ new_n5938;
  assign new_n5983 = new_n5981 & new_n5982;
  assign new_n5984 = new_n5983 ^ new_n5980;
  assign new_n5985 = new_n5984 ^ new_n5938;
  assign new_n5986 = new_n5965 ^ new_n5938;
  assign new_n5987 = new_n5977 ^ new_n5957;
  assign new_n5988 = new_n5986 & new_n5987;
  assign new_n5989 = new_n5945 & new_n5971;
  assign new_n5990 = new_n5989 ^ new_n5988;
  assign new_n5991 = new_n5990 ^ new_n5981;
  assign new_n5992 = new_n5991 ^ new_n5985;
  assign new_n5993 = ~new_n5955 & ~new_n5978;
  assign new_n5994 = new_n5993 ^ new_n5955;
  assign new_n5995 = new_n5994 ^ new_n5983;
  assign new_n5996 = new_n5995 ^ new_n5986;
  assign new_n5997 = new_n5976 ^ new_n5944;
  assign new_n5998 = new_n5997 ^ new_n5986;
  assign new_n5999 = new_n5965 ^ new_n5944;
  assign new_n6000 = new_n5998 & new_n5999;
  assign new_n6001 = new_n6000 ^ new_n5989;
  assign new_n6002 = new_n5976 ^ new_n5950;
  assign new_n6003 = new_n6002 ^ new_n6001;
  assign new_n6004 = new_n6003 ^ new_n5996;
  assign new_n6005 = new_n5955 ^ new_n5944;
  assign new_n6006 = new_n6005 ^ new_n5986;
  assign new_n6007 = new_n5957 & new_n6006;
  assign new_n6008 = new_n6007 ^ new_n5970;
  assign new_n6009 = new_n6008 ^ new_n5957;
  assign new_n6010 = new_n5978 ^ new_n5955;
  assign new_n6011 = new_n6010 ^ new_n5986;
  assign new_n6012 = new_n5961 & new_n6011;
  assign new_n6013 = new_n6012 ^ new_n5989;
  assign new_n6014 = new_n6000 ^ new_n5965;
  assign new_n6015 = new_n6014 ^ new_n6013;
  assign new_n6016 = new_n6015 ^ new_n6009;
  assign new_n6017 = ~new_n6004 & new_n6016;
  assign new_n6018 = new_n6017 ^ new_n5992;
  assign new_n6019 = new_n5978 ^ new_n5944;
  assign new_n6020 = new_n5960 & new_n6019;
  assign new_n6021 = new_n6020 ^ new_n5944;
  assign new_n6022 = new_n6021 ^ new_n6008;
  assign new_n6023 = new_n6022 ^ new_n6017;
  assign new_n6024 = new_n6023 ^ new_n5991;
  assign new_n6025 = new_n6000 ^ new_n5988;
  assign new_n6026 = new_n5993 ^ new_n5980;
  assign new_n6027 = new_n6026 ^ new_n6025;
  assign new_n6028 = ~new_n6027 & new_n6024;
  assign new_n6029 = new_n6028 ^ new_n6017;
  assign new_n6030 = ~new_n5992 & ~new_n6029;
  assign new_n6031 = new_n6030 ^ new_n6028;
  assign new_n6032 = new_n6031 ^ new_n6018;
  assign new_n6033 = new_n6032 ^ new_n6028;
  assign new_n6034 = new_n6033 ^ new_n6027;
  assign new_n6035 = new_n5961 & new_n6034;
  assign new_n6036 = new_n6032 ^ new_n6004;
  assign new_n6037 = new_n5957 & new_n6036;
  assign new_n6038 = new_n6037 ^ new_n6035;
  assign new_n6039 = new_n6006 & new_n6036;
  assign new_n6040 = new_n6039 ^ new_n6038;
  assign new_n6041 = new_n5976 ^ new_n5938;
  assign new_n6042 = new_n6020 ^ new_n6012;
  assign new_n6043 = new_n6042 ^ new_n6025;
  assign new_n6044 = new_n6043 ^ new_n6041;
  assign new_n6045 = new_n6018 & new_n6044;
  assign new_n6046 = new_n6045 ^ new_n6022;
  assign new_n6047 = new_n6046 ^ new_n5991;
  assign new_n6048 = ~new_n6031 & new_n6047;
  assign new_n6049 = new_n6048 ^ new_n6045;
  assign new_n6050 = new_n6049 ^ new_n6016;
  assign new_n6051 = new_n5981 & new_n6050;
  assign new_n6052 = new_n6011 & new_n6034;
  assign new_n6053 = new_n6045 ^ new_n6028;
  assign new_n6054 = new_n6022 ^ new_n5985;
  assign new_n6055 = new_n6054 ^ new_n6053;
  assign new_n6056 = new_n5945 & new_n6055;
  assign new_n6057 = new_n5976 ^ new_n5955;
  assign new_n6058 = new_n6012 ^ new_n5994;
  assign new_n6059 = new_n6048 ^ new_n6032;
  assign new_n6060 = new_n6059 ^ new_n6058;
  assign new_n6061 = new_n6060 ^ new_n6057;
  assign new_n6062 = new_n6061 ^ new_n5944;
  assign new_n6063 = new_n6045 ^ new_n5983;
  assign new_n6064 = new_n6063 ^ new_n6008;
  assign new_n6065 = new_n6064 ^ new_n6062;
  assign new_n6066 = new_n5999 & new_n6065;
  assign new_n6067 = new_n6066 ^ new_n6056;
  assign new_n6068 = new_n6067 ^ new_n6052;
  assign new_n6069 = new_n6048 ^ new_n6044;
  assign new_n6070 = new_n5978 & new_n6069;
  assign new_n6071 = new_n6070 ^ new_n6068;
  assign new_n6072 = new_n6071 ^ new_n6051;
  assign new_n6073 = new_n6072 ^ new_n6040;
  assign new_n6074 = new_n6073 ^ new_n5934;
  assign new_n6075 = new_n3421 ^ n31;
  assign new_n6076 = new_n3594 ^ n29;
  assign new_n6077 = new_n6076 ^ new_n6075;
  assign new_n6078 = new_n3474 ^ n25;
  assign new_n6079 = new_n3553 ^ n28;
  assign new_n6080 = new_n6079 ^ new_n6078;
  assign new_n6081 = new_n6080 ^ new_n6077;
  assign new_n6082 = new_n3529 ^ n30;
  assign new_n6083 = new_n6082 ^ new_n6077;
  assign new_n6084 = new_n3621 ^ n26;
  assign new_n6085 = new_n6084 ^ new_n6083;
  assign new_n6086 = new_n6080 & new_n6085;
  assign new_n6087 = new_n6082 ^ new_n6078;
  assign new_n6088 = new_n3646 ^ n27;
  assign new_n6089 = new_n6088 ^ new_n6084;
  assign new_n6090 = new_n6089 ^ new_n6081;
  assign new_n6091 = ~new_n6090 & new_n6087;
  assign new_n6092 = new_n6091 ^ new_n6086;
  assign new_n6093 = new_n6088 ^ new_n6083;
  assign new_n6094 = new_n6093 ^ new_n6092;
  assign new_n6095 = new_n6078 ^ new_n6075;
  assign new_n6096 = ~new_n6095 & new_n6093;
  assign new_n6097 = new_n3661 ^ n32;
  assign new_n6098 = new_n6097 ^ new_n6089;
  assign new_n6099 = new_n6098 ^ new_n6078;
  assign new_n6100 = new_n6097 ^ new_n6085;
  assign new_n6101 = new_n6099 & new_n6100;
  assign new_n6102 = new_n6101 ^ new_n6096;
  assign new_n6103 = new_n6102 ^ new_n6078;
  assign new_n6104 = new_n6103 ^ new_n6094;
  assign new_n6105 = new_n6098 ^ new_n6079;
  assign new_n6106 = new_n6097 & new_n6105;
  assign new_n6107 = new_n6106 ^ new_n6079;
  assign new_n6108 = new_n6079 ^ new_n6075;
  assign new_n6109 = new_n6108 ^ new_n6087;
  assign new_n6110 = ~new_n6081 & ~new_n6109;
  assign new_n6111 = new_n6110 ^ new_n6084;
  assign new_n6112 = new_n6111 ^ new_n6107;
  assign new_n6113 = ~new_n6098 & new_n6075;
  assign new_n6114 = new_n6113 ^ new_n6075;
  assign new_n6115 = new_n6114 ^ new_n6096;
  assign new_n6116 = new_n6115 ^ new_n6087;
  assign new_n6117 = new_n6088 ^ new_n6079;
  assign new_n6118 = new_n6117 ^ new_n6087;
  assign new_n6119 = new_n6082 ^ new_n6079;
  assign new_n6120 = ~new_n6118 & new_n6119;
  assign new_n6121 = new_n6120 ^ new_n6086;
  assign new_n6122 = new_n6088 ^ new_n6076;
  assign new_n6123 = new_n6122 ^ new_n6121;
  assign new_n6124 = new_n6123 ^ new_n6116;
  assign new_n6125 = new_n6111 ^ new_n6081;
  assign new_n6126 = new_n6097 ^ new_n6081;
  assign new_n6127 = new_n6098 ^ new_n6075;
  assign new_n6128 = new_n6127 ^ new_n6087;
  assign new_n6129 = ~new_n6126 & ~new_n6128;
  assign new_n6130 = new_n6129 ^ new_n6082;
  assign new_n6131 = new_n6130 ^ new_n6121;
  assign new_n6132 = new_n6131 ^ new_n6125;
  assign new_n6133 = ~new_n6124 & new_n6132;
  assign new_n6134 = new_n6133 ^ new_n6112;
  assign new_n6135 = new_n6134 ^ new_n6094;
  assign new_n6136 = new_n6113 ^ new_n6101;
  assign new_n6137 = new_n6120 ^ new_n6091;
  assign new_n6138 = new_n6137 ^ new_n6136;
  assign new_n6139 = ~new_n6135 & ~new_n6138;
  assign new_n6140 = new_n6139 ^ new_n6133;
  assign new_n6141 = new_n6104 & new_n6140;
  assign new_n6142 = new_n6141 ^ new_n6124;
  assign new_n6143 = ~new_n6081 & ~new_n6142;
  assign new_n6144 = new_n6141 ^ new_n6139;
  assign new_n6145 = new_n6144 ^ new_n6138;
  assign new_n6146 = ~new_n6126 & ~new_n6145;
  assign new_n6147 = new_n6146 ^ new_n6143;
  assign new_n6148 = ~new_n6109 & ~new_n6142;
  assign new_n6149 = new_n6148 ^ new_n6147;
  assign new_n6150 = new_n6088 ^ new_n6078;
  assign new_n6151 = new_n6129 ^ new_n6106;
  assign new_n6152 = new_n6151 ^ new_n6137;
  assign new_n6153 = new_n6152 ^ new_n6150;
  assign new_n6154 = new_n6133 ^ new_n6104;
  assign new_n6155 = ~new_n6153 & new_n6154;
  assign new_n6156 = new_n6155 ^ new_n6112;
  assign new_n6157 = new_n6156 ^ new_n6094;
  assign new_n6158 = new_n6154 ^ new_n6141;
  assign new_n6159 = ~new_n6157 & new_n6158;
  assign new_n6160 = new_n6159 ^ new_n6155;
  assign new_n6161 = new_n6160 ^ new_n6132;
  assign new_n6162 = new_n6093 & new_n6161;
  assign new_n6163 = ~new_n6128 & ~new_n6145;
  assign new_n6164 = new_n6155 ^ new_n6139;
  assign new_n6165 = new_n6112 ^ new_n6103;
  assign new_n6166 = new_n6165 ^ new_n6164;
  assign new_n6167 = ~new_n6166 & new_n6080;
  assign new_n6168 = new_n6088 ^ new_n6075;
  assign new_n6169 = new_n6129 ^ new_n6114;
  assign new_n6170 = new_n6159 ^ new_n6141;
  assign new_n6171 = new_n6170 ^ new_n6169;
  assign new_n6172 = new_n6171 ^ new_n6168;
  assign new_n6173 = new_n6172 ^ new_n6079;
  assign new_n6174 = new_n6155 ^ new_n6096;
  assign new_n6175 = new_n6174 ^ new_n6111;
  assign new_n6176 = new_n6175 ^ new_n6173;
  assign new_n6177 = ~new_n6176 & new_n6119;
  assign new_n6178 = new_n6177 ^ new_n6167;
  assign new_n6179 = new_n6178 ^ new_n6163;
  assign new_n6180 = new_n6159 ^ new_n6153;
  assign new_n6181 = ~new_n6180 & new_n6098;
  assign new_n6182 = new_n6181 ^ new_n6179;
  assign new_n6183 = new_n6182 ^ new_n6162;
  assign new_n6184 = new_n6183 ^ new_n6149;
  assign new_n6185 = new_n6184 ^ new_n6074;
  assign new_n6186 = new_n5314 ^ new_n2076;
  assign new_n6187 = new_n6186 ^ new_n1991;
  assign new_n6188 = new_n2005 ^ new_n1928;
  assign new_n6189 = new_n6188 ^ new_n390;
  assign new_n6190 = new_n6189 ^ new_n6187;
  assign new_n6191 = new_n1991 ^ new_n370;
  assign new_n6192 = new_n6191 ^ new_n1894;
  assign new_n6193 = new_n2058 ^ n100;
  assign new_n6194 = new_n6193 ^ new_n5334;
  assign new_n6195 = new_n6194 ^ new_n6192;
  assign new_n6196 = new_n6195 ^ new_n6190;
  assign new_n6197 = new_n2015 ^ new_n1765;
  assign new_n6198 = new_n6197 ^ new_n2026;
  assign new_n6199 = new_n1947 ^ new_n1919;
  assign new_n6200 = new_n421 ^ n102;
  assign new_n6201 = new_n6200 ^ new_n6199;
  assign new_n6202 = new_n6201 ^ new_n6198;
  assign new_n6203 = new_n361 ^ n97;
  assign new_n6204 = new_n6203 ^ new_n2047;
  assign new_n6205 = new_n5322 ^ new_n1770;
  assign new_n6206 = new_n6205 ^ new_n6204;
  assign new_n6207 = new_n6206 ^ new_n6202;
  assign new_n6208 = new_n6207 ^ new_n6196;
  assign new_n6209 = new_n6206 ^ new_n6195;
  assign new_n6210 = new_n1955 ^ new_n1887;
  assign new_n6211 = new_n1514 ^ n101;
  assign new_n6212 = new_n6211 ^ new_n6210;
  assign new_n6213 = new_n1991 ^ new_n399;
  assign new_n6214 = new_n6213 ^ new_n2016;
  assign new_n6215 = new_n6214 ^ new_n6212;
  assign new_n6216 = new_n6215 ^ new_n6190;
  assign new_n6217 = new_n6216 ^ new_n6202;
  assign new_n6218 = new_n2033 ^ new_n430;
  assign new_n6219 = new_n2046 ^ new_n1982;
  assign new_n6220 = new_n6219 ^ new_n2064;
  assign new_n6221 = new_n6220 ^ new_n6218;
  assign new_n6222 = new_n6221 ^ new_n6217;
  assign new_n6223 = new_n6209 & new_n6222;
  assign new_n6224 = new_n6216 ^ new_n6209;
  assign new_n6225 = new_n2056 ^ new_n441;
  assign new_n6226 = new_n2063 ^ new_n2042;
  assign new_n6227 = new_n6226 ^ new_n1967;
  assign new_n6228 = new_n6227 ^ new_n6225;
  assign new_n6229 = new_n6228 ^ new_n6221;
  assign new_n6230 = new_n6229 ^ new_n6224;
  assign new_n6231 = new_n6207 & new_n6230;
  assign new_n6232 = new_n6231 ^ new_n6223;
  assign new_n6233 = new_n6228 ^ new_n6217;
  assign new_n6234 = new_n6233 ^ new_n6232;
  assign new_n6235 = new_n6206 ^ new_n6190;
  assign new_n6236 = new_n6233 & new_n6235;
  assign new_n6237 = new_n2076 ^ new_n410;
  assign new_n6238 = new_n2079 ^ new_n1926;
  assign new_n6239 = new_n6238 ^ new_n1991;
  assign new_n6240 = new_n6239 ^ new_n6237;
  assign new_n6241 = new_n6240 ^ new_n6222;
  assign new_n6242 = new_n6240 ^ new_n6229;
  assign new_n6243 = new_n6242 ^ new_n6206;
  assign new_n6244 = new_n6241 & new_n6243;
  assign new_n6245 = new_n6244 ^ new_n6236;
  assign new_n6246 = new_n6245 ^ new_n6206;
  assign new_n6247 = new_n6246 ^ new_n6234;
  assign new_n6248 = new_n6242 ^ new_n6195;
  assign new_n6249 = new_n6240 & new_n6248;
  assign new_n6250 = new_n6249 ^ new_n6195;
  assign new_n6251 = new_n6208 & new_n6224;
  assign new_n6252 = new_n6251 ^ new_n6221;
  assign new_n6253 = new_n6252 ^ new_n6250;
  assign new_n6254 = ~new_n6190 & ~new_n6242;
  assign new_n6255 = new_n6254 ^ new_n6190;
  assign new_n6256 = new_n6255 ^ new_n6236;
  assign new_n6257 = new_n6256 ^ new_n6207;
  assign new_n6258 = new_n6228 ^ new_n6195;
  assign new_n6259 = new_n6258 ^ new_n6207;
  assign new_n6260 = new_n6202 ^ new_n6195;
  assign new_n6261 = new_n6259 & new_n6260;
  assign new_n6262 = new_n6261 ^ new_n6223;
  assign new_n6263 = new_n6228 ^ new_n6215;
  assign new_n6264 = new_n6263 ^ new_n6262;
  assign new_n6265 = new_n6264 ^ new_n6257;
  assign new_n6266 = new_n6252 ^ new_n6224;
  assign new_n6267 = new_n6240 ^ new_n6224;
  assign new_n6268 = new_n6242 ^ new_n6190;
  assign new_n6269 = new_n6268 ^ new_n6207;
  assign new_n6270 = new_n6267 & new_n6269;
  assign new_n6271 = new_n6270 ^ new_n6262;
  assign new_n6272 = new_n6271 ^ new_n6202;
  assign new_n6273 = new_n6272 ^ new_n6266;
  assign new_n6274 = ~new_n6265 & new_n6273;
  assign new_n6275 = new_n6274 ^ new_n6253;
  assign new_n6276 = new_n6275 ^ new_n6234;
  assign new_n6277 = new_n6254 ^ new_n6244;
  assign new_n6278 = new_n6261 ^ new_n6231;
  assign new_n6279 = new_n6278 ^ new_n6277;
  assign new_n6280 = ~new_n6279 & new_n6276;
  assign new_n6281 = new_n6280 ^ new_n6274;
  assign new_n6282 = new_n6247 & new_n6281;
  assign new_n6283 = new_n6282 ^ new_n6265;
  assign new_n6284 = ~new_n6283 & new_n6208;
  assign new_n6285 = new_n6228 ^ new_n6206;
  assign new_n6286 = new_n6270 ^ new_n6249;
  assign new_n6287 = new_n6286 ^ new_n6278;
  assign new_n6288 = new_n6287 ^ new_n6285;
  assign new_n6289 = new_n6274 ^ new_n6247;
  assign new_n6290 = new_n6288 & new_n6289;
  assign new_n6291 = new_n6290 ^ new_n6280;
  assign new_n6292 = new_n6253 ^ new_n6246;
  assign new_n6293 = new_n6292 ^ new_n6291;
  assign new_n6294 = new_n6222 & new_n6293;
  assign new_n6295 = new_n6294 ^ new_n6284;
  assign new_n6296 = new_n6290 ^ new_n6253;
  assign new_n6297 = new_n6296 ^ new_n6234;
  assign new_n6298 = new_n6289 ^ new_n6282;
  assign new_n6299 = new_n6297 & new_n6298;
  assign new_n6300 = new_n6299 ^ new_n6290;
  assign new_n6301 = new_n6300 ^ new_n6273;
  assign new_n6302 = new_n6233 & new_n6301;
  assign new_n6303 = new_n6282 ^ new_n6280;
  assign new_n6304 = new_n6303 ^ new_n6279;
  assign new_n6305 = ~new_n6304 & new_n6269;
  assign new_n6306 = new_n6228 ^ new_n6190;
  assign new_n6307 = new_n6270 ^ new_n6255;
  assign new_n6308 = new_n6299 ^ new_n6282;
  assign new_n6309 = new_n6308 ^ new_n6307;
  assign new_n6310 = new_n6309 ^ new_n6306;
  assign new_n6311 = new_n6310 ^ new_n6195;
  assign new_n6312 = new_n6290 ^ new_n6236;
  assign new_n6313 = new_n6312 ^ new_n6252;
  assign new_n6314 = new_n6313 ^ new_n6311;
  assign new_n6315 = ~new_n6314 & new_n6260;
  assign new_n6316 = new_n6209 & new_n6293;
  assign new_n6317 = new_n6316 ^ new_n6315;
  assign new_n6318 = new_n6317 ^ new_n6305;
  assign new_n6319 = new_n6299 ^ new_n6288;
  assign new_n6320 = new_n6242 & new_n6319;
  assign new_n6321 = new_n6320 ^ new_n6318;
  assign new_n6322 = new_n6321 ^ new_n6302;
  assign new_n6323 = ~new_n6314 & new_n6259;
  assign new_n6324 = new_n6323 ^ new_n6322;
  assign new_n6325 = new_n6324 ^ new_n6295;
  assign new_n6326 = new_n4928 ^ new_n2759;
  assign new_n6327 = new_n3473 ^ new_n2748;
  assign new_n6328 = new_n6327 ^ new_n2797;
  assign new_n6329 = new_n6328 ^ new_n6326;
  assign new_n6330 = new_n4910 ^ new_n2655;
  assign new_n6331 = new_n2748 ^ new_n2618;
  assign new_n6332 = new_n6331 ^ new_n6330;
  assign new_n6333 = new_n3420 ^ new_n2395;
  assign new_n6334 = new_n6333 ^ new_n2838;
  assign new_n6335 = new_n6334 ^ new_n6332;
  assign new_n6336 = new_n6335 ^ new_n6329;
  assign new_n6337 = new_n4907 ^ new_n2647;
  assign new_n6338 = new_n3528 ^ new_n2781;
  assign new_n6339 = new_n6338 ^ new_n2395;
  assign new_n6340 = new_n6339 ^ new_n6337;
  assign new_n6341 = new_n4936 ^ new_n3552;
  assign new_n6342 = new_n6341 ^ new_n6331;
  assign new_n6343 = new_n2726 ^ new_n2709;
  assign new_n6344 = new_n6343 ^ new_n2673;
  assign new_n6345 = new_n6344 ^ new_n6342;
  assign new_n6346 = new_n6345 ^ new_n6340;
  assign new_n6347 = new_n6346 ^ new_n6336;
  assign new_n6348 = new_n3660 ^ new_n2838;
  assign new_n6349 = new_n6331 ^ new_n4933;
  assign new_n6350 = new_n6349 ^ new_n6348;
  assign new_n6351 = new_n4924 ^ new_n2821;
  assign new_n6352 = new_n2737 ^ new_n2726;
  assign new_n6353 = new_n6352 ^ new_n3645;
  assign new_n6354 = new_n6353 ^ new_n6351;
  assign new_n6355 = new_n4903 ^ new_n2808;
  assign new_n6356 = new_n3620 ^ new_n2797;
  assign new_n6357 = new_n6356 ^ new_n2821;
  assign new_n6358 = new_n6357 ^ new_n6355;
  assign new_n6359 = new_n6358 ^ new_n6354;
  assign new_n6360 = new_n6359 ^ new_n6350;
  assign new_n6361 = new_n6360 ^ new_n6329;
  assign new_n6362 = new_n2781 ^ new_n2709;
  assign new_n6363 = new_n6362 ^ new_n2680;
  assign new_n6364 = new_n4917 ^ new_n3593;
  assign new_n6365 = new_n6364 ^ new_n6331;
  assign new_n6366 = new_n6365 ^ new_n6363;
  assign new_n6367 = new_n6366 ^ new_n6335;
  assign new_n6368 = new_n6367 ^ new_n6340;
  assign new_n6369 = new_n6368 ^ new_n6358;
  assign new_n6370 = new_n6369 ^ new_n6350;
  assign new_n6371 = ~new_n6361 & ~new_n6370;
  assign new_n6372 = new_n6368 ^ new_n6354;
  assign new_n6373 = new_n6336 & new_n6372;
  assign new_n6374 = new_n6373 ^ new_n6371;
  assign new_n6375 = new_n6374 ^ new_n6329;
  assign new_n6376 = new_n6340 ^ new_n6329;
  assign new_n6377 = new_n6345 ^ new_n6329;
  assign new_n6378 = new_n6377 ^ new_n6367;
  assign new_n6379 = new_n6378 ^ new_n6359;
  assign new_n6380 = new_n6376 & new_n6379;
  assign new_n6381 = new_n6369 & new_n6377;
  assign new_n6382 = new_n6381 ^ new_n6380;
  assign new_n6383 = new_n6382 ^ new_n6372;
  assign new_n6384 = new_n6383 ^ new_n6375;
  assign new_n6385 = ~new_n6335 & new_n6360;
  assign new_n6386 = new_n6385 ^ new_n6335;
  assign new_n6387 = new_n6386 ^ new_n6373;
  assign new_n6388 = new_n6387 ^ new_n6376;
  assign new_n6389 = new_n6354 ^ new_n6345;
  assign new_n6390 = new_n6389 ^ new_n6376;
  assign new_n6391 = new_n6346 & new_n6390;
  assign new_n6392 = new_n6391 ^ new_n6381;
  assign new_n6393 = new_n6366 ^ new_n6354;
  assign new_n6394 = new_n6393 ^ new_n6392;
  assign new_n6395 = new_n6394 ^ new_n6388;
  assign new_n6396 = new_n6347 & new_n6378;
  assign new_n6397 = new_n6396 ^ new_n6358;
  assign new_n6398 = new_n6397 ^ new_n6378;
  assign new_n6399 = new_n6378 ^ new_n6350;
  assign new_n6400 = new_n6360 ^ new_n6335;
  assign new_n6401 = new_n6400 ^ new_n6376;
  assign new_n6402 = ~new_n6399 & ~new_n6401;
  assign new_n6403 = new_n6402 ^ new_n6392;
  assign new_n6404 = new_n6403 ^ new_n6340;
  assign new_n6405 = new_n6404 ^ new_n6398;
  assign new_n6406 = ~new_n6395 & new_n6405;
  assign new_n6407 = new_n6360 ^ new_n6345;
  assign new_n6408 = ~new_n6350 & ~new_n6407;
  assign new_n6409 = new_n6408 ^ new_n6345;
  assign new_n6410 = new_n6409 ^ new_n6397;
  assign new_n6411 = new_n6410 ^ new_n6406;
  assign new_n6412 = new_n6411 ^ new_n6383;
  assign new_n6413 = new_n6385 ^ new_n6371;
  assign new_n6414 = new_n6391 ^ new_n6380;
  assign new_n6415 = new_n6414 ^ new_n6413;
  assign new_n6416 = ~new_n6415 & new_n6412;
  assign new_n6417 = new_n6416 ^ new_n6406;
  assign new_n6418 = ~new_n6384 & ~new_n6417;
  assign new_n6419 = new_n6418 ^ new_n6416;
  assign new_n6420 = new_n6406 ^ new_n6384;
  assign new_n6421 = new_n6420 ^ new_n6419;
  assign new_n6422 = new_n6421 ^ new_n6395;
  assign new_n6423 = new_n6347 & new_n6422;
  assign new_n6424 = new_n6354 ^ new_n6329;
  assign new_n6425 = new_n6408 ^ new_n6402;
  assign new_n6426 = new_n6425 ^ new_n6414;
  assign new_n6427 = new_n6426 ^ new_n6424;
  assign new_n6428 = new_n6420 & new_n6427;
  assign new_n6429 = new_n6428 ^ new_n6416;
  assign new_n6430 = new_n6410 ^ new_n6375;
  assign new_n6431 = new_n6430 ^ new_n6429;
  assign new_n6432 = new_n6369 & new_n6431;
  assign new_n6433 = new_n6432 ^ new_n6423;
  assign new_n6434 = new_n6428 ^ new_n6410;
  assign new_n6435 = new_n6434 ^ new_n6383;
  assign new_n6436 = ~new_n6419 & new_n6435;
  assign new_n6437 = new_n6436 ^ new_n6428;
  assign new_n6438 = new_n6437 ^ new_n6405;
  assign new_n6439 = new_n6372 & new_n6438;
  assign new_n6440 = new_n6436 ^ new_n6427;
  assign new_n6441 = ~new_n6360 & new_n6440;
  assign new_n6442 = new_n6354 ^ new_n6335;
  assign new_n6443 = new_n6402 ^ new_n6386;
  assign new_n6444 = new_n6436 ^ new_n6421;
  assign new_n6445 = new_n6444 ^ new_n6443;
  assign new_n6446 = new_n6445 ^ new_n6442;
  assign new_n6447 = new_n6446 ^ new_n6345;
  assign new_n6448 = new_n6428 ^ new_n6373;
  assign new_n6449 = new_n6448 ^ new_n6397;
  assign new_n6450 = new_n6449 ^ new_n6447;
  assign new_n6451 = new_n6346 & new_n6450;
  assign new_n6452 = new_n6377 & new_n6431;
  assign new_n6453 = new_n6452 ^ new_n6451;
  assign new_n6454 = new_n6421 ^ new_n6416;
  assign new_n6455 = new_n6454 ^ new_n6415;
  assign new_n6456 = ~new_n6401 & new_n6455;
  assign new_n6457 = new_n6456 ^ new_n6453;
  assign new_n6458 = new_n6457 ^ new_n6441;
  assign new_n6459 = new_n6458 ^ new_n6439;
  assign new_n6460 = new_n6390 & new_n6450;
  assign new_n6461 = new_n6460 ^ new_n6459;
  assign new_n6462 = new_n6461 ^ new_n6433;
  assign new_n6463 = new_n6462 ^ new_n6325;
  assign new_n6464 = new_n6463 ^ new_n6185;
  assign new_n6465 = new_n6241 & new_n6297;
  assign new_n6466 = new_n6465 ^ new_n6284;
  assign new_n6467 = ~new_n6304 & new_n6267;
  assign new_n6468 = new_n6280 ^ new_n6247;
  assign new_n6469 = new_n6240 & new_n6468;
  assign new_n6470 = new_n6469 ^ new_n6467;
  assign new_n6471 = new_n6470 ^ new_n6321;
  assign new_n6472 = new_n6471 ^ new_n6466;
  assign new_n6473 = ~new_n6399 & new_n6455;
  assign new_n6474 = new_n6378 & new_n6422;
  assign new_n6475 = new_n6474 ^ new_n6473;
  assign new_n6476 = new_n6475 ^ new_n6423;
  assign new_n6477 = new_n6476 ^ new_n6459;
  assign new_n6478 = new_n6477 ^ new_n6472;
  assign new_n6479 = ~new_n6370 & new_n6435;
  assign new_n6480 = new_n6479 ^ new_n6423;
  assign new_n6481 = new_n6416 ^ new_n6384;
  assign new_n6482 = ~new_n6350 & new_n6481;
  assign new_n6483 = new_n6482 ^ new_n6473;
  assign new_n6484 = new_n6483 ^ new_n6458;
  assign new_n6485 = new_n6484 ^ new_n6480;
  assign new_n6486 = new_n6485 ^ n68;
  assign new_n6487 = new_n6486 ^ new_n6478;
  assign new_n6488 = new_n6487 ^ new_n6464;
  assign new_n6489 = ~new_n6283 & new_n6224;
  assign new_n6490 = new_n6489 ^ new_n6467;
  assign new_n6491 = new_n6490 ^ new_n6284;
  assign new_n6492 = new_n6491 ^ new_n6322;
  assign new_n6493 = new_n6492 ^ new_n6477;
  assign new_n6494 = new_n6493 ^ n67;
  assign new_n6495 = new_n5833 & new_n5916;
  assign new_n6496 = new_n6495 ^ new_n5917;
  assign new_n6497 = new_n5889 ^ new_n5801;
  assign new_n6498 = new_n5856 ^ new_n5851;
  assign new_n6499 = new_n6498 ^ new_n5922;
  assign new_n6500 = new_n6499 ^ new_n6497;
  assign new_n6501 = ~new_n6500 & new_n5835;
  assign new_n6502 = new_n5850 & new_n5907;
  assign new_n6503 = ~new_n6500 & new_n5841;
  assign new_n6504 = new_n6503 ^ new_n6502;
  assign new_n6505 = new_n5889 ^ new_n5854;
  assign new_n6506 = new_n5822 & new_n6505;
  assign new_n6507 = new_n6506 ^ new_n5896;
  assign new_n6508 = new_n5846 & new_n5911;
  assign new_n6509 = new_n6508 ^ new_n6507;
  assign new_n6510 = new_n6509 ^ new_n6504;
  assign new_n6511 = new_n6510 ^ new_n6501;
  assign new_n6512 = new_n6511 ^ new_n6496;
  assign new_n6513 = new_n5971 & new_n6055;
  assign new_n6514 = new_n6513 ^ new_n6056;
  assign new_n6515 = new_n6028 ^ new_n5938;
  assign new_n6516 = new_n6020 ^ new_n5980;
  assign new_n6517 = new_n6516 ^ new_n6061;
  assign new_n6518 = new_n6517 ^ new_n6515;
  assign new_n6519 = new_n5986 & new_n6518;
  assign new_n6520 = new_n5979 & new_n6047;
  assign new_n6521 = new_n5987 & new_n6518;
  assign new_n6522 = new_n6521 ^ new_n6520;
  assign new_n6523 = new_n6028 ^ new_n5992;
  assign new_n6524 = new_n5960 & new_n6523;
  assign new_n6525 = new_n6524 ^ new_n6037;
  assign new_n6526 = new_n5982 & new_n6050;
  assign new_n6527 = new_n6526 ^ new_n6525;
  assign new_n6528 = new_n6527 ^ new_n6522;
  assign new_n6529 = new_n6528 ^ new_n6519;
  assign new_n6530 = new_n6529 ^ new_n6514;
  assign new_n6531 = new_n6530 ^ new_n6512;
  assign new_n6532 = new_n6452 ^ new_n6432;
  assign new_n6533 = new_n6416 ^ new_n6329;
  assign new_n6534 = new_n6408 ^ new_n6371;
  assign new_n6535 = new_n6534 ^ new_n6446;
  assign new_n6536 = new_n6535 ^ new_n6533;
  assign new_n6537 = new_n6376 & new_n6536;
  assign new_n6538 = new_n6336 & new_n6438;
  assign new_n6539 = new_n6482 ^ new_n6474;
  assign new_n6540 = new_n6539 ^ new_n6538;
  assign new_n6541 = new_n6379 & new_n6536;
  assign new_n6542 = ~new_n6361 & new_n6435;
  assign new_n6543 = new_n6542 ^ new_n6541;
  assign new_n6544 = new_n6543 ^ new_n6540;
  assign new_n6545 = new_n6544 ^ new_n6537;
  assign new_n6546 = new_n6545 ^ new_n6532;
  assign new_n6547 = ~new_n6166 & new_n6085;
  assign new_n6548 = new_n6547 ^ new_n6167;
  assign new_n6549 = ~new_n6157 & new_n6099;
  assign new_n6550 = new_n6139 ^ new_n6078;
  assign new_n6551 = new_n6106 ^ new_n6101;
  assign new_n6552 = new_n6551 ^ new_n6172;
  assign new_n6553 = new_n6552 ^ new_n6550;
  assign new_n6554 = ~new_n6090 & new_n6553;
  assign new_n6555 = new_n6554 ^ new_n6549;
  assign new_n6556 = new_n6139 ^ new_n6104;
  assign new_n6557 = new_n6097 & new_n6556;
  assign new_n6558 = new_n6557 ^ new_n6143;
  assign new_n6559 = ~new_n6095 & new_n6161;
  assign new_n6560 = new_n6559 ^ new_n6558;
  assign new_n6561 = new_n6560 ^ new_n6555;
  assign new_n6562 = new_n6087 & new_n6553;
  assign new_n6563 = new_n6562 ^ new_n6561;
  assign new_n6564 = new_n6563 ^ new_n6548;
  assign new_n6565 = new_n6564 ^ new_n6546;
  assign new_n6566 = new_n6565 ^ new_n6531;
  assign new_n6567 = new_n6566 ^ new_n6494;
  assign new_n6568 = new_n6460 ^ new_n6432;
  assign new_n6569 = new_n6476 ^ new_n6457;
  assign new_n6570 = new_n6569 ^ new_n6568;
  assign new_n6571 = ~new_n6118 & ~new_n6176;
  assign new_n6572 = new_n6571 ^ new_n6547;
  assign new_n6573 = new_n6179 ^ new_n6149;
  assign new_n6574 = new_n6573 ^ new_n6572;
  assign new_n6575 = new_n6574 ^ n66;
  assign new_n6576 = new_n6575 ^ new_n6570;
  assign new_n6577 = new_n5998 & new_n6065;
  assign new_n6578 = new_n6577 ^ new_n6513;
  assign new_n6579 = new_n6068 ^ new_n6040;
  assign new_n6580 = new_n6579 ^ new_n6578;
  assign new_n6581 = ~new_n5926 & new_n5868;
  assign new_n6582 = new_n6581 ^ new_n6495;
  assign new_n6583 = new_n5929 ^ new_n5899;
  assign new_n6584 = new_n6583 ^ new_n6582;
  assign new_n6585 = new_n6584 ^ new_n6580;
  assign new_n6586 = new_n6316 ^ new_n6294;
  assign new_n6587 = new_n6280 ^ new_n6206;
  assign new_n6588 = new_n6249 ^ new_n6244;
  assign new_n6589 = new_n6588 ^ new_n6310;
  assign new_n6590 = new_n6589 ^ new_n6587;
  assign new_n6591 = ~new_n6590 & new_n6207;
  assign new_n6592 = new_n6489 ^ new_n6469;
  assign new_n6593 = new_n6235 & new_n6301;
  assign new_n6594 = new_n6593 ^ new_n6592;
  assign new_n6595 = new_n6243 & new_n6297;
  assign new_n6596 = ~new_n6590 & new_n6230;
  assign new_n6597 = new_n6596 ^ new_n6595;
  assign new_n6598 = new_n6597 ^ new_n6594;
  assign new_n6599 = new_n6598 ^ new_n6591;
  assign new_n6600 = new_n6599 ^ new_n6586;
  assign new_n6601 = new_n6600 ^ new_n6546;
  assign new_n6602 = new_n6601 ^ new_n6585;
  assign new_n6603 = new_n6602 ^ new_n6576;
  assign new_n6604 = new_n6603 ^ new_n6567;
  assign new_n6605 = new_n6527 ^ new_n6051;
  assign new_n6606 = new_n6010 & new_n6069;
  assign new_n6607 = new_n5972 & new_n6047;
  assign new_n6608 = new_n6607 ^ new_n6606;
  assign new_n6609 = new_n6608 ^ new_n6067;
  assign new_n6610 = new_n6609 ^ new_n6605;
  assign new_n6611 = new_n6509 ^ new_n5912;
  assign new_n6612 = new_n5876 & new_n5930;
  assign new_n6613 = new_n5848 & new_n5907;
  assign new_n6614 = new_n6613 ^ new_n6612;
  assign new_n6615 = new_n6614 ^ new_n5928;
  assign new_n6616 = new_n6615 ^ new_n6611;
  assign new_n6617 = new_n6616 ^ new_n6610;
  assign new_n6618 = new_n6617 ^ new_n6463;
  assign new_n6619 = new_n6540 ^ new_n6439;
  assign new_n6620 = ~new_n6400 & new_n6440;
  assign new_n6621 = new_n6620 ^ new_n6479;
  assign new_n6622 = new_n6621 ^ new_n6453;
  assign new_n6623 = new_n6622 ^ new_n6619;
  assign new_n6624 = new_n6560 ^ new_n6162;
  assign new_n6625 = ~new_n6127 & ~new_n6180;
  assign new_n6626 = ~new_n6157 & new_n6100;
  assign new_n6627 = new_n6626 ^ new_n6625;
  assign new_n6628 = new_n6627 ^ new_n6178;
  assign new_n6629 = new_n6628 ^ new_n6624;
  assign new_n6630 = new_n6629 ^ n72;
  assign new_n6631 = new_n6630 ^ new_n6623;
  assign new_n6632 = new_n6631 ^ new_n6618;
  assign new_n6633 = new_n6632 ^ new_n6604;
  assign new_n6634 = new_n6633 ^ new_n6488;
  assign new_n6635 = new_n6508 ^ new_n6503;
  assign new_n6636 = new_n6581 ^ new_n5931;
  assign new_n6637 = new_n6636 ^ new_n6615;
  assign new_n6638 = new_n6637 ^ new_n6635;
  assign new_n6639 = new_n6526 ^ new_n6521;
  assign new_n6640 = new_n6577 ^ new_n6070;
  assign new_n6641 = new_n6640 ^ new_n6609;
  assign new_n6642 = new_n6641 ^ new_n6639;
  assign new_n6643 = new_n6642 ^ new_n6638;
  assign new_n6644 = new_n6594 ^ new_n6302;
  assign new_n6645 = new_n6268 & new_n6319;
  assign new_n6646 = new_n6645 ^ new_n6465;
  assign new_n6647 = new_n6646 ^ new_n6317;
  assign new_n6648 = new_n6647 ^ new_n6644;
  assign new_n6649 = new_n6648 ^ new_n6463;
  assign new_n6650 = new_n6649 ^ new_n6643;
  assign new_n6651 = new_n6541 ^ new_n6538;
  assign new_n6652 = new_n6460 ^ new_n6441;
  assign new_n6653 = new_n6652 ^ new_n6622;
  assign new_n6654 = new_n6653 ^ new_n6651;
  assign new_n6655 = new_n6654 ^ new_n6623;
  assign new_n6656 = new_n6559 ^ new_n6554;
  assign new_n6657 = new_n6571 ^ new_n6181;
  assign new_n6658 = new_n6657 ^ new_n6628;
  assign new_n6659 = new_n6658 ^ new_n6656;
  assign new_n6660 = new_n6659 ^ n71;
  assign new_n6661 = new_n6660 ^ new_n6655;
  assign new_n6662 = new_n6661 ^ new_n6650;
  assign new_n6663 = ~new_n6633 & ~new_n6662;
  assign new_n6664 = new_n6663 ^ new_n6662;
  assign new_n6665 = new_n6495 ^ new_n5898;
  assign new_n6666 = new_n6581 ^ new_n5933;
  assign new_n6667 = new_n6666 ^ new_n6665;
  assign new_n6668 = new_n6513 ^ new_n6039;
  assign new_n6669 = new_n6577 ^ new_n6072;
  assign new_n6670 = new_n6669 ^ new_n6668;
  assign new_n6671 = new_n6670 ^ new_n6667;
  assign new_n6672 = new_n6323 ^ new_n6294;
  assign new_n6673 = new_n6491 ^ new_n6318;
  assign new_n6674 = new_n6673 ^ new_n6672;
  assign new_n6675 = new_n6674 ^ new_n6570;
  assign new_n6676 = new_n6675 ^ new_n6671;
  assign new_n6677 = new_n6571 ^ new_n6183;
  assign new_n6678 = new_n6547 ^ new_n6148;
  assign new_n6679 = new_n6678 ^ new_n6677;
  assign new_n6680 = new_n6679 ^ n65;
  assign new_n6681 = new_n6680 ^ new_n6462;
  assign new_n6682 = new_n6681 ^ new_n6676;
  assign new_n6683 = new_n6682 ^ new_n6662;
  assign new_n6684 = new_n6248 & new_n6468;
  assign new_n6685 = new_n6684 ^ new_n6324;
  assign new_n6686 = new_n6685 ^ new_n6598;
  assign new_n6687 = new_n6686 ^ new_n6485;
  assign new_n6688 = ~new_n6407 & new_n6481;
  assign new_n6689 = new_n6688 ^ new_n6461;
  assign new_n6690 = new_n6689 ^ new_n6544;
  assign new_n6691 = new_n6690 ^ n69;
  assign new_n6692 = new_n6691 ^ new_n6687;
  assign new_n6693 = new_n6607 ^ new_n6039;
  assign new_n6694 = new_n6524 ^ new_n6035;
  assign new_n6695 = new_n6694 ^ new_n6071;
  assign new_n6696 = new_n6695 ^ new_n6693;
  assign new_n6697 = new_n6613 ^ new_n5898;
  assign new_n6698 = new_n6506 ^ new_n5894;
  assign new_n6699 = new_n6698 ^ new_n5932;
  assign new_n6700 = new_n6699 ^ new_n6697;
  assign new_n6701 = new_n6700 ^ new_n6696;
  assign new_n6702 = new_n6626 ^ new_n6148;
  assign new_n6703 = new_n6557 ^ new_n6146;
  assign new_n6704 = new_n6703 ^ new_n6182;
  assign new_n6705 = new_n6704 ^ new_n6702;
  assign new_n6706 = new_n6705 ^ new_n6463;
  assign new_n6707 = new_n6706 ^ new_n6701;
  assign new_n6708 = new_n6707 ^ new_n6692;
  assign new_n6709 = new_n6708 ^ new_n6662;
  assign new_n6710 = new_n5855 & new_n6505;
  assign new_n6711 = new_n6710 ^ new_n6666;
  assign new_n6712 = new_n6711 ^ new_n6510;
  assign new_n6713 = new_n6019 & new_n6523;
  assign new_n6714 = new_n6713 ^ new_n6669;
  assign new_n6715 = new_n6714 ^ new_n6528;
  assign new_n6716 = new_n6715 ^ new_n6712;
  assign new_n6717 = new_n6596 ^ new_n6593;
  assign new_n6718 = new_n6323 ^ new_n6320;
  assign new_n6719 = new_n6718 ^ new_n6647;
  assign new_n6720 = new_n6719 ^ new_n6717;
  assign new_n6721 = new_n6720 ^ new_n6654;
  assign new_n6722 = new_n6721 ^ new_n6716;
  assign new_n6723 = new_n6105 & new_n6556;
  assign new_n6724 = new_n6723 ^ new_n6677;
  assign new_n6725 = new_n6724 ^ new_n6561;
  assign new_n6726 = new_n6725 ^ n70;
  assign new_n6727 = new_n6726 ^ new_n6690;
  assign new_n6728 = new_n6727 ^ new_n6722;
  assign new_n6729 = new_n6728 ^ new_n6709;
  assign new_n6730 = new_n6729 ^ new_n6567;
  assign new_n6731 = new_n6683 & new_n6730;
  assign new_n6732 = new_n6731 ^ new_n6664;
  assign new_n6733 = new_n6728 ^ new_n6682;
  assign new_n6734 = new_n6733 ^ new_n6732;
  assign new_n6735 = new_n6728 ^ new_n6488;
  assign new_n6736 = new_n6567 ^ new_n6488;
  assign new_n6737 = new_n6736 ^ new_n6733;
  assign new_n6738 = new_n6735 & new_n6737;
  assign new_n6739 = new_n6729 ^ new_n6603;
  assign new_n6740 = new_n6682 ^ new_n6488;
  assign new_n6741 = new_n6739 & new_n6740;
  assign new_n6742 = new_n6741 ^ new_n6738;
  assign new_n6743 = new_n6708 ^ new_n6567;
  assign new_n6744 = new_n6743 ^ new_n6742;
  assign new_n6745 = new_n6744 ^ new_n6734;
  assign new_n6746 = new_n6740 ^ new_n6709;
  assign new_n6747 = new_n6662 ^ new_n6488;
  assign new_n6748 = new_n6747 ^ new_n6733;
  assign new_n6749 = new_n6746 & new_n6748;
  assign new_n6750 = new_n6749 ^ new_n6603;
  assign new_n6751 = new_n6750 ^ new_n6746;
  assign new_n6752 = new_n6746 ^ new_n6632;
  assign new_n6753 = new_n6662 ^ new_n6633;
  assign new_n6754 = new_n6753 ^ new_n6733;
  assign new_n6755 = new_n6752 & new_n6754;
  assign new_n6756 = new_n6755 ^ new_n6742;
  assign new_n6757 = new_n6756 ^ new_n6728;
  assign new_n6758 = new_n6757 ^ new_n6751;
  assign new_n6759 = ~new_n6745 & new_n6758;
  assign new_n6760 = new_n6632 & new_n6634;
  assign new_n6761 = new_n6760 ^ new_n6488;
  assign new_n6762 = new_n6761 ^ new_n6750;
  assign new_n6763 = new_n6762 ^ new_n6759;
  assign new_n6764 = new_n6746 ^ new_n6604;
  assign new_n6765 = new_n6733 & new_n6764;
  assign new_n6766 = new_n6765 ^ new_n6741;
  assign new_n6767 = new_n6766 ^ new_n6730;
  assign new_n6768 = new_n6767 ^ new_n6763;
  assign new_n6769 = new_n6739 ^ new_n6632;
  assign new_n6770 = new_n6682 ^ new_n6633;
  assign new_n6771 = new_n6769 & new_n6770;
  assign new_n6772 = new_n6771 ^ new_n6663;
  assign new_n6773 = new_n6765 ^ new_n6738;
  assign new_n6774 = new_n6773 ^ new_n6772;
  assign new_n6775 = ~new_n6774 & new_n6768;
  assign new_n6776 = new_n6771 ^ new_n6731;
  assign new_n6777 = new_n6776 ^ new_n6682;
  assign new_n6778 = new_n6777 ^ new_n6767;
  assign new_n6779 = new_n6778 ^ new_n6775;
  assign new_n6780 = new_n6634 & new_n6779;
  assign new_n6781 = new_n6662 ^ new_n6567;
  assign new_n6782 = new_n6755 ^ new_n6664;
  assign new_n6783 = new_n6775 ^ new_n6759;
  assign new_n6784 = ~new_n6778 & ~new_n6783;
  assign new_n6785 = new_n6784 ^ new_n6775;
  assign new_n6786 = new_n6778 ^ new_n6759;
  assign new_n6787 = new_n6682 ^ new_n6567;
  assign new_n6788 = new_n6760 ^ new_n6755;
  assign new_n6789 = new_n6788 ^ new_n6773;
  assign new_n6790 = new_n6789 ^ new_n6787;
  assign new_n6791 = new_n6786 & new_n6790;
  assign new_n6792 = new_n6791 ^ new_n6762;
  assign new_n6793 = new_n6792 ^ new_n6767;
  assign new_n6794 = ~new_n6785 & new_n6793;
  assign new_n6795 = new_n6786 ^ new_n6785;
  assign new_n6796 = new_n6795 ^ new_n6794;
  assign new_n6797 = new_n6796 ^ new_n6782;
  assign new_n6798 = new_n6797 ^ new_n6781;
  assign new_n6799 = new_n6798 ^ new_n6488;
  assign new_n6800 = new_n6791 ^ new_n6731;
  assign new_n6801 = new_n6800 ^ new_n6750;
  assign new_n6802 = new_n6801 ^ new_n6799;
  assign new_n6803 = new_n6737 & new_n6802;
  assign new_n6804 = new_n6794 ^ new_n6790;
  assign new_n6805 = new_n6633 & new_n6804;
  assign new_n6806 = new_n6791 ^ new_n6775;
  assign new_n6807 = new_n6777 ^ new_n6762;
  assign new_n6808 = new_n6807 ^ new_n6806;
  assign new_n6809 = new_n6740 & new_n6808;
  assign new_n6810 = new_n6735 & new_n6802;
  assign new_n6811 = new_n6810 ^ new_n6809;
  assign new_n6812 = new_n6795 ^ new_n6775;
  assign new_n6813 = new_n6812 ^ new_n6774;
  assign new_n6814 = new_n6754 & new_n6813;
  assign new_n6815 = new_n6814 ^ new_n6811;
  assign new_n6816 = new_n6815 ^ new_n6805;
  assign new_n6817 = new_n6794 ^ new_n6791;
  assign new_n6818 = new_n6817 ^ new_n6758;
  assign new_n6819 = new_n6730 & new_n6818;
  assign new_n6820 = new_n6819 ^ new_n6816;
  assign new_n6821 = new_n6820 ^ new_n6803;
  assign new_n6822 = new_n6821 ^ new_n6780;
  assign new_n6823 = new_n6770 & new_n6793;
  assign new_n6824 = new_n6775 ^ new_n6682;
  assign new_n6825 = new_n6771 ^ new_n6760;
  assign new_n6826 = new_n6825 ^ new_n6798;
  assign new_n6827 = new_n6826 ^ new_n6824;
  assign new_n6828 = new_n6764 & new_n6827;
  assign new_n6829 = new_n6828 ^ new_n6823;
  assign new_n6830 = new_n6632 & new_n6779;
  assign new_n6831 = new_n6795 ^ new_n6745;
  assign new_n6832 = new_n6746 & new_n6831;
  assign new_n6833 = new_n6832 ^ new_n6830;
  assign new_n6834 = new_n6683 & new_n6818;
  assign new_n6835 = new_n6834 ^ new_n6833;
  assign new_n6836 = new_n6835 ^ new_n6829;
  assign new_n6837 = new_n6836 ^ new_n6822;
  assign new_n6838 = new_n6837 ^ new_n5797;
  assign new_n6839 = ~new_n970 & new_n922;
  assign new_n6840 = ~new_n906 & new_n1005;
  assign new_n6841 = new_n6840 ^ new_n6839;
  assign new_n6842 = new_n6841 ^ new_n995;
  assign new_n6843 = new_n6842 ^ n81;
  assign new_n6844 = new_n6843 ^ n17;
  assign new_n6845 = new_n5808 ^ new_n4282;
  assign new_n6846 = new_n6082 ^ new_n4011;
  assign new_n6847 = new_n6846 ^ new_n4326;
  assign new_n6848 = new_n6847 ^ new_n6845;
  assign new_n6849 = new_n5799 ^ new_n4402;
  assign new_n6850 = new_n6849 ^ new_n5825;
  assign new_n6851 = new_n6075 ^ new_n4326;
  assign new_n6852 = new_n6851 ^ new_n4249;
  assign new_n6853 = new_n6852 ^ new_n6850;
  assign new_n6854 = new_n4386 ^ new_n4309;
  assign new_n6855 = new_n6854 ^ new_n4011;
  assign new_n6856 = new_n6076 ^ new_n5802;
  assign new_n6857 = new_n6856 ^ new_n5799;
  assign new_n6858 = new_n6857 ^ new_n6855;
  assign new_n6859 = new_n6858 ^ new_n6853;
  assign new_n6860 = new_n6859 ^ new_n6848;
  assign new_n6861 = new_n4409 ^ new_n4359;
  assign new_n6862 = new_n6084 ^ new_n4371;
  assign new_n6863 = new_n6862 ^ new_n4346;
  assign new_n6864 = new_n6863 ^ new_n6861;
  assign new_n6865 = new_n6864 ^ new_n6860;
  assign new_n6866 = new_n4375 ^ new_n4337;
  assign new_n6867 = new_n6078 ^ new_n4016;
  assign new_n6868 = new_n6867 ^ new_n4371;
  assign new_n6869 = new_n6868 ^ new_n6866;
  assign new_n6870 = new_n4417 ^ new_n4346;
  assign new_n6871 = new_n4411 ^ new_n4388;
  assign new_n6872 = new_n6871 ^ new_n6088;
  assign new_n6873 = new_n6872 ^ new_n6870;
  assign new_n6874 = new_n6873 ^ new_n6869;
  assign new_n6875 = new_n6079 ^ new_n5799;
  assign new_n6876 = new_n6875 ^ new_n4381;
  assign new_n6877 = new_n4411 ^ new_n4130;
  assign new_n6878 = new_n6877 ^ new_n4386;
  assign new_n6879 = new_n6878 ^ new_n6876;
  assign new_n6880 = new_n6879 ^ new_n6869;
  assign new_n6881 = new_n6880 ^ new_n6859;
  assign new_n6882 = new_n6097 ^ new_n4249;
  assign new_n6883 = new_n5814 ^ new_n5799;
  assign new_n6884 = new_n6883 ^ new_n6882;
  assign new_n6885 = new_n6884 ^ new_n6881;
  assign new_n6886 = new_n6873 ^ new_n6864;
  assign new_n6887 = new_n6886 ^ new_n6884;
  assign new_n6888 = new_n6887 ^ new_n6853;
  assign new_n6889 = new_n6869 ^ new_n6848;
  assign new_n6890 = new_n6889 ^ new_n6888;
  assign new_n6891 = ~new_n6885 & ~new_n6890;
  assign new_n6892 = new_n6887 ^ new_n6879;
  assign new_n6893 = ~new_n6884 & ~new_n6892;
  assign new_n6894 = new_n6893 ^ new_n6891;
  assign new_n6895 = new_n6886 ^ new_n6881;
  assign new_n6896 = new_n6889 & new_n6895;
  assign new_n6897 = new_n6879 ^ new_n6848;
  assign new_n6898 = new_n6879 ^ new_n6873;
  assign new_n6899 = new_n6898 ^ new_n6889;
  assign new_n6900 = new_n6897 & new_n6899;
  assign new_n6901 = new_n6900 ^ new_n6896;
  assign new_n6902 = new_n6901 ^ new_n6894;
  assign new_n6903 = new_n6902 ^ new_n6874;
  assign new_n6904 = new_n6884 ^ new_n6865;
  assign new_n6905 = new_n6887 ^ new_n6869;
  assign new_n6906 = ~new_n6904 & ~new_n6905;
  assign new_n6907 = new_n6869 ^ new_n6853;
  assign new_n6908 = new_n6873 ^ new_n6860;
  assign new_n6909 = new_n6907 & new_n6908;
  assign new_n6910 = new_n6909 ^ new_n6906;
  assign new_n6911 = new_n6910 ^ new_n6869;
  assign new_n6912 = new_n6865 & new_n6880;
  assign new_n6913 = new_n6912 ^ new_n6896;
  assign new_n6914 = new_n6913 ^ new_n6908;
  assign new_n6915 = new_n6914 ^ new_n6911;
  assign new_n6916 = ~new_n6853 & new_n6887;
  assign new_n6917 = new_n6916 ^ new_n6853;
  assign new_n6918 = new_n6917 ^ new_n6909;
  assign new_n6919 = new_n6918 ^ new_n6889;
  assign new_n6920 = new_n6912 ^ new_n6900;
  assign new_n6921 = new_n6873 ^ new_n6858;
  assign new_n6922 = new_n6921 ^ new_n6920;
  assign new_n6923 = new_n6922 ^ new_n6919;
  assign new_n6924 = new_n6907 ^ new_n6897;
  assign new_n6925 = new_n6881 & new_n6924;
  assign new_n6926 = new_n6925 ^ new_n6864;
  assign new_n6927 = new_n6926 ^ new_n6881;
  assign new_n6928 = new_n6912 ^ new_n6891;
  assign new_n6929 = new_n6900 ^ new_n6848;
  assign new_n6930 = new_n6929 ^ new_n6928;
  assign new_n6931 = new_n6930 ^ new_n6927;
  assign new_n6932 = ~new_n6923 & new_n6931;
  assign new_n6933 = new_n6932 ^ new_n6915;
  assign new_n6934 = new_n6903 & new_n6933;
  assign new_n6935 = new_n6893 ^ new_n6879;
  assign new_n6936 = new_n6935 ^ new_n6926;
  assign new_n6937 = new_n6936 ^ new_n6932;
  assign new_n6938 = new_n6937 ^ new_n6914;
  assign new_n6939 = new_n6916 ^ new_n6906;
  assign new_n6940 = new_n6939 ^ new_n6901;
  assign new_n6941 = ~new_n6940 & new_n6938;
  assign new_n6942 = new_n6941 ^ new_n6934;
  assign new_n6943 = new_n6936 ^ new_n6911;
  assign new_n6944 = new_n6943 ^ new_n6942;
  assign new_n6945 = new_n6865 & new_n6944;
  assign new_n6946 = new_n6941 ^ new_n6932;
  assign new_n6947 = ~new_n6946 & new_n6915;
  assign new_n6948 = new_n6947 ^ new_n6915;
  assign new_n6949 = new_n6948 ^ new_n6923;
  assign new_n6950 = ~new_n6949 & new_n6924;
  assign new_n6951 = new_n6950 ^ new_n6945;
  assign new_n6952 = new_n6936 ^ new_n6934;
  assign new_n6953 = new_n6952 ^ new_n6914;
  assign new_n6954 = new_n6947 ^ new_n6932;
  assign new_n6955 = new_n6953 & new_n6954;
  assign new_n6956 = new_n6955 ^ new_n6903;
  assign new_n6957 = ~new_n6887 & new_n6956;
  assign new_n6958 = new_n6948 ^ new_n6941;
  assign new_n6959 = new_n6958 ^ new_n6940;
  assign new_n6960 = ~new_n6890 & ~new_n6959;
  assign new_n6961 = new_n6880 & new_n6944;
  assign new_n6962 = new_n6873 ^ new_n6853;
  assign new_n6963 = new_n6917 ^ new_n6891;
  assign new_n6964 = new_n6955 ^ new_n6948;
  assign new_n6965 = new_n6964 ^ new_n6963;
  assign new_n6966 = new_n6965 ^ new_n6962;
  assign new_n6967 = new_n6966 ^ new_n6879;
  assign new_n6968 = new_n6934 ^ new_n6909;
  assign new_n6969 = new_n6968 ^ new_n6926;
  assign new_n6970 = new_n6969 ^ new_n6967;
  assign new_n6971 = ~new_n6970 & new_n6897;
  assign new_n6972 = new_n6971 ^ new_n6961;
  assign new_n6973 = new_n6972 ^ new_n6960;
  assign new_n6974 = new_n6973 ^ new_n6957;
  assign new_n6975 = new_n6955 ^ new_n6934;
  assign new_n6976 = new_n6975 ^ new_n6931;
  assign new_n6977 = new_n6908 & new_n6976;
  assign new_n6978 = new_n6977 ^ new_n6974;
  assign new_n6979 = ~new_n6970 & new_n6899;
  assign new_n6980 = new_n6979 ^ new_n6978;
  assign new_n6981 = new_n6980 ^ new_n6951;
  assign new_n6982 = new_n6981 ^ new_n6844;
  assign new_n6983 = new_n2781 ^ new_n2668;
  assign new_n6984 = new_n6983 ^ new_n2680;
  assign new_n6985 = new_n4910 ^ new_n902;
  assign new_n6986 = new_n6985 ^ new_n6984;
  assign new_n6987 = new_n4928 ^ new_n2786;
  assign new_n6988 = new_n6987 ^ new_n4933;
  assign new_n6989 = new_n2395 ^ new_n891;
  assign new_n6990 = new_n6989 ^ new_n2647;
  assign new_n6991 = new_n6990 ^ new_n6988;
  assign new_n6992 = new_n2734 ^ new_n2709;
  assign new_n6993 = new_n6992 ^ new_n2673;
  assign new_n6994 = new_n4928 ^ new_n883;
  assign new_n6995 = new_n6994 ^ new_n4907;
  assign new_n6996 = new_n6995 ^ new_n6993;
  assign new_n6997 = new_n6996 ^ new_n6991;
  assign new_n6998 = new_n6997 ^ new_n6986;
  assign new_n6999 = new_n4924 ^ new_n2754;
  assign new_n7000 = new_n2797 ^ new_n819;
  assign new_n7001 = new_n7000 ^ new_n2759;
  assign new_n7002 = new_n7001 ^ new_n6999;
  assign new_n7003 = new_n7002 ^ new_n6998;
  assign new_n7004 = new_n4903 ^ new_n874;
  assign new_n7005 = new_n2748 ^ new_n2619;
  assign new_n7006 = new_n7005 ^ new_n7004;
  assign new_n7007 = new_n7006 ^ new_n6991;
  assign new_n7008 = new_n4936 ^ new_n2802;
  assign new_n7009 = new_n2821 ^ new_n842;
  assign new_n7010 = new_n7009 ^ new_n2808;
  assign new_n7011 = new_n7010 ^ new_n7008;
  assign new_n7012 = new_n7011 ^ new_n6998;
  assign new_n7013 = new_n7007 & new_n7012;
  assign new_n7014 = new_n4928 ^ new_n2631;
  assign new_n7015 = new_n2838 ^ new_n855;
  assign new_n7016 = new_n7015 ^ new_n2655;
  assign new_n7017 = new_n7016 ^ new_n7014;
  assign new_n7018 = new_n7011 ^ new_n7002;
  assign new_n7019 = new_n7018 ^ new_n7017;
  assign new_n7020 = ~new_n6991 & ~new_n7019;
  assign new_n7021 = new_n7020 ^ new_n6991;
  assign new_n7022 = new_n7021 ^ new_n7013;
  assign new_n7023 = new_n7006 ^ new_n6986;
  assign new_n7024 = new_n7023 ^ new_n7022;
  assign new_n7025 = new_n4928 ^ new_n864;
  assign new_n7026 = new_n7025 ^ new_n4917;
  assign new_n7027 = new_n2825 ^ new_n2726;
  assign new_n7028 = new_n7027 ^ new_n7026;
  assign new_n7029 = new_n7028 ^ new_n7006;
  assign new_n7030 = new_n7003 & new_n7029;
  assign new_n7031 = new_n7028 ^ new_n6986;
  assign new_n7032 = new_n7028 ^ new_n7011;
  assign new_n7033 = new_n7032 ^ new_n7023;
  assign new_n7034 = new_n7031 & new_n7033;
  assign new_n7035 = new_n7034 ^ new_n7030;
  assign new_n7036 = new_n7011 ^ new_n6996;
  assign new_n7037 = new_n7036 ^ new_n7035;
  assign new_n7038 = new_n7037 ^ new_n7024;
  assign new_n7039 = new_n7029 ^ new_n6997;
  assign new_n7040 = new_n7031 ^ new_n7007;
  assign new_n7041 = new_n7039 & new_n7040;
  assign new_n7042 = new_n7041 ^ new_n7002;
  assign new_n7043 = new_n7042 ^ new_n7039;
  assign new_n7044 = new_n7039 ^ new_n7017;
  assign new_n7045 = new_n7019 ^ new_n6991;
  assign new_n7046 = new_n7045 ^ new_n7023;
  assign new_n7047 = new_n7044 & new_n7046;
  assign new_n7048 = new_n7047 ^ new_n7035;
  assign new_n7049 = new_n7048 ^ new_n6986;
  assign new_n7050 = new_n7049 ^ new_n7043;
  assign new_n7051 = ~new_n7038 & new_n7050;
  assign new_n7052 = new_n7028 ^ new_n7019;
  assign new_n7053 = new_n7017 & new_n7052;
  assign new_n7054 = new_n7053 ^ new_n7028;
  assign new_n7055 = new_n7054 ^ new_n7042;
  assign new_n7056 = new_n7055 ^ new_n7051;
  assign new_n7057 = new_n7039 ^ new_n7018;
  assign new_n7058 = new_n7023 & new_n7057;
  assign new_n7059 = new_n7058 ^ new_n7030;
  assign new_n7060 = new_n7059 ^ new_n7012;
  assign new_n7061 = new_n7060 ^ new_n7056;
  assign new_n7062 = new_n7017 ^ new_n7003;
  assign new_n7063 = new_n7019 ^ new_n7006;
  assign new_n7064 = new_n7062 & new_n7063;
  assign new_n7065 = new_n7064 ^ new_n7020;
  assign new_n7066 = new_n7058 ^ new_n7034;
  assign new_n7067 = new_n7066 ^ new_n7065;
  assign new_n7068 = ~new_n7067 & new_n7061;
  assign new_n7069 = new_n7011 ^ new_n7006;
  assign new_n7070 = new_n7053 ^ new_n7047;
  assign new_n7071 = new_n7070 ^ new_n7066;
  assign new_n7072 = new_n7071 ^ new_n7069;
  assign new_n7073 = new_n7064 ^ new_n7013;
  assign new_n7074 = new_n7073 ^ new_n7006;
  assign new_n7075 = new_n7074 ^ new_n7060;
  assign new_n7076 = new_n7075 ^ new_n7051;
  assign new_n7077 = new_n7072 & new_n7076;
  assign new_n7078 = new_n7077 ^ new_n7068;
  assign new_n7079 = new_n7074 ^ new_n7055;
  assign new_n7080 = new_n7079 ^ new_n7078;
  assign new_n7081 = new_n7003 & new_n7080;
  assign new_n7082 = new_n7011 ^ new_n6991;
  assign new_n7083 = new_n7047 ^ new_n7021;
  assign new_n7084 = new_n7077 ^ new_n7055;
  assign new_n7085 = new_n7084 ^ new_n7060;
  assign new_n7086 = new_n7068 ^ new_n7051;
  assign new_n7087 = new_n7075 & new_n7086;
  assign new_n7088 = new_n7087 ^ new_n7076;
  assign new_n7089 = new_n7085 & new_n7088;
  assign new_n7090 = new_n7089 ^ new_n7087;
  assign new_n7091 = new_n7090 ^ new_n7083;
  assign new_n7092 = new_n7091 ^ new_n7082;
  assign new_n7093 = new_n7092 ^ new_n7028;
  assign new_n7094 = new_n7077 ^ new_n7013;
  assign new_n7095 = new_n7094 ^ new_n7042;
  assign new_n7096 = new_n7095 ^ new_n7093;
  assign new_n7097 = ~new_n7096 & new_n7033;
  assign new_n7098 = new_n7097 ^ new_n7081;
  assign new_n7099 = new_n7087 ^ new_n7068;
  assign new_n7100 = new_n7099 ^ new_n7067;
  assign new_n7101 = ~new_n7100 & new_n7044;
  assign new_n7102 = new_n7087 ^ new_n7038;
  assign new_n7103 = ~new_n7102 & new_n7039;
  assign new_n7104 = new_n7103 ^ new_n7101;
  assign new_n7105 = ~new_n7102 & new_n7040;
  assign new_n7106 = new_n7105 ^ new_n7104;
  assign new_n7107 = ~new_n7100 & new_n7046;
  assign new_n7108 = new_n7029 & new_n7080;
  assign new_n7109 = ~new_n7096 & new_n7031;
  assign new_n7110 = new_n7109 ^ new_n7108;
  assign new_n7111 = new_n7110 ^ new_n7107;
  assign new_n7112 = new_n7111 ^ new_n7106;
  assign new_n7113 = new_n7112 ^ new_n7098;
  assign new_n7114 = new_n2058 ^ new_n1974;
  assign new_n7115 = new_n7114 ^ n115;
  assign new_n7116 = new_n2042 ^ new_n1138;
  assign new_n7117 = new_n7116 ^ new_n2064;
  assign new_n7118 = new_n7117 ^ new_n7115;
  assign new_n7119 = new_n1996 ^ new_n1770;
  assign new_n7120 = new_n7119 ^ new_n1160;
  assign new_n7121 = new_n7120 ^ new_n1967;
  assign new_n7122 = new_n2058 ^ new_n1955;
  assign new_n7123 = new_n1514 ^ n116;
  assign new_n7124 = new_n7123 ^ new_n7122;
  assign new_n7125 = new_n7124 ^ new_n7121;
  assign new_n7126 = new_n7125 ^ new_n7118;
  assign new_n7127 = new_n2005 ^ new_n1912;
  assign new_n7128 = new_n7127 ^ new_n2016;
  assign new_n7129 = new_n1765 ^ n118;
  assign new_n7130 = new_n7129 ^ new_n1198;
  assign new_n7131 = new_n7130 ^ new_n7128;
  assign new_n7132 = new_n2033 ^ new_n1982;
  assign new_n7133 = new_n7132 ^ new_n1991;
  assign new_n7134 = new_n1770 ^ n113;
  assign new_n7135 = new_n7134 ^ new_n1187;
  assign new_n7136 = new_n7135 ^ new_n7133;
  assign new_n7137 = new_n7136 ^ new_n7131;
  assign new_n7138 = new_n7137 ^ new_n7126;
  assign new_n7139 = new_n6238 ^ new_n6199;
  assign new_n7140 = new_n7139 ^ new_n7119;
  assign new_n7141 = new_n2005 ^ new_n1180;
  assign new_n7142 = new_n7141 ^ new_n7140;
  assign new_n7143 = new_n7142 ^ new_n7118;
  assign new_n7144 = new_n7136 ^ new_n7125;
  assign new_n7145 = new_n1955 ^ new_n1765;
  assign new_n7146 = new_n2026 ^ n117;
  assign new_n7147 = new_n7146 ^ new_n7145;
  assign new_n7148 = new_n7119 ^ new_n1171;
  assign new_n7149 = new_n7148 ^ new_n1894;
  assign new_n7150 = new_n7149 ^ new_n7147;
  assign new_n7151 = new_n7150 ^ new_n7142;
  assign new_n7152 = new_n7151 ^ new_n7144;
  assign new_n7153 = new_n2076 ^ new_n1152;
  assign new_n7154 = new_n7119 ^ new_n1929;
  assign new_n7155 = new_n7154 ^ new_n7153;
  assign new_n7156 = new_n7155 ^ new_n7152;
  assign new_n7157 = new_n2056 ^ new_n1116;
  assign new_n7158 = new_n2042 ^ new_n1982;
  assign new_n7159 = new_n7158 ^ new_n2047;
  assign new_n7160 = new_n7159 ^ new_n7157;
  assign new_n7161 = new_n7160 ^ new_n7118;
  assign new_n7162 = new_n7161 ^ new_n7155;
  assign new_n7163 = new_n7162 ^ new_n7142;
  assign new_n7164 = new_n7163 ^ new_n7137;
  assign new_n7165 = new_n7156 & new_n7164;
  assign new_n7166 = ~new_n7142 & ~new_n7162;
  assign new_n7167 = new_n7166 ^ new_n7142;
  assign new_n7168 = new_n7167 ^ new_n7165;
  assign new_n7169 = new_n7136 ^ new_n7118;
  assign new_n7170 = ~new_n7161 & new_n7155;
  assign new_n7171 = ~new_n7155 & new_n7125;
  assign new_n7172 = new_n7171 ^ new_n7170;
  assign new_n7173 = new_n7172 ^ new_n7125;
  assign new_n7174 = new_n7173 ^ new_n7165;
  assign new_n7175 = new_n7131 ^ new_n7125;
  assign new_n7176 = new_n7138 & new_n7175;
  assign new_n7177 = new_n7161 ^ new_n7152;
  assign new_n7178 = new_n7137 & new_n7177;
  assign new_n7179 = new_n7178 ^ new_n7176;
  assign new_n7180 = new_n7179 ^ new_n7174;
  assign new_n7181 = new_n7180 ^ new_n7169;
  assign new_n7182 = new_n7151 ^ new_n7131;
  assign new_n7183 = new_n7182 ^ new_n7118;
  assign new_n7184 = new_n7142 ^ new_n7136;
  assign new_n7185 = new_n7183 & new_n7184;
  assign new_n7186 = new_n7185 ^ new_n7167;
  assign new_n7187 = new_n7186 ^ new_n7137;
  assign new_n7188 = new_n7182 ^ new_n7160;
  assign new_n7189 = new_n7144 & new_n7188;
  assign new_n7190 = new_n7189 ^ new_n7176;
  assign new_n7191 = new_n7150 ^ new_n7118;
  assign new_n7192 = new_n7191 ^ new_n7190;
  assign new_n7193 = new_n7192 ^ new_n7187;
  assign new_n7194 = new_n7142 ^ new_n7125;
  assign new_n7195 = new_n7194 ^ new_n7137;
  assign new_n7196 = new_n7152 & new_n7195;
  assign new_n7197 = new_n7196 ^ new_n7160;
  assign new_n7198 = new_n7197 ^ new_n7152;
  assign new_n7199 = new_n7190 ^ new_n7165;
  assign new_n7200 = new_n7199 ^ new_n7131;
  assign new_n7201 = new_n7200 ^ new_n7198;
  assign new_n7202 = ~new_n7193 & new_n7201;
  assign new_n7203 = new_n7189 ^ new_n7178;
  assign new_n7204 = new_n7203 ^ new_n7183;
  assign new_n7205 = new_n7162 ^ new_n7136;
  assign new_n7206 = new_n7188 ^ new_n7155;
  assign new_n7207 = new_n7205 & new_n7206;
  assign new_n7208 = new_n7207 ^ new_n7185;
  assign new_n7209 = new_n7208 ^ new_n7136;
  assign new_n7210 = new_n7209 ^ new_n7204;
  assign new_n7211 = new_n7210 ^ new_n7202;
  assign new_n7212 = new_n7181 & new_n7211;
  assign new_n7213 = new_n7197 ^ new_n7172;
  assign new_n7214 = new_n7213 ^ new_n7212;
  assign new_n7215 = new_n7214 ^ new_n7204;
  assign new_n7216 = new_n7213 ^ new_n7202;
  assign new_n7217 = new_n7216 ^ new_n7204;
  assign new_n7218 = new_n7207 ^ new_n7166;
  assign new_n7219 = new_n7218 ^ new_n7179;
  assign new_n7220 = ~new_n7219 & new_n7217;
  assign new_n7221 = new_n7220 ^ new_n7202;
  assign new_n7222 = new_n7210 & new_n7221;
  assign new_n7223 = new_n7222 ^ new_n7211;
  assign new_n7224 = new_n7215 & new_n7223;
  assign new_n7225 = new_n7224 ^ new_n7222;
  assign new_n7226 = new_n7225 ^ new_n7168;
  assign new_n7227 = new_n7226 ^ new_n7143;
  assign new_n7228 = new_n7227 ^ new_n7125;
  assign new_n7229 = new_n7212 ^ new_n7185;
  assign new_n7230 = new_n7229 ^ new_n7197;
  assign new_n7231 = new_n7230 ^ new_n7228;
  assign new_n7232 = ~new_n7231 & new_n7138;
  assign new_n7233 = new_n7220 ^ new_n7212;
  assign new_n7234 = new_n7213 ^ new_n7209;
  assign new_n7235 = new_n7234 ^ new_n7233;
  assign new_n7236 = new_n7188 & new_n7235;
  assign new_n7237 = new_n7236 ^ new_n7232;
  assign new_n7238 = new_n7222 ^ new_n7220;
  assign new_n7239 = new_n7238 ^ new_n7219;
  assign new_n7240 = ~new_n7239 & new_n7156;
  assign new_n7241 = new_n7222 ^ new_n7193;
  assign new_n7242 = ~new_n7241 & new_n7152;
  assign new_n7243 = new_n7242 ^ new_n7240;
  assign new_n7244 = ~new_n7241 & new_n7195;
  assign new_n7245 = new_n7244 ^ new_n7243;
  assign new_n7246 = new_n7144 & new_n7235;
  assign new_n7247 = ~new_n7231 & new_n7175;
  assign new_n7248 = new_n7247 ^ new_n7246;
  assign new_n7249 = ~new_n7239 & new_n7164;
  assign new_n7250 = new_n7249 ^ new_n7248;
  assign new_n7251 = new_n7250 ^ new_n7245;
  assign new_n7252 = new_n7251 ^ new_n7237;
  assign new_n7253 = new_n7252 ^ new_n7113;
  assign new_n7254 = new_n5936 ^ new_n3631;
  assign new_n7255 = new_n3481 ^ new_n432;
  assign new_n7256 = new_n7255 ^ new_n3615;
  assign new_n7257 = new_n7256 ^ new_n7254;
  assign new_n7258 = new_n5040 ^ new_n3666;
  assign new_n7259 = new_n7258 ^ new_n5963;
  assign new_n7260 = new_n3539 ^ new_n392;
  assign new_n7261 = new_n7260 ^ new_n3403;
  assign new_n7262 = new_n7261 ^ new_n7259;
  assign new_n7263 = new_n3565 ^ new_n3495;
  assign new_n7264 = new_n7263 ^ new_n3577;
  assign new_n7265 = new_n5040 ^ new_n402;
  assign new_n7266 = new_n7265 ^ new_n5939;
  assign new_n7267 = new_n7266 ^ new_n7264;
  assign new_n7268 = new_n7267 ^ new_n7262;
  assign new_n7269 = new_n5948 ^ new_n3153;
  assign new_n7270 = new_n3577 ^ new_n424;
  assign new_n7271 = new_n7270 ^ new_n3539;
  assign new_n7272 = new_n7271 ^ new_n7269;
  assign new_n7273 = new_n7272 ^ new_n7268;
  assign new_n7274 = new_n7273 ^ new_n7257;
  assign new_n7275 = new_n5942 ^ new_n3602;
  assign new_n7276 = new_n3376 ^ new_n364;
  assign new_n7277 = new_n7276 ^ new_n3481;
  assign new_n7278 = new_n7277 ^ new_n7275;
  assign new_n7279 = new_n5968 ^ new_n3615;
  assign new_n7280 = new_n5045 ^ new_n443;
  assign new_n7281 = new_n7280 ^ new_n7279;
  assign new_n7282 = new_n7281 ^ new_n7278;
  assign new_n7283 = new_n5974 ^ new_n373;
  assign new_n7284 = new_n7283 ^ new_n5040;
  assign new_n7285 = new_n3638 ^ new_n3582;
  assign new_n7286 = new_n7285 ^ new_n3565;
  assign new_n7287 = new_n7286 ^ new_n7284;
  assign new_n7288 = new_n7287 ^ new_n7278;
  assign new_n7289 = new_n7288 ^ new_n7268;
  assign new_n7290 = new_n3403 ^ new_n412;
  assign new_n7291 = new_n5951 ^ new_n5040;
  assign new_n7292 = new_n7291 ^ new_n7290;
  assign new_n7293 = new_n7292 ^ new_n7289;
  assign new_n7294 = new_n7281 ^ new_n7257;
  assign new_n7295 = new_n7294 ^ new_n7292;
  assign new_n7296 = new_n7295 ^ new_n7262;
  assign new_n7297 = new_n7278 ^ new_n7272;
  assign new_n7298 = new_n7297 ^ new_n7296;
  assign new_n7299 = new_n7293 & new_n7298;
  assign new_n7300 = new_n7295 ^ new_n7287;
  assign new_n7301 = new_n7292 & new_n7300;
  assign new_n7302 = new_n7301 ^ new_n7299;
  assign new_n7303 = new_n7287 ^ new_n7272;
  assign new_n7304 = new_n7287 ^ new_n7281;
  assign new_n7305 = new_n7304 ^ new_n7297;
  assign new_n7306 = new_n7303 & new_n7305;
  assign new_n7307 = new_n7294 ^ new_n7289;
  assign new_n7308 = new_n7297 & new_n7307;
  assign new_n7309 = new_n7308 ^ new_n7306;
  assign new_n7310 = new_n7309 ^ new_n7302;
  assign new_n7311 = new_n7310 ^ new_n7282;
  assign new_n7312 = ~new_n7262 & ~new_n7295;
  assign new_n7313 = new_n7312 ^ new_n7262;
  assign new_n7314 = new_n7278 ^ new_n7262;
  assign new_n7315 = new_n7281 ^ new_n7273;
  assign new_n7316 = new_n7314 & new_n7315;
  assign new_n7317 = new_n7316 ^ new_n7313;
  assign new_n7318 = new_n7317 ^ new_n7297;
  assign new_n7319 = new_n7274 & new_n7288;
  assign new_n7320 = new_n7319 ^ new_n7306;
  assign new_n7321 = new_n7281 ^ new_n7267;
  assign new_n7322 = new_n7321 ^ new_n7320;
  assign new_n7323 = new_n7322 ^ new_n7318;
  assign new_n7324 = new_n7314 ^ new_n7303;
  assign new_n7325 = new_n7289 & new_n7324;
  assign new_n7326 = new_n7325 ^ new_n7257;
  assign new_n7327 = new_n7326 ^ new_n7289;
  assign new_n7328 = new_n7319 ^ new_n7299;
  assign new_n7329 = new_n7306 ^ new_n7272;
  assign new_n7330 = new_n7329 ^ new_n7328;
  assign new_n7331 = new_n7330 ^ new_n7327;
  assign new_n7332 = ~new_n7323 & new_n7331;
  assign new_n7333 = new_n7319 ^ new_n7308;
  assign new_n7334 = new_n7333 ^ new_n7315;
  assign new_n7335 = new_n7292 ^ new_n7274;
  assign new_n7336 = new_n7295 ^ new_n7278;
  assign new_n7337 = new_n7335 & new_n7336;
  assign new_n7338 = new_n7337 ^ new_n7316;
  assign new_n7339 = new_n7338 ^ new_n7278;
  assign new_n7340 = new_n7339 ^ new_n7334;
  assign new_n7341 = new_n7340 ^ new_n7332;
  assign new_n7342 = new_n7311 & new_n7341;
  assign new_n7343 = new_n7301 ^ new_n7287;
  assign new_n7344 = new_n7343 ^ new_n7326;
  assign new_n7345 = new_n7344 ^ new_n7332;
  assign new_n7346 = new_n7345 ^ new_n7334;
  assign new_n7347 = new_n7337 ^ new_n7312;
  assign new_n7348 = new_n7347 ^ new_n7309;
  assign new_n7349 = ~new_n7348 & new_n7346;
  assign new_n7350 = new_n7349 ^ new_n7342;
  assign new_n7351 = new_n7344 ^ new_n7339;
  assign new_n7352 = new_n7351 ^ new_n7350;
  assign new_n7353 = new_n7274 & new_n7352;
  assign new_n7354 = new_n7349 ^ new_n7332;
  assign new_n7355 = ~new_n7354 & new_n7340;
  assign new_n7356 = new_n7355 ^ new_n7340;
  assign new_n7357 = new_n7356 ^ new_n7323;
  assign new_n7358 = ~new_n7357 & new_n7324;
  assign new_n7359 = new_n7358 ^ new_n7353;
  assign new_n7360 = new_n7344 ^ new_n7342;
  assign new_n7361 = new_n7360 ^ new_n7334;
  assign new_n7362 = new_n7355 ^ new_n7332;
  assign new_n7363 = new_n7361 & new_n7362;
  assign new_n7364 = new_n7363 ^ new_n7311;
  assign new_n7365 = new_n7295 & new_n7364;
  assign new_n7366 = new_n7356 ^ new_n7349;
  assign new_n7367 = new_n7366 ^ new_n7348;
  assign new_n7368 = ~new_n7367 & new_n7298;
  assign new_n7369 = new_n7288 & new_n7352;
  assign new_n7370 = new_n7281 ^ new_n7262;
  assign new_n7371 = new_n7313 ^ new_n7299;
  assign new_n7372 = new_n7363 ^ new_n7356;
  assign new_n7373 = new_n7372 ^ new_n7371;
  assign new_n7374 = new_n7373 ^ new_n7370;
  assign new_n7375 = new_n7374 ^ new_n7287;
  assign new_n7376 = new_n7342 ^ new_n7316;
  assign new_n7377 = new_n7376 ^ new_n7326;
  assign new_n7378 = new_n7377 ^ new_n7375;
  assign new_n7379 = ~new_n7378 & new_n7303;
  assign new_n7380 = new_n7379 ^ new_n7369;
  assign new_n7381 = new_n7380 ^ new_n7368;
  assign new_n7382 = new_n7381 ^ new_n7365;
  assign new_n7383 = new_n7363 ^ new_n7342;
  assign new_n7384 = new_n7383 ^ new_n7331;
  assign new_n7385 = new_n7315 & new_n7384;
  assign new_n7386 = new_n7385 ^ new_n7382;
  assign new_n7387 = ~new_n7378 & new_n7305;
  assign new_n7388 = new_n7387 ^ new_n7386;
  assign new_n7389 = new_n7388 ^ new_n7359;
  assign new_n7390 = new_n7105 ^ new_n7081;
  assign new_n7391 = new_n7089 ^ new_n7077;
  assign new_n7392 = new_n7391 ^ new_n7050;
  assign new_n7393 = new_n7012 & new_n7392;
  assign new_n7394 = new_n7089 ^ new_n7072;
  assign new_n7395 = new_n7019 & new_n7394;
  assign new_n7396 = new_n7395 ^ new_n7111;
  assign new_n7397 = new_n7396 ^ new_n7393;
  assign new_n7398 = new_n7397 ^ new_n7097;
  assign new_n7399 = new_n7398 ^ new_n7390;
  assign new_n7400 = new_n7399 ^ new_n7389;
  assign new_n7401 = new_n7400 ^ new_n7253;
  assign new_n7402 = new_n7401 ^ new_n6982;
  assign new_n7403 = new_n7220 ^ new_n7210;
  assign new_n7404 = new_n7155 & new_n7403;
  assign new_n7405 = new_n7404 ^ new_n7242;
  assign new_n7406 = new_n7224 ^ new_n7212;
  assign new_n7407 = new_n7406 ^ new_n7201;
  assign new_n7408 = new_n7184 & new_n7407;
  assign new_n7409 = new_n7408 ^ new_n7405;
  assign new_n7410 = new_n7183 & new_n7407;
  assign new_n7411 = new_n7410 ^ new_n7409;
  assign new_n7412 = new_n7224 ^ new_n7181;
  assign new_n7413 = new_n7163 & new_n7412;
  assign new_n7414 = new_n7206 & new_n7215;
  assign new_n7415 = new_n7414 ^ new_n7413;
  assign new_n7416 = new_n7415 ^ new_n7248;
  assign new_n7417 = new_n7416 ^ new_n7411;
  assign new_n7418 = new_n7162 & new_n7412;
  assign new_n7419 = new_n7418 ^ new_n7250;
  assign new_n7420 = new_n7419 ^ new_n7410;
  assign new_n7421 = new_n7420 ^ new_n7232;
  assign new_n7422 = new_n7244 ^ new_n7236;
  assign new_n7423 = new_n7422 ^ new_n7421;
  assign new_n7424 = new_n7423 ^ new_n7399;
  assign new_n7425 = new_n7424 ^ new_n7417;
  assign new_n7426 = new_n6941 ^ new_n6869;
  assign new_n7427 = new_n6906 ^ new_n6893;
  assign new_n7428 = new_n7427 ^ new_n6966;
  assign new_n7429 = new_n7428 ^ new_n7426;
  assign new_n7430 = ~new_n7429 & new_n6895;
  assign new_n7431 = new_n6907 & new_n6976;
  assign new_n7432 = new_n7431 ^ new_n7430;
  assign new_n7433 = new_n6979 ^ new_n6957;
  assign new_n7434 = ~new_n6888 & new_n6956;
  assign new_n7435 = ~new_n6904 & new_n6953;
  assign new_n7436 = new_n7435 ^ new_n7434;
  assign new_n7437 = new_n7436 ^ new_n6972;
  assign new_n7438 = new_n7437 ^ new_n7433;
  assign new_n7439 = new_n7438 ^ new_n7432;
  assign new_n7440 = new_n7349 ^ new_n7278;
  assign new_n7441 = new_n7337 ^ new_n7301;
  assign new_n7442 = new_n7441 ^ new_n7374;
  assign new_n7443 = new_n7442 ^ new_n7440;
  assign new_n7444 = ~new_n7443 & new_n7307;
  assign new_n7445 = new_n7314 & new_n7384;
  assign new_n7446 = new_n7445 ^ new_n7444;
  assign new_n7447 = new_n7387 ^ new_n7365;
  assign new_n7448 = new_n7296 & new_n7364;
  assign new_n7449 = new_n7335 & new_n7361;
  assign new_n7450 = new_n7449 ^ new_n7448;
  assign new_n7451 = new_n7450 ^ new_n7380;
  assign new_n7452 = new_n7451 ^ new_n7447;
  assign new_n7453 = new_n7452 ^ new_n7446;
  assign new_n7454 = new_n7453 ^ new_n7439;
  assign new_n7455 = new_n7454 ^ new_n7425;
  assign new_n7456 = new_n1008 ^ new_n1002;
  assign new_n7457 = new_n994 ^ new_n988;
  assign new_n7458 = ~new_n987 & new_n930;
  assign new_n7459 = ~new_n944 & ~new_n975;
  assign new_n7460 = new_n7459 ^ new_n7458;
  assign new_n7461 = new_n7460 ^ new_n985;
  assign new_n7462 = new_n7461 ^ new_n7457;
  assign new_n7463 = new_n7462 ^ new_n7456;
  assign new_n7464 = new_n7463 ^ n87;
  assign new_n7465 = new_n7464 ^ n23;
  assign new_n7466 = new_n7068 ^ new_n7006;
  assign new_n7467 = new_n7064 ^ new_n7053;
  assign new_n7468 = new_n7467 ^ new_n7092;
  assign new_n7469 = new_n7468 ^ new_n7466;
  assign new_n7470 = ~new_n7469 & new_n7057;
  assign new_n7471 = new_n7007 & new_n7392;
  assign new_n7472 = new_n7471 ^ new_n7470;
  assign new_n7473 = new_n7395 ^ new_n7097;
  assign new_n7474 = new_n7045 & new_n7394;
  assign new_n7475 = new_n7062 & new_n7085;
  assign new_n7476 = new_n7475 ^ new_n7474;
  assign new_n7477 = new_n7476 ^ new_n7110;
  assign new_n7478 = new_n7477 ^ new_n7473;
  assign new_n7479 = new_n7478 ^ new_n7472;
  assign new_n7480 = new_n7479 ^ new_n7465;
  assign new_n7481 = new_n7075 ^ new_n7068;
  assign new_n7482 = new_n7017 & new_n7481;
  assign new_n7483 = new_n7482 ^ new_n7103;
  assign new_n7484 = new_n7483 ^ new_n7471;
  assign new_n7485 = new_n7484 ^ new_n7393;
  assign new_n7486 = new_n7485 ^ new_n7477;
  assign new_n7487 = new_n7486 ^ new_n7480;
  assign new_n7488 = new_n7487 ^ new_n7455;
  assign new_n7489 = new_n7488 ^ new_n7402;
  assign new_n7490 = new_n6941 ^ new_n6915;
  assign new_n7491 = ~new_n6892 & new_n7490;
  assign new_n7492 = new_n7491 ^ new_n6980;
  assign new_n7493 = ~new_n6905 & new_n6953;
  assign new_n7494 = new_n7493 ^ new_n7430;
  assign new_n7495 = ~new_n6949 & new_n6881;
  assign new_n7496 = ~new_n6884 & new_n7490;
  assign new_n7497 = new_n7496 ^ new_n7495;
  assign new_n7498 = new_n7497 ^ new_n7431;
  assign new_n7499 = new_n7498 ^ new_n7494;
  assign new_n7500 = new_n7499 ^ new_n7492;
  assign new_n7501 = new_n7349 ^ new_n7340;
  assign new_n7502 = new_n7300 & new_n7501;
  assign new_n7503 = new_n7502 ^ new_n7388;
  assign new_n7504 = new_n7336 & new_n7361;
  assign new_n7505 = new_n7504 ^ new_n7444;
  assign new_n7506 = ~new_n7357 & new_n7289;
  assign new_n7507 = new_n7292 & new_n7501;
  assign new_n7508 = new_n7507 ^ new_n7506;
  assign new_n7509 = new_n7508 ^ new_n7445;
  assign new_n7510 = new_n7509 ^ new_n7505;
  assign new_n7511 = new_n7510 ^ new_n7503;
  assign new_n7512 = new_n7511 ^ new_n7500;
  assign new_n7513 = new_n7220 ^ new_n7136;
  assign new_n7514 = new_n7207 ^ new_n7173;
  assign new_n7515 = new_n7514 ^ new_n7227;
  assign new_n7516 = new_n7515 ^ new_n7513;
  assign new_n7517 = ~new_n7516 & new_n7177;
  assign new_n7518 = new_n7517 ^ new_n7408;
  assign new_n7519 = new_n7418 ^ new_n7232;
  assign new_n7520 = new_n7519 ^ new_n7416;
  assign new_n7521 = new_n7520 ^ new_n7518;
  assign new_n7522 = new_n7521 ^ new_n7512;
  assign new_n7523 = new_n1012 ^ n22;
  assign new_n7524 = new_n7063 & new_n7085;
  assign new_n7525 = new_n7524 ^ new_n7470;
  assign new_n7526 = new_n7525 ^ new_n7484;
  assign new_n7527 = new_n7052 & new_n7481;
  assign new_n7528 = new_n7527 ^ new_n7398;
  assign new_n7529 = new_n7528 ^ new_n7526;
  assign new_n7530 = new_n7529 ^ new_n7523;
  assign new_n7531 = new_n7530 ^ new_n7479;
  assign new_n7532 = new_n7531 ^ new_n7522;
  assign new_n7533 = new_n7532 ^ new_n7402;
  assign new_n7534 = new_n6839 ^ new_n994;
  assign new_n7535 = new_n929 & new_n961;
  assign new_n7536 = new_n7535 ^ new_n1006;
  assign new_n7537 = new_n7536 ^ new_n6840;
  assign new_n7538 = new_n7537 ^ new_n986;
  assign new_n7539 = new_n7538 ^ new_n7534;
  assign new_n7540 = new_n7539 ^ n82;
  assign new_n7541 = new_n7540 ^ n18;
  assign new_n7542 = new_n6979 ^ new_n6945;
  assign new_n7543 = ~new_n6885 & ~new_n6959;
  assign new_n7544 = new_n7543 ^ new_n7495;
  assign new_n7545 = new_n7544 ^ new_n6950;
  assign new_n7546 = new_n7545 ^ new_n6973;
  assign new_n7547 = new_n7546 ^ new_n7542;
  assign new_n7548 = new_n7547 ^ new_n7541;
  assign new_n7549 = new_n7246 ^ new_n7236;
  assign new_n7550 = ~new_n7516 & new_n7137;
  assign new_n7551 = new_n7205 & new_n7215;
  assign new_n7552 = new_n7551 ^ new_n7517;
  assign new_n7553 = new_n7552 ^ new_n7409;
  assign new_n7554 = new_n7553 ^ new_n7550;
  assign new_n7555 = new_n7554 ^ new_n7549;
  assign new_n7556 = new_n7108 ^ new_n7081;
  assign new_n7557 = ~new_n7469 & new_n7023;
  assign new_n7558 = new_n7557 ^ new_n7526;
  assign new_n7559 = new_n7558 ^ new_n7556;
  assign new_n7560 = new_n7559 ^ new_n7555;
  assign new_n7561 = new_n7387 ^ new_n7353;
  assign new_n7562 = ~new_n7367 & new_n7293;
  assign new_n7563 = new_n7562 ^ new_n7506;
  assign new_n7564 = new_n7563 ^ new_n7358;
  assign new_n7565 = new_n7564 ^ new_n7381;
  assign new_n7566 = new_n7565 ^ new_n7561;
  assign new_n7567 = new_n7566 ^ new_n7113;
  assign new_n7568 = new_n7567 ^ new_n7560;
  assign new_n7569 = new_n7568 ^ new_n7548;
  assign new_n7570 = new_n6839 ^ new_n971;
  assign new_n7571 = ~new_n1001 & new_n905;
  assign new_n7572 = new_n7571 ^ new_n1010;
  assign new_n7573 = new_n7572 ^ new_n7570;
  assign new_n7574 = new_n7573 ^ n83;
  assign new_n7575 = new_n7574 ^ n19;
  assign new_n7576 = new_n6961 ^ new_n6945;
  assign new_n7577 = ~new_n7429 & new_n6889;
  assign new_n7578 = new_n7577 ^ new_n7499;
  assign new_n7579 = new_n7578 ^ new_n7576;
  assign new_n7580 = new_n7579 ^ new_n7575;
  assign new_n7581 = new_n7420 ^ new_n7245;
  assign new_n7582 = new_n7397 ^ new_n7106;
  assign new_n7583 = new_n7582 ^ new_n7581;
  assign new_n7584 = new_n7369 ^ new_n7353;
  assign new_n7585 = ~new_n7443 & new_n7297;
  assign new_n7586 = new_n7585 ^ new_n7510;
  assign new_n7587 = new_n7586 ^ new_n7584;
  assign new_n7588 = new_n7587 ^ new_n7559;
  assign new_n7589 = new_n7588 ^ new_n7583;
  assign new_n7590 = new_n7589 ^ new_n7580;
  assign new_n7591 = new_n7590 ^ new_n7569;
  assign new_n7592 = new_n7537 ^ new_n993;
  assign new_n7593 = new_n7592 ^ n84;
  assign new_n7594 = new_n7593 ^ n20;
  assign new_n7595 = new_n7594 ^ new_n7424;
  assign new_n7596 = new_n7564 ^ new_n7386;
  assign new_n7597 = new_n7596 ^ new_n7582;
  assign new_n7598 = new_n7597 ^ new_n7595;
  assign new_n7599 = new_n7414 ^ new_n7244;
  assign new_n7600 = new_n7404 ^ new_n7240;
  assign new_n7601 = new_n7600 ^ new_n7419;
  assign new_n7602 = new_n7601 ^ new_n7599;
  assign new_n7603 = new_n7475 ^ new_n7105;
  assign new_n7604 = new_n7482 ^ new_n7101;
  assign new_n7605 = new_n7604 ^ new_n7396;
  assign new_n7606 = new_n7605 ^ new_n7603;
  assign new_n7607 = new_n7606 ^ new_n7602;
  assign new_n7608 = new_n7545 ^ new_n6978;
  assign new_n7609 = new_n7608 ^ new_n7607;
  assign new_n7610 = new_n7609 ^ new_n7598;
  assign new_n7611 = new_n7610 ^ new_n7402;
  assign new_n7612 = new_n7606 ^ new_n7529;
  assign new_n7613 = new_n7162 ^ new_n7125;
  assign new_n7614 = new_n7403 & new_n7613;
  assign new_n7615 = new_n7614 ^ new_n7421;
  assign new_n7616 = new_n7615 ^ new_n7553;
  assign new_n7617 = new_n7616 ^ new_n7612;
  assign new_n7618 = new_n7459 ^ new_n6840;
  assign new_n7619 = new_n7535 ^ new_n1004;
  assign new_n7620 = new_n7619 ^ new_n989;
  assign new_n7621 = new_n7620 ^ new_n7618;
  assign new_n7622 = new_n7621 ^ n85;
  assign new_n7623 = new_n7622 ^ n21;
  assign new_n7624 = new_n7623 ^ new_n7424;
  assign new_n7625 = new_n7435 ^ new_n6950;
  assign new_n7626 = new_n7543 ^ new_n7496;
  assign new_n7627 = new_n7626 ^ new_n6974;
  assign new_n7628 = new_n7627 ^ new_n7625;
  assign new_n7629 = new_n7449 ^ new_n7358;
  assign new_n7630 = new_n7562 ^ new_n7507;
  assign new_n7631 = new_n7630 ^ new_n7382;
  assign new_n7632 = new_n7631 ^ new_n7629;
  assign new_n7633 = new_n7632 ^ new_n7628;
  assign new_n7634 = new_n7633 ^ new_n7624;
  assign new_n7635 = new_n7634 ^ new_n7617;
  assign new_n7636 = new_n7635 ^ new_n7488;
  assign new_n7637 = new_n7636 ^ new_n7611;
  assign new_n7638 = new_n7637 ^ new_n7591;
  assign new_n7639 = new_n7533 & new_n7638;
  assign new_n7640 = new_n7636 ^ new_n7532;
  assign new_n7641 = new_n7640 ^ new_n7569;
  assign new_n7642 = new_n7611 & new_n7641;
  assign new_n7643 = new_n7642 ^ new_n7639;
  assign new_n7644 = new_n7640 ^ new_n7590;
  assign new_n7645 = new_n7644 ^ new_n7643;
  assign new_n7646 = new_n1009 ^ new_n992;
  assign new_n7647 = new_n7646 ^ new_n7461;
  assign new_n7648 = new_n7647 ^ n88;
  assign new_n7649 = new_n7648 ^ n24;
  assign new_n7650 = new_n7649 ^ new_n7486;
  assign new_n7651 = new_n7498 ^ new_n6977;
  assign new_n7652 = new_n7651 ^ new_n7437;
  assign new_n7653 = new_n7509 ^ new_n7385;
  assign new_n7654 = new_n7653 ^ new_n7451;
  assign new_n7655 = new_n7654 ^ new_n7652;
  assign new_n7656 = new_n7655 ^ new_n7424;
  assign new_n7657 = new_n7656 ^ new_n7650;
  assign new_n7658 = new_n7657 ^ new_n7591;
  assign new_n7659 = new_n7658 ^ new_n7402;
  assign new_n7660 = new_n7657 ^ new_n7641;
  assign new_n7661 = new_n7659 & new_n7660;
  assign new_n7662 = new_n7489 & new_n7644;
  assign new_n7663 = new_n7662 ^ new_n7661;
  assign new_n7664 = new_n7663 ^ new_n7402;
  assign new_n7665 = new_n7664 ^ new_n7645;
  assign new_n7666 = new_n7658 ^ new_n7610;
  assign new_n7667 = new_n7657 & new_n7666;
  assign new_n7668 = new_n7667 ^ new_n7610;
  assign new_n7669 = new_n7610 ^ new_n7532;
  assign new_n7670 = new_n7669 ^ new_n7489;
  assign new_n7671 = new_n7637 & new_n7670;
  assign new_n7672 = new_n7671 ^ new_n7569;
  assign new_n7673 = new_n7672 ^ new_n7668;
  assign new_n7674 = ~new_n7488 & ~new_n7658;
  assign new_n7675 = new_n7674 ^ new_n7488;
  assign new_n7676 = new_n7675 ^ new_n7662;
  assign new_n7677 = new_n7676 ^ new_n7533;
  assign new_n7678 = new_n7610 ^ new_n7590;
  assign new_n7679 = new_n7678 ^ new_n7533;
  assign new_n7680 = new_n7669 & new_n7679;
  assign new_n7681 = new_n7680 ^ new_n7642;
  assign new_n7682 = new_n7635 ^ new_n7590;
  assign new_n7683 = new_n7682 ^ new_n7681;
  assign new_n7684 = new_n7683 ^ new_n7677;
  assign new_n7685 = new_n7672 ^ new_n7637;
  assign new_n7686 = new_n7657 ^ new_n7637;
  assign new_n7687 = new_n7658 ^ new_n7488;
  assign new_n7688 = new_n7687 ^ new_n7533;
  assign new_n7689 = new_n7686 & new_n7688;
  assign new_n7690 = new_n7689 ^ new_n7681;
  assign new_n7691 = new_n7690 ^ new_n7532;
  assign new_n7692 = new_n7691 ^ new_n7685;
  assign new_n7693 = ~new_n7684 & new_n7692;
  assign new_n7694 = new_n7693 ^ new_n7673;
  assign new_n7695 = new_n7694 ^ new_n7645;
  assign new_n7696 = new_n7680 ^ new_n7639;
  assign new_n7697 = new_n7674 ^ new_n7661;
  assign new_n7698 = new_n7697 ^ new_n7696;
  assign new_n7699 = ~new_n7698 & new_n7695;
  assign new_n7700 = new_n7699 ^ new_n7693;
  assign new_n7701 = ~new_n7665 & ~new_n7700;
  assign new_n7702 = new_n7701 ^ new_n7699;
  assign new_n7703 = new_n7693 ^ new_n7665;
  assign new_n7704 = new_n7590 ^ new_n7402;
  assign new_n7705 = new_n7689 ^ new_n7667;
  assign new_n7706 = new_n7705 ^ new_n7696;
  assign new_n7707 = new_n7706 ^ new_n7704;
  assign new_n7708 = new_n7703 & new_n7707;
  assign new_n7709 = new_n7708 ^ new_n7673;
  assign new_n7710 = new_n7709 ^ new_n7645;
  assign new_n7711 = ~new_n7702 & new_n7710;
  assign new_n7712 = new_n7711 ^ new_n7708;
  assign new_n7713 = new_n7712 ^ new_n7692;
  assign new_n7714 = new_n7489 & new_n7713;
  assign new_n7715 = new_n7699 ^ new_n7402;
  assign new_n7716 = new_n7667 ^ new_n7661;
  assign new_n7717 = new_n7590 ^ new_n7488;
  assign new_n7718 = new_n7689 ^ new_n7675;
  assign new_n7719 = new_n7703 ^ new_n7702;
  assign new_n7720 = new_n7719 ^ new_n7711;
  assign new_n7721 = new_n7720 ^ new_n7718;
  assign new_n7722 = new_n7721 ^ new_n7717;
  assign new_n7723 = new_n7722 ^ new_n7716;
  assign new_n7724 = new_n7723 ^ new_n7715;
  assign new_n7725 = new_n7638 & new_n7724;
  assign new_n7726 = new_n7725 ^ new_n7714;
  assign new_n7727 = new_n7722 ^ new_n7610;
  assign new_n7728 = new_n7708 ^ new_n7662;
  assign new_n7729 = new_n7728 ^ new_n7672;
  assign new_n7730 = new_n7729 ^ new_n7727;
  assign new_n7731 = new_n7679 & new_n7730;
  assign new_n7732 = new_n7711 ^ new_n7707;
  assign new_n7733 = new_n7658 & new_n7732;
  assign new_n7734 = new_n7733 ^ new_n7731;
  assign new_n7735 = new_n7687 & new_n7732;
  assign new_n7736 = new_n7660 & new_n7710;
  assign new_n7737 = new_n7736 ^ new_n7735;
  assign new_n7738 = new_n7708 ^ new_n7699;
  assign new_n7739 = new_n7673 ^ new_n7664;
  assign new_n7740 = new_n7739 ^ new_n7738;
  assign new_n7741 = new_n7611 & new_n7740;
  assign new_n7742 = new_n7669 & new_n7730;
  assign new_n7743 = new_n7742 ^ new_n7741;
  assign new_n7744 = new_n7743 ^ new_n7737;
  assign new_n7745 = new_n7744 ^ new_n7734;
  assign new_n7746 = new_n7745 ^ new_n7726;
  assign new_n7747 = new_n5794 ^ new_n5788;
  assign new_n7748 = ~new_n5756 & new_n5716;
  assign new_n7749 = ~new_n5731 & ~new_n5751;
  assign new_n7750 = new_n7749 ^ new_n7748;
  assign new_n7751 = new_n7750 ^ new_n5773;
  assign new_n7752 = new_n5780 ^ new_n5757;
  assign new_n7753 = new_n7752 ^ new_n7751;
  assign new_n7754 = new_n7753 ^ new_n7747;
  assign new_n7755 = new_n7754 ^ new_n7746;
  assign new_n7756 = new_n7755 ^ new_n6838;
  assign new_n7757 = new_n7756 ^ new_n4900;
  assign new_n7758 = new_n6834 ^ new_n6828;
  assign new_n7759 = new_n6805 ^ new_n6803;
  assign new_n7760 = new_n6753 & new_n6804;
  assign new_n7761 = new_n6769 & new_n6793;
  assign new_n7762 = new_n7761 ^ new_n7760;
  assign new_n7763 = new_n7762 ^ new_n6811;
  assign new_n7764 = new_n7763 ^ new_n7759;
  assign new_n7765 = new_n7764 ^ new_n7758;
  assign new_n7766 = new_n7765 ^ new_n7754;
  assign new_n7767 = new_n5795 ^ new_n5755;
  assign new_n7768 = new_n7767 ^ new_n7751;
  assign new_n7769 = new_n7719 ^ new_n7684;
  assign new_n7770 = new_n7637 & new_n7769;
  assign new_n7771 = new_n7699 ^ new_n7665;
  assign new_n7772 = new_n7657 & new_n7771;
  assign new_n7773 = new_n7772 ^ new_n7770;
  assign new_n7774 = new_n7773 ^ new_n7714;
  assign new_n7775 = new_n7644 & new_n7713;
  assign new_n7776 = new_n7775 ^ new_n7774;
  assign new_n7777 = new_n7776 ^ new_n7744;
  assign new_n7778 = new_n7777 ^ new_n7768;
  assign new_n7779 = new_n7778 ^ new_n7766;
  assign new_n7780 = new_n710 ^ new_n704;
  assign new_n7781 = new_n681 ^ new_n679;
  assign new_n7782 = ~new_n680 & new_n632;
  assign new_n7783 = ~new_n647 & ~new_n669;
  assign new_n7784 = new_n7783 ^ new_n7782;
  assign new_n7785 = new_n7784 ^ new_n687;
  assign new_n7786 = new_n7785 ^ new_n7781;
  assign new_n7787 = new_n7786 ^ new_n7780;
  assign new_n7788 = new_n7787 ^ n55;
  assign new_n7789 = new_n7788 ^ new_n7464;
  assign new_n7790 = new_n4896 ^ new_n4890;
  assign new_n7791 = new_n4867 ^ new_n4865;
  assign new_n7792 = ~new_n4866 & new_n4815;
  assign new_n7793 = ~new_n4832 & new_n4852;
  assign new_n7794 = new_n7793 ^ new_n7792;
  assign new_n7795 = new_n7794 ^ new_n4873;
  assign new_n7796 = new_n7795 ^ new_n7791;
  assign new_n7797 = new_n7796 ^ new_n7790;
  assign new_n7798 = new_n7797 ^ new_n7789;
  assign new_n7799 = new_n7641 & new_n7740;
  assign new_n7800 = new_n7670 & new_n7769;
  assign new_n7801 = new_n7800 ^ new_n7799;
  assign new_n7802 = new_n7719 ^ new_n7699;
  assign new_n7803 = new_n7802 ^ new_n7698;
  assign new_n7804 = new_n7688 & new_n7803;
  assign new_n7805 = new_n7804 ^ new_n7743;
  assign new_n7806 = new_n7805 ^ new_n7733;
  assign new_n7807 = new_n7806 ^ new_n7775;
  assign new_n7808 = new_n7807 ^ new_n7731;
  assign new_n7809 = new_n7808 ^ new_n7801;
  assign new_n7810 = ~new_n5760 & new_n5704;
  assign new_n7811 = ~new_n5692 & new_n5790;
  assign new_n7812 = new_n7811 ^ new_n7810;
  assign new_n7813 = new_n7812 ^ new_n5781;
  assign new_n7814 = new_n7813 ^ new_n7809;
  assign new_n7815 = new_n7814 ^ new_n7798;
  assign new_n7816 = new_n7815 ^ new_n7779;
  assign new_n7817 = ~new_n608 & new_n707;
  assign new_n7818 = new_n7817 ^ new_n7783;
  assign new_n7819 = new_n631 & new_n689;
  assign new_n7820 = new_n7819 ^ new_n706;
  assign new_n7821 = new_n7820 ^ new_n692;
  assign new_n7822 = new_n7821 ^ new_n7818;
  assign new_n7823 = new_n7822 ^ n53;
  assign new_n7824 = new_n7823 ^ new_n7622;
  assign new_n7825 = ~new_n4892 & new_n4810;
  assign new_n7826 = new_n7825 ^ new_n7793;
  assign new_n7827 = new_n4814 & new_n4875;
  assign new_n7828 = new_n7827 ^ new_n4894;
  assign new_n7829 = new_n7828 ^ new_n4878;
  assign new_n7830 = new_n7829 ^ new_n7826;
  assign new_n7831 = new_n7830 ^ new_n7824;
  assign new_n7832 = new_n7831 ^ new_n7814;
  assign new_n7833 = new_n6748 & new_n6831;
  assign new_n7834 = new_n7833 ^ new_n7761;
  assign new_n7835 = new_n6752 & new_n6813;
  assign new_n7836 = new_n7835 ^ new_n6830;
  assign new_n7837 = new_n7836 ^ new_n6816;
  assign new_n7838 = new_n7837 ^ new_n7834;
  assign new_n7839 = new_n7811 ^ new_n7749;
  assign new_n7840 = new_n5715 & new_n5775;
  assign new_n7841 = new_n7840 ^ new_n5792;
  assign new_n7842 = new_n7841 ^ new_n5778;
  assign new_n7843 = new_n7842 ^ new_n7839;
  assign new_n7844 = new_n7843 ^ new_n7838;
  assign new_n7845 = new_n7666 & new_n7771;
  assign new_n7846 = new_n7845 ^ new_n7808;
  assign new_n7847 = new_n7659 & new_n7710;
  assign new_n7848 = new_n7847 ^ new_n7725;
  assign new_n7849 = new_n7848 ^ new_n7774;
  assign new_n7850 = new_n7849 ^ new_n7846;
  assign new_n7851 = new_n7850 ^ new_n5797;
  assign new_n7852 = new_n7851 ^ new_n7844;
  assign new_n7853 = new_n7852 ^ new_n7832;
  assign new_n7854 = new_n7853 ^ new_n7816;
  assign new_n7855 = new_n7854 ^ new_n7757;
  assign new_n7856 = ~new_n685 & new_n624;
  assign new_n7857 = new_n7856 ^ new_n679;
  assign new_n7858 = new_n7819 ^ new_n708;
  assign new_n7859 = new_n7858 ^ new_n7817;
  assign new_n7860 = new_n7859 ^ new_n691;
  assign new_n7861 = new_n7860 ^ new_n7857;
  assign new_n7862 = new_n7861 ^ n50;
  assign new_n7863 = new_n7862 ^ new_n7540;
  assign new_n7864 = ~new_n4797 & ~new_n4871;
  assign new_n7865 = new_n7864 ^ new_n4865;
  assign new_n7866 = new_n7827 ^ new_n4893;
  assign new_n7867 = new_n7866 ^ new_n7825;
  assign new_n7868 = new_n7867 ^ new_n4877;
  assign new_n7869 = new_n7868 ^ new_n7865;
  assign new_n7870 = new_n7869 ^ new_n7863;
  assign new_n7871 = new_n7810 ^ new_n5780;
  assign new_n7872 = new_n7840 ^ new_n5791;
  assign new_n7873 = new_n7872 ^ new_n7811;
  assign new_n7874 = new_n7873 ^ new_n5777;
  assign new_n7875 = new_n7874 ^ new_n7871;
  assign new_n7876 = new_n6739 & new_n6808;
  assign new_n7877 = new_n7876 ^ new_n6803;
  assign new_n7878 = new_n7835 ^ new_n6832;
  assign new_n7879 = new_n7878 ^ new_n7833;
  assign new_n7880 = new_n7879 ^ new_n6815;
  assign new_n7881 = new_n7880 ^ new_n7877;
  assign new_n7882 = new_n7881 ^ new_n7875;
  assign new_n7883 = new_n7810 ^ new_n5761;
  assign new_n7884 = ~new_n5787 & new_n5691;
  assign new_n7885 = new_n7884 ^ new_n5796;
  assign new_n7886 = new_n7885 ^ new_n7883;
  assign new_n7887 = new_n7799 ^ new_n7741;
  assign new_n7888 = new_n7533 & new_n7724;
  assign new_n7889 = new_n7888 ^ new_n7849;
  assign new_n7890 = new_n7889 ^ new_n7887;
  assign new_n7891 = new_n7890 ^ new_n7886;
  assign new_n7892 = new_n7891 ^ new_n7882;
  assign new_n7893 = new_n7892 ^ new_n7870;
  assign new_n7894 = new_n7893 ^ new_n7855;
  assign new_n7895 = new_n711 ^ new_n695;
  assign new_n7896 = new_n7895 ^ new_n7785;
  assign new_n7897 = new_n7896 ^ n56;
  assign new_n7898 = new_n7897 ^ new_n7648;
  assign new_n7899 = new_n4897 ^ new_n4881;
  assign new_n7900 = new_n7899 ^ new_n7795;
  assign new_n7901 = new_n7900 ^ new_n7898;
  assign new_n7902 = new_n6835 ^ new_n6819;
  assign new_n7903 = new_n7902 ^ new_n7763;
  assign new_n7904 = new_n7903 ^ new_n7768;
  assign new_n7905 = new_n7904 ^ new_n7814;
  assign new_n7906 = new_n7905 ^ new_n7901;
  assign new_n7907 = new_n7856 ^ new_n686;
  assign new_n7908 = ~new_n703 & new_n607;
  assign new_n7909 = new_n7908 ^ new_n712;
  assign new_n7910 = new_n7909 ^ new_n7907;
  assign new_n7911 = new_n7910 ^ n51;
  assign new_n7912 = new_n7911 ^ new_n7574;
  assign new_n7913 = new_n7864 ^ new_n4872;
  assign new_n7914 = ~new_n4889 & new_n4795;
  assign new_n7915 = new_n7914 ^ new_n4898;
  assign new_n7916 = new_n7915 ^ new_n7913;
  assign new_n7917 = new_n7916 ^ new_n7912;
  assign new_n7918 = new_n7876 ^ new_n6809;
  assign new_n7919 = new_n6733 & new_n6827;
  assign new_n7920 = new_n7919 ^ new_n6836;
  assign new_n7921 = new_n7920 ^ new_n7918;
  assign new_n7922 = new_n7921 ^ new_n7886;
  assign new_n7923 = new_n7686 & new_n7803;
  assign new_n7924 = new_n7923 ^ new_n7770;
  assign new_n7925 = new_n7924 ^ new_n7800;
  assign new_n7926 = new_n7925 ^ new_n7807;
  assign new_n7927 = new_n7873 ^ new_n5779;
  assign new_n7928 = new_n7927 ^ new_n7926;
  assign new_n7929 = new_n7928 ^ new_n7922;
  assign new_n7930 = new_n7929 ^ new_n7917;
  assign new_n7931 = new_n7930 ^ new_n7893;
  assign new_n7932 = new_n7931 ^ new_n7906;
  assign new_n7933 = new_n7816 & new_n7932;
  assign new_n7934 = new_n7933 ^ new_n7816;
  assign new_n7935 = new_n7930 ^ new_n7855;
  assign new_n7936 = new_n7856 ^ new_n7817;
  assign new_n7937 = new_n7936 ^ new_n697;
  assign new_n7938 = new_n7937 ^ n49;
  assign new_n7939 = new_n7938 ^ new_n6843;
  assign new_n7940 = new_n7864 ^ new_n7825;
  assign new_n7941 = new_n7940 ^ new_n4883;
  assign new_n7942 = new_n7941 ^ new_n7939;
  assign new_n7943 = new_n7876 ^ new_n7833;
  assign new_n7944 = new_n7943 ^ new_n6821;
  assign new_n7945 = new_n7944 ^ new_n7813;
  assign new_n7946 = new_n7799 ^ new_n7731;
  assign new_n7947 = new_n7925 ^ new_n7805;
  assign new_n7948 = new_n7947 ^ new_n7946;
  assign new_n7949 = new_n7948 ^ new_n7875;
  assign new_n7950 = new_n7949 ^ new_n7945;
  assign new_n7951 = new_n7950 ^ new_n7942;
  assign new_n7952 = new_n7951 ^ new_n7816;
  assign new_n7953 = ~new_n7952 & new_n7935;
  assign new_n7954 = new_n7953 ^ new_n7934;
  assign new_n7955 = new_n7951 ^ new_n7757;
  assign new_n7956 = new_n7955 ^ new_n7954;
  assign new_n7957 = new_n7879 ^ new_n6820;
  assign new_n7958 = new_n7957 ^ new_n7927;
  assign new_n7959 = new_n7800 ^ new_n7736;
  assign new_n7960 = new_n7923 ^ new_n7772;
  assign new_n7961 = new_n7960 ^ new_n7806;
  assign new_n7962 = new_n7961 ^ new_n7959;
  assign new_n7963 = new_n7962 ^ new_n7843;
  assign new_n7964 = new_n7963 ^ new_n7958;
  assign new_n7965 = new_n7859 ^ new_n696;
  assign new_n7966 = new_n7965 ^ n52;
  assign new_n7967 = new_n7966 ^ new_n7593;
  assign new_n7968 = new_n7867 ^ new_n4882;
  assign new_n7969 = new_n7968 ^ new_n7967;
  assign new_n7970 = new_n7969 ^ new_n7814;
  assign new_n7971 = new_n7970 ^ new_n7964;
  assign new_n7972 = new_n7971 ^ new_n7951;
  assign new_n7973 = new_n7894 & new_n7972;
  assign new_n7974 = new_n7971 ^ new_n7930;
  assign new_n7975 = new_n7974 ^ new_n7955;
  assign new_n7976 = new_n7971 ^ new_n7757;
  assign new_n7977 = ~new_n7975 & new_n7976;
  assign new_n7978 = new_n7977 ^ new_n7973;
  assign new_n7979 = new_n7930 ^ new_n7853;
  assign new_n7980 = new_n7979 ^ new_n7978;
  assign new_n7981 = new_n7980 ^ new_n7956;
  assign new_n7982 = new_n7972 ^ new_n7854;
  assign new_n7983 = new_n7971 ^ new_n7816;
  assign new_n7984 = new_n7983 ^ new_n7955;
  assign new_n7985 = ~new_n7982 & ~new_n7984;
  assign new_n7986 = new_n7985 ^ new_n7893;
  assign new_n7987 = new_n7986 ^ new_n7982;
  assign new_n7988 = new_n7982 ^ new_n7906;
  assign new_n7989 = new_n7932 ^ new_n7816;
  assign new_n7990 = new_n7989 ^ new_n7955;
  assign new_n7991 = new_n7988 & new_n7990;
  assign new_n7992 = new_n7991 ^ new_n7973;
  assign new_n7993 = new_n7977 ^ new_n7757;
  assign new_n7994 = new_n7993 ^ new_n7992;
  assign new_n7995 = new_n7994 ^ new_n7987;
  assign new_n7996 = ~new_n7981 & new_n7995;
  assign new_n7997 = new_n7971 ^ new_n7932;
  assign new_n7998 = ~new_n7906 & ~new_n7997;
  assign new_n7999 = new_n7998 ^ new_n7971;
  assign new_n8000 = new_n7999 ^ new_n7986;
  assign new_n8001 = new_n8000 ^ new_n7996;
  assign new_n8002 = new_n7982 ^ new_n7931;
  assign new_n8003 = ~new_n8002 & new_n7955;
  assign new_n8004 = new_n8003 ^ new_n7973;
  assign new_n8005 = new_n8004 ^ new_n7935;
  assign new_n8006 = new_n8005 ^ new_n8001;
  assign new_n8007 = new_n7951 ^ new_n7932;
  assign new_n8008 = new_n7906 ^ new_n7894;
  assign new_n8009 = ~new_n8007 & ~new_n8008;
  assign new_n8010 = new_n8009 ^ new_n7933;
  assign new_n8011 = new_n8003 ^ new_n7977;
  assign new_n8012 = new_n8011 ^ new_n8010;
  assign new_n8013 = ~new_n8006 & ~new_n8012;
  assign new_n8014 = new_n7951 ^ new_n7930;
  assign new_n8015 = new_n7998 ^ new_n7991;
  assign new_n8016 = new_n8015 ^ new_n8011;
  assign new_n8017 = new_n8016 ^ new_n8014;
  assign new_n8018 = new_n8009 ^ new_n7953;
  assign new_n8019 = new_n8018 ^ new_n7951;
  assign new_n8020 = new_n8019 ^ new_n8005;
  assign new_n8021 = new_n8020 ^ new_n7996;
  assign new_n8022 = ~new_n8017 & new_n8021;
  assign new_n8023 = new_n8022 ^ new_n8013;
  assign new_n8024 = new_n8019 ^ new_n8000;
  assign new_n8025 = new_n8024 ^ new_n8023;
  assign new_n8026 = ~new_n8025 & new_n7894;
  assign new_n8027 = ~new_n8025 & new_n7972;
  assign new_n8028 = new_n8027 ^ new_n8026;
  assign new_n8029 = new_n8013 ^ new_n7951;
  assign new_n8030 = new_n8009 ^ new_n7998;
  assign new_n8031 = new_n7930 ^ new_n7816;
  assign new_n8032 = new_n7991 ^ new_n7934;
  assign new_n8033 = new_n8013 ^ new_n7996;
  assign new_n8034 = ~new_n8033 & new_n8020;
  assign new_n8035 = new_n8034 ^ new_n8020;
  assign new_n8036 = new_n8022 ^ new_n8000;
  assign new_n8037 = new_n8036 ^ new_n8005;
  assign new_n8038 = new_n8034 ^ new_n7996;
  assign new_n8039 = ~new_n8037 & new_n8038;
  assign new_n8040 = new_n8039 ^ new_n8035;
  assign new_n8041 = new_n8040 ^ new_n8032;
  assign new_n8042 = new_n8041 ^ new_n8031;
  assign new_n8043 = new_n8042 ^ new_n8030;
  assign new_n8044 = new_n8043 ^ new_n8029;
  assign new_n8045 = new_n7955 & new_n8044;
  assign new_n8046 = ~new_n8007 & ~new_n8037;
  assign new_n8047 = ~new_n8002 & new_n8044;
  assign new_n8048 = new_n8047 ^ new_n8046;
  assign new_n8049 = new_n8035 ^ new_n7981;
  assign new_n8050 = ~new_n7982 & ~new_n8049;
  assign new_n8051 = new_n8020 ^ new_n8013;
  assign new_n8052 = ~new_n7906 & new_n8051;
  assign new_n8053 = new_n8052 ^ new_n8050;
  assign new_n8054 = new_n8039 ^ new_n8022;
  assign new_n8055 = new_n8054 ^ new_n7995;
  assign new_n8056 = ~new_n7952 & new_n8055;
  assign new_n8057 = new_n8056 ^ new_n8053;
  assign new_n8058 = new_n8057 ^ new_n8048;
  assign new_n8059 = new_n8058 ^ new_n8045;
  assign new_n8060 = new_n8059 ^ new_n8028;
  assign new_n8061 = new_n7592 ^ new_n1160;
  assign new_n8062 = new_n8061 ^ n116;
  assign new_n8063 = new_n5612 ^ new_n5560;
  assign new_n8064 = new_n8063 ^ new_n8062;
  assign new_n8065 = new_n8064 ^ new_n5594;
  assign new_n8066 = new_n5584 ^ new_n5513;
  assign new_n8067 = new_n8066 ^ new_n5654;
  assign new_n8068 = new_n8067 ^ new_n8065;
  assign new_n8069 = new_n5540 ^ new_n5173;
  assign new_n8070 = new_n5601 ^ new_n5513;
  assign new_n8071 = new_n7573 ^ new_n1138;
  assign new_n8072 = new_n8071 ^ n115;
  assign new_n8073 = new_n8072 ^ new_n8070;
  assign new_n8074 = new_n8073 ^ new_n8069;
  assign new_n8075 = new_n5470 ^ new_n5173;
  assign new_n8076 = new_n7539 ^ new_n1116;
  assign new_n8077 = new_n8076 ^ new_n5492;
  assign new_n8078 = new_n8077 ^ new_n5616;
  assign new_n8079 = new_n8078 ^ new_n8075;
  assign new_n8080 = new_n8079 ^ new_n8074;
  assign new_n8081 = new_n7647 ^ new_n1152;
  assign new_n8082 = new_n8081 ^ new_n5552;
  assign new_n8083 = new_n8063 ^ new_n5640;
  assign new_n8084 = new_n8083 ^ new_n8082;
  assign new_n8085 = new_n8084 ^ new_n8080;
  assign new_n8086 = new_n8085 ^ new_n8068;
  assign new_n8087 = new_n5645 ^ new_n5628;
  assign new_n8088 = new_n8087 ^ new_n8063;
  assign new_n8089 = new_n7463 ^ new_n1180;
  assign new_n8090 = new_n8089 ^ new_n5677;
  assign new_n8091 = new_n5639 ^ new_n5575;
  assign new_n8092 = new_n8091 ^ new_n8090;
  assign new_n8093 = new_n8092 ^ new_n8088;
  assign new_n8094 = new_n8085 & new_n8093;
  assign new_n8095 = new_n8094 ^ new_n8093;
  assign new_n8096 = new_n5621 ^ new_n5616;
  assign new_n8097 = new_n6842 ^ new_n1187;
  assign new_n8098 = new_n8097 ^ n113;
  assign new_n8099 = new_n8098 ^ new_n5560;
  assign new_n8100 = new_n8099 ^ new_n5037;
  assign new_n8101 = new_n8100 ^ new_n8096;
  assign new_n8102 = new_n8101 ^ new_n8093;
  assign new_n8103 = new_n5662 ^ new_n5584;
  assign new_n8104 = new_n8103 ^ new_n5687;
  assign new_n8105 = new_n7621 ^ new_n1171;
  assign new_n8106 = new_n8105 ^ n117;
  assign new_n8107 = new_n8106 ^ new_n8063;
  assign new_n8108 = new_n8107 ^ new_n5668;
  assign new_n8109 = new_n8108 ^ new_n8104;
  assign new_n8110 = new_n8109 ^ new_n8093;
  assign new_n8111 = new_n1198 ^ new_n1011;
  assign new_n8112 = new_n8111 ^ n118;
  assign new_n8113 = new_n8112 ^ new_n5662;
  assign new_n8114 = new_n8113 ^ new_n5632;
  assign new_n8115 = new_n8114 ^ new_n5682;
  assign new_n8116 = new_n8115 ^ new_n8110;
  assign new_n8117 = new_n8116 ^ new_n8074;
  assign new_n8118 = ~new_n8102 & new_n8117;
  assign new_n8119 = new_n8118 ^ new_n8095;
  assign new_n8120 = new_n8115 ^ new_n8101;
  assign new_n8121 = new_n8120 ^ new_n8119;
  assign new_n8122 = new_n8074 ^ new_n8068;
  assign new_n8123 = new_n8122 ^ new_n8120;
  assign new_n8124 = new_n8115 ^ new_n8068;
  assign new_n8125 = ~new_n8123 & new_n8124;
  assign new_n8126 = new_n8116 ^ new_n8079;
  assign new_n8127 = new_n8101 ^ new_n8068;
  assign new_n8128 = new_n8126 & new_n8127;
  assign new_n8129 = new_n8128 ^ new_n8125;
  assign new_n8130 = new_n8109 ^ new_n8074;
  assign new_n8131 = new_n8130 ^ new_n8129;
  assign new_n8132 = new_n8131 ^ new_n8121;
  assign new_n8133 = new_n8127 ^ new_n8110;
  assign new_n8134 = new_n8093 ^ new_n8068;
  assign new_n8135 = new_n8134 ^ new_n8120;
  assign new_n8136 = ~new_n8133 & ~new_n8135;
  assign new_n8137 = new_n8136 ^ new_n8079;
  assign new_n8138 = new_n8137 ^ new_n8133;
  assign new_n8139 = new_n8133 ^ new_n8084;
  assign new_n8140 = new_n8093 ^ new_n8085;
  assign new_n8141 = new_n8140 ^ new_n8120;
  assign new_n8142 = new_n8139 & new_n8141;
  assign new_n8143 = new_n8142 ^ new_n8129;
  assign new_n8144 = new_n8143 ^ new_n8115;
  assign new_n8145 = new_n8144 ^ new_n8138;
  assign new_n8146 = ~new_n8132 & new_n8145;
  assign new_n8147 = ~new_n8084 & ~new_n8086;
  assign new_n8148 = new_n8147 ^ new_n8068;
  assign new_n8149 = new_n8148 ^ new_n8137;
  assign new_n8150 = new_n8149 ^ new_n8146;
  assign new_n8151 = new_n8133 ^ new_n8080;
  assign new_n8152 = ~new_n8151 & new_n8120;
  assign new_n8153 = new_n8152 ^ new_n8128;
  assign new_n8154 = new_n8153 ^ new_n8117;
  assign new_n8155 = new_n8154 ^ new_n8150;
  assign new_n8156 = new_n8101 ^ new_n8085;
  assign new_n8157 = new_n8126 ^ new_n8084;
  assign new_n8158 = ~new_n8156 & ~new_n8157;
  assign new_n8159 = new_n8158 ^ new_n8094;
  assign new_n8160 = new_n8152 ^ new_n8125;
  assign new_n8161 = new_n8160 ^ new_n8159;
  assign new_n8162 = ~new_n8155 & ~new_n8161;
  assign new_n8163 = new_n8158 ^ new_n8118;
  assign new_n8164 = new_n8163 ^ new_n8101;
  assign new_n8165 = new_n8164 ^ new_n8154;
  assign new_n8166 = new_n8165 ^ new_n8162;
  assign new_n8167 = ~new_n8086 & new_n8166;
  assign new_n8168 = new_n8093 ^ new_n8074;
  assign new_n8169 = new_n8142 ^ new_n8095;
  assign new_n8170 = new_n8162 ^ new_n8146;
  assign new_n8171 = ~new_n8165 & ~new_n8170;
  assign new_n8172 = new_n8171 ^ new_n8162;
  assign new_n8173 = new_n8165 ^ new_n8146;
  assign new_n8174 = new_n8101 ^ new_n8074;
  assign new_n8175 = new_n8147 ^ new_n8142;
  assign new_n8176 = new_n8175 ^ new_n8160;
  assign new_n8177 = new_n8176 ^ new_n8174;
  assign new_n8178 = ~new_n8177 & new_n8173;
  assign new_n8179 = new_n8178 ^ new_n8149;
  assign new_n8180 = new_n8179 ^ new_n8154;
  assign new_n8181 = ~new_n8172 & ~new_n8180;
  assign new_n8182 = new_n8173 ^ new_n8172;
  assign new_n8183 = new_n8182 ^ new_n8181;
  assign new_n8184 = new_n8183 ^ new_n8169;
  assign new_n8185 = new_n8184 ^ new_n8168;
  assign new_n8186 = new_n8185 ^ new_n8068;
  assign new_n8187 = new_n8178 ^ new_n8118;
  assign new_n8188 = new_n8187 ^ new_n8137;
  assign new_n8189 = new_n8188 ^ new_n8186;
  assign new_n8190 = ~new_n8123 & new_n8189;
  assign new_n8191 = new_n8181 ^ new_n8177;
  assign new_n8192 = ~new_n8085 & ~new_n8191;
  assign new_n8193 = new_n8124 & new_n8189;
  assign new_n8194 = new_n8178 ^ new_n8162;
  assign new_n8195 = new_n8164 ^ new_n8149;
  assign new_n8196 = new_n8195 ^ new_n8194;
  assign new_n8197 = ~new_n8196 & new_n8127;
  assign new_n8198 = new_n8197 ^ new_n8193;
  assign new_n8199 = new_n8182 ^ new_n8162;
  assign new_n8200 = new_n8199 ^ new_n8161;
  assign new_n8201 = new_n8141 & new_n8200;
  assign new_n8202 = new_n8201 ^ new_n8198;
  assign new_n8203 = new_n8202 ^ new_n8192;
  assign new_n8204 = new_n8181 ^ new_n8178;
  assign new_n8205 = new_n8204 ^ new_n8145;
  assign new_n8206 = new_n8117 & new_n8205;
  assign new_n8207 = new_n8206 ^ new_n8203;
  assign new_n8208 = new_n8207 ^ new_n8190;
  assign new_n8209 = new_n8208 ^ new_n8167;
  assign new_n8210 = ~new_n8156 & ~new_n8180;
  assign new_n8211 = new_n8162 ^ new_n8101;
  assign new_n8212 = new_n8158 ^ new_n8147;
  assign new_n8213 = new_n8212 ^ new_n8185;
  assign new_n8214 = new_n8213 ^ new_n8211;
  assign new_n8215 = ~new_n8151 & ~new_n8214;
  assign new_n8216 = new_n8215 ^ new_n8210;
  assign new_n8217 = new_n8182 ^ new_n8132;
  assign new_n8218 = ~new_n8133 & new_n8217;
  assign new_n8219 = ~new_n8084 & new_n8166;
  assign new_n8220 = new_n8219 ^ new_n8218;
  assign new_n8221 = ~new_n8102 & new_n8205;
  assign new_n8222 = new_n8221 ^ new_n8220;
  assign new_n8223 = new_n8222 ^ new_n8216;
  assign new_n8224 = new_n8223 ^ new_n8209;
  assign new_n8225 = new_n6575 ^ n2;
  assign new_n8226 = new_n6564 ^ n67;
  assign new_n8227 = new_n8226 ^ n3;
  assign new_n8228 = new_n8227 ^ new_n8225;
  assign new_n8229 = new_n6630 ^ n8;
  assign new_n8230 = new_n8229 ^ new_n8228;
  assign new_n8231 = new_n6680 ^ n1;
  assign new_n8232 = new_n8231 ^ new_n8230;
  assign new_n8233 = new_n6660 ^ n7;
  assign new_n8234 = new_n6705 ^ n69;
  assign new_n8235 = new_n8234 ^ n5;
  assign new_n8236 = new_n8235 ^ new_n8233;
  assign new_n8237 = new_n6184 ^ n68;
  assign new_n8238 = new_n8237 ^ n4;
  assign new_n8239 = new_n8238 ^ new_n8231;
  assign new_n8240 = new_n8239 ^ new_n8236;
  assign new_n8241 = new_n8238 ^ new_n8233;
  assign new_n8242 = new_n6726 ^ n6;
  assign new_n8243 = new_n8242 ^ new_n8231;
  assign new_n8244 = new_n8243 ^ new_n8241;
  assign new_n8245 = ~new_n8240 & ~new_n8244;
  assign new_n8246 = new_n8245 ^ new_n8225;
  assign new_n8247 = new_n8246 ^ new_n8240;
  assign new_n8248 = new_n8238 ^ new_n8227;
  assign new_n8249 = new_n8248 ^ new_n8243;
  assign new_n8250 = new_n8242 ^ new_n8238;
  assign new_n8251 = ~new_n8249 & new_n8250;
  assign new_n8252 = new_n8242 ^ new_n8236;
  assign new_n8253 = new_n8252 ^ new_n8225;
  assign new_n8254 = new_n8239 & new_n8253;
  assign new_n8255 = new_n8254 ^ new_n8251;
  assign new_n8256 = new_n8240 ^ new_n8229;
  assign new_n8257 = new_n8233 ^ new_n8230;
  assign new_n8258 = new_n8257 ^ new_n8243;
  assign new_n8259 = new_n8256 & new_n8258;
  assign new_n8260 = new_n8259 ^ new_n8242;
  assign new_n8261 = new_n8260 ^ new_n8255;
  assign new_n8262 = new_n8261 ^ new_n8247;
  assign new_n8263 = new_n8230 & new_n8233;
  assign new_n8264 = new_n8263 ^ new_n8233;
  assign new_n8265 = new_n8252 ^ new_n8227;
  assign new_n8266 = new_n8233 ^ new_n8231;
  assign new_n8267 = ~new_n8266 & new_n8265;
  assign new_n8268 = new_n8267 ^ new_n8264;
  assign new_n8269 = new_n8268 ^ new_n8243;
  assign new_n8270 = new_n8235 ^ new_n8227;
  assign new_n8271 = new_n8270 ^ new_n8255;
  assign new_n8272 = new_n8271 ^ new_n8269;
  assign new_n8273 = ~new_n8272 & new_n8262;
  assign new_n8274 = new_n8240 ^ new_n8228;
  assign new_n8275 = ~new_n8274 & new_n8243;
  assign new_n8276 = new_n8275 ^ new_n8254;
  assign new_n8277 = new_n8276 ^ new_n8265;
  assign new_n8278 = new_n8253 ^ new_n8229;
  assign new_n8279 = ~new_n8232 & ~new_n8278;
  assign new_n8280 = new_n8279 ^ new_n8267;
  assign new_n8281 = new_n8280 ^ new_n8231;
  assign new_n8282 = new_n8281 ^ new_n8277;
  assign new_n8283 = new_n8282 ^ new_n8273;
  assign new_n8284 = new_n8231 ^ new_n8227;
  assign new_n8285 = new_n8238 ^ new_n8230;
  assign new_n8286 = ~new_n8229 & ~new_n8285;
  assign new_n8287 = new_n8286 ^ new_n8259;
  assign new_n8288 = new_n8275 ^ new_n8251;
  assign new_n8289 = new_n8288 ^ new_n8287;
  assign new_n8290 = new_n8289 ^ new_n8284;
  assign new_n8291 = ~new_n8290 & new_n8283;
  assign new_n8292 = new_n8286 ^ new_n8238;
  assign new_n8293 = new_n8292 ^ new_n8246;
  assign new_n8294 = new_n8293 ^ new_n8291;
  assign new_n8295 = new_n8294 ^ new_n8277;
  assign new_n8296 = ~new_n8232 & ~new_n8295;
  assign new_n8297 = new_n8293 ^ new_n8273;
  assign new_n8298 = new_n8297 ^ new_n8277;
  assign new_n8299 = new_n8279 ^ new_n8263;
  assign new_n8300 = new_n8299 ^ new_n8288;
  assign new_n8301 = ~new_n8298 & ~new_n8300;
  assign new_n8302 = new_n8301 ^ new_n8231;
  assign new_n8303 = new_n8286 ^ new_n8279;
  assign new_n8304 = new_n8233 ^ new_n8227;
  assign new_n8305 = new_n8264 ^ new_n8259;
  assign new_n8306 = new_n8301 ^ new_n8273;
  assign new_n8307 = ~new_n8282 & ~new_n8306;
  assign new_n8308 = new_n8307 ^ new_n8301;
  assign new_n8309 = ~new_n8295 & ~new_n8308;
  assign new_n8310 = new_n8308 ^ new_n8283;
  assign new_n8311 = new_n8310 ^ new_n8309;
  assign new_n8312 = new_n8311 ^ new_n8305;
  assign new_n8313 = new_n8312 ^ new_n8304;
  assign new_n8314 = new_n8313 ^ new_n8303;
  assign new_n8315 = new_n8314 ^ new_n8302;
  assign new_n8316 = ~new_n8274 & ~new_n8315;
  assign new_n8317 = new_n8316 ^ new_n8296;
  assign new_n8318 = new_n8301 ^ new_n8282;
  assign new_n8319 = ~new_n8229 & new_n8318;
  assign new_n8320 = new_n8310 ^ new_n8272;
  assign new_n8321 = ~new_n8240 & new_n8320;
  assign new_n8322 = new_n8321 ^ new_n8319;
  assign new_n8323 = new_n8309 ^ new_n8291;
  assign new_n8324 = new_n8323 ^ new_n8262;
  assign new_n8325 = ~new_n8266 & new_n8324;
  assign new_n8326 = new_n8325 ^ new_n8322;
  assign new_n8327 = new_n8326 ^ new_n8317;
  assign new_n8328 = ~new_n8285 & new_n8318;
  assign new_n8329 = new_n8313 ^ new_n8238;
  assign new_n8330 = new_n8291 ^ new_n8267;
  assign new_n8331 = new_n8330 ^ new_n8246;
  assign new_n8332 = new_n8331 ^ new_n8329;
  assign new_n8333 = ~new_n8249 & new_n8332;
  assign new_n8334 = new_n8309 ^ new_n8290;
  assign new_n8335 = ~new_n8230 & ~new_n8334;
  assign new_n8336 = new_n8250 & new_n8332;
  assign new_n8337 = new_n8301 ^ new_n8291;
  assign new_n8338 = new_n8293 ^ new_n8281;
  assign new_n8339 = new_n8338 ^ new_n8337;
  assign new_n8340 = ~new_n8339 & new_n8239;
  assign new_n8341 = new_n8340 ^ new_n8336;
  assign new_n8342 = new_n8310 ^ new_n8301;
  assign new_n8343 = new_n8342 ^ new_n8300;
  assign new_n8344 = new_n8258 & new_n8343;
  assign new_n8345 = new_n8344 ^ new_n8341;
  assign new_n8346 = new_n8345 ^ new_n8335;
  assign new_n8347 = new_n8265 & new_n8324;
  assign new_n8348 = new_n8347 ^ new_n8346;
  assign new_n8349 = new_n8348 ^ new_n8333;
  assign new_n8350 = new_n8349 ^ new_n8328;
  assign new_n8351 = new_n8350 ^ new_n8327;
  assign new_n8352 = new_n8351 ^ n46;
  assign new_n8353 = new_n8352 ^ n14;
  assign new_n8354 = new_n8353 ^ new_n8224;
  assign new_n8355 = new_n4653 ^ new_n4626;
  assign new_n8356 = new_n8355 ^ new_n4573;
  assign new_n8357 = new_n6574 ^ new_n430;
  assign new_n8358 = new_n8357 ^ n34;
  assign new_n8359 = new_n8358 ^ new_n4736;
  assign new_n8360 = new_n8359 ^ new_n4649;
  assign new_n8361 = new_n8360 ^ new_n8356;
  assign new_n8362 = new_n4589 ^ new_n4555;
  assign new_n8363 = new_n8362 ^ new_n4649;
  assign new_n8364 = new_n6564 ^ new_n441;
  assign new_n8365 = new_n8364 ^ n35;
  assign new_n8366 = new_n4594 ^ new_n2929;
  assign new_n8367 = new_n8366 ^ new_n8365;
  assign new_n8368 = new_n8367 ^ new_n8363;
  assign new_n8369 = new_n8368 ^ new_n8361;
  assign new_n8370 = new_n6629 ^ new_n410;
  assign new_n8371 = new_n8370 ^ n40;
  assign new_n8372 = new_n8371 ^ new_n4709;
  assign new_n8373 = new_n4721 ^ new_n3755;
  assign new_n8374 = new_n4682 ^ new_n4669;
  assign new_n8375 = new_n8374 ^ new_n8373;
  assign new_n8376 = new_n8375 ^ new_n8372;
  assign new_n8377 = new_n8376 ^ new_n8369;
  assign new_n8378 = new_n6184 ^ new_n370;
  assign new_n8379 = new_n8378 ^ n100;
  assign new_n8380 = new_n8379 ^ n36;
  assign new_n8381 = new_n4519 ^ new_n2169;
  assign new_n8382 = new_n8381 ^ new_n8380;
  assign new_n8383 = new_n8382 ^ new_n8373;
  assign new_n8384 = new_n4781 ^ new_n4594;
  assign new_n8385 = new_n8384 ^ new_n4535;
  assign new_n8386 = new_n8385 ^ new_n8383;
  assign new_n8387 = new_n8386 ^ new_n8377;
  assign new_n8388 = ~new_n8376 & ~new_n8387;
  assign new_n8389 = new_n8388 ^ new_n8386;
  assign new_n8390 = new_n8373 ^ new_n4676;
  assign new_n8391 = new_n4714 ^ new_n4695;
  assign new_n8392 = new_n8391 ^ new_n8390;
  assign new_n8393 = new_n6659 ^ new_n390;
  assign new_n8394 = new_n8393 ^ n39;
  assign new_n8395 = new_n8394 ^ new_n4762;
  assign new_n8396 = new_n8395 ^ new_n4709;
  assign new_n8397 = new_n8396 ^ new_n8392;
  assign new_n8398 = new_n4745 ^ new_n4535;
  assign new_n8399 = new_n8398 ^ new_n4769;
  assign new_n8400 = new_n6705 ^ new_n399;
  assign new_n8401 = new_n8400 ^ n101;
  assign new_n8402 = new_n8401 ^ n37;
  assign new_n8403 = new_n8402 ^ new_n8373;
  assign new_n8404 = new_n4785 ^ new_n4526;
  assign new_n8405 = new_n8404 ^ new_n8403;
  assign new_n8406 = new_n8405 ^ new_n8399;
  assign new_n8407 = new_n8406 ^ new_n8397;
  assign new_n8408 = new_n4724 ^ new_n4512;
  assign new_n8409 = new_n8408 ^ new_n4622;
  assign new_n8410 = new_n6679 ^ new_n6203;
  assign new_n8411 = new_n8410 ^ n33;
  assign new_n8412 = new_n8411 ^ new_n3755;
  assign new_n8413 = new_n8412 ^ new_n4736;
  assign new_n8414 = new_n8413 ^ new_n8409;
  assign new_n8415 = new_n8414 ^ new_n8386;
  assign new_n8416 = new_n8415 ^ new_n8407;
  assign new_n8417 = new_n8414 ^ new_n8397;
  assign new_n8418 = new_n4757 ^ new_n4742;
  assign new_n8419 = new_n8418 ^ new_n4691;
  assign new_n8420 = new_n6725 ^ new_n6200;
  assign new_n8421 = new_n8420 ^ n38;
  assign new_n8422 = new_n8421 ^ new_n4769;
  assign new_n8423 = new_n8422 ^ new_n4762;
  assign new_n8424 = new_n8423 ^ new_n8419;
  assign new_n8425 = new_n8424 ^ new_n8386;
  assign new_n8426 = new_n8425 ^ new_n8417;
  assign new_n8427 = ~new_n8416 & ~new_n8426;
  assign new_n8428 = new_n8427 ^ new_n8361;
  assign new_n8429 = new_n8428 ^ new_n8389;
  assign new_n8430 = new_n8424 ^ new_n8407;
  assign new_n8431 = new_n8430 ^ new_n8368;
  assign new_n8432 = ~new_n8417 & new_n8431;
  assign new_n8433 = new_n8377 & new_n8397;
  assign new_n8434 = new_n8433 ^ new_n8397;
  assign new_n8435 = new_n8434 ^ new_n8432;
  assign new_n8436 = new_n8424 ^ new_n8414;
  assign new_n8437 = new_n8436 ^ new_n8435;
  assign new_n8438 = new_n8430 ^ new_n8361;
  assign new_n8439 = new_n8415 & new_n8438;
  assign new_n8440 = new_n8386 ^ new_n8368;
  assign new_n8441 = new_n8440 ^ new_n8436;
  assign new_n8442 = ~new_n8441 & new_n8425;
  assign new_n8443 = new_n8442 ^ new_n8439;
  assign new_n8444 = new_n8406 ^ new_n8368;
  assign new_n8445 = new_n8444 ^ new_n8443;
  assign new_n8446 = new_n8445 ^ new_n8437;
  assign new_n8447 = new_n8428 ^ new_n8416;
  assign new_n8448 = new_n8416 ^ new_n8376;
  assign new_n8449 = new_n8397 ^ new_n8377;
  assign new_n8450 = new_n8449 ^ new_n8436;
  assign new_n8451 = new_n8448 & new_n8450;
  assign new_n8452 = new_n8451 ^ new_n8443;
  assign new_n8453 = new_n8452 ^ new_n8424;
  assign new_n8454 = new_n8453 ^ new_n8447;
  assign new_n8455 = ~new_n8446 & new_n8454;
  assign new_n8456 = new_n8455 ^ new_n8429;
  assign new_n8457 = new_n8416 ^ new_n8369;
  assign new_n8458 = ~new_n8457 & new_n8436;
  assign new_n8459 = new_n8458 ^ new_n8439;
  assign new_n8460 = new_n8459 ^ new_n8431;
  assign new_n8461 = new_n8460 ^ new_n8456;
  assign new_n8462 = new_n8458 ^ new_n8442;
  assign new_n8463 = new_n8414 ^ new_n8377;
  assign new_n8464 = new_n8438 ^ new_n8376;
  assign new_n8465 = ~new_n8463 & ~new_n8464;
  assign new_n8466 = new_n8465 ^ new_n8433;
  assign new_n8467 = new_n8466 ^ new_n8462;
  assign new_n8468 = ~new_n8461 & ~new_n8467;
  assign new_n8469 = new_n8465 ^ new_n8432;
  assign new_n8470 = new_n8469 ^ new_n8414;
  assign new_n8471 = new_n8470 ^ new_n8460;
  assign new_n8472 = new_n8471 ^ new_n8468;
  assign new_n8473 = ~new_n8387 & new_n8472;
  assign new_n8474 = new_n8468 ^ new_n8455;
  assign new_n8475 = ~new_n8471 & ~new_n8474;
  assign new_n8476 = new_n8475 ^ new_n8468;
  assign new_n8477 = new_n8471 ^ new_n8455;
  assign new_n8478 = new_n8414 ^ new_n8368;
  assign new_n8479 = new_n8451 ^ new_n8388;
  assign new_n8480 = new_n8479 ^ new_n8462;
  assign new_n8481 = new_n8480 ^ new_n8478;
  assign new_n8482 = ~new_n8481 & new_n8477;
  assign new_n8483 = new_n8482 ^ new_n8429;
  assign new_n8484 = new_n8483 ^ new_n8460;
  assign new_n8485 = ~new_n8476 & ~new_n8484;
  assign new_n8486 = new_n8485 ^ new_n8482;
  assign new_n8487 = new_n8486 ^ new_n8454;
  assign new_n8488 = new_n8431 & new_n8487;
  assign new_n8489 = new_n8485 ^ new_n8481;
  assign new_n8490 = ~new_n8377 & ~new_n8489;
  assign new_n8491 = new_n8482 ^ new_n8468;
  assign new_n8492 = new_n8470 ^ new_n8429;
  assign new_n8493 = new_n8492 ^ new_n8491;
  assign new_n8494 = ~new_n8493 & new_n8415;
  assign new_n8495 = new_n8397 ^ new_n8368;
  assign new_n8496 = new_n8451 ^ new_n8434;
  assign new_n8497 = new_n8477 ^ new_n8476;
  assign new_n8498 = new_n8497 ^ new_n8485;
  assign new_n8499 = new_n8498 ^ new_n8496;
  assign new_n8500 = new_n8499 ^ new_n8495;
  assign new_n8501 = new_n8500 ^ new_n8386;
  assign new_n8502 = new_n8482 ^ new_n8432;
  assign new_n8503 = new_n8502 ^ new_n8428;
  assign new_n8504 = new_n8503 ^ new_n8501;
  assign new_n8505 = new_n8425 & new_n8504;
  assign new_n8506 = new_n8505 ^ new_n8494;
  assign new_n8507 = new_n8497 ^ new_n8468;
  assign new_n8508 = new_n8507 ^ new_n8467;
  assign new_n8509 = new_n8450 & new_n8508;
  assign new_n8510 = new_n8509 ^ new_n8506;
  assign new_n8511 = new_n8510 ^ new_n8490;
  assign new_n8512 = new_n8511 ^ new_n8488;
  assign new_n8513 = ~new_n8441 & new_n8504;
  assign new_n8514 = new_n8513 ^ new_n8512;
  assign new_n8515 = new_n8514 ^ new_n8473;
  assign new_n8516 = ~new_n8463 & ~new_n8484;
  assign new_n8517 = new_n8468 ^ new_n8414;
  assign new_n8518 = new_n8465 ^ new_n8388;
  assign new_n8519 = new_n8518 ^ new_n8500;
  assign new_n8520 = new_n8519 ^ new_n8517;
  assign new_n8521 = ~new_n8457 & ~new_n8520;
  assign new_n8522 = new_n8521 ^ new_n8516;
  assign new_n8523 = new_n8497 ^ new_n8446;
  assign new_n8524 = ~new_n8416 & new_n8523;
  assign new_n8525 = ~new_n8376 & new_n8472;
  assign new_n8526 = new_n8525 ^ new_n8524;
  assign new_n8527 = ~new_n8417 & new_n8487;
  assign new_n8528 = new_n8527 ^ new_n8526;
  assign new_n8529 = new_n8528 ^ new_n8522;
  assign new_n8530 = new_n8529 ^ new_n8515;
  assign new_n8531 = new_n7423 ^ new_n6981;
  assign new_n8532 = new_n1295 ^ n92;
  assign new_n8533 = new_n8532 ^ n28;
  assign new_n8534 = new_n8533 ^ new_n8531;
  assign new_n8535 = new_n8534 ^ new_n7597;
  assign new_n8536 = new_n7628 ^ new_n7581;
  assign new_n8537 = new_n8536 ^ new_n7602;
  assign new_n8538 = new_n8537 ^ new_n8535;
  assign new_n8539 = new_n7588 ^ new_n7555;
  assign new_n8540 = new_n7608 ^ new_n7581;
  assign new_n8541 = new_n4613 ^ n91;
  assign new_n8542 = new_n8541 ^ n27;
  assign new_n8543 = new_n8542 ^ new_n8540;
  assign new_n8544 = new_n8543 ^ new_n8539;
  assign new_n8545 = new_n7579 ^ new_n7567;
  assign new_n8546 = new_n4632 ^ n90;
  assign new_n8547 = new_n8546 ^ n26;
  assign new_n8548 = new_n8547 ^ new_n7252;
  assign new_n8549 = new_n8548 ^ new_n7555;
  assign new_n8550 = new_n8549 ^ new_n8545;
  assign new_n8551 = new_n8550 ^ new_n8544;
  assign new_n8552 = new_n4662 ^ n96;
  assign new_n8553 = new_n8552 ^ n32;
  assign new_n8554 = new_n8553 ^ new_n7417;
  assign new_n8555 = new_n7654 ^ new_n7486;
  assign new_n8556 = new_n8555 ^ new_n8531;
  assign new_n8557 = new_n8556 ^ new_n8554;
  assign new_n8558 = new_n8557 ^ new_n8551;
  assign new_n8559 = new_n8558 ^ new_n8538;
  assign new_n8560 = new_n8531 ^ new_n7652;
  assign new_n8561 = new_n7479 ^ new_n7453;
  assign new_n8562 = new_n8561 ^ new_n8560;
  assign new_n8563 = new_n4702 ^ n95;
  assign new_n8564 = new_n8563 ^ n31;
  assign new_n8565 = new_n8564 ^ new_n7521;
  assign new_n8566 = new_n8565 ^ new_n7417;
  assign new_n8567 = new_n8566 ^ new_n8562;
  assign new_n8568 = ~new_n8558 & new_n8567;
  assign new_n8569 = new_n8568 ^ new_n8567;
  assign new_n8570 = new_n7547 ^ new_n7400;
  assign new_n8571 = new_n4729 ^ n89;
  assign new_n8572 = new_n8571 ^ n25;
  assign new_n8573 = new_n8572 ^ new_n7423;
  assign new_n8574 = new_n8573 ^ new_n7252;
  assign new_n8575 = new_n8574 ^ new_n8570;
  assign new_n8576 = new_n8575 ^ new_n8567;
  assign new_n8577 = new_n7602 ^ new_n7500;
  assign new_n8578 = new_n8577 ^ new_n7616;
  assign new_n8579 = new_n7632 ^ new_n7606;
  assign new_n8580 = new_n4774 ^ n93;
  assign new_n8581 = new_n8580 ^ n29;
  assign new_n8582 = new_n8581 ^ new_n8579;
  assign new_n8583 = new_n8582 ^ new_n8531;
  assign new_n8584 = new_n8583 ^ new_n8578;
  assign new_n8585 = new_n8584 ^ new_n8567;
  assign new_n8586 = new_n7529 ^ new_n7511;
  assign new_n8587 = new_n8586 ^ new_n7439;
  assign new_n8588 = new_n4750 ^ n94;
  assign new_n8589 = new_n8588 ^ n30;
  assign new_n8590 = new_n8589 ^ new_n7616;
  assign new_n8591 = new_n8590 ^ new_n7521;
  assign new_n8592 = new_n8591 ^ new_n8587;
  assign new_n8593 = new_n8592 ^ new_n8585;
  assign new_n8594 = new_n8593 ^ new_n8544;
  assign new_n8595 = ~new_n8576 & ~new_n8594;
  assign new_n8596 = new_n8595 ^ new_n8569;
  assign new_n8597 = new_n8592 ^ new_n8575;
  assign new_n8598 = new_n8597 ^ new_n8596;
  assign new_n8599 = new_n8592 ^ new_n8538;
  assign new_n8600 = new_n8544 ^ new_n8538;
  assign new_n8601 = new_n8600 ^ new_n8597;
  assign new_n8602 = new_n8599 & new_n8601;
  assign new_n8603 = new_n8593 ^ new_n8550;
  assign new_n8604 = new_n8575 ^ new_n8538;
  assign new_n8605 = ~new_n8603 & new_n8604;
  assign new_n8606 = new_n8605 ^ new_n8602;
  assign new_n8607 = new_n8584 ^ new_n8544;
  assign new_n8608 = new_n8607 ^ new_n8606;
  assign new_n8609 = new_n8608 ^ new_n8598;
  assign new_n8610 = new_n8604 ^ new_n8585;
  assign new_n8611 = new_n8567 ^ new_n8538;
  assign new_n8612 = new_n8611 ^ new_n8597;
  assign new_n8613 = ~new_n8610 & ~new_n8612;
  assign new_n8614 = new_n8613 ^ new_n8550;
  assign new_n8615 = new_n8614 ^ new_n8610;
  assign new_n8616 = new_n8610 ^ new_n8557;
  assign new_n8617 = new_n8567 ^ new_n8558;
  assign new_n8618 = new_n8617 ^ new_n8597;
  assign new_n8619 = ~new_n8616 & ~new_n8618;
  assign new_n8620 = new_n8619 ^ new_n8606;
  assign new_n8621 = new_n8620 ^ new_n8592;
  assign new_n8622 = new_n8621 ^ new_n8615;
  assign new_n8623 = ~new_n8622 & new_n8609;
  assign new_n8624 = new_n8557 & new_n8559;
  assign new_n8625 = new_n8624 ^ new_n8538;
  assign new_n8626 = new_n8625 ^ new_n8614;
  assign new_n8627 = new_n8626 ^ new_n8623;
  assign new_n8628 = new_n8610 ^ new_n8551;
  assign new_n8629 = ~new_n8628 & new_n8597;
  assign new_n8630 = new_n8629 ^ new_n8605;
  assign new_n8631 = new_n8630 ^ new_n8594;
  assign new_n8632 = new_n8631 ^ new_n8627;
  assign new_n8633 = new_n8575 ^ new_n8558;
  assign new_n8634 = new_n8603 ^ new_n8557;
  assign new_n8635 = ~new_n8634 & new_n8633;
  assign new_n8636 = new_n8635 ^ new_n8568;
  assign new_n8637 = new_n8629 ^ new_n8602;
  assign new_n8638 = new_n8637 ^ new_n8636;
  assign new_n8639 = ~new_n8632 & ~new_n8638;
  assign new_n8640 = new_n8635 ^ new_n8595;
  assign new_n8641 = new_n8640 ^ new_n8575;
  assign new_n8642 = new_n8641 ^ new_n8631;
  assign new_n8643 = new_n8642 ^ new_n8639;
  assign new_n8644 = ~new_n8643 & new_n8559;
  assign new_n8645 = new_n8567 ^ new_n8544;
  assign new_n8646 = new_n8619 ^ new_n8569;
  assign new_n8647 = new_n8639 ^ new_n8623;
  assign new_n8648 = ~new_n8647 & new_n8642;
  assign new_n8649 = new_n8648 ^ new_n8639;
  assign new_n8650 = new_n8642 ^ new_n8623;
  assign new_n8651 = new_n8575 ^ new_n8544;
  assign new_n8652 = new_n8624 ^ new_n8619;
  assign new_n8653 = new_n8652 ^ new_n8637;
  assign new_n8654 = new_n8653 ^ new_n8651;
  assign new_n8655 = ~new_n8650 & new_n8654;
  assign new_n8656 = new_n8655 ^ new_n8626;
  assign new_n8657 = new_n8656 ^ new_n8631;
  assign new_n8658 = ~new_n8649 & ~new_n8657;
  assign new_n8659 = new_n8650 ^ new_n8649;
  assign new_n8660 = new_n8659 ^ new_n8658;
  assign new_n8661 = new_n8660 ^ new_n8646;
  assign new_n8662 = new_n8661 ^ new_n8645;
  assign new_n8663 = new_n8662 ^ new_n8538;
  assign new_n8664 = new_n8655 ^ new_n8595;
  assign new_n8665 = new_n8664 ^ new_n8614;
  assign new_n8666 = new_n8665 ^ new_n8663;
  assign new_n8667 = ~new_n8666 & new_n8601;
  assign new_n8668 = new_n8658 ^ new_n8654;
  assign new_n8669 = new_n8558 & new_n8668;
  assign new_n8670 = new_n8655 ^ new_n8639;
  assign new_n8671 = new_n8641 ^ new_n8626;
  assign new_n8672 = new_n8671 ^ new_n8670;
  assign new_n8673 = new_n8604 & new_n8672;
  assign new_n8674 = ~new_n8666 & new_n8599;
  assign new_n8675 = new_n8674 ^ new_n8673;
  assign new_n8676 = new_n8659 ^ new_n8639;
  assign new_n8677 = new_n8676 ^ new_n8638;
  assign new_n8678 = ~new_n8618 & ~new_n8677;
  assign new_n8679 = new_n8678 ^ new_n8675;
  assign new_n8680 = new_n8679 ^ new_n8669;
  assign new_n8681 = new_n8658 ^ new_n8655;
  assign new_n8682 = new_n8681 ^ new_n8622;
  assign new_n8683 = ~new_n8594 & ~new_n8682;
  assign new_n8684 = new_n8683 ^ new_n8680;
  assign new_n8685 = new_n8684 ^ new_n8667;
  assign new_n8686 = new_n8685 ^ new_n8644;
  assign new_n8687 = ~new_n8657 & new_n8633;
  assign new_n8688 = new_n8639 ^ new_n8575;
  assign new_n8689 = new_n8635 ^ new_n8624;
  assign new_n8690 = new_n8689 ^ new_n8662;
  assign new_n8691 = new_n8690 ^ new_n8688;
  assign new_n8692 = ~new_n8628 & ~new_n8691;
  assign new_n8693 = new_n8692 ^ new_n8687;
  assign new_n8694 = ~new_n8643 & new_n8557;
  assign new_n8695 = new_n8659 ^ new_n8609;
  assign new_n8696 = ~new_n8610 & new_n8695;
  assign new_n8697 = new_n8696 ^ new_n8694;
  assign new_n8698 = ~new_n8576 & ~new_n8682;
  assign new_n8699 = new_n8698 ^ new_n8697;
  assign new_n8700 = new_n8699 ^ new_n8693;
  assign new_n8701 = new_n8700 ^ new_n8686;
  assign new_n8702 = new_n8701 ^ new_n8530;
  assign new_n8703 = new_n6667 ^ new_n6325;
  assign new_n8704 = new_n8703 ^ new_n6720;
  assign new_n8705 = new_n6648 ^ new_n6616;
  assign new_n8706 = new_n8705 ^ new_n8704;
  assign new_n8707 = new_n6654 ^ new_n6642;
  assign new_n8708 = new_n8707 ^ new_n591;
  assign new_n8709 = new_n8708 ^ new_n8706;
  assign new_n8710 = new_n6674 ^ new_n6584;
  assign new_n8711 = new_n8710 ^ new_n584;
  assign new_n8712 = new_n6670 ^ new_n6462;
  assign new_n8713 = new_n8712 ^ new_n6325;
  assign new_n8714 = new_n8713 ^ new_n8711;
  assign new_n8715 = new_n8714 ^ new_n8709;
  assign new_n8716 = new_n6530 ^ new_n560;
  assign new_n8717 = new_n6492 ^ new_n5934;
  assign new_n8718 = new_n8717 ^ new_n6601;
  assign new_n8719 = new_n8718 ^ new_n8716;
  assign new_n8720 = new_n8719 ^ new_n8714;
  assign new_n8721 = new_n6610 ^ new_n575;
  assign new_n8722 = new_n6648 ^ new_n6623;
  assign new_n8723 = new_n8722 ^ new_n8703;
  assign new_n8724 = new_n8723 ^ new_n8721;
  assign new_n8725 = new_n6696 ^ new_n6472;
  assign new_n8726 = new_n6485 ^ n77;
  assign new_n8727 = new_n8726 ^ new_n8725;
  assign new_n8728 = new_n8703 ^ new_n596;
  assign new_n8729 = new_n6712 ^ new_n6686;
  assign new_n8730 = new_n8729 ^ new_n8728;
  assign new_n8731 = new_n8730 ^ new_n8727;
  assign new_n8732 = new_n8731 ^ new_n8709;
  assign new_n8733 = new_n8703 ^ new_n539;
  assign new_n8734 = new_n6700 ^ new_n6472;
  assign new_n8735 = new_n8734 ^ new_n8733;
  assign new_n8736 = new_n6073 ^ n76;
  assign new_n8737 = new_n8736 ^ new_n6493;
  assign new_n8738 = new_n8737 ^ new_n8735;
  assign new_n8739 = new_n8738 ^ new_n8714;
  assign new_n8740 = new_n8739 ^ new_n8732;
  assign new_n8741 = new_n8740 ^ new_n8724;
  assign new_n8742 = new_n6580 ^ new_n566;
  assign new_n8743 = new_n6600 ^ new_n6512;
  assign new_n8744 = new_n8743 ^ new_n6675;
  assign new_n8745 = new_n8744 ^ new_n8742;
  assign new_n8746 = new_n8745 ^ new_n8719;
  assign new_n8747 = new_n8746 ^ new_n8724;
  assign new_n8748 = new_n8747 ^ new_n8709;
  assign new_n8749 = new_n6715 ^ new_n6686;
  assign new_n8750 = new_n8749 ^ new_n6690;
  assign new_n8751 = new_n6720 ^ new_n6638;
  assign new_n8752 = new_n8751 ^ new_n605;
  assign new_n8753 = new_n8752 ^ new_n8750;
  assign new_n8754 = new_n8753 ^ new_n8714;
  assign new_n8755 = new_n8754 ^ new_n8748;
  assign new_n8756 = new_n8741 & new_n8755;
  assign new_n8757 = new_n8747 ^ new_n8738;
  assign new_n8758 = new_n8724 & new_n8757;
  assign new_n8759 = new_n8758 ^ new_n8756;
  assign new_n8760 = new_n8753 ^ new_n8738;
  assign new_n8761 = new_n8738 ^ new_n8719;
  assign new_n8762 = new_n8761 ^ new_n8754;
  assign new_n8763 = new_n8760 & new_n8762;
  assign new_n8764 = new_n8746 ^ new_n8740;
  assign new_n8765 = new_n8754 & new_n8764;
  assign new_n8766 = new_n8765 ^ new_n8763;
  assign new_n8767 = new_n8766 ^ new_n8759;
  assign new_n8768 = new_n8767 ^ new_n8720;
  assign new_n8769 = ~new_n8709 & ~new_n8747;
  assign new_n8770 = new_n8769 ^ new_n8709;
  assign new_n8771 = new_n8753 ^ new_n8732;
  assign new_n8772 = new_n8771 ^ new_n8719;
  assign new_n8773 = new_n8715 & new_n8772;
  assign new_n8774 = new_n8773 ^ new_n8770;
  assign new_n8775 = new_n8774 ^ new_n8754;
  assign new_n8776 = new_n8771 ^ new_n8745;
  assign new_n8777 = new_n8739 & new_n8776;
  assign new_n8778 = new_n8777 ^ new_n8763;
  assign new_n8779 = new_n8731 ^ new_n8719;
  assign new_n8780 = new_n8779 ^ new_n8778;
  assign new_n8781 = new_n8780 ^ new_n8775;
  assign new_n8782 = new_n8738 ^ new_n8709;
  assign new_n8783 = new_n8782 ^ new_n8754;
  assign new_n8784 = new_n8740 & new_n8783;
  assign new_n8785 = new_n8784 ^ new_n8745;
  assign new_n8786 = new_n8785 ^ new_n8740;
  assign new_n8787 = new_n8778 ^ new_n8756;
  assign new_n8788 = new_n8787 ^ new_n8753;
  assign new_n8789 = new_n8788 ^ new_n8786;
  assign new_n8790 = ~new_n8781 & new_n8789;
  assign new_n8791 = new_n8777 ^ new_n8765;
  assign new_n8792 = new_n8791 ^ new_n8772;
  assign new_n8793 = new_n8747 ^ new_n8714;
  assign new_n8794 = new_n8776 ^ new_n8724;
  assign new_n8795 = new_n8793 & new_n8794;
  assign new_n8796 = new_n8795 ^ new_n8773;
  assign new_n8797 = new_n8796 ^ new_n8714;
  assign new_n8798 = new_n8797 ^ new_n8792;
  assign new_n8799 = new_n8798 ^ new_n8790;
  assign new_n8800 = new_n8768 & new_n8799;
  assign new_n8801 = new_n8758 ^ new_n8738;
  assign new_n8802 = new_n8801 ^ new_n8785;
  assign new_n8803 = new_n8802 ^ new_n8800;
  assign new_n8804 = new_n8803 ^ new_n8792;
  assign new_n8805 = new_n8802 ^ new_n8790;
  assign new_n8806 = new_n8805 ^ new_n8792;
  assign new_n8807 = new_n8795 ^ new_n8769;
  assign new_n8808 = new_n8807 ^ new_n8766;
  assign new_n8809 = ~new_n8808 & new_n8806;
  assign new_n8810 = new_n8809 ^ new_n8790;
  assign new_n8811 = ~new_n8810 & new_n8798;
  assign new_n8812 = new_n8811 ^ new_n8790;
  assign new_n8813 = new_n8804 & new_n8812;
  assign new_n8814 = new_n8813 ^ new_n8800;
  assign new_n8815 = new_n8814 ^ new_n8789;
  assign new_n8816 = new_n8715 & new_n8815;
  assign new_n8817 = new_n8809 ^ new_n8714;
  assign new_n8818 = new_n8795 ^ new_n8758;
  assign new_n8819 = new_n8719 ^ new_n8709;
  assign new_n8820 = new_n8770 ^ new_n8756;
  assign new_n8821 = new_n8811 ^ new_n8798;
  assign new_n8822 = new_n8821 ^ new_n8813;
  assign new_n8823 = new_n8822 ^ new_n8820;
  assign new_n8824 = new_n8823 ^ new_n8819;
  assign new_n8825 = new_n8824 ^ new_n8818;
  assign new_n8826 = new_n8825 ^ new_n8817;
  assign new_n8827 = ~new_n8826 & new_n8764;
  assign new_n8828 = new_n8827 ^ new_n8816;
  assign new_n8829 = new_n8824 ^ new_n8738;
  assign new_n8830 = new_n8800 ^ new_n8773;
  assign new_n8831 = new_n8830 ^ new_n8785;
  assign new_n8832 = new_n8831 ^ new_n8829;
  assign new_n8833 = ~new_n8832 & new_n8762;
  assign new_n8834 = new_n8813 ^ new_n8768;
  assign new_n8835 = new_n8747 & new_n8834;
  assign new_n8836 = new_n8835 ^ new_n8833;
  assign new_n8837 = new_n8748 & new_n8834;
  assign new_n8838 = new_n8794 & new_n8804;
  assign new_n8839 = new_n8838 ^ new_n8837;
  assign new_n8840 = ~new_n8832 & new_n8760;
  assign new_n8841 = new_n8809 ^ new_n8800;
  assign new_n8842 = new_n8802 ^ new_n8797;
  assign new_n8843 = new_n8842 ^ new_n8841;
  assign new_n8844 = new_n8739 & new_n8843;
  assign new_n8845 = new_n8844 ^ new_n8840;
  assign new_n8846 = new_n8845 ^ new_n8839;
  assign new_n8847 = new_n8846 ^ new_n8836;
  assign new_n8848 = new_n8847 ^ new_n8828;
  assign new_n8849 = new_n8527 ^ new_n8521;
  assign new_n8850 = new_n8513 ^ new_n8490;
  assign new_n8851 = ~new_n8489 & new_n8449;
  assign new_n8852 = ~new_n8464 & ~new_n8484;
  assign new_n8853 = new_n8852 ^ new_n8851;
  assign new_n8854 = new_n8853 ^ new_n8506;
  assign new_n8855 = new_n8854 ^ new_n8850;
  assign new_n8856 = new_n8855 ^ new_n8849;
  assign new_n8857 = new_n8856 ^ new_n8848;
  assign new_n8858 = new_n8857 ^ new_n8702;
  assign new_n8859 = new_n8858 ^ new_n8354;
  assign new_n8860 = new_n8698 ^ new_n8692;
  assign new_n8861 = new_n8669 ^ new_n8667;
  assign new_n8862 = ~new_n8617 & new_n8668;
  assign new_n8863 = ~new_n8634 & ~new_n8657;
  assign new_n8864 = new_n8863 ^ new_n8862;
  assign new_n8865 = new_n8864 ^ new_n8675;
  assign new_n8866 = new_n8865 ^ new_n8861;
  assign new_n8867 = new_n8866 ^ new_n8860;
  assign new_n8868 = new_n8867 ^ new_n8856;
  assign new_n8869 = new_n8776 & new_n8843;
  assign new_n8870 = new_n8821 ^ new_n8781;
  assign new_n8871 = ~new_n8870 & new_n8783;
  assign new_n8872 = new_n8871 ^ new_n8869;
  assign new_n8873 = new_n8772 & new_n8815;
  assign new_n8874 = new_n8821 ^ new_n8809;
  assign new_n8875 = new_n8874 ^ new_n8808;
  assign new_n8876 = ~new_n8875 & new_n8755;
  assign new_n8877 = new_n8876 ^ new_n8845;
  assign new_n8878 = new_n8877 ^ new_n8835;
  assign new_n8879 = new_n8878 ^ new_n8873;
  assign new_n8880 = new_n8879 ^ new_n8833;
  assign new_n8881 = new_n8880 ^ new_n8872;
  assign new_n8882 = ~new_n8493 & new_n8438;
  assign new_n8883 = ~new_n8426 & new_n8523;
  assign new_n8884 = new_n8883 ^ new_n8882;
  assign new_n8885 = new_n8884 ^ new_n8514;
  assign new_n8886 = new_n8885 ^ new_n8881;
  assign new_n8887 = new_n8886 ^ new_n8868;
  assign new_n8888 = new_n8221 ^ new_n8215;
  assign new_n8889 = new_n8192 ^ new_n8190;
  assign new_n8890 = ~new_n8191 & new_n8140;
  assign new_n8891 = ~new_n8157 & ~new_n8180;
  assign new_n8892 = new_n8891 ^ new_n8890;
  assign new_n8893 = new_n8892 ^ new_n8198;
  assign new_n8894 = new_n8893 ^ new_n8889;
  assign new_n8895 = new_n8894 ^ new_n8888;
  assign new_n8896 = new_n8325 ^ new_n8316;
  assign new_n8897 = new_n8335 ^ new_n8333;
  assign new_n8898 = ~new_n8334 & new_n8257;
  assign new_n8899 = ~new_n8278 & ~new_n8295;
  assign new_n8900 = new_n8899 ^ new_n8898;
  assign new_n8901 = new_n8900 ^ new_n8341;
  assign new_n8902 = new_n8901 ^ new_n8897;
  assign new_n8903 = new_n8902 ^ new_n8896;
  assign new_n8904 = new_n8903 ^ n47;
  assign new_n8905 = new_n8904 ^ n15;
  assign new_n8906 = new_n8905 ^ new_n8895;
  assign new_n8907 = new_n8528 ^ new_n8488;
  assign new_n8908 = new_n8907 ^ new_n8854;
  assign new_n8909 = ~new_n8870 & new_n8740;
  assign new_n8910 = new_n8809 ^ new_n8798;
  assign new_n8911 = new_n8724 & new_n8910;
  assign new_n8912 = new_n8911 ^ new_n8909;
  assign new_n8913 = new_n8912 ^ new_n8816;
  assign new_n8914 = new_n8913 ^ new_n8873;
  assign new_n8915 = new_n8914 ^ new_n8846;
  assign new_n8916 = new_n8915 ^ new_n8908;
  assign new_n8917 = new_n8916 ^ new_n8906;
  assign new_n8918 = new_n8917 ^ new_n8887;
  assign new_n8919 = ~new_n8135 & new_n8217;
  assign new_n8920 = new_n8919 ^ new_n8891;
  assign new_n8921 = new_n8139 & new_n8200;
  assign new_n8922 = new_n8921 ^ new_n8219;
  assign new_n8923 = new_n8922 ^ new_n8203;
  assign new_n8924 = new_n8923 ^ new_n8920;
  assign new_n8925 = ~new_n8244 & new_n8320;
  assign new_n8926 = new_n8925 ^ new_n8899;
  assign new_n8927 = new_n8256 & new_n8343;
  assign new_n8928 = new_n8927 ^ new_n8319;
  assign new_n8929 = new_n8928 ^ new_n8346;
  assign new_n8930 = new_n8929 ^ new_n8926;
  assign new_n8931 = new_n8930 ^ n45;
  assign new_n8932 = new_n8931 ^ n13;
  assign new_n8933 = new_n8932 ^ new_n8924;
  assign new_n8934 = new_n8757 & new_n8910;
  assign new_n8935 = new_n8934 ^ new_n8880;
  assign new_n8936 = new_n8793 & new_n8804;
  assign new_n8937 = new_n8936 ^ new_n8827;
  assign new_n8938 = new_n8937 ^ new_n8913;
  assign new_n8939 = new_n8938 ^ new_n8935;
  assign new_n8940 = new_n8939 ^ new_n8530;
  assign new_n8941 = new_n8940 ^ new_n8933;
  assign new_n8942 = ~new_n8612 & new_n8695;
  assign new_n8943 = new_n8942 ^ new_n8863;
  assign new_n8944 = ~new_n8616 & ~new_n8677;
  assign new_n8945 = new_n8944 ^ new_n8694;
  assign new_n8946 = new_n8945 ^ new_n8680;
  assign new_n8947 = new_n8946 ^ new_n8943;
  assign new_n8948 = new_n8883 ^ new_n8852;
  assign new_n8949 = new_n8448 & new_n8508;
  assign new_n8950 = new_n8949 ^ new_n8525;
  assign new_n8951 = new_n8950 ^ new_n8511;
  assign new_n8952 = new_n8951 ^ new_n8948;
  assign new_n8953 = new_n8952 ^ new_n8947;
  assign new_n8954 = new_n8953 ^ new_n8886;
  assign new_n8955 = new_n8954 ^ new_n8941;
  assign new_n8956 = new_n8955 ^ new_n8918;
  assign new_n8957 = new_n8956 ^ new_n8859;
  assign new_n8958 = new_n8882 ^ new_n8494;
  assign new_n8959 = ~new_n8520 & new_n8436;
  assign new_n8960 = new_n8959 ^ new_n8529;
  assign new_n8961 = new_n8960 ^ new_n8958;
  assign new_n8962 = new_n8869 ^ new_n8844;
  assign new_n8963 = ~new_n8826 & new_n8754;
  assign new_n8964 = new_n8963 ^ new_n8938;
  assign new_n8965 = new_n8964 ^ new_n8962;
  assign new_n8966 = new_n8965 ^ new_n8961;
  assign new_n8967 = new_n8882 ^ new_n8513;
  assign new_n8968 = new_n8949 ^ new_n8524;
  assign new_n8969 = new_n8968 ^ new_n8883;
  assign new_n8970 = new_n8969 ^ new_n8510;
  assign new_n8971 = new_n8970 ^ new_n8967;
  assign new_n8972 = new_n8971 ^ new_n8966;
  assign new_n8973 = ~new_n8196 & new_n8126;
  assign new_n8974 = new_n8973 ^ new_n8190;
  assign new_n8975 = new_n8921 ^ new_n8218;
  assign new_n8976 = new_n8975 ^ new_n8919;
  assign new_n8977 = new_n8976 ^ new_n8202;
  assign new_n8978 = new_n8977 ^ new_n8974;
  assign new_n8979 = ~new_n8339 & new_n8253;
  assign new_n8980 = new_n8979 ^ new_n8333;
  assign new_n8981 = new_n8927 ^ new_n8321;
  assign new_n8982 = new_n8981 ^ new_n8925;
  assign new_n8983 = new_n8982 ^ new_n8345;
  assign new_n8984 = new_n8983 ^ new_n8980;
  assign new_n8985 = new_n8984 ^ n42;
  assign new_n8986 = new_n8985 ^ n10;
  assign new_n8987 = new_n8986 ^ new_n8978;
  assign new_n8988 = ~new_n8603 & new_n8672;
  assign new_n8989 = new_n8988 ^ new_n8667;
  assign new_n8990 = new_n8944 ^ new_n8696;
  assign new_n8991 = new_n8990 ^ new_n8942;
  assign new_n8992 = new_n8991 ^ new_n8679;
  assign new_n8993 = new_n8992 ^ new_n8989;
  assign new_n8994 = new_n8993 ^ new_n8987;
  assign new_n8995 = new_n8994 ^ new_n8972;
  assign new_n8996 = new_n8995 ^ new_n8957;
  assign new_n8997 = new_n8222 ^ new_n8206;
  assign new_n8998 = new_n8997 ^ new_n8893;
  assign new_n8999 = new_n8347 ^ new_n8326;
  assign new_n9000 = new_n8999 ^ new_n8901;
  assign new_n9001 = new_n9000 ^ n48;
  assign new_n9002 = new_n9001 ^ n16;
  assign new_n9003 = new_n9002 ^ new_n8998;
  assign new_n9004 = new_n8699 ^ new_n8683;
  assign new_n9005 = new_n9004 ^ new_n8865;
  assign new_n9006 = new_n9005 ^ new_n8908;
  assign new_n9007 = new_n9006 ^ new_n8886;
  assign new_n9008 = new_n9007 ^ new_n9003;
  assign new_n9009 = ~new_n8875 & new_n8741;
  assign new_n9010 = new_n9009 ^ new_n8909;
  assign new_n9011 = new_n9010 ^ new_n8871;
  assign new_n9012 = new_n9011 ^ new_n8879;
  assign new_n9013 = new_n8969 ^ new_n8512;
  assign new_n9014 = new_n9013 ^ new_n9012;
  assign new_n9015 = new_n9014 ^ new_n8961;
  assign new_n9016 = new_n8973 ^ new_n8197;
  assign new_n9017 = ~new_n8214 & new_n8120;
  assign new_n9018 = new_n9017 ^ new_n8223;
  assign new_n9019 = new_n9018 ^ new_n9016;
  assign new_n9020 = new_n8979 ^ new_n8340;
  assign new_n9021 = ~new_n8315 & new_n8243;
  assign new_n9022 = new_n9021 ^ new_n8327;
  assign new_n9023 = new_n9022 ^ new_n9020;
  assign new_n9024 = new_n9023 ^ n43;
  assign new_n9025 = new_n9024 ^ n11;
  assign new_n9026 = new_n9025 ^ new_n9019;
  assign new_n9027 = new_n8988 ^ new_n8673;
  assign new_n9028 = ~new_n8691 & new_n8597;
  assign new_n9029 = new_n9028 ^ new_n8700;
  assign new_n9030 = new_n9029 ^ new_n9027;
  assign new_n9031 = new_n9030 ^ new_n9026;
  assign new_n9032 = new_n9031 ^ new_n9015;
  assign new_n9033 = new_n9032 ^ new_n8995;
  assign new_n9034 = new_n9033 ^ new_n9008;
  assign new_n9035 = ~new_n8918 & ~new_n9034;
  assign new_n9036 = new_n9035 ^ new_n8918;
  assign new_n9037 = new_n9032 ^ new_n8957;
  assign new_n9038 = new_n8869 ^ new_n8833;
  assign new_n9039 = new_n9011 ^ new_n8877;
  assign new_n9040 = new_n9039 ^ new_n9038;
  assign new_n9041 = new_n9040 ^ new_n8971;
  assign new_n9042 = new_n8979 ^ new_n8925;
  assign new_n9043 = new_n9042 ^ new_n8349;
  assign new_n9044 = new_n9043 ^ n41;
  assign new_n9045 = new_n9044 ^ n9;
  assign new_n9046 = new_n9045 ^ new_n9041;
  assign new_n9047 = new_n8973 ^ new_n8919;
  assign new_n9048 = new_n9047 ^ new_n8208;
  assign new_n9049 = new_n8988 ^ new_n8942;
  assign new_n9050 = new_n9049 ^ new_n8685;
  assign new_n9051 = new_n9050 ^ new_n9048;
  assign new_n9052 = new_n9051 ^ new_n8885;
  assign new_n9053 = new_n9052 ^ new_n9046;
  assign new_n9054 = new_n9053 ^ new_n8918;
  assign new_n9055 = new_n9037 & new_n9054;
  assign new_n9056 = new_n9055 ^ new_n9036;
  assign new_n9057 = new_n9053 ^ new_n8859;
  assign new_n9058 = new_n9057 ^ new_n9056;
  assign new_n9059 = new_n8871 ^ new_n8838;
  assign new_n9060 = new_n9009 ^ new_n8911;
  assign new_n9061 = new_n9060 ^ new_n8878;
  assign new_n9062 = new_n9061 ^ new_n9059;
  assign new_n9063 = new_n9062 ^ new_n8952;
  assign new_n9064 = new_n8982 ^ new_n8348;
  assign new_n9065 = new_n9064 ^ n44;
  assign new_n9066 = new_n9065 ^ n12;
  assign new_n9067 = new_n9066 ^ new_n9063;
  assign new_n9068 = new_n9067 ^ new_n8886;
  assign new_n9069 = new_n8991 ^ new_n8684;
  assign new_n9070 = new_n9069 ^ new_n9013;
  assign new_n9071 = new_n8976 ^ new_n8207;
  assign new_n9072 = new_n9071 ^ new_n9070;
  assign new_n9073 = new_n9072 ^ new_n9068;
  assign new_n9074 = new_n9073 ^ new_n9053;
  assign new_n9075 = new_n8996 & new_n9074;
  assign new_n9076 = new_n9073 ^ new_n9032;
  assign new_n9077 = new_n9076 ^ new_n9057;
  assign new_n9078 = new_n9073 ^ new_n8859;
  assign new_n9079 = new_n9077 & new_n9078;
  assign new_n9080 = new_n9079 ^ new_n9075;
  assign new_n9081 = new_n9032 ^ new_n8955;
  assign new_n9082 = new_n9081 ^ new_n9080;
  assign new_n9083 = new_n9082 ^ new_n9058;
  assign new_n9084 = new_n9074 ^ new_n8956;
  assign new_n9085 = new_n9073 ^ new_n8918;
  assign new_n9086 = new_n9085 ^ new_n9057;
  assign new_n9087 = new_n9084 & new_n9086;
  assign new_n9088 = new_n9087 ^ new_n8995;
  assign new_n9089 = new_n9088 ^ new_n9084;
  assign new_n9090 = new_n9084 ^ new_n9008;
  assign new_n9091 = new_n9034 ^ new_n8918;
  assign new_n9092 = new_n9091 ^ new_n9057;
  assign new_n9093 = new_n9090 & new_n9092;
  assign new_n9094 = new_n9093 ^ new_n9080;
  assign new_n9095 = new_n9094 ^ new_n8859;
  assign new_n9096 = new_n9095 ^ new_n9089;
  assign new_n9097 = ~new_n9083 & new_n9096;
  assign new_n9098 = new_n9073 ^ new_n9034;
  assign new_n9099 = new_n9008 & new_n9098;
  assign new_n9100 = new_n9099 ^ new_n9073;
  assign new_n9101 = new_n9100 ^ new_n9088;
  assign new_n9102 = new_n9101 ^ new_n9097;
  assign new_n9103 = new_n9084 ^ new_n9033;
  assign new_n9104 = new_n9057 & new_n9103;
  assign new_n9105 = new_n9104 ^ new_n9075;
  assign new_n9106 = new_n9105 ^ new_n9037;
  assign new_n9107 = new_n9106 ^ new_n9102;
  assign new_n9108 = new_n9053 ^ new_n9034;
  assign new_n9109 = new_n9008 ^ new_n8996;
  assign new_n9110 = new_n9108 & new_n9109;
  assign new_n9111 = new_n9110 ^ new_n9035;
  assign new_n9112 = new_n9104 ^ new_n9079;
  assign new_n9113 = new_n9112 ^ new_n9111;
  assign new_n9114 = ~new_n9113 & new_n9107;
  assign new_n9115 = new_n9053 ^ new_n9032;
  assign new_n9116 = new_n9099 ^ new_n9093;
  assign new_n9117 = new_n9116 ^ new_n9112;
  assign new_n9118 = new_n9117 ^ new_n9115;
  assign new_n9119 = new_n9110 ^ new_n9055;
  assign new_n9120 = new_n9119 ^ new_n9053;
  assign new_n9121 = new_n9120 ^ new_n9106;
  assign new_n9122 = new_n9121 ^ new_n9097;
  assign new_n9123 = new_n9118 & new_n9122;
  assign new_n9124 = new_n9123 ^ new_n9114;
  assign new_n9125 = new_n9120 ^ new_n9101;
  assign new_n9126 = new_n9125 ^ new_n9124;
  assign new_n9127 = new_n8996 & new_n9126;
  assign new_n9128 = new_n9074 & new_n9126;
  assign new_n9129 = new_n9128 ^ new_n9127;
  assign new_n9130 = new_n9114 ^ new_n9053;
  assign new_n9131 = new_n9110 ^ new_n9099;
  assign new_n9132 = new_n9032 ^ new_n8918;
  assign new_n9133 = new_n9093 ^ new_n9036;
  assign new_n9134 = new_n9114 ^ new_n9097;
  assign new_n9135 = ~new_n9134 & new_n9121;
  assign new_n9136 = new_n9135 ^ new_n9121;
  assign new_n9137 = new_n9123 ^ new_n9101;
  assign new_n9138 = new_n9137 ^ new_n9106;
  assign new_n9139 = new_n9135 ^ new_n9097;
  assign new_n9140 = new_n9138 & new_n9139;
  assign new_n9141 = new_n9140 ^ new_n9136;
  assign new_n9142 = new_n9141 ^ new_n9133;
  assign new_n9143 = new_n9142 ^ new_n9132;
  assign new_n9144 = new_n9143 ^ new_n9131;
  assign new_n9145 = new_n9144 ^ new_n9130;
  assign new_n9146 = ~new_n9145 & new_n9057;
  assign new_n9147 = new_n9108 & new_n9138;
  assign new_n9148 = ~new_n9145 & new_n9103;
  assign new_n9149 = new_n9148 ^ new_n9147;
  assign new_n9150 = new_n9136 ^ new_n9083;
  assign new_n9151 = ~new_n9150 & new_n9084;
  assign new_n9152 = new_n9121 ^ new_n9114;
  assign new_n9153 = new_n9008 & new_n9152;
  assign new_n9154 = new_n9153 ^ new_n9151;
  assign new_n9155 = new_n9140 ^ new_n9123;
  assign new_n9156 = new_n9155 ^ new_n9096;
  assign new_n9157 = new_n9054 & new_n9156;
  assign new_n9158 = new_n9157 ^ new_n9154;
  assign new_n9159 = new_n9158 ^ new_n9149;
  assign new_n9160 = new_n9159 ^ new_n9146;
  assign new_n9161 = new_n9160 ^ new_n9129;
  assign new_n9162 = new_n9161 ^ new_n8060;
  assign new_n9163 = new_n8112 ^ n54;
  assign new_n9164 = new_n9163 ^ new_n4769;
  assign new_n9165 = new_n8391 ^ new_n4746;
  assign new_n9166 = new_n9165 ^ new_n9164;
  assign new_n9167 = new_n8374 ^ new_n4696;
  assign new_n9168 = new_n8089 ^ n55;
  assign new_n9169 = new_n9168 ^ new_n4762;
  assign new_n9170 = new_n9169 ^ new_n8408;
  assign new_n9171 = new_n9170 ^ new_n9167;
  assign new_n9172 = new_n8106 ^ n53;
  assign new_n9173 = new_n9172 ^ new_n4535;
  assign new_n9174 = new_n9173 ^ new_n8408;
  assign new_n9175 = new_n8418 ^ new_n4786;
  assign new_n9176 = new_n9175 ^ new_n9174;
  assign new_n9177 = new_n9176 ^ new_n9171;
  assign new_n9178 = new_n9177 ^ new_n9166;
  assign new_n9179 = new_n8076 ^ n50;
  assign new_n9180 = new_n9179 ^ new_n4736;
  assign new_n9181 = new_n8362 ^ new_n4627;
  assign new_n9182 = new_n9181 ^ new_n9180;
  assign new_n9183 = new_n9182 ^ new_n9178;
  assign new_n9184 = new_n8081 ^ n56;
  assign new_n9185 = new_n9184 ^ new_n4709;
  assign new_n9186 = new_n8408 ^ new_n4683;
  assign new_n9187 = new_n9186 ^ new_n9185;
  assign new_n9188 = new_n9187 ^ new_n9183;
  assign new_n9189 = new_n8404 ^ new_n2930;
  assign new_n9190 = new_n8062 ^ n52;
  assign new_n9191 = new_n9190 ^ new_n4594;
  assign new_n9192 = new_n9191 ^ new_n8408;
  assign new_n9193 = new_n9192 ^ new_n9189;
  assign new_n9194 = new_n8098 ^ n49;
  assign new_n9195 = new_n9194 ^ new_n3755;
  assign new_n9196 = new_n8355 ^ new_n4725;
  assign new_n9197 = new_n9196 ^ new_n9195;
  assign new_n9198 = new_n9197 ^ new_n9193;
  assign new_n9199 = new_n9198 ^ new_n9177;
  assign new_n9200 = new_n9193 ^ new_n9171;
  assign new_n9201 = new_n9197 ^ new_n9166;
  assign new_n9202 = new_n9201 ^ new_n9200;
  assign new_n9203 = ~new_n9199 & ~new_n9202;
  assign new_n9204 = new_n9203 ^ new_n9182;
  assign new_n9205 = new_n9204 ^ new_n9199;
  assign new_n9206 = new_n9199 ^ new_n9187;
  assign new_n9207 = new_n8072 ^ n51;
  assign new_n9208 = new_n9207 ^ new_n4649;
  assign new_n9209 = new_n8381 ^ new_n4574;
  assign new_n9210 = new_n9209 ^ new_n9208;
  assign new_n9211 = new_n9210 ^ new_n9182;
  assign new_n9212 = new_n9211 ^ new_n9187;
  assign new_n9213 = new_n9212 ^ new_n9171;
  assign new_n9214 = new_n9213 ^ new_n9201;
  assign new_n9215 = new_n9206 & new_n9214;
  assign new_n9216 = new_n9183 & new_n9198;
  assign new_n9217 = new_n9216 ^ new_n9215;
  assign new_n9218 = new_n9210 ^ new_n9193;
  assign new_n9219 = new_n9218 ^ new_n9201;
  assign new_n9220 = new_n9193 ^ new_n9166;
  assign new_n9221 = ~new_n9219 & new_n9220;
  assign new_n9222 = new_n9221 ^ new_n9166;
  assign new_n9223 = new_n9222 ^ new_n9217;
  assign new_n9224 = new_n9223 ^ new_n9205;
  assign new_n9225 = new_n9171 & new_n9212;
  assign new_n9226 = new_n9225 ^ new_n9171;
  assign new_n9227 = new_n9210 ^ new_n9178;
  assign new_n9228 = new_n9197 ^ new_n9171;
  assign new_n9229 = ~new_n9228 & new_n9227;
  assign new_n9230 = new_n9229 ^ new_n9226;
  assign new_n9231 = new_n9230 ^ new_n9201;
  assign new_n9232 = new_n9221 ^ new_n9216;
  assign new_n9233 = new_n9210 ^ new_n9176;
  assign new_n9234 = new_n9233 ^ new_n9232;
  assign new_n9235 = new_n9234 ^ new_n9231;
  assign new_n9236 = ~new_n9235 & new_n9224;
  assign new_n9237 = new_n9211 ^ new_n9199;
  assign new_n9238 = ~new_n9237 & new_n9201;
  assign new_n9239 = new_n9238 ^ new_n9216;
  assign new_n9240 = new_n9239 ^ new_n9227;
  assign new_n9241 = new_n9212 ^ new_n9197;
  assign new_n9242 = ~new_n9188 & ~new_n9241;
  assign new_n9243 = new_n9242 ^ new_n9229;
  assign new_n9244 = new_n9243 ^ new_n9197;
  assign new_n9245 = new_n9244 ^ new_n9240;
  assign new_n9246 = new_n9245 ^ new_n9236;
  assign new_n9247 = new_n9210 ^ new_n9197;
  assign new_n9248 = new_n9212 ^ new_n9193;
  assign new_n9249 = ~new_n9187 & ~new_n9248;
  assign new_n9250 = new_n9249 ^ new_n9215;
  assign new_n9251 = new_n9238 ^ new_n9221;
  assign new_n9252 = new_n9251 ^ new_n9250;
  assign new_n9253 = new_n9252 ^ new_n9247;
  assign new_n9254 = ~new_n9253 & new_n9246;
  assign new_n9255 = new_n9249 ^ new_n9193;
  assign new_n9256 = new_n9255 ^ new_n9204;
  assign new_n9257 = new_n9256 ^ new_n9254;
  assign new_n9258 = new_n9257 ^ new_n9240;
  assign new_n9259 = ~new_n9188 & ~new_n9258;
  assign new_n9260 = new_n9256 ^ new_n9236;
  assign new_n9261 = new_n9260 ^ new_n9240;
  assign new_n9262 = new_n9242 ^ new_n9225;
  assign new_n9263 = new_n9262 ^ new_n9251;
  assign new_n9264 = ~new_n9261 & ~new_n9263;
  assign new_n9265 = new_n9264 ^ new_n9236;
  assign new_n9266 = ~new_n9245 & ~new_n9265;
  assign new_n9267 = new_n9266 ^ new_n9264;
  assign new_n9268 = new_n9267 ^ new_n9246;
  assign new_n9269 = new_n9268 ^ new_n9235;
  assign new_n9270 = ~new_n9202 & new_n9269;
  assign new_n9271 = new_n9270 ^ new_n9259;
  assign new_n9272 = new_n9264 ^ new_n9245;
  assign new_n9273 = ~new_n9187 & new_n9272;
  assign new_n9274 = new_n9268 ^ new_n9264;
  assign new_n9275 = new_n9274 ^ new_n9263;
  assign new_n9276 = new_n9206 & new_n9275;
  assign new_n9277 = new_n9276 ^ new_n9273;
  assign new_n9278 = new_n9214 & new_n9275;
  assign new_n9279 = new_n9210 ^ new_n9171;
  assign new_n9280 = new_n9226 ^ new_n9215;
  assign new_n9281 = ~new_n9258 & ~new_n9267;
  assign new_n9282 = new_n9281 ^ new_n9268;
  assign new_n9283 = new_n9282 ^ new_n9280;
  assign new_n9284 = new_n9283 ^ new_n9279;
  assign new_n9285 = new_n9284 ^ new_n9193;
  assign new_n9286 = new_n9254 ^ new_n9229;
  assign new_n9287 = new_n9286 ^ new_n9204;
  assign new_n9288 = new_n9287 ^ new_n9285;
  assign new_n9289 = new_n9220 & new_n9288;
  assign new_n9290 = new_n9264 ^ new_n9254;
  assign new_n9291 = new_n9256 ^ new_n9244;
  assign new_n9292 = new_n9291 ^ new_n9290;
  assign new_n9293 = ~new_n9292 & new_n9198;
  assign new_n9294 = new_n9293 ^ new_n9289;
  assign new_n9295 = new_n9294 ^ new_n9278;
  assign new_n9296 = new_n9281 ^ new_n9253;
  assign new_n9297 = ~new_n9212 & ~new_n9296;
  assign new_n9298 = new_n9297 ^ new_n9295;
  assign new_n9299 = new_n9298 ^ new_n9277;
  assign new_n9300 = new_n9299 ^ new_n9271;
  assign new_n9301 = ~new_n9248 & new_n9272;
  assign new_n9302 = ~new_n9219 & new_n9288;
  assign new_n9303 = new_n9281 ^ new_n9254;
  assign new_n9304 = new_n9303 ^ new_n9224;
  assign new_n9305 = new_n9227 & new_n9304;
  assign new_n9306 = new_n9305 ^ new_n9298;
  assign new_n9307 = new_n9306 ^ new_n9302;
  assign new_n9308 = new_n9307 ^ new_n9301;
  assign new_n9309 = ~new_n9241 & ~new_n9258;
  assign new_n9310 = new_n9264 ^ new_n9197;
  assign new_n9311 = new_n9249 ^ new_n9242;
  assign new_n9312 = new_n9311 ^ new_n9284;
  assign new_n9313 = new_n9312 ^ new_n9310;
  assign new_n9314 = ~new_n9237 & ~new_n9313;
  assign new_n9315 = new_n9314 ^ new_n9309;
  assign new_n9316 = ~new_n9199 & new_n9269;
  assign new_n9317 = new_n9316 ^ new_n9273;
  assign new_n9318 = ~new_n9228 & new_n9304;
  assign new_n9319 = new_n9318 ^ new_n9317;
  assign new_n9320 = new_n9319 ^ new_n9315;
  assign new_n9321 = new_n9320 ^ new_n9308;
  assign new_n9322 = new_n9321 ^ new_n9300;
  assign new_n9323 = new_n6477 ^ new_n6073;
  assign new_n9324 = new_n9323 ^ n91;
  assign new_n9325 = new_n6530 ^ new_n4613;
  assign new_n9326 = new_n9325 ^ new_n8743;
  assign new_n9327 = new_n9326 ^ new_n9324;
  assign new_n9328 = new_n8546 ^ new_n6580;
  assign new_n9329 = new_n6546 ^ new_n6530;
  assign new_n9330 = new_n9329 ^ new_n8710;
  assign new_n9331 = new_n9330 ^ new_n9328;
  assign new_n9332 = new_n9331 ^ new_n9327;
  assign new_n9333 = new_n8552 ^ new_n6610;
  assign new_n9334 = new_n8712 ^ new_n8705;
  assign new_n9335 = new_n9334 ^ new_n9333;
  assign new_n9336 = new_n9335 ^ new_n9332;
  assign new_n9337 = new_n8717 ^ new_n1295;
  assign new_n9338 = new_n9337 ^ new_n8712;
  assign new_n9339 = new_n6696 ^ new_n6073;
  assign new_n9340 = new_n6485 ^ n92;
  assign new_n9341 = new_n9340 ^ new_n9339;
  assign new_n9342 = new_n9341 ^ new_n9338;
  assign new_n9343 = new_n9342 ^ new_n9336;
  assign new_n9344 = new_n9335 & new_n9343;
  assign new_n9345 = new_n9344 ^ new_n9342;
  assign new_n9346 = new_n6580 ^ new_n6570;
  assign new_n9347 = new_n9346 ^ new_n8703;
  assign new_n9348 = new_n8571 ^ new_n6670;
  assign new_n9349 = new_n9348 ^ new_n9347;
  assign new_n9350 = new_n9349 ^ new_n9342;
  assign new_n9351 = new_n8751 ^ new_n6623;
  assign new_n9352 = new_n9351 ^ new_n8712;
  assign new_n9353 = new_n6642 ^ new_n6610;
  assign new_n9354 = new_n9353 ^ new_n8563;
  assign new_n9355 = new_n9354 ^ new_n9352;
  assign new_n9356 = new_n6715 ^ new_n6696;
  assign new_n9357 = new_n6690 ^ n93;
  assign new_n9358 = new_n9357 ^ new_n9356;
  assign new_n9359 = new_n8734 ^ new_n4774;
  assign new_n9360 = new_n9359 ^ new_n8712;
  assign new_n9361 = new_n9360 ^ new_n9358;
  assign new_n9362 = new_n9361 ^ new_n9355;
  assign new_n9363 = new_n9362 ^ new_n9350;
  assign new_n9364 = new_n8729 ^ new_n8707;
  assign new_n9365 = new_n8588 ^ new_n6715;
  assign new_n9366 = new_n9365 ^ new_n9364;
  assign new_n9367 = new_n9366 ^ new_n9342;
  assign new_n9368 = new_n9355 ^ new_n9349;
  assign new_n9369 = new_n9368 ^ new_n9367;
  assign new_n9370 = ~new_n9363 & ~new_n9369;
  assign new_n9371 = new_n9370 ^ new_n9331;
  assign new_n9372 = new_n9371 ^ new_n9345;
  assign new_n9373 = ~new_n9336 & new_n9355;
  assign new_n9374 = new_n9373 ^ new_n9355;
  assign new_n9375 = new_n9366 ^ new_n9362;
  assign new_n9376 = new_n9375 ^ new_n9327;
  assign new_n9377 = ~new_n9368 & ~new_n9376;
  assign new_n9378 = new_n9377 ^ new_n9374;
  assign new_n9379 = new_n9366 ^ new_n9349;
  assign new_n9380 = new_n9379 ^ new_n9378;
  assign new_n9381 = new_n9342 ^ new_n9327;
  assign new_n9382 = new_n9381 ^ new_n9379;
  assign new_n9383 = new_n9367 & new_n9382;
  assign new_n9384 = new_n9375 ^ new_n9331;
  assign new_n9385 = ~new_n9384 & new_n9350;
  assign new_n9386 = new_n9385 ^ new_n9383;
  assign new_n9387 = new_n9361 ^ new_n9327;
  assign new_n9388 = new_n9387 ^ new_n9386;
  assign new_n9389 = new_n9388 ^ new_n9380;
  assign new_n9390 = new_n9371 ^ new_n9363;
  assign new_n9391 = new_n9363 ^ new_n9335;
  assign new_n9392 = new_n9355 ^ new_n9336;
  assign new_n9393 = new_n9392 ^ new_n9379;
  assign new_n9394 = ~new_n9391 & ~new_n9393;
  assign new_n9395 = new_n9394 ^ new_n9385;
  assign new_n9396 = new_n9383 ^ new_n9366;
  assign new_n9397 = new_n9396 ^ new_n9395;
  assign new_n9398 = new_n9397 ^ new_n9390;
  assign new_n9399 = ~new_n9398 & new_n9389;
  assign new_n9400 = new_n9399 ^ new_n9372;
  assign new_n9401 = new_n9363 ^ new_n9332;
  assign new_n9402 = ~new_n9401 & new_n9379;
  assign new_n9403 = new_n9402 ^ new_n9385;
  assign new_n9404 = new_n9403 ^ new_n9376;
  assign new_n9405 = new_n9404 ^ new_n9400;
  assign new_n9406 = new_n9349 ^ new_n9336;
  assign new_n9407 = new_n9384 ^ new_n9335;
  assign new_n9408 = ~new_n9407 & new_n9406;
  assign new_n9409 = new_n9408 ^ new_n9373;
  assign new_n9410 = new_n9402 ^ new_n9383;
  assign new_n9411 = new_n9410 ^ new_n9409;
  assign new_n9412 = ~new_n9405 & ~new_n9411;
  assign new_n9413 = new_n9408 ^ new_n9377;
  assign new_n9414 = new_n9413 ^ new_n9349;
  assign new_n9415 = new_n9414 ^ new_n9404;
  assign new_n9416 = new_n9415 ^ new_n9412;
  assign new_n9417 = ~new_n9416 & new_n9343;
  assign new_n9418 = new_n9355 ^ new_n9327;
  assign new_n9419 = new_n9394 ^ new_n9374;
  assign new_n9420 = new_n9412 ^ new_n9399;
  assign new_n9421 = ~new_n9420 & new_n9415;
  assign new_n9422 = new_n9421 ^ new_n9412;
  assign new_n9423 = new_n9415 ^ new_n9399;
  assign new_n9424 = new_n9349 ^ new_n9327;
  assign new_n9425 = new_n9394 ^ new_n9344;
  assign new_n9426 = new_n9425 ^ new_n9410;
  assign new_n9427 = new_n9426 ^ new_n9424;
  assign new_n9428 = ~new_n9423 & new_n9427;
  assign new_n9429 = new_n9428 ^ new_n9372;
  assign new_n9430 = new_n9429 ^ new_n9404;
  assign new_n9431 = ~new_n9422 & ~new_n9430;
  assign new_n9432 = new_n9423 ^ new_n9422;
  assign new_n9433 = new_n9432 ^ new_n9431;
  assign new_n9434 = new_n9433 ^ new_n9419;
  assign new_n9435 = new_n9434 ^ new_n9418;
  assign new_n9436 = new_n9435 ^ new_n9342;
  assign new_n9437 = new_n9428 ^ new_n9377;
  assign new_n9438 = new_n9437 ^ new_n9371;
  assign new_n9439 = new_n9438 ^ new_n9436;
  assign new_n9440 = ~new_n9439 & new_n9382;
  assign new_n9441 = new_n9431 ^ new_n9427;
  assign new_n9442 = new_n9336 & new_n9441;
  assign new_n9443 = ~new_n9439 & new_n9367;
  assign new_n9444 = new_n9428 ^ new_n9412;
  assign new_n9445 = new_n9414 ^ new_n9372;
  assign new_n9446 = new_n9445 ^ new_n9444;
  assign new_n9447 = new_n9350 & new_n9446;
  assign new_n9448 = new_n9447 ^ new_n9443;
  assign new_n9449 = new_n9432 ^ new_n9412;
  assign new_n9450 = new_n9449 ^ new_n9411;
  assign new_n9451 = ~new_n9393 & ~new_n9450;
  assign new_n9452 = new_n9451 ^ new_n9448;
  assign new_n9453 = new_n9452 ^ new_n9442;
  assign new_n9454 = new_n9431 ^ new_n9428;
  assign new_n9455 = new_n9454 ^ new_n9398;
  assign new_n9456 = ~new_n9376 & ~new_n9455;
  assign new_n9457 = new_n9456 ^ new_n9453;
  assign new_n9458 = new_n9457 ^ new_n9440;
  assign new_n9459 = new_n9458 ^ new_n9417;
  assign new_n9460 = new_n9412 ^ new_n9349;
  assign new_n9461 = new_n9408 ^ new_n9344;
  assign new_n9462 = new_n9461 ^ new_n9435;
  assign new_n9463 = new_n9462 ^ new_n9460;
  assign new_n9464 = ~new_n9401 & ~new_n9463;
  assign new_n9465 = ~new_n9430 & new_n9406;
  assign new_n9466 = new_n9465 ^ new_n9464;
  assign new_n9467 = ~new_n9368 & ~new_n9455;
  assign new_n9468 = ~new_n9416 & new_n9335;
  assign new_n9469 = new_n9432 ^ new_n9389;
  assign new_n9470 = ~new_n9363 & new_n9469;
  assign new_n9471 = new_n9470 ^ new_n9468;
  assign new_n9472 = new_n9471 ^ new_n9467;
  assign new_n9473 = new_n9472 ^ new_n9466;
  assign new_n9474 = new_n9473 ^ new_n9459;
  assign new_n9475 = new_n9474 ^ new_n9322;
  assign new_n9476 = new_n7623 ^ new_n7465;
  assign new_n9477 = new_n9476 ^ new_n7523;
  assign new_n9478 = new_n9477 ^ new_n7541;
  assign new_n9479 = new_n9478 ^ new_n7649;
  assign new_n9480 = new_n7575 ^ new_n7541;
  assign new_n9481 = new_n9480 ^ new_n7649;
  assign new_n9482 = new_n7465 & new_n9481;
  assign new_n9483 = new_n9482 ^ new_n7465;
  assign new_n9484 = new_n7465 ^ new_n6844;
  assign new_n9485 = new_n9477 ^ new_n7575;
  assign new_n9486 = ~new_n9484 & new_n9485;
  assign new_n9487 = new_n9486 ^ new_n9483;
  assign new_n9488 = new_n7523 ^ new_n6844;
  assign new_n9489 = new_n9488 ^ new_n9487;
  assign new_n9490 = new_n7594 ^ new_n7575;
  assign new_n9491 = new_n9490 ^ new_n9488;
  assign new_n9492 = new_n7594 ^ new_n7523;
  assign new_n9493 = ~new_n9491 & new_n9492;
  assign new_n9494 = new_n7594 ^ new_n6844;
  assign new_n9495 = new_n9478 & new_n9494;
  assign new_n9496 = new_n9495 ^ new_n9493;
  assign new_n9497 = new_n7623 ^ new_n7575;
  assign new_n9498 = new_n9497 ^ new_n9496;
  assign new_n9499 = new_n9498 ^ new_n9489;
  assign new_n9500 = new_n9494 ^ new_n9476;
  assign new_n9501 = new_n7594 ^ new_n7465;
  assign new_n9502 = new_n9501 ^ new_n9488;
  assign new_n9503 = ~new_n9500 & ~new_n9502;
  assign new_n9504 = new_n9503 ^ new_n7541;
  assign new_n9505 = new_n9504 ^ new_n9500;
  assign new_n9506 = new_n9500 ^ new_n7649;
  assign new_n9507 = new_n9481 ^ new_n7465;
  assign new_n9508 = new_n9507 ^ new_n9488;
  assign new_n9509 = new_n9506 & new_n9508;
  assign new_n9510 = new_n9509 ^ new_n7523;
  assign new_n9511 = new_n9510 ^ new_n9496;
  assign new_n9512 = new_n9511 ^ new_n9505;
  assign new_n9513 = ~new_n9499 & new_n9512;
  assign new_n9514 = new_n9500 ^ new_n9480;
  assign new_n9515 = ~new_n9514 & new_n9488;
  assign new_n9516 = new_n9515 ^ new_n9495;
  assign new_n9517 = new_n9516 ^ new_n9485;
  assign new_n9518 = new_n9481 ^ new_n6844;
  assign new_n9519 = ~new_n9479 & ~new_n9518;
  assign new_n9520 = new_n9519 ^ new_n9486;
  assign new_n9521 = new_n9520 ^ new_n6844;
  assign new_n9522 = new_n9521 ^ new_n9517;
  assign new_n9523 = new_n9522 ^ new_n9513;
  assign new_n9524 = new_n7575 ^ new_n6844;
  assign new_n9525 = ~new_n7649 & ~new_n9480;
  assign new_n9526 = new_n7594 & new_n7649;
  assign new_n9527 = new_n9526 ^ new_n9525;
  assign new_n9528 = new_n9527 ^ new_n7594;
  assign new_n9529 = new_n9528 ^ new_n9509;
  assign new_n9530 = new_n9515 ^ new_n9493;
  assign new_n9531 = new_n9530 ^ new_n9529;
  assign new_n9532 = new_n9531 ^ new_n9524;
  assign new_n9533 = ~new_n9532 & new_n9523;
  assign new_n9534 = new_n9527 ^ new_n9504;
  assign new_n9535 = new_n9534 ^ new_n9533;
  assign new_n9536 = new_n9535 ^ new_n9517;
  assign new_n9537 = ~new_n9479 & ~new_n9536;
  assign new_n9538 = new_n9534 ^ new_n9513;
  assign new_n9539 = new_n9538 ^ new_n9517;
  assign new_n9540 = new_n9519 ^ new_n9482;
  assign new_n9541 = new_n9540 ^ new_n9530;
  assign new_n9542 = ~new_n9539 & ~new_n9541;
  assign new_n9543 = new_n9542 ^ new_n9513;
  assign new_n9544 = ~new_n9522 & ~new_n9543;
  assign new_n9545 = new_n9544 ^ new_n9542;
  assign new_n9546 = new_n9545 ^ new_n9523;
  assign new_n9547 = new_n9546 ^ new_n9499;
  assign new_n9548 = ~new_n9502 & new_n9547;
  assign new_n9549 = new_n9548 ^ new_n9537;
  assign new_n9550 = ~new_n9536 & ~new_n9545;
  assign new_n9551 = new_n9550 ^ new_n9532;
  assign new_n9552 = ~new_n9481 & ~new_n9551;
  assign new_n9553 = new_n9546 ^ new_n9542;
  assign new_n9554 = new_n9553 ^ new_n9541;
  assign new_n9555 = new_n9508 & new_n9554;
  assign new_n9556 = new_n7575 ^ new_n7465;
  assign new_n9557 = new_n9509 ^ new_n9483;
  assign new_n9558 = new_n9550 ^ new_n9546;
  assign new_n9559 = new_n9558 ^ new_n9557;
  assign new_n9560 = new_n9559 ^ new_n9556;
  assign new_n9561 = new_n9560 ^ new_n7594;
  assign new_n9562 = new_n9533 ^ new_n9486;
  assign new_n9563 = new_n9562 ^ new_n9504;
  assign new_n9564 = new_n9563 ^ new_n9561;
  assign new_n9565 = new_n9492 & new_n9564;
  assign new_n9566 = new_n9542 ^ new_n9533;
  assign new_n9567 = new_n9534 ^ new_n9521;
  assign new_n9568 = new_n9567 ^ new_n9566;
  assign new_n9569 = ~new_n9568 & new_n9494;
  assign new_n9570 = new_n9569 ^ new_n9565;
  assign new_n9571 = new_n9570 ^ new_n9555;
  assign new_n9572 = new_n9571 ^ new_n9552;
  assign new_n9573 = new_n9542 ^ new_n9522;
  assign new_n9574 = ~new_n7649 & new_n9573;
  assign new_n9575 = new_n9506 & new_n9554;
  assign new_n9576 = new_n9575 ^ new_n9574;
  assign new_n9577 = new_n9576 ^ new_n9572;
  assign new_n9578 = new_n9577 ^ new_n9549;
  assign new_n9579 = new_n9578 ^ new_n3593;
  assign new_n9580 = new_n5540 ^ new_n5451;
  assign new_n9581 = new_n8357 ^ new_n5037;
  assign new_n9582 = new_n9581 ^ new_n5616;
  assign new_n9583 = new_n9582 ^ new_n9580;
  assign new_n9584 = new_n5680 ^ new_n5662;
  assign new_n9585 = new_n9584 ^ new_n5687;
  assign new_n9586 = new_n8420 ^ new_n8087;
  assign new_n9587 = new_n9586 ^ new_n9585;
  assign new_n9588 = new_n5645 ^ new_n5632;
  assign new_n9589 = new_n9588 ^ new_n5552;
  assign new_n9590 = new_n9589 ^ new_n5621;
  assign new_n9591 = new_n8393 ^ new_n5567;
  assign new_n9592 = new_n9591 ^ new_n5677;
  assign new_n9593 = new_n9592 ^ new_n9590;
  assign new_n9594 = new_n5667 ^ new_n5584;
  assign new_n9595 = new_n9594 ^ new_n5654;
  assign new_n9596 = new_n8401 ^ new_n5621;
  assign new_n9597 = new_n9596 ^ new_n5681;
  assign new_n9598 = new_n9597 ^ new_n9595;
  assign new_n9599 = new_n9598 ^ new_n9593;
  assign new_n9600 = new_n9599 ^ new_n9587;
  assign new_n9601 = new_n9600 ^ new_n9583;
  assign new_n9602 = new_n8370 ^ new_n5552;
  assign new_n9603 = new_n8091 ^ new_n5621;
  assign new_n9604 = new_n9603 ^ new_n9602;
  assign new_n9605 = new_n9604 ^ new_n9601;
  assign new_n9606 = new_n5594 ^ new_n5539;
  assign new_n9607 = new_n8364 ^ new_n5492;
  assign new_n9608 = new_n9607 ^ new_n5173;
  assign new_n9609 = new_n9608 ^ new_n9606;
  assign new_n9610 = new_n8410 ^ new_n5470;
  assign new_n9611 = new_n5620 ^ new_n5612;
  assign new_n9612 = new_n9611 ^ new_n5560;
  assign new_n9613 = new_n9612 ^ new_n9610;
  assign new_n9614 = new_n9613 ^ new_n9609;
  assign new_n9615 = new_n9609 ^ new_n9583;
  assign new_n9616 = ~new_n9604 & ~new_n9615;
  assign new_n9617 = new_n8379 ^ new_n5621;
  assign new_n9618 = new_n9617 ^ new_n5668;
  assign new_n9619 = new_n5601 ^ new_n5593;
  assign new_n9620 = new_n9619 ^ new_n5513;
  assign new_n9621 = new_n9620 ^ new_n9618;
  assign new_n9622 = new_n9604 & new_n9621;
  assign new_n9623 = new_n9622 ^ new_n9616;
  assign new_n9624 = new_n9623 ^ new_n9621;
  assign new_n9625 = new_n9621 ^ new_n9613;
  assign new_n9626 = new_n9625 ^ new_n9599;
  assign new_n9627 = new_n9626 ^ new_n9604;
  assign new_n9628 = new_n9615 ^ new_n9604;
  assign new_n9629 = new_n9628 ^ new_n9593;
  assign new_n9630 = new_n9613 ^ new_n9587;
  assign new_n9631 = new_n9630 ^ new_n9629;
  assign new_n9632 = new_n9627 & new_n9631;
  assign new_n9633 = new_n9632 ^ new_n9624;
  assign new_n9634 = new_n9621 ^ new_n9587;
  assign new_n9635 = new_n9621 ^ new_n9609;
  assign new_n9636 = new_n9635 ^ new_n9630;
  assign new_n9637 = ~new_n9636 & new_n9634;
  assign new_n9638 = new_n9626 ^ new_n9615;
  assign new_n9639 = ~new_n9638 & new_n9630;
  assign new_n9640 = new_n9639 ^ new_n9637;
  assign new_n9641 = new_n9640 ^ new_n9633;
  assign new_n9642 = new_n9641 ^ new_n9614;
  assign new_n9643 = new_n9593 & new_n9628;
  assign new_n9644 = new_n9643 ^ new_n9593;
  assign new_n9645 = new_n9609 ^ new_n9600;
  assign new_n9646 = new_n9613 ^ new_n9593;
  assign new_n9647 = ~new_n9646 & new_n9645;
  assign new_n9648 = new_n9647 ^ new_n9644;
  assign new_n9649 = new_n9648 ^ new_n9630;
  assign new_n9650 = new_n9601 & new_n9625;
  assign new_n9651 = new_n9650 ^ new_n9637;
  assign new_n9652 = new_n9609 ^ new_n9598;
  assign new_n9653 = new_n9652 ^ new_n9651;
  assign new_n9654 = new_n9653 ^ new_n9649;
  assign new_n9655 = new_n9646 ^ new_n9634;
  assign new_n9656 = ~new_n9626 & ~new_n9655;
  assign new_n9657 = new_n9656 ^ new_n9583;
  assign new_n9658 = new_n9657 ^ new_n9626;
  assign new_n9659 = new_n9651 ^ new_n9632;
  assign new_n9660 = new_n9659 ^ new_n9587;
  assign new_n9661 = new_n9660 ^ new_n9658;
  assign new_n9662 = ~new_n9654 & new_n9661;
  assign new_n9663 = new_n9650 ^ new_n9639;
  assign new_n9664 = new_n9663 ^ new_n9645;
  assign new_n9665 = new_n9628 ^ new_n9613;
  assign new_n9666 = ~new_n9605 & ~new_n9665;
  assign new_n9667 = new_n9666 ^ new_n9647;
  assign new_n9668 = new_n9667 ^ new_n9613;
  assign new_n9669 = new_n9668 ^ new_n9664;
  assign new_n9670 = new_n9669 ^ new_n9662;
  assign new_n9671 = ~new_n9642 & new_n9670;
  assign new_n9672 = new_n9657 ^ new_n9623;
  assign new_n9673 = new_n9672 ^ new_n9671;
  assign new_n9674 = new_n9673 ^ new_n9664;
  assign new_n9675 = ~new_n9605 & ~new_n9674;
  assign new_n9676 = new_n9672 ^ new_n9662;
  assign new_n9677 = new_n9676 ^ new_n9664;
  assign new_n9678 = new_n9666 ^ new_n9643;
  assign new_n9679 = new_n9678 ^ new_n9640;
  assign new_n9680 = ~new_n9677 & ~new_n9679;
  assign new_n9681 = new_n9680 ^ new_n9662;
  assign new_n9682 = ~new_n9681 & new_n9669;
  assign new_n9683 = new_n9682 ^ new_n9669;
  assign new_n9684 = new_n9683 ^ new_n9654;
  assign new_n9685 = ~new_n9655 & ~new_n9684;
  assign new_n9686 = new_n9685 ^ new_n9675;
  assign new_n9687 = new_n9680 ^ new_n9669;
  assign new_n9688 = ~new_n9604 & new_n9687;
  assign new_n9689 = new_n9683 ^ new_n9680;
  assign new_n9690 = new_n9689 ^ new_n9679;
  assign new_n9691 = ~new_n9690 & new_n9627;
  assign new_n9692 = new_n9691 ^ new_n9688;
  assign new_n9693 = new_n9682 ^ new_n9662;
  assign new_n9694 = ~new_n9674 & new_n9693;
  assign new_n9695 = new_n9694 ^ new_n9642;
  assign new_n9696 = ~new_n9628 & ~new_n9695;
  assign new_n9697 = ~new_n9690 & new_n9631;
  assign new_n9698 = new_n9609 ^ new_n9593;
  assign new_n9699 = new_n9644 ^ new_n9632;
  assign new_n9700 = new_n9694 ^ new_n9683;
  assign new_n9701 = new_n9700 ^ new_n9699;
  assign new_n9702 = new_n9701 ^ new_n9698;
  assign new_n9703 = new_n9702 ^ new_n9621;
  assign new_n9704 = new_n9671 ^ new_n9647;
  assign new_n9705 = new_n9704 ^ new_n9657;
  assign new_n9706 = new_n9705 ^ new_n9703;
  assign new_n9707 = ~new_n9706 & new_n9634;
  assign new_n9708 = new_n9680 ^ new_n9671;
  assign new_n9709 = new_n9672 ^ new_n9668;
  assign new_n9710 = new_n9709 ^ new_n9708;
  assign new_n9711 = ~new_n9710 & new_n9625;
  assign new_n9712 = new_n9711 ^ new_n9707;
  assign new_n9713 = new_n9712 ^ new_n9697;
  assign new_n9714 = new_n9713 ^ new_n9696;
  assign new_n9715 = new_n9714 ^ new_n9692;
  assign new_n9716 = new_n9715 ^ new_n9686;
  assign new_n9717 = new_n7417 ^ new_n576;
  assign new_n9718 = new_n7655 ^ new_n7400;
  assign new_n9719 = new_n9718 ^ new_n9717;
  assign new_n9720 = new_n7588 ^ new_n7566;
  assign new_n9721 = new_n7252 ^ new_n567;
  assign new_n9722 = new_n9721 ^ new_n7547;
  assign new_n9723 = new_n9722 ^ new_n9720;
  assign new_n9724 = new_n7602 ^ new_n598;
  assign new_n9725 = new_n9724 ^ new_n8586;
  assign new_n9726 = new_n7633 ^ new_n7400;
  assign new_n9727 = new_n9726 ^ new_n9725;
  assign new_n9728 = new_n7454 ^ new_n7400;
  assign new_n9729 = new_n7521 ^ new_n592;
  assign new_n9730 = new_n9729 ^ new_n8555;
  assign new_n9731 = new_n9730 ^ new_n9728;
  assign new_n9732 = new_n9731 ^ new_n9727;
  assign new_n9733 = new_n7616 ^ new_n606;
  assign new_n9734 = new_n8561 ^ new_n7512;
  assign new_n9735 = new_n9734 ^ new_n9733;
  assign new_n9736 = new_n9735 ^ new_n9732;
  assign new_n9737 = new_n9736 ^ new_n9723;
  assign new_n9738 = new_n9737 ^ new_n9719;
  assign new_n9739 = new_n7597 ^ new_n7587;
  assign new_n9740 = new_n7555 ^ new_n561;
  assign new_n9741 = new_n9740 ^ new_n7579;
  assign new_n9742 = new_n9741 ^ new_n9739;
  assign new_n9743 = new_n9742 ^ new_n9723;
  assign new_n9744 = new_n9743 ^ new_n9719;
  assign new_n9745 = ~new_n9731 & ~new_n9744;
  assign new_n9746 = new_n9745 ^ new_n9731;
  assign new_n9747 = new_n7567 ^ new_n585;
  assign new_n9748 = new_n7389 ^ new_n6981;
  assign new_n9749 = new_n9748 ^ new_n7423;
  assign new_n9750 = new_n9749 ^ new_n9747;
  assign new_n9751 = new_n9750 ^ new_n9731;
  assign new_n9752 = new_n9742 ^ new_n9736;
  assign new_n9753 = new_n9751 & new_n9752;
  assign new_n9754 = new_n9753 ^ new_n9746;
  assign new_n9755 = new_n9750 ^ new_n9735;
  assign new_n9756 = new_n9755 ^ new_n9754;
  assign new_n9757 = new_n8579 ^ new_n541;
  assign new_n9758 = new_n9757 ^ new_n7400;
  assign new_n9759 = new_n7608 ^ new_n7596;
  assign new_n9760 = new_n9759 ^ new_n7581;
  assign new_n9761 = new_n9760 ^ new_n9758;
  assign new_n9762 = new_n9761 ^ new_n9742;
  assign new_n9763 = new_n9762 ^ new_n9755;
  assign new_n9764 = new_n9761 ^ new_n9735;
  assign new_n9765 = new_n9763 & new_n9764;
  assign new_n9766 = new_n9761 ^ new_n9750;
  assign new_n9767 = new_n9737 & new_n9766;
  assign new_n9768 = new_n9767 ^ new_n9765;
  assign new_n9769 = new_n9742 ^ new_n9727;
  assign new_n9770 = new_n9769 ^ new_n9768;
  assign new_n9771 = new_n9770 ^ new_n9756;
  assign new_n9772 = new_n9766 ^ new_n9732;
  assign new_n9773 = new_n9761 ^ new_n9731;
  assign new_n9774 = new_n9773 ^ new_n9755;
  assign new_n9775 = new_n9772 & new_n9774;
  assign new_n9776 = new_n9775 ^ new_n9723;
  assign new_n9777 = new_n9776 ^ new_n9772;
  assign new_n9778 = new_n9772 ^ new_n9719;
  assign new_n9779 = new_n9744 ^ new_n9731;
  assign new_n9780 = new_n9779 ^ new_n9755;
  assign new_n9781 = new_n9778 & new_n9780;
  assign new_n9782 = new_n9781 ^ new_n9768;
  assign new_n9783 = new_n9782 ^ new_n9735;
  assign new_n9784 = new_n9783 ^ new_n9777;
  assign new_n9785 = ~new_n9771 & new_n9784;
  assign new_n9786 = new_n9772 ^ new_n9743;
  assign new_n9787 = new_n9755 & new_n9786;
  assign new_n9788 = new_n9787 ^ new_n9767;
  assign new_n9789 = new_n9788 ^ new_n9752;
  assign new_n9790 = new_n9750 ^ new_n9744;
  assign new_n9791 = new_n9738 & new_n9790;
  assign new_n9792 = new_n9791 ^ new_n9753;
  assign new_n9793 = new_n9792 ^ new_n9750;
  assign new_n9794 = new_n9793 ^ new_n9789;
  assign new_n9795 = new_n9794 ^ new_n9785;
  assign new_n9796 = new_n9750 ^ new_n9742;
  assign new_n9797 = new_n9787 ^ new_n9765;
  assign new_n9798 = ~new_n9743 & new_n9719;
  assign new_n9799 = ~new_n9719 & new_n9761;
  assign new_n9800 = new_n9799 ^ new_n9798;
  assign new_n9801 = new_n9800 ^ new_n9761;
  assign new_n9802 = new_n9801 ^ new_n9781;
  assign new_n9803 = new_n9802 ^ new_n9797;
  assign new_n9804 = new_n9803 ^ new_n9796;
  assign new_n9805 = new_n9795 & new_n9804;
  assign new_n9806 = new_n9800 ^ new_n9776;
  assign new_n9807 = new_n9806 ^ new_n9805;
  assign new_n9808 = new_n9807 ^ new_n9789;
  assign new_n9809 = new_n9738 & new_n9808;
  assign new_n9810 = new_n9806 ^ new_n9785;
  assign new_n9811 = new_n9810 ^ new_n9789;
  assign new_n9812 = new_n9791 ^ new_n9745;
  assign new_n9813 = new_n9812 ^ new_n9797;
  assign new_n9814 = ~new_n9813 & new_n9811;
  assign new_n9815 = new_n9814 ^ new_n9785;
  assign new_n9816 = ~new_n9794 & ~new_n9815;
  assign new_n9817 = new_n9816 ^ new_n9814;
  assign new_n9818 = new_n9817 ^ new_n9795;
  assign new_n9819 = new_n9818 ^ new_n9771;
  assign new_n9820 = new_n9774 & new_n9819;
  assign new_n9821 = new_n9820 ^ new_n9809;
  assign new_n9822 = new_n9814 ^ new_n9794;
  assign new_n9823 = new_n9719 & new_n9822;
  assign new_n9824 = new_n9818 ^ new_n9814;
  assign new_n9825 = new_n9824 ^ new_n9813;
  assign new_n9826 = new_n9778 & new_n9825;
  assign new_n9827 = new_n9826 ^ new_n9823;
  assign new_n9828 = ~new_n9817 & new_n9808;
  assign new_n9829 = new_n9828 ^ new_n9804;
  assign new_n9830 = new_n9744 & new_n9829;
  assign new_n9831 = new_n9780 & new_n9825;
  assign new_n9832 = new_n9742 ^ new_n9731;
  assign new_n9833 = new_n9781 ^ new_n9746;
  assign new_n9834 = new_n9828 ^ new_n9818;
  assign new_n9835 = new_n9834 ^ new_n9833;
  assign new_n9836 = new_n9835 ^ new_n9832;
  assign new_n9837 = new_n9836 ^ new_n9761;
  assign new_n9838 = new_n9805 ^ new_n9753;
  assign new_n9839 = new_n9838 ^ new_n9776;
  assign new_n9840 = new_n9839 ^ new_n9837;
  assign new_n9841 = new_n9764 & new_n9840;
  assign new_n9842 = new_n9814 ^ new_n9805;
  assign new_n9843 = new_n9806 ^ new_n9793;
  assign new_n9844 = new_n9843 ^ new_n9842;
  assign new_n9845 = new_n9766 & new_n9844;
  assign new_n9846 = new_n9845 ^ new_n9841;
  assign new_n9847 = new_n9846 ^ new_n9831;
  assign new_n9848 = new_n9847 ^ new_n9830;
  assign new_n9849 = new_n9848 ^ new_n9827;
  assign new_n9850 = new_n9849 ^ new_n9821;
  assign new_n9851 = new_n9850 ^ new_n9716;
  assign new_n9852 = new_n9851 ^ new_n9579;
  assign new_n9853 = ~new_n9292 & new_n9183;
  assign new_n9854 = new_n9853 ^ new_n9270;
  assign new_n9855 = new_n9854 ^ new_n9307;
  assign new_n9856 = ~new_n9384 & new_n9446;
  assign new_n9857 = ~new_n9369 & new_n9469;
  assign new_n9858 = new_n9857 ^ new_n9856;
  assign new_n9859 = new_n9858 ^ new_n9458;
  assign new_n9860 = new_n9859 ^ new_n9855;
  assign new_n9861 = new_n9860 ^ new_n9852;
  assign new_n9862 = new_n9861 ^ new_n9475;
  assign new_n9863 = new_n9472 ^ new_n9456;
  assign new_n9864 = ~new_n9392 & new_n9441;
  assign new_n9865 = ~new_n9407 & ~new_n9430;
  assign new_n9866 = new_n9865 ^ new_n9864;
  assign new_n9867 = new_n9866 ^ new_n9448;
  assign new_n9868 = new_n9867 ^ new_n9863;
  assign new_n9869 = new_n9680 ^ new_n9613;
  assign new_n9870 = new_n9666 ^ new_n9624;
  assign new_n9871 = new_n9870 ^ new_n9702;
  assign new_n9872 = new_n9871 ^ new_n9869;
  assign new_n9873 = ~new_n9638 & new_n9872;
  assign new_n9874 = new_n9694 ^ new_n9671;
  assign new_n9875 = new_n9874 ^ new_n9661;
  assign new_n9876 = ~new_n9646 & new_n9875;
  assign new_n9877 = new_n9876 ^ new_n9873;
  assign new_n9878 = ~new_n9636 & ~new_n9706;
  assign new_n9879 = new_n9878 ^ new_n9696;
  assign new_n9880 = ~new_n9695 & new_n9629;
  assign new_n9881 = new_n9880 ^ new_n9675;
  assign new_n9882 = new_n9881 ^ new_n9712;
  assign new_n9883 = new_n9882 ^ new_n9879;
  assign new_n9884 = new_n9883 ^ new_n9877;
  assign new_n9885 = new_n9814 ^ new_n9750;
  assign new_n9886 = new_n9801 ^ new_n9791;
  assign new_n9887 = new_n9886 ^ new_n9836;
  assign new_n9888 = new_n9887 ^ new_n9885;
  assign new_n9889 = new_n9786 & new_n9888;
  assign new_n9890 = new_n9828 ^ new_n9805;
  assign new_n9891 = new_n9890 ^ new_n9784;
  assign new_n9892 = new_n9751 & new_n9891;
  assign new_n9893 = new_n9892 ^ new_n9889;
  assign new_n9894 = new_n9763 & new_n9840;
  assign new_n9895 = new_n9894 ^ new_n9830;
  assign new_n9896 = new_n9779 & new_n9829;
  assign new_n9897 = new_n9896 ^ new_n9809;
  assign new_n9898 = new_n9897 ^ new_n9846;
  assign new_n9899 = new_n9898 ^ new_n9895;
  assign new_n9900 = new_n9899 ^ new_n9893;
  assign new_n9901 = new_n9900 ^ new_n9884;
  assign new_n9902 = new_n9901 ^ new_n9868;
  assign new_n9903 = new_n9902 ^ new_n9860;
  assign new_n9904 = new_n9542 ^ new_n6844;
  assign new_n9905 = new_n9528 ^ new_n9519;
  assign new_n9906 = new_n9905 ^ new_n9560;
  assign new_n9907 = new_n9906 ^ new_n9904;
  assign new_n9908 = ~new_n9514 & ~new_n9907;
  assign new_n9909 = new_n9550 ^ new_n9533;
  assign new_n9910 = new_n9909 ^ new_n9512;
  assign new_n9911 = ~new_n9484 & new_n9910;
  assign new_n9912 = new_n9911 ^ new_n9908;
  assign new_n9913 = ~new_n9491 & new_n9564;
  assign new_n9914 = new_n9913 ^ new_n9552;
  assign new_n9915 = ~new_n9551 & new_n9507;
  assign new_n9916 = new_n9915 ^ new_n9537;
  assign new_n9917 = new_n9916 ^ new_n9570;
  assign new_n9918 = new_n9917 ^ new_n9914;
  assign new_n9919 = new_n9918 ^ new_n9912;
  assign new_n9920 = new_n9919 ^ new_n3420;
  assign new_n9921 = new_n9318 ^ new_n9314;
  assign new_n9922 = new_n9302 ^ new_n9297;
  assign new_n9923 = ~new_n9296 & new_n9213;
  assign new_n9924 = new_n9923 ^ new_n9259;
  assign new_n9925 = new_n9924 ^ new_n9294;
  assign new_n9926 = new_n9925 ^ new_n9922;
  assign new_n9927 = new_n9926 ^ new_n9921;
  assign new_n9928 = new_n9927 ^ new_n9920;
  assign new_n9929 = new_n9319 ^ new_n9305;
  assign new_n9930 = new_n9929 ^ new_n9925;
  assign new_n9931 = new_n9930 ^ new_n9928;
  assign new_n9932 = new_n9931 ^ new_n9903;
  assign new_n9933 = new_n9932 ^ new_n9862;
  assign new_n9934 = new_n9761 ^ new_n9744;
  assign new_n9935 = new_n9822 & new_n9934;
  assign new_n9936 = new_n9752 & new_n9891;
  assign new_n9937 = new_n9936 ^ new_n9848;
  assign new_n9938 = new_n9937 ^ new_n9894;
  assign new_n9939 = new_n9938 ^ new_n9935;
  assign new_n9940 = new_n9790 & new_n9808;
  assign new_n9941 = new_n9940 ^ new_n9889;
  assign new_n9942 = new_n9772 & new_n9819;
  assign new_n9943 = new_n9942 ^ new_n9823;
  assign new_n9944 = new_n9943 ^ new_n9892;
  assign new_n9945 = new_n9944 ^ new_n9941;
  assign new_n9946 = new_n9945 ^ new_n9939;
  assign new_n9947 = new_n9628 ^ new_n9621;
  assign new_n9948 = ~new_n9947 & new_n9687;
  assign new_n9949 = new_n9645 & new_n9875;
  assign new_n9950 = new_n9949 ^ new_n9714;
  assign new_n9951 = new_n9950 ^ new_n9878;
  assign new_n9952 = new_n9951 ^ new_n9948;
  assign new_n9953 = ~new_n9665 & ~new_n9674;
  assign new_n9954 = new_n9953 ^ new_n9873;
  assign new_n9955 = ~new_n9626 & ~new_n9684;
  assign new_n9956 = new_n9955 ^ new_n9688;
  assign new_n9957 = new_n9956 ^ new_n9876;
  assign new_n9958 = new_n9957 ^ new_n9954;
  assign new_n9959 = new_n9958 ^ new_n9952;
  assign new_n9960 = new_n9959 ^ new_n9946;
  assign new_n9961 = new_n9467 ^ new_n9464;
  assign new_n9962 = new_n9442 ^ new_n9440;
  assign new_n9963 = new_n9962 ^ new_n9867;
  assign new_n9964 = new_n9963 ^ new_n9961;
  assign new_n9965 = new_n9964 ^ new_n9960;
  assign new_n9966 = new_n9481 ^ new_n7594;
  assign new_n9967 = ~new_n9966 & new_n9573;
  assign new_n9968 = new_n9485 & new_n9910;
  assign new_n9969 = new_n9968 ^ new_n9572;
  assign new_n9970 = new_n9969 ^ new_n9913;
  assign new_n9971 = new_n9970 ^ new_n9967;
  assign new_n9972 = ~new_n9518 & ~new_n9536;
  assign new_n9973 = new_n9972 ^ new_n9908;
  assign new_n9974 = ~new_n9500 & new_n9547;
  assign new_n9975 = new_n9974 ^ new_n9574;
  assign new_n9976 = new_n9975 ^ new_n9911;
  assign new_n9977 = new_n9976 ^ new_n9973;
  assign new_n9978 = new_n9977 ^ new_n9971;
  assign new_n9979 = new_n9978 ^ new_n3528;
  assign new_n9980 = new_n9979 ^ new_n9321;
  assign new_n9981 = new_n9980 ^ new_n9927;
  assign new_n9982 = new_n9981 ^ new_n9965;
  assign new_n9983 = new_n9982 ^ new_n9933;
  assign new_n9984 = ~new_n9710 & new_n9601;
  assign new_n9985 = new_n9984 ^ new_n9878;
  assign new_n9986 = new_n9955 ^ new_n9691;
  assign new_n9987 = new_n9986 ^ new_n9685;
  assign new_n9988 = new_n9987 ^ new_n9713;
  assign new_n9989 = new_n9988 ^ new_n9985;
  assign new_n9990 = new_n9737 & new_n9844;
  assign new_n9991 = new_n9990 ^ new_n9894;
  assign new_n9992 = new_n9942 ^ new_n9826;
  assign new_n9993 = new_n9992 ^ new_n9820;
  assign new_n9994 = new_n9993 ^ new_n9847;
  assign new_n9995 = new_n9994 ^ new_n9991;
  assign new_n9996 = new_n9995 ^ new_n9989;
  assign new_n9997 = new_n9856 ^ new_n9447;
  assign new_n9998 = ~new_n9463 & new_n9379;
  assign new_n9999 = new_n9998 ^ new_n9473;
  assign new_n10000 = new_n9999 ^ new_n9997;
  assign new_n10001 = new_n10000 ^ new_n9996;
  assign new_n10002 = ~new_n9568 & new_n9478;
  assign new_n10003 = new_n10002 ^ new_n9913;
  assign new_n10004 = new_n9974 ^ new_n9575;
  assign new_n10005 = new_n10004 ^ new_n9548;
  assign new_n10006 = new_n10005 ^ new_n9571;
  assign new_n10007 = new_n10006 ^ new_n10003;
  assign new_n10008 = new_n10007 ^ new_n3620;
  assign new_n10009 = new_n9853 ^ new_n9302;
  assign new_n10010 = new_n9316 ^ new_n9276;
  assign new_n10011 = new_n10010 ^ new_n9270;
  assign new_n10012 = new_n10011 ^ new_n9295;
  assign new_n10013 = new_n10012 ^ new_n10009;
  assign new_n10014 = new_n10013 ^ new_n10008;
  assign new_n10015 = new_n9853 ^ new_n9293;
  assign new_n10016 = ~new_n9313 & new_n9201;
  assign new_n10017 = new_n10016 ^ new_n9320;
  assign new_n10018 = new_n10017 ^ new_n10015;
  assign new_n10019 = new_n10018 ^ new_n10014;
  assign new_n10020 = new_n10019 ^ new_n10001;
  assign new_n10021 = new_n10020 ^ new_n9983;
  assign new_n10022 = new_n9976 ^ new_n9968;
  assign new_n10023 = new_n10022 ^ new_n9917;
  assign new_n10024 = new_n10023 ^ new_n3660;
  assign new_n10025 = new_n10024 ^ new_n9930;
  assign new_n10026 = new_n9944 ^ new_n9936;
  assign new_n10027 = new_n10026 ^ new_n9898;
  assign new_n10028 = new_n9957 ^ new_n9949;
  assign new_n10029 = new_n10028 ^ new_n9882;
  assign new_n10030 = new_n10029 ^ new_n10027;
  assign new_n10031 = new_n10030 ^ new_n9860;
  assign new_n10032 = new_n10031 ^ new_n10025;
  assign new_n10033 = new_n9990 ^ new_n9845;
  assign new_n10034 = new_n9755 & new_n9888;
  assign new_n10035 = new_n10034 ^ new_n9945;
  assign new_n10036 = new_n10035 ^ new_n10033;
  assign new_n10037 = new_n9984 ^ new_n9711;
  assign new_n10038 = new_n9630 & new_n9872;
  assign new_n10039 = new_n10038 ^ new_n9958;
  assign new_n10040 = new_n10039 ^ new_n10037;
  assign new_n10041 = new_n10040 ^ new_n10036;
  assign new_n10042 = new_n10041 ^ new_n10018;
  assign new_n10043 = new_n10002 ^ new_n9569;
  assign new_n10044 = ~new_n9907 & new_n9488;
  assign new_n10045 = new_n10044 ^ new_n9977;
  assign new_n10046 = new_n10045 ^ new_n10043;
  assign new_n10047 = new_n10046 ^ new_n3645;
  assign new_n10048 = new_n10011 ^ new_n9306;
  assign new_n10049 = ~new_n9391 & ~new_n9450;
  assign new_n10050 = new_n10049 ^ new_n9470;
  assign new_n10051 = new_n10050 ^ new_n9857;
  assign new_n10052 = new_n10051 ^ new_n9457;
  assign new_n10053 = new_n10052 ^ new_n10048;
  assign new_n10054 = new_n10053 ^ new_n10047;
  assign new_n10055 = new_n10054 ^ new_n10042;
  assign new_n10056 = new_n10055 ^ new_n10020;
  assign new_n10057 = new_n10056 ^ new_n10032;
  assign new_n10058 = new_n10005 ^ new_n9969;
  assign new_n10059 = new_n10058 ^ new_n3552;
  assign new_n10060 = new_n9993 ^ new_n9937;
  assign new_n10061 = new_n9987 ^ new_n9950;
  assign new_n10062 = new_n10061 ^ new_n10060;
  assign new_n10063 = new_n10062 ^ new_n10059;
  assign new_n10064 = new_n10063 ^ new_n9860;
  assign new_n10065 = new_n10048 ^ new_n9300;
  assign new_n10066 = new_n9865 ^ new_n9857;
  assign new_n10067 = new_n10049 ^ new_n9468;
  assign new_n10068 = new_n10067 ^ new_n9453;
  assign new_n10069 = new_n10068 ^ new_n10066;
  assign new_n10070 = new_n10069 ^ new_n10065;
  assign new_n10071 = new_n10070 ^ new_n10064;
  assign new_n10072 = new_n10071 ^ new_n10057;
  assign new_n10073 = new_n10032 & new_n10072;
  assign new_n10074 = new_n10073 ^ new_n10071;
  assign new_n10075 = new_n9856 ^ new_n9440;
  assign new_n10076 = new_n10051 ^ new_n9452;
  assign new_n10077 = new_n10076 ^ new_n10075;
  assign new_n10078 = new_n9984 ^ new_n9685;
  assign new_n10079 = new_n10078 ^ new_n9951;
  assign new_n10080 = new_n9990 ^ new_n9820;
  assign new_n10081 = new_n10080 ^ new_n9938;
  assign new_n10082 = new_n10081 ^ new_n10079;
  assign new_n10083 = new_n10082 ^ new_n10077;
  assign new_n10084 = new_n10002 ^ new_n9548;
  assign new_n10085 = new_n10084 ^ new_n9970;
  assign new_n10086 = new_n10085 ^ new_n3473;
  assign new_n10087 = new_n10086 ^ new_n9855;
  assign new_n10088 = new_n10087 ^ new_n10013;
  assign new_n10089 = new_n10088 ^ new_n10083;
  assign new_n10090 = new_n10089 ^ new_n10071;
  assign new_n10091 = new_n10090 ^ new_n9933;
  assign new_n10092 = new_n10071 ^ new_n9932;
  assign new_n10093 = new_n10089 ^ new_n9982;
  assign new_n10094 = new_n10093 ^ new_n10092;
  assign new_n10095 = ~new_n10091 & new_n10094;
  assign new_n10096 = new_n10095 ^ new_n10020;
  assign new_n10097 = new_n10096 ^ new_n10074;
  assign new_n10098 = new_n10055 ^ new_n9983;
  assign new_n10099 = new_n10089 ^ new_n9932;
  assign new_n10100 = ~new_n10098 & ~new_n10099;
  assign new_n10101 = ~new_n10057 & new_n9932;
  assign new_n10102 = new_n10101 ^ new_n9932;
  assign new_n10103 = new_n10102 ^ new_n10100;
  assign new_n10104 = new_n10103 ^ new_n10093;
  assign new_n10105 = ~new_n10021 & new_n10090;
  assign new_n10106 = new_n10071 ^ new_n10055;
  assign new_n10107 = new_n10106 ^ new_n10093;
  assign new_n10108 = new_n10071 ^ new_n9982;
  assign new_n10109 = ~new_n10108 & new_n10107;
  assign new_n10110 = new_n10109 ^ new_n10105;
  assign new_n10111 = new_n10055 ^ new_n9862;
  assign new_n10112 = new_n10111 ^ new_n10110;
  assign new_n10113 = new_n10112 ^ new_n10104;
  assign new_n10114 = new_n10096 ^ new_n10091;
  assign new_n10115 = new_n10091 ^ new_n10032;
  assign new_n10116 = new_n10057 ^ new_n9932;
  assign new_n10117 = new_n10116 ^ new_n10093;
  assign new_n10118 = ~new_n10115 & new_n10117;
  assign new_n10119 = new_n10118 ^ new_n9982;
  assign new_n10120 = new_n10119 ^ new_n10110;
  assign new_n10121 = new_n10120 ^ new_n10114;
  assign new_n10122 = ~new_n10121 & new_n10113;
  assign new_n10123 = new_n10122 ^ new_n10097;
  assign new_n10124 = new_n10091 ^ new_n10056;
  assign new_n10125 = ~new_n10093 & ~new_n10124;
  assign new_n10126 = new_n10125 ^ new_n10105;
  assign new_n10127 = new_n10126 ^ new_n10098;
  assign new_n10128 = new_n10127 ^ new_n10123;
  assign new_n10129 = new_n10089 ^ new_n10057;
  assign new_n10130 = new_n10032 ^ new_n10021;
  assign new_n10131 = ~new_n10130 & new_n10129;
  assign new_n10132 = new_n10131 ^ new_n10101;
  assign new_n10133 = new_n10125 ^ new_n10109;
  assign new_n10134 = new_n10133 ^ new_n10132;
  assign new_n10135 = ~new_n10134 & new_n10128;
  assign new_n10136 = new_n10089 ^ new_n10055;
  assign new_n10137 = new_n10118 ^ new_n10073;
  assign new_n10138 = new_n10137 ^ new_n10133;
  assign new_n10139 = new_n10138 ^ new_n10136;
  assign new_n10140 = new_n10131 ^ new_n10100;
  assign new_n10141 = new_n10140 ^ new_n10089;
  assign new_n10142 = new_n10141 ^ new_n10127;
  assign new_n10143 = new_n10142 ^ new_n10122;
  assign new_n10144 = ~new_n10139 & ~new_n10143;
  assign new_n10145 = new_n10144 ^ new_n10135;
  assign new_n10146 = new_n10141 ^ new_n10097;
  assign new_n10147 = new_n10146 ^ new_n10145;
  assign new_n10148 = ~new_n10021 & ~new_n10147;
  assign new_n10149 = ~new_n10147 & new_n10090;
  assign new_n10150 = new_n10149 ^ new_n10148;
  assign new_n10151 = new_n10135 ^ new_n10089;
  assign new_n10152 = new_n10131 ^ new_n10073;
  assign new_n10153 = new_n10055 ^ new_n9932;
  assign new_n10154 = new_n10118 ^ new_n10102;
  assign new_n10155 = new_n10144 ^ new_n10097;
  assign new_n10156 = new_n10155 ^ new_n10127;
  assign new_n10157 = new_n10135 ^ new_n10122;
  assign new_n10158 = ~new_n10142 & new_n10157;
  assign new_n10159 = new_n10158 ^ new_n10143;
  assign new_n10160 = ~new_n10159 & new_n10156;
  assign new_n10161 = new_n10160 ^ new_n10158;
  assign new_n10162 = new_n10161 ^ new_n10154;
  assign new_n10163 = new_n10162 ^ new_n10153;
  assign new_n10164 = new_n10163 ^ new_n10152;
  assign new_n10165 = new_n10164 ^ new_n10151;
  assign new_n10166 = ~new_n10093 & new_n10165;
  assign new_n10167 = new_n10129 & new_n10156;
  assign new_n10168 = ~new_n10124 & new_n10165;
  assign new_n10169 = new_n10168 ^ new_n10167;
  assign new_n10170 = new_n10142 ^ new_n10135;
  assign new_n10171 = ~new_n10170 & new_n10032;
  assign new_n10172 = new_n10158 ^ new_n10113;
  assign new_n10173 = ~new_n10091 & new_n10172;
  assign new_n10174 = new_n10173 ^ new_n10171;
  assign new_n10175 = new_n10160 ^ new_n10144;
  assign new_n10176 = new_n10175 ^ new_n10121;
  assign new_n10177 = ~new_n10099 & ~new_n10176;
  assign new_n10178 = new_n10177 ^ new_n10174;
  assign new_n10179 = new_n10178 ^ new_n10169;
  assign new_n10180 = new_n10179 ^ new_n10166;
  assign new_n10181 = new_n10180 ^ new_n10150;
  assign new_n10182 = new_n10181 ^ new_n9162;
  assign new_n10183 = new_n10085 ^ n57;
  assign new_n10184 = new_n10183 ^ n25;
  assign new_n10185 = new_n10058 ^ n60;
  assign new_n10186 = new_n10185 ^ n28;
  assign new_n10187 = new_n10186 ^ new_n10184;
  assign new_n10188 = new_n10023 ^ n64;
  assign new_n10189 = new_n10188 ^ n32;
  assign new_n10190 = new_n10046 ^ n59;
  assign new_n10191 = new_n10190 ^ n27;
  assign new_n10192 = new_n10007 ^ n58;
  assign new_n10193 = new_n10192 ^ n26;
  assign new_n10194 = new_n10193 ^ new_n10191;
  assign new_n10195 = ~new_n10189 & ~new_n10194;
  assign new_n10196 = new_n10186 & new_n10189;
  assign new_n10197 = new_n10196 ^ new_n10195;
  assign new_n10198 = new_n10197 ^ new_n10186;
  assign new_n10199 = new_n10194 ^ new_n10189;
  assign new_n10200 = new_n9919 ^ n63;
  assign new_n10201 = new_n10200 ^ n31;
  assign new_n10202 = new_n10201 ^ new_n10199;
  assign new_n10203 = new_n9978 ^ n62;
  assign new_n10204 = new_n10203 ^ n30;
  assign new_n10205 = new_n10204 ^ new_n10184;
  assign new_n10206 = new_n10205 ^ new_n10202;
  assign new_n10207 = new_n9578 ^ n61;
  assign new_n10208 = new_n10207 ^ n29;
  assign new_n10209 = new_n10208 ^ new_n10201;
  assign new_n10210 = new_n10209 ^ new_n10187;
  assign new_n10211 = new_n10210 ^ new_n10189;
  assign new_n10212 = ~new_n10206 & new_n10211;
  assign new_n10213 = new_n10212 ^ new_n10198;
  assign new_n10214 = new_n10204 ^ new_n10186;
  assign new_n10215 = new_n10191 ^ new_n10184;
  assign new_n10216 = new_n10215 ^ new_n10214;
  assign new_n10217 = ~new_n10214 & new_n10216;
  assign new_n10218 = new_n10210 ^ new_n10194;
  assign new_n10219 = ~new_n10205 & ~new_n10218;
  assign new_n10220 = new_n10219 ^ new_n10217;
  assign new_n10221 = new_n10220 ^ new_n10213;
  assign new_n10222 = new_n10221 ^ new_n10215;
  assign new_n10223 = new_n10199 & new_n10201;
  assign new_n10224 = new_n10223 ^ new_n10201;
  assign new_n10225 = new_n10209 ^ new_n10204;
  assign new_n10226 = new_n10225 ^ new_n10191;
  assign new_n10227 = new_n10201 ^ new_n10184;
  assign new_n10228 = ~new_n10226 & ~new_n10227;
  assign new_n10229 = new_n10228 ^ new_n10224;
  assign new_n10230 = new_n10229 ^ new_n10205;
  assign new_n10231 = new_n10225 ^ new_n10193;
  assign new_n10232 = ~new_n10231 & new_n10187;
  assign new_n10233 = new_n10232 ^ new_n10217;
  assign new_n10234 = new_n10208 ^ new_n10191;
  assign new_n10235 = new_n10234 ^ new_n10233;
  assign new_n10236 = new_n10235 ^ new_n10230;
  assign new_n10237 = new_n10201 ^ new_n10186;
  assign new_n10238 = new_n10237 ^ new_n10205;
  assign new_n10239 = ~new_n10210 & new_n10238;
  assign new_n10240 = new_n10239 ^ new_n10193;
  assign new_n10241 = new_n10240 ^ new_n10210;
  assign new_n10242 = new_n10232 ^ new_n10212;
  assign new_n10243 = new_n10217 ^ new_n10204;
  assign new_n10244 = new_n10243 ^ new_n10242;
  assign new_n10245 = new_n10244 ^ new_n10241;
  assign new_n10246 = ~new_n10245 & new_n10236;
  assign new_n10247 = new_n10232 ^ new_n10219;
  assign new_n10248 = new_n10247 ^ new_n10226;
  assign new_n10249 = new_n10199 ^ new_n10184;
  assign new_n10250 = new_n10231 ^ new_n10189;
  assign new_n10251 = ~new_n10249 & new_n10250;
  assign new_n10252 = new_n10251 ^ new_n10228;
  assign new_n10253 = new_n10252 ^ new_n10184;
  assign new_n10254 = new_n10253 ^ new_n10248;
  assign new_n10255 = new_n10254 ^ new_n10246;
  assign new_n10256 = ~new_n10222 & ~new_n10255;
  assign new_n10257 = new_n10240 ^ new_n10197;
  assign new_n10258 = new_n10257 ^ new_n10246;
  assign new_n10259 = new_n10258 ^ new_n10248;
  assign new_n10260 = new_n10251 ^ new_n10223;
  assign new_n10261 = new_n10260 ^ new_n10220;
  assign new_n10262 = ~new_n10261 & new_n10259;
  assign new_n10263 = new_n10262 ^ new_n10256;
  assign new_n10264 = new_n10257 ^ new_n10253;
  assign new_n10265 = new_n10264 ^ new_n10263;
  assign new_n10266 = ~new_n10265 & new_n10187;
  assign new_n10267 = ~new_n10231 & ~new_n10265;
  assign new_n10268 = new_n10267 ^ new_n10266;
  assign new_n10269 = new_n10251 ^ new_n10198;
  assign new_n10270 = new_n10201 ^ new_n10191;
  assign new_n10271 = new_n10224 ^ new_n10212;
  assign new_n10272 = new_n10257 ^ new_n10256;
  assign new_n10273 = new_n10272 ^ new_n10248;
  assign new_n10274 = new_n10262 ^ new_n10246;
  assign new_n10275 = ~new_n10254 & new_n10274;
  assign new_n10276 = new_n10275 ^ new_n10255;
  assign new_n10277 = ~new_n10276 & new_n10273;
  assign new_n10278 = new_n10277 ^ new_n10275;
  assign new_n10279 = new_n10278 ^ new_n10271;
  assign new_n10280 = new_n10279 ^ new_n10270;
  assign new_n10281 = new_n10280 ^ new_n10184;
  assign new_n10282 = new_n10281 ^ new_n10262;
  assign new_n10283 = new_n10282 ^ new_n10269;
  assign new_n10284 = ~new_n10205 & new_n10283;
  assign new_n10285 = ~new_n10249 & new_n10273;
  assign new_n10286 = ~new_n10218 & new_n10283;
  assign new_n10287 = new_n10286 ^ new_n10285;
  assign new_n10288 = new_n10262 ^ new_n10254;
  assign new_n10289 = ~new_n10189 & ~new_n10288;
  assign new_n10290 = new_n10275 ^ new_n10236;
  assign new_n10291 = ~new_n10210 & new_n10290;
  assign new_n10292 = new_n10291 ^ new_n10289;
  assign new_n10293 = new_n10277 ^ new_n10256;
  assign new_n10294 = new_n10293 ^ new_n10245;
  assign new_n10295 = ~new_n10227 & ~new_n10294;
  assign new_n10296 = new_n10295 ^ new_n10292;
  assign new_n10297 = new_n10296 ^ new_n10287;
  assign new_n10298 = new_n10297 ^ new_n10284;
  assign new_n10299 = new_n10298 ^ new_n10268;
  assign new_n10300 = new_n10299 ^ new_n8226;
  assign new_n10301 = new_n5520 ^ new_n1402;
  assign new_n10302 = new_n10301 ^ new_n9611;
  assign new_n10303 = new_n5667 ^ new_n5601;
  assign new_n10304 = new_n10303 ^ new_n5654;
  assign new_n10305 = new_n10304 ^ new_n10302;
  assign new_n10306 = new_n5492 ^ new_n5309;
  assign new_n10307 = new_n9619 ^ new_n4615;
  assign new_n10308 = new_n10307 ^ new_n10306;
  assign new_n10309 = new_n10308 ^ new_n10305;
  assign new_n10310 = new_n5561 ^ new_n5451;
  assign new_n10311 = new_n5612 ^ new_n4731;
  assign new_n10312 = new_n10311 ^ new_n5037;
  assign new_n10313 = new_n10312 ^ new_n10310;
  assign new_n10314 = new_n5687 ^ new_n4752;
  assign new_n10315 = new_n9588 ^ new_n5663;
  assign new_n10316 = new_n10315 ^ new_n10314;
  assign new_n10317 = new_n10316 ^ new_n10313;
  assign new_n10318 = new_n10317 ^ new_n10309;
  assign new_n10319 = new_n9611 ^ new_n5552;
  assign new_n10320 = new_n10319 ^ new_n5633;
  assign new_n10321 = new_n5575 ^ new_n4703;
  assign new_n10322 = new_n10321 ^ new_n5677;
  assign new_n10323 = new_n10322 ^ new_n10320;
  assign new_n10324 = new_n10323 ^ new_n10308;
  assign new_n10325 = new_n5617 ^ new_n5539;
  assign new_n10326 = new_n5037 ^ new_n4633;
  assign new_n10327 = new_n10326 ^ new_n5492;
  assign new_n10328 = new_n10327 ^ new_n10325;
  assign new_n10329 = new_n10328 ^ new_n10308;
  assign new_n10330 = new_n5639 ^ new_n4663;
  assign new_n10331 = new_n9611 ^ new_n5576;
  assign new_n10332 = new_n10331 ^ new_n10330;
  assign new_n10333 = new_n10332 ^ new_n10329;
  assign new_n10334 = new_n10333 ^ new_n10323;
  assign new_n10335 = new_n10334 ^ new_n10317;
  assign new_n10336 = new_n10313 ^ new_n10305;
  assign new_n10337 = new_n5680 ^ new_n5654;
  assign new_n10338 = new_n10337 ^ new_n5687;
  assign new_n10339 = new_n9611 ^ new_n4776;
  assign new_n10340 = new_n10339 ^ new_n5589;
  assign new_n10341 = new_n10340 ^ new_n10338;
  assign new_n10342 = new_n10341 ^ new_n10323;
  assign new_n10343 = new_n10342 ^ new_n10336;
  assign new_n10344 = new_n10343 ^ new_n10332;
  assign new_n10345 = new_n10335 & new_n10344;
  assign new_n10346 = ~new_n10323 & ~new_n10333;
  assign new_n10347 = new_n10346 ^ new_n10323;
  assign new_n10348 = new_n10347 ^ new_n10345;
  assign new_n10349 = new_n10313 ^ new_n10308;
  assign new_n10350 = new_n10333 ^ new_n10305;
  assign new_n10351 = new_n10332 & new_n10350;
  assign new_n10352 = new_n10351 ^ new_n10345;
  assign new_n10353 = new_n10316 ^ new_n10305;
  assign new_n10354 = ~new_n10318 & new_n10353;
  assign new_n10355 = new_n10343 ^ new_n10329;
  assign new_n10356 = new_n10317 & new_n10355;
  assign new_n10357 = new_n10356 ^ new_n10354;
  assign new_n10358 = new_n10357 ^ new_n10352;
  assign new_n10359 = new_n10358 ^ new_n10349;
  assign new_n10360 = new_n10342 ^ new_n10316;
  assign new_n10361 = new_n10360 ^ new_n10308;
  assign new_n10362 = new_n10323 ^ new_n10313;
  assign new_n10363 = ~new_n10361 & new_n10362;
  assign new_n10364 = new_n10363 ^ new_n10347;
  assign new_n10365 = new_n10364 ^ new_n10317;
  assign new_n10366 = new_n10360 ^ new_n10328;
  assign new_n10367 = ~new_n10366 & new_n10336;
  assign new_n10368 = new_n10367 ^ new_n10354;
  assign new_n10369 = new_n10341 ^ new_n10308;
  assign new_n10370 = new_n10369 ^ new_n10368;
  assign new_n10371 = new_n10370 ^ new_n10365;
  assign new_n10372 = new_n10323 ^ new_n10305;
  assign new_n10373 = new_n10372 ^ new_n10317;
  assign new_n10374 = new_n10343 & new_n10373;
  assign new_n10375 = new_n10374 ^ new_n10328;
  assign new_n10376 = new_n10375 ^ new_n10343;
  assign new_n10377 = new_n10368 ^ new_n10345;
  assign new_n10378 = new_n10377 ^ new_n10316;
  assign new_n10379 = new_n10378 ^ new_n10376;
  assign new_n10380 = ~new_n10379 & new_n10371;
  assign new_n10381 = new_n10367 ^ new_n10356;
  assign new_n10382 = new_n10381 ^ new_n10361;
  assign new_n10383 = new_n10366 ^ new_n10332;
  assign new_n10384 = new_n10333 ^ new_n10313;
  assign new_n10385 = ~new_n10383 & new_n10384;
  assign new_n10386 = new_n10385 ^ new_n10363;
  assign new_n10387 = new_n10386 ^ new_n10313;
  assign new_n10388 = new_n10387 ^ new_n10382;
  assign new_n10389 = new_n10388 ^ new_n10380;
  assign new_n10390 = ~new_n10359 & ~new_n10389;
  assign new_n10391 = new_n10351 ^ new_n10305;
  assign new_n10392 = new_n10391 ^ new_n10375;
  assign new_n10393 = new_n10392 ^ new_n10390;
  assign new_n10394 = new_n10393 ^ new_n10382;
  assign new_n10395 = new_n10392 ^ new_n10380;
  assign new_n10396 = new_n10395 ^ new_n10382;
  assign new_n10397 = new_n10385 ^ new_n10346;
  assign new_n10398 = new_n10397 ^ new_n10357;
  assign new_n10399 = ~new_n10398 & new_n10396;
  assign new_n10400 = new_n10399 ^ new_n10380;
  assign new_n10401 = ~new_n10388 & ~new_n10400;
  assign new_n10402 = new_n10401 ^ new_n10380;
  assign new_n10403 = new_n10394 & new_n10402;
  assign new_n10404 = new_n10401 ^ new_n10388;
  assign new_n10405 = new_n10404 ^ new_n10403;
  assign new_n10406 = new_n10405 ^ new_n10348;
  assign new_n10407 = new_n10406 ^ new_n10324;
  assign new_n10408 = new_n10407 ^ new_n10305;
  assign new_n10409 = new_n10390 ^ new_n10363;
  assign new_n10410 = new_n10409 ^ new_n10375;
  assign new_n10411 = new_n10410 ^ new_n10408;
  assign new_n10412 = ~new_n10318 & new_n10411;
  assign new_n10413 = new_n10399 ^ new_n10390;
  assign new_n10414 = new_n10392 ^ new_n10387;
  assign new_n10415 = new_n10414 ^ new_n10413;
  assign new_n10416 = ~new_n10366 & ~new_n10415;
  assign new_n10417 = new_n10416 ^ new_n10412;
  assign new_n10418 = new_n10353 & new_n10411;
  assign new_n10419 = ~new_n10415 & new_n10336;
  assign new_n10420 = new_n10419 ^ new_n10418;
  assign new_n10421 = new_n10404 ^ new_n10399;
  assign new_n10422 = new_n10421 ^ new_n10398;
  assign new_n10423 = new_n10335 & new_n10422;
  assign new_n10424 = new_n10423 ^ new_n10420;
  assign new_n10425 = new_n10404 ^ new_n10371;
  assign new_n10426 = ~new_n10425 & new_n10373;
  assign new_n10427 = new_n10344 & new_n10422;
  assign new_n10428 = ~new_n10425 & new_n10343;
  assign new_n10429 = new_n10428 ^ new_n10427;
  assign new_n10430 = new_n10429 ^ new_n10426;
  assign new_n10431 = new_n10430 ^ new_n10424;
  assign new_n10432 = new_n10431 ^ new_n10417;
  assign new_n10433 = new_n9748 ^ new_n7439;
  assign new_n10434 = new_n10433 ^ new_n7655;
  assign new_n10435 = new_n8233 ^ new_n7479;
  assign new_n10436 = new_n10435 ^ new_n7521;
  assign new_n10437 = new_n10436 ^ new_n10434;
  assign new_n10438 = new_n9748 ^ new_n8235;
  assign new_n10439 = new_n10438 ^ new_n7512;
  assign new_n10440 = new_n7628 ^ new_n7607;
  assign new_n10441 = new_n10440 ^ new_n10439;
  assign new_n10442 = new_n10441 ^ new_n10437;
  assign new_n10443 = new_n8242 ^ new_n7454;
  assign new_n10444 = new_n7529 ^ new_n7500;
  assign new_n10445 = new_n10444 ^ new_n7616;
  assign new_n10446 = new_n10445 ^ new_n10443;
  assign new_n10447 = new_n10446 ^ new_n10442;
  assign new_n10448 = new_n7587 ^ new_n7253;
  assign new_n10449 = new_n8225 ^ new_n7547;
  assign new_n10450 = new_n10449 ^ new_n7579;
  assign new_n10451 = new_n10450 ^ new_n10448;
  assign new_n10452 = new_n10451 ^ new_n10447;
  assign new_n10453 = new_n9748 ^ new_n7583;
  assign new_n10454 = new_n8238 ^ new_n7608;
  assign new_n10455 = new_n10454 ^ new_n7633;
  assign new_n10456 = new_n10455 ^ new_n10453;
  assign new_n10457 = new_n7566 ^ new_n7424;
  assign new_n10458 = new_n8231 ^ new_n6981;
  assign new_n10459 = new_n10458 ^ new_n7547;
  assign new_n10460 = new_n10459 ^ new_n10457;
  assign new_n10461 = new_n10460 ^ new_n10456;
  assign new_n10462 = new_n10461 ^ new_n10442;
  assign new_n10463 = new_n10456 ^ new_n10437;
  assign new_n10464 = new_n10460 ^ new_n10446;
  assign new_n10465 = new_n10464 ^ new_n10463;
  assign new_n10466 = new_n10462 & new_n10465;
  assign new_n10467 = new_n10466 ^ new_n10451;
  assign new_n10468 = new_n9748 ^ new_n7652;
  assign new_n10469 = new_n8229 ^ new_n7486;
  assign new_n10470 = new_n10469 ^ new_n7417;
  assign new_n10471 = new_n10470 ^ new_n10468;
  assign new_n10472 = new_n7579 ^ new_n7560;
  assign new_n10473 = new_n9759 ^ new_n8227;
  assign new_n10474 = new_n10473 ^ new_n10472;
  assign new_n10475 = new_n10474 ^ new_n10451;
  assign new_n10476 = ~new_n10475 & new_n10471;
  assign new_n10477 = ~new_n10471 & new_n10456;
  assign new_n10478 = new_n10477 ^ new_n10476;
  assign new_n10479 = new_n10478 ^ new_n10467;
  assign new_n10480 = new_n10474 ^ new_n10447;
  assign new_n10481 = new_n10460 ^ new_n10437;
  assign new_n10482 = new_n10480 & new_n10481;
  assign new_n10483 = new_n10475 ^ new_n10471;
  assign new_n10484 = ~new_n10437 & ~new_n10483;
  assign new_n10485 = new_n10484 ^ new_n10437;
  assign new_n10486 = new_n10485 ^ new_n10482;
  assign new_n10487 = new_n10486 ^ new_n10464;
  assign new_n10488 = new_n10452 & new_n10461;
  assign new_n10489 = new_n10474 ^ new_n10456;
  assign new_n10490 = new_n10489 ^ new_n10464;
  assign new_n10491 = new_n10456 ^ new_n10446;
  assign new_n10492 = new_n10490 & new_n10491;
  assign new_n10493 = new_n10492 ^ new_n10488;
  assign new_n10494 = new_n10474 ^ new_n10441;
  assign new_n10495 = new_n10494 ^ new_n10493;
  assign new_n10496 = new_n10495 ^ new_n10487;
  assign new_n10497 = new_n10467 ^ new_n10462;
  assign new_n10498 = new_n10471 ^ new_n10462;
  assign new_n10499 = new_n10483 ^ new_n10437;
  assign new_n10500 = new_n10499 ^ new_n10464;
  assign new_n10501 = new_n10498 & new_n10500;
  assign new_n10502 = new_n10501 ^ new_n10493;
  assign new_n10503 = new_n10502 ^ new_n10446;
  assign new_n10504 = new_n10503 ^ new_n10497;
  assign new_n10505 = ~new_n10496 & new_n10504;
  assign new_n10506 = new_n10505 ^ new_n10479;
  assign new_n10507 = new_n10475 ^ new_n10462;
  assign new_n10508 = new_n10464 & new_n10507;
  assign new_n10509 = new_n10508 ^ new_n10488;
  assign new_n10510 = new_n10509 ^ new_n10480;
  assign new_n10511 = new_n10510 ^ new_n10506;
  assign new_n10512 = new_n10483 ^ new_n10460;
  assign new_n10513 = new_n10471 ^ new_n10452;
  assign new_n10514 = new_n10512 & new_n10513;
  assign new_n10515 = new_n10514 ^ new_n10484;
  assign new_n10516 = new_n10508 ^ new_n10492;
  assign new_n10517 = new_n10516 ^ new_n10515;
  assign new_n10518 = ~new_n10517 & new_n10511;
  assign new_n10519 = new_n10474 ^ new_n10460;
  assign new_n10520 = new_n10478 ^ new_n10456;
  assign new_n10521 = new_n10520 ^ new_n10501;
  assign new_n10522 = new_n10521 ^ new_n10516;
  assign new_n10523 = new_n10522 ^ new_n10519;
  assign new_n10524 = new_n10514 ^ new_n10482;
  assign new_n10525 = new_n10524 ^ new_n10460;
  assign new_n10526 = new_n10525 ^ new_n10510;
  assign new_n10527 = new_n10526 ^ new_n10505;
  assign new_n10528 = new_n10523 & new_n10527;
  assign new_n10529 = new_n10528 ^ new_n10518;
  assign new_n10530 = new_n10525 ^ new_n10479;
  assign new_n10531 = new_n10530 ^ new_n10529;
  assign new_n10532 = new_n10452 & new_n10531;
  assign new_n10533 = new_n10461 & new_n10531;
  assign new_n10534 = new_n10533 ^ new_n10532;
  assign new_n10535 = new_n10528 ^ new_n10479;
  assign new_n10536 = new_n10535 ^ new_n10510;
  assign new_n10537 = new_n10518 ^ new_n10505;
  assign new_n10538 = new_n10526 & new_n10537;
  assign new_n10539 = new_n10538 ^ new_n10527;
  assign new_n10540 = new_n10536 & new_n10539;
  assign new_n10541 = new_n10540 ^ new_n10528;
  assign new_n10542 = new_n10541 ^ new_n10504;
  assign new_n10543 = new_n10481 & new_n10542;
  assign new_n10544 = new_n10526 ^ new_n10518;
  assign new_n10545 = new_n10471 & new_n10544;
  assign new_n10546 = new_n10538 ^ new_n10496;
  assign new_n10547 = ~new_n10546 & new_n10462;
  assign new_n10548 = new_n10547 ^ new_n10545;
  assign new_n10549 = new_n10548 ^ new_n10543;
  assign new_n10550 = new_n10518 ^ new_n10460;
  assign new_n10551 = new_n10474 ^ new_n10437;
  assign new_n10552 = new_n10501 ^ new_n10485;
  assign new_n10553 = new_n10540 ^ new_n10538;
  assign new_n10554 = new_n10553 ^ new_n10552;
  assign new_n10555 = new_n10554 ^ new_n10551;
  assign new_n10556 = new_n10520 ^ new_n10514;
  assign new_n10557 = new_n10556 ^ new_n10555;
  assign new_n10558 = new_n10557 ^ new_n10550;
  assign new_n10559 = ~new_n10558 & new_n10507;
  assign new_n10560 = new_n10512 & new_n10536;
  assign new_n10561 = new_n10560 ^ new_n10559;
  assign new_n10562 = new_n10561 ^ new_n10549;
  assign new_n10563 = ~new_n10558 & new_n10464;
  assign new_n10564 = new_n10563 ^ new_n10562;
  assign new_n10565 = new_n10564 ^ new_n10534;
  assign new_n10566 = new_n10419 ^ new_n10416;
  assign new_n10567 = new_n10403 ^ new_n10390;
  assign new_n10568 = new_n10567 ^ new_n10379;
  assign new_n10569 = ~new_n10568 & new_n10362;
  assign new_n10570 = new_n10399 ^ new_n10388;
  assign new_n10571 = ~new_n10570 & new_n10332;
  assign new_n10572 = new_n10571 ^ new_n10428;
  assign new_n10573 = new_n10572 ^ new_n10569;
  assign new_n10574 = new_n10399 ^ new_n10313;
  assign new_n10575 = new_n10385 ^ new_n10351;
  assign new_n10576 = new_n10575 ^ new_n10407;
  assign new_n10577 = new_n10576 ^ new_n10574;
  assign new_n10578 = ~new_n10577 & new_n10355;
  assign new_n10579 = new_n10384 & new_n10394;
  assign new_n10580 = new_n10579 ^ new_n10578;
  assign new_n10581 = new_n10580 ^ new_n10573;
  assign new_n10582 = ~new_n10577 & new_n10317;
  assign new_n10583 = new_n10582 ^ new_n10581;
  assign new_n10584 = new_n10583 ^ new_n10566;
  assign new_n10585 = new_n10584 ^ new_n10565;
  assign new_n10586 = new_n10585 ^ new_n10432;
  assign new_n10587 = new_n8581 ^ new_n8564;
  assign new_n10588 = new_n10587 ^ new_n8589;
  assign new_n10589 = new_n10588 ^ new_n8547;
  assign new_n10590 = new_n8547 ^ new_n8542;
  assign new_n10591 = new_n10590 ^ new_n8553;
  assign new_n10592 = ~new_n8564 & new_n10591;
  assign new_n10593 = new_n10592 ^ new_n8564;
  assign new_n10594 = new_n10588 ^ new_n8542;
  assign new_n10595 = new_n8572 ^ new_n8564;
  assign new_n10596 = ~new_n10594 & new_n10595;
  assign new_n10597 = new_n10596 ^ new_n10593;
  assign new_n10598 = new_n8589 ^ new_n8572;
  assign new_n10599 = new_n10598 ^ new_n10597;
  assign new_n10600 = new_n8542 ^ new_n8533;
  assign new_n10601 = new_n10600 ^ new_n10598;
  assign new_n10602 = new_n8589 ^ new_n8533;
  assign new_n10603 = ~new_n10601 & new_n10602;
  assign new_n10604 = new_n8572 ^ new_n8533;
  assign new_n10605 = ~new_n10589 & new_n10604;
  assign new_n10606 = new_n10605 ^ new_n10603;
  assign new_n10607 = new_n8581 ^ new_n8542;
  assign new_n10608 = new_n10607 ^ new_n10606;
  assign new_n10609 = new_n10608 ^ new_n10599;
  assign new_n10610 = new_n10604 ^ new_n10587;
  assign new_n10611 = new_n8564 ^ new_n8533;
  assign new_n10612 = new_n10611 ^ new_n10598;
  assign new_n10613 = new_n10610 & new_n10612;
  assign new_n10614 = new_n10613 ^ new_n8547;
  assign new_n10615 = new_n10614 ^ new_n10610;
  assign new_n10616 = new_n10591 ^ new_n8564;
  assign new_n10617 = new_n10616 ^ new_n10598;
  assign new_n10618 = new_n10610 ^ new_n8553;
  assign new_n10619 = ~new_n10617 & ~new_n10618;
  assign new_n10620 = new_n10619 ^ new_n8589;
  assign new_n10621 = new_n10620 ^ new_n10606;
  assign new_n10622 = new_n10621 ^ new_n10615;
  assign new_n10623 = ~new_n10622 & new_n10609;
  assign new_n10624 = new_n10610 ^ new_n10590;
  assign new_n10625 = new_n10598 & new_n10624;
  assign new_n10626 = new_n10625 ^ new_n10605;
  assign new_n10627 = new_n10626 ^ new_n10594;
  assign new_n10628 = new_n10589 ^ new_n8553;
  assign new_n10629 = new_n10591 ^ new_n8572;
  assign new_n10630 = ~new_n10629 & new_n10628;
  assign new_n10631 = new_n10630 ^ new_n10596;
  assign new_n10632 = new_n10631 ^ new_n8572;
  assign new_n10633 = new_n10632 ^ new_n10627;
  assign new_n10634 = new_n10633 ^ new_n10623;
  assign new_n10635 = new_n8572 ^ new_n8542;
  assign new_n10636 = new_n10591 ^ new_n8533;
  assign new_n10637 = ~new_n8553 & ~new_n10636;
  assign new_n10638 = new_n10637 ^ new_n10619;
  assign new_n10639 = new_n10625 ^ new_n10603;
  assign new_n10640 = new_n10639 ^ new_n10638;
  assign new_n10641 = new_n10640 ^ new_n10635;
  assign new_n10642 = ~new_n10634 & ~new_n10641;
  assign new_n10643 = new_n10637 ^ new_n8533;
  assign new_n10644 = new_n10643 ^ new_n10614;
  assign new_n10645 = new_n10644 ^ new_n10623;
  assign new_n10646 = new_n10645 ^ new_n10627;
  assign new_n10647 = new_n10630 ^ new_n10592;
  assign new_n10648 = new_n10647 ^ new_n10639;
  assign new_n10649 = ~new_n10648 & new_n10646;
  assign new_n10650 = new_n10649 ^ new_n10642;
  assign new_n10651 = new_n10644 ^ new_n10632;
  assign new_n10652 = new_n10651 ^ new_n10650;
  assign new_n10653 = ~new_n10589 & ~new_n10652;
  assign new_n10654 = new_n8564 ^ new_n8542;
  assign new_n10655 = new_n10619 ^ new_n10593;
  assign new_n10656 = new_n10649 ^ new_n10623;
  assign new_n10657 = ~new_n10656 & new_n10633;
  assign new_n10658 = new_n10657 ^ new_n10649;
  assign new_n10659 = new_n10644 ^ new_n10642;
  assign new_n10660 = new_n10659 ^ new_n10627;
  assign new_n10661 = ~new_n10658 & new_n10660;
  assign new_n10662 = new_n10658 ^ new_n10634;
  assign new_n10663 = new_n10662 ^ new_n10661;
  assign new_n10664 = new_n10663 ^ new_n10655;
  assign new_n10665 = new_n10664 ^ new_n10654;
  assign new_n10666 = new_n10665 ^ new_n8533;
  assign new_n10667 = new_n10642 ^ new_n10596;
  assign new_n10668 = new_n10667 ^ new_n10614;
  assign new_n10669 = new_n10668 ^ new_n10666;
  assign new_n10670 = ~new_n10601 & ~new_n10669;
  assign new_n10671 = new_n10670 ^ new_n10653;
  assign new_n10672 = new_n10662 ^ new_n10609;
  assign new_n10673 = new_n10610 & new_n10672;
  assign new_n10674 = new_n10662 ^ new_n10649;
  assign new_n10675 = new_n10674 ^ new_n10648;
  assign new_n10676 = ~new_n10618 & ~new_n10675;
  assign new_n10677 = new_n10676 ^ new_n10673;
  assign new_n10678 = new_n10612 & new_n10672;
  assign new_n10679 = new_n10678 ^ new_n10677;
  assign new_n10680 = ~new_n10669 & new_n10602;
  assign new_n10681 = ~new_n10652 & new_n10604;
  assign new_n10682 = new_n10681 ^ new_n10680;
  assign new_n10683 = ~new_n10617 & ~new_n10675;
  assign new_n10684 = new_n10683 ^ new_n10682;
  assign new_n10685 = new_n10684 ^ new_n10679;
  assign new_n10686 = new_n10685 ^ new_n10671;
  assign new_n10687 = new_n10686 ^ new_n8357;
  assign new_n10688 = new_n7540 ^ new_n6570;
  assign new_n10689 = new_n8710 ^ new_n6531;
  assign new_n10690 = new_n10689 ^ new_n10688;
  assign new_n10691 = new_n8729 ^ new_n6643;
  assign new_n10692 = new_n6690 ^ new_n1012;
  assign new_n10693 = new_n10692 ^ new_n10691;
  assign new_n10694 = new_n6671 ^ new_n6617;
  assign new_n10695 = new_n10694 ^ new_n8751;
  assign new_n10696 = new_n7464 ^ new_n6654;
  assign new_n10697 = new_n10696 ^ new_n10695;
  assign new_n10698 = new_n6716 ^ new_n6671;
  assign new_n10699 = new_n10698 ^ new_n8734;
  assign new_n10700 = new_n7622 ^ new_n6485;
  assign new_n10701 = new_n10700 ^ new_n10699;
  assign new_n10702 = new_n10701 ^ new_n10697;
  assign new_n10703 = new_n10702 ^ new_n10693;
  assign new_n10704 = new_n10703 ^ new_n10690;
  assign new_n10705 = new_n7574 ^ new_n6546;
  assign new_n10706 = new_n8743 ^ new_n6074;
  assign new_n10707 = new_n10706 ^ new_n10705;
  assign new_n10708 = new_n10707 ^ new_n10690;
  assign new_n10709 = new_n7648 ^ new_n6623;
  assign new_n10710 = new_n8705 ^ new_n6671;
  assign new_n10711 = new_n10710 ^ new_n10709;
  assign new_n10712 = new_n10711 ^ new_n10708;
  assign new_n10713 = ~new_n10697 & ~new_n10712;
  assign new_n10714 = new_n10713 ^ new_n10697;
  assign new_n10715 = new_n10707 ^ new_n10703;
  assign new_n10716 = new_n8703 ^ new_n6585;
  assign new_n10717 = new_n6843 ^ new_n6462;
  assign new_n10718 = new_n10717 ^ new_n10716;
  assign new_n10719 = new_n10718 ^ new_n10697;
  assign new_n10720 = new_n10715 & new_n10719;
  assign new_n10721 = new_n10720 ^ new_n10714;
  assign new_n10722 = new_n10718 ^ new_n10693;
  assign new_n10723 = new_n10722 ^ new_n10721;
  assign new_n10724 = new_n6701 ^ new_n6671;
  assign new_n10725 = new_n10724 ^ new_n8717;
  assign new_n10726 = new_n7593 ^ new_n6477;
  assign new_n10727 = new_n10726 ^ new_n10725;
  assign new_n10728 = new_n10727 ^ new_n10707;
  assign new_n10729 = new_n10728 ^ new_n10722;
  assign new_n10730 = new_n10727 ^ new_n10693;
  assign new_n10731 = new_n10729 & new_n10730;
  assign new_n10732 = new_n10727 ^ new_n10718;
  assign new_n10733 = new_n10704 & new_n10732;
  assign new_n10734 = new_n10733 ^ new_n10731;
  assign new_n10735 = new_n10707 ^ new_n10701;
  assign new_n10736 = new_n10735 ^ new_n10734;
  assign new_n10737 = new_n10736 ^ new_n10723;
  assign new_n10738 = new_n10732 ^ new_n10702;
  assign new_n10739 = new_n10727 ^ new_n10697;
  assign new_n10740 = new_n10739 ^ new_n10722;
  assign new_n10741 = new_n10738 & new_n10740;
  assign new_n10742 = new_n10741 ^ new_n10690;
  assign new_n10743 = new_n10742 ^ new_n10738;
  assign new_n10744 = new_n10738 ^ new_n10711;
  assign new_n10745 = new_n10712 ^ new_n10697;
  assign new_n10746 = new_n10745 ^ new_n10722;
  assign new_n10747 = new_n10744 & new_n10746;
  assign new_n10748 = new_n10747 ^ new_n10734;
  assign new_n10749 = new_n10748 ^ new_n10693;
  assign new_n10750 = new_n10749 ^ new_n10743;
  assign new_n10751 = ~new_n10737 & new_n10750;
  assign new_n10752 = new_n10738 ^ new_n10708;
  assign new_n10753 = new_n10722 & new_n10752;
  assign new_n10754 = new_n10753 ^ new_n10733;
  assign new_n10755 = new_n10754 ^ new_n10715;
  assign new_n10756 = new_n10711 ^ new_n10704;
  assign new_n10757 = new_n10718 ^ new_n10712;
  assign new_n10758 = new_n10756 & new_n10757;
  assign new_n10759 = new_n10758 ^ new_n10720;
  assign new_n10760 = new_n10759 ^ new_n10718;
  assign new_n10761 = new_n10760 ^ new_n10755;
  assign new_n10762 = new_n10761 ^ new_n10751;
  assign new_n10763 = new_n10718 ^ new_n10707;
  assign new_n10764 = new_n10727 ^ new_n10712;
  assign new_n10765 = new_n10711 & new_n10764;
  assign new_n10766 = new_n10765 ^ new_n10747;
  assign new_n10767 = new_n10753 ^ new_n10731;
  assign new_n10768 = new_n10767 ^ new_n10766;
  assign new_n10769 = new_n10768 ^ new_n10763;
  assign new_n10770 = new_n10762 & new_n10769;
  assign new_n10771 = new_n10765 ^ new_n10727;
  assign new_n10772 = new_n10771 ^ new_n10742;
  assign new_n10773 = new_n10772 ^ new_n10751;
  assign new_n10774 = new_n10773 ^ new_n10755;
  assign new_n10775 = new_n10758 ^ new_n10713;
  assign new_n10776 = new_n10775 ^ new_n10767;
  assign new_n10777 = ~new_n10776 & new_n10774;
  assign new_n10778 = new_n10777 ^ new_n10770;
  assign new_n10779 = new_n10772 ^ new_n10760;
  assign new_n10780 = new_n10779 ^ new_n10778;
  assign new_n10781 = new_n10704 & new_n10780;
  assign new_n10782 = new_n10707 ^ new_n10697;
  assign new_n10783 = new_n10747 ^ new_n10714;
  assign new_n10784 = new_n10777 ^ new_n10751;
  assign new_n10785 = ~new_n10761 & ~new_n10784;
  assign new_n10786 = new_n10785 ^ new_n10777;
  assign new_n10787 = new_n10772 ^ new_n10770;
  assign new_n10788 = new_n10787 ^ new_n10755;
  assign new_n10789 = ~new_n10786 & new_n10788;
  assign new_n10790 = new_n10786 ^ new_n10762;
  assign new_n10791 = new_n10790 ^ new_n10789;
  assign new_n10792 = new_n10791 ^ new_n10783;
  assign new_n10793 = new_n10792 ^ new_n10782;
  assign new_n10794 = new_n10793 ^ new_n10727;
  assign new_n10795 = new_n10770 ^ new_n10720;
  assign new_n10796 = new_n10795 ^ new_n10742;
  assign new_n10797 = new_n10796 ^ new_n10794;
  assign new_n10798 = new_n10729 & new_n10797;
  assign new_n10799 = new_n10798 ^ new_n10781;
  assign new_n10800 = new_n10730 & new_n10797;
  assign new_n10801 = new_n10732 & new_n10780;
  assign new_n10802 = new_n10801 ^ new_n10800;
  assign new_n10803 = new_n10790 ^ new_n10777;
  assign new_n10804 = new_n10803 ^ new_n10776;
  assign new_n10805 = new_n10746 & new_n10804;
  assign new_n10806 = new_n10805 ^ new_n10802;
  assign new_n10807 = new_n10790 ^ new_n10737;
  assign new_n10808 = new_n10740 & new_n10807;
  assign new_n10809 = new_n10744 & new_n10804;
  assign new_n10810 = new_n10738 & new_n10807;
  assign new_n10811 = new_n10810 ^ new_n10809;
  assign new_n10812 = new_n10811 ^ new_n10808;
  assign new_n10813 = new_n10812 ^ new_n10806;
  assign new_n10814 = new_n10813 ^ new_n10799;
  assign new_n10815 = new_n10814 ^ new_n10687;
  assign new_n10816 = new_n4589 ^ new_n2930;
  assign new_n10817 = new_n5473 ^ n43;
  assign new_n10818 = new_n10817 ^ new_n4649;
  assign new_n10819 = new_n10818 ^ new_n4573;
  assign new_n10820 = new_n10819 ^ new_n10816;
  assign new_n10821 = new_n5597 ^ n44;
  assign new_n10822 = new_n10821 ^ new_n4725;
  assign new_n10823 = new_n10822 ^ new_n4786;
  assign new_n10824 = new_n4595 ^ new_n2929;
  assign new_n10825 = new_n10824 ^ new_n10823;
  assign new_n10826 = new_n10825 ^ new_n10820;
  assign new_n10827 = new_n4757 ^ new_n4745;
  assign new_n10828 = new_n10827 ^ new_n4769;
  assign new_n10829 = new_n5684 ^ n46;
  assign new_n10830 = new_n10829 ^ new_n4696;
  assign new_n10831 = new_n10830 ^ new_n10828;
  assign new_n10832 = new_n5609 ^ n41;
  assign new_n10833 = new_n10832 ^ new_n4627;
  assign new_n10834 = new_n4721 ^ new_n4513;
  assign new_n10835 = new_n10834 ^ new_n10833;
  assign new_n10836 = new_n10835 ^ new_n10831;
  assign new_n10837 = new_n10836 ^ new_n10826;
  assign new_n10838 = new_n4725 ^ new_n4714;
  assign new_n10839 = new_n10838 ^ new_n4683;
  assign new_n10840 = new_n5641 ^ n47;
  assign new_n10841 = new_n10840 ^ new_n4762;
  assign new_n10842 = new_n10841 ^ new_n4691;
  assign new_n10843 = new_n10842 ^ new_n10839;
  assign new_n10844 = new_n10843 ^ new_n10820;
  assign new_n10845 = new_n4653 ^ new_n4574;
  assign new_n10846 = new_n4901 ^ n42;
  assign new_n10847 = new_n10846 ^ new_n4736;
  assign new_n10848 = new_n10847 ^ new_n4622;
  assign new_n10849 = new_n10848 ^ new_n10845;
  assign new_n10850 = new_n10849 ^ new_n10820;
  assign new_n10851 = new_n4725 ^ new_n4669;
  assign new_n10852 = new_n5544 ^ n48;
  assign new_n10853 = new_n10852 ^ new_n4709;
  assign new_n10854 = new_n10853 ^ new_n4676;
  assign new_n10855 = new_n10854 ^ new_n10851;
  assign new_n10856 = new_n10855 ^ new_n10850;
  assign new_n10857 = new_n10856 ^ new_n10843;
  assign new_n10858 = new_n10857 ^ new_n10836;
  assign new_n10859 = new_n4781 ^ new_n4526;
  assign new_n10860 = new_n10859 ^ new_n4535;
  assign new_n10861 = new_n5650 ^ n45;
  assign new_n10862 = new_n10861 ^ new_n4725;
  assign new_n10863 = new_n10862 ^ new_n4746;
  assign new_n10864 = new_n10863 ^ new_n10860;
  assign new_n10865 = new_n10864 ^ new_n10843;
  assign new_n10866 = new_n10835 ^ new_n10825;
  assign new_n10867 = new_n10866 ^ new_n10865;
  assign new_n10868 = new_n10867 ^ new_n10855;
  assign new_n10869 = new_n10858 & new_n10868;
  assign new_n10870 = new_n10843 & new_n10856;
  assign new_n10871 = new_n10870 ^ new_n10843;
  assign new_n10872 = new_n10871 ^ new_n10869;
  assign new_n10873 = new_n10865 ^ new_n10831;
  assign new_n10874 = new_n10873 ^ new_n10849;
  assign new_n10875 = new_n10866 & new_n10874;
  assign new_n10876 = new_n10867 ^ new_n10850;
  assign new_n10877 = ~new_n10876 & new_n10836;
  assign new_n10878 = new_n10877 ^ new_n10875;
  assign new_n10879 = new_n10873 ^ new_n10820;
  assign new_n10880 = new_n10879 ^ new_n10878;
  assign new_n10881 = new_n10843 ^ new_n10835;
  assign new_n10882 = ~new_n10881 & new_n10879;
  assign new_n10883 = new_n10874 ^ new_n10855;
  assign new_n10884 = new_n10856 ^ new_n10835;
  assign new_n10885 = ~new_n10883 & ~new_n10884;
  assign new_n10886 = new_n10885 ^ new_n10882;
  assign new_n10887 = new_n10886 ^ new_n10835;
  assign new_n10888 = new_n10887 ^ new_n10880;
  assign new_n10889 = new_n10856 ^ new_n10825;
  assign new_n10890 = ~new_n10855 & ~new_n10889;
  assign new_n10891 = new_n10890 ^ new_n10825;
  assign new_n10892 = new_n10831 ^ new_n10825;
  assign new_n10893 = new_n10892 ^ new_n10881;
  assign new_n10894 = ~new_n10867 & ~new_n10893;
  assign new_n10895 = new_n10894 ^ new_n10849;
  assign new_n10896 = new_n10895 ^ new_n10891;
  assign new_n10897 = new_n10882 ^ new_n10871;
  assign new_n10898 = new_n10897 ^ new_n10836;
  assign new_n10899 = ~new_n10837 & new_n10892;
  assign new_n10900 = new_n10899 ^ new_n10875;
  assign new_n10901 = new_n10864 ^ new_n10820;
  assign new_n10902 = new_n10901 ^ new_n10900;
  assign new_n10903 = new_n10902 ^ new_n10898;
  assign new_n10904 = new_n10895 ^ new_n10867;
  assign new_n10905 = new_n10900 ^ new_n10869;
  assign new_n10906 = new_n10905 ^ new_n10831;
  assign new_n10907 = new_n10906 ^ new_n10904;
  assign new_n10908 = ~new_n10903 & new_n10907;
  assign new_n10909 = new_n10908 ^ new_n10896;
  assign new_n10910 = new_n10909 ^ new_n10880;
  assign new_n10911 = new_n10899 ^ new_n10877;
  assign new_n10912 = new_n10885 ^ new_n10870;
  assign new_n10913 = new_n10912 ^ new_n10911;
  assign new_n10914 = ~new_n10910 & ~new_n10913;
  assign new_n10915 = new_n10914 ^ new_n10908;
  assign new_n10916 = ~new_n10888 & ~new_n10915;
  assign new_n10917 = new_n10916 ^ new_n10914;
  assign new_n10918 = new_n10908 ^ new_n10888;
  assign new_n10919 = new_n10835 ^ new_n10820;
  assign new_n10920 = new_n10890 ^ new_n10869;
  assign new_n10921 = new_n10920 ^ new_n10911;
  assign new_n10922 = new_n10921 ^ new_n10919;
  assign new_n10923 = ~new_n10922 & new_n10918;
  assign new_n10924 = new_n10923 ^ new_n10896;
  assign new_n10925 = new_n10924 ^ new_n10880;
  assign new_n10926 = ~new_n10917 & ~new_n10925;
  assign new_n10927 = new_n10918 ^ new_n10917;
  assign new_n10928 = new_n10927 ^ new_n10926;
  assign new_n10929 = new_n10928 ^ new_n10872;
  assign new_n10930 = new_n10929 ^ new_n10844;
  assign new_n10931 = new_n10930 ^ new_n10825;
  assign new_n10932 = new_n10923 ^ new_n10882;
  assign new_n10933 = new_n10932 ^ new_n10895;
  assign new_n10934 = new_n10933 ^ new_n10931;
  assign new_n10935 = ~new_n10837 & new_n10934;
  assign new_n10936 = new_n10923 ^ new_n10914;
  assign new_n10937 = new_n10896 ^ new_n10887;
  assign new_n10938 = new_n10937 ^ new_n10936;
  assign new_n10939 = ~new_n10938 & new_n10874;
  assign new_n10940 = new_n10939 ^ new_n10935;
  assign new_n10941 = new_n10892 & new_n10934;
  assign new_n10942 = ~new_n10938 & new_n10866;
  assign new_n10943 = new_n10942 ^ new_n10941;
  assign new_n10944 = new_n10927 ^ new_n10914;
  assign new_n10945 = new_n10944 ^ new_n10913;
  assign new_n10946 = new_n10858 & new_n10945;
  assign new_n10947 = new_n10946 ^ new_n10943;
  assign new_n10948 = new_n10927 ^ new_n10903;
  assign new_n10949 = ~new_n10893 & new_n10948;
  assign new_n10950 = new_n10868 & new_n10945;
  assign new_n10951 = ~new_n10867 & new_n10948;
  assign new_n10952 = new_n10951 ^ new_n10950;
  assign new_n10953 = new_n10952 ^ new_n10949;
  assign new_n10954 = new_n10953 ^ new_n10947;
  assign new_n10955 = new_n10954 ^ new_n10940;
  assign new_n10956 = new_n10955 ^ new_n10815;
  assign new_n10957 = new_n10956 ^ new_n10586;
  assign new_n10958 = ~new_n10361 & ~new_n10568;
  assign new_n10959 = new_n10403 ^ new_n10359;
  assign new_n10960 = ~new_n10959 & new_n10333;
  assign new_n10961 = new_n10960 ^ new_n10424;
  assign new_n10962 = new_n10961 ^ new_n10958;
  assign new_n10963 = new_n10962 ^ new_n10430;
  assign new_n10964 = new_n10540 ^ new_n10523;
  assign new_n10965 = new_n10483 & new_n10964;
  assign new_n10966 = new_n10538 ^ new_n10518;
  assign new_n10967 = new_n10966 ^ new_n10517;
  assign new_n10968 = ~new_n10967 & new_n10500;
  assign new_n10969 = new_n10555 ^ new_n10456;
  assign new_n10970 = new_n10528 ^ new_n10482;
  assign new_n10971 = new_n10970 ^ new_n10467;
  assign new_n10972 = new_n10971 ^ new_n10969;
  assign new_n10973 = ~new_n10972 & new_n10491;
  assign new_n10974 = new_n10973 ^ new_n10533;
  assign new_n10975 = new_n10974 ^ new_n10968;
  assign new_n10976 = new_n10975 ^ new_n10965;
  assign new_n10977 = new_n10480 & new_n10542;
  assign new_n10978 = new_n10977 ^ new_n10976;
  assign new_n10979 = ~new_n10546 & new_n10465;
  assign new_n10980 = ~new_n10967 & new_n10498;
  assign new_n10981 = new_n10980 ^ new_n10547;
  assign new_n10982 = new_n10981 ^ new_n10979;
  assign new_n10983 = new_n10982 ^ new_n10978;
  assign new_n10984 = new_n10983 ^ new_n10963;
  assign new_n10985 = new_n10984 ^ new_n10584;
  assign new_n10986 = new_n10681 ^ new_n10653;
  assign new_n10987 = ~new_n10629 & new_n10660;
  assign new_n10988 = new_n10649 ^ new_n8572;
  assign new_n10989 = new_n10637 ^ new_n10630;
  assign new_n10990 = new_n10989 ^ new_n10665;
  assign new_n10991 = new_n10990 ^ new_n10988;
  assign new_n10992 = new_n10624 & new_n10991;
  assign new_n10993 = new_n10992 ^ new_n10987;
  assign new_n10994 = new_n10649 ^ new_n10633;
  assign new_n10995 = ~new_n8553 & ~new_n10994;
  assign new_n10996 = new_n10995 ^ new_n10673;
  assign new_n10997 = new_n10661 ^ new_n10642;
  assign new_n10998 = new_n10997 ^ new_n10622;
  assign new_n10999 = ~new_n10998 & new_n10595;
  assign new_n11000 = new_n10999 ^ new_n10996;
  assign new_n11001 = new_n11000 ^ new_n10993;
  assign new_n11002 = new_n10598 & new_n10991;
  assign new_n11003 = new_n11002 ^ new_n11001;
  assign new_n11004 = new_n11003 ^ new_n10986;
  assign new_n11005 = new_n11004 ^ new_n8364;
  assign new_n11006 = new_n10801 ^ new_n10781;
  assign new_n11007 = new_n10777 ^ new_n10718;
  assign new_n11008 = new_n10765 ^ new_n10758;
  assign new_n11009 = new_n11008 ^ new_n10793;
  assign new_n11010 = new_n11009 ^ new_n11007;
  assign new_n11011 = new_n10722 & new_n11010;
  assign new_n11012 = new_n10757 & new_n10788;
  assign new_n11013 = new_n10752 & new_n11010;
  assign new_n11014 = new_n11013 ^ new_n11012;
  assign new_n11015 = new_n10777 ^ new_n10761;
  assign new_n11016 = new_n10711 & new_n11015;
  assign new_n11017 = new_n11016 ^ new_n10810;
  assign new_n11018 = new_n10789 ^ new_n10770;
  assign new_n11019 = new_n11018 ^ new_n10750;
  assign new_n11020 = new_n10719 & new_n11019;
  assign new_n11021 = new_n11020 ^ new_n11017;
  assign new_n11022 = new_n11021 ^ new_n11014;
  assign new_n11023 = new_n11022 ^ new_n11011;
  assign new_n11024 = new_n11023 ^ new_n11006;
  assign new_n11025 = new_n11024 ^ new_n11005;
  assign new_n11026 = new_n10942 ^ new_n10939;
  assign new_n11027 = new_n10914 ^ new_n10835;
  assign new_n11028 = new_n10890 ^ new_n10885;
  assign new_n11029 = new_n11028 ^ new_n10930;
  assign new_n11030 = new_n11029 ^ new_n11027;
  assign new_n11031 = ~new_n10876 & ~new_n11030;
  assign new_n11032 = ~new_n10884 & ~new_n10925;
  assign new_n11033 = new_n11032 ^ new_n11031;
  assign new_n11034 = new_n10926 ^ new_n10923;
  assign new_n11035 = new_n11034 ^ new_n10907;
  assign new_n11036 = ~new_n10881 & new_n11035;
  assign new_n11037 = new_n10914 ^ new_n10888;
  assign new_n11038 = ~new_n10855 & new_n11037;
  assign new_n11039 = new_n11038 ^ new_n10951;
  assign new_n11040 = new_n11039 ^ new_n11036;
  assign new_n11041 = new_n11040 ^ new_n11033;
  assign new_n11042 = ~new_n11030 & new_n10836;
  assign new_n11043 = new_n11042 ^ new_n11041;
  assign new_n11044 = new_n11043 ^ new_n11026;
  assign new_n11045 = new_n11044 ^ new_n11025;
  assign new_n11046 = new_n11045 ^ new_n10985;
  assign new_n11047 = new_n11046 ^ new_n10957;
  assign new_n11048 = ~new_n10594 & ~new_n10998;
  assign new_n11049 = new_n11048 ^ new_n11000;
  assign new_n11050 = new_n10661 ^ new_n10641;
  assign new_n11051 = ~new_n10616 & ~new_n11050;
  assign new_n11052 = new_n10628 & new_n10660;
  assign new_n11053 = new_n11052 ^ new_n11051;
  assign new_n11054 = new_n11053 ^ new_n10682;
  assign new_n11055 = new_n11054 ^ new_n11049;
  assign new_n11056 = new_n11055 ^ new_n8370;
  assign new_n11057 = new_n10958 ^ new_n10573;
  assign new_n11058 = ~new_n10959 & new_n10334;
  assign new_n11059 = ~new_n10383 & new_n10394;
  assign new_n11060 = new_n11059 ^ new_n11058;
  assign new_n11061 = new_n11060 ^ new_n10420;
  assign new_n11062 = new_n11061 ^ new_n11057;
  assign new_n11063 = new_n11062 ^ new_n11056;
  assign new_n11064 = new_n10879 & new_n11035;
  assign new_n11065 = new_n11064 ^ new_n11040;
  assign new_n11066 = new_n10926 ^ new_n10922;
  assign new_n11067 = ~new_n11066 & new_n10857;
  assign new_n11068 = ~new_n10883 & ~new_n10925;
  assign new_n11069 = new_n11068 ^ new_n11067;
  assign new_n11070 = new_n11069 ^ new_n10943;
  assign new_n11071 = new_n11070 ^ new_n11065;
  assign new_n11072 = new_n10715 & new_n11019;
  assign new_n11073 = new_n11072 ^ new_n11021;
  assign new_n11074 = new_n10789 ^ new_n10769;
  assign new_n11075 = new_n10745 & new_n11074;
  assign new_n11076 = new_n10756 & new_n10788;
  assign new_n11077 = new_n11076 ^ new_n11075;
  assign new_n11078 = new_n11077 ^ new_n10802;
  assign new_n11079 = new_n11078 ^ new_n11073;
  assign new_n11080 = new_n11079 ^ new_n11071;
  assign new_n11081 = new_n10979 ^ new_n10532;
  assign new_n11082 = ~new_n10972 & new_n10490;
  assign new_n11083 = new_n11082 ^ new_n10978;
  assign new_n11084 = new_n11083 ^ new_n11081;
  assign new_n11085 = new_n10426 ^ new_n10416;
  assign new_n11086 = new_n10962 ^ new_n10412;
  assign new_n11087 = new_n11086 ^ new_n11085;
  assign new_n11088 = new_n11087 ^ new_n11084;
  assign new_n11089 = new_n11088 ^ new_n11080;
  assign new_n11090 = new_n11089 ^ new_n11063;
  assign new_n11091 = new_n11090 ^ new_n11047;
  assign new_n11092 = ~new_n10591 & ~new_n11050;
  assign new_n11093 = new_n11092 ^ new_n10684;
  assign new_n11094 = new_n11093 ^ new_n11048;
  assign new_n11095 = new_n11094 ^ new_n10679;
  assign new_n11096 = new_n11095 ^ new_n8379;
  assign new_n11097 = new_n11096 ^ new_n11088;
  assign new_n11098 = new_n11059 ^ new_n10426;
  assign new_n11099 = new_n10571 ^ new_n10427;
  assign new_n11100 = new_n11099 ^ new_n10961;
  assign new_n11101 = new_n11100 ^ new_n11098;
  assign new_n11102 = new_n10513 & new_n10536;
  assign new_n11103 = new_n11102 ^ new_n10979;
  assign new_n11104 = new_n10980 ^ new_n10545;
  assign new_n11105 = new_n11104 ^ new_n10976;
  assign new_n11106 = new_n11105 ^ new_n11103;
  assign new_n11107 = new_n11106 ^ new_n11101;
  assign new_n11108 = new_n11107 ^ new_n11097;
  assign new_n11109 = new_n10712 & new_n11074;
  assign new_n11110 = new_n11109 ^ new_n10806;
  assign new_n11111 = new_n11110 ^ new_n11072;
  assign new_n11112 = new_n11111 ^ new_n10812;
  assign new_n11113 = new_n11112 ^ new_n10963;
  assign new_n11114 = ~new_n10856 & ~new_n11066;
  assign new_n11115 = new_n11114 ^ new_n10947;
  assign new_n11116 = new_n11115 ^ new_n11064;
  assign new_n11117 = new_n11116 ^ new_n10953;
  assign new_n11118 = new_n11117 ^ new_n11113;
  assign new_n11119 = new_n11118 ^ new_n11108;
  assign new_n11120 = new_n11119 ^ new_n11091;
  assign new_n11121 = new_n11090 & new_n11120;
  assign new_n11122 = new_n11121 ^ new_n11119;
  assign new_n11123 = new_n10578 ^ new_n10569;
  assign new_n11124 = new_n10960 ^ new_n10412;
  assign new_n11125 = new_n11124 ^ new_n11061;
  assign new_n11126 = new_n11125 ^ new_n11123;
  assign new_n11127 = new_n11020 ^ new_n11013;
  assign new_n11128 = new_n11109 ^ new_n10798;
  assign new_n11129 = new_n11128 ^ new_n11078;
  assign new_n11130 = new_n11129 ^ new_n11127;
  assign new_n11131 = new_n11130 ^ new_n11126;
  assign new_n11132 = new_n11131 ^ new_n11062;
  assign new_n11133 = new_n11132 ^ new_n11088;
  assign new_n11134 = new_n10999 ^ new_n10992;
  assign new_n11135 = new_n11092 ^ new_n10670;
  assign new_n11136 = new_n11135 ^ new_n11054;
  assign new_n11137 = new_n11136 ^ new_n11134;
  assign new_n11138 = new_n11137 ^ new_n8393;
  assign new_n11139 = new_n10977 ^ new_n10549;
  assign new_n11140 = new_n10499 & new_n10964;
  assign new_n11141 = new_n11140 ^ new_n11102;
  assign new_n11142 = new_n11141 ^ new_n10974;
  assign new_n11143 = new_n11142 ^ new_n11139;
  assign new_n11144 = new_n11143 ^ new_n11138;
  assign new_n11145 = new_n11036 ^ new_n11031;
  assign new_n11146 = new_n11114 ^ new_n10935;
  assign new_n11147 = new_n11146 ^ new_n11070;
  assign new_n11148 = new_n11147 ^ new_n11145;
  assign new_n11149 = new_n11148 ^ new_n11144;
  assign new_n11150 = new_n11149 ^ new_n11133;
  assign new_n11151 = new_n11068 ^ new_n10949;
  assign new_n11152 = new_n11038 ^ new_n10950;
  assign new_n11153 = new_n11152 ^ new_n11115;
  assign new_n11154 = new_n11153 ^ new_n11151;
  assign new_n11155 = new_n11154 ^ new_n11101;
  assign new_n11156 = new_n11076 ^ new_n10808;
  assign new_n11157 = new_n11016 ^ new_n10809;
  assign new_n11158 = new_n11157 ^ new_n11110;
  assign new_n11159 = new_n11158 ^ new_n11156;
  assign new_n11160 = new_n11159 ^ new_n11155;
  assign new_n11161 = new_n11052 ^ new_n10678;
  assign new_n11162 = new_n10995 ^ new_n10676;
  assign new_n11163 = new_n11162 ^ new_n11093;
  assign new_n11164 = new_n11163 ^ new_n11161;
  assign new_n11165 = new_n11164 ^ new_n8401;
  assign new_n11166 = new_n11165 ^ new_n11088;
  assign new_n11167 = ~new_n10570 & new_n10350;
  assign new_n11168 = new_n11167 ^ new_n11086;
  assign new_n11169 = new_n11168 ^ new_n10581;
  assign new_n11170 = new_n10483 ^ new_n10456;
  assign new_n11171 = new_n10544 & new_n11170;
  assign new_n11172 = new_n11171 ^ new_n11083;
  assign new_n11173 = new_n11172 ^ new_n10562;
  assign new_n11174 = new_n11173 ^ new_n11169;
  assign new_n11175 = new_n11174 ^ new_n11166;
  assign new_n11176 = new_n11175 ^ new_n11160;
  assign new_n11177 = new_n11176 ^ new_n11150;
  assign new_n11178 = new_n10678 ^ new_n10653;
  assign new_n11179 = new_n11094 ^ new_n10670;
  assign new_n11180 = new_n11179 ^ new_n11178;
  assign new_n11181 = new_n11180 ^ new_n8410;
  assign new_n11182 = new_n11082 ^ new_n10532;
  assign new_n11183 = new_n10982 ^ new_n10975;
  assign new_n11184 = new_n11183 ^ new_n11182;
  assign new_n11185 = new_n11184 ^ new_n10432;
  assign new_n11186 = new_n11185 ^ new_n11181;
  assign new_n11187 = new_n10808 ^ new_n10781;
  assign new_n11188 = new_n11111 ^ new_n10798;
  assign new_n11189 = new_n11188 ^ new_n11187;
  assign new_n11190 = new_n11189 ^ new_n11087;
  assign new_n11191 = new_n10949 ^ new_n10939;
  assign new_n11192 = new_n11116 ^ new_n10935;
  assign new_n11193 = new_n11192 ^ new_n11191;
  assign new_n11194 = new_n11193 ^ new_n11190;
  assign new_n11195 = new_n11194 ^ new_n11186;
  assign new_n11196 = new_n11195 ^ new_n11119;
  assign new_n11197 = new_n11196 ^ new_n11177;
  assign new_n11198 = new_n11195 ^ new_n11150;
  assign new_n11199 = ~new_n10889 & new_n11037;
  assign new_n11200 = new_n11199 ^ new_n11192;
  assign new_n11201 = new_n11200 ^ new_n11041;
  assign new_n11202 = new_n11201 ^ new_n11169;
  assign new_n11203 = new_n10764 & new_n11015;
  assign new_n11204 = new_n11203 ^ new_n11188;
  assign new_n11205 = new_n11204 ^ new_n11022;
  assign new_n11206 = new_n11205 ^ new_n11202;
  assign new_n11207 = ~new_n10636 & ~new_n10994;
  assign new_n11208 = new_n11207 ^ new_n11179;
  assign new_n11209 = new_n11208 ^ new_n11001;
  assign new_n11210 = new_n11209 ^ new_n8420;
  assign new_n11211 = new_n10559 ^ new_n10543;
  assign new_n11212 = new_n11082 ^ new_n10965;
  assign new_n11213 = new_n11212 ^ new_n11142;
  assign new_n11214 = new_n11213 ^ new_n11211;
  assign new_n11215 = new_n11214 ^ new_n11126;
  assign new_n11216 = new_n11215 ^ new_n11210;
  assign new_n11217 = new_n11216 ^ new_n11206;
  assign new_n11218 = new_n11217 ^ new_n11119;
  assign new_n11219 = new_n11218 ^ new_n11198;
  assign new_n11220 = new_n11197 & new_n11219;
  assign new_n11221 = new_n11220 ^ new_n10957;
  assign new_n11222 = new_n11221 ^ new_n11122;
  assign new_n11223 = new_n11195 ^ new_n11046;
  assign new_n11224 = new_n11217 ^ new_n11195;
  assign new_n11225 = new_n11197 ^ new_n11047;
  assign new_n11226 = new_n11224 & new_n11225;
  assign new_n11227 = new_n11119 ^ new_n11046;
  assign new_n11228 = new_n11227 ^ new_n11224;
  assign new_n11229 = new_n11218 & new_n11228;
  assign new_n11230 = new_n11229 ^ new_n11226;
  assign new_n11231 = new_n11197 ^ new_n11090;
  assign new_n11232 = new_n11150 ^ new_n11091;
  assign new_n11233 = new_n11232 ^ new_n11224;
  assign new_n11234 = new_n11231 & new_n11233;
  assign new_n11235 = new_n11234 ^ new_n11121;
  assign new_n11236 = new_n11235 ^ new_n11230;
  assign new_n11237 = new_n11236 ^ new_n11223;
  assign new_n11238 = new_n11195 ^ new_n11091;
  assign new_n11239 = new_n11217 ^ new_n11177;
  assign new_n11240 = new_n11239 ^ new_n10957;
  assign new_n11241 = new_n11240 ^ new_n11090;
  assign new_n11242 = new_n11238 & new_n11241;
  assign new_n11243 = new_n11239 ^ new_n11046;
  assign new_n11244 = new_n11198 & new_n11243;
  assign new_n11245 = new_n11244 ^ new_n11242;
  assign new_n11246 = new_n11245 ^ new_n11195;
  assign new_n11247 = new_n11196 & new_n11240;
  assign new_n11248 = new_n11247 ^ new_n11226;
  assign new_n11249 = new_n11248 ^ new_n11243;
  assign new_n11250 = new_n11249 ^ new_n11246;
  assign new_n11251 = ~new_n11091 & ~new_n11150;
  assign new_n11252 = new_n11251 ^ new_n11150;
  assign new_n11253 = new_n11252 ^ new_n11244;
  assign new_n11254 = new_n11253 ^ new_n11224;
  assign new_n11255 = new_n11247 ^ new_n11229;
  assign new_n11256 = new_n11176 ^ new_n11046;
  assign new_n11257 = new_n11256 ^ new_n11255;
  assign new_n11258 = new_n11257 ^ new_n11254;
  assign new_n11259 = new_n11221 ^ new_n11197;
  assign new_n11260 = new_n11255 ^ new_n11234;
  assign new_n11261 = new_n11260 ^ new_n11217;
  assign new_n11262 = new_n11261 ^ new_n11259;
  assign new_n11263 = ~new_n11258 & new_n11262;
  assign new_n11264 = new_n11263 ^ new_n11250;
  assign new_n11265 = new_n11237 & new_n11264;
  assign new_n11266 = new_n11265 ^ new_n11222;
  assign new_n11267 = new_n11266 ^ new_n11249;
  assign new_n11268 = new_n11263 ^ new_n11222;
  assign new_n11269 = new_n11268 ^ new_n11249;
  assign new_n11270 = new_n11251 ^ new_n11242;
  assign new_n11271 = new_n11270 ^ new_n11230;
  assign new_n11272 = ~new_n11271 & new_n11269;
  assign new_n11273 = new_n11272 ^ new_n11263;
  assign new_n11274 = ~new_n11273 & new_n11250;
  assign new_n11275 = new_n11274 ^ new_n11263;
  assign new_n11276 = new_n11267 & new_n11275;
  assign new_n11277 = new_n11276 ^ new_n11237;
  assign new_n11278 = new_n11091 & new_n11277;
  assign new_n11279 = new_n11274 ^ new_n11250;
  assign new_n11280 = new_n11279 ^ new_n11272;
  assign new_n11281 = new_n11280 ^ new_n11271;
  assign new_n11282 = ~new_n11281 & new_n11233;
  assign new_n11283 = new_n11272 ^ new_n11265;
  assign new_n11284 = new_n11246 ^ new_n11222;
  assign new_n11285 = new_n11284 ^ new_n11283;
  assign new_n11286 = new_n11196 & new_n11285;
  assign new_n11287 = new_n11150 ^ new_n11046;
  assign new_n11288 = new_n11252 ^ new_n11234;
  assign new_n11289 = new_n11279 ^ new_n11276;
  assign new_n11290 = new_n11289 ^ new_n11288;
  assign new_n11291 = new_n11290 ^ new_n11287;
  assign new_n11292 = new_n11291 ^ new_n11119;
  assign new_n11293 = new_n11265 ^ new_n11244;
  assign new_n11294 = new_n11293 ^ new_n11221;
  assign new_n11295 = new_n11294 ^ new_n11292;
  assign new_n11296 = ~new_n11295 & new_n11218;
  assign new_n11297 = new_n11296 ^ new_n11286;
  assign new_n11298 = new_n11297 ^ new_n11282;
  assign new_n11299 = new_n11298 ^ new_n11278;
  assign new_n11300 = new_n11276 ^ new_n11265;
  assign new_n11301 = new_n11300 ^ new_n11262;
  assign new_n11302 = new_n11243 & new_n11301;
  assign new_n11303 = new_n11302 ^ new_n11299;
  assign new_n11304 = new_n11279 ^ new_n11258;
  assign new_n11305 = ~new_n11304 & new_n11197;
  assign new_n11306 = ~new_n11281 & new_n11231;
  assign new_n11307 = new_n11306 ^ new_n11305;
  assign new_n11308 = ~new_n11304 & new_n11219;
  assign new_n11309 = new_n11308 ^ new_n11307;
  assign new_n11310 = new_n11309 ^ new_n11303;
  assign new_n11311 = new_n10158 ^ new_n10135;
  assign new_n11312 = new_n11311 ^ new_n10134;
  assign new_n11313 = ~new_n10115 & ~new_n11312;
  assign new_n11314 = new_n11313 ^ new_n10173;
  assign new_n11315 = new_n10094 & new_n10172;
  assign new_n11316 = new_n11315 ^ new_n11314;
  assign new_n11317 = ~new_n11312 & new_n10117;
  assign new_n11318 = new_n10163 ^ new_n10071;
  assign new_n11319 = new_n10144 ^ new_n10100;
  assign new_n11320 = new_n11319 ^ new_n10096;
  assign new_n11321 = new_n11320 ^ new_n11318;
  assign new_n11322 = ~new_n10108 & ~new_n11321;
  assign new_n11323 = new_n11322 ^ new_n10149;
  assign new_n11324 = new_n11323 ^ new_n11317;
  assign new_n11325 = new_n10160 ^ new_n10139;
  assign new_n11326 = ~new_n11325 & new_n10057;
  assign new_n11327 = new_n11326 ^ new_n11324;
  assign new_n11328 = ~new_n10098 & ~new_n10176;
  assign new_n11329 = new_n11328 ^ new_n11327;
  assign new_n11330 = new_n11329 ^ new_n11316;
  assign new_n11331 = new_n11330 ^ new_n11310;
  assign new_n11332 = new_n11331 ^ new_n10300;
  assign new_n11333 = new_n11332 ^ new_n10182;
  assign new_n11334 = new_n9143 ^ new_n9073;
  assign new_n11335 = new_n9123 ^ new_n9055;
  assign new_n11336 = new_n11335 ^ new_n9088;
  assign new_n11337 = new_n11336 ^ new_n11334;
  assign new_n11338 = ~new_n11337 & new_n9077;
  assign new_n11339 = new_n11338 ^ new_n9127;
  assign new_n11340 = new_n9136 ^ new_n9114;
  assign new_n11341 = new_n11340 ^ new_n9113;
  assign new_n11342 = ~new_n11341 & new_n9090;
  assign new_n11343 = new_n11342 ^ new_n9151;
  assign new_n11344 = ~new_n9150 & new_n9086;
  assign new_n11345 = new_n11344 ^ new_n11343;
  assign new_n11346 = ~new_n11337 & new_n9078;
  assign new_n11347 = new_n11346 ^ new_n9128;
  assign new_n11348 = ~new_n11341 & new_n9092;
  assign new_n11349 = new_n11348 ^ new_n11347;
  assign new_n11350 = new_n11349 ^ new_n11345;
  assign new_n11351 = new_n11350 ^ new_n11339;
  assign new_n11352 = new_n8042 ^ new_n7971;
  assign new_n11353 = new_n8022 ^ new_n7953;
  assign new_n11354 = new_n11353 ^ new_n7986;
  assign new_n11355 = new_n11354 ^ new_n11352;
  assign new_n11356 = ~new_n7975 & ~new_n11355;
  assign new_n11357 = new_n11356 ^ new_n8026;
  assign new_n11358 = new_n8035 ^ new_n8013;
  assign new_n11359 = new_n11358 ^ new_n8012;
  assign new_n11360 = ~new_n11359 & new_n7988;
  assign new_n11361 = new_n11360 ^ new_n8050;
  assign new_n11362 = ~new_n7984 & ~new_n8049;
  assign new_n11363 = new_n11362 ^ new_n11361;
  assign new_n11364 = ~new_n11355 & new_n7976;
  assign new_n11365 = new_n11364 ^ new_n8027;
  assign new_n11366 = ~new_n11359 & new_n7990;
  assign new_n11367 = new_n11366 ^ new_n11365;
  assign new_n11368 = new_n11367 ^ new_n11363;
  assign new_n11369 = new_n11368 ^ new_n11357;
  assign new_n11370 = new_n11369 ^ new_n11351;
  assign new_n11371 = new_n11240 & new_n11285;
  assign new_n11372 = new_n11371 ^ new_n11286;
  assign new_n11373 = new_n11272 ^ new_n11195;
  assign new_n11374 = new_n11242 ^ new_n11121;
  assign new_n11375 = new_n11374 ^ new_n11291;
  assign new_n11376 = new_n11375 ^ new_n11373;
  assign new_n11377 = ~new_n11376 & new_n11224;
  assign new_n11378 = new_n11238 & new_n11267;
  assign new_n11379 = ~new_n11376 & new_n11225;
  assign new_n11380 = new_n11379 ^ new_n11378;
  assign new_n11381 = new_n11272 ^ new_n11250;
  assign new_n11382 = new_n11090 & new_n11381;
  assign new_n11383 = new_n11382 ^ new_n11305;
  assign new_n11384 = new_n11198 & new_n11301;
  assign new_n11385 = new_n11384 ^ new_n11383;
  assign new_n11386 = new_n11385 ^ new_n11380;
  assign new_n11387 = new_n11386 ^ new_n11377;
  assign new_n11388 = new_n11387 ^ new_n11372;
  assign new_n11389 = new_n11388 ^ new_n11370;
  assign new_n11390 = new_n10280 ^ new_n10186;
  assign new_n11391 = new_n10256 ^ new_n10228;
  assign new_n11392 = new_n11391 ^ new_n10240;
  assign new_n11393 = new_n11392 ^ new_n11390;
  assign new_n11394 = ~new_n11393 & new_n10216;
  assign new_n11395 = new_n11394 ^ new_n10267;
  assign new_n11396 = new_n10275 ^ new_n10262;
  assign new_n11397 = new_n11396 ^ new_n10261;
  assign new_n11398 = ~new_n11397 & new_n10211;
  assign new_n11399 = new_n11398 ^ new_n10291;
  assign new_n11400 = new_n10238 & new_n10290;
  assign new_n11401 = new_n11400 ^ new_n11399;
  assign new_n11402 = ~new_n10206 & ~new_n11397;
  assign new_n11403 = ~new_n10214 & ~new_n11393;
  assign new_n11404 = new_n11403 ^ new_n10266;
  assign new_n11405 = new_n11404 ^ new_n11402;
  assign new_n11406 = new_n11405 ^ new_n11401;
  assign new_n11407 = new_n11406 ^ new_n11395;
  assign new_n11408 = new_n11407 ^ new_n6575;
  assign new_n11409 = ~new_n11321 & new_n10107;
  assign new_n11410 = new_n11409 ^ new_n10148;
  assign new_n11411 = new_n11324 ^ new_n11316;
  assign new_n11412 = new_n11411 ^ new_n11410;
  assign new_n11413 = new_n11412 ^ new_n11408;
  assign new_n11414 = new_n11413 ^ new_n10181;
  assign new_n11415 = new_n11414 ^ new_n11389;
  assign new_n11416 = new_n11415 ^ new_n11333;
  assign new_n11417 = ~new_n10226 & ~new_n10294;
  assign new_n11418 = new_n11417 ^ new_n10296;
  assign new_n11419 = new_n10277 ^ new_n10222;
  assign new_n11420 = ~new_n11419 & new_n10202;
  assign new_n11421 = new_n10250 & new_n10273;
  assign new_n11422 = new_n11421 ^ new_n11420;
  assign new_n11423 = new_n11422 ^ new_n11404;
  assign new_n11424 = new_n11423 ^ new_n11418;
  assign new_n11425 = new_n11424 ^ new_n6630;
  assign new_n11426 = new_n11328 ^ new_n10178;
  assign new_n11427 = ~new_n10130 & new_n10156;
  assign new_n11428 = ~new_n10116 & ~new_n11325;
  assign new_n11429 = new_n11428 ^ new_n11427;
  assign new_n11430 = new_n11429 ^ new_n11323;
  assign new_n11431 = new_n11430 ^ new_n11426;
  assign new_n11432 = new_n11431 ^ new_n11425;
  assign new_n11433 = new_n9037 & new_n9156;
  assign new_n11434 = new_n11433 ^ new_n9158;
  assign new_n11435 = new_n9140 ^ new_n9118;
  assign new_n11436 = new_n9091 & new_n11435;
  assign new_n11437 = new_n9109 & new_n9138;
  assign new_n11438 = new_n11437 ^ new_n11436;
  assign new_n11439 = new_n11438 ^ new_n11347;
  assign new_n11440 = new_n11439 ^ new_n11434;
  assign new_n11441 = new_n7935 & new_n8055;
  assign new_n11442 = new_n11441 ^ new_n8057;
  assign new_n11443 = new_n8039 ^ new_n8017;
  assign new_n11444 = ~new_n11443 & new_n7989;
  assign new_n11445 = ~new_n8008 & ~new_n8037;
  assign new_n11446 = new_n11445 ^ new_n11444;
  assign new_n11447 = new_n11446 ^ new_n11365;
  assign new_n11448 = new_n11447 ^ new_n11442;
  assign new_n11449 = new_n11448 ^ new_n11440;
  assign new_n11450 = new_n11371 ^ new_n11308;
  assign new_n11451 = ~new_n11295 & new_n11228;
  assign new_n11452 = new_n11451 ^ new_n11303;
  assign new_n11453 = new_n11452 ^ new_n11450;
  assign new_n11454 = new_n11315 ^ new_n10148;
  assign new_n11455 = new_n11409 ^ new_n11329;
  assign new_n11456 = new_n11455 ^ new_n11454;
  assign new_n11457 = new_n11456 ^ new_n11453;
  assign new_n11458 = new_n11457 ^ new_n11449;
  assign new_n11459 = new_n11458 ^ new_n11432;
  assign new_n11460 = new_n11459 ^ new_n11416;
  assign new_n11461 = ~new_n10199 & ~new_n11419;
  assign new_n11462 = new_n11461 ^ new_n11405;
  assign new_n11463 = new_n11462 ^ new_n11417;
  assign new_n11464 = new_n11463 ^ new_n11401;
  assign new_n11465 = new_n11464 ^ new_n8237;
  assign new_n11466 = new_n9034 & new_n11435;
  assign new_n11467 = new_n11466 ^ new_n11349;
  assign new_n11468 = new_n11467 ^ new_n11433;
  assign new_n11469 = new_n11468 ^ new_n11345;
  assign new_n11470 = ~new_n7932 & ~new_n11443;
  assign new_n11471 = new_n11470 ^ new_n11367;
  assign new_n11472 = new_n11471 ^ new_n11441;
  assign new_n11473 = new_n11472 ^ new_n11363;
  assign new_n11474 = new_n11473 ^ new_n11469;
  assign new_n11475 = new_n11474 ^ new_n11465;
  assign new_n11476 = new_n11475 ^ new_n11457;
  assign new_n11477 = new_n11241 & new_n11267;
  assign new_n11478 = new_n11477 ^ new_n11308;
  assign new_n11479 = new_n11382 ^ new_n11306;
  assign new_n11480 = new_n11479 ^ new_n11299;
  assign new_n11481 = new_n11480 ^ new_n11478;
  assign new_n11482 = new_n11481 ^ new_n11330;
  assign new_n11483 = new_n11427 ^ new_n11315;
  assign new_n11484 = new_n11313 ^ new_n10171;
  assign new_n11485 = new_n11484 ^ new_n11327;
  assign new_n11486 = new_n11485 ^ new_n11483;
  assign new_n11487 = new_n11486 ^ new_n11482;
  assign new_n11488 = new_n11487 ^ new_n11476;
  assign new_n11489 = new_n11488 ^ new_n11460;
  assign new_n11490 = ~new_n11459 & ~new_n11489;
  assign new_n11491 = new_n11490 ^ new_n11488;
  assign new_n11492 = ~new_n10170 & new_n10072;
  assign new_n11493 = new_n11492 ^ new_n11455;
  assign new_n11494 = new_n11493 ^ new_n10179;
  assign new_n11495 = new_n11120 & new_n11381;
  assign new_n11496 = new_n11495 ^ new_n11452;
  assign new_n11497 = new_n11496 ^ new_n11386;
  assign new_n11498 = new_n11497 ^ new_n11486;
  assign new_n11499 = new_n11498 ^ new_n11494;
  assign new_n11500 = new_n11421 ^ new_n11400;
  assign new_n11501 = new_n11398 ^ new_n10289;
  assign new_n11502 = new_n11501 ^ new_n11462;
  assign new_n11503 = new_n11502 ^ new_n11500;
  assign new_n11504 = new_n11503 ^ new_n8234;
  assign new_n11505 = new_n11504 ^ new_n11457;
  assign new_n11506 = new_n11437 ^ new_n11344;
  assign new_n11507 = new_n11342 ^ new_n9153;
  assign new_n11508 = new_n11507 ^ new_n11467;
  assign new_n11509 = new_n11508 ^ new_n11506;
  assign new_n11510 = new_n11445 ^ new_n11362;
  assign new_n11511 = new_n11360 ^ new_n8052;
  assign new_n11512 = new_n11511 ^ new_n11471;
  assign new_n11513 = new_n11512 ^ new_n11510;
  assign new_n11514 = new_n11513 ^ new_n11509;
  assign new_n11515 = new_n11514 ^ new_n11505;
  assign new_n11516 = new_n11515 ^ new_n11499;
  assign new_n11517 = new_n11385 ^ new_n11302;
  assign new_n11518 = new_n11232 & new_n11277;
  assign new_n11519 = new_n11518 ^ new_n11477;
  assign new_n11520 = new_n11519 ^ new_n11297;
  assign new_n11521 = new_n11520 ^ new_n11517;
  assign new_n11522 = new_n11521 ^ new_n11457;
  assign new_n11523 = new_n9157 ^ new_n9148;
  assign new_n11524 = new_n11466 ^ new_n11338;
  assign new_n11525 = new_n11524 ^ new_n11439;
  assign new_n11526 = new_n11525 ^ new_n11523;
  assign new_n11527 = new_n8056 ^ new_n8047;
  assign new_n11528 = new_n11470 ^ new_n11356;
  assign new_n11529 = new_n11528 ^ new_n11447;
  assign new_n11530 = new_n11529 ^ new_n11527;
  assign new_n11531 = new_n11530 ^ new_n11526;
  assign new_n11532 = new_n11531 ^ new_n11522;
  assign new_n11533 = new_n10295 ^ new_n10286;
  assign new_n11534 = new_n11461 ^ new_n11394;
  assign new_n11535 = new_n11534 ^ new_n11423;
  assign new_n11536 = new_n11535 ^ new_n11533;
  assign new_n11537 = new_n11536 ^ new_n6660;
  assign new_n11538 = new_n10177 ^ new_n10168;
  assign new_n11539 = new_n11409 ^ new_n11326;
  assign new_n11540 = new_n11539 ^ new_n11430;
  assign new_n11541 = new_n11540 ^ new_n11538;
  assign new_n11542 = new_n11541 ^ new_n11537;
  assign new_n11543 = new_n11542 ^ new_n11431;
  assign new_n11544 = new_n11543 ^ new_n11532;
  assign new_n11545 = new_n11544 ^ new_n11516;
  assign new_n11546 = new_n11344 ^ new_n9127;
  assign new_n11547 = new_n11468 ^ new_n11338;
  assign new_n11548 = new_n11547 ^ new_n11546;
  assign new_n11549 = new_n11362 ^ new_n8026;
  assign new_n11550 = new_n11472 ^ new_n11356;
  assign new_n11551 = new_n11550 ^ new_n11549;
  assign new_n11552 = new_n11551 ^ new_n11548;
  assign new_n11553 = new_n11451 ^ new_n11371;
  assign new_n11554 = new_n11309 ^ new_n11298;
  assign new_n11555 = new_n11554 ^ new_n11553;
  assign new_n11556 = new_n11555 ^ new_n11552;
  assign new_n11557 = new_n11463 ^ new_n11394;
  assign new_n11558 = new_n11400 ^ new_n10267;
  assign new_n11559 = new_n11558 ^ new_n11557;
  assign new_n11560 = new_n11559 ^ new_n6680;
  assign new_n11561 = new_n11560 ^ new_n11456;
  assign new_n11562 = new_n11561 ^ new_n11412;
  assign new_n11563 = new_n11562 ^ new_n11556;
  assign new_n11564 = new_n11563 ^ new_n11488;
  assign new_n11565 = new_n11564 ^ new_n11545;
  assign new_n11566 = new_n9098 & new_n9152;
  assign new_n11567 = new_n11566 ^ new_n11547;
  assign new_n11568 = new_n11567 ^ new_n9159;
  assign new_n11569 = ~new_n7997 & new_n8051;
  assign new_n11570 = new_n11569 ^ new_n11550;
  assign new_n11571 = new_n11570 ^ new_n8058;
  assign new_n11572 = new_n11571 ^ new_n11568;
  assign new_n11573 = new_n11384 ^ new_n11379;
  assign new_n11574 = new_n11451 ^ new_n11278;
  assign new_n11575 = new_n11574 ^ new_n11520;
  assign new_n11576 = new_n11575 ^ new_n11573;
  assign new_n11577 = new_n11576 ^ new_n11572;
  assign new_n11578 = new_n10199 ^ new_n10186;
  assign new_n11579 = ~new_n10288 & ~new_n11578;
  assign new_n11580 = new_n11579 ^ new_n11557;
  assign new_n11581 = new_n11580 ^ new_n10297;
  assign new_n11582 = new_n11581 ^ new_n6726;
  assign new_n11583 = new_n11582 ^ new_n11494;
  assign new_n11584 = new_n11583 ^ new_n11541;
  assign new_n11585 = new_n11584 ^ new_n11577;
  assign new_n11586 = new_n11585 ^ new_n11488;
  assign new_n11587 = new_n11563 ^ new_n11544;
  assign new_n11588 = new_n11587 ^ new_n11586;
  assign new_n11589 = ~new_n11565 & ~new_n11588;
  assign new_n11590 = new_n11589 ^ new_n11415;
  assign new_n11591 = new_n11590 ^ new_n11491;
  assign new_n11592 = new_n11460 & new_n11544;
  assign new_n11593 = new_n11592 ^ new_n11544;
  assign new_n11594 = new_n11585 ^ new_n11545;
  assign new_n11595 = new_n11594 ^ new_n11333;
  assign new_n11596 = ~new_n11587 & new_n11595;
  assign new_n11597 = new_n11596 ^ new_n11593;
  assign new_n11598 = new_n11585 ^ new_n11563;
  assign new_n11599 = new_n11598 ^ new_n11597;
  assign new_n11600 = new_n11594 ^ new_n11415;
  assign new_n11601 = new_n11564 & new_n11600;
  assign new_n11602 = new_n11488 ^ new_n11333;
  assign new_n11603 = new_n11602 ^ new_n11598;
  assign new_n11604 = ~new_n11603 & new_n11586;
  assign new_n11605 = new_n11604 ^ new_n11601;
  assign new_n11606 = new_n11516 ^ new_n11333;
  assign new_n11607 = new_n11606 ^ new_n11605;
  assign new_n11608 = new_n11607 ^ new_n11599;
  assign new_n11609 = new_n11590 ^ new_n11565;
  assign new_n11610 = new_n11565 ^ new_n11459;
  assign new_n11611 = new_n11544 ^ new_n11460;
  assign new_n11612 = new_n11611 ^ new_n11598;
  assign new_n11613 = new_n11610 & new_n11612;
  assign new_n11614 = new_n11613 ^ new_n11605;
  assign new_n11615 = new_n11614 ^ new_n11585;
  assign new_n11616 = new_n11615 ^ new_n11609;
  assign new_n11617 = ~new_n11608 & new_n11616;
  assign new_n11618 = new_n11617 ^ new_n11591;
  assign new_n11619 = new_n11565 ^ new_n11416;
  assign new_n11620 = ~new_n11619 & new_n11598;
  assign new_n11621 = new_n11620 ^ new_n11601;
  assign new_n11622 = new_n11621 ^ new_n11595;
  assign new_n11623 = new_n11622 ^ new_n11618;
  assign new_n11624 = new_n11600 ^ new_n11459;
  assign new_n11625 = new_n11563 ^ new_n11460;
  assign new_n11626 = ~new_n11624 & ~new_n11625;
  assign new_n11627 = new_n11626 ^ new_n11592;
  assign new_n11628 = new_n11620 ^ new_n11604;
  assign new_n11629 = new_n11628 ^ new_n11627;
  assign new_n11630 = ~new_n11623 & ~new_n11629;
  assign new_n11631 = new_n11626 ^ new_n11596;
  assign new_n11632 = new_n11631 ^ new_n11563;
  assign new_n11633 = new_n11632 ^ new_n11622;
  assign new_n11634 = new_n11633 ^ new_n11630;
  assign new_n11635 = ~new_n11489 & new_n11634;
  assign new_n11636 = new_n11563 ^ new_n11333;
  assign new_n11637 = new_n11613 ^ new_n11490;
  assign new_n11638 = new_n11637 ^ new_n11628;
  assign new_n11639 = new_n11638 ^ new_n11636;
  assign new_n11640 = new_n11633 ^ new_n11617;
  assign new_n11641 = ~new_n11639 & new_n11640;
  assign new_n11642 = new_n11641 ^ new_n11591;
  assign new_n11643 = new_n11642 ^ new_n11622;
  assign new_n11644 = new_n11630 ^ new_n11617;
  assign new_n11645 = ~new_n11644 & new_n11633;
  assign new_n11646 = new_n11645 ^ new_n11617;
  assign new_n11647 = ~new_n11643 & new_n11646;
  assign new_n11648 = new_n11647 ^ new_n11639;
  assign new_n11649 = ~new_n11460 & ~new_n11648;
  assign new_n11650 = new_n11645 ^ new_n11633;
  assign new_n11651 = new_n11650 ^ new_n11630;
  assign new_n11652 = new_n11651 ^ new_n11629;
  assign new_n11653 = ~new_n11652 & new_n11612;
  assign new_n11654 = new_n11544 ^ new_n11333;
  assign new_n11655 = new_n11613 ^ new_n11593;
  assign new_n11656 = new_n11650 ^ new_n11647;
  assign new_n11657 = new_n11656 ^ new_n11655;
  assign new_n11658 = new_n11657 ^ new_n11654;
  assign new_n11659 = new_n11658 ^ new_n11488;
  assign new_n11660 = new_n11641 ^ new_n11596;
  assign new_n11661 = new_n11660 ^ new_n11590;
  assign new_n11662 = new_n11661 ^ new_n11659;
  assign new_n11663 = ~new_n11662 & new_n11586;
  assign new_n11664 = new_n11641 ^ new_n11630;
  assign new_n11665 = new_n11632 ^ new_n11591;
  assign new_n11666 = new_n11665 ^ new_n11664;
  assign new_n11667 = ~new_n11666 & new_n11564;
  assign new_n11668 = new_n11667 ^ new_n11663;
  assign new_n11669 = new_n11668 ^ new_n11653;
  assign new_n11670 = new_n11669 ^ new_n11649;
  assign new_n11671 = new_n11647 ^ new_n11641;
  assign new_n11672 = new_n11671 ^ new_n11616;
  assign new_n11673 = new_n11595 & new_n11672;
  assign new_n11674 = new_n11673 ^ new_n11670;
  assign new_n11675 = ~new_n11603 & ~new_n11662;
  assign new_n11676 = new_n11675 ^ new_n11674;
  assign new_n11677 = new_n11676 ^ new_n11635;
  assign new_n11678 = ~new_n11625 & ~new_n11643;
  assign new_n11679 = new_n11630 ^ new_n11563;
  assign new_n11680 = new_n11626 ^ new_n11490;
  assign new_n11681 = new_n11680 ^ new_n11658;
  assign new_n11682 = new_n11681 ^ new_n11679;
  assign new_n11683 = ~new_n11619 & new_n11682;
  assign new_n11684 = new_n11683 ^ new_n11678;
  assign new_n11685 = ~new_n11459 & new_n11634;
  assign new_n11686 = new_n11650 ^ new_n11608;
  assign new_n11687 = ~new_n11565 & ~new_n11686;
  assign new_n11688 = new_n11687 ^ new_n11685;
  assign new_n11689 = ~new_n11587 & new_n11672;
  assign new_n11690 = new_n11689 ^ new_n11688;
  assign new_n11691 = new_n11690 ^ new_n11684;
  assign new_n11692 = new_n11691 ^ new_n11677;
  assign new_n11693 = new_n11095 ^ n36;
  assign new_n11694 = new_n11693 ^ new_n8237;
  assign new_n11695 = new_n11694 ^ new_n7928;
  assign new_n11696 = new_n7944 ^ new_n7941;
  assign new_n11697 = new_n11696 ^ new_n11695;
  assign new_n11698 = new_n7968 ^ new_n7838;
  assign new_n11699 = new_n11698 ^ new_n7830;
  assign new_n11700 = new_n11699 ^ new_n11697;
  assign new_n11701 = new_n7881 ^ new_n7814;
  assign new_n11702 = new_n11180 ^ n33;
  assign new_n11703 = new_n11702 ^ new_n6680;
  assign new_n11704 = new_n11703 ^ new_n7941;
  assign new_n11705 = new_n11704 ^ new_n7869;
  assign new_n11706 = new_n11705 ^ new_n11701;
  assign new_n11707 = new_n11706 ^ new_n11700;
  assign new_n11708 = new_n11696 ^ new_n7903;
  assign new_n11709 = new_n11708 ^ new_n7755;
  assign new_n11710 = new_n11137 ^ n39;
  assign new_n11711 = new_n11710 ^ new_n6660;
  assign new_n11712 = new_n11711 ^ new_n7797;
  assign new_n11713 = new_n11712 ^ new_n7900;
  assign new_n11714 = new_n11713 ^ new_n11709;
  assign new_n11715 = new_n7830 ^ new_n6837;
  assign new_n11716 = new_n11715 ^ new_n4899;
  assign new_n11717 = new_n11164 ^ n37;
  assign new_n11718 = new_n11717 ^ new_n8234;
  assign new_n11719 = new_n11718 ^ new_n11696;
  assign new_n11720 = new_n11719 ^ new_n7963;
  assign new_n11721 = new_n11720 ^ new_n11716;
  assign new_n11722 = new_n11721 ^ new_n11714;
  assign new_n11723 = new_n11722 ^ new_n11707;
  assign new_n11724 = new_n7851 ^ new_n7765;
  assign new_n11725 = new_n11209 ^ n38;
  assign new_n11726 = new_n11725 ^ new_n6726;
  assign new_n11727 = new_n11726 ^ new_n4899;
  assign new_n11728 = new_n11727 ^ new_n7797;
  assign new_n11729 = new_n11728 ^ new_n11724;
  assign new_n11730 = new_n11729 ^ new_n11706;
  assign new_n11731 = new_n7916 ^ new_n7891;
  assign new_n11732 = new_n11004 ^ n35;
  assign new_n11733 = new_n11732 ^ new_n8226;
  assign new_n11734 = new_n7968 ^ new_n7957;
  assign new_n11735 = new_n11734 ^ new_n11733;
  assign new_n11736 = new_n11735 ^ new_n11731;
  assign new_n11737 = new_n7949 ^ new_n7921;
  assign new_n11738 = new_n10686 ^ n34;
  assign new_n11739 = new_n11738 ^ new_n6575;
  assign new_n11740 = new_n11739 ^ new_n7869;
  assign new_n11741 = new_n11740 ^ new_n7916;
  assign new_n11742 = new_n11741 ^ new_n11737;
  assign new_n11743 = new_n11742 ^ new_n11736;
  assign new_n11744 = new_n11743 ^ new_n11723;
  assign new_n11745 = ~new_n11744 & new_n11730;
  assign new_n11746 = new_n11729 ^ new_n11722;
  assign new_n11747 = new_n11746 ^ new_n11742;
  assign new_n11748 = new_n11707 & new_n11747;
  assign new_n11749 = new_n11748 ^ new_n11745;
  assign new_n11750 = new_n11746 ^ new_n11736;
  assign new_n11751 = new_n11750 ^ new_n11749;
  assign new_n11752 = new_n11714 ^ new_n11706;
  assign new_n11753 = ~new_n11752 & new_n11750;
  assign new_n11754 = new_n11055 ^ n40;
  assign new_n11755 = new_n11754 ^ new_n6630;
  assign new_n11756 = new_n11755 ^ new_n7900;
  assign new_n11757 = new_n11696 ^ new_n7778;
  assign new_n11758 = new_n11757 ^ new_n11756;
  assign new_n11759 = new_n11758 ^ new_n11743;
  assign new_n11760 = new_n11759 ^ new_n11706;
  assign new_n11761 = new_n11758 ^ new_n11747;
  assign new_n11762 = ~new_n11760 & ~new_n11761;
  assign new_n11763 = new_n11762 ^ new_n11753;
  assign new_n11764 = new_n11763 ^ new_n11706;
  assign new_n11765 = new_n11764 ^ new_n11751;
  assign new_n11766 = new_n11714 & new_n11759;
  assign new_n11767 = new_n11766 ^ new_n11714;
  assign new_n11768 = new_n11767 ^ new_n11753;
  assign new_n11769 = new_n11768 ^ new_n11730;
  assign new_n11770 = new_n11729 ^ new_n11700;
  assign new_n11771 = new_n11736 ^ new_n11700;
  assign new_n11772 = new_n11771 ^ new_n11730;
  assign new_n11773 = ~new_n11772 & new_n11770;
  assign new_n11774 = new_n11773 ^ new_n11748;
  assign new_n11775 = new_n11736 ^ new_n11721;
  assign new_n11776 = new_n11775 ^ new_n11774;
  assign new_n11777 = new_n11776 ^ new_n11769;
  assign new_n11778 = new_n11770 ^ new_n11752;
  assign new_n11779 = ~new_n11723 & ~new_n11778;
  assign new_n11780 = new_n11779 ^ new_n11742;
  assign new_n11781 = new_n11780 ^ new_n11723;
  assign new_n11782 = new_n11758 ^ new_n11723;
  assign new_n11783 = new_n11759 ^ new_n11714;
  assign new_n11784 = new_n11783 ^ new_n11730;
  assign new_n11785 = new_n11782 & new_n11784;
  assign new_n11786 = new_n11785 ^ new_n11774;
  assign new_n11787 = new_n11786 ^ new_n11729;
  assign new_n11788 = new_n11787 ^ new_n11781;
  assign new_n11789 = ~new_n11777 & new_n11788;
  assign new_n11790 = new_n11759 ^ new_n11700;
  assign new_n11791 = ~new_n11758 & ~new_n11790;
  assign new_n11792 = new_n11791 ^ new_n11700;
  assign new_n11793 = new_n11792 ^ new_n11780;
  assign new_n11794 = new_n11793 ^ new_n11789;
  assign new_n11795 = new_n11794 ^ new_n11751;
  assign new_n11796 = new_n11773 ^ new_n11745;
  assign new_n11797 = new_n11766 ^ new_n11762;
  assign new_n11798 = new_n11797 ^ new_n11796;
  assign new_n11799 = ~new_n11795 & ~new_n11798;
  assign new_n11800 = new_n11799 ^ new_n11789;
  assign new_n11801 = ~new_n11800 & new_n11765;
  assign new_n11802 = new_n11801 ^ new_n11765;
  assign new_n11803 = new_n11802 ^ new_n11777;
  assign new_n11804 = ~new_n11723 & ~new_n11803;
  assign new_n11805 = new_n11802 ^ new_n11799;
  assign new_n11806 = new_n11805 ^ new_n11798;
  assign new_n11807 = ~new_n11806 & new_n11782;
  assign new_n11808 = new_n11807 ^ new_n11804;
  assign new_n11809 = ~new_n11778 & ~new_n11803;
  assign new_n11810 = new_n11809 ^ new_n11808;
  assign new_n11811 = new_n11736 ^ new_n11706;
  assign new_n11812 = new_n11791 ^ new_n11785;
  assign new_n11813 = new_n11812 ^ new_n11796;
  assign new_n11814 = new_n11813 ^ new_n11811;
  assign new_n11815 = new_n11789 ^ new_n11765;
  assign new_n11816 = ~new_n11814 & new_n11815;
  assign new_n11817 = new_n11816 ^ new_n11793;
  assign new_n11818 = new_n11817 ^ new_n11751;
  assign new_n11819 = new_n11801 ^ new_n11789;
  assign new_n11820 = ~new_n11818 & new_n11819;
  assign new_n11821 = new_n11820 ^ new_n11816;
  assign new_n11822 = new_n11821 ^ new_n11788;
  assign new_n11823 = new_n11750 & new_n11822;
  assign new_n11824 = new_n11816 ^ new_n11799;
  assign new_n11825 = new_n11793 ^ new_n11764;
  assign new_n11826 = new_n11825 ^ new_n11824;
  assign new_n11827 = ~new_n11826 & new_n11707;
  assign new_n11828 = new_n11736 ^ new_n11714;
  assign new_n11829 = new_n11785 ^ new_n11767;
  assign new_n11830 = new_n11820 ^ new_n11802;
  assign new_n11831 = new_n11830 ^ new_n11829;
  assign new_n11832 = new_n11831 ^ new_n11828;
  assign new_n11833 = new_n11832 ^ new_n11700;
  assign new_n11834 = new_n11816 ^ new_n11753;
  assign new_n11835 = new_n11834 ^ new_n11780;
  assign new_n11836 = new_n11835 ^ new_n11833;
  assign new_n11837 = ~new_n11836 & new_n11770;
  assign new_n11838 = new_n11837 ^ new_n11827;
  assign new_n11839 = ~new_n11806 & new_n11784;
  assign new_n11840 = new_n11839 ^ new_n11838;
  assign new_n11841 = new_n11820 ^ new_n11814;
  assign new_n11842 = ~new_n11759 & ~new_n11841;
  assign new_n11843 = new_n11842 ^ new_n11840;
  assign new_n11844 = new_n11843 ^ new_n11823;
  assign new_n11845 = new_n11844 ^ new_n11810;
  assign new_n11846 = new_n10082 ^ new_n10029;
  assign new_n11847 = new_n9000 ^ new_n855;
  assign new_n11848 = new_n11847 ^ new_n9930;
  assign new_n11849 = new_n11848 ^ new_n9868;
  assign new_n11850 = new_n11849 ^ new_n11846;
  assign new_n11851 = new_n9716 ^ new_n9300;
  assign new_n11852 = new_n11851 ^ new_n10069;
  assign new_n11853 = new_n8930 ^ new_n883;
  assign new_n11854 = new_n11853 ^ new_n10082;
  assign new_n11855 = new_n11854 ^ new_n9960;
  assign new_n11856 = new_n11855 ^ new_n11852;
  assign new_n11857 = new_n10082 ^ new_n9884;
  assign new_n11858 = new_n11857 ^ new_n10030;
  assign new_n11859 = new_n8903 ^ new_n891;
  assign new_n11860 = new_n11859 ^ new_n9927;
  assign new_n11861 = new_n11860 ^ new_n9964;
  assign new_n11862 = new_n11861 ^ new_n11858;
  assign new_n11863 = new_n11862 ^ new_n11856;
  assign new_n11864 = new_n9043 ^ new_n874;
  assign new_n11865 = new_n11864 ^ new_n9996;
  assign new_n11866 = new_n10079 ^ new_n9859;
  assign new_n11867 = new_n11866 ^ new_n9855;
  assign new_n11868 = new_n11867 ^ new_n11865;
  assign new_n11869 = new_n9064 ^ new_n864;
  assign new_n11870 = new_n11869 ^ new_n10082;
  assign new_n11871 = new_n11870 ^ new_n9851;
  assign new_n11872 = new_n10061 ^ new_n10052;
  assign new_n11873 = new_n11872 ^ new_n10048;
  assign new_n11874 = new_n11873 ^ new_n11871;
  assign new_n11875 = new_n11874 ^ new_n11868;
  assign new_n11876 = new_n11875 ^ new_n11863;
  assign new_n11877 = new_n11876 ^ new_n11850;
  assign new_n11878 = new_n9959 ^ new_n9321;
  assign new_n11879 = new_n11878 ^ new_n9474;
  assign new_n11880 = new_n8351 ^ new_n902;
  assign new_n11881 = new_n11880 ^ new_n9901;
  assign new_n11882 = new_n11881 ^ new_n11879;
  assign new_n11883 = new_n11882 ^ new_n11863;
  assign new_n11884 = new_n10041 ^ new_n9989;
  assign new_n11885 = new_n8984 ^ new_n819;
  assign new_n11886 = new_n11885 ^ new_n10013;
  assign new_n11887 = new_n11886 ^ new_n10077;
  assign new_n11888 = new_n11887 ^ new_n11884;
  assign new_n11889 = new_n11888 ^ new_n11883;
  assign new_n11890 = new_n11875 & new_n11889;
  assign new_n11891 = new_n11882 ^ new_n11868;
  assign new_n11892 = new_n10062 ^ new_n10040;
  assign new_n11893 = new_n9023 ^ new_n842;
  assign new_n11894 = new_n11893 ^ new_n10018;
  assign new_n11895 = new_n11894 ^ new_n10000;
  assign new_n11896 = new_n11895 ^ new_n11892;
  assign new_n11897 = new_n11896 ^ new_n11888;
  assign new_n11898 = new_n11897 ^ new_n11876;
  assign new_n11899 = ~new_n11898 & new_n11891;
  assign new_n11900 = new_n11899 ^ new_n11890;
  assign new_n11901 = new_n11896 ^ new_n11883;
  assign new_n11902 = new_n11901 ^ new_n11900;
  assign new_n11903 = new_n11868 ^ new_n11862;
  assign new_n11904 = ~new_n11903 & new_n11901;
  assign new_n11905 = new_n11897 ^ new_n11850;
  assign new_n11906 = new_n11905 ^ new_n11868;
  assign new_n11907 = new_n11889 ^ new_n11850;
  assign new_n11908 = ~new_n11906 & ~new_n11907;
  assign new_n11909 = new_n11908 ^ new_n11904;
  assign new_n11910 = new_n11909 ^ new_n11868;
  assign new_n11911 = new_n11910 ^ new_n11902;
  assign new_n11912 = new_n11905 ^ new_n11874;
  assign new_n11913 = ~new_n11850 & ~new_n11912;
  assign new_n11914 = new_n11913 ^ new_n11874;
  assign new_n11915 = new_n11882 ^ new_n11874;
  assign new_n11916 = new_n11915 ^ new_n11903;
  assign new_n11917 = ~new_n11876 & ~new_n11916;
  assign new_n11918 = new_n11917 ^ new_n11888;
  assign new_n11919 = new_n11918 ^ new_n11914;
  assign new_n11920 = new_n11918 ^ new_n11876;
  assign new_n11921 = new_n11905 ^ new_n11862;
  assign new_n11922 = new_n11921 ^ new_n11891;
  assign new_n11923 = new_n11877 & new_n11922;
  assign new_n11924 = new_n11923 ^ new_n11890;
  assign new_n11925 = new_n11896 ^ new_n11874;
  assign new_n11926 = new_n11925 ^ new_n11891;
  assign new_n11927 = ~new_n11926 & new_n11915;
  assign new_n11928 = new_n11927 ^ new_n11882;
  assign new_n11929 = new_n11928 ^ new_n11924;
  assign new_n11930 = new_n11929 ^ new_n11920;
  assign new_n11931 = new_n11862 & new_n11905;
  assign new_n11932 = new_n11931 ^ new_n11862;
  assign new_n11933 = new_n11932 ^ new_n11904;
  assign new_n11934 = new_n11933 ^ new_n11891;
  assign new_n11935 = new_n11927 ^ new_n11890;
  assign new_n11936 = new_n11896 ^ new_n11856;
  assign new_n11937 = new_n11936 ^ new_n11935;
  assign new_n11938 = new_n11937 ^ new_n11934;
  assign new_n11939 = ~new_n11938 & new_n11930;
  assign new_n11940 = new_n11939 ^ new_n11919;
  assign new_n11941 = new_n11940 ^ new_n11902;
  assign new_n11942 = new_n11931 ^ new_n11908;
  assign new_n11943 = new_n11927 ^ new_n11899;
  assign new_n11944 = new_n11943 ^ new_n11942;
  assign new_n11945 = ~new_n11941 & ~new_n11944;
  assign new_n11946 = new_n11945 ^ new_n11939;
  assign new_n11947 = new_n11911 & new_n11946;
  assign new_n11948 = new_n11947 ^ new_n11945;
  assign new_n11949 = new_n11948 ^ new_n11944;
  assign new_n11950 = ~new_n11949 & new_n11877;
  assign new_n11951 = new_n11947 ^ new_n11938;
  assign new_n11952 = ~new_n11876 & ~new_n11951;
  assign new_n11953 = new_n11952 ^ new_n11950;
  assign new_n11954 = ~new_n11916 & ~new_n11951;
  assign new_n11955 = new_n11954 ^ new_n11953;
  assign new_n11956 = new_n11896 ^ new_n11868;
  assign new_n11957 = new_n11923 ^ new_n11913;
  assign new_n11958 = new_n11957 ^ new_n11943;
  assign new_n11959 = new_n11958 ^ new_n11956;
  assign new_n11960 = new_n11939 ^ new_n11911;
  assign new_n11961 = ~new_n11959 & new_n11960;
  assign new_n11962 = new_n11961 ^ new_n11919;
  assign new_n11963 = new_n11962 ^ new_n11902;
  assign new_n11964 = new_n11960 ^ new_n11947;
  assign new_n11965 = ~new_n11963 & new_n11964;
  assign new_n11966 = new_n11965 ^ new_n11961;
  assign new_n11967 = new_n11966 ^ new_n11930;
  assign new_n11968 = new_n11901 & new_n11967;
  assign new_n11969 = new_n11965 ^ new_n11959;
  assign new_n11970 = ~new_n11905 & ~new_n11969;
  assign new_n11971 = ~new_n11949 & new_n11922;
  assign new_n11972 = new_n11947 ^ new_n11931;
  assign new_n11973 = new_n11965 ^ new_n11896;
  assign new_n11974 = new_n11973 ^ new_n11923;
  assign new_n11975 = new_n11974 ^ new_n11972;
  assign new_n11976 = new_n11975 ^ new_n11874;
  assign new_n11977 = new_n11961 ^ new_n11904;
  assign new_n11978 = new_n11977 ^ new_n11918;
  assign new_n11979 = new_n11978 ^ new_n11976;
  assign new_n11980 = ~new_n11979 & new_n11915;
  assign new_n11981 = new_n11961 ^ new_n11945;
  assign new_n11982 = new_n11919 ^ new_n11910;
  assign new_n11983 = new_n11982 ^ new_n11981;
  assign new_n11984 = ~new_n11983 & new_n11875;
  assign new_n11985 = new_n11984 ^ new_n11980;
  assign new_n11986 = new_n11985 ^ new_n11971;
  assign new_n11987 = new_n11986 ^ new_n11970;
  assign new_n11988 = new_n11987 ^ new_n11968;
  assign new_n11989 = new_n11988 ^ new_n11955;
  assign new_n11990 = new_n11989 ^ new_n11845;
  assign new_n11991 = ~new_n11983 & new_n11889;
  assign new_n11992 = new_n11991 ^ new_n11954;
  assign new_n11993 = ~new_n11926 & ~new_n11979;
  assign new_n11994 = new_n11993 ^ new_n11988;
  assign new_n11995 = new_n11994 ^ new_n11992;
  assign new_n11996 = new_n11193 ^ new_n11189;
  assign new_n11997 = new_n11996 ^ new_n11215;
  assign new_n11998 = new_n8089 ^ new_n7787;
  assign new_n11999 = new_n11998 ^ new_n11148;
  assign new_n12000 = new_n11999 ^ new_n11080;
  assign new_n12001 = new_n12000 ^ new_n11997;
  assign new_n12002 = new_n8062 ^ new_n7965;
  assign new_n12003 = new_n12002 ^ new_n11996;
  assign new_n12004 = new_n12003 ^ new_n10984;
  assign new_n12005 = new_n11154 ^ new_n11117;
  assign new_n12006 = new_n12005 ^ new_n11159;
  assign new_n12007 = new_n12006 ^ new_n12004;
  assign new_n12008 = new_n12007 ^ new_n12001;
  assign new_n12009 = new_n11088 ^ new_n10955;
  assign new_n12010 = new_n8098 ^ new_n7937;
  assign new_n12011 = new_n12010 ^ new_n11193;
  assign new_n12012 = new_n12011 ^ new_n10814;
  assign new_n12013 = new_n12012 ^ new_n12009;
  assign new_n12014 = new_n8112 ^ new_n713;
  assign new_n12015 = new_n12014 ^ new_n11201;
  assign new_n12016 = new_n12015 ^ new_n11130;
  assign new_n12017 = new_n11174 ^ new_n11148;
  assign new_n12018 = new_n12017 ^ new_n12016;
  assign new_n12019 = new_n12018 ^ new_n12013;
  assign new_n12020 = new_n12019 ^ new_n12008;
  assign new_n12021 = new_n8081 ^ new_n7896;
  assign new_n12022 = new_n12021 ^ new_n11062;
  assign new_n12023 = new_n11143 ^ new_n11071;
  assign new_n12024 = new_n12023 ^ new_n11996;
  assign new_n12025 = new_n12024 ^ new_n12022;
  assign new_n12026 = new_n11185 ^ new_n11044;
  assign new_n12027 = new_n8076 ^ new_n7861;
  assign new_n12028 = new_n12027 ^ new_n11024;
  assign new_n12029 = new_n12028 ^ new_n10955;
  assign new_n12030 = new_n12029 ^ new_n12026;
  assign new_n12031 = new_n11044 ^ new_n10585;
  assign new_n12032 = new_n8072 ^ new_n7910;
  assign new_n12033 = new_n11117 ^ new_n11112;
  assign new_n12034 = new_n12033 ^ new_n12032;
  assign new_n12035 = new_n12034 ^ new_n12031;
  assign new_n12036 = new_n12035 ^ new_n12030;
  assign new_n12037 = new_n12036 ^ new_n12025;
  assign new_n12038 = new_n12037 ^ new_n12013;
  assign new_n12039 = new_n11201 ^ new_n11154;
  assign new_n12040 = new_n12039 ^ new_n11205;
  assign new_n12041 = new_n8106 ^ new_n7822;
  assign new_n12042 = new_n12041 ^ new_n11996;
  assign new_n12043 = new_n12042 ^ new_n11107;
  assign new_n12044 = new_n12043 ^ new_n12040;
  assign new_n12045 = new_n12044 ^ new_n12001;
  assign new_n12046 = new_n12045 ^ new_n12018;
  assign new_n12047 = new_n12046 ^ new_n12030;
  assign new_n12048 = new_n12047 ^ new_n12025;
  assign new_n12049 = new_n12038 & new_n12048;
  assign new_n12050 = new_n12046 ^ new_n12035;
  assign new_n12051 = new_n12013 ^ new_n12001;
  assign new_n12052 = new_n12050 & new_n12051;
  assign new_n12053 = new_n12052 ^ new_n12049;
  assign new_n12054 = new_n12053 ^ new_n12013;
  assign new_n12055 = new_n12013 ^ new_n12007;
  assign new_n12056 = new_n12055 ^ new_n12045;
  assign new_n12057 = new_n12056 ^ new_n12036;
  assign new_n12058 = new_n12019 & new_n12057;
  assign new_n12059 = new_n12047 & new_n12055;
  assign new_n12060 = new_n12059 ^ new_n12058;
  assign new_n12061 = new_n12060 ^ new_n12050;
  assign new_n12062 = new_n12061 ^ new_n12054;
  assign new_n12063 = ~new_n12001 & ~new_n12037;
  assign new_n12064 = new_n12063 ^ new_n12049;
  assign new_n12065 = new_n12035 ^ new_n12007;
  assign new_n12066 = new_n12065 ^ new_n12019;
  assign new_n12067 = new_n12018 ^ new_n12007;
  assign new_n12068 = new_n12066 & new_n12067;
  assign new_n12069 = new_n12068 ^ new_n12058;
  assign new_n12070 = new_n12069 ^ new_n12064;
  assign new_n12071 = ~new_n12036 & new_n12025;
  assign new_n12072 = ~new_n12025 & new_n12007;
  assign new_n12073 = new_n12072 ^ new_n12071;
  assign new_n12074 = new_n12020 & new_n12056;
  assign new_n12075 = new_n12074 ^ new_n12030;
  assign new_n12076 = new_n12075 ^ new_n12073;
  assign new_n12077 = new_n12063 ^ new_n12001;
  assign new_n12078 = new_n12077 ^ new_n12052;
  assign new_n12079 = new_n12078 ^ new_n12019;
  assign new_n12080 = new_n12068 ^ new_n12059;
  assign new_n12081 = new_n12044 ^ new_n12035;
  assign new_n12082 = new_n12081 ^ new_n12080;
  assign new_n12083 = new_n12082 ^ new_n12079;
  assign new_n12084 = new_n12075 ^ new_n12056;
  assign new_n12085 = new_n12056 ^ new_n12025;
  assign new_n12086 = new_n12037 ^ new_n12001;
  assign new_n12087 = new_n12086 ^ new_n12019;
  assign new_n12088 = new_n12085 & new_n12087;
  assign new_n12089 = new_n12088 ^ new_n12059;
  assign new_n12090 = new_n12068 ^ new_n12018;
  assign new_n12091 = new_n12090 ^ new_n12089;
  assign new_n12092 = new_n12091 ^ new_n12084;
  assign new_n12093 = ~new_n12083 & new_n12092;
  assign new_n12094 = new_n12093 ^ new_n12076;
  assign new_n12095 = new_n12094 ^ new_n12061;
  assign new_n12096 = ~new_n12070 & new_n12095;
  assign new_n12097 = new_n12096 ^ new_n12093;
  assign new_n12098 = ~new_n12062 & ~new_n12097;
  assign new_n12099 = new_n12098 ^ new_n12096;
  assign new_n12100 = new_n12093 ^ new_n12062;
  assign new_n12101 = new_n12100 ^ new_n12099;
  assign new_n12102 = new_n12101 ^ new_n12083;
  assign new_n12103 = new_n12020 & new_n12102;
  assign new_n12104 = new_n12035 ^ new_n12013;
  assign new_n12105 = new_n12073 ^ new_n12007;
  assign new_n12106 = new_n12105 ^ new_n12088;
  assign new_n12107 = new_n12106 ^ new_n12069;
  assign new_n12108 = new_n12107 ^ new_n12104;
  assign new_n12109 = new_n12100 & new_n12108;
  assign new_n12110 = new_n12109 ^ new_n12096;
  assign new_n12111 = new_n12076 ^ new_n12054;
  assign new_n12112 = new_n12111 ^ new_n12110;
  assign new_n12113 = new_n12047 & new_n12112;
  assign new_n12114 = new_n12113 ^ new_n12103;
  assign new_n12115 = new_n12109 ^ new_n12076;
  assign new_n12116 = new_n12115 ^ new_n12061;
  assign new_n12117 = ~new_n12099 & new_n12116;
  assign new_n12118 = new_n12117 ^ new_n12108;
  assign new_n12119 = new_n12037 & new_n12118;
  assign new_n12120 = new_n12101 ^ new_n12096;
  assign new_n12121 = new_n12120 ^ new_n12070;
  assign new_n12122 = new_n12087 & new_n12121;
  assign new_n12123 = new_n12035 ^ new_n12001;
  assign new_n12124 = new_n12088 ^ new_n12077;
  assign new_n12125 = new_n12117 ^ new_n12101;
  assign new_n12126 = new_n12125 ^ new_n12124;
  assign new_n12127 = new_n12126 ^ new_n12123;
  assign new_n12128 = new_n12127 ^ new_n12007;
  assign new_n12129 = new_n12109 ^ new_n12052;
  assign new_n12130 = new_n12129 ^ new_n12075;
  assign new_n12131 = new_n12130 ^ new_n12128;
  assign new_n12132 = new_n12067 & new_n12131;
  assign new_n12133 = new_n12055 & new_n12112;
  assign new_n12134 = new_n12133 ^ new_n12132;
  assign new_n12135 = new_n12134 ^ new_n12122;
  assign new_n12136 = new_n12135 ^ new_n12119;
  assign new_n12137 = new_n12117 ^ new_n12109;
  assign new_n12138 = new_n12137 ^ new_n12092;
  assign new_n12139 = new_n12050 & new_n12138;
  assign new_n12140 = new_n12139 ^ new_n12136;
  assign new_n12141 = new_n12066 & new_n12131;
  assign new_n12142 = new_n12141 ^ new_n12140;
  assign new_n12143 = new_n12142 ^ new_n12114;
  assign new_n12144 = new_n12143 ^ new_n11995;
  assign new_n12145 = new_n12144 ^ new_n11990;
  assign new_n12146 = new_n9066 ^ new_n9045;
  assign new_n12147 = new_n8932 ^ new_n8905;
  assign new_n12148 = new_n12147 ^ new_n12146;
  assign new_n12149 = new_n9025 ^ new_n8986;
  assign new_n12150 = new_n12149 ^ new_n9002;
  assign new_n12151 = new_n8905 & new_n12150;
  assign new_n12152 = new_n12151 ^ new_n8905;
  assign new_n12153 = new_n12147 ^ new_n8353;
  assign new_n12154 = new_n12153 ^ new_n9025;
  assign new_n12155 = new_n9045 ^ new_n8905;
  assign new_n12156 = ~new_n12155 & new_n12154;
  assign new_n12157 = new_n12156 ^ new_n12152;
  assign new_n12158 = new_n9045 ^ new_n8353;
  assign new_n12159 = new_n12158 ^ new_n12157;
  assign new_n12160 = new_n9066 ^ new_n9025;
  assign new_n12161 = new_n12160 ^ new_n12158;
  assign new_n12162 = new_n9066 ^ new_n8353;
  assign new_n12163 = ~new_n12161 & new_n12162;
  assign new_n12164 = new_n12153 ^ new_n8986;
  assign new_n12165 = new_n12146 & new_n12164;
  assign new_n12166 = new_n12165 ^ new_n12163;
  assign new_n12167 = new_n9025 ^ new_n8932;
  assign new_n12168 = new_n12167 ^ new_n12166;
  assign new_n12169 = new_n12168 ^ new_n12159;
  assign new_n12170 = new_n9066 ^ new_n8905;
  assign new_n12171 = new_n12170 ^ new_n12158;
  assign new_n12172 = ~new_n12148 & ~new_n12171;
  assign new_n12173 = new_n12172 ^ new_n8986;
  assign new_n12174 = new_n12173 ^ new_n12148;
  assign new_n12175 = new_n12148 ^ new_n9002;
  assign new_n12176 = new_n12150 ^ new_n8905;
  assign new_n12177 = new_n12176 ^ new_n12158;
  assign new_n12178 = new_n12175 & new_n12177;
  assign new_n12179 = new_n12178 ^ new_n8353;
  assign new_n12180 = new_n12179 ^ new_n12166;
  assign new_n12181 = new_n12180 ^ new_n12174;
  assign new_n12182 = ~new_n12169 & new_n12181;
  assign new_n12183 = new_n12149 ^ new_n12148;
  assign new_n12184 = ~new_n12183 & new_n12158;
  assign new_n12185 = new_n12184 ^ new_n12165;
  assign new_n12186 = new_n12185 ^ new_n12154;
  assign new_n12187 = new_n12164 ^ new_n9002;
  assign new_n12188 = new_n12150 ^ new_n9045;
  assign new_n12189 = ~new_n12187 & ~new_n12188;
  assign new_n12190 = new_n12189 ^ new_n12156;
  assign new_n12191 = new_n12190 ^ new_n9045;
  assign new_n12192 = new_n12191 ^ new_n12186;
  assign new_n12193 = new_n12192 ^ new_n12182;
  assign new_n12194 = new_n12150 ^ new_n9066;
  assign new_n12195 = ~new_n9002 & ~new_n12194;
  assign new_n12196 = new_n12195 ^ new_n9066;
  assign new_n12197 = new_n12196 ^ new_n12173;
  assign new_n12198 = new_n12197 ^ new_n12182;
  assign new_n12199 = new_n12198 ^ new_n12186;
  assign new_n12200 = new_n12184 ^ new_n12163;
  assign new_n12201 = new_n12189 ^ new_n12151;
  assign new_n12202 = new_n12201 ^ new_n12200;
  assign new_n12203 = ~new_n12199 & ~new_n12202;
  assign new_n12204 = new_n12203 ^ new_n12182;
  assign new_n12205 = ~new_n12192 & ~new_n12204;
  assign new_n12206 = new_n12205 ^ new_n12203;
  assign new_n12207 = new_n12206 ^ new_n12193;
  assign new_n12208 = new_n12207 ^ new_n12169;
  assign new_n12209 = ~new_n12148 & new_n12208;
  assign new_n12210 = new_n12207 ^ new_n12203;
  assign new_n12211 = new_n12210 ^ new_n12202;
  assign new_n12212 = new_n12175 & new_n12211;
  assign new_n12213 = new_n12212 ^ new_n12209;
  assign new_n12214 = ~new_n12171 & new_n12208;
  assign new_n12215 = new_n12214 ^ new_n12213;
  assign new_n12216 = new_n9045 ^ new_n9025;
  assign new_n12217 = new_n12195 ^ new_n12178;
  assign new_n12218 = new_n12217 ^ new_n12200;
  assign new_n12219 = new_n12218 ^ new_n12216;
  assign new_n12220 = ~new_n12219 & new_n12193;
  assign new_n12221 = new_n12220 ^ new_n12197;
  assign new_n12222 = new_n12221 ^ new_n12186;
  assign new_n12223 = ~new_n12206 & ~new_n12222;
  assign new_n12224 = new_n12223 ^ new_n12220;
  assign new_n12225 = new_n12224 ^ new_n12181;
  assign new_n12226 = new_n12154 & new_n12225;
  assign new_n12227 = new_n12220 ^ new_n12203;
  assign new_n12228 = new_n12197 ^ new_n12191;
  assign new_n12229 = new_n12228 ^ new_n12227;
  assign new_n12230 = ~new_n12229 & new_n12146;
  assign new_n12231 = new_n9025 ^ new_n8905;
  assign new_n12232 = new_n12178 ^ new_n12152;
  assign new_n12233 = new_n12223 ^ new_n12207;
  assign new_n12234 = new_n12233 ^ new_n12232;
  assign new_n12235 = new_n12234 ^ new_n12231;
  assign new_n12236 = new_n12235 ^ new_n9066;
  assign new_n12237 = new_n12220 ^ new_n12156;
  assign new_n12238 = new_n12237 ^ new_n12173;
  assign new_n12239 = new_n12238 ^ new_n12236;
  assign new_n12240 = new_n12162 & new_n12239;
  assign new_n12241 = new_n12240 ^ new_n12230;
  assign new_n12242 = new_n12177 & new_n12211;
  assign new_n12243 = new_n12242 ^ new_n12241;
  assign new_n12244 = new_n12223 ^ new_n12219;
  assign new_n12245 = ~new_n12150 & ~new_n12244;
  assign new_n12246 = new_n12245 ^ new_n12243;
  assign new_n12247 = new_n12246 ^ new_n12226;
  assign new_n12248 = new_n12247 ^ new_n12215;
  assign new_n12249 = new_n12248 ^ n20;
  assign new_n12250 = new_n12249 ^ new_n12145;
  assign new_n12251 = new_n12048 & new_n12116;
  assign new_n12252 = new_n12251 ^ new_n12103;
  assign new_n12253 = new_n12085 & new_n12121;
  assign new_n12254 = new_n12096 ^ new_n12062;
  assign new_n12255 = new_n12025 & new_n12254;
  assign new_n12256 = new_n12255 ^ new_n12253;
  assign new_n12257 = new_n12256 ^ new_n12136;
  assign new_n12258 = new_n12257 ^ new_n12252;
  assign new_n12259 = ~new_n11907 & ~new_n11963;
  assign new_n12260 = new_n12259 ^ new_n11954;
  assign new_n12261 = new_n11945 ^ new_n11911;
  assign new_n12262 = ~new_n11850 & new_n12261;
  assign new_n12263 = new_n12262 ^ new_n11950;
  assign new_n12264 = new_n12263 ^ new_n11987;
  assign new_n12265 = new_n12264 ^ new_n12260;
  assign new_n12266 = new_n12265 ^ new_n12258;
  assign new_n12267 = new_n8993 ^ new_n8886;
  assign new_n12268 = new_n10184 ^ new_n9048;
  assign new_n12269 = new_n12268 ^ new_n8978;
  assign new_n12270 = new_n12269 ^ new_n12267;
  assign new_n12271 = new_n10186 ^ new_n9051;
  assign new_n12272 = new_n12271 ^ new_n9014;
  assign new_n12273 = new_n9071 ^ new_n8947;
  assign new_n12274 = new_n12273 ^ new_n8924;
  assign new_n12275 = new_n12274 ^ new_n12272;
  assign new_n12276 = new_n12275 ^ new_n12270;
  assign new_n12277 = new_n9051 ^ new_n9005;
  assign new_n12278 = new_n12277 ^ new_n8857;
  assign new_n12279 = new_n10201 ^ new_n8895;
  assign new_n12280 = new_n12279 ^ new_n8998;
  assign new_n12281 = new_n12280 ^ new_n12278;
  assign new_n12282 = new_n8924 ^ new_n8701;
  assign new_n12283 = new_n12282 ^ new_n8224;
  assign new_n12284 = new_n10208 ^ new_n9063;
  assign new_n12285 = new_n12284 ^ new_n9051;
  assign new_n12286 = new_n12285 ^ new_n12283;
  assign new_n12287 = new_n12286 ^ new_n12281;
  assign new_n12288 = new_n12287 ^ new_n12276;
  assign new_n12289 = new_n8940 ^ new_n8867;
  assign new_n12290 = new_n10204 ^ new_n8224;
  assign new_n12291 = new_n12290 ^ new_n8895;
  assign new_n12292 = new_n12291 ^ new_n12289;
  assign new_n12293 = new_n12292 ^ new_n12270;
  assign new_n12294 = new_n9019 ^ new_n8966;
  assign new_n12295 = new_n9071 ^ new_n9069;
  assign new_n12296 = new_n12295 ^ new_n10191;
  assign new_n12297 = new_n12296 ^ new_n12294;
  assign new_n12298 = new_n9041 ^ new_n9030;
  assign new_n12299 = new_n10193 ^ new_n8978;
  assign new_n12300 = new_n12299 ^ new_n9019;
  assign new_n12301 = new_n12300 ^ new_n12298;
  assign new_n12302 = new_n12301 ^ new_n12297;
  assign new_n12303 = new_n12302 ^ new_n12288;
  assign new_n12304 = ~new_n12293 & new_n12303;
  assign new_n12305 = new_n12292 ^ new_n12287;
  assign new_n12306 = new_n12305 ^ new_n12301;
  assign new_n12307 = ~new_n12306 & new_n12276;
  assign new_n12308 = new_n12307 ^ new_n12304;
  assign new_n12309 = new_n12305 ^ new_n12297;
  assign new_n12310 = new_n12309 ^ new_n12308;
  assign new_n12311 = new_n12281 ^ new_n12270;
  assign new_n12312 = ~new_n12309 & new_n12311;
  assign new_n12313 = new_n10189 ^ new_n8998;
  assign new_n12314 = new_n9051 ^ new_n8916;
  assign new_n12315 = new_n12314 ^ new_n12313;
  assign new_n12316 = new_n12315 ^ new_n12306;
  assign new_n12317 = new_n12315 ^ new_n12302;
  assign new_n12318 = new_n12317 ^ new_n12270;
  assign new_n12319 = ~new_n12316 & new_n12318;
  assign new_n12320 = new_n12319 ^ new_n12312;
  assign new_n12321 = new_n12320 ^ new_n12270;
  assign new_n12322 = new_n12321 ^ new_n12310;
  assign new_n12323 = ~new_n12281 & ~new_n12317;
  assign new_n12324 = new_n12323 ^ new_n12281;
  assign new_n12325 = new_n12324 ^ new_n12312;
  assign new_n12326 = new_n12325 ^ new_n12293;
  assign new_n12327 = new_n12297 ^ new_n12275;
  assign new_n12328 = new_n12327 ^ new_n12293;
  assign new_n12329 = new_n12292 ^ new_n12275;
  assign new_n12330 = ~new_n12328 & ~new_n12329;
  assign new_n12331 = new_n12330 ^ new_n12307;
  assign new_n12332 = new_n12297 ^ new_n12286;
  assign new_n12333 = new_n12332 ^ new_n12331;
  assign new_n12334 = new_n12333 ^ new_n12326;
  assign new_n12335 = new_n12281 ^ new_n12275;
  assign new_n12336 = new_n12335 ^ new_n12293;
  assign new_n12337 = ~new_n12336 & new_n12288;
  assign new_n12338 = new_n12337 ^ new_n12301;
  assign new_n12339 = new_n12338 ^ new_n12288;
  assign new_n12340 = new_n12315 ^ new_n12288;
  assign new_n12341 = new_n12317 ^ new_n12281;
  assign new_n12342 = new_n12341 ^ new_n12293;
  assign new_n12343 = ~new_n12342 & new_n12340;
  assign new_n12344 = new_n12343 ^ new_n12292;
  assign new_n12345 = new_n12344 ^ new_n12331;
  assign new_n12346 = new_n12345 ^ new_n12339;
  assign new_n12347 = ~new_n12346 & new_n12334;
  assign new_n12348 = new_n12317 ^ new_n12275;
  assign new_n12349 = new_n12315 & new_n12348;
  assign new_n12350 = new_n12349 ^ new_n12275;
  assign new_n12351 = new_n12350 ^ new_n12338;
  assign new_n12352 = new_n12351 ^ new_n12347;
  assign new_n12353 = new_n12352 ^ new_n12310;
  assign new_n12354 = new_n12330 ^ new_n12304;
  assign new_n12355 = new_n12323 ^ new_n12319;
  assign new_n12356 = new_n12355 ^ new_n12354;
  assign new_n12357 = ~new_n12353 & ~new_n12356;
  assign new_n12358 = new_n12357 ^ new_n12347;
  assign new_n12359 = ~new_n12322 & ~new_n12358;
  assign new_n12360 = new_n12359 ^ new_n12322;
  assign new_n12361 = new_n12360 ^ new_n12334;
  assign new_n12362 = ~new_n12361 & new_n12288;
  assign new_n12363 = new_n12360 ^ new_n12357;
  assign new_n12364 = new_n12363 ^ new_n12356;
  assign new_n12365 = new_n12340 & new_n12364;
  assign new_n12366 = new_n12365 ^ new_n12362;
  assign new_n12367 = ~new_n12336 & ~new_n12361;
  assign new_n12368 = new_n12367 ^ new_n12366;
  assign new_n12369 = new_n12297 ^ new_n12270;
  assign new_n12370 = new_n12349 ^ new_n12343;
  assign new_n12371 = new_n12370 ^ new_n12354;
  assign new_n12372 = new_n12371 ^ new_n12369;
  assign new_n12373 = new_n12347 ^ new_n12322;
  assign new_n12374 = ~new_n12373 & new_n12372;
  assign new_n12375 = new_n12374 ^ new_n12351;
  assign new_n12376 = new_n12375 ^ new_n12310;
  assign new_n12377 = new_n12359 ^ new_n12347;
  assign new_n12378 = ~new_n12376 & new_n12377;
  assign new_n12379 = new_n12378 ^ new_n12374;
  assign new_n12380 = new_n12379 ^ new_n12346;
  assign new_n12381 = ~new_n12309 & ~new_n12380;
  assign new_n12382 = new_n12374 ^ new_n12357;
  assign new_n12383 = new_n12351 ^ new_n12321;
  assign new_n12384 = new_n12383 ^ new_n12382;
  assign new_n12385 = new_n12276 & new_n12384;
  assign new_n12386 = new_n12297 ^ new_n12281;
  assign new_n12387 = new_n12343 ^ new_n12324;
  assign new_n12388 = new_n12378 ^ new_n12360;
  assign new_n12389 = new_n12388 ^ new_n12387;
  assign new_n12390 = new_n12389 ^ new_n12386;
  assign new_n12391 = new_n12390 ^ new_n12275;
  assign new_n12392 = new_n12374 ^ new_n12312;
  assign new_n12393 = new_n12392 ^ new_n12338;
  assign new_n12394 = new_n12393 ^ new_n12391;
  assign new_n12395 = ~new_n12329 & new_n12394;
  assign new_n12396 = new_n12395 ^ new_n12385;
  assign new_n12397 = ~new_n12342 & new_n12364;
  assign new_n12398 = new_n12397 ^ new_n12396;
  assign new_n12399 = new_n12378 ^ new_n12372;
  assign new_n12400 = new_n12317 & new_n12399;
  assign new_n12401 = new_n12400 ^ new_n12398;
  assign new_n12402 = new_n12401 ^ new_n12381;
  assign new_n12403 = new_n12402 ^ new_n12368;
  assign new_n12404 = new_n12403 ^ new_n12266;
  assign new_n12405 = new_n12404 ^ new_n12250;
  assign new_n12406 = new_n12056 & new_n12102;
  assign new_n12407 = new_n12406 ^ new_n12253;
  assign new_n12408 = new_n12407 ^ new_n12103;
  assign new_n12409 = new_n12408 ^ new_n12140;
  assign new_n12410 = new_n12409 ^ new_n11989;
  assign new_n12411 = ~new_n12306 & new_n12384;
  assign new_n12412 = new_n12411 ^ new_n12385;
  assign new_n12413 = new_n12357 ^ new_n12270;
  assign new_n12414 = new_n12349 ^ new_n12319;
  assign new_n12415 = new_n12414 ^ new_n12390;
  assign new_n12416 = new_n12415 ^ new_n12413;
  assign new_n12417 = ~new_n12293 & new_n12416;
  assign new_n12418 = ~new_n12376 & new_n12318;
  assign new_n12419 = new_n12303 & new_n12416;
  assign new_n12420 = new_n12419 ^ new_n12418;
  assign new_n12421 = new_n12357 ^ new_n12322;
  assign new_n12422 = ~new_n12421 & new_n12315;
  assign new_n12423 = new_n12422 ^ new_n12362;
  assign new_n12424 = ~new_n12380 & new_n12311;
  assign new_n12425 = new_n12424 ^ new_n12423;
  assign new_n12426 = new_n12425 ^ new_n12420;
  assign new_n12427 = new_n12426 ^ new_n12417;
  assign new_n12428 = new_n12427 ^ new_n12412;
  assign new_n12429 = new_n12428 ^ new_n12410;
  assign new_n12430 = ~new_n11826 & new_n11747;
  assign new_n12431 = new_n12430 ^ new_n11827;
  assign new_n12432 = new_n11799 ^ new_n11706;
  assign new_n12433 = new_n11791 ^ new_n11762;
  assign new_n12434 = new_n12433 ^ new_n11832;
  assign new_n12435 = new_n12434 ^ new_n12432;
  assign new_n12436 = new_n11730 & new_n12435;
  assign new_n12437 = new_n11799 ^ new_n11765;
  assign new_n12438 = ~new_n11758 & new_n12437;
  assign new_n12439 = new_n12438 ^ new_n11804;
  assign new_n12440 = ~new_n11752 & new_n11822;
  assign new_n12441 = new_n12440 ^ new_n12439;
  assign new_n12442 = ~new_n11760 & ~new_n11818;
  assign new_n12443 = ~new_n11744 & new_n12435;
  assign new_n12444 = new_n12443 ^ new_n12442;
  assign new_n12445 = new_n12444 ^ new_n12441;
  assign new_n12446 = new_n12445 ^ new_n12436;
  assign new_n12447 = new_n12446 ^ new_n12431;
  assign new_n12448 = new_n11991 ^ new_n11984;
  assign new_n12449 = new_n11945 ^ new_n11868;
  assign new_n12450 = new_n11913 ^ new_n11908;
  assign new_n12451 = new_n12450 ^ new_n11975;
  assign new_n12452 = new_n12451 ^ new_n12449;
  assign new_n12453 = new_n11891 & new_n12452;
  assign new_n12454 = ~new_n11903 & new_n11967;
  assign new_n12455 = new_n12262 ^ new_n11952;
  assign new_n12456 = new_n12455 ^ new_n12454;
  assign new_n12457 = ~new_n11898 & new_n12452;
  assign new_n12458 = ~new_n11906 & ~new_n11963;
  assign new_n12459 = new_n12458 ^ new_n12457;
  assign new_n12460 = new_n12459 ^ new_n12456;
  assign new_n12461 = new_n12460 ^ new_n12453;
  assign new_n12462 = new_n12461 ^ new_n12448;
  assign new_n12463 = new_n12462 ^ new_n12447;
  assign new_n12464 = ~new_n12229 & new_n12164;
  assign new_n12465 = new_n12464 ^ new_n12230;
  assign new_n12466 = ~new_n12188 & ~new_n12222;
  assign new_n12467 = new_n12203 ^ new_n9045;
  assign new_n12468 = new_n12195 ^ new_n12189;
  assign new_n12469 = new_n12468 ^ new_n12235;
  assign new_n12470 = new_n12469 ^ new_n12467;
  assign new_n12471 = ~new_n12183 & ~new_n12470;
  assign new_n12472 = new_n12471 ^ new_n12466;
  assign new_n12473 = new_n12203 ^ new_n12192;
  assign new_n12474 = ~new_n9002 & new_n12473;
  assign new_n12475 = new_n12474 ^ new_n12209;
  assign new_n12476 = ~new_n12155 & new_n12225;
  assign new_n12477 = new_n12476 ^ new_n12475;
  assign new_n12478 = new_n12477 ^ new_n12472;
  assign new_n12479 = ~new_n12470 & new_n12158;
  assign new_n12480 = new_n12479 ^ new_n12478;
  assign new_n12481 = new_n12480 ^ new_n12465;
  assign new_n12482 = new_n12481 ^ n19;
  assign new_n12483 = new_n12482 ^ new_n12463;
  assign new_n12484 = new_n12483 ^ new_n12429;
  assign new_n12485 = new_n12133 ^ new_n12113;
  assign new_n12486 = new_n12096 ^ new_n12013;
  assign new_n12487 = new_n12105 ^ new_n12049;
  assign new_n12488 = new_n12487 ^ new_n12127;
  assign new_n12489 = new_n12488 ^ new_n12486;
  assign new_n12490 = new_n12019 & new_n12489;
  assign new_n12491 = new_n12038 & new_n12116;
  assign new_n12492 = new_n12057 & new_n12489;
  assign new_n12493 = new_n12492 ^ new_n12491;
  assign new_n12494 = new_n12406 ^ new_n12255;
  assign new_n12495 = new_n12051 & new_n12138;
  assign new_n12496 = new_n12495 ^ new_n12494;
  assign new_n12497 = new_n12496 ^ new_n12493;
  assign new_n12498 = new_n12497 ^ new_n12490;
  assign new_n12499 = new_n12498 ^ new_n12485;
  assign new_n12500 = new_n12499 ^ new_n12462;
  assign new_n12501 = ~new_n12328 & new_n12394;
  assign new_n12502 = new_n12501 ^ new_n12411;
  assign new_n12503 = new_n12398 ^ new_n12368;
  assign new_n12504 = new_n12503 ^ new_n12502;
  assign new_n12505 = new_n12504 ^ new_n12500;
  assign new_n12506 = ~new_n11772 & ~new_n11836;
  assign new_n12507 = new_n12506 ^ new_n12430;
  assign new_n12508 = new_n11840 ^ new_n11810;
  assign new_n12509 = new_n12508 ^ new_n12507;
  assign new_n12510 = new_n11993 ^ new_n11991;
  assign new_n12511 = new_n11986 ^ new_n11955;
  assign new_n12512 = new_n12511 ^ new_n12510;
  assign new_n12513 = new_n12512 ^ new_n12509;
  assign new_n12514 = ~new_n12161 & new_n12239;
  assign new_n12515 = new_n12514 ^ new_n12464;
  assign new_n12516 = new_n12243 ^ new_n12215;
  assign new_n12517 = new_n12516 ^ new_n12515;
  assign new_n12518 = new_n12517 ^ n18;
  assign new_n12519 = new_n12518 ^ new_n12513;
  assign new_n12520 = new_n12519 ^ new_n12505;
  assign new_n12521 = new_n12520 ^ new_n12484;
  assign new_n12522 = new_n12456 ^ new_n11968;
  assign new_n12523 = ~new_n11969 & new_n11921;
  assign new_n12524 = new_n12523 ^ new_n12259;
  assign new_n12525 = new_n12524 ^ new_n11985;
  assign new_n12526 = new_n12525 ^ new_n12522;
  assign new_n12527 = new_n12526 ^ new_n12144;
  assign new_n12528 = new_n12425 ^ new_n12381;
  assign new_n12529 = new_n12341 & new_n12399;
  assign new_n12530 = ~new_n12316 & ~new_n12376;
  assign new_n12531 = new_n12530 ^ new_n12529;
  assign new_n12532 = new_n12531 ^ new_n12396;
  assign new_n12533 = new_n12532 ^ new_n12528;
  assign new_n12534 = new_n12441 ^ new_n11823;
  assign new_n12535 = ~new_n11841 & new_n11783;
  assign new_n12536 = ~new_n11761 & ~new_n11818;
  assign new_n12537 = new_n12536 ^ new_n12535;
  assign new_n12538 = new_n12537 ^ new_n11838;
  assign new_n12539 = new_n12538 ^ new_n12534;
  assign new_n12540 = new_n12539 ^ new_n12533;
  assign new_n12541 = new_n12477 ^ new_n12226;
  assign new_n12542 = ~new_n12244 & new_n12176;
  assign new_n12543 = ~new_n12187 & ~new_n12222;
  assign new_n12544 = new_n12543 ^ new_n12542;
  assign new_n12545 = new_n12544 ^ new_n12241;
  assign new_n12546 = new_n12545 ^ new_n12541;
  assign new_n12547 = new_n12546 ^ n24;
  assign new_n12548 = new_n12547 ^ new_n12540;
  assign new_n12549 = new_n12548 ^ new_n12527;
  assign new_n12550 = new_n12549 ^ new_n12521;
  assign new_n12551 = new_n12550 ^ new_n12405;
  assign new_n12552 = new_n12443 ^ new_n12440;
  assign new_n12553 = new_n12506 ^ new_n11842;
  assign new_n12554 = new_n12553 ^ new_n12538;
  assign new_n12555 = new_n12554 ^ new_n12552;
  assign new_n12556 = new_n12424 ^ new_n12419;
  assign new_n12557 = new_n12501 ^ new_n12400;
  assign new_n12558 = new_n12557 ^ new_n12532;
  assign new_n12559 = new_n12558 ^ new_n12556;
  assign new_n12560 = new_n12559 ^ new_n12555;
  assign new_n12561 = new_n12560 ^ new_n12144;
  assign new_n12562 = new_n12476 ^ new_n12471;
  assign new_n12563 = new_n12514 ^ new_n12245;
  assign new_n12564 = new_n12563 ^ new_n12545;
  assign new_n12565 = new_n12564 ^ new_n12562;
  assign new_n12566 = new_n12565 ^ n23;
  assign new_n12567 = new_n12566 ^ new_n12561;
  assign new_n12568 = new_n12496 ^ new_n12139;
  assign new_n12569 = new_n12086 & new_n12118;
  assign new_n12570 = new_n12569 ^ new_n12251;
  assign new_n12571 = new_n12570 ^ new_n12134;
  assign new_n12572 = new_n12571 ^ new_n12568;
  assign new_n12573 = new_n12572 ^ new_n12526;
  assign new_n12574 = new_n12457 ^ new_n12454;
  assign new_n12575 = new_n11993 ^ new_n11970;
  assign new_n12576 = new_n12575 ^ new_n12525;
  assign new_n12577 = new_n12576 ^ new_n12574;
  assign new_n12578 = new_n12577 ^ new_n12573;
  assign new_n12579 = new_n12578 ^ new_n12567;
  assign new_n12580 = ~new_n12550 & ~new_n12579;
  assign new_n12581 = new_n12580 ^ new_n12579;
  assign new_n12582 = ~new_n12421 & new_n12348;
  assign new_n12583 = new_n12501 ^ new_n12402;
  assign new_n12584 = new_n12583 ^ new_n12582;
  assign new_n12585 = new_n12584 ^ new_n12426;
  assign new_n12586 = ~new_n11790 & new_n12437;
  assign new_n12587 = new_n12506 ^ new_n11844;
  assign new_n12588 = new_n12587 ^ new_n12586;
  assign new_n12589 = new_n12588 ^ new_n12445;
  assign new_n12590 = new_n12589 ^ new_n12585;
  assign new_n12591 = ~new_n12194 & new_n12473;
  assign new_n12592 = new_n12514 ^ new_n12247;
  assign new_n12593 = new_n12592 ^ new_n12591;
  assign new_n12594 = new_n12593 ^ new_n12478;
  assign new_n12595 = new_n12594 ^ n22;
  assign new_n12596 = new_n12595 ^ new_n12590;
  assign new_n12597 = new_n12495 ^ new_n12492;
  assign new_n12598 = new_n12141 ^ new_n12119;
  assign new_n12599 = new_n12598 ^ new_n12571;
  assign new_n12600 = new_n12599 ^ new_n12597;
  assign new_n12601 = new_n12600 ^ new_n12577;
  assign new_n12602 = ~new_n11912 & new_n12261;
  assign new_n12603 = new_n12602 ^ new_n11994;
  assign new_n12604 = new_n12603 ^ new_n12460;
  assign new_n12605 = new_n12604 ^ new_n12601;
  assign new_n12606 = new_n12605 ^ new_n12596;
  assign new_n12607 = new_n12604 ^ new_n12265;
  assign new_n12608 = new_n12037 ^ new_n12007;
  assign new_n12609 = new_n12254 & new_n12608;
  assign new_n12610 = new_n12609 ^ new_n12142;
  assign new_n12611 = new_n12610 ^ new_n12497;
  assign new_n12612 = new_n12611 ^ new_n12607;
  assign new_n12613 = new_n12530 ^ new_n12367;
  assign new_n12614 = new_n12422 ^ new_n12365;
  assign new_n12615 = new_n12614 ^ new_n12401;
  assign new_n12616 = new_n12615 ^ new_n12613;
  assign new_n12617 = new_n12536 ^ new_n11809;
  assign new_n12618 = new_n12438 ^ new_n11807;
  assign new_n12619 = new_n12618 ^ new_n11843;
  assign new_n12620 = new_n12619 ^ new_n12617;
  assign new_n12621 = new_n12620 ^ new_n12616;
  assign new_n12622 = new_n12621 ^ new_n12144;
  assign new_n12623 = new_n12543 ^ new_n12214;
  assign new_n12624 = new_n12474 ^ new_n12212;
  assign new_n12625 = new_n12624 ^ new_n12246;
  assign new_n12626 = new_n12625 ^ new_n12623;
  assign new_n12627 = new_n12626 ^ n21;
  assign new_n12628 = new_n12627 ^ new_n12622;
  assign new_n12629 = new_n12628 ^ new_n12612;
  assign new_n12630 = new_n12629 ^ new_n12579;
  assign new_n12631 = new_n12630 ^ new_n12606;
  assign new_n12632 = new_n12631 ^ new_n12484;
  assign new_n12633 = new_n12141 ^ new_n12113;
  assign new_n12634 = new_n12408 ^ new_n12135;
  assign new_n12635 = new_n12634 ^ new_n12633;
  assign new_n12636 = new_n12635 ^ new_n12512;
  assign new_n12637 = new_n12411 ^ new_n12367;
  assign new_n12638 = new_n12637 ^ new_n12583;
  assign new_n12639 = new_n12638 ^ new_n12636;
  assign new_n12640 = new_n12430 ^ new_n11809;
  assign new_n12641 = new_n12640 ^ new_n12587;
  assign new_n12642 = new_n12641 ^ new_n11995;
  assign new_n12643 = new_n12464 ^ new_n12214;
  assign new_n12644 = new_n12643 ^ new_n12592;
  assign new_n12645 = new_n12644 ^ n17;
  assign new_n12646 = new_n12645 ^ new_n12642;
  assign new_n12647 = new_n12646 ^ new_n12639;
  assign new_n12648 = new_n12647 ^ new_n12579;
  assign new_n12649 = new_n12632 & new_n12648;
  assign new_n12650 = new_n12649 ^ new_n12581;
  assign new_n12651 = new_n12647 ^ new_n12606;
  assign new_n12652 = new_n12651 ^ new_n12650;
  assign new_n12653 = new_n12631 ^ new_n12520;
  assign new_n12654 = new_n12647 ^ new_n12405;
  assign new_n12655 = new_n12653 & new_n12654;
  assign new_n12656 = new_n12484 ^ new_n12405;
  assign new_n12657 = new_n12656 ^ new_n12651;
  assign new_n12658 = new_n12606 ^ new_n12405;
  assign new_n12659 = new_n12657 & new_n12658;
  assign new_n12660 = new_n12659 ^ new_n12655;
  assign new_n12661 = new_n12629 ^ new_n12484;
  assign new_n12662 = new_n12661 ^ new_n12660;
  assign new_n12663 = new_n12662 ^ new_n12652;
  assign new_n12664 = new_n12654 ^ new_n12630;
  assign new_n12665 = new_n12579 ^ new_n12405;
  assign new_n12666 = new_n12665 ^ new_n12651;
  assign new_n12667 = new_n12664 & new_n12666;
  assign new_n12668 = new_n12667 ^ new_n12520;
  assign new_n12669 = new_n12668 ^ new_n12664;
  assign new_n12670 = new_n12664 ^ new_n12549;
  assign new_n12671 = new_n12579 ^ new_n12550;
  assign new_n12672 = new_n12671 ^ new_n12651;
  assign new_n12673 = new_n12670 & new_n12672;
  assign new_n12674 = new_n12673 ^ new_n12655;
  assign new_n12675 = new_n12659 ^ new_n12606;
  assign new_n12676 = new_n12675 ^ new_n12674;
  assign new_n12677 = new_n12676 ^ new_n12669;
  assign new_n12678 = ~new_n12663 & new_n12677;
  assign new_n12679 = new_n12549 & new_n12551;
  assign new_n12680 = new_n12679 ^ new_n12405;
  assign new_n12681 = new_n12680 ^ new_n12668;
  assign new_n12682 = new_n12681 ^ new_n12678;
  assign new_n12683 = new_n12664 ^ new_n12521;
  assign new_n12684 = new_n12651 & new_n12683;
  assign new_n12685 = new_n12684 ^ new_n12655;
  assign new_n12686 = new_n12685 ^ new_n12632;
  assign new_n12687 = new_n12686 ^ new_n12682;
  assign new_n12688 = new_n12653 ^ new_n12549;
  assign new_n12689 = new_n12647 ^ new_n12550;
  assign new_n12690 = new_n12688 & new_n12689;
  assign new_n12691 = new_n12690 ^ new_n12580;
  assign new_n12692 = new_n12684 ^ new_n12659;
  assign new_n12693 = new_n12692 ^ new_n12691;
  assign new_n12694 = ~new_n12693 & new_n12687;
  assign new_n12695 = new_n12690 ^ new_n12649;
  assign new_n12696 = new_n12695 ^ new_n12647;
  assign new_n12697 = new_n12696 ^ new_n12686;
  assign new_n12698 = new_n12697 ^ new_n12694;
  assign new_n12699 = new_n12551 & new_n12698;
  assign new_n12700 = new_n12579 ^ new_n12484;
  assign new_n12701 = new_n12673 ^ new_n12581;
  assign new_n12702 = new_n12647 ^ new_n12484;
  assign new_n12703 = new_n12679 ^ new_n12673;
  assign new_n12704 = new_n12703 ^ new_n12692;
  assign new_n12705 = new_n12704 ^ new_n12702;
  assign new_n12706 = new_n12697 ^ new_n12678;
  assign new_n12707 = new_n12705 & new_n12706;
  assign new_n12708 = new_n12707 ^ new_n12681;
  assign new_n12709 = new_n12708 ^ new_n12686;
  assign new_n12710 = new_n12694 ^ new_n12678;
  assign new_n12711 = ~new_n12710 & new_n12697;
  assign new_n12712 = new_n12711 ^ new_n12678;
  assign new_n12713 = new_n12709 & new_n12712;
  assign new_n12714 = new_n12711 ^ new_n12697;
  assign new_n12715 = new_n12714 ^ new_n12713;
  assign new_n12716 = new_n12715 ^ new_n12701;
  assign new_n12717 = new_n12716 ^ new_n12700;
  assign new_n12718 = new_n12717 ^ new_n12405;
  assign new_n12719 = new_n12707 ^ new_n12649;
  assign new_n12720 = new_n12719 ^ new_n12668;
  assign new_n12721 = new_n12720 ^ new_n12718;
  assign new_n12722 = ~new_n12721 & new_n12657;
  assign new_n12723 = new_n12713 ^ new_n12705;
  assign new_n12724 = new_n12550 & new_n12723;
  assign new_n12725 = new_n12714 ^ new_n12694;
  assign new_n12726 = new_n12725 ^ new_n12693;
  assign new_n12727 = ~new_n12726 & new_n12672;
  assign new_n12728 = ~new_n12721 & new_n12658;
  assign new_n12729 = new_n12707 ^ new_n12694;
  assign new_n12730 = new_n12696 ^ new_n12681;
  assign new_n12731 = new_n12730 ^ new_n12729;
  assign new_n12732 = new_n12654 & new_n12731;
  assign new_n12733 = new_n12732 ^ new_n12728;
  assign new_n12734 = new_n12733 ^ new_n12727;
  assign new_n12735 = new_n12734 ^ new_n12724;
  assign new_n12736 = new_n12713 ^ new_n12707;
  assign new_n12737 = new_n12736 ^ new_n12677;
  assign new_n12738 = new_n12632 & new_n12737;
  assign new_n12739 = new_n12738 ^ new_n12735;
  assign new_n12740 = new_n12739 ^ new_n12722;
  assign new_n12741 = new_n12740 ^ new_n12699;
  assign new_n12742 = new_n12689 & new_n12709;
  assign new_n12743 = new_n12694 ^ new_n12647;
  assign new_n12744 = new_n12690 ^ new_n12679;
  assign new_n12745 = new_n12744 ^ new_n12717;
  assign new_n12746 = new_n12745 ^ new_n12743;
  assign new_n12747 = ~new_n12746 & new_n12683;
  assign new_n12748 = new_n12747 ^ new_n12742;
  assign new_n12749 = new_n12549 & new_n12698;
  assign new_n12750 = new_n12714 ^ new_n12663;
  assign new_n12751 = ~new_n12750 & new_n12664;
  assign new_n12752 = new_n12751 ^ new_n12749;
  assign new_n12753 = new_n12648 & new_n12737;
  assign new_n12754 = new_n12753 ^ new_n12752;
  assign new_n12755 = new_n12754 ^ new_n12748;
  assign new_n12756 = new_n12755 ^ new_n12741;
  assign new_n12757 = new_n12756 ^ new_n11692;
  assign new_n12758 = new_n7823 ^ n21;
  assign new_n12759 = new_n7788 ^ n23;
  assign new_n12760 = new_n12759 ^ new_n12758;
  assign new_n12761 = new_n7938 ^ n17;
  assign new_n12762 = new_n7966 ^ n20;
  assign new_n12763 = new_n12762 ^ new_n12761;
  assign new_n12764 = new_n12763 ^ new_n12760;
  assign new_n12765 = new_n714 ^ n22;
  assign new_n12766 = new_n12765 ^ new_n12761;
  assign new_n12767 = new_n7911 ^ n19;
  assign new_n12768 = new_n7862 ^ n18;
  assign new_n12769 = new_n12768 ^ new_n12767;
  assign new_n12770 = new_n12769 ^ new_n12764;
  assign new_n12771 = ~new_n12770 & new_n12766;
  assign new_n12772 = new_n12765 ^ new_n12760;
  assign new_n12773 = new_n12772 ^ new_n12768;
  assign new_n12774 = new_n12763 & new_n12773;
  assign new_n12775 = new_n12774 ^ new_n12771;
  assign new_n12776 = new_n12772 ^ new_n12767;
  assign new_n12777 = new_n12776 ^ new_n12775;
  assign new_n12778 = new_n12761 ^ new_n12759;
  assign new_n12779 = ~new_n12778 & new_n12776;
  assign new_n12780 = new_n7897 ^ n24;
  assign new_n12781 = new_n12780 ^ new_n12769;
  assign new_n12782 = new_n12781 ^ new_n12761;
  assign new_n12783 = new_n12780 ^ new_n12773;
  assign new_n12784 = ~new_n12782 & ~new_n12783;
  assign new_n12785 = new_n12784 ^ new_n12779;
  assign new_n12786 = new_n12785 ^ new_n12761;
  assign new_n12787 = new_n12786 ^ new_n12777;
  assign new_n12788 = new_n12762 ^ new_n12759;
  assign new_n12789 = new_n12788 ^ new_n12766;
  assign new_n12790 = ~new_n12764 & ~new_n12789;
  assign new_n12791 = new_n12790 ^ new_n12768;
  assign new_n12792 = new_n12791 ^ new_n12764;
  assign new_n12793 = new_n12767 ^ new_n12762;
  assign new_n12794 = new_n12793 ^ new_n12766;
  assign new_n12795 = new_n12765 ^ new_n12762;
  assign new_n12796 = ~new_n12794 & new_n12795;
  assign new_n12797 = new_n12796 ^ new_n12774;
  assign new_n12798 = new_n12780 ^ new_n12764;
  assign new_n12799 = new_n12781 ^ new_n12759;
  assign new_n12800 = new_n12799 ^ new_n12766;
  assign new_n12801 = new_n12798 & new_n12800;
  assign new_n12802 = new_n12801 ^ new_n12765;
  assign new_n12803 = new_n12802 ^ new_n12797;
  assign new_n12804 = new_n12803 ^ new_n12792;
  assign new_n12805 = new_n12759 & new_n12781;
  assign new_n12806 = new_n12805 ^ new_n12759;
  assign new_n12807 = new_n12806 ^ new_n12779;
  assign new_n12808 = new_n12807 ^ new_n12766;
  assign new_n12809 = new_n12767 ^ new_n12758;
  assign new_n12810 = new_n12809 ^ new_n12797;
  assign new_n12811 = new_n12810 ^ new_n12808;
  assign new_n12812 = ~new_n12811 & new_n12804;
  assign new_n12813 = new_n12781 ^ new_n12762;
  assign new_n12814 = ~new_n12780 & ~new_n12813;
  assign new_n12815 = new_n12814 ^ new_n12762;
  assign new_n12816 = new_n12815 ^ new_n12791;
  assign new_n12817 = new_n12816 ^ new_n12812;
  assign new_n12818 = new_n12817 ^ new_n12777;
  assign new_n12819 = new_n12796 ^ new_n12771;
  assign new_n12820 = new_n12805 ^ new_n12784;
  assign new_n12821 = new_n12820 ^ new_n12819;
  assign new_n12822 = ~new_n12818 & ~new_n12821;
  assign new_n12823 = new_n12822 ^ new_n12812;
  assign new_n12824 = ~new_n12823 & new_n12787;
  assign new_n12825 = new_n12824 ^ new_n12787;
  assign new_n12826 = new_n12825 ^ new_n12811;
  assign new_n12827 = ~new_n12764 & ~new_n12826;
  assign new_n12828 = new_n12825 ^ new_n12822;
  assign new_n12829 = new_n12828 ^ new_n12821;
  assign new_n12830 = ~new_n12829 & new_n12798;
  assign new_n12831 = new_n12830 ^ new_n12827;
  assign new_n12832 = ~new_n12789 & ~new_n12826;
  assign new_n12833 = new_n12832 ^ new_n12831;
  assign new_n12834 = new_n12767 ^ new_n12761;
  assign new_n12835 = new_n12814 ^ new_n12801;
  assign new_n12836 = new_n12835 ^ new_n12819;
  assign new_n12837 = new_n12836 ^ new_n12834;
  assign new_n12838 = new_n12812 ^ new_n12787;
  assign new_n12839 = ~new_n12837 & new_n12838;
  assign new_n12840 = new_n12839 ^ new_n12816;
  assign new_n12841 = new_n12840 ^ new_n12777;
  assign new_n12842 = new_n12824 ^ new_n12812;
  assign new_n12843 = ~new_n12841 & new_n12842;
  assign new_n12844 = new_n12843 ^ new_n12839;
  assign new_n12845 = new_n12844 ^ new_n12804;
  assign new_n12846 = new_n12776 & new_n12845;
  assign new_n12847 = new_n12839 ^ new_n12822;
  assign new_n12848 = new_n12816 ^ new_n12786;
  assign new_n12849 = new_n12848 ^ new_n12847;
  assign new_n12850 = ~new_n12849 & new_n12763;
  assign new_n12851 = new_n12767 ^ new_n12759;
  assign new_n12852 = new_n12806 ^ new_n12801;
  assign new_n12853 = new_n12843 ^ new_n12825;
  assign new_n12854 = new_n12853 ^ new_n12852;
  assign new_n12855 = new_n12854 ^ new_n12851;
  assign new_n12856 = new_n12855 ^ new_n12762;
  assign new_n12857 = new_n12839 ^ new_n12779;
  assign new_n12858 = new_n12857 ^ new_n12791;
  assign new_n12859 = new_n12858 ^ new_n12856;
  assign new_n12860 = ~new_n12859 & new_n12795;
  assign new_n12861 = new_n12860 ^ new_n12850;
  assign new_n12862 = ~new_n12829 & new_n12800;
  assign new_n12863 = new_n12862 ^ new_n12861;
  assign new_n12864 = new_n12843 ^ new_n12837;
  assign new_n12865 = ~new_n12781 & ~new_n12864;
  assign new_n12866 = new_n12865 ^ new_n12863;
  assign new_n12867 = new_n12866 ^ new_n12846;
  assign new_n12868 = new_n12867 ^ new_n12833;
  assign new_n12869 = new_n12868 ^ new_n10185;
  assign new_n12870 = new_n9043 ^ new_n5609;
  assign new_n12871 = new_n12870 ^ new_n11189;
  assign new_n12872 = new_n11184 ^ new_n10955;
  assign new_n12873 = new_n12872 ^ new_n11088;
  assign new_n12874 = new_n12873 ^ new_n12871;
  assign new_n12875 = new_n11154 ^ new_n11106;
  assign new_n12876 = new_n12875 ^ new_n10984;
  assign new_n12877 = new_n9064 ^ new_n5597;
  assign new_n12878 = new_n12877 ^ new_n11112;
  assign new_n12879 = new_n11193 ^ new_n11084;
  assign new_n12880 = new_n12879 ^ new_n12878;
  assign new_n12881 = new_n12880 ^ new_n12876;
  assign new_n12882 = new_n12881 ^ new_n12874;
  assign new_n12883 = new_n11214 ^ new_n11130;
  assign new_n12884 = new_n12883 ^ new_n12879;
  assign new_n12885 = new_n8903 ^ new_n5641;
  assign new_n12886 = new_n12885 ^ new_n11126;
  assign new_n12887 = new_n12886 ^ new_n12023;
  assign new_n12888 = new_n12887 ^ new_n12884;
  assign new_n12889 = new_n8930 ^ new_n5650;
  assign new_n12890 = new_n12889 ^ new_n11159;
  assign new_n12891 = new_n12890 ^ new_n12879;
  assign new_n12892 = new_n11201 ^ new_n11173;
  assign new_n12893 = new_n12892 ^ new_n11107;
  assign new_n12894 = new_n12893 ^ new_n12891;
  assign new_n12895 = new_n12894 ^ new_n12888;
  assign new_n12896 = new_n12895 ^ new_n12882;
  assign new_n12897 = new_n9023 ^ new_n5473;
  assign new_n12898 = new_n12897 ^ new_n11024;
  assign new_n12899 = new_n11117 ^ new_n10983;
  assign new_n12900 = new_n12899 ^ new_n10585;
  assign new_n12901 = new_n12900 ^ new_n12898;
  assign new_n12902 = new_n8984 ^ new_n4901;
  assign new_n12903 = new_n12902 ^ new_n10814;
  assign new_n12904 = new_n11044 ^ new_n10565;
  assign new_n12905 = new_n12904 ^ new_n11185;
  assign new_n12906 = new_n12905 ^ new_n12903;
  assign new_n12907 = new_n12906 ^ new_n12901;
  assign new_n12908 = new_n9000 ^ new_n5544;
  assign new_n12909 = new_n12908 ^ new_n11062;
  assign new_n12910 = new_n11143 ^ new_n11079;
  assign new_n12911 = new_n12910 ^ new_n12879;
  assign new_n12912 = new_n12911 ^ new_n12909;
  assign new_n12913 = new_n12912 ^ new_n12907;
  assign new_n12914 = ~new_n12888 & ~new_n12913;
  assign new_n12915 = new_n12914 ^ new_n12888;
  assign new_n12916 = new_n8351 ^ new_n5684;
  assign new_n12917 = new_n12916 ^ new_n11205;
  assign new_n12918 = new_n12917 ^ new_n11214;
  assign new_n12919 = new_n12918 ^ new_n12017;
  assign new_n12920 = new_n12919 ^ new_n12895;
  assign new_n12921 = new_n12920 ^ new_n12901;
  assign new_n12922 = new_n12888 ^ new_n12874;
  assign new_n12923 = new_n12921 & new_n12922;
  assign new_n12924 = new_n12923 ^ new_n12915;
  assign new_n12925 = new_n12919 ^ new_n12874;
  assign new_n12926 = new_n12925 ^ new_n12924;
  assign new_n12927 = new_n12901 ^ new_n12881;
  assign new_n12928 = new_n12927 ^ new_n12925;
  assign new_n12929 = new_n12919 ^ new_n12881;
  assign new_n12930 = new_n12928 & new_n12929;
  assign new_n12931 = new_n12920 ^ new_n12906;
  assign new_n12932 = new_n12882 & new_n12931;
  assign new_n12933 = new_n12932 ^ new_n12930;
  assign new_n12934 = new_n12901 ^ new_n12894;
  assign new_n12935 = new_n12934 ^ new_n12933;
  assign new_n12936 = new_n12935 ^ new_n12926;
  assign new_n12937 = new_n12888 ^ new_n12881;
  assign new_n12938 = new_n12937 ^ new_n12925;
  assign new_n12939 = new_n12896 & new_n12938;
  assign new_n12940 = new_n12939 ^ new_n12906;
  assign new_n12941 = new_n12940 ^ new_n12896;
  assign new_n12942 = new_n12912 ^ new_n12896;
  assign new_n12943 = new_n12913 ^ new_n12888;
  assign new_n12944 = new_n12943 ^ new_n12925;
  assign new_n12945 = new_n12942 & new_n12944;
  assign new_n12946 = new_n12945 ^ new_n12932;
  assign new_n12947 = new_n12930 ^ new_n12919;
  assign new_n12948 = new_n12947 ^ new_n12946;
  assign new_n12949 = new_n12948 ^ new_n12941;
  assign new_n12950 = ~new_n12936 & new_n12949;
  assign new_n12951 = new_n12907 ^ new_n12896;
  assign new_n12952 = new_n12925 & new_n12951;
  assign new_n12953 = new_n12952 ^ new_n12932;
  assign new_n12954 = new_n12953 ^ new_n12921;
  assign new_n12955 = new_n12913 ^ new_n12874;
  assign new_n12956 = new_n12931 ^ new_n12912;
  assign new_n12957 = new_n12955 & new_n12956;
  assign new_n12958 = new_n12957 ^ new_n12923;
  assign new_n12959 = new_n12958 ^ new_n12874;
  assign new_n12960 = new_n12959 ^ new_n12954;
  assign new_n12961 = new_n12960 ^ new_n12950;
  assign new_n12962 = new_n12913 ^ new_n12881;
  assign new_n12963 = new_n12912 & new_n12962;
  assign new_n12964 = new_n12963 ^ new_n12881;
  assign new_n12965 = new_n12964 ^ new_n12940;
  assign new_n12966 = new_n12965 ^ new_n12950;
  assign new_n12967 = new_n12966 ^ new_n12954;
  assign new_n12968 = new_n12952 ^ new_n12930;
  assign new_n12969 = new_n12957 ^ new_n12914;
  assign new_n12970 = new_n12969 ^ new_n12968;
  assign new_n12971 = ~new_n12970 & new_n12967;
  assign new_n12972 = new_n12971 ^ new_n12950;
  assign new_n12973 = ~new_n12960 & ~new_n12972;
  assign new_n12974 = new_n12973 ^ new_n12971;
  assign new_n12975 = new_n12974 ^ new_n12961;
  assign new_n12976 = new_n12975 ^ new_n12936;
  assign new_n12977 = new_n12896 & new_n12976;
  assign new_n12978 = new_n12975 ^ new_n12971;
  assign new_n12979 = new_n12978 ^ new_n12970;
  assign new_n12980 = new_n12942 & new_n12979;
  assign new_n12981 = new_n12980 ^ new_n12977;
  assign new_n12982 = new_n12938 & new_n12976;
  assign new_n12983 = new_n12982 ^ new_n12981;
  assign new_n12984 = new_n12901 ^ new_n12874;
  assign new_n12985 = new_n12963 ^ new_n12945;
  assign new_n12986 = new_n12985 ^ new_n12968;
  assign new_n12987 = new_n12986 ^ new_n12984;
  assign new_n12988 = new_n12961 & new_n12987;
  assign new_n12989 = new_n12988 ^ new_n12965;
  assign new_n12990 = new_n12989 ^ new_n12954;
  assign new_n12991 = ~new_n12974 & new_n12990;
  assign new_n12992 = new_n12991 ^ new_n12988;
  assign new_n12993 = new_n12992 ^ new_n12949;
  assign new_n12994 = new_n12921 & new_n12993;
  assign new_n12995 = new_n12988 ^ new_n12971;
  assign new_n12996 = new_n12965 ^ new_n12959;
  assign new_n12997 = new_n12996 ^ new_n12995;
  assign new_n12998 = new_n12882 & new_n12997;
  assign new_n12999 = new_n12901 ^ new_n12888;
  assign new_n13000 = new_n12945 ^ new_n12915;
  assign new_n13001 = new_n12991 ^ new_n12975;
  assign new_n13002 = new_n13001 ^ new_n13000;
  assign new_n13003 = new_n13002 ^ new_n12999;
  assign new_n13004 = new_n13003 ^ new_n12881;
  assign new_n13005 = new_n12988 ^ new_n12923;
  assign new_n13006 = new_n13005 ^ new_n12940;
  assign new_n13007 = new_n13006 ^ new_n13004;
  assign new_n13008 = new_n12929 & new_n13007;
  assign new_n13009 = new_n13008 ^ new_n12998;
  assign new_n13010 = new_n12944 & new_n12979;
  assign new_n13011 = new_n13010 ^ new_n13009;
  assign new_n13012 = new_n12991 ^ new_n12987;
  assign new_n13013 = new_n12913 & new_n13012;
  assign new_n13014 = new_n13013 ^ new_n13011;
  assign new_n13015 = new_n13014 ^ new_n12994;
  assign new_n13016 = new_n13015 ^ new_n12983;
  assign new_n13017 = new_n10069 ^ new_n9959;
  assign new_n13018 = new_n13017 ^ new_n9474;
  assign new_n13019 = new_n11164 ^ new_n401;
  assign new_n13020 = new_n13019 ^ new_n11866;
  assign new_n13021 = new_n9850 ^ new_n9300;
  assign new_n13022 = new_n13021 ^ new_n13020;
  assign new_n13023 = new_n13022 ^ new_n13018;
  assign new_n13024 = new_n11866 ^ new_n10029;
  assign new_n13025 = new_n9927 ^ new_n9900;
  assign new_n13026 = new_n13025 ^ new_n13024;
  assign new_n13027 = new_n11137 ^ new_n391;
  assign new_n13028 = new_n13027 ^ new_n9964;
  assign new_n13029 = new_n13028 ^ new_n9868;
  assign new_n13030 = new_n13029 ^ new_n13026;
  assign new_n13031 = new_n13030 ^ new_n13023;
  assign new_n13032 = new_n10081 ^ new_n9855;
  assign new_n13033 = new_n13032 ^ new_n9989;
  assign new_n13034 = new_n11180 ^ new_n363;
  assign new_n13035 = new_n13034 ^ new_n9859;
  assign new_n13036 = new_n13035 ^ new_n10077;
  assign new_n13037 = new_n13036 ^ new_n13033;
  assign new_n13038 = new_n11095 ^ new_n372;
  assign new_n13039 = new_n10060 ^ new_n10048;
  assign new_n13040 = new_n13039 ^ new_n13038;
  assign new_n13041 = new_n13040 ^ new_n11866;
  assign new_n13042 = new_n10052 ^ new_n9716;
  assign new_n13043 = new_n13042 ^ new_n10069;
  assign new_n13044 = new_n13043 ^ new_n13041;
  assign new_n13045 = new_n13044 ^ new_n13037;
  assign new_n13046 = new_n13045 ^ new_n13031;
  assign new_n13047 = new_n9946 ^ new_n9321;
  assign new_n13048 = new_n13047 ^ new_n9884;
  assign new_n13049 = new_n11209 ^ new_n423;
  assign new_n13050 = new_n13049 ^ new_n9474;
  assign new_n13051 = new_n13050 ^ new_n9964;
  assign new_n13052 = new_n13051 ^ new_n13048;
  assign new_n13053 = new_n13052 ^ new_n13037;
  assign new_n13054 = new_n10013 ^ new_n9995;
  assign new_n13055 = new_n13054 ^ new_n10040;
  assign new_n13056 = new_n10686 ^ new_n431;
  assign new_n13057 = new_n13056 ^ new_n10077;
  assign new_n13058 = new_n13057 ^ new_n10000;
  assign new_n13059 = new_n13058 ^ new_n13055;
  assign new_n13060 = new_n10036 ^ new_n10018;
  assign new_n13061 = new_n13060 ^ new_n10000;
  assign new_n13062 = new_n11004 ^ new_n442;
  assign new_n13063 = new_n13062 ^ new_n11872;
  assign new_n13064 = new_n13063 ^ new_n13061;
  assign new_n13065 = new_n13064 ^ new_n13059;
  assign new_n13066 = new_n13065 ^ new_n13046;
  assign new_n13067 = ~new_n13066 & new_n13053;
  assign new_n13068 = new_n13052 ^ new_n13031;
  assign new_n13069 = new_n13068 ^ new_n13059;
  assign new_n13070 = new_n13045 & new_n13069;
  assign new_n13071 = new_n13070 ^ new_n13067;
  assign new_n13072 = new_n13068 ^ new_n13064;
  assign new_n13073 = new_n13072 ^ new_n13071;
  assign new_n13074 = new_n13037 ^ new_n13030;
  assign new_n13075 = ~new_n13074 & new_n13072;
  assign new_n13076 = new_n11055 ^ new_n411;
  assign new_n13077 = new_n13076 ^ new_n9868;
  assign new_n13078 = new_n10027 ^ new_n9930;
  assign new_n13079 = new_n13078 ^ new_n11866;
  assign new_n13080 = new_n13079 ^ new_n13077;
  assign new_n13081 = new_n13080 ^ new_n13065;
  assign new_n13082 = new_n13081 ^ new_n13037;
  assign new_n13083 = new_n13080 ^ new_n13069;
  assign new_n13084 = ~new_n13082 & ~new_n13083;
  assign new_n13085 = new_n13084 ^ new_n13075;
  assign new_n13086 = new_n13085 ^ new_n13037;
  assign new_n13087 = new_n13086 ^ new_n13073;
  assign new_n13088 = new_n13030 & new_n13081;
  assign new_n13089 = new_n13088 ^ new_n13030;
  assign new_n13090 = new_n13089 ^ new_n13075;
  assign new_n13091 = new_n13090 ^ new_n13053;
  assign new_n13092 = new_n13052 ^ new_n13044;
  assign new_n13093 = new_n13064 ^ new_n13044;
  assign new_n13094 = new_n13093 ^ new_n13053;
  assign new_n13095 = ~new_n13094 & new_n13092;
  assign new_n13096 = new_n13095 ^ new_n13070;
  assign new_n13097 = new_n13064 ^ new_n13023;
  assign new_n13098 = new_n13097 ^ new_n13096;
  assign new_n13099 = new_n13098 ^ new_n13091;
  assign new_n13100 = new_n13092 ^ new_n13074;
  assign new_n13101 = ~new_n13046 & ~new_n13100;
  assign new_n13102 = new_n13101 ^ new_n13059;
  assign new_n13103 = new_n13102 ^ new_n13046;
  assign new_n13104 = new_n13080 ^ new_n13046;
  assign new_n13105 = new_n13081 ^ new_n13030;
  assign new_n13106 = new_n13105 ^ new_n13053;
  assign new_n13107 = new_n13104 & new_n13106;
  assign new_n13108 = new_n13107 ^ new_n13070;
  assign new_n13109 = new_n13095 ^ new_n13052;
  assign new_n13110 = new_n13109 ^ new_n13108;
  assign new_n13111 = new_n13110 ^ new_n13103;
  assign new_n13112 = ~new_n13099 & new_n13111;
  assign new_n13113 = new_n13081 ^ new_n13044;
  assign new_n13114 = ~new_n13080 & ~new_n13113;
  assign new_n13115 = new_n13114 ^ new_n13044;
  assign new_n13116 = new_n13115 ^ new_n13102;
  assign new_n13117 = new_n13116 ^ new_n13112;
  assign new_n13118 = new_n13117 ^ new_n13073;
  assign new_n13119 = new_n13095 ^ new_n13067;
  assign new_n13120 = new_n13088 ^ new_n13084;
  assign new_n13121 = new_n13120 ^ new_n13119;
  assign new_n13122 = ~new_n13118 & ~new_n13121;
  assign new_n13123 = new_n13122 ^ new_n13112;
  assign new_n13124 = ~new_n13123 & new_n13087;
  assign new_n13125 = new_n13124 ^ new_n13087;
  assign new_n13126 = new_n13125 ^ new_n13099;
  assign new_n13127 = ~new_n13046 & ~new_n13126;
  assign new_n13128 = new_n13125 ^ new_n13122;
  assign new_n13129 = new_n13128 ^ new_n13121;
  assign new_n13130 = ~new_n13129 & new_n13104;
  assign new_n13131 = new_n13130 ^ new_n13127;
  assign new_n13132 = ~new_n13100 & ~new_n13126;
  assign new_n13133 = new_n13132 ^ new_n13131;
  assign new_n13134 = new_n13064 ^ new_n13037;
  assign new_n13135 = new_n13114 ^ new_n13107;
  assign new_n13136 = new_n13135 ^ new_n13119;
  assign new_n13137 = new_n13136 ^ new_n13134;
  assign new_n13138 = new_n13112 ^ new_n13087;
  assign new_n13139 = ~new_n13137 & new_n13138;
  assign new_n13140 = new_n13139 ^ new_n13116;
  assign new_n13141 = new_n13140 ^ new_n13073;
  assign new_n13142 = new_n13124 ^ new_n13112;
  assign new_n13143 = ~new_n13141 & new_n13142;
  assign new_n13144 = new_n13143 ^ new_n13139;
  assign new_n13145 = new_n13144 ^ new_n13111;
  assign new_n13146 = new_n13072 & new_n13145;
  assign new_n13147 = new_n13139 ^ new_n13122;
  assign new_n13148 = new_n13116 ^ new_n13086;
  assign new_n13149 = new_n13148 ^ new_n13147;
  assign new_n13150 = ~new_n13149 & new_n13045;
  assign new_n13151 = new_n13064 ^ new_n13030;
  assign new_n13152 = new_n13107 ^ new_n13089;
  assign new_n13153 = new_n13143 ^ new_n13125;
  assign new_n13154 = new_n13153 ^ new_n13152;
  assign new_n13155 = new_n13154 ^ new_n13151;
  assign new_n13156 = new_n13155 ^ new_n13044;
  assign new_n13157 = new_n13139 ^ new_n13075;
  assign new_n13158 = new_n13157 ^ new_n13102;
  assign new_n13159 = new_n13158 ^ new_n13156;
  assign new_n13160 = ~new_n13159 & new_n13092;
  assign new_n13161 = new_n13160 ^ new_n13150;
  assign new_n13162 = ~new_n13129 & new_n13106;
  assign new_n13163 = new_n13162 ^ new_n13161;
  assign new_n13164 = new_n13143 ^ new_n13137;
  assign new_n13165 = ~new_n13081 & ~new_n13164;
  assign new_n13166 = new_n13165 ^ new_n13163;
  assign new_n13167 = new_n13166 ^ new_n13146;
  assign new_n13168 = new_n13167 ^ new_n13133;
  assign new_n13169 = new_n13168 ^ new_n13016;
  assign new_n13170 = new_n13169 ^ new_n12869;
  assign new_n13171 = new_n7746 ^ new_n6838;
  assign new_n13172 = new_n10203 ^ new_n8588;
  assign new_n13173 = new_n13172 ^ new_n7850;
  assign new_n13174 = new_n13173 ^ new_n7797;
  assign new_n13175 = new_n13174 ^ new_n13171;
  assign new_n13176 = new_n7948 ^ new_n7945;
  assign new_n13177 = new_n10183 ^ new_n8571;
  assign new_n13178 = new_n13177 ^ new_n7809;
  assign new_n13179 = new_n13178 ^ new_n7869;
  assign new_n13180 = new_n13179 ^ new_n13176;
  assign new_n13181 = new_n13180 ^ new_n13175;
  assign new_n13182 = new_n7777 ^ new_n7766;
  assign new_n13183 = new_n7941 ^ new_n7809;
  assign new_n13184 = new_n13183 ^ new_n13182;
  assign new_n13185 = new_n10200 ^ new_n8563;
  assign new_n13186 = new_n13185 ^ new_n7900;
  assign new_n13187 = new_n13186 ^ new_n7746;
  assign new_n13188 = new_n13187 ^ new_n13184;
  assign new_n13189 = new_n10185 ^ new_n8532;
  assign new_n13190 = new_n13189 ^ new_n7958;
  assign new_n13191 = new_n13190 ^ new_n13183;
  assign new_n13192 = new_n7962 ^ new_n7926;
  assign new_n13193 = new_n13192 ^ new_n7830;
  assign new_n13194 = new_n13193 ^ new_n13191;
  assign new_n13195 = new_n13194 ^ new_n13188;
  assign new_n13196 = new_n13195 ^ new_n13181;
  assign new_n13197 = new_n10188 ^ new_n8552;
  assign new_n13198 = new_n13197 ^ new_n7777;
  assign new_n13199 = new_n13183 ^ new_n7904;
  assign new_n13200 = new_n13199 ^ new_n13198;
  assign new_n13201 = new_n7922 ^ new_n7890;
  assign new_n13202 = new_n10190 ^ new_n8541;
  assign new_n13203 = new_n7968 ^ new_n7926;
  assign new_n13204 = new_n13203 ^ new_n13202;
  assign new_n13205 = new_n13204 ^ new_n13201;
  assign new_n13206 = new_n7890 ^ new_n7882;
  assign new_n13207 = new_n10192 ^ new_n8546;
  assign new_n13208 = new_n13207 ^ new_n7916;
  assign new_n13209 = new_n13208 ^ new_n7948;
  assign new_n13210 = new_n13209 ^ new_n13206;
  assign new_n13211 = new_n13210 ^ new_n13205;
  assign new_n13212 = new_n13211 ^ new_n13200;
  assign new_n13213 = new_n13212 ^ new_n13180;
  assign new_n13214 = new_n7962 ^ new_n7850;
  assign new_n13215 = new_n13214 ^ new_n4899;
  assign new_n13216 = new_n10207 ^ new_n8580;
  assign new_n13217 = new_n13216 ^ new_n7844;
  assign new_n13218 = new_n13217 ^ new_n13183;
  assign new_n13219 = new_n13218 ^ new_n13215;
  assign new_n13220 = new_n13219 ^ new_n13188;
  assign new_n13221 = new_n13220 ^ new_n13175;
  assign new_n13222 = new_n13221 ^ new_n13210;
  assign new_n13223 = new_n13222 ^ new_n13200;
  assign new_n13224 = ~new_n13213 & ~new_n13223;
  assign new_n13225 = new_n13221 ^ new_n13205;
  assign new_n13226 = new_n13188 ^ new_n13180;
  assign new_n13227 = new_n13225 & new_n13226;
  assign new_n13228 = new_n13227 ^ new_n13224;
  assign new_n13229 = new_n13228 ^ new_n13180;
  assign new_n13230 = new_n13194 ^ new_n13180;
  assign new_n13231 = new_n13230 ^ new_n13220;
  assign new_n13232 = new_n13231 ^ new_n13211;
  assign new_n13233 = ~new_n13181 & new_n13232;
  assign new_n13234 = new_n13222 & new_n13230;
  assign new_n13235 = new_n13234 ^ new_n13233;
  assign new_n13236 = new_n13235 ^ new_n13225;
  assign new_n13237 = new_n13236 ^ new_n13229;
  assign new_n13238 = ~new_n13188 & new_n13212;
  assign new_n13239 = new_n13238 ^ new_n13188;
  assign new_n13240 = new_n13239 ^ new_n13227;
  assign new_n13241 = new_n13240 ^ new_n13181;
  assign new_n13242 = new_n13205 ^ new_n13194;
  assign new_n13243 = new_n13242 ^ new_n13181;
  assign new_n13244 = new_n13194 ^ new_n13175;
  assign new_n13245 = ~new_n13244 & new_n13243;
  assign new_n13246 = new_n13245 ^ new_n13234;
  assign new_n13247 = new_n13219 ^ new_n13205;
  assign new_n13248 = new_n13247 ^ new_n13246;
  assign new_n13249 = new_n13248 ^ new_n13241;
  assign new_n13250 = ~new_n13196 & new_n13231;
  assign new_n13251 = new_n13250 ^ new_n13210;
  assign new_n13252 = new_n13251 ^ new_n13231;
  assign new_n13253 = new_n13231 ^ new_n13200;
  assign new_n13254 = new_n13212 ^ new_n13188;
  assign new_n13255 = new_n13254 ^ new_n13181;
  assign new_n13256 = ~new_n13253 & new_n13255;
  assign new_n13257 = new_n13256 ^ new_n13175;
  assign new_n13258 = new_n13257 ^ new_n13246;
  assign new_n13259 = new_n13258 ^ new_n13252;
  assign new_n13260 = ~new_n13249 & new_n13259;
  assign new_n13261 = new_n13212 ^ new_n13194;
  assign new_n13262 = ~new_n13200 & ~new_n13261;
  assign new_n13263 = new_n13262 ^ new_n13194;
  assign new_n13264 = new_n13263 ^ new_n13251;
  assign new_n13265 = new_n13264 ^ new_n13260;
  assign new_n13266 = new_n13265 ^ new_n13236;
  assign new_n13267 = new_n13245 ^ new_n13233;
  assign new_n13268 = new_n13238 ^ new_n13224;
  assign new_n13269 = new_n13268 ^ new_n13267;
  assign new_n13270 = ~new_n13266 & ~new_n13269;
  assign new_n13271 = new_n13270 ^ new_n13260;
  assign new_n13272 = ~new_n13271 & new_n13237;
  assign new_n13273 = new_n13272 ^ new_n13237;
  assign new_n13274 = new_n13273 ^ new_n13249;
  assign new_n13275 = ~new_n13196 & ~new_n13274;
  assign new_n13276 = new_n13205 ^ new_n13180;
  assign new_n13277 = new_n13262 ^ new_n13256;
  assign new_n13278 = new_n13277 ^ new_n13267;
  assign new_n13279 = new_n13278 ^ new_n13276;
  assign new_n13280 = new_n13260 ^ new_n13237;
  assign new_n13281 = ~new_n13279 & new_n13280;
  assign new_n13282 = new_n13281 ^ new_n13270;
  assign new_n13283 = new_n13264 ^ new_n13229;
  assign new_n13284 = new_n13283 ^ new_n13282;
  assign new_n13285 = ~new_n13284 & new_n13222;
  assign new_n13286 = new_n13285 ^ new_n13275;
  assign new_n13287 = new_n13281 ^ new_n13264;
  assign new_n13288 = new_n13287 ^ new_n13236;
  assign new_n13289 = new_n13272 ^ new_n13260;
  assign new_n13290 = ~new_n13288 & new_n13289;
  assign new_n13291 = new_n13290 ^ new_n13281;
  assign new_n13292 = new_n13291 ^ new_n13259;
  assign new_n13293 = new_n13225 & new_n13292;
  assign new_n13294 = new_n13290 ^ new_n13279;
  assign new_n13295 = ~new_n13212 & ~new_n13294;
  assign new_n13296 = new_n13205 ^ new_n13188;
  assign new_n13297 = new_n13256 ^ new_n13239;
  assign new_n13298 = new_n13290 ^ new_n13273;
  assign new_n13299 = new_n13298 ^ new_n13297;
  assign new_n13300 = new_n13299 ^ new_n13296;
  assign new_n13301 = new_n13300 ^ new_n13194;
  assign new_n13302 = new_n13281 ^ new_n13227;
  assign new_n13303 = new_n13302 ^ new_n13251;
  assign new_n13304 = new_n13303 ^ new_n13301;
  assign new_n13305 = ~new_n13244 & ~new_n13304;
  assign new_n13306 = ~new_n13284 & new_n13230;
  assign new_n13307 = new_n13306 ^ new_n13305;
  assign new_n13308 = new_n13273 ^ new_n13270;
  assign new_n13309 = new_n13308 ^ new_n13269;
  assign new_n13310 = ~new_n13309 & new_n13255;
  assign new_n13311 = new_n13310 ^ new_n13307;
  assign new_n13312 = new_n13311 ^ new_n13295;
  assign new_n13313 = new_n13312 ^ new_n13293;
  assign new_n13314 = ~new_n13304 & new_n13243;
  assign new_n13315 = new_n13314 ^ new_n13313;
  assign new_n13316 = new_n13315 ^ new_n13286;
  assign new_n13317 = new_n9062 ^ new_n8939;
  assign new_n13318 = new_n13317 ^ new_n8224;
  assign new_n13319 = new_n9048 ^ new_n8881;
  assign new_n13320 = new_n13319 ^ new_n12758;
  assign new_n13321 = new_n13320 ^ new_n8953;
  assign new_n13322 = new_n13321 ^ new_n13318;
  assign new_n13323 = new_n13319 ^ new_n8998;
  assign new_n13324 = new_n13323 ^ new_n8868;
  assign new_n13325 = new_n12759 ^ new_n8848;
  assign new_n13326 = new_n13325 ^ new_n8915;
  assign new_n13327 = new_n13326 ^ new_n13324;
  assign new_n13328 = new_n13327 ^ new_n13322;
  assign new_n13329 = new_n8895 ^ new_n8702;
  assign new_n13330 = new_n12765 ^ new_n8939;
  assign new_n13331 = new_n13330 ^ new_n8848;
  assign new_n13332 = new_n13331 ^ new_n13329;
  assign new_n13333 = new_n13332 ^ new_n13328;
  assign new_n13334 = new_n12768 ^ new_n8993;
  assign new_n13335 = new_n9019 ^ new_n8965;
  assign new_n13336 = new_n13335 ^ new_n9041;
  assign new_n13337 = new_n13336 ^ new_n13334;
  assign new_n13338 = new_n13337 ^ new_n13333;
  assign new_n13339 = new_n12761 ^ new_n9050;
  assign new_n13340 = new_n9040 ^ new_n8978;
  assign new_n13341 = new_n13340 ^ new_n8886;
  assign new_n13342 = new_n13341 ^ new_n13339;
  assign new_n13343 = new_n12780 ^ new_n8915;
  assign new_n13344 = new_n13319 ^ new_n9006;
  assign new_n13345 = new_n13344 ^ new_n13343;
  assign new_n13346 = new_n12767 ^ new_n9030;
  assign new_n13347 = new_n9071 ^ new_n9012;
  assign new_n13348 = new_n13347 ^ new_n8966;
  assign new_n13349 = new_n13348 ^ new_n13346;
  assign new_n13350 = new_n13349 ^ new_n13337;
  assign new_n13351 = new_n13350 ^ new_n13345;
  assign new_n13352 = new_n13351 ^ new_n13342;
  assign new_n13353 = new_n13345 ^ new_n13338;
  assign new_n13354 = new_n13352 & new_n13353;
  assign new_n13355 = new_n13342 ^ new_n13327;
  assign new_n13356 = new_n13349 ^ new_n13333;
  assign new_n13357 = new_n13355 & new_n13356;
  assign new_n13358 = new_n13357 ^ new_n13354;
  assign new_n13359 = new_n13358 ^ new_n13342;
  assign new_n13360 = new_n13342 ^ new_n13332;
  assign new_n13361 = new_n13319 ^ new_n12762;
  assign new_n13362 = new_n13361 ^ new_n9014;
  assign new_n13363 = new_n9062 ^ new_n8924;
  assign new_n13364 = new_n13363 ^ new_n9069;
  assign new_n13365 = new_n13364 ^ new_n13362;
  assign new_n13366 = new_n13365 ^ new_n13342;
  assign new_n13367 = new_n13366 ^ new_n13328;
  assign new_n13368 = new_n13367 ^ new_n13350;
  assign new_n13369 = new_n13360 & new_n13368;
  assign new_n13370 = new_n13338 & new_n13366;
  assign new_n13371 = new_n13370 ^ new_n13369;
  assign new_n13372 = new_n13371 ^ new_n13356;
  assign new_n13373 = new_n13372 ^ new_n13359;
  assign new_n13374 = ~new_n13327 & ~new_n13351;
  assign new_n13375 = new_n13374 ^ new_n13327;
  assign new_n13376 = new_n13375 ^ new_n13357;
  assign new_n13377 = new_n13376 ^ new_n13360;
  assign new_n13378 = new_n13365 ^ new_n13332;
  assign new_n13379 = new_n13365 ^ new_n13349;
  assign new_n13380 = new_n13379 ^ new_n13360;
  assign new_n13381 = new_n13378 & new_n13380;
  assign new_n13382 = new_n13381 ^ new_n13370;
  assign new_n13383 = new_n13349 ^ new_n13322;
  assign new_n13384 = new_n13383 ^ new_n13382;
  assign new_n13385 = new_n13384 ^ new_n13377;
  assign new_n13386 = new_n13378 ^ new_n13355;
  assign new_n13387 = new_n13367 & new_n13386;
  assign new_n13388 = new_n13387 ^ new_n13337;
  assign new_n13389 = new_n13388 ^ new_n13367;
  assign new_n13390 = new_n13351 ^ new_n13327;
  assign new_n13391 = new_n13390 ^ new_n13360;
  assign new_n13392 = new_n13367 ^ new_n13345;
  assign new_n13393 = new_n13391 & new_n13392;
  assign new_n13394 = new_n13393 ^ new_n13370;
  assign new_n13395 = new_n13381 ^ new_n13332;
  assign new_n13396 = new_n13395 ^ new_n13394;
  assign new_n13397 = new_n13396 ^ new_n13389;
  assign new_n13398 = ~new_n13385 & new_n13397;
  assign new_n13399 = new_n13398 ^ new_n13373;
  assign new_n13400 = new_n13349 ^ new_n13342;
  assign new_n13401 = new_n13365 ^ new_n13351;
  assign new_n13402 = new_n13345 & new_n13401;
  assign new_n13403 = new_n13402 ^ new_n13393;
  assign new_n13404 = new_n13381 ^ new_n13369;
  assign new_n13405 = new_n13404 ^ new_n13403;
  assign new_n13406 = new_n13405 ^ new_n13400;
  assign new_n13407 = new_n13399 & new_n13406;
  assign new_n13408 = new_n13402 ^ new_n13365;
  assign new_n13409 = new_n13408 ^ new_n13388;
  assign new_n13410 = new_n13409 ^ new_n13398;
  assign new_n13411 = new_n13410 ^ new_n13372;
  assign new_n13412 = new_n13374 ^ new_n13354;
  assign new_n13413 = new_n13412 ^ new_n13404;
  assign new_n13414 = ~new_n13413 & new_n13411;
  assign new_n13415 = new_n13414 ^ new_n13407;
  assign new_n13416 = new_n13409 ^ new_n13359;
  assign new_n13417 = new_n13416 ^ new_n13415;
  assign new_n13418 = new_n13338 & new_n13417;
  assign new_n13419 = new_n13414 ^ new_n13398;
  assign new_n13420 = ~new_n13373 & ~new_n13419;
  assign new_n13421 = new_n13420 ^ new_n13414;
  assign new_n13422 = new_n13421 ^ new_n13399;
  assign new_n13423 = new_n13422 ^ new_n13385;
  assign new_n13424 = new_n13386 & new_n13423;
  assign new_n13425 = new_n13424 ^ new_n13418;
  assign new_n13426 = new_n13409 ^ new_n13407;
  assign new_n13427 = new_n13426 ^ new_n13372;
  assign new_n13428 = ~new_n13421 & new_n13427;
  assign new_n13429 = new_n13428 ^ new_n13407;
  assign new_n13430 = new_n13429 ^ new_n13397;
  assign new_n13431 = new_n13356 & new_n13430;
  assign new_n13432 = new_n13428 ^ new_n13406;
  assign new_n13433 = new_n13351 & new_n13432;
  assign new_n13434 = new_n13366 & new_n13417;
  assign new_n13435 = new_n13349 ^ new_n13327;
  assign new_n13436 = new_n13393 ^ new_n13375;
  assign new_n13437 = new_n13428 ^ new_n13422;
  assign new_n13438 = new_n13437 ^ new_n13436;
  assign new_n13439 = new_n13438 ^ new_n13435;
  assign new_n13440 = new_n13439 ^ new_n13365;
  assign new_n13441 = new_n13407 ^ new_n13357;
  assign new_n13442 = new_n13441 ^ new_n13388;
  assign new_n13443 = new_n13442 ^ new_n13440;
  assign new_n13444 = new_n13378 & new_n13443;
  assign new_n13445 = new_n13444 ^ new_n13434;
  assign new_n13446 = new_n13422 ^ new_n13414;
  assign new_n13447 = new_n13446 ^ new_n13413;
  assign new_n13448 = new_n13391 & new_n13447;
  assign new_n13449 = new_n13448 ^ new_n13445;
  assign new_n13450 = new_n13449 ^ new_n13433;
  assign new_n13451 = new_n13450 ^ new_n13431;
  assign new_n13452 = new_n13380 & new_n13443;
  assign new_n13453 = new_n13452 ^ new_n13451;
  assign new_n13454 = new_n13453 ^ new_n13425;
  assign new_n13455 = new_n13454 ^ new_n13316;
  assign new_n13456 = new_n13455 ^ new_n13170;
  assign new_n13457 = new_n13392 & new_n13447;
  assign new_n13458 = new_n13367 & new_n13423;
  assign new_n13459 = new_n13458 ^ new_n13457;
  assign new_n13460 = new_n13459 ^ new_n13424;
  assign new_n13461 = new_n13460 ^ new_n13451;
  assign new_n13462 = new_n13353 & new_n13427;
  assign new_n13463 = new_n13462 ^ new_n13424;
  assign new_n13464 = new_n13414 ^ new_n13373;
  assign new_n13465 = new_n13345 & new_n13464;
  assign new_n13466 = new_n13465 ^ new_n13457;
  assign new_n13467 = new_n13466 ^ new_n13450;
  assign new_n13468 = new_n13467 ^ new_n13463;
  assign new_n13469 = new_n13468 ^ new_n13461;
  assign new_n13470 = ~new_n13223 & ~new_n13288;
  assign new_n13471 = new_n13470 ^ new_n13275;
  assign new_n13472 = ~new_n13253 & ~new_n13309;
  assign new_n13473 = new_n13270 ^ new_n13237;
  assign new_n13474 = ~new_n13200 & new_n13473;
  assign new_n13475 = new_n13474 ^ new_n13472;
  assign new_n13476 = new_n13475 ^ new_n13312;
  assign new_n13477 = new_n13476 ^ new_n13471;
  assign new_n13478 = new_n13477 ^ new_n13469;
  assign new_n13479 = new_n13478 ^ new_n13456;
  assign new_n13480 = ~new_n13149 & new_n13069;
  assign new_n13481 = new_n13480 ^ new_n13150;
  assign new_n13482 = new_n13122 ^ new_n13037;
  assign new_n13483 = new_n13114 ^ new_n13084;
  assign new_n13484 = new_n13483 ^ new_n13155;
  assign new_n13485 = new_n13484 ^ new_n13482;
  assign new_n13486 = new_n13053 & new_n13485;
  assign new_n13487 = ~new_n13082 & ~new_n13141;
  assign new_n13488 = ~new_n13066 & new_n13485;
  assign new_n13489 = new_n13488 ^ new_n13487;
  assign new_n13490 = new_n13122 ^ new_n13087;
  assign new_n13491 = ~new_n13080 & new_n13490;
  assign new_n13492 = new_n13491 ^ new_n13127;
  assign new_n13493 = ~new_n13074 & new_n13145;
  assign new_n13494 = new_n13493 ^ new_n13492;
  assign new_n13495 = new_n13494 ^ new_n13489;
  assign new_n13496 = new_n13495 ^ new_n13486;
  assign new_n13497 = new_n13496 ^ new_n13481;
  assign new_n13498 = new_n12931 & new_n12997;
  assign new_n13499 = new_n13498 ^ new_n12998;
  assign new_n13500 = new_n12971 ^ new_n12874;
  assign new_n13501 = new_n12963 ^ new_n12957;
  assign new_n13502 = new_n13501 ^ new_n13003;
  assign new_n13503 = new_n13502 ^ new_n13500;
  assign new_n13504 = new_n12925 & new_n13503;
  assign new_n13505 = new_n12955 & new_n12990;
  assign new_n13506 = new_n12951 & new_n13503;
  assign new_n13507 = new_n13506 ^ new_n13505;
  assign new_n13508 = new_n12971 ^ new_n12960;
  assign new_n13509 = new_n12912 & new_n13508;
  assign new_n13510 = new_n13509 ^ new_n12977;
  assign new_n13511 = new_n12922 & new_n12993;
  assign new_n13512 = new_n13511 ^ new_n13510;
  assign new_n13513 = new_n13512 ^ new_n13507;
  assign new_n13514 = new_n13513 ^ new_n13504;
  assign new_n13515 = new_n13514 ^ new_n13499;
  assign new_n13516 = new_n13515 ^ new_n13497;
  assign new_n13517 = new_n13434 ^ new_n13418;
  assign new_n13518 = new_n13414 ^ new_n13342;
  assign new_n13519 = new_n13402 ^ new_n13354;
  assign new_n13520 = new_n13519 ^ new_n13439;
  assign new_n13521 = new_n13520 ^ new_n13518;
  assign new_n13522 = new_n13360 & new_n13521;
  assign new_n13523 = new_n13355 & new_n13430;
  assign new_n13524 = new_n13465 ^ new_n13458;
  assign new_n13525 = new_n13524 ^ new_n13523;
  assign new_n13526 = new_n13368 & new_n13521;
  assign new_n13527 = new_n13352 & new_n13427;
  assign new_n13528 = new_n13527 ^ new_n13526;
  assign new_n13529 = new_n13528 ^ new_n13525;
  assign new_n13530 = new_n13529 ^ new_n13522;
  assign new_n13531 = new_n13530 ^ new_n13517;
  assign new_n13532 = new_n13531 ^ new_n13516;
  assign new_n13533 = ~new_n12849 & new_n12773;
  assign new_n13534 = new_n13533 ^ new_n12850;
  assign new_n13535 = new_n12822 ^ new_n12761;
  assign new_n13536 = new_n12814 ^ new_n12784;
  assign new_n13537 = new_n13536 ^ new_n12855;
  assign new_n13538 = new_n13537 ^ new_n13535;
  assign new_n13539 = new_n12766 & new_n13538;
  assign new_n13540 = ~new_n12782 & ~new_n12841;
  assign new_n13541 = ~new_n12770 & new_n13538;
  assign new_n13542 = new_n13541 ^ new_n13540;
  assign new_n13543 = new_n12822 ^ new_n12787;
  assign new_n13544 = ~new_n12780 & new_n13543;
  assign new_n13545 = new_n13544 ^ new_n12827;
  assign new_n13546 = ~new_n12778 & new_n12845;
  assign new_n13547 = new_n13546 ^ new_n13545;
  assign new_n13548 = new_n13547 ^ new_n13542;
  assign new_n13549 = new_n13548 ^ new_n13539;
  assign new_n13550 = new_n13549 ^ new_n13534;
  assign new_n13551 = new_n13550 ^ new_n10190;
  assign new_n13552 = ~new_n13274 & new_n13231;
  assign new_n13553 = new_n13552 ^ new_n13472;
  assign new_n13554 = new_n13553 ^ new_n13275;
  assign new_n13555 = new_n13554 ^ new_n13313;
  assign new_n13556 = new_n13555 ^ new_n13461;
  assign new_n13557 = new_n13556 ^ new_n13551;
  assign new_n13558 = new_n13557 ^ new_n13532;
  assign new_n13559 = ~new_n13094 & ~new_n13159;
  assign new_n13560 = new_n13559 ^ new_n13480;
  assign new_n13561 = new_n13163 ^ new_n13133;
  assign new_n13562 = new_n13561 ^ new_n13560;
  assign new_n13563 = new_n12928 & new_n13007;
  assign new_n13564 = new_n13563 ^ new_n13498;
  assign new_n13565 = new_n13011 ^ new_n12983;
  assign new_n13566 = new_n13565 ^ new_n13564;
  assign new_n13567 = new_n13566 ^ new_n13562;
  assign new_n13568 = new_n13567 ^ new_n13531;
  assign new_n13569 = ~new_n12794 & ~new_n12859;
  assign new_n13570 = new_n13569 ^ new_n13533;
  assign new_n13571 = new_n12863 ^ new_n12833;
  assign new_n13572 = new_n13571 ^ new_n13570;
  assign new_n13573 = new_n13572 ^ new_n10192;
  assign new_n13574 = new_n13306 ^ new_n13285;
  assign new_n13575 = new_n13270 ^ new_n13180;
  assign new_n13576 = new_n13262 ^ new_n13224;
  assign new_n13577 = new_n13576 ^ new_n13300;
  assign new_n13578 = new_n13577 ^ new_n13575;
  assign new_n13579 = ~new_n13181 & new_n13578;
  assign new_n13580 = ~new_n13213 & ~new_n13288;
  assign new_n13581 = new_n13232 & new_n13578;
  assign new_n13582 = new_n13581 ^ new_n13580;
  assign new_n13583 = new_n13552 ^ new_n13474;
  assign new_n13584 = new_n13226 & new_n13292;
  assign new_n13585 = new_n13584 ^ new_n13583;
  assign new_n13586 = new_n13585 ^ new_n13582;
  assign new_n13587 = new_n13586 ^ new_n13579;
  assign new_n13588 = new_n13587 ^ new_n13574;
  assign new_n13589 = new_n13588 ^ new_n13573;
  assign new_n13590 = new_n13452 ^ new_n13418;
  assign new_n13591 = new_n13460 ^ new_n13449;
  assign new_n13592 = new_n13591 ^ new_n13590;
  assign new_n13593 = new_n13592 ^ new_n13589;
  assign new_n13594 = new_n13593 ^ new_n13568;
  assign new_n13595 = new_n13594 ^ new_n13558;
  assign new_n13596 = new_n13547 ^ new_n12846;
  assign new_n13597 = ~new_n12864 & new_n12799;
  assign new_n13598 = ~new_n12783 & ~new_n12841;
  assign new_n13599 = new_n13598 ^ new_n13597;
  assign new_n13600 = new_n13599 ^ new_n12861;
  assign new_n13601 = new_n13600 ^ new_n13596;
  assign new_n13602 = new_n13601 ^ new_n10188;
  assign new_n13603 = new_n13525 ^ new_n13431;
  assign new_n13604 = new_n13390 & new_n13432;
  assign new_n13605 = new_n13604 ^ new_n13462;
  assign new_n13606 = new_n13605 ^ new_n13445;
  assign new_n13607 = new_n13606 ^ new_n13603;
  assign new_n13608 = new_n13607 ^ new_n13602;
  assign new_n13609 = new_n13494 ^ new_n13146;
  assign new_n13610 = ~new_n13164 & new_n13105;
  assign new_n13611 = ~new_n13083 & ~new_n13141;
  assign new_n13612 = new_n13611 ^ new_n13610;
  assign new_n13613 = new_n13612 ^ new_n13161;
  assign new_n13614 = new_n13613 ^ new_n13609;
  assign new_n13615 = new_n13512 ^ new_n12994;
  assign new_n13616 = new_n12943 & new_n13012;
  assign new_n13617 = new_n12956 & new_n12990;
  assign new_n13618 = new_n13617 ^ new_n13616;
  assign new_n13619 = new_n13618 ^ new_n13009;
  assign new_n13620 = new_n13619 ^ new_n13615;
  assign new_n13621 = new_n13620 ^ new_n13614;
  assign new_n13622 = new_n13621 ^ new_n13455;
  assign new_n13623 = new_n13622 ^ new_n13608;
  assign new_n13624 = new_n13623 ^ new_n13595;
  assign new_n13625 = new_n13624 ^ new_n13479;
  assign new_n13626 = new_n13511 ^ new_n13506;
  assign new_n13627 = new_n13563 ^ new_n13013;
  assign new_n13628 = new_n13627 ^ new_n13619;
  assign new_n13629 = new_n13628 ^ new_n13626;
  assign new_n13630 = new_n13493 ^ new_n13488;
  assign new_n13631 = new_n13559 ^ new_n13165;
  assign new_n13632 = new_n13631 ^ new_n13613;
  assign new_n13633 = new_n13632 ^ new_n13630;
  assign new_n13634 = new_n13633 ^ new_n13629;
  assign new_n13635 = new_n13634 ^ new_n13607;
  assign new_n13636 = new_n13635 ^ new_n13455;
  assign new_n13637 = new_n13546 ^ new_n13541;
  assign new_n13638 = new_n13569 ^ new_n12865;
  assign new_n13639 = new_n13638 ^ new_n13600;
  assign new_n13640 = new_n13639 ^ new_n13637;
  assign new_n13641 = new_n13640 ^ new_n10200;
  assign new_n13642 = new_n13585 ^ new_n13293;
  assign new_n13643 = ~new_n13254 & ~new_n13294;
  assign new_n13644 = new_n13643 ^ new_n13470;
  assign new_n13645 = new_n13644 ^ new_n13307;
  assign new_n13646 = new_n13645 ^ new_n13642;
  assign new_n13647 = new_n13646 ^ new_n13641;
  assign new_n13648 = new_n13526 ^ new_n13523;
  assign new_n13649 = new_n13452 ^ new_n13433;
  assign new_n13650 = new_n13649 ^ new_n13606;
  assign new_n13651 = new_n13650 ^ new_n13648;
  assign new_n13652 = new_n13651 ^ new_n13647;
  assign new_n13653 = new_n13652 ^ new_n13636;
  assign new_n13654 = new_n13624 & new_n13653;
  assign new_n13655 = new_n13654 ^ new_n13653;
  assign new_n13656 = ~new_n13113 & new_n13490;
  assign new_n13657 = new_n13559 ^ new_n13167;
  assign new_n13658 = new_n13657 ^ new_n13656;
  assign new_n13659 = new_n13658 ^ new_n13495;
  assign new_n13660 = new_n12962 & new_n13508;
  assign new_n13661 = new_n13563 ^ new_n13015;
  assign new_n13662 = new_n13661 ^ new_n13660;
  assign new_n13663 = new_n13662 ^ new_n13513;
  assign new_n13664 = new_n13663 ^ new_n13659;
  assign new_n13665 = new_n13664 ^ new_n13651;
  assign new_n13666 = ~new_n12813 & new_n13543;
  assign new_n13667 = new_n13569 ^ new_n12867;
  assign new_n13668 = new_n13667 ^ new_n13666;
  assign new_n13669 = new_n13668 ^ new_n13548;
  assign new_n13670 = new_n13669 ^ new_n10203;
  assign new_n13671 = new_n13401 & new_n13464;
  assign new_n13672 = new_n13671 ^ new_n13453;
  assign new_n13673 = new_n13672 ^ new_n13529;
  assign new_n13674 = new_n13673 ^ new_n13670;
  assign new_n13675 = new_n13584 ^ new_n13581;
  assign new_n13676 = new_n13314 ^ new_n13295;
  assign new_n13677 = new_n13676 ^ new_n13645;
  assign new_n13678 = new_n13677 ^ new_n13675;
  assign new_n13679 = new_n13678 ^ new_n13674;
  assign new_n13680 = new_n13679 ^ new_n13665;
  assign new_n13681 = new_n13598 ^ new_n12832;
  assign new_n13682 = new_n13544 ^ new_n12830;
  assign new_n13683 = new_n13682 ^ new_n12866;
  assign new_n13684 = new_n13683 ^ new_n13681;
  assign new_n13685 = new_n13684 ^ new_n10207;
  assign new_n13686 = new_n13611 ^ new_n13132;
  assign new_n13687 = new_n13491 ^ new_n13130;
  assign new_n13688 = new_n13687 ^ new_n13166;
  assign new_n13689 = new_n13688 ^ new_n13686;
  assign new_n13690 = new_n13617 ^ new_n12982;
  assign new_n13691 = new_n13509 ^ new_n12980;
  assign new_n13692 = new_n13691 ^ new_n13014;
  assign new_n13693 = new_n13692 ^ new_n13690;
  assign new_n13694 = new_n13693 ^ new_n13689;
  assign new_n13695 = new_n13694 ^ new_n13685;
  assign new_n13696 = new_n13695 ^ new_n13455;
  assign new_n13697 = new_n13673 ^ new_n13468;
  assign new_n13698 = ~new_n13261 & new_n13473;
  assign new_n13699 = new_n13698 ^ new_n13315;
  assign new_n13700 = new_n13699 ^ new_n13586;
  assign new_n13701 = new_n13700 ^ new_n13697;
  assign new_n13702 = new_n13701 ^ new_n13696;
  assign new_n13703 = new_n13702 ^ new_n13653;
  assign new_n13704 = new_n13703 ^ new_n13680;
  assign new_n13705 = new_n13704 ^ new_n13558;
  assign new_n13706 = new_n13480 ^ new_n13132;
  assign new_n13707 = new_n13706 ^ new_n13657;
  assign new_n13708 = new_n13498 ^ new_n12982;
  assign new_n13709 = new_n13708 ^ new_n13661;
  assign new_n13710 = new_n13709 ^ new_n13707;
  assign new_n13711 = new_n13710 ^ new_n13592;
  assign new_n13712 = new_n13533 ^ new_n12832;
  assign new_n13713 = new_n13712 ^ new_n13667;
  assign new_n13714 = new_n13713 ^ new_n10183;
  assign new_n13715 = new_n13714 ^ new_n13454;
  assign new_n13716 = new_n13314 ^ new_n13285;
  assign new_n13717 = new_n13554 ^ new_n13311;
  assign new_n13718 = new_n13717 ^ new_n13716;
  assign new_n13719 = new_n13718 ^ new_n13715;
  assign new_n13720 = new_n13719 ^ new_n13711;
  assign new_n13721 = new_n13720 ^ new_n13653;
  assign new_n13722 = ~new_n13721 & new_n13705;
  assign new_n13723 = new_n13722 ^ new_n13655;
  assign new_n13724 = new_n13720 ^ new_n13680;
  assign new_n13725 = new_n13724 ^ new_n13723;
  assign new_n13726 = new_n13704 ^ new_n13594;
  assign new_n13727 = new_n13720 ^ new_n13479;
  assign new_n13728 = new_n13726 & new_n13727;
  assign new_n13729 = new_n13558 ^ new_n13479;
  assign new_n13730 = new_n13729 ^ new_n13724;
  assign new_n13731 = new_n13680 ^ new_n13479;
  assign new_n13732 = ~new_n13731 & new_n13730;
  assign new_n13733 = new_n13732 ^ new_n13728;
  assign new_n13734 = new_n13702 ^ new_n13558;
  assign new_n13735 = new_n13734 ^ new_n13733;
  assign new_n13736 = new_n13735 ^ new_n13725;
  assign new_n13737 = new_n13727 ^ new_n13703;
  assign new_n13738 = new_n13653 ^ new_n13479;
  assign new_n13739 = new_n13738 ^ new_n13724;
  assign new_n13740 = new_n13737 & new_n13739;
  assign new_n13741 = new_n13740 ^ new_n13594;
  assign new_n13742 = new_n13741 ^ new_n13737;
  assign new_n13743 = new_n13737 ^ new_n13623;
  assign new_n13744 = new_n13653 ^ new_n13624;
  assign new_n13745 = new_n13744 ^ new_n13724;
  assign new_n13746 = ~new_n13743 & ~new_n13745;
  assign new_n13747 = new_n13746 ^ new_n13680;
  assign new_n13748 = new_n13747 ^ new_n13733;
  assign new_n13749 = new_n13748 ^ new_n13742;
  assign new_n13750 = ~new_n13736 & new_n13749;
  assign new_n13751 = ~new_n13623 & ~new_n13625;
  assign new_n13752 = new_n13751 ^ new_n13479;
  assign new_n13753 = new_n13752 ^ new_n13741;
  assign new_n13754 = new_n13753 ^ new_n13750;
  assign new_n13755 = new_n13737 ^ new_n13595;
  assign new_n13756 = ~new_n13724 & new_n13755;
  assign new_n13757 = new_n13756 ^ new_n13728;
  assign new_n13758 = new_n13757 ^ new_n13705;
  assign new_n13759 = new_n13758 ^ new_n13754;
  assign new_n13760 = new_n13726 ^ new_n13623;
  assign new_n13761 = new_n13720 ^ new_n13624;
  assign new_n13762 = ~new_n13760 & ~new_n13761;
  assign new_n13763 = new_n13762 ^ new_n13654;
  assign new_n13764 = new_n13756 ^ new_n13732;
  assign new_n13765 = new_n13764 ^ new_n13763;
  assign new_n13766 = ~new_n13759 & ~new_n13765;
  assign new_n13767 = new_n13762 ^ new_n13722;
  assign new_n13768 = new_n13767 ^ new_n13720;
  assign new_n13769 = new_n13768 ^ new_n13758;
  assign new_n13770 = new_n13769 ^ new_n13766;
  assign new_n13771 = ~new_n13625 & new_n13770;
  assign new_n13772 = new_n13653 ^ new_n13558;
  assign new_n13773 = new_n13746 ^ new_n13655;
  assign new_n13774 = new_n13720 ^ new_n13558;
  assign new_n13775 = new_n13751 ^ new_n13746;
  assign new_n13776 = new_n13775 ^ new_n13764;
  assign new_n13777 = new_n13776 ^ new_n13774;
  assign new_n13778 = new_n13769 ^ new_n13750;
  assign new_n13779 = ~new_n13777 & new_n13778;
  assign new_n13780 = new_n13779 ^ new_n13753;
  assign new_n13781 = new_n13780 ^ new_n13758;
  assign new_n13782 = new_n13766 ^ new_n13750;
  assign new_n13783 = ~new_n13782 & new_n13769;
  assign new_n13784 = new_n13783 ^ new_n13750;
  assign new_n13785 = ~new_n13781 & new_n13784;
  assign new_n13786 = new_n13783 ^ new_n13769;
  assign new_n13787 = new_n13786 ^ new_n13785;
  assign new_n13788 = new_n13787 ^ new_n13773;
  assign new_n13789 = new_n13788 ^ new_n13772;
  assign new_n13790 = new_n13789 ^ new_n13479;
  assign new_n13791 = new_n13779 ^ new_n13722;
  assign new_n13792 = new_n13791 ^ new_n13741;
  assign new_n13793 = new_n13792 ^ new_n13790;
  assign new_n13794 = ~new_n13793 & new_n13730;
  assign new_n13795 = new_n13785 ^ new_n13779;
  assign new_n13796 = new_n13795 ^ new_n13749;
  assign new_n13797 = new_n13705 & new_n13796;
  assign new_n13798 = new_n13785 ^ new_n13777;
  assign new_n13799 = ~new_n13624 & ~new_n13798;
  assign new_n13800 = ~new_n13731 & ~new_n13793;
  assign new_n13801 = new_n13779 ^ new_n13766;
  assign new_n13802 = new_n13768 ^ new_n13753;
  assign new_n13803 = new_n13802 ^ new_n13801;
  assign new_n13804 = ~new_n13803 & new_n13727;
  assign new_n13805 = new_n13804 ^ new_n13800;
  assign new_n13806 = new_n13786 ^ new_n13766;
  assign new_n13807 = new_n13806 ^ new_n13765;
  assign new_n13808 = ~new_n13745 & ~new_n13807;
  assign new_n13809 = new_n13808 ^ new_n13805;
  assign new_n13810 = new_n13809 ^ new_n13799;
  assign new_n13811 = new_n13810 ^ new_n13797;
  assign new_n13812 = new_n13811 ^ new_n13794;
  assign new_n13813 = new_n13812 ^ new_n13771;
  assign new_n13814 = new_n13766 ^ new_n13720;
  assign new_n13815 = new_n13762 ^ new_n13751;
  assign new_n13816 = new_n13815 ^ new_n13789;
  assign new_n13817 = new_n13816 ^ new_n13814;
  assign new_n13818 = new_n13755 & new_n13817;
  assign new_n13819 = ~new_n13761 & ~new_n13781;
  assign new_n13820 = new_n13819 ^ new_n13818;
  assign new_n13821 = ~new_n13721 & new_n13796;
  assign new_n13822 = ~new_n13623 & new_n13770;
  assign new_n13823 = new_n13786 ^ new_n13736;
  assign new_n13824 = ~new_n13823 & new_n13737;
  assign new_n13825 = new_n13824 ^ new_n13822;
  assign new_n13826 = new_n13825 ^ new_n13821;
  assign new_n13827 = new_n13826 ^ new_n13820;
  assign new_n13828 = new_n13827 ^ new_n13813;
  assign new_n13829 = new_n13828 ^ new_n12757;
  assign new_n13830 = new_n11424 ^ n8;
  assign new_n13831 = new_n10299 ^ n3;
  assign new_n13832 = new_n11407 ^ n2;
  assign new_n13833 = new_n13832 ^ new_n13831;
  assign new_n13834 = ~new_n13830 & ~new_n13833;
  assign new_n13835 = new_n11464 ^ n4;
  assign new_n13836 = new_n13830 & new_n13835;
  assign new_n13837 = new_n13836 ^ new_n13834;
  assign new_n13838 = new_n11559 ^ n1;
  assign new_n13839 = new_n13838 ^ new_n13835;
  assign new_n13840 = new_n11536 ^ n7;
  assign new_n13841 = new_n11503 ^ n5;
  assign new_n13842 = new_n13841 ^ new_n13840;
  assign new_n13843 = new_n13842 ^ new_n13839;
  assign new_n13844 = new_n13840 ^ new_n13835;
  assign new_n13845 = new_n11581 ^ n6;
  assign new_n13846 = new_n13845 ^ new_n13838;
  assign new_n13847 = new_n13846 ^ new_n13844;
  assign new_n13848 = ~new_n13843 & ~new_n13847;
  assign new_n13849 = new_n13848 ^ new_n13832;
  assign new_n13850 = new_n13849 ^ new_n13837;
  assign new_n13851 = new_n13833 ^ new_n13830;
  assign new_n13852 = new_n13840 & new_n13851;
  assign new_n13853 = new_n13852 ^ new_n13840;
  assign new_n13854 = new_n13845 ^ new_n13842;
  assign new_n13855 = new_n13854 ^ new_n13831;
  assign new_n13856 = new_n13840 ^ new_n13838;
  assign new_n13857 = ~new_n13856 & new_n13855;
  assign new_n13858 = new_n13857 ^ new_n13853;
  assign new_n13859 = new_n13858 ^ new_n13846;
  assign new_n13860 = new_n13835 ^ new_n13831;
  assign new_n13861 = new_n13860 ^ new_n13846;
  assign new_n13862 = new_n13845 ^ new_n13835;
  assign new_n13863 = ~new_n13861 & new_n13862;
  assign new_n13864 = new_n13854 ^ new_n13832;
  assign new_n13865 = new_n13839 & new_n13864;
  assign new_n13866 = new_n13865 ^ new_n13863;
  assign new_n13867 = new_n13841 ^ new_n13831;
  assign new_n13868 = new_n13867 ^ new_n13866;
  assign new_n13869 = new_n13868 ^ new_n13859;
  assign new_n13870 = new_n13849 ^ new_n13843;
  assign new_n13871 = new_n13851 ^ new_n13840;
  assign new_n13872 = new_n13871 ^ new_n13846;
  assign new_n13873 = new_n13843 ^ new_n13830;
  assign new_n13874 = new_n13872 & new_n13873;
  assign new_n13875 = new_n13874 ^ new_n13845;
  assign new_n13876 = new_n13875 ^ new_n13866;
  assign new_n13877 = new_n13876 ^ new_n13870;
  assign new_n13878 = ~new_n13869 & new_n13877;
  assign new_n13879 = new_n13878 ^ new_n13850;
  assign new_n13880 = new_n13843 ^ new_n13833;
  assign new_n13881 = ~new_n13880 & new_n13846;
  assign new_n13882 = new_n13881 ^ new_n13865;
  assign new_n13883 = new_n13882 ^ new_n13855;
  assign new_n13884 = new_n13883 ^ new_n13879;
  assign new_n13885 = new_n13864 ^ new_n13830;
  assign new_n13886 = new_n13851 ^ new_n13838;
  assign new_n13887 = ~new_n13885 & ~new_n13886;
  assign new_n13888 = new_n13887 ^ new_n13852;
  assign new_n13889 = new_n13881 ^ new_n13863;
  assign new_n13890 = new_n13889 ^ new_n13888;
  assign new_n13891 = ~new_n13884 & ~new_n13890;
  assign new_n13892 = new_n13887 ^ new_n13857;
  assign new_n13893 = new_n13892 ^ new_n13838;
  assign new_n13894 = new_n13893 ^ new_n13883;
  assign new_n13895 = new_n13894 ^ new_n13891;
  assign new_n13896 = new_n13851 ^ new_n13835;
  assign new_n13897 = ~new_n13896 & new_n13895;
  assign new_n13898 = new_n13838 ^ new_n13831;
  assign new_n13899 = new_n13837 ^ new_n13835;
  assign new_n13900 = new_n13899 ^ new_n13874;
  assign new_n13901 = new_n13900 ^ new_n13889;
  assign new_n13902 = new_n13901 ^ new_n13898;
  assign new_n13903 = new_n13894 ^ new_n13878;
  assign new_n13904 = ~new_n13902 & new_n13903;
  assign new_n13905 = new_n13904 ^ new_n13850;
  assign new_n13906 = new_n13905 ^ new_n13883;
  assign new_n13907 = new_n13891 ^ new_n13878;
  assign new_n13908 = ~new_n13907 & new_n13894;
  assign new_n13909 = new_n13908 ^ new_n13878;
  assign new_n13910 = ~new_n13906 & new_n13909;
  assign new_n13911 = new_n13910 ^ new_n13902;
  assign new_n13912 = ~new_n13851 & ~new_n13911;
  assign new_n13913 = new_n13908 ^ new_n13894;
  assign new_n13914 = new_n13913 ^ new_n13891;
  assign new_n13915 = new_n13914 ^ new_n13890;
  assign new_n13916 = ~new_n13915 & new_n13872;
  assign new_n13917 = new_n13840 ^ new_n13831;
  assign new_n13918 = new_n13874 ^ new_n13853;
  assign new_n13919 = new_n13913 ^ new_n13910;
  assign new_n13920 = new_n13919 ^ new_n13918;
  assign new_n13921 = new_n13920 ^ new_n13917;
  assign new_n13922 = new_n13921 ^ new_n13835;
  assign new_n13923 = new_n13904 ^ new_n13857;
  assign new_n13924 = new_n13923 ^ new_n13849;
  assign new_n13925 = new_n13924 ^ new_n13922;
  assign new_n13926 = ~new_n13925 & new_n13862;
  assign new_n13927 = new_n13904 ^ new_n13891;
  assign new_n13928 = new_n13893 ^ new_n13850;
  assign new_n13929 = new_n13928 ^ new_n13927;
  assign new_n13930 = ~new_n13929 & new_n13839;
  assign new_n13931 = new_n13930 ^ new_n13926;
  assign new_n13932 = new_n13931 ^ new_n13916;
  assign new_n13933 = new_n13932 ^ new_n13912;
  assign new_n13934 = new_n13910 ^ new_n13904;
  assign new_n13935 = new_n13934 ^ new_n13877;
  assign new_n13936 = new_n13855 & new_n13935;
  assign new_n13937 = new_n13936 ^ new_n13933;
  assign new_n13938 = ~new_n13861 & ~new_n13925;
  assign new_n13939 = new_n13938 ^ new_n13937;
  assign new_n13940 = new_n13939 ^ new_n13897;
  assign new_n13941 = new_n13891 ^ new_n13838;
  assign new_n13942 = new_n13899 ^ new_n13887;
  assign new_n13943 = new_n13942 ^ new_n13921;
  assign new_n13944 = new_n13943 ^ new_n13941;
  assign new_n13945 = ~new_n13880 & new_n13944;
  assign new_n13946 = ~new_n13886 & ~new_n13906;
  assign new_n13947 = new_n13946 ^ new_n13945;
  assign new_n13948 = ~new_n13856 & new_n13935;
  assign new_n13949 = ~new_n13830 & new_n13895;
  assign new_n13950 = new_n13913 ^ new_n13869;
  assign new_n13951 = ~new_n13843 & ~new_n13950;
  assign new_n13952 = new_n13951 ^ new_n13949;
  assign new_n13953 = new_n13952 ^ new_n13948;
  assign new_n13954 = new_n13953 ^ new_n13947;
  assign new_n13955 = new_n13954 ^ new_n13940;
  assign new_n13956 = new_n11738 ^ n2;
  assign new_n13957 = new_n11732 ^ n3;
  assign new_n13958 = new_n13957 ^ new_n13956;
  assign new_n13959 = new_n11754 ^ n8;
  assign new_n13960 = new_n13959 ^ new_n13958;
  assign new_n13961 = new_n11693 ^ n4;
  assign new_n13962 = new_n13961 ^ new_n13960;
  assign new_n13963 = ~new_n13959 & ~new_n13962;
  assign new_n13964 = new_n13963 ^ new_n13961;
  assign new_n13965 = new_n11710 ^ n7;
  assign new_n13966 = new_n13965 ^ new_n13961;
  assign new_n13967 = new_n11702 ^ n1;
  assign new_n13968 = new_n11725 ^ n6;
  assign new_n13969 = new_n13968 ^ new_n13967;
  assign new_n13970 = new_n13969 ^ new_n13966;
  assign new_n13971 = new_n13967 ^ new_n13961;
  assign new_n13972 = new_n11717 ^ n5;
  assign new_n13973 = new_n13972 ^ new_n13965;
  assign new_n13974 = new_n13973 ^ new_n13971;
  assign new_n13975 = ~new_n13970 & ~new_n13974;
  assign new_n13976 = new_n13975 ^ new_n13956;
  assign new_n13977 = new_n13976 ^ new_n13964;
  assign new_n13978 = new_n13960 & new_n13965;
  assign new_n13979 = new_n13978 ^ new_n13965;
  assign new_n13980 = new_n13973 ^ new_n13968;
  assign new_n13981 = new_n13980 ^ new_n13957;
  assign new_n13982 = new_n13967 ^ new_n13965;
  assign new_n13983 = ~new_n13982 & new_n13981;
  assign new_n13984 = new_n13983 ^ new_n13979;
  assign new_n13985 = new_n13984 ^ new_n13969;
  assign new_n13986 = new_n13961 ^ new_n13957;
  assign new_n13987 = new_n13986 ^ new_n13969;
  assign new_n13988 = new_n13968 ^ new_n13961;
  assign new_n13989 = ~new_n13987 & new_n13988;
  assign new_n13990 = new_n13980 ^ new_n13956;
  assign new_n13991 = new_n13971 & new_n13990;
  assign new_n13992 = new_n13991 ^ new_n13989;
  assign new_n13993 = new_n13972 ^ new_n13957;
  assign new_n13994 = new_n13993 ^ new_n13992;
  assign new_n13995 = new_n13994 ^ new_n13985;
  assign new_n13996 = new_n13976 ^ new_n13974;
  assign new_n13997 = new_n13974 ^ new_n13959;
  assign new_n13998 = new_n13965 ^ new_n13960;
  assign new_n13999 = new_n13998 ^ new_n13969;
  assign new_n14000 = new_n13997 & new_n13999;
  assign new_n14001 = new_n14000 ^ new_n13968;
  assign new_n14002 = new_n14001 ^ new_n13992;
  assign new_n14003 = new_n14002 ^ new_n13996;
  assign new_n14004 = ~new_n13995 & new_n14003;
  assign new_n14005 = new_n14004 ^ new_n13977;
  assign new_n14006 = new_n13974 ^ new_n13958;
  assign new_n14007 = ~new_n14006 & new_n13969;
  assign new_n14008 = new_n14007 ^ new_n13991;
  assign new_n14009 = new_n14008 ^ new_n13981;
  assign new_n14010 = new_n14009 ^ new_n14005;
  assign new_n14011 = new_n13990 ^ new_n13959;
  assign new_n14012 = new_n13967 ^ new_n13960;
  assign new_n14013 = ~new_n14011 & ~new_n14012;
  assign new_n14014 = new_n14013 ^ new_n13978;
  assign new_n14015 = new_n14007 ^ new_n13989;
  assign new_n14016 = new_n14015 ^ new_n14014;
  assign new_n14017 = ~new_n14010 & ~new_n14016;
  assign new_n14018 = new_n14013 ^ new_n13983;
  assign new_n14019 = new_n14018 ^ new_n13967;
  assign new_n14020 = new_n14019 ^ new_n14009;
  assign new_n14021 = new_n14020 ^ new_n14017;
  assign new_n14022 = ~new_n13962 & new_n14021;
  assign new_n14023 = new_n13965 ^ new_n13957;
  assign new_n14024 = new_n14000 ^ new_n13979;
  assign new_n14025 = new_n13967 ^ new_n13957;
  assign new_n14026 = new_n14000 ^ new_n13963;
  assign new_n14027 = new_n14026 ^ new_n14015;
  assign new_n14028 = new_n14027 ^ new_n14025;
  assign new_n14029 = new_n14020 ^ new_n14004;
  assign new_n14030 = ~new_n14028 & new_n14029;
  assign new_n14031 = new_n14030 ^ new_n13977;
  assign new_n14032 = new_n14031 ^ new_n14009;
  assign new_n14033 = new_n14017 ^ new_n14004;
  assign new_n14034 = ~new_n14033 & new_n14020;
  assign new_n14035 = new_n14034 ^ new_n14004;
  assign new_n14036 = ~new_n14032 & new_n14035;
  assign new_n14037 = new_n14034 ^ new_n14020;
  assign new_n14038 = new_n14037 ^ new_n14036;
  assign new_n14039 = new_n14038 ^ new_n14024;
  assign new_n14040 = new_n14039 ^ new_n14023;
  assign new_n14041 = new_n14040 ^ new_n13961;
  assign new_n14042 = new_n14030 ^ new_n13983;
  assign new_n14043 = new_n14042 ^ new_n13976;
  assign new_n14044 = new_n14043 ^ new_n14041;
  assign new_n14045 = ~new_n13987 & ~new_n14044;
  assign new_n14046 = new_n14036 ^ new_n14028;
  assign new_n14047 = ~new_n13960 & ~new_n14046;
  assign new_n14048 = new_n14037 ^ new_n14017;
  assign new_n14049 = new_n14048 ^ new_n14016;
  assign new_n14050 = ~new_n14049 & new_n13999;
  assign new_n14051 = ~new_n14044 & new_n13988;
  assign new_n14052 = new_n14030 ^ new_n14017;
  assign new_n14053 = new_n14019 ^ new_n13977;
  assign new_n14054 = new_n14053 ^ new_n14052;
  assign new_n14055 = ~new_n14054 & new_n13971;
  assign new_n14056 = new_n14055 ^ new_n14051;
  assign new_n14057 = new_n14056 ^ new_n14050;
  assign new_n14058 = new_n14057 ^ new_n14047;
  assign new_n14059 = new_n14036 ^ new_n14030;
  assign new_n14060 = new_n14059 ^ new_n14003;
  assign new_n14061 = new_n13981 & new_n14060;
  assign new_n14062 = new_n14061 ^ new_n14058;
  assign new_n14063 = new_n14062 ^ new_n14045;
  assign new_n14064 = new_n14063 ^ new_n14022;
  assign new_n14065 = ~new_n14012 & ~new_n14032;
  assign new_n14066 = new_n14017 ^ new_n13967;
  assign new_n14067 = new_n14013 ^ new_n13963;
  assign new_n14068 = new_n14067 ^ new_n14040;
  assign new_n14069 = new_n14068 ^ new_n14066;
  assign new_n14070 = ~new_n14006 & new_n14069;
  assign new_n14071 = new_n14070 ^ new_n14065;
  assign new_n14072 = ~new_n13959 & new_n14021;
  assign new_n14073 = new_n14037 ^ new_n13995;
  assign new_n14074 = ~new_n13974 & ~new_n14073;
  assign new_n14075 = new_n14074 ^ new_n14072;
  assign new_n14076 = ~new_n13982 & new_n14060;
  assign new_n14077 = new_n14076 ^ new_n14075;
  assign new_n14078 = new_n14077 ^ new_n14071;
  assign new_n14079 = new_n14078 ^ new_n14064;
  assign new_n14080 = new_n14079 ^ new_n13955;
  assign new_n14081 = new_n14080 ^ new_n903;
  assign new_n14082 = new_n11689 ^ new_n11683;
  assign new_n14083 = new_n11675 ^ new_n11649;
  assign new_n14084 = ~new_n11624 & ~new_n11643;
  assign new_n14085 = ~new_n11648 & new_n11611;
  assign new_n14086 = new_n14085 ^ new_n14084;
  assign new_n14087 = new_n14086 ^ new_n11668;
  assign new_n14088 = new_n14087 ^ new_n14083;
  assign new_n14089 = new_n14088 ^ new_n14082;
  assign new_n14090 = ~new_n14054 & new_n13990;
  assign new_n14091 = new_n14090 ^ new_n14045;
  assign new_n14092 = ~new_n14049 & new_n13997;
  assign new_n14093 = new_n14092 ^ new_n14074;
  assign new_n14094 = ~new_n13970 & ~new_n14073;
  assign new_n14095 = new_n14094 ^ new_n14093;
  assign new_n14096 = new_n14095 ^ new_n14057;
  assign new_n14097 = new_n14096 ^ new_n14091;
  assign new_n14098 = new_n14097 ^ new_n12902;
  assign new_n14099 = new_n7861 ^ new_n1117;
  assign new_n14100 = new_n14099 ^ new_n10077;
  assign new_n14101 = new_n13060 ^ new_n9996;
  assign new_n14102 = new_n14101 ^ new_n14100;
  assign new_n14103 = new_n1200 ^ new_n713;
  assign new_n14104 = new_n14103 ^ new_n9474;
  assign new_n14105 = new_n13025 ^ new_n9960;
  assign new_n14106 = new_n14105 ^ new_n14104;
  assign new_n14107 = new_n13078 ^ new_n9901;
  assign new_n14108 = new_n7787 ^ new_n1181;
  assign new_n14109 = new_n14108 ^ new_n9964;
  assign new_n14110 = new_n14109 ^ new_n13032;
  assign new_n14111 = new_n14110 ^ new_n14107;
  assign new_n14112 = new_n7822 ^ new_n1173;
  assign new_n14113 = new_n14112 ^ new_n10069;
  assign new_n14114 = new_n14113 ^ new_n13032;
  assign new_n14115 = new_n13047 ^ new_n9851;
  assign new_n14116 = new_n14115 ^ new_n14114;
  assign new_n14117 = new_n14116 ^ new_n14111;
  assign new_n14118 = new_n14117 ^ new_n14106;
  assign new_n14119 = new_n14118 ^ new_n14102;
  assign new_n14120 = new_n7937 ^ new_n1189;
  assign new_n14121 = new_n14120 ^ new_n9859;
  assign new_n14122 = new_n13054 ^ new_n10082;
  assign new_n14123 = new_n14122 ^ new_n14121;
  assign new_n14124 = new_n13021 ^ new_n10062;
  assign new_n14125 = new_n7965 ^ new_n1162;
  assign new_n14126 = new_n14125 ^ new_n10052;
  assign new_n14127 = new_n14126 ^ new_n13032;
  assign new_n14128 = new_n14127 ^ new_n14124;
  assign new_n14129 = new_n14128 ^ new_n14123;
  assign new_n14130 = new_n14129 ^ new_n14117;
  assign new_n14131 = new_n14128 ^ new_n14111;
  assign new_n14132 = new_n14123 ^ new_n14106;
  assign new_n14133 = new_n14132 ^ new_n14131;
  assign new_n14134 = ~new_n14130 & ~new_n14133;
  assign new_n14135 = new_n14134 ^ new_n14102;
  assign new_n14136 = new_n7896 ^ new_n1153;
  assign new_n14137 = new_n14136 ^ new_n9868;
  assign new_n14138 = new_n13032 ^ new_n10030;
  assign new_n14139 = new_n14138 ^ new_n14137;
  assign new_n14140 = new_n7910 ^ new_n1140;
  assign new_n14141 = new_n14140 ^ new_n10000;
  assign new_n14142 = new_n13039 ^ new_n10041;
  assign new_n14143 = new_n14142 ^ new_n14141;
  assign new_n14144 = new_n14143 ^ new_n14102;
  assign new_n14145 = ~new_n14139 & ~new_n14144;
  assign new_n14146 = new_n14128 & new_n14139;
  assign new_n14147 = new_n14146 ^ new_n14145;
  assign new_n14148 = new_n14147 ^ new_n14135;
  assign new_n14149 = new_n14144 ^ new_n14139;
  assign new_n14150 = new_n14111 & new_n14149;
  assign new_n14151 = new_n14150 ^ new_n14111;
  assign new_n14152 = new_n14143 ^ new_n14118;
  assign new_n14153 = new_n14123 ^ new_n14111;
  assign new_n14154 = ~new_n14153 & new_n14152;
  assign new_n14155 = new_n14154 ^ new_n14151;
  assign new_n14156 = new_n14155 ^ new_n14132;
  assign new_n14157 = new_n14119 & new_n14129;
  assign new_n14158 = new_n14143 ^ new_n14128;
  assign new_n14159 = new_n14158 ^ new_n14132;
  assign new_n14160 = new_n14128 ^ new_n14106;
  assign new_n14161 = ~new_n14159 & new_n14160;
  assign new_n14162 = new_n14161 ^ new_n14157;
  assign new_n14163 = new_n14143 ^ new_n14116;
  assign new_n14164 = new_n14163 ^ new_n14162;
  assign new_n14165 = new_n14164 ^ new_n14156;
  assign new_n14166 = new_n14135 ^ new_n14130;
  assign new_n14167 = new_n14139 ^ new_n14130;
  assign new_n14168 = new_n14149 ^ new_n14111;
  assign new_n14169 = new_n14168 ^ new_n14132;
  assign new_n14170 = new_n14167 & new_n14169;
  assign new_n14171 = new_n14170 ^ new_n14157;
  assign new_n14172 = new_n14161 ^ new_n14106;
  assign new_n14173 = new_n14172 ^ new_n14171;
  assign new_n14174 = new_n14173 ^ new_n14166;
  assign new_n14175 = ~new_n14165 & new_n14174;
  assign new_n14176 = new_n14175 ^ new_n14148;
  assign new_n14177 = new_n14144 ^ new_n14130;
  assign new_n14178 = ~new_n14177 & new_n14132;
  assign new_n14179 = new_n14178 ^ new_n14157;
  assign new_n14180 = new_n14179 ^ new_n14152;
  assign new_n14181 = new_n14180 ^ new_n14176;
  assign new_n14182 = new_n14149 ^ new_n14123;
  assign new_n14183 = new_n14139 ^ new_n14119;
  assign new_n14184 = ~new_n14182 & ~new_n14183;
  assign new_n14185 = new_n14184 ^ new_n14150;
  assign new_n14186 = new_n14178 ^ new_n14161;
  assign new_n14187 = new_n14186 ^ new_n14185;
  assign new_n14188 = ~new_n14181 & ~new_n14187;
  assign new_n14189 = new_n14143 ^ new_n14123;
  assign new_n14190 = new_n14147 ^ new_n14128;
  assign new_n14191 = new_n14190 ^ new_n14170;
  assign new_n14192 = new_n14191 ^ new_n14186;
  assign new_n14193 = new_n14192 ^ new_n14189;
  assign new_n14194 = new_n14184 ^ new_n14154;
  assign new_n14195 = new_n14194 ^ new_n14123;
  assign new_n14196 = new_n14195 ^ new_n14180;
  assign new_n14197 = new_n14196 ^ new_n14175;
  assign new_n14198 = ~new_n14193 & new_n14197;
  assign new_n14199 = new_n14198 ^ new_n14188;
  assign new_n14200 = new_n14195 ^ new_n14148;
  assign new_n14201 = new_n14200 ^ new_n14199;
  assign new_n14202 = ~new_n14201 & new_n14119;
  assign new_n14203 = new_n14143 ^ new_n14111;
  assign new_n14204 = new_n14170 ^ new_n14151;
  assign new_n14205 = new_n14198 ^ new_n14148;
  assign new_n14206 = new_n14205 ^ new_n14180;
  assign new_n14207 = new_n14188 ^ new_n14175;
  assign new_n14208 = new_n14196 & new_n14207;
  assign new_n14209 = new_n14208 ^ new_n14197;
  assign new_n14210 = ~new_n14206 & new_n14209;
  assign new_n14211 = new_n14210 ^ new_n14208;
  assign new_n14212 = new_n14211 ^ new_n14204;
  assign new_n14213 = new_n14212 ^ new_n14203;
  assign new_n14214 = new_n14213 ^ new_n14128;
  assign new_n14215 = new_n14198 ^ new_n14154;
  assign new_n14216 = new_n14215 ^ new_n14135;
  assign new_n14217 = new_n14216 ^ new_n14214;
  assign new_n14218 = ~new_n14159 & ~new_n14217;
  assign new_n14219 = new_n14218 ^ new_n14202;
  assign new_n14220 = new_n14208 ^ new_n14188;
  assign new_n14221 = new_n14220 ^ new_n14187;
  assign new_n14222 = ~new_n14221 & new_n14167;
  assign new_n14223 = new_n14208 ^ new_n14165;
  assign new_n14224 = ~new_n14130 & ~new_n14223;
  assign new_n14225 = new_n14224 ^ new_n14222;
  assign new_n14226 = ~new_n14133 & ~new_n14223;
  assign new_n14227 = new_n14226 ^ new_n14225;
  assign new_n14228 = ~new_n14221 & new_n14169;
  assign new_n14229 = ~new_n14201 & new_n14129;
  assign new_n14230 = ~new_n14217 & new_n14160;
  assign new_n14231 = new_n14230 ^ new_n14229;
  assign new_n14232 = new_n14231 ^ new_n14228;
  assign new_n14233 = new_n14232 ^ new_n14227;
  assign new_n14234 = new_n14233 ^ new_n14219;
  assign new_n14235 = new_n14234 ^ new_n14098;
  assign new_n14236 = new_n7850 ^ new_n6837;
  assign new_n14237 = new_n14236 ^ new_n4899;
  assign new_n14238 = new_n8352 ^ new_n605;
  assign new_n14239 = new_n14238 ^ new_n7766;
  assign new_n14240 = new_n14239 ^ new_n14237;
  assign new_n14241 = new_n7962 ^ new_n7838;
  assign new_n14242 = new_n14241 ^ new_n7830;
  assign new_n14243 = new_n8931 ^ new_n597;
  assign new_n14244 = new_n14243 ^ new_n7945;
  assign new_n14245 = new_n14244 ^ new_n6838;
  assign new_n14246 = new_n14245 ^ new_n14242;
  assign new_n14247 = new_n7945 ^ new_n7746;
  assign new_n14248 = new_n14247 ^ new_n7904;
  assign new_n14249 = new_n8904 ^ new_n591;
  assign new_n14250 = new_n14249 ^ new_n7797;
  assign new_n14251 = new_n14250 ^ new_n7765;
  assign new_n14252 = new_n14251 ^ new_n14248;
  assign new_n14253 = new_n14252 ^ new_n14246;
  assign new_n14254 = new_n14253 ^ new_n14240;
  assign new_n14255 = new_n7948 ^ new_n7922;
  assign new_n14256 = new_n8985 ^ new_n566;
  assign new_n14257 = new_n14256 ^ new_n7869;
  assign new_n14258 = new_n14257 ^ new_n7881;
  assign new_n14259 = new_n14258 ^ new_n14255;
  assign new_n14260 = new_n14259 ^ new_n14254;
  assign new_n14261 = new_n7958 ^ new_n7890;
  assign new_n14262 = new_n9024 ^ new_n560;
  assign new_n14263 = new_n14262 ^ new_n7916;
  assign new_n14264 = new_n14263 ^ new_n7921;
  assign new_n14265 = new_n14264 ^ new_n14261;
  assign new_n14266 = new_n14265 ^ new_n14259;
  assign new_n14267 = new_n7945 ^ new_n7777;
  assign new_n14268 = new_n9001 ^ new_n575;
  assign new_n14269 = new_n14268 ^ new_n7900;
  assign new_n14270 = new_n14269 ^ new_n7903;
  assign new_n14271 = new_n14270 ^ new_n14267;
  assign new_n14272 = new_n14271 ^ new_n14266;
  assign new_n14273 = new_n14252 & new_n14272;
  assign new_n14274 = new_n14273 ^ new_n14252;
  assign new_n14275 = new_n9044 ^ new_n584;
  assign new_n14276 = new_n14275 ^ new_n7882;
  assign new_n14277 = new_n13183 ^ new_n7944;
  assign new_n14278 = new_n14277 ^ new_n14276;
  assign new_n14279 = new_n14278 ^ new_n14252;
  assign new_n14280 = new_n14265 ^ new_n14254;
  assign new_n14281 = ~new_n14279 & new_n14280;
  assign new_n14282 = new_n14281 ^ new_n14274;
  assign new_n14283 = new_n14278 ^ new_n14240;
  assign new_n14284 = new_n14283 ^ new_n14282;
  assign new_n14285 = new_n9065 ^ new_n540;
  assign new_n14286 = new_n14285 ^ new_n7945;
  assign new_n14287 = new_n14286 ^ new_n7844;
  assign new_n14288 = new_n13203 ^ new_n7957;
  assign new_n14289 = new_n14288 ^ new_n14287;
  assign new_n14290 = new_n14289 ^ new_n14240;
  assign new_n14291 = new_n14289 ^ new_n14265;
  assign new_n14292 = new_n14291 ^ new_n14283;
  assign new_n14293 = ~new_n14292 & new_n14290;
  assign new_n14294 = new_n14289 ^ new_n14278;
  assign new_n14295 = new_n14260 & new_n14294;
  assign new_n14296 = new_n14295 ^ new_n14293;
  assign new_n14297 = new_n14265 ^ new_n14246;
  assign new_n14298 = new_n14297 ^ new_n14296;
  assign new_n14299 = new_n14298 ^ new_n14284;
  assign new_n14300 = new_n14294 ^ new_n14253;
  assign new_n14301 = new_n14290 ^ new_n14279;
  assign new_n14302 = ~new_n14300 & ~new_n14301;
  assign new_n14303 = new_n14302 ^ new_n14259;
  assign new_n14304 = new_n14303 ^ new_n14300;
  assign new_n14305 = new_n14300 ^ new_n14271;
  assign new_n14306 = new_n14272 ^ new_n14252;
  assign new_n14307 = new_n14306 ^ new_n14283;
  assign new_n14308 = new_n14305 & new_n14307;
  assign new_n14309 = new_n14308 ^ new_n14295;
  assign new_n14310 = new_n14293 ^ new_n14240;
  assign new_n14311 = new_n14310 ^ new_n14309;
  assign new_n14312 = new_n14311 ^ new_n14304;
  assign new_n14313 = ~new_n14299 & new_n14312;
  assign new_n14314 = new_n14300 ^ new_n14266;
  assign new_n14315 = ~new_n14314 & new_n14283;
  assign new_n14316 = new_n14315 ^ new_n14295;
  assign new_n14317 = new_n14316 ^ new_n14280;
  assign new_n14318 = new_n14278 ^ new_n14272;
  assign new_n14319 = new_n14271 ^ new_n14260;
  assign new_n14320 = ~new_n14318 & ~new_n14319;
  assign new_n14321 = new_n14320 ^ new_n14281;
  assign new_n14322 = new_n14321 ^ new_n14278;
  assign new_n14323 = new_n14322 ^ new_n14317;
  assign new_n14324 = new_n14323 ^ new_n14313;
  assign new_n14325 = new_n14278 ^ new_n14265;
  assign new_n14326 = new_n14289 ^ new_n14272;
  assign new_n14327 = ~new_n14271 & ~new_n14326;
  assign new_n14328 = new_n14327 ^ new_n14308;
  assign new_n14329 = new_n14315 ^ new_n14293;
  assign new_n14330 = new_n14329 ^ new_n14328;
  assign new_n14331 = new_n14330 ^ new_n14325;
  assign new_n14332 = ~new_n14331 & new_n14324;
  assign new_n14333 = new_n14327 ^ new_n14289;
  assign new_n14334 = new_n14333 ^ new_n14303;
  assign new_n14335 = new_n14334 ^ new_n14313;
  assign new_n14336 = new_n14335 ^ new_n14317;
  assign new_n14337 = new_n14320 ^ new_n14273;
  assign new_n14338 = new_n14337 ^ new_n14329;
  assign new_n14339 = ~new_n14336 & ~new_n14338;
  assign new_n14340 = new_n14339 ^ new_n14332;
  assign new_n14341 = new_n14334 ^ new_n14322;
  assign new_n14342 = new_n14341 ^ new_n14340;
  assign new_n14343 = ~new_n14342 & new_n14260;
  assign new_n14344 = ~new_n14342 & new_n14294;
  assign new_n14345 = new_n14344 ^ new_n14343;
  assign new_n14346 = new_n14339 ^ new_n14278;
  assign new_n14347 = new_n14327 ^ new_n14320;
  assign new_n14348 = new_n14265 ^ new_n14252;
  assign new_n14349 = new_n14308 ^ new_n14274;
  assign new_n14350 = new_n14339 ^ new_n14313;
  assign new_n14351 = ~new_n14323 & ~new_n14350;
  assign new_n14352 = new_n14351 ^ new_n14339;
  assign new_n14353 = new_n14334 ^ new_n14332;
  assign new_n14354 = new_n14353 ^ new_n14317;
  assign new_n14355 = ~new_n14352 & ~new_n14354;
  assign new_n14356 = new_n14352 ^ new_n14324;
  assign new_n14357 = new_n14356 ^ new_n14355;
  assign new_n14358 = new_n14357 ^ new_n14349;
  assign new_n14359 = new_n14358 ^ new_n14348;
  assign new_n14360 = new_n14359 ^ new_n14347;
  assign new_n14361 = new_n14360 ^ new_n14346;
  assign new_n14362 = ~new_n14361 & new_n14283;
  assign new_n14363 = ~new_n14318 & ~new_n14354;
  assign new_n14364 = ~new_n14314 & ~new_n14361;
  assign new_n14365 = new_n14364 ^ new_n14363;
  assign new_n14366 = new_n14339 ^ new_n14323;
  assign new_n14367 = ~new_n14271 & new_n14366;
  assign new_n14368 = new_n14356 ^ new_n14299;
  assign new_n14369 = ~new_n14300 & new_n14368;
  assign new_n14370 = new_n14369 ^ new_n14367;
  assign new_n14371 = new_n14355 ^ new_n14332;
  assign new_n14372 = new_n14371 ^ new_n14312;
  assign new_n14373 = ~new_n14279 & new_n14372;
  assign new_n14374 = new_n14373 ^ new_n14370;
  assign new_n14375 = new_n14374 ^ new_n14365;
  assign new_n14376 = new_n14375 ^ new_n14362;
  assign new_n14377 = new_n14376 ^ new_n14345;
  assign new_n14378 = new_n13340 ^ new_n8961;
  assign new_n14379 = new_n13956 ^ new_n8993;
  assign new_n14380 = new_n14379 ^ new_n9030;
  assign new_n14381 = new_n14380 ^ new_n14378;
  assign new_n14382 = new_n9050 ^ new_n8885;
  assign new_n14383 = new_n14382 ^ new_n13972;
  assign new_n14384 = new_n14383 ^ new_n8702;
  assign new_n14385 = new_n13363 ^ new_n8947;
  assign new_n14386 = new_n14385 ^ new_n14384;
  assign new_n14387 = new_n14382 ^ new_n8867;
  assign new_n14388 = new_n14387 ^ new_n9006;
  assign new_n14389 = new_n13965 ^ new_n8848;
  assign new_n14390 = new_n14389 ^ new_n8895;
  assign new_n14391 = new_n14390 ^ new_n14388;
  assign new_n14392 = new_n14391 ^ new_n14386;
  assign new_n14393 = new_n13968 ^ new_n8868;
  assign new_n14394 = new_n8939 ^ new_n8701;
  assign new_n14395 = new_n14394 ^ new_n8224;
  assign new_n14396 = new_n14395 ^ new_n14393;
  assign new_n14397 = new_n14396 ^ new_n14392;
  assign new_n14398 = new_n14397 ^ new_n14381;
  assign new_n14399 = new_n14382 ^ new_n9005;
  assign new_n14400 = new_n13959 ^ new_n8915;
  assign new_n14401 = new_n14400 ^ new_n8998;
  assign new_n14402 = new_n14401 ^ new_n14399;
  assign new_n14403 = new_n14382 ^ new_n13347;
  assign new_n14404 = new_n13961 ^ new_n9069;
  assign new_n14405 = new_n14404 ^ new_n8953;
  assign new_n14406 = new_n14405 ^ new_n14403;
  assign new_n14407 = new_n13335 ^ new_n9030;
  assign new_n14408 = new_n13957 ^ new_n9070;
  assign new_n14409 = new_n14408 ^ new_n14407;
  assign new_n14410 = new_n14409 ^ new_n14381;
  assign new_n14411 = new_n14410 ^ new_n14402;
  assign new_n14412 = new_n14411 ^ new_n14406;
  assign new_n14413 = new_n14402 & new_n14412;
  assign new_n14414 = new_n14413 ^ new_n14406;
  assign new_n14415 = new_n13319 ^ new_n8971;
  assign new_n14416 = new_n13967 ^ new_n9050;
  assign new_n14417 = new_n14416 ^ new_n8993;
  assign new_n14418 = new_n14417 ^ new_n14415;
  assign new_n14419 = new_n14418 ^ new_n14406;
  assign new_n14420 = new_n14419 ^ new_n14392;
  assign new_n14421 = new_n14406 ^ new_n14391;
  assign new_n14422 = new_n14418 ^ new_n14396;
  assign new_n14423 = new_n14422 ^ new_n14421;
  assign new_n14424 = new_n14420 & new_n14423;
  assign new_n14425 = new_n14424 ^ new_n14381;
  assign new_n14426 = new_n14425 ^ new_n14414;
  assign new_n14427 = ~new_n14391 & ~new_n14411;
  assign new_n14428 = new_n14427 ^ new_n14391;
  assign new_n14429 = new_n14409 ^ new_n14397;
  assign new_n14430 = new_n14418 ^ new_n14391;
  assign new_n14431 = new_n14429 & new_n14430;
  assign new_n14432 = new_n14431 ^ new_n14428;
  assign new_n14433 = new_n14432 ^ new_n14422;
  assign new_n14434 = new_n14398 & new_n14419;
  assign new_n14435 = new_n14409 ^ new_n14406;
  assign new_n14436 = new_n14435 ^ new_n14422;
  assign new_n14437 = new_n14406 ^ new_n14396;
  assign new_n14438 = new_n14436 & new_n14437;
  assign new_n14439 = new_n14438 ^ new_n14434;
  assign new_n14440 = new_n14409 ^ new_n14386;
  assign new_n14441 = new_n14440 ^ new_n14439;
  assign new_n14442 = new_n14441 ^ new_n14433;
  assign new_n14443 = new_n14425 ^ new_n14420;
  assign new_n14444 = new_n14411 ^ new_n14391;
  assign new_n14445 = new_n14444 ^ new_n14422;
  assign new_n14446 = new_n14420 ^ new_n14402;
  assign new_n14447 = new_n14445 & new_n14446;
  assign new_n14448 = new_n14447 ^ new_n14439;
  assign new_n14449 = new_n14448 ^ new_n14396;
  assign new_n14450 = new_n14449 ^ new_n14443;
  assign new_n14451 = ~new_n14442 & new_n14450;
  assign new_n14452 = new_n14451 ^ new_n14426;
  assign new_n14453 = new_n14420 ^ new_n14410;
  assign new_n14454 = new_n14422 & new_n14453;
  assign new_n14455 = new_n14454 ^ new_n14434;
  assign new_n14456 = new_n14455 ^ new_n14429;
  assign new_n14457 = new_n14456 ^ new_n14452;
  assign new_n14458 = new_n14402 ^ new_n14398;
  assign new_n14459 = new_n14418 ^ new_n14411;
  assign new_n14460 = new_n14458 & new_n14459;
  assign new_n14461 = new_n14460 ^ new_n14427;
  assign new_n14462 = new_n14454 ^ new_n14438;
  assign new_n14463 = new_n14462 ^ new_n14461;
  assign new_n14464 = ~new_n14463 & new_n14457;
  assign new_n14465 = new_n14418 ^ new_n14409;
  assign new_n14466 = new_n14447 ^ new_n14413;
  assign new_n14467 = new_n14466 ^ new_n14462;
  assign new_n14468 = new_n14467 ^ new_n14465;
  assign new_n14469 = new_n14460 ^ new_n14431;
  assign new_n14470 = new_n14469 ^ new_n14418;
  assign new_n14471 = new_n14470 ^ new_n14456;
  assign new_n14472 = new_n14471 ^ new_n14451;
  assign new_n14473 = new_n14468 & new_n14472;
  assign new_n14474 = new_n14473 ^ new_n14464;
  assign new_n14475 = new_n14470 ^ new_n14426;
  assign new_n14476 = new_n14475 ^ new_n14474;
  assign new_n14477 = new_n14398 & new_n14476;
  assign new_n14478 = new_n14419 & new_n14476;
  assign new_n14479 = new_n14478 ^ new_n14477;
  assign new_n14480 = new_n14464 ^ new_n14418;
  assign new_n14481 = new_n14460 ^ new_n14413;
  assign new_n14482 = new_n14409 ^ new_n14391;
  assign new_n14483 = new_n14447 ^ new_n14428;
  assign new_n14484 = new_n14473 ^ new_n14426;
  assign new_n14485 = new_n14484 ^ new_n14456;
  assign new_n14486 = new_n14464 ^ new_n14451;
  assign new_n14487 = new_n14471 & new_n14486;
  assign new_n14488 = new_n14487 ^ new_n14472;
  assign new_n14489 = new_n14485 & new_n14488;
  assign new_n14490 = new_n14489 ^ new_n14487;
  assign new_n14491 = new_n14490 ^ new_n14483;
  assign new_n14492 = new_n14491 ^ new_n14482;
  assign new_n14493 = new_n14492 ^ new_n14481;
  assign new_n14494 = new_n14493 ^ new_n14480;
  assign new_n14495 = ~new_n14494 & new_n14422;
  assign new_n14496 = new_n14489 ^ new_n14473;
  assign new_n14497 = new_n14496 ^ new_n14450;
  assign new_n14498 = new_n14430 & new_n14497;
  assign new_n14499 = new_n14471 ^ new_n14464;
  assign new_n14500 = new_n14402 & new_n14499;
  assign new_n14501 = new_n14487 ^ new_n14442;
  assign new_n14502 = ~new_n14501 & new_n14420;
  assign new_n14503 = new_n14502 ^ new_n14500;
  assign new_n14504 = new_n14503 ^ new_n14498;
  assign new_n14505 = ~new_n14494 & new_n14453;
  assign new_n14506 = new_n14459 & new_n14485;
  assign new_n14507 = new_n14506 ^ new_n14505;
  assign new_n14508 = new_n14507 ^ new_n14504;
  assign new_n14509 = new_n14508 ^ new_n14495;
  assign new_n14510 = new_n14509 ^ new_n14479;
  assign new_n14511 = new_n14510 ^ new_n14377;
  assign new_n14512 = new_n12872 ^ new_n10584;
  assign new_n14513 = new_n10007 ^ new_n4633;
  assign new_n14514 = new_n14513 ^ new_n10814;
  assign new_n14515 = new_n14514 ^ new_n11024;
  assign new_n14516 = new_n14515 ^ new_n14512;
  assign new_n14517 = new_n11169 ^ new_n11159;
  assign new_n14518 = new_n14517 ^ new_n11205;
  assign new_n14519 = new_n9578 ^ new_n4776;
  assign new_n14520 = new_n14519 ^ new_n11190;
  assign new_n14521 = new_n14520 ^ new_n12875;
  assign new_n14522 = new_n14521 ^ new_n14518;
  assign new_n14523 = new_n11190 ^ new_n11062;
  assign new_n14524 = new_n14523 ^ new_n12883;
  assign new_n14525 = new_n9919 ^ new_n4703;
  assign new_n14526 = new_n14525 ^ new_n11079;
  assign new_n14527 = new_n14526 ^ new_n11148;
  assign new_n14528 = new_n14527 ^ new_n14524;
  assign new_n14529 = new_n14528 ^ new_n14522;
  assign new_n14530 = new_n9978 ^ new_n4752;
  assign new_n14531 = new_n14530 ^ new_n11205;
  assign new_n14532 = new_n12892 ^ new_n11131;
  assign new_n14533 = new_n14532 ^ new_n14531;
  assign new_n14534 = new_n14533 ^ new_n14529;
  assign new_n14535 = new_n14534 ^ new_n14516;
  assign new_n14536 = new_n10023 ^ new_n4663;
  assign new_n14537 = new_n14536 ^ new_n11071;
  assign new_n14538 = new_n12910 ^ new_n11190;
  assign new_n14539 = new_n14538 ^ new_n14537;
  assign new_n14540 = new_n12904 ^ new_n11024;
  assign new_n14541 = new_n10046 ^ new_n4615;
  assign new_n14542 = new_n14541 ^ new_n11113;
  assign new_n14543 = new_n14542 ^ new_n14540;
  assign new_n14544 = new_n14543 ^ new_n14516;
  assign new_n14545 = new_n14544 ^ new_n14539;
  assign new_n14546 = new_n10058 ^ new_n1402;
  assign new_n14547 = new_n14546 ^ new_n12899;
  assign new_n14548 = new_n14547 ^ new_n11190;
  assign new_n14549 = new_n11112 ^ new_n11101;
  assign new_n14550 = new_n14549 ^ new_n11159;
  assign new_n14551 = new_n14550 ^ new_n14548;
  assign new_n14552 = new_n14551 ^ new_n14545;
  assign new_n14553 = ~new_n14539 & ~new_n14552;
  assign new_n14554 = new_n14553 ^ new_n14551;
  assign new_n14555 = new_n12879 ^ new_n10432;
  assign new_n14556 = new_n10085 ^ new_n4731;
  assign new_n14557 = new_n14556 ^ new_n11189;
  assign new_n14558 = new_n14557 ^ new_n10814;
  assign new_n14559 = new_n14558 ^ new_n14555;
  assign new_n14560 = new_n14559 ^ new_n14551;
  assign new_n14561 = new_n14560 ^ new_n14529;
  assign new_n14562 = new_n14551 ^ new_n14528;
  assign new_n14563 = new_n14559 ^ new_n14533;
  assign new_n14564 = new_n14563 ^ new_n14562;
  assign new_n14565 = ~new_n14561 & new_n14564;
  assign new_n14566 = new_n14565 ^ new_n14516;
  assign new_n14567 = new_n14566 ^ new_n14554;
  assign new_n14568 = new_n14528 & new_n14545;
  assign new_n14569 = new_n14568 ^ new_n14528;
  assign new_n14570 = new_n14543 ^ new_n14534;
  assign new_n14571 = new_n14559 ^ new_n14528;
  assign new_n14572 = ~new_n14571 & new_n14570;
  assign new_n14573 = new_n14572 ^ new_n14569;
  assign new_n14574 = new_n14573 ^ new_n14563;
  assign new_n14575 = new_n14535 & new_n14560;
  assign new_n14576 = new_n14551 ^ new_n14543;
  assign new_n14577 = new_n14576 ^ new_n14563;
  assign new_n14578 = new_n14551 ^ new_n14533;
  assign new_n14579 = ~new_n14577 & ~new_n14578;
  assign new_n14580 = new_n14579 ^ new_n14575;
  assign new_n14581 = new_n14543 ^ new_n14522;
  assign new_n14582 = new_n14581 ^ new_n14580;
  assign new_n14583 = new_n14582 ^ new_n14574;
  assign new_n14584 = new_n14566 ^ new_n14561;
  assign new_n14585 = new_n14561 ^ new_n14539;
  assign new_n14586 = new_n14545 ^ new_n14528;
  assign new_n14587 = new_n14586 ^ new_n14563;
  assign new_n14588 = ~new_n14587 & new_n14585;
  assign new_n14589 = new_n14588 ^ new_n14533;
  assign new_n14590 = new_n14589 ^ new_n14580;
  assign new_n14591 = new_n14590 ^ new_n14584;
  assign new_n14592 = ~new_n14583 & new_n14591;
  assign new_n14593 = new_n14592 ^ new_n14567;
  assign new_n14594 = new_n14561 ^ new_n14544;
  assign new_n14595 = ~new_n14563 & ~new_n14594;
  assign new_n14596 = new_n14595 ^ new_n14575;
  assign new_n14597 = new_n14596 ^ new_n14570;
  assign new_n14598 = new_n14597 ^ new_n14593;
  assign new_n14599 = new_n14539 ^ new_n14535;
  assign new_n14600 = new_n14559 ^ new_n14545;
  assign new_n14601 = ~new_n14599 & ~new_n14600;
  assign new_n14602 = new_n14601 ^ new_n14568;
  assign new_n14603 = new_n14595 ^ new_n14579;
  assign new_n14604 = new_n14603 ^ new_n14602;
  assign new_n14605 = ~new_n14604 & new_n14598;
  assign new_n14606 = new_n14559 ^ new_n14543;
  assign new_n14607 = new_n14588 ^ new_n14553;
  assign new_n14608 = new_n14607 ^ new_n14603;
  assign new_n14609 = new_n14608 ^ new_n14606;
  assign new_n14610 = new_n14601 ^ new_n14572;
  assign new_n14611 = new_n14610 ^ new_n14559;
  assign new_n14612 = new_n14611 ^ new_n14597;
  assign new_n14613 = new_n14612 ^ new_n14592;
  assign new_n14614 = new_n14609 & new_n14613;
  assign new_n14615 = new_n14614 ^ new_n14605;
  assign new_n14616 = new_n14611 ^ new_n14567;
  assign new_n14617 = new_n14616 ^ new_n14615;
  assign new_n14618 = new_n14535 & new_n14617;
  assign new_n14619 = new_n14543 ^ new_n14528;
  assign new_n14620 = new_n14588 ^ new_n14569;
  assign new_n14621 = new_n14614 ^ new_n14567;
  assign new_n14622 = new_n14621 ^ new_n14597;
  assign new_n14623 = new_n14605 ^ new_n14592;
  assign new_n14624 = new_n14612 & new_n14623;
  assign new_n14625 = new_n14624 ^ new_n14613;
  assign new_n14626 = new_n14622 & new_n14625;
  assign new_n14627 = new_n14626 ^ new_n14624;
  assign new_n14628 = new_n14627 ^ new_n14620;
  assign new_n14629 = new_n14628 ^ new_n14619;
  assign new_n14630 = new_n14629 ^ new_n14551;
  assign new_n14631 = new_n14614 ^ new_n14572;
  assign new_n14632 = new_n14631 ^ new_n14566;
  assign new_n14633 = new_n14632 ^ new_n14630;
  assign new_n14634 = ~new_n14577 & ~new_n14633;
  assign new_n14635 = new_n14634 ^ new_n14618;
  assign new_n14636 = new_n14624 ^ new_n14605;
  assign new_n14637 = new_n14636 ^ new_n14604;
  assign new_n14638 = ~new_n14637 & new_n14585;
  assign new_n14639 = new_n14624 ^ new_n14583;
  assign new_n14640 = ~new_n14561 & ~new_n14639;
  assign new_n14641 = new_n14640 ^ new_n14638;
  assign new_n14642 = ~new_n14639 & new_n14564;
  assign new_n14643 = new_n14642 ^ new_n14641;
  assign new_n14644 = new_n14560 & new_n14617;
  assign new_n14645 = ~new_n14578 & ~new_n14633;
  assign new_n14646 = new_n14645 ^ new_n14644;
  assign new_n14647 = ~new_n14587 & ~new_n14637;
  assign new_n14648 = new_n14647 ^ new_n14646;
  assign new_n14649 = new_n14648 ^ new_n14643;
  assign new_n14650 = new_n14649 ^ new_n14635;
  assign new_n14651 = new_n14492 ^ new_n14406;
  assign new_n14652 = new_n14473 ^ new_n14431;
  assign new_n14653 = new_n14652 ^ new_n14425;
  assign new_n14654 = new_n14653 ^ new_n14651;
  assign new_n14655 = ~new_n14654 & new_n14436;
  assign new_n14656 = new_n14655 ^ new_n14477;
  assign new_n14657 = new_n14487 ^ new_n14464;
  assign new_n14658 = new_n14657 ^ new_n14463;
  assign new_n14659 = ~new_n14658 & new_n14446;
  assign new_n14660 = new_n14659 ^ new_n14502;
  assign new_n14661 = ~new_n14501 & new_n14423;
  assign new_n14662 = new_n14661 ^ new_n14660;
  assign new_n14663 = ~new_n14658 & new_n14445;
  assign new_n14664 = ~new_n14654 & new_n14437;
  assign new_n14665 = new_n14664 ^ new_n14478;
  assign new_n14666 = new_n14665 ^ new_n14663;
  assign new_n14667 = new_n14666 ^ new_n14662;
  assign new_n14668 = new_n14667 ^ new_n14656;
  assign new_n14669 = new_n14668 ^ new_n14650;
  assign new_n14670 = new_n14669 ^ new_n14511;
  assign new_n14671 = new_n14670 ^ new_n14235;
  assign new_n14672 = new_n14090 ^ new_n14055;
  assign new_n14673 = new_n13969 & new_n14069;
  assign new_n14674 = new_n14673 ^ new_n14078;
  assign new_n14675 = new_n14674 ^ new_n14672;
  assign new_n14676 = new_n14675 ^ new_n12897;
  assign new_n14677 = new_n14229 ^ new_n14202;
  assign new_n14678 = new_n14188 ^ new_n14123;
  assign new_n14679 = new_n14190 ^ new_n14184;
  assign new_n14680 = new_n14679 ^ new_n14213;
  assign new_n14681 = new_n14680 ^ new_n14678;
  assign new_n14682 = new_n14132 & new_n14681;
  assign new_n14683 = ~new_n14182 & ~new_n14206;
  assign new_n14684 = ~new_n14177 & new_n14681;
  assign new_n14685 = new_n14684 ^ new_n14683;
  assign new_n14686 = new_n14196 ^ new_n14188;
  assign new_n14687 = ~new_n14139 & new_n14686;
  assign new_n14688 = new_n14687 ^ new_n14224;
  assign new_n14689 = new_n14210 ^ new_n14198;
  assign new_n14690 = new_n14689 ^ new_n14174;
  assign new_n14691 = ~new_n14153 & new_n14690;
  assign new_n14692 = new_n14691 ^ new_n14688;
  assign new_n14693 = new_n14692 ^ new_n14685;
  assign new_n14694 = new_n14693 ^ new_n14682;
  assign new_n14695 = new_n14694 ^ new_n14677;
  assign new_n14696 = new_n14695 ^ new_n14676;
  assign new_n14697 = new_n14355 ^ new_n14331;
  assign new_n14698 = ~new_n14272 & ~new_n14697;
  assign new_n14699 = new_n14356 ^ new_n14339;
  assign new_n14700 = new_n14699 ^ new_n14338;
  assign new_n14701 = new_n14307 & new_n14700;
  assign new_n14702 = new_n14359 ^ new_n14289;
  assign new_n14703 = new_n14332 ^ new_n14281;
  assign new_n14704 = new_n14703 ^ new_n14303;
  assign new_n14705 = new_n14704 ^ new_n14702;
  assign new_n14706 = new_n14290 & new_n14705;
  assign new_n14707 = new_n14706 ^ new_n14344;
  assign new_n14708 = new_n14707 ^ new_n14701;
  assign new_n14709 = new_n14708 ^ new_n14698;
  assign new_n14710 = new_n14280 & new_n14372;
  assign new_n14711 = new_n14710 ^ new_n14709;
  assign new_n14712 = ~new_n14301 & new_n14368;
  assign new_n14713 = new_n14305 & new_n14700;
  assign new_n14714 = new_n14713 ^ new_n14369;
  assign new_n14715 = new_n14714 ^ new_n14712;
  assign new_n14716 = new_n14715 ^ new_n14711;
  assign new_n14717 = new_n14489 ^ new_n14468;
  assign new_n14718 = new_n14411 & new_n14717;
  assign new_n14719 = new_n14718 ^ new_n14666;
  assign new_n14720 = new_n14429 & new_n14497;
  assign new_n14721 = new_n14720 ^ new_n14719;
  assign new_n14722 = new_n14721 ^ new_n14662;
  assign new_n14723 = new_n14722 ^ new_n14716;
  assign new_n14724 = new_n14644 ^ new_n14618;
  assign new_n14725 = new_n14605 ^ new_n14559;
  assign new_n14726 = new_n14601 ^ new_n14553;
  assign new_n14727 = new_n14726 ^ new_n14629;
  assign new_n14728 = new_n14727 ^ new_n14725;
  assign new_n14729 = ~new_n14563 & ~new_n14728;
  assign new_n14730 = ~new_n14600 & new_n14622;
  assign new_n14731 = ~new_n14594 & ~new_n14728;
  assign new_n14732 = new_n14731 ^ new_n14730;
  assign new_n14733 = new_n14612 ^ new_n14605;
  assign new_n14734 = ~new_n14539 & new_n14733;
  assign new_n14735 = new_n14734 ^ new_n14640;
  assign new_n14736 = new_n14626 ^ new_n14614;
  assign new_n14737 = new_n14736 ^ new_n14591;
  assign new_n14738 = ~new_n14571 & new_n14737;
  assign new_n14739 = new_n14738 ^ new_n14735;
  assign new_n14740 = new_n14739 ^ new_n14732;
  assign new_n14741 = new_n14740 ^ new_n14729;
  assign new_n14742 = new_n14741 ^ new_n14724;
  assign new_n14743 = new_n14742 ^ new_n14510;
  assign new_n14744 = new_n14743 ^ new_n14723;
  assign new_n14745 = new_n14744 ^ new_n14696;
  assign new_n14746 = new_n14745 ^ new_n14671;
  assign new_n14747 = new_n14505 ^ new_n14498;
  assign new_n14748 = new_n14718 ^ new_n14655;
  assign new_n14749 = new_n14444 & new_n14717;
  assign new_n14750 = new_n14458 & new_n14485;
  assign new_n14751 = new_n14750 ^ new_n14749;
  assign new_n14752 = new_n14751 ^ new_n14665;
  assign new_n14753 = new_n14752 ^ new_n14748;
  assign new_n14754 = new_n14753 ^ new_n14747;
  assign new_n14755 = new_n14691 ^ new_n14684;
  assign new_n14756 = new_n14210 ^ new_n14193;
  assign new_n14757 = ~new_n14149 & ~new_n14756;
  assign new_n14758 = new_n14757 ^ new_n14218;
  assign new_n14759 = ~new_n14756 & new_n14168;
  assign new_n14760 = ~new_n14183 & ~new_n14206;
  assign new_n14761 = new_n14760 ^ new_n14759;
  assign new_n14762 = new_n14761 ^ new_n14231;
  assign new_n14763 = new_n14762 ^ new_n14758;
  assign new_n14764 = new_n14763 ^ new_n14755;
  assign new_n14765 = new_n14764 ^ new_n14754;
  assign new_n14766 = new_n14712 ^ new_n14343;
  assign new_n14767 = ~new_n14292 & new_n14705;
  assign new_n14768 = new_n14767 ^ new_n14711;
  assign new_n14769 = new_n14768 ^ new_n14766;
  assign new_n14770 = new_n14661 ^ new_n14477;
  assign new_n14771 = new_n14721 ^ new_n14655;
  assign new_n14772 = new_n14771 ^ new_n14770;
  assign new_n14773 = new_n14772 ^ new_n14769;
  assign new_n14774 = new_n14773 ^ new_n14765;
  assign new_n14775 = new_n14710 ^ new_n14374;
  assign new_n14776 = ~new_n14697 & new_n14306;
  assign new_n14777 = ~new_n14319 & ~new_n14354;
  assign new_n14778 = new_n14777 ^ new_n14776;
  assign new_n14779 = new_n14778 ^ new_n14707;
  assign new_n14780 = new_n14779 ^ new_n14775;
  assign new_n14781 = new_n14720 ^ new_n14504;
  assign new_n14782 = new_n14781 ^ new_n14752;
  assign new_n14783 = new_n14782 ^ new_n14780;
  assign new_n14784 = new_n14076 ^ new_n14070;
  assign new_n14785 = new_n14047 ^ new_n14045;
  assign new_n14786 = ~new_n14046 & new_n13998;
  assign new_n14787 = ~new_n14011 & ~new_n14032;
  assign new_n14788 = new_n14787 ^ new_n14786;
  assign new_n14789 = new_n14788 ^ new_n14056;
  assign new_n14790 = new_n14789 ^ new_n14785;
  assign new_n14791 = new_n14790 ^ new_n14784;
  assign new_n14792 = new_n14791 ^ new_n12885;
  assign new_n14793 = new_n14738 ^ new_n14731;
  assign new_n14794 = new_n14626 ^ new_n14609;
  assign new_n14795 = ~new_n14545 & new_n14794;
  assign new_n14796 = new_n14795 ^ new_n14634;
  assign new_n14797 = new_n14586 & new_n14794;
  assign new_n14798 = ~new_n14599 & new_n14622;
  assign new_n14799 = new_n14798 ^ new_n14797;
  assign new_n14800 = new_n14799 ^ new_n14646;
  assign new_n14801 = new_n14800 ^ new_n14796;
  assign new_n14802 = new_n14801 ^ new_n14793;
  assign new_n14803 = new_n14802 ^ new_n14792;
  assign new_n14804 = new_n14803 ^ new_n14783;
  assign new_n14805 = new_n14804 ^ new_n14774;
  assign new_n14806 = new_n14787 ^ new_n14094;
  assign new_n14807 = new_n14092 ^ new_n14072;
  assign new_n14808 = new_n14807 ^ new_n14058;
  assign new_n14809 = new_n14808 ^ new_n14806;
  assign new_n14810 = new_n14809 ^ new_n12889;
  assign new_n14811 = new_n14760 ^ new_n14226;
  assign new_n14812 = new_n14687 ^ new_n14222;
  assign new_n14813 = new_n14757 ^ new_n14232;
  assign new_n14814 = new_n14813 ^ new_n14812;
  assign new_n14815 = new_n14814 ^ new_n14811;
  assign new_n14816 = new_n14815 ^ new_n14810;
  assign new_n14817 = new_n14816 ^ new_n14773;
  assign new_n14818 = ~new_n14326 & new_n14366;
  assign new_n14819 = new_n14818 ^ new_n14768;
  assign new_n14820 = new_n14819 ^ new_n14375;
  assign new_n14821 = new_n14412 & new_n14499;
  assign new_n14822 = new_n14821 ^ new_n14771;
  assign new_n14823 = new_n14822 ^ new_n14508;
  assign new_n14824 = new_n14823 ^ new_n14820;
  assign new_n14825 = new_n14798 ^ new_n14642;
  assign new_n14826 = new_n14734 ^ new_n14638;
  assign new_n14827 = new_n14795 ^ new_n14648;
  assign new_n14828 = new_n14827 ^ new_n14826;
  assign new_n14829 = new_n14828 ^ new_n14825;
  assign new_n14830 = new_n14750 ^ new_n14661;
  assign new_n14831 = new_n14659 ^ new_n14500;
  assign new_n14832 = new_n14831 ^ new_n14719;
  assign new_n14833 = new_n14832 ^ new_n14830;
  assign new_n14834 = new_n14833 ^ new_n14829;
  assign new_n14835 = new_n14834 ^ new_n14824;
  assign new_n14836 = new_n14835 ^ new_n14817;
  assign new_n14837 = new_n14836 ^ new_n14805;
  assign new_n14838 = new_n14777 ^ new_n14712;
  assign new_n14839 = new_n14713 ^ new_n14367;
  assign new_n14840 = new_n14839 ^ new_n14709;
  assign new_n14841 = new_n14840 ^ new_n14838;
  assign new_n14842 = new_n14841 ^ new_n14833;
  assign new_n14843 = new_n14570 & new_n14737;
  assign new_n14844 = new_n14843 ^ new_n14827;
  assign new_n14845 = new_n14844 ^ new_n14643;
  assign new_n14846 = new_n14845 ^ new_n14722;
  assign new_n14847 = new_n14846 ^ new_n14842;
  assign new_n14848 = new_n14095 ^ new_n14062;
  assign new_n14849 = new_n14848 ^ new_n12877;
  assign new_n14850 = new_n14152 & new_n14690;
  assign new_n14851 = new_n14850 ^ new_n14813;
  assign new_n14852 = new_n14851 ^ new_n14227;
  assign new_n14853 = new_n14852 ^ new_n14849;
  assign new_n14854 = new_n14853 ^ new_n14773;
  assign new_n14855 = new_n14854 ^ new_n14847;
  assign new_n14856 = new_n14094 ^ new_n14090;
  assign new_n14857 = new_n14856 ^ new_n14063;
  assign new_n14858 = new_n14857 ^ new_n12870;
  assign new_n14859 = new_n14226 ^ new_n14202;
  assign new_n14860 = new_n14851 ^ new_n14218;
  assign new_n14861 = new_n14860 ^ new_n14859;
  assign new_n14862 = new_n14861 ^ new_n14858;
  assign new_n14863 = new_n14767 ^ new_n14343;
  assign new_n14864 = new_n14715 ^ new_n14708;
  assign new_n14865 = new_n14864 ^ new_n14863;
  assign new_n14866 = new_n14865 ^ new_n14668;
  assign new_n14867 = new_n14642 ^ new_n14618;
  assign new_n14868 = new_n14844 ^ new_n14634;
  assign new_n14869 = new_n14868 ^ new_n14867;
  assign new_n14870 = new_n14869 ^ new_n14772;
  assign new_n14871 = new_n14870 ^ new_n14866;
  assign new_n14872 = new_n14871 ^ new_n14862;
  assign new_n14873 = new_n14872 ^ new_n14855;
  assign new_n14874 = new_n14873 ^ new_n14837;
  assign new_n14875 = new_n14874 ^ new_n14746;
  assign new_n14876 = new_n14077 ^ new_n14061;
  assign new_n14877 = new_n14876 ^ new_n14789;
  assign new_n14878 = new_n14877 ^ new_n12908;
  assign new_n14879 = new_n14843 ^ new_n14739;
  assign new_n14880 = new_n14879 ^ new_n14800;
  assign new_n14881 = new_n14880 ^ new_n14878;
  assign new_n14882 = new_n14850 ^ new_n14692;
  assign new_n14883 = new_n14882 ^ new_n14762;
  assign new_n14884 = new_n14883 ^ new_n14782;
  assign new_n14885 = new_n14884 ^ new_n14773;
  assign new_n14886 = new_n14885 ^ new_n14881;
  assign new_n14887 = new_n14886 ^ new_n14746;
  assign new_n14888 = new_n14887 ^ new_n14855;
  assign new_n14889 = ~new_n14886 & ~new_n14888;
  assign new_n14890 = new_n14889 ^ new_n14855;
  assign new_n14891 = new_n14855 ^ new_n14805;
  assign new_n14892 = new_n14373 ^ new_n14364;
  assign new_n14893 = new_n14767 ^ new_n14698;
  assign new_n14894 = new_n14893 ^ new_n14779;
  assign new_n14895 = new_n14894 ^ new_n14892;
  assign new_n14896 = ~new_n14552 & new_n14733;
  assign new_n14897 = new_n14896 ^ new_n14868;
  assign new_n14898 = new_n14897 ^ new_n14740;
  assign new_n14899 = new_n14898 ^ new_n14823;
  assign new_n14900 = new_n14899 ^ new_n14895;
  assign new_n14901 = new_n14079 ^ new_n12916;
  assign new_n14902 = new_n14149 ^ new_n14128;
  assign new_n14903 = ~new_n14902 & new_n14686;
  assign new_n14904 = new_n14903 ^ new_n14860;
  assign new_n14905 = new_n14904 ^ new_n14693;
  assign new_n14906 = new_n14905 ^ new_n14901;
  assign new_n14907 = new_n14906 ^ new_n14754;
  assign new_n14908 = new_n14907 ^ new_n14900;
  assign new_n14909 = new_n14908 ^ new_n14872;
  assign new_n14910 = new_n14909 ^ new_n14891;
  assign new_n14911 = ~new_n14874 & ~new_n14910;
  assign new_n14912 = new_n14911 ^ new_n14671;
  assign new_n14913 = new_n14912 ^ new_n14890;
  assign new_n14914 = new_n14805 & new_n14887;
  assign new_n14915 = new_n14914 ^ new_n14805;
  assign new_n14916 = new_n14908 ^ new_n14837;
  assign new_n14917 = new_n14916 ^ new_n14745;
  assign new_n14918 = new_n14872 ^ new_n14805;
  assign new_n14919 = ~new_n14918 & new_n14917;
  assign new_n14920 = new_n14919 ^ new_n14915;
  assign new_n14921 = new_n14920 ^ new_n14909;
  assign new_n14922 = new_n14855 ^ new_n14745;
  assign new_n14923 = new_n14922 ^ new_n14909;
  assign new_n14924 = new_n14908 ^ new_n14855;
  assign new_n14925 = ~new_n14923 & new_n14924;
  assign new_n14926 = new_n14916 ^ new_n14671;
  assign new_n14927 = new_n14873 & new_n14926;
  assign new_n14928 = new_n14927 ^ new_n14925;
  assign new_n14929 = new_n14836 ^ new_n14745;
  assign new_n14930 = new_n14929 ^ new_n14928;
  assign new_n14931 = new_n14930 ^ new_n14921;
  assign new_n14932 = new_n14912 ^ new_n14874;
  assign new_n14933 = new_n14886 ^ new_n14874;
  assign new_n14934 = new_n14887 ^ new_n14805;
  assign new_n14935 = new_n14934 ^ new_n14909;
  assign new_n14936 = new_n14933 & new_n14935;
  assign new_n14937 = new_n14936 ^ new_n14927;
  assign new_n14938 = new_n14925 ^ new_n14908;
  assign new_n14939 = new_n14938 ^ new_n14937;
  assign new_n14940 = new_n14939 ^ new_n14932;
  assign new_n14941 = ~new_n14931 & new_n14940;
  assign new_n14942 = new_n14941 ^ new_n14913;
  assign new_n14943 = ~new_n14875 & new_n14909;
  assign new_n14944 = new_n14943 ^ new_n14927;
  assign new_n14945 = new_n14944 ^ new_n14917;
  assign new_n14946 = new_n14945 ^ new_n14942;
  assign new_n14947 = new_n14887 ^ new_n14872;
  assign new_n14948 = new_n14926 ^ new_n14886;
  assign new_n14949 = ~new_n14947 & ~new_n14948;
  assign new_n14950 = new_n14949 ^ new_n14914;
  assign new_n14951 = new_n14943 ^ new_n14925;
  assign new_n14952 = new_n14951 ^ new_n14950;
  assign new_n14953 = ~new_n14946 & ~new_n14952;
  assign new_n14954 = new_n14953 ^ new_n14872;
  assign new_n14955 = new_n14949 ^ new_n14889;
  assign new_n14956 = new_n14805 ^ new_n14745;
  assign new_n14957 = new_n14936 ^ new_n14915;
  assign new_n14958 = new_n14949 ^ new_n14919;
  assign new_n14959 = new_n14958 ^ new_n14872;
  assign new_n14960 = new_n14959 ^ new_n14945;
  assign new_n14961 = new_n14953 ^ new_n14941;
  assign new_n14962 = ~new_n14960 & ~new_n14961;
  assign new_n14963 = new_n14962 ^ new_n14953;
  assign new_n14964 = new_n14960 ^ new_n14941;
  assign new_n14965 = new_n14872 ^ new_n14745;
  assign new_n14966 = new_n14936 ^ new_n14889;
  assign new_n14967 = new_n14966 ^ new_n14951;
  assign new_n14968 = new_n14967 ^ new_n14965;
  assign new_n14969 = ~new_n14968 & new_n14964;
  assign new_n14970 = new_n14969 ^ new_n14913;
  assign new_n14971 = new_n14970 ^ new_n14945;
  assign new_n14972 = ~new_n14963 & ~new_n14971;
  assign new_n14973 = new_n14964 ^ new_n14963;
  assign new_n14974 = new_n14973 ^ new_n14972;
  assign new_n14975 = new_n14974 ^ new_n14957;
  assign new_n14976 = new_n14975 ^ new_n14956;
  assign new_n14977 = new_n14976 ^ new_n14955;
  assign new_n14978 = new_n14977 ^ new_n14954;
  assign new_n14979 = ~new_n14875 & ~new_n14978;
  assign new_n14980 = new_n14972 ^ new_n14969;
  assign new_n14981 = new_n14980 ^ new_n14940;
  assign new_n14982 = ~new_n14918 & new_n14981;
  assign new_n14983 = new_n14982 ^ new_n14979;
  assign new_n14984 = new_n14972 ^ new_n14968;
  assign new_n14985 = ~new_n14887 & ~new_n14984;
  assign new_n14986 = new_n14976 ^ new_n14855;
  assign new_n14987 = new_n14969 ^ new_n14919;
  assign new_n14988 = new_n14987 ^ new_n14912;
  assign new_n14989 = new_n14988 ^ new_n14986;
  assign new_n14990 = ~new_n14923 & new_n14989;
  assign new_n14991 = new_n14990 ^ new_n14985;
  assign new_n14992 = ~new_n14948 & ~new_n14971;
  assign new_n14993 = ~new_n14984 & new_n14934;
  assign new_n14994 = new_n14993 ^ new_n14992;
  assign new_n14995 = new_n14924 & new_n14989;
  assign new_n14996 = new_n14969 ^ new_n14953;
  assign new_n14997 = new_n14959 ^ new_n14913;
  assign new_n14998 = new_n14997 ^ new_n14996;
  assign new_n14999 = ~new_n14998 & new_n14873;
  assign new_n15000 = new_n14999 ^ new_n14995;
  assign new_n15001 = new_n15000 ^ new_n14994;
  assign new_n15002 = new_n15001 ^ new_n14991;
  assign new_n15003 = new_n15002 ^ new_n14983;
  assign new_n15004 = new_n15003 ^ new_n14089;
  assign new_n15005 = new_n15004 ^ new_n14081;
  assign new_n15006 = new_n15005 ^ new_n13829;
  assign new_n15007 = ~new_n11588 & ~new_n11686;
  assign new_n15008 = new_n15007 ^ new_n14084;
  assign new_n15009 = ~new_n11652 & new_n11610;
  assign new_n15010 = new_n15009 ^ new_n11685;
  assign new_n15011 = new_n15010 ^ new_n11670;
  assign new_n15012 = new_n15011 ^ new_n15008;
  assign new_n15013 = new_n12688 & new_n12709;
  assign new_n15014 = ~new_n12750 & new_n12666;
  assign new_n15015 = new_n15014 ^ new_n15013;
  assign new_n15016 = ~new_n12726 & new_n12670;
  assign new_n15017 = new_n15016 ^ new_n12749;
  assign new_n15018 = new_n15017 ^ new_n12735;
  assign new_n15019 = new_n15018 ^ new_n15015;
  assign new_n15020 = new_n15019 ^ new_n15012;
  assign new_n15021 = ~new_n13760 & ~new_n13781;
  assign new_n15022 = ~new_n13823 & new_n13739;
  assign new_n15023 = new_n15022 ^ new_n15021;
  assign new_n15024 = ~new_n13743 & ~new_n13807;
  assign new_n15025 = new_n15024 ^ new_n13822;
  assign new_n15026 = new_n15025 ^ new_n13810;
  assign new_n15027 = new_n15026 ^ new_n15023;
  assign new_n15028 = new_n15027 ^ new_n15020;
  assign new_n15029 = ~new_n13847 & ~new_n13950;
  assign new_n15030 = ~new_n13885 & ~new_n13906;
  assign new_n15031 = new_n15030 ^ new_n15029;
  assign new_n15032 = ~new_n13915 & new_n13873;
  assign new_n15033 = new_n15032 ^ new_n13949;
  assign new_n15034 = new_n15033 ^ new_n13933;
  assign new_n15035 = new_n15034 ^ new_n15031;
  assign new_n15036 = new_n15035 ^ new_n14809;
  assign new_n15037 = new_n15036 ^ new_n884;
  assign new_n15038 = new_n14973 ^ new_n14931;
  assign new_n15039 = ~new_n14910 & new_n15038;
  assign new_n15040 = ~new_n14998 & new_n14926;
  assign new_n15041 = new_n15040 ^ new_n15039;
  assign new_n15042 = new_n14973 ^ new_n14953;
  assign new_n15043 = new_n15042 ^ new_n14952;
  assign new_n15044 = new_n14935 & new_n15043;
  assign new_n15045 = new_n15044 ^ new_n15000;
  assign new_n15046 = new_n15045 ^ new_n14985;
  assign new_n15047 = new_n14917 & new_n14981;
  assign new_n15048 = new_n15047 ^ new_n15046;
  assign new_n15049 = new_n15048 ^ new_n14990;
  assign new_n15050 = new_n15049 ^ new_n15041;
  assign new_n15051 = ~new_n11666 & new_n11600;
  assign new_n15052 = new_n15051 ^ new_n15007;
  assign new_n15053 = new_n15052 ^ new_n11676;
  assign new_n15054 = new_n15053 ^ new_n15050;
  assign new_n15055 = new_n15054 ^ new_n15037;
  assign new_n15056 = new_n14960 ^ new_n14953;
  assign new_n15057 = ~new_n14888 & new_n15056;
  assign new_n15058 = new_n15057 ^ new_n15049;
  assign new_n15059 = ~new_n14947 & ~new_n14971;
  assign new_n15060 = new_n15059 ^ new_n14979;
  assign new_n15061 = ~new_n14886 & new_n15056;
  assign new_n15062 = ~new_n14874 & new_n15038;
  assign new_n15063 = new_n15062 ^ new_n15061;
  assign new_n15064 = new_n15063 ^ new_n14982;
  assign new_n15065 = new_n15064 ^ new_n15060;
  assign new_n15066 = new_n15065 ^ new_n15058;
  assign new_n15067 = new_n15066 ^ new_n11692;
  assign new_n15068 = new_n15067 ^ new_n15055;
  assign new_n15069 = new_n15068 ^ new_n15028;
  assign new_n15070 = new_n12753 ^ new_n12747;
  assign new_n15071 = new_n12724 ^ new_n12722;
  assign new_n15072 = new_n12671 & new_n12723;
  assign new_n15073 = new_n15072 ^ new_n15013;
  assign new_n15074 = new_n15073 ^ new_n12733;
  assign new_n15075 = new_n15074 ^ new_n15071;
  assign new_n15076 = new_n15075 ^ new_n15070;
  assign new_n15077 = new_n15076 ^ new_n15054;
  assign new_n15078 = new_n11690 ^ new_n11673;
  assign new_n15079 = new_n15078 ^ new_n14087;
  assign new_n15080 = new_n15064 ^ new_n15047;
  assign new_n15081 = new_n15080 ^ new_n15001;
  assign new_n15082 = new_n15081 ^ new_n15079;
  assign new_n15083 = new_n15082 ^ new_n15077;
  assign new_n15084 = new_n13948 ^ new_n13945;
  assign new_n15085 = new_n13938 ^ new_n13912;
  assign new_n15086 = ~new_n13911 & new_n13871;
  assign new_n15087 = new_n15086 ^ new_n15030;
  assign new_n15088 = new_n15087 ^ new_n13931;
  assign new_n15089 = new_n15088 ^ new_n15085;
  assign new_n15090 = new_n15089 ^ new_n15084;
  assign new_n15091 = new_n15090 ^ new_n14791;
  assign new_n15092 = new_n15091 ^ new_n892;
  assign new_n15093 = new_n13821 ^ new_n13818;
  assign new_n15094 = new_n13799 ^ new_n13794;
  assign new_n15095 = ~new_n13798 & new_n13744;
  assign new_n15096 = new_n15095 ^ new_n15021;
  assign new_n15097 = new_n15096 ^ new_n13805;
  assign new_n15098 = new_n15097 ^ new_n15094;
  assign new_n15099 = new_n15098 ^ new_n15093;
  assign new_n15100 = new_n15099 ^ new_n15092;
  assign new_n15101 = new_n15100 ^ new_n14089;
  assign new_n15102 = new_n15101 ^ new_n15083;
  assign new_n15103 = new_n15102 ^ new_n15069;
  assign new_n15104 = new_n15103 ^ new_n15006;
  assign new_n15105 = new_n12653 & new_n12731;
  assign new_n15106 = new_n15105 ^ new_n12722;
  assign new_n15107 = new_n15016 ^ new_n12751;
  assign new_n15108 = new_n15107 ^ new_n15014;
  assign new_n15109 = new_n15108 ^ new_n12734;
  assign new_n15110 = new_n15109 ^ new_n15106;
  assign new_n15111 = new_n15051 ^ new_n11667;
  assign new_n15112 = new_n11598 & new_n11682;
  assign new_n15113 = new_n15112 ^ new_n11691;
  assign new_n15114 = new_n15113 ^ new_n15111;
  assign new_n15115 = new_n15040 ^ new_n14999;
  assign new_n15116 = ~new_n14978 & new_n14909;
  assign new_n15117 = new_n15116 ^ new_n15065;
  assign new_n15118 = new_n15117 ^ new_n15115;
  assign new_n15119 = new_n15118 ^ new_n15114;
  assign new_n15120 = new_n15119 ^ new_n15110;
  assign new_n15121 = ~new_n13929 & new_n13864;
  assign new_n15122 = new_n15121 ^ new_n13938;
  assign new_n15123 = new_n15032 ^ new_n13951;
  assign new_n15124 = new_n15123 ^ new_n15029;
  assign new_n15125 = new_n15124 ^ new_n13932;
  assign new_n15126 = new_n15125 ^ new_n15122;
  assign new_n15127 = new_n15126 ^ new_n14097;
  assign new_n15128 = new_n15127 ^ new_n820;
  assign new_n15129 = ~new_n13803 & new_n13726;
  assign new_n15130 = new_n15129 ^ new_n13794;
  assign new_n15131 = new_n15024 ^ new_n13824;
  assign new_n15132 = new_n15131 ^ new_n15022;
  assign new_n15133 = new_n15132 ^ new_n13809;
  assign new_n15134 = new_n15133 ^ new_n15130;
  assign new_n15135 = new_n15134 ^ new_n15128;
  assign new_n15136 = new_n15051 ^ new_n11675;
  assign new_n15137 = new_n15009 ^ new_n11687;
  assign new_n15138 = new_n15137 ^ new_n15007;
  assign new_n15139 = new_n15138 ^ new_n11669;
  assign new_n15140 = new_n15139 ^ new_n15136;
  assign new_n15141 = new_n15140 ^ new_n15135;
  assign new_n15142 = new_n15141 ^ new_n15120;
  assign new_n15143 = new_n15142 ^ new_n15104;
  assign new_n15144 = new_n15121 ^ new_n15029;
  assign new_n15145 = new_n15144 ^ new_n13939;
  assign new_n15146 = new_n15145 ^ new_n14857;
  assign new_n15147 = new_n15146 ^ new_n875;
  assign new_n15148 = new_n15040 ^ new_n14990;
  assign new_n15149 = new_n14933 & new_n15043;
  assign new_n15150 = new_n15149 ^ new_n15062;
  assign new_n15151 = new_n15150 ^ new_n15039;
  assign new_n15152 = new_n15151 ^ new_n15045;
  assign new_n15153 = new_n15152 ^ new_n15148;
  assign new_n15154 = new_n15153 ^ new_n15140;
  assign new_n15155 = new_n15154 ^ new_n15147;
  assign new_n15156 = new_n15129 ^ new_n15022;
  assign new_n15157 = new_n15156 ^ new_n13812;
  assign new_n15158 = new_n15105 ^ new_n15014;
  assign new_n15159 = new_n15158 ^ new_n12740;
  assign new_n15160 = new_n15159 ^ new_n15157;
  assign new_n15161 = new_n15160 ^ new_n15053;
  assign new_n15162 = new_n15161 ^ new_n15155;
  assign new_n15163 = new_n15138 ^ new_n11674;
  assign new_n15164 = new_n15151 ^ new_n15048;
  assign new_n15165 = new_n15164 ^ new_n15163;
  assign new_n15166 = new_n15105 ^ new_n12732;
  assign new_n15167 = ~new_n12746 & new_n12651;
  assign new_n15168 = new_n15167 ^ new_n12755;
  assign new_n15169 = new_n15168 ^ new_n15166;
  assign new_n15170 = new_n15169 ^ new_n15165;
  assign new_n15171 = new_n15121 ^ new_n13930;
  assign new_n15172 = new_n13846 & new_n13944;
  assign new_n15173 = new_n15172 ^ new_n13954;
  assign new_n15174 = new_n15173 ^ new_n15171;
  assign new_n15175 = new_n15174 ^ new_n14675;
  assign new_n15176 = new_n15175 ^ new_n843;
  assign new_n15177 = new_n15129 ^ new_n13804;
  assign new_n15178 = ~new_n13724 & new_n13817;
  assign new_n15179 = new_n15178 ^ new_n13827;
  assign new_n15180 = new_n15179 ^ new_n15177;
  assign new_n15181 = new_n15180 ^ new_n15176;
  assign new_n15182 = new_n15181 ^ new_n15114;
  assign new_n15183 = new_n15182 ^ new_n15170;
  assign new_n15184 = new_n15183 ^ new_n15162;
  assign new_n15185 = new_n15124 ^ new_n13937;
  assign new_n15186 = new_n15185 ^ new_n14848;
  assign new_n15187 = new_n15186 ^ new_n865;
  assign new_n15188 = new_n15187 ^ new_n15054;
  assign new_n15189 = new_n15039 ^ new_n14992;
  assign new_n15190 = new_n15149 ^ new_n15061;
  assign new_n15191 = new_n15190 ^ new_n15046;
  assign new_n15192 = new_n15191 ^ new_n15189;
  assign new_n15193 = new_n15192 ^ new_n15012;
  assign new_n15194 = new_n15193 ^ new_n15188;
  assign new_n15195 = new_n15132 ^ new_n13811;
  assign new_n15196 = new_n15195 ^ new_n15163;
  assign new_n15197 = new_n15108 ^ new_n12739;
  assign new_n15198 = new_n15197 ^ new_n15196;
  assign new_n15199 = new_n15198 ^ new_n15194;
  assign new_n15200 = new_n15199 ^ new_n15162;
  assign new_n15201 = new_n15200 ^ new_n15103;
  assign new_n15202 = new_n12754 ^ new_n12738;
  assign new_n15203 = new_n15202 ^ new_n15074;
  assign new_n15204 = new_n15203 ^ new_n15054;
  assign new_n15205 = new_n13953 ^ new_n13936;
  assign new_n15206 = new_n15205 ^ new_n15088;
  assign new_n15207 = new_n15206 ^ new_n14877;
  assign new_n15208 = new_n15207 ^ new_n856;
  assign new_n15209 = new_n13826 ^ new_n13797;
  assign new_n15210 = new_n15209 ^ new_n15097;
  assign new_n15211 = new_n15210 ^ new_n15208;
  assign new_n15212 = new_n15211 ^ new_n15079;
  assign new_n15213 = new_n15212 ^ new_n15204;
  assign new_n15214 = new_n15213 ^ new_n15201;
  assign new_n15215 = new_n15183 ^ new_n15142;
  assign new_n15216 = new_n15215 ^ new_n15213;
  assign new_n15217 = new_n15216 ^ new_n15102;
  assign new_n15218 = new_n15162 ^ new_n15006;
  assign new_n15219 = new_n15218 ^ new_n15217;
  assign new_n15220 = new_n15214 & new_n15219;
  assign new_n15221 = new_n15216 ^ new_n15199;
  assign new_n15222 = new_n15213 & new_n15221;
  assign new_n15223 = new_n15222 ^ new_n15220;
  assign new_n15224 = new_n15215 ^ new_n15201;
  assign new_n15225 = new_n15218 & new_n15224;
  assign new_n15226 = new_n15199 ^ new_n15006;
  assign new_n15227 = new_n15199 ^ new_n15183;
  assign new_n15228 = new_n15227 ^ new_n15218;
  assign new_n15229 = new_n15226 & new_n15228;
  assign new_n15230 = new_n15229 ^ new_n15225;
  assign new_n15231 = new_n15230 ^ new_n15223;
  assign new_n15232 = new_n15231 ^ new_n15184;
  assign new_n15233 = new_n15216 ^ new_n15162;
  assign new_n15234 = new_n15213 ^ new_n15143;
  assign new_n15235 = new_n15233 & new_n15234;
  assign new_n15236 = new_n15162 ^ new_n15102;
  assign new_n15237 = new_n15183 ^ new_n15104;
  assign new_n15238 = new_n15236 & new_n15237;
  assign new_n15239 = new_n15238 ^ new_n15235;
  assign new_n15240 = new_n15239 ^ new_n15162;
  assign new_n15241 = new_n15143 & new_n15200;
  assign new_n15242 = new_n15241 ^ new_n15225;
  assign new_n15243 = new_n15242 ^ new_n15237;
  assign new_n15244 = new_n15243 ^ new_n15240;
  assign new_n15245 = ~new_n15102 & ~new_n15216;
  assign new_n15246 = new_n15245 ^ new_n15102;
  assign new_n15247 = new_n15246 ^ new_n15238;
  assign new_n15248 = new_n15247 ^ new_n15218;
  assign new_n15249 = new_n15241 ^ new_n15229;
  assign new_n15250 = new_n15183 ^ new_n15069;
  assign new_n15251 = new_n15250 ^ new_n15249;
  assign new_n15252 = new_n15251 ^ new_n15248;
  assign new_n15253 = new_n15236 ^ new_n15226;
  assign new_n15254 = new_n15201 & new_n15253;
  assign new_n15255 = new_n15254 ^ new_n15142;
  assign new_n15256 = new_n15255 ^ new_n15201;
  assign new_n15257 = new_n15249 ^ new_n15220;
  assign new_n15258 = new_n15257 ^ new_n15006;
  assign new_n15259 = new_n15258 ^ new_n15256;
  assign new_n15260 = ~new_n15252 & new_n15259;
  assign new_n15261 = new_n15260 ^ new_n15244;
  assign new_n15262 = new_n15232 & new_n15261;
  assign new_n15263 = new_n15222 ^ new_n15199;
  assign new_n15264 = new_n15263 ^ new_n15255;
  assign new_n15265 = new_n15264 ^ new_n15260;
  assign new_n15266 = new_n15265 ^ new_n15243;
  assign new_n15267 = new_n15245 ^ new_n15235;
  assign new_n15268 = new_n15267 ^ new_n15230;
  assign new_n15269 = ~new_n15268 & new_n15266;
  assign new_n15270 = new_n15269 ^ new_n15262;
  assign new_n15271 = new_n15264 ^ new_n15240;
  assign new_n15272 = new_n15271 ^ new_n15270;
  assign new_n15273 = new_n15143 & new_n15272;
  assign new_n15274 = new_n15269 ^ new_n15260;
  assign new_n15275 = ~new_n15274 & new_n15244;
  assign new_n15276 = new_n15275 ^ new_n15244;
  assign new_n15277 = new_n15276 ^ new_n15252;
  assign new_n15278 = ~new_n15277 & new_n15253;
  assign new_n15279 = new_n15278 ^ new_n15273;
  assign new_n15280 = new_n15276 ^ new_n15269;
  assign new_n15281 = new_n15280 ^ new_n15268;
  assign new_n15282 = ~new_n15281 & new_n15219;
  assign new_n15283 = new_n15183 ^ new_n15102;
  assign new_n15284 = new_n15246 ^ new_n15220;
  assign new_n15285 = new_n15264 ^ new_n15262;
  assign new_n15286 = new_n15285 ^ new_n15243;
  assign new_n15287 = new_n15275 ^ new_n15260;
  assign new_n15288 = new_n15286 & new_n15287;
  assign new_n15289 = new_n15288 ^ new_n15276;
  assign new_n15290 = new_n15289 ^ new_n15284;
  assign new_n15291 = new_n15290 ^ new_n15283;
  assign new_n15292 = new_n15291 ^ new_n15199;
  assign new_n15293 = new_n15262 ^ new_n15238;
  assign new_n15294 = new_n15293 ^ new_n15255;
  assign new_n15295 = new_n15294 ^ new_n15292;
  assign new_n15296 = ~new_n15295 & new_n15226;
  assign new_n15297 = new_n15200 & new_n15272;
  assign new_n15298 = new_n15297 ^ new_n15296;
  assign new_n15299 = new_n15298 ^ new_n15282;
  assign new_n15300 = new_n15288 ^ new_n15232;
  assign new_n15301 = new_n15216 & new_n15300;
  assign new_n15302 = new_n15301 ^ new_n15299;
  assign new_n15303 = new_n15288 ^ new_n15262;
  assign new_n15304 = new_n15303 ^ new_n15259;
  assign new_n15305 = new_n15237 & new_n15304;
  assign new_n15306 = new_n15305 ^ new_n15302;
  assign new_n15307 = ~new_n15295 & new_n15228;
  assign new_n15308 = new_n15307 ^ new_n15306;
  assign new_n15309 = new_n15308 ^ new_n15279;
  assign new_n15310 = new_n12409 ^ new_n12403;
  assign new_n15311 = new_n15310 ^ new_n12499;
  assign new_n15312 = new_n13550 ^ n27;
  assign new_n15313 = new_n15312 ^ new_n12463;
  assign new_n15314 = new_n15313 ^ new_n15311;
  assign new_n15315 = new_n13572 ^ n26;
  assign new_n15316 = new_n15315 ^ new_n12513;
  assign new_n15317 = new_n12499 ^ new_n12428;
  assign new_n15318 = new_n15317 ^ new_n12635;
  assign new_n15319 = new_n15318 ^ new_n15316;
  assign new_n15320 = new_n15319 ^ new_n15314;
  assign new_n15321 = new_n12638 ^ new_n12143;
  assign new_n15322 = new_n13640 ^ n31;
  assign new_n15323 = new_n15322 ^ new_n15321;
  assign new_n15324 = new_n12577 ^ new_n12555;
  assign new_n15325 = new_n15324 ^ new_n15323;
  assign new_n15326 = new_n12600 ^ new_n12572;
  assign new_n15327 = new_n15326 ^ new_n12533;
  assign new_n15328 = new_n15327 ^ new_n15325;
  assign new_n15329 = new_n13684 ^ n29;
  assign new_n15330 = new_n15329 ^ new_n15321;
  assign new_n15331 = new_n12620 ^ new_n12265;
  assign new_n15332 = new_n15331 ^ new_n15330;
  assign new_n15333 = new_n12585 ^ new_n12258;
  assign new_n15334 = new_n15333 ^ new_n12611;
  assign new_n15335 = new_n15334 ^ new_n15332;
  assign new_n15336 = new_n15335 ^ new_n15328;
  assign new_n15337 = new_n13713 ^ n25;
  assign new_n15338 = new_n15337 ^ new_n12642;
  assign new_n15339 = new_n12635 ^ new_n12504;
  assign new_n15340 = new_n15339 ^ new_n12143;
  assign new_n15341 = new_n15340 ^ new_n15338;
  assign new_n15342 = new_n15321 ^ new_n11990;
  assign new_n15343 = new_n12868 ^ n28;
  assign new_n15344 = new_n15343 ^ new_n15342;
  assign new_n15345 = new_n12616 ^ new_n12409;
  assign new_n15346 = new_n15345 ^ new_n12258;
  assign new_n15347 = new_n15346 ^ new_n15344;
  assign new_n15348 = new_n15347 ^ new_n15341;
  assign new_n15349 = new_n15348 ^ new_n15336;
  assign new_n15350 = new_n15349 ^ new_n15320;
  assign new_n15351 = new_n15321 ^ new_n12572;
  assign new_n15352 = new_n12539 ^ new_n12526;
  assign new_n15353 = new_n13601 ^ n32;
  assign new_n15354 = new_n15353 ^ new_n15352;
  assign new_n15355 = new_n15354 ^ new_n15351;
  assign new_n15356 = new_n15355 ^ new_n15320;
  assign new_n15357 = new_n15356 ^ new_n15347;
  assign new_n15358 = new_n15355 & new_n15357;
  assign new_n15359 = new_n15358 ^ new_n15347;
  assign new_n15360 = new_n15347 ^ new_n15328;
  assign new_n15361 = new_n12611 ^ new_n12600;
  assign new_n15362 = new_n15361 ^ new_n12559;
  assign new_n15363 = new_n12604 ^ new_n12589;
  assign new_n15364 = new_n13669 ^ n30;
  assign new_n15365 = new_n15364 ^ new_n15363;
  assign new_n15366 = new_n15365 ^ new_n15362;
  assign new_n15367 = new_n15366 ^ new_n15341;
  assign new_n15368 = new_n15367 ^ new_n15360;
  assign new_n15369 = ~new_n15349 & new_n15368;
  assign new_n15370 = new_n15369 ^ new_n15319;
  assign new_n15371 = new_n15370 ^ new_n15359;
  assign new_n15372 = ~new_n15328 & ~new_n15356;
  assign new_n15373 = new_n15372 ^ new_n15328;
  assign new_n15374 = new_n15366 ^ new_n15336;
  assign new_n15375 = new_n15374 ^ new_n15314;
  assign new_n15376 = new_n15341 ^ new_n15328;
  assign new_n15377 = ~new_n15375 & new_n15376;
  assign new_n15378 = new_n15377 ^ new_n15373;
  assign new_n15379 = new_n15378 ^ new_n15367;
  assign new_n15380 = new_n15347 ^ new_n15314;
  assign new_n15381 = new_n15380 ^ new_n15367;
  assign new_n15382 = new_n15366 ^ new_n15347;
  assign new_n15383 = new_n15381 & new_n15382;
  assign new_n15384 = new_n15374 ^ new_n15319;
  assign new_n15385 = ~new_n15384 & new_n15348;
  assign new_n15386 = new_n15385 ^ new_n15383;
  assign new_n15387 = new_n15335 ^ new_n15314;
  assign new_n15388 = new_n15387 ^ new_n15386;
  assign new_n15389 = new_n15388 ^ new_n15379;
  assign new_n15390 = new_n15370 ^ new_n15349;
  assign new_n15391 = new_n15355 ^ new_n15349;
  assign new_n15392 = new_n15356 ^ new_n15328;
  assign new_n15393 = new_n15392 ^ new_n15367;
  assign new_n15394 = ~new_n15391 & new_n15393;
  assign new_n15395 = new_n15394 ^ new_n15386;
  assign new_n15396 = new_n15395 ^ new_n15366;
  assign new_n15397 = new_n15396 ^ new_n15390;
  assign new_n15398 = ~new_n15397 & new_n15389;
  assign new_n15399 = new_n15398 ^ new_n15371;
  assign new_n15400 = ~new_n15350 & new_n15367;
  assign new_n15401 = new_n15400 ^ new_n15385;
  assign new_n15402 = new_n15401 ^ new_n15375;
  assign new_n15403 = new_n15402 ^ new_n15399;
  assign new_n15404 = new_n15400 ^ new_n15383;
  assign new_n15405 = new_n15384 ^ new_n15355;
  assign new_n15406 = new_n15356 ^ new_n15341;
  assign new_n15407 = ~new_n15405 & new_n15406;
  assign new_n15408 = new_n15407 ^ new_n15372;
  assign new_n15409 = new_n15408 ^ new_n15404;
  assign new_n15410 = ~new_n15403 & ~new_n15409;
  assign new_n15411 = new_n15410 ^ new_n15341;
  assign new_n15412 = new_n15407 ^ new_n15358;
  assign new_n15413 = new_n15328 ^ new_n15314;
  assign new_n15414 = new_n15394 ^ new_n15373;
  assign new_n15415 = new_n15407 ^ new_n15377;
  assign new_n15416 = new_n15415 ^ new_n15341;
  assign new_n15417 = new_n15416 ^ new_n15402;
  assign new_n15418 = new_n15410 ^ new_n15398;
  assign new_n15419 = ~new_n15418 & new_n15417;
  assign new_n15420 = new_n15419 ^ new_n15410;
  assign new_n15421 = new_n15417 ^ new_n15398;
  assign new_n15422 = new_n15341 ^ new_n15314;
  assign new_n15423 = new_n15394 ^ new_n15358;
  assign new_n15424 = new_n15423 ^ new_n15404;
  assign new_n15425 = new_n15424 ^ new_n15422;
  assign new_n15426 = ~new_n15421 & new_n15425;
  assign new_n15427 = new_n15426 ^ new_n15371;
  assign new_n15428 = new_n15427 ^ new_n15402;
  assign new_n15429 = ~new_n15420 & ~new_n15428;
  assign new_n15430 = new_n15421 ^ new_n15420;
  assign new_n15431 = new_n15430 ^ new_n15429;
  assign new_n15432 = new_n15431 ^ new_n15414;
  assign new_n15433 = new_n15432 ^ new_n15413;
  assign new_n15434 = new_n15433 ^ new_n15412;
  assign new_n15435 = new_n15434 ^ new_n15411;
  assign new_n15436 = ~new_n15350 & ~new_n15435;
  assign new_n15437 = new_n15429 ^ new_n15426;
  assign new_n15438 = new_n15437 ^ new_n15397;
  assign new_n15439 = ~new_n15438 & new_n15376;
  assign new_n15440 = new_n15439 ^ new_n15436;
  assign new_n15441 = new_n15429 ^ new_n15425;
  assign new_n15442 = new_n15356 & new_n15441;
  assign new_n15443 = new_n15433 ^ new_n15347;
  assign new_n15444 = new_n15426 ^ new_n15377;
  assign new_n15445 = new_n15444 ^ new_n15370;
  assign new_n15446 = new_n15445 ^ new_n15443;
  assign new_n15447 = ~new_n15446 & new_n15381;
  assign new_n15448 = new_n15447 ^ new_n15442;
  assign new_n15449 = new_n15392 & new_n15441;
  assign new_n15450 = ~new_n15405 & ~new_n15428;
  assign new_n15451 = new_n15450 ^ new_n15449;
  assign new_n15452 = ~new_n15446 & new_n15382;
  assign new_n15453 = new_n15426 ^ new_n15410;
  assign new_n15454 = new_n15416 ^ new_n15371;
  assign new_n15455 = new_n15454 ^ new_n15453;
  assign new_n15456 = new_n15348 & new_n15455;
  assign new_n15457 = new_n15456 ^ new_n15452;
  assign new_n15458 = new_n15457 ^ new_n15451;
  assign new_n15459 = new_n15458 ^ new_n15448;
  assign new_n15460 = new_n15459 ^ new_n15440;
  assign new_n15461 = new_n13531 ^ new_n13515;
  assign new_n15462 = new_n15461 ^ new_n13588;
  assign new_n15463 = new_n11732 ^ new_n10299;
  assign new_n15464 = new_n13555 ^ new_n13168;
  assign new_n15465 = new_n15464 ^ new_n15463;
  assign new_n15466 = new_n15465 ^ new_n15462;
  assign new_n15467 = new_n13592 ^ new_n13566;
  assign new_n15468 = new_n15467 ^ new_n13497;
  assign new_n15469 = new_n11738 ^ new_n11407;
  assign new_n15470 = new_n15469 ^ new_n13718;
  assign new_n15471 = new_n15470 ^ new_n13588;
  assign new_n15472 = new_n15471 ^ new_n15468;
  assign new_n15473 = new_n15472 ^ new_n15466;
  assign new_n15474 = new_n13707 ^ new_n13316;
  assign new_n15475 = new_n15474 ^ new_n13614;
  assign new_n15476 = new_n13651 ^ new_n13629;
  assign new_n15477 = new_n15476 ^ new_n15475;
  assign new_n15478 = new_n11710 ^ new_n11536;
  assign new_n15479 = new_n15478 ^ new_n13678;
  assign new_n15480 = new_n15479 ^ new_n13646;
  assign new_n15481 = new_n15480 ^ new_n15477;
  assign new_n15482 = new_n13659 ^ new_n13477;
  assign new_n15483 = new_n15482 ^ new_n13700;
  assign new_n15484 = new_n11717 ^ new_n11503;
  assign new_n15485 = new_n15484 ^ new_n15474;
  assign new_n15486 = new_n13693 ^ new_n13468;
  assign new_n15487 = new_n15486 ^ new_n15485;
  assign new_n15488 = new_n15487 ^ new_n15483;
  assign new_n15489 = new_n15488 ^ new_n15481;
  assign new_n15490 = new_n13709 ^ new_n13454;
  assign new_n15491 = new_n15490 ^ new_n13562;
  assign new_n15492 = new_n11702 ^ new_n11559;
  assign new_n15493 = new_n15492 ^ new_n13316;
  assign new_n15494 = new_n15493 ^ new_n13718;
  assign new_n15495 = new_n15494 ^ new_n15491;
  assign new_n15496 = new_n11693 ^ new_n11464;
  assign new_n15497 = new_n13461 ^ new_n13016;
  assign new_n15498 = new_n15497 ^ new_n15496;
  assign new_n15499 = new_n15498 ^ new_n15474;
  assign new_n15500 = new_n13689 ^ new_n13555;
  assign new_n15501 = new_n15500 ^ new_n13477;
  assign new_n15502 = new_n15501 ^ new_n15499;
  assign new_n15503 = new_n15502 ^ new_n15495;
  assign new_n15504 = new_n15503 ^ new_n15489;
  assign new_n15505 = new_n15504 ^ new_n15473;
  assign new_n15506 = new_n13673 ^ new_n13663;
  assign new_n15507 = new_n15506 ^ new_n13633;
  assign new_n15508 = new_n11725 ^ new_n11581;
  assign new_n15509 = new_n15508 ^ new_n13700;
  assign new_n15510 = new_n15509 ^ new_n13678;
  assign new_n15511 = new_n15510 ^ new_n15507;
  assign new_n15512 = new_n15511 ^ new_n15502;
  assign new_n15513 = new_n15495 ^ new_n15481;
  assign new_n15514 = new_n15513 ^ new_n15512;
  assign new_n15515 = ~new_n15504 & ~new_n15514;
  assign new_n15516 = new_n15515 ^ new_n15472;
  assign new_n15517 = new_n15516 ^ new_n15504;
  assign new_n15518 = new_n11754 ^ new_n11424;
  assign new_n15519 = new_n15518 ^ new_n13646;
  assign new_n15520 = new_n13620 ^ new_n13607;
  assign new_n15521 = new_n15520 ^ new_n15474;
  assign new_n15522 = new_n15521 ^ new_n15519;
  assign new_n15523 = new_n15522 ^ new_n15504;
  assign new_n15524 = new_n15522 ^ new_n15473;
  assign new_n15525 = new_n15524 ^ new_n15481;
  assign new_n15526 = new_n15511 ^ new_n15495;
  assign new_n15527 = new_n15526 ^ new_n15525;
  assign new_n15528 = new_n15523 & new_n15527;
  assign new_n15529 = new_n15511 ^ new_n15489;
  assign new_n15530 = new_n15529 ^ new_n15472;
  assign new_n15531 = new_n15503 & new_n15530;
  assign new_n15532 = new_n15531 ^ new_n15528;
  assign new_n15533 = new_n15502 ^ new_n15466;
  assign new_n15534 = new_n15533 ^ new_n15526;
  assign new_n15535 = ~new_n15534 & new_n15512;
  assign new_n15536 = new_n15535 ^ new_n15511;
  assign new_n15537 = new_n15536 ^ new_n15532;
  assign new_n15538 = new_n15537 ^ new_n15517;
  assign new_n15539 = new_n15481 & new_n15524;
  assign new_n15540 = new_n15539 ^ new_n15481;
  assign new_n15541 = new_n15529 ^ new_n15466;
  assign new_n15542 = ~new_n15513 & new_n15541;
  assign new_n15543 = new_n15542 ^ new_n15540;
  assign new_n15544 = new_n15543 ^ new_n15526;
  assign new_n15545 = new_n15535 ^ new_n15531;
  assign new_n15546 = new_n15488 ^ new_n15466;
  assign new_n15547 = new_n15546 ^ new_n15545;
  assign new_n15548 = new_n15547 ^ new_n15544;
  assign new_n15549 = ~new_n15548 & new_n15538;
  assign new_n15550 = new_n15524 ^ new_n15502;
  assign new_n15551 = ~new_n15522 & ~new_n15550;
  assign new_n15552 = new_n15551 ^ new_n15502;
  assign new_n15553 = new_n15552 ^ new_n15516;
  assign new_n15554 = new_n15553 ^ new_n15549;
  assign new_n15555 = ~new_n15505 & new_n15526;
  assign new_n15556 = new_n15555 ^ new_n15531;
  assign new_n15557 = new_n15556 ^ new_n15541;
  assign new_n15558 = new_n15557 ^ new_n15554;
  assign new_n15559 = new_n15555 ^ new_n15535;
  assign new_n15560 = new_n15530 ^ new_n15522;
  assign new_n15561 = new_n15524 ^ new_n15495;
  assign new_n15562 = ~new_n15560 & ~new_n15561;
  assign new_n15563 = new_n15562 ^ new_n15539;
  assign new_n15564 = new_n15563 ^ new_n15559;
  assign new_n15565 = ~new_n15558 & ~new_n15564;
  assign new_n15566 = new_n15565 ^ new_n15495;
  assign new_n15567 = new_n15562 ^ new_n15551;
  assign new_n15568 = new_n15481 ^ new_n15466;
  assign new_n15569 = new_n15540 ^ new_n15528;
  assign new_n15570 = new_n15495 ^ new_n15466;
  assign new_n15571 = new_n15551 ^ new_n15528;
  assign new_n15572 = new_n15571 ^ new_n15559;
  assign new_n15573 = new_n15572 ^ new_n15570;
  assign new_n15574 = new_n15562 ^ new_n15542;
  assign new_n15575 = new_n15574 ^ new_n15495;
  assign new_n15576 = new_n15575 ^ new_n15557;
  assign new_n15577 = new_n15576 ^ new_n15549;
  assign new_n15578 = ~new_n15573 & new_n15577;
  assign new_n15579 = new_n15578 ^ new_n15553;
  assign new_n15580 = new_n15579 ^ new_n15557;
  assign new_n15581 = new_n15565 ^ new_n15549;
  assign new_n15582 = ~new_n15581 & new_n15576;
  assign new_n15583 = new_n15582 ^ new_n15549;
  assign new_n15584 = ~new_n15580 & new_n15583;
  assign new_n15585 = new_n15582 ^ new_n15576;
  assign new_n15586 = new_n15585 ^ new_n15584;
  assign new_n15587 = new_n15586 ^ new_n15569;
  assign new_n15588 = new_n15587 ^ new_n15568;
  assign new_n15589 = new_n15588 ^ new_n15567;
  assign new_n15590 = new_n15589 ^ new_n15566;
  assign new_n15591 = ~new_n15505 & new_n15590;
  assign new_n15592 = new_n15584 ^ new_n15578;
  assign new_n15593 = new_n15592 ^ new_n15538;
  assign new_n15594 = ~new_n15513 & new_n15593;
  assign new_n15595 = new_n15594 ^ new_n15591;
  assign new_n15596 = new_n15584 ^ new_n15573;
  assign new_n15597 = ~new_n15524 & ~new_n15596;
  assign new_n15598 = new_n15588 ^ new_n15502;
  assign new_n15599 = new_n15578 ^ new_n15542;
  assign new_n15600 = new_n15599 ^ new_n15516;
  assign new_n15601 = new_n15600 ^ new_n15598;
  assign new_n15602 = ~new_n15534 & ~new_n15601;
  assign new_n15603 = new_n15602 ^ new_n15597;
  assign new_n15604 = ~new_n15596 & new_n15525;
  assign new_n15605 = ~new_n15560 & ~new_n15580;
  assign new_n15606 = new_n15605 ^ new_n15604;
  assign new_n15607 = ~new_n15601 & new_n15512;
  assign new_n15608 = new_n15578 ^ new_n15565;
  assign new_n15609 = new_n15575 ^ new_n15553;
  assign new_n15610 = new_n15609 ^ new_n15608;
  assign new_n15611 = ~new_n15610 & new_n15503;
  assign new_n15612 = new_n15611 ^ new_n15607;
  assign new_n15613 = new_n15612 ^ new_n15606;
  assign new_n15614 = new_n15613 ^ new_n15603;
  assign new_n15615 = new_n15614 ^ new_n15595;
  assign new_n15616 = new_n15615 ^ new_n15460;
  assign new_n15617 = new_n15315 ^ new_n15312;
  assign new_n15618 = new_n15617 ^ new_n15353;
  assign new_n15619 = new_n15618 ^ new_n15343;
  assign new_n15620 = new_n15322 & new_n15618;
  assign new_n15621 = new_n15620 ^ new_n15322;
  assign new_n15622 = new_n15337 ^ new_n15322;
  assign new_n15623 = new_n15329 ^ new_n15322;
  assign new_n15624 = new_n15623 ^ new_n15364;
  assign new_n15625 = new_n15624 ^ new_n15312;
  assign new_n15626 = ~new_n15622 & ~new_n15625;
  assign new_n15627 = new_n15626 ^ new_n15621;
  assign new_n15628 = new_n15364 ^ new_n15337;
  assign new_n15629 = new_n15628 ^ new_n15627;
  assign new_n15630 = new_n15343 ^ new_n15312;
  assign new_n15631 = new_n15630 ^ new_n15628;
  assign new_n15632 = new_n15364 ^ new_n15343;
  assign new_n15633 = ~new_n15631 & new_n15632;
  assign new_n15634 = new_n15343 ^ new_n15337;
  assign new_n15635 = new_n15624 ^ new_n15315;
  assign new_n15636 = ~new_n15635 & new_n15634;
  assign new_n15637 = new_n15636 ^ new_n15633;
  assign new_n15638 = new_n15329 ^ new_n15312;
  assign new_n15639 = new_n15638 ^ new_n15637;
  assign new_n15640 = new_n15639 ^ new_n15629;
  assign new_n15641 = new_n15634 ^ new_n15623;
  assign new_n15642 = new_n15343 ^ new_n15322;
  assign new_n15643 = new_n15642 ^ new_n15628;
  assign new_n15644 = ~new_n15643 & new_n15641;
  assign new_n15645 = new_n15644 ^ new_n15315;
  assign new_n15646 = new_n15645 ^ new_n15641;
  assign new_n15647 = new_n15641 ^ new_n15353;
  assign new_n15648 = new_n15618 ^ new_n15322;
  assign new_n15649 = new_n15648 ^ new_n15628;
  assign new_n15650 = ~new_n15647 & new_n15649;
  assign new_n15651 = new_n15650 ^ new_n15364;
  assign new_n15652 = new_n15651 ^ new_n15637;
  assign new_n15653 = new_n15652 ^ new_n15646;
  assign new_n15654 = ~new_n15653 & new_n15640;
  assign new_n15655 = ~new_n15353 & ~new_n15619;
  assign new_n15656 = new_n15655 ^ new_n15343;
  assign new_n15657 = new_n15656 ^ new_n15645;
  assign new_n15658 = new_n15657 ^ new_n15654;
  assign new_n15659 = new_n15641 ^ new_n15617;
  assign new_n15660 = new_n15628 & new_n15659;
  assign new_n15661 = new_n15660 ^ new_n15636;
  assign new_n15662 = new_n15661 ^ new_n15625;
  assign new_n15663 = new_n15662 ^ new_n15658;
  assign new_n15664 = new_n15660 ^ new_n15633;
  assign new_n15665 = new_n15618 ^ new_n15337;
  assign new_n15666 = new_n15635 ^ new_n15353;
  assign new_n15667 = ~new_n15665 & new_n15666;
  assign new_n15668 = new_n15667 ^ new_n15620;
  assign new_n15669 = new_n15668 ^ new_n15664;
  assign new_n15670 = ~new_n15669 & new_n15663;
  assign new_n15671 = new_n15667 ^ new_n15626;
  assign new_n15672 = new_n15671 ^ new_n15337;
  assign new_n15673 = new_n15672 ^ new_n15662;
  assign new_n15674 = new_n15673 ^ new_n15670;
  assign new_n15675 = ~new_n15619 & ~new_n15674;
  assign new_n15676 = new_n15337 ^ new_n15312;
  assign new_n15677 = new_n15655 ^ new_n15650;
  assign new_n15678 = new_n15677 ^ new_n15664;
  assign new_n15679 = new_n15678 ^ new_n15676;
  assign new_n15680 = new_n15673 ^ new_n15654;
  assign new_n15681 = ~new_n15679 & ~new_n15680;
  assign new_n15682 = new_n15681 ^ new_n15657;
  assign new_n15683 = new_n15682 ^ new_n15662;
  assign new_n15684 = new_n15670 ^ new_n15654;
  assign new_n15685 = ~new_n15673 & ~new_n15684;
  assign new_n15686 = new_n15685 ^ new_n15654;
  assign new_n15687 = new_n15683 & new_n15686;
  assign new_n15688 = new_n15687 ^ new_n15679;
  assign new_n15689 = ~new_n15618 & ~new_n15688;
  assign new_n15690 = new_n15685 ^ new_n15673;
  assign new_n15691 = new_n15690 ^ new_n15670;
  assign new_n15692 = new_n15691 ^ new_n15669;
  assign new_n15693 = new_n15649 & new_n15692;
  assign new_n15694 = new_n15322 ^ new_n15312;
  assign new_n15695 = new_n15650 ^ new_n15621;
  assign new_n15696 = new_n15690 ^ new_n15687;
  assign new_n15697 = new_n15696 ^ new_n15695;
  assign new_n15698 = new_n15697 ^ new_n15694;
  assign new_n15699 = new_n15698 ^ new_n15343;
  assign new_n15700 = new_n15681 ^ new_n15626;
  assign new_n15701 = new_n15700 ^ new_n15645;
  assign new_n15702 = new_n15701 ^ new_n15699;
  assign new_n15703 = new_n15632 & new_n15702;
  assign new_n15704 = new_n15681 ^ new_n15670;
  assign new_n15705 = new_n15672 ^ new_n15657;
  assign new_n15706 = new_n15705 ^ new_n15704;
  assign new_n15707 = ~new_n15706 & new_n15634;
  assign new_n15708 = new_n15707 ^ new_n15703;
  assign new_n15709 = new_n15708 ^ new_n15693;
  assign new_n15710 = new_n15709 ^ new_n15689;
  assign new_n15711 = new_n15687 ^ new_n15681;
  assign new_n15712 = new_n15711 ^ new_n15653;
  assign new_n15713 = ~new_n15625 & ~new_n15712;
  assign new_n15714 = new_n15713 ^ new_n15710;
  assign new_n15715 = ~new_n15631 & new_n15702;
  assign new_n15716 = new_n15715 ^ new_n15714;
  assign new_n15717 = new_n15716 ^ new_n15675;
  assign new_n15718 = new_n15670 ^ new_n15337;
  assign new_n15719 = new_n15667 ^ new_n15655;
  assign new_n15720 = new_n15719 ^ new_n15698;
  assign new_n15721 = new_n15720 ^ new_n15718;
  assign new_n15722 = ~new_n15721 & new_n15659;
  assign new_n15723 = ~new_n15665 & new_n15683;
  assign new_n15724 = new_n15723 ^ new_n15722;
  assign new_n15725 = ~new_n15622 & ~new_n15712;
  assign new_n15726 = ~new_n15353 & ~new_n15674;
  assign new_n15727 = new_n15690 ^ new_n15640;
  assign new_n15728 = ~new_n15727 & new_n15641;
  assign new_n15729 = new_n15728 ^ new_n15726;
  assign new_n15730 = new_n15729 ^ new_n15725;
  assign new_n15731 = new_n15730 ^ new_n15724;
  assign new_n15732 = new_n15731 ^ new_n15717;
  assign new_n15733 = new_n15732 ^ new_n425;
  assign new_n15734 = new_n15733 ^ new_n15616;
  assign new_n15735 = new_n15417 ^ new_n15410;
  assign new_n15736 = ~new_n15735 & new_n15357;
  assign new_n15737 = new_n15430 ^ new_n15410;
  assign new_n15738 = new_n15737 ^ new_n15409;
  assign new_n15739 = ~new_n15738 & new_n15393;
  assign new_n15740 = new_n15739 ^ new_n15457;
  assign new_n15741 = new_n15740 ^ new_n15442;
  assign new_n15742 = ~new_n15375 & ~new_n15438;
  assign new_n15743 = new_n15742 ^ new_n15741;
  assign new_n15744 = new_n15743 ^ new_n15447;
  assign new_n15745 = new_n15744 ^ new_n15736;
  assign new_n15746 = ~new_n15428 & new_n15406;
  assign new_n15747 = new_n15746 ^ new_n15436;
  assign new_n15748 = ~new_n15735 & new_n15355;
  assign new_n15749 = new_n15430 ^ new_n15389;
  assign new_n15750 = ~new_n15349 & new_n15749;
  assign new_n15751 = new_n15750 ^ new_n15748;
  assign new_n15752 = new_n15751 ^ new_n15439;
  assign new_n15753 = new_n15752 ^ new_n15747;
  assign new_n15754 = new_n15753 ^ new_n15745;
  assign new_n15755 = new_n14848 ^ new_n540;
  assign new_n15756 = new_n11548 ^ new_n11453;
  assign new_n15757 = new_n15756 ^ new_n15755;
  assign new_n15758 = new_n11509 ^ new_n11481;
  assign new_n15759 = new_n15758 ^ new_n15757;
  assign new_n15760 = new_n11473 ^ new_n11330;
  assign new_n15761 = new_n15760 ^ new_n11310;
  assign new_n15762 = new_n15761 ^ new_n15759;
  assign new_n15763 = new_n11469 ^ new_n11310;
  assign new_n15764 = new_n15763 ^ new_n11388;
  assign new_n15765 = new_n14675 ^ new_n560;
  assign new_n15766 = new_n15765 ^ new_n8060;
  assign new_n15767 = new_n15766 ^ new_n10181;
  assign new_n15768 = new_n15767 ^ new_n15764;
  assign new_n15769 = new_n11388 ^ new_n9161;
  assign new_n15770 = new_n15769 ^ new_n11555;
  assign new_n15771 = new_n14097 ^ new_n566;
  assign new_n15772 = new_n15771 ^ new_n11369;
  assign new_n15773 = new_n15772 ^ new_n11412;
  assign new_n15774 = new_n15773 ^ new_n15770;
  assign new_n15775 = new_n15774 ^ new_n15768;
  assign new_n15776 = new_n15756 ^ new_n11521;
  assign new_n15777 = new_n14877 ^ new_n575;
  assign new_n15778 = new_n15777 ^ new_n11448;
  assign new_n15779 = new_n15778 ^ new_n11431;
  assign new_n15780 = new_n15779 ^ new_n15776;
  assign new_n15781 = new_n15780 ^ new_n15775;
  assign new_n15782 = new_n15781 ^ new_n15762;
  assign new_n15783 = new_n14857 ^ new_n584;
  assign new_n15784 = new_n11555 ^ new_n11351;
  assign new_n15785 = new_n15784 ^ new_n15783;
  assign new_n15786 = new_n11551 ^ new_n11456;
  assign new_n15787 = new_n15786 ^ new_n11453;
  assign new_n15788 = new_n15787 ^ new_n15785;
  assign new_n15789 = new_n15788 ^ new_n15762;
  assign new_n15790 = new_n11513 ^ new_n11481;
  assign new_n15791 = new_n15790 ^ new_n11486;
  assign new_n15792 = new_n14809 ^ new_n597;
  assign new_n15793 = new_n15792 ^ new_n15756;
  assign new_n15794 = new_n11568 ^ new_n11497;
  assign new_n15795 = new_n15794 ^ new_n15793;
  assign new_n15796 = new_n15795 ^ new_n15791;
  assign new_n15797 = new_n15756 ^ new_n11576;
  assign new_n15798 = new_n11521 ^ new_n11440;
  assign new_n15799 = new_n15798 ^ new_n15797;
  assign new_n15800 = new_n14791 ^ new_n591;
  assign new_n15801 = new_n15800 ^ new_n11530;
  assign new_n15802 = new_n15801 ^ new_n11541;
  assign new_n15803 = new_n15802 ^ new_n15799;
  assign new_n15804 = new_n15803 ^ new_n15796;
  assign new_n15805 = new_n15804 ^ new_n15789;
  assign new_n15806 = new_n11571 ^ new_n11497;
  assign new_n15807 = new_n15806 ^ new_n11494;
  assign new_n15808 = new_n14079 ^ new_n605;
  assign new_n15809 = new_n11576 ^ new_n11526;
  assign new_n15810 = new_n15809 ^ new_n15808;
  assign new_n15811 = new_n15810 ^ new_n15807;
  assign new_n15812 = new_n15811 ^ new_n15762;
  assign new_n15813 = new_n15803 ^ new_n15788;
  assign new_n15814 = new_n15813 ^ new_n15812;
  assign new_n15815 = ~new_n15805 & ~new_n15814;
  assign new_n15816 = new_n15815 ^ new_n15774;
  assign new_n15817 = new_n15816 ^ new_n15805;
  assign new_n15818 = new_n15811 ^ new_n15804;
  assign new_n15819 = new_n15818 ^ new_n15774;
  assign new_n15820 = new_n15789 & new_n15819;
  assign new_n15821 = new_n15805 ^ new_n15780;
  assign new_n15822 = new_n15803 ^ new_n15781;
  assign new_n15823 = new_n15811 ^ new_n15788;
  assign new_n15824 = new_n15823 ^ new_n15822;
  assign new_n15825 = new_n15821 & new_n15824;
  assign new_n15826 = new_n15825 ^ new_n15820;
  assign new_n15827 = new_n15768 ^ new_n15762;
  assign new_n15828 = new_n15827 ^ new_n15823;
  assign new_n15829 = ~new_n15828 & new_n15812;
  assign new_n15830 = new_n15829 ^ new_n15811;
  assign new_n15831 = new_n15830 ^ new_n15826;
  assign new_n15832 = new_n15831 ^ new_n15817;
  assign new_n15833 = new_n15781 & new_n15803;
  assign new_n15834 = new_n15833 ^ new_n15803;
  assign new_n15835 = new_n15818 ^ new_n15768;
  assign new_n15836 = ~new_n15813 & new_n15835;
  assign new_n15837 = new_n15836 ^ new_n15834;
  assign new_n15838 = new_n15837 ^ new_n15823;
  assign new_n15839 = new_n15829 ^ new_n15820;
  assign new_n15840 = new_n15796 ^ new_n15768;
  assign new_n15841 = new_n15840 ^ new_n15839;
  assign new_n15842 = new_n15841 ^ new_n15838;
  assign new_n15843 = ~new_n15842 & new_n15832;
  assign new_n15844 = ~new_n15780 & ~new_n15782;
  assign new_n15845 = new_n15844 ^ new_n15762;
  assign new_n15846 = new_n15845 ^ new_n15816;
  assign new_n15847 = new_n15846 ^ new_n15843;
  assign new_n15848 = new_n15805 ^ new_n15775;
  assign new_n15849 = ~new_n15848 & new_n15823;
  assign new_n15850 = new_n15849 ^ new_n15820;
  assign new_n15851 = new_n15850 ^ new_n15835;
  assign new_n15852 = new_n15851 ^ new_n15847;
  assign new_n15853 = new_n15819 ^ new_n15780;
  assign new_n15854 = new_n15788 ^ new_n15781;
  assign new_n15855 = ~new_n15853 & ~new_n15854;
  assign new_n15856 = new_n15855 ^ new_n15833;
  assign new_n15857 = new_n15849 ^ new_n15829;
  assign new_n15858 = new_n15857 ^ new_n15856;
  assign new_n15859 = ~new_n15852 & ~new_n15858;
  assign new_n15860 = new_n15855 ^ new_n15836;
  assign new_n15861 = new_n15860 ^ new_n15788;
  assign new_n15862 = new_n15861 ^ new_n15851;
  assign new_n15863 = new_n15862 ^ new_n15859;
  assign new_n15864 = ~new_n15782 & new_n15863;
  assign new_n15865 = new_n15803 ^ new_n15768;
  assign new_n15866 = new_n15834 ^ new_n15825;
  assign new_n15867 = new_n15788 ^ new_n15768;
  assign new_n15868 = new_n15844 ^ new_n15825;
  assign new_n15869 = new_n15868 ^ new_n15857;
  assign new_n15870 = new_n15869 ^ new_n15867;
  assign new_n15871 = new_n15862 ^ new_n15843;
  assign new_n15872 = ~new_n15870 & new_n15871;
  assign new_n15873 = new_n15872 ^ new_n15846;
  assign new_n15874 = new_n15873 ^ new_n15851;
  assign new_n15875 = new_n15859 ^ new_n15843;
  assign new_n15876 = ~new_n15875 & new_n15862;
  assign new_n15877 = new_n15876 ^ new_n15843;
  assign new_n15878 = ~new_n15874 & new_n15877;
  assign new_n15879 = new_n15876 ^ new_n15862;
  assign new_n15880 = new_n15879 ^ new_n15878;
  assign new_n15881 = new_n15880 ^ new_n15866;
  assign new_n15882 = new_n15881 ^ new_n15865;
  assign new_n15883 = new_n15882 ^ new_n15762;
  assign new_n15884 = new_n15872 ^ new_n15836;
  assign new_n15885 = new_n15884 ^ new_n15816;
  assign new_n15886 = new_n15885 ^ new_n15883;
  assign new_n15887 = ~new_n15828 & ~new_n15886;
  assign new_n15888 = new_n15878 ^ new_n15872;
  assign new_n15889 = new_n15888 ^ new_n15832;
  assign new_n15890 = new_n15835 & new_n15889;
  assign new_n15891 = new_n15878 ^ new_n15870;
  assign new_n15892 = ~new_n15781 & ~new_n15891;
  assign new_n15893 = ~new_n15886 & new_n15812;
  assign new_n15894 = new_n15872 ^ new_n15859;
  assign new_n15895 = new_n15861 ^ new_n15846;
  assign new_n15896 = new_n15895 ^ new_n15894;
  assign new_n15897 = ~new_n15896 & new_n15789;
  assign new_n15898 = new_n15897 ^ new_n15893;
  assign new_n15899 = new_n15879 ^ new_n15859;
  assign new_n15900 = new_n15899 ^ new_n15858;
  assign new_n15901 = ~new_n15900 & new_n15824;
  assign new_n15902 = new_n15901 ^ new_n15898;
  assign new_n15903 = new_n15902 ^ new_n15892;
  assign new_n15904 = new_n15903 ^ new_n15890;
  assign new_n15905 = new_n15904 ^ new_n15887;
  assign new_n15906 = new_n15905 ^ new_n15864;
  assign new_n15907 = ~new_n15854 & ~new_n15874;
  assign new_n15908 = new_n15859 ^ new_n15788;
  assign new_n15909 = new_n15855 ^ new_n15844;
  assign new_n15910 = new_n15909 ^ new_n15882;
  assign new_n15911 = new_n15910 ^ new_n15908;
  assign new_n15912 = ~new_n15848 & new_n15911;
  assign new_n15913 = new_n15912 ^ new_n15907;
  assign new_n15914 = new_n15879 ^ new_n15842;
  assign new_n15915 = ~new_n15805 & ~new_n15914;
  assign new_n15916 = ~new_n15780 & new_n15863;
  assign new_n15917 = new_n15916 ^ new_n15915;
  assign new_n15918 = ~new_n15813 & new_n15889;
  assign new_n15919 = new_n15918 ^ new_n15917;
  assign new_n15920 = new_n15919 ^ new_n15913;
  assign new_n15921 = new_n15920 ^ new_n15906;
  assign new_n15922 = new_n15921 ^ new_n15754;
  assign new_n15923 = new_n12248 ^ new_n12002;
  assign new_n15924 = new_n14861 ^ new_n14769;
  assign new_n15925 = new_n15924 ^ new_n15923;
  assign new_n15926 = new_n15925 ^ new_n14846;
  assign new_n15927 = new_n14841 ^ new_n14716;
  assign new_n15928 = new_n15927 ^ new_n14815;
  assign new_n15929 = new_n15928 ^ new_n15926;
  assign new_n15930 = new_n14743 ^ new_n14377;
  assign new_n15931 = new_n12481 ^ new_n12032;
  assign new_n15932 = new_n14852 ^ new_n14716;
  assign new_n15933 = new_n15932 ^ new_n15931;
  assign new_n15934 = new_n15933 ^ new_n15930;
  assign new_n15935 = new_n14669 ^ new_n14377;
  assign new_n15936 = new_n12517 ^ new_n12027;
  assign new_n15937 = new_n15936 ^ new_n14695;
  assign new_n15938 = new_n15937 ^ new_n14865;
  assign new_n15939 = new_n15938 ^ new_n15935;
  assign new_n15940 = new_n15939 ^ new_n15934;
  assign new_n15941 = new_n12546 ^ new_n12021;
  assign new_n15942 = new_n15941 ^ new_n14880;
  assign new_n15943 = new_n15924 ^ new_n14783;
  assign new_n15944 = new_n15943 ^ new_n15942;
  assign new_n15945 = new_n15944 ^ new_n15940;
  assign new_n15946 = new_n15945 ^ new_n15929;
  assign new_n15947 = new_n14802 ^ new_n14754;
  assign new_n15948 = new_n15947 ^ new_n15924;
  assign new_n15949 = new_n12565 ^ new_n11998;
  assign new_n15950 = new_n15949 ^ new_n14895;
  assign new_n15951 = new_n14883 ^ new_n14780;
  assign new_n15952 = new_n15951 ^ new_n15950;
  assign new_n15953 = new_n15952 ^ new_n15948;
  assign new_n15954 = new_n15945 & new_n15953;
  assign new_n15955 = new_n15954 ^ new_n15953;
  assign new_n15956 = new_n12594 ^ new_n12014;
  assign new_n15957 = new_n15956 ^ new_n14820;
  assign new_n15958 = new_n15957 ^ new_n14764;
  assign new_n15959 = new_n15958 ^ new_n14900;
  assign new_n15960 = new_n14841 ^ new_n14820;
  assign new_n15961 = new_n15960 ^ new_n14905;
  assign new_n15962 = new_n12626 ^ new_n12041;
  assign new_n15963 = new_n15962 ^ new_n15924;
  assign new_n15964 = new_n15963 ^ new_n14834;
  assign new_n15965 = new_n15964 ^ new_n15961;
  assign new_n15966 = new_n15965 ^ new_n15953;
  assign new_n15967 = new_n15966 ^ new_n15959;
  assign new_n15968 = new_n15967 ^ new_n15934;
  assign new_n15969 = new_n14870 ^ new_n14865;
  assign new_n15970 = new_n12644 ^ new_n12010;
  assign new_n15971 = new_n15970 ^ new_n14769;
  assign new_n15972 = new_n15971 ^ new_n14234;
  assign new_n15973 = new_n15972 ^ new_n15969;
  assign new_n15974 = new_n15973 ^ new_n15953;
  assign new_n15975 = ~new_n15974 & new_n15968;
  assign new_n15976 = new_n15975 ^ new_n15955;
  assign new_n15977 = new_n15973 ^ new_n15959;
  assign new_n15978 = new_n15977 ^ new_n15976;
  assign new_n15979 = new_n15967 ^ new_n15939;
  assign new_n15980 = new_n15973 ^ new_n15929;
  assign new_n15981 = new_n15979 & new_n15980;
  assign new_n15982 = new_n15959 ^ new_n15929;
  assign new_n15983 = new_n15934 ^ new_n15929;
  assign new_n15984 = new_n15983 ^ new_n15977;
  assign new_n15985 = ~new_n15984 & new_n15982;
  assign new_n15986 = new_n15985 ^ new_n15981;
  assign new_n15987 = new_n15965 ^ new_n15934;
  assign new_n15988 = new_n15987 ^ new_n15986;
  assign new_n15989 = new_n15988 ^ new_n15978;
  assign new_n15990 = new_n15980 ^ new_n15966;
  assign new_n15991 = new_n15953 ^ new_n15929;
  assign new_n15992 = new_n15991 ^ new_n15977;
  assign new_n15993 = ~new_n15990 & ~new_n15992;
  assign new_n15994 = new_n15993 ^ new_n15939;
  assign new_n15995 = new_n15994 ^ new_n15990;
  assign new_n15996 = new_n15990 ^ new_n15944;
  assign new_n15997 = new_n15953 ^ new_n15945;
  assign new_n15998 = new_n15997 ^ new_n15977;
  assign new_n15999 = new_n15996 & new_n15998;
  assign new_n16000 = new_n15999 ^ new_n15981;
  assign new_n16001 = new_n15985 ^ new_n15959;
  assign new_n16002 = new_n16001 ^ new_n16000;
  assign new_n16003 = new_n16002 ^ new_n15995;
  assign new_n16004 = ~new_n15989 & new_n16003;
  assign new_n16005 = ~new_n15944 & ~new_n15946;
  assign new_n16006 = new_n16005 ^ new_n15929;
  assign new_n16007 = new_n16006 ^ new_n15994;
  assign new_n16008 = new_n16007 ^ new_n16004;
  assign new_n16009 = new_n15990 ^ new_n15940;
  assign new_n16010 = ~new_n16009 & new_n15977;
  assign new_n16011 = new_n16010 ^ new_n15981;
  assign new_n16012 = new_n16011 ^ new_n15968;
  assign new_n16013 = new_n16012 ^ new_n16008;
  assign new_n16014 = new_n15973 ^ new_n15945;
  assign new_n16015 = new_n15979 ^ new_n15944;
  assign new_n16016 = ~new_n16014 & ~new_n16015;
  assign new_n16017 = new_n16016 ^ new_n15954;
  assign new_n16018 = new_n16010 ^ new_n15985;
  assign new_n16019 = new_n16018 ^ new_n16017;
  assign new_n16020 = ~new_n16013 & ~new_n16019;
  assign new_n16021 = new_n16016 ^ new_n15975;
  assign new_n16022 = new_n16021 ^ new_n15973;
  assign new_n16023 = new_n16022 ^ new_n16012;
  assign new_n16024 = new_n16023 ^ new_n16020;
  assign new_n16025 = ~new_n15946 & new_n16024;
  assign new_n16026 = new_n15953 ^ new_n15934;
  assign new_n16027 = new_n15999 ^ new_n15955;
  assign new_n16028 = new_n15973 ^ new_n15934;
  assign new_n16029 = new_n16005 ^ new_n15999;
  assign new_n16030 = new_n16029 ^ new_n16018;
  assign new_n16031 = new_n16030 ^ new_n16028;
  assign new_n16032 = new_n16023 ^ new_n16004;
  assign new_n16033 = ~new_n16031 & new_n16032;
  assign new_n16034 = new_n16033 ^ new_n16007;
  assign new_n16035 = new_n16034 ^ new_n16012;
  assign new_n16036 = new_n16020 ^ new_n16004;
  assign new_n16037 = ~new_n16036 & new_n16023;
  assign new_n16038 = new_n16037 ^ new_n16004;
  assign new_n16039 = ~new_n16035 & new_n16038;
  assign new_n16040 = new_n16037 ^ new_n16023;
  assign new_n16041 = new_n16040 ^ new_n16039;
  assign new_n16042 = new_n16041 ^ new_n16027;
  assign new_n16043 = new_n16042 ^ new_n16026;
  assign new_n16044 = new_n16043 ^ new_n15929;
  assign new_n16045 = new_n16033 ^ new_n15975;
  assign new_n16046 = new_n16045 ^ new_n15994;
  assign new_n16047 = new_n16046 ^ new_n16044;
  assign new_n16048 = ~new_n15984 & ~new_n16047;
  assign new_n16049 = new_n16039 ^ new_n16033;
  assign new_n16050 = new_n16049 ^ new_n16003;
  assign new_n16051 = new_n15968 & new_n16050;
  assign new_n16052 = new_n16039 ^ new_n16031;
  assign new_n16053 = ~new_n15945 & ~new_n16052;
  assign new_n16054 = new_n16033 ^ new_n16020;
  assign new_n16055 = new_n16022 ^ new_n16007;
  assign new_n16056 = new_n16055 ^ new_n16054;
  assign new_n16057 = ~new_n16056 & new_n15980;
  assign new_n16058 = ~new_n16047 & new_n15982;
  assign new_n16059 = new_n16058 ^ new_n16057;
  assign new_n16060 = new_n16040 ^ new_n16020;
  assign new_n16061 = new_n16060 ^ new_n16019;
  assign new_n16062 = ~new_n16061 & new_n15998;
  assign new_n16063 = new_n16062 ^ new_n16059;
  assign new_n16064 = new_n16063 ^ new_n16053;
  assign new_n16065 = new_n16064 ^ new_n16051;
  assign new_n16066 = new_n16065 ^ new_n16048;
  assign new_n16067 = new_n16066 ^ new_n16025;
  assign new_n16068 = new_n16020 ^ new_n15973;
  assign new_n16069 = new_n16016 ^ new_n16005;
  assign new_n16070 = new_n16069 ^ new_n16043;
  assign new_n16071 = new_n16070 ^ new_n16068;
  assign new_n16072 = ~new_n16009 & new_n16071;
  assign new_n16073 = ~new_n16014 & ~new_n16035;
  assign new_n16074 = new_n16073 ^ new_n16072;
  assign new_n16075 = ~new_n15974 & new_n16050;
  assign new_n16076 = ~new_n15944 & new_n16024;
  assign new_n16077 = new_n16040 ^ new_n15989;
  assign new_n16078 = ~new_n15990 & ~new_n16077;
  assign new_n16079 = new_n16078 ^ new_n16076;
  assign new_n16080 = new_n16079 ^ new_n16075;
  assign new_n16081 = new_n16080 ^ new_n16074;
  assign new_n16082 = new_n16081 ^ new_n16067;
  assign new_n16083 = new_n16082 ^ new_n15922;
  assign new_n16084 = new_n16083 ^ new_n15734;
  assign new_n16085 = new_n15368 & new_n15749;
  assign new_n16086 = ~new_n15384 & new_n15455;
  assign new_n16087 = new_n16086 ^ new_n16085;
  assign new_n16088 = new_n16087 ^ new_n15744;
  assign new_n16089 = new_n15585 ^ new_n15548;
  assign new_n16090 = ~new_n15514 & ~new_n16089;
  assign new_n16091 = ~new_n15610 & new_n15530;
  assign new_n16092 = new_n16091 ^ new_n16090;
  assign new_n16093 = new_n15585 ^ new_n15565;
  assign new_n16094 = new_n16093 ^ new_n15564;
  assign new_n16095 = ~new_n16094 & new_n15527;
  assign new_n16096 = new_n16095 ^ new_n15612;
  assign new_n16097 = new_n16096 ^ new_n15597;
  assign new_n16098 = new_n15541 & new_n15593;
  assign new_n16099 = new_n16098 ^ new_n16097;
  assign new_n16100 = new_n16099 ^ new_n15602;
  assign new_n16101 = new_n16100 ^ new_n16092;
  assign new_n16102 = new_n16101 ^ new_n16088;
  assign new_n16103 = new_n16102 ^ new_n15460;
  assign new_n16104 = new_n15752 ^ new_n15742;
  assign new_n16105 = new_n16104 ^ new_n15458;
  assign new_n16106 = new_n15576 ^ new_n15565;
  assign new_n16107 = ~new_n15522 & new_n16106;
  assign new_n16108 = ~new_n15504 & ~new_n16089;
  assign new_n16109 = new_n16108 ^ new_n16107;
  assign new_n16110 = new_n16109 ^ new_n15594;
  assign new_n16111 = new_n16110 ^ new_n16098;
  assign new_n16112 = new_n16111 ^ new_n15613;
  assign new_n16113 = new_n16112 ^ new_n16105;
  assign new_n16114 = new_n16113 ^ new_n16103;
  assign new_n16115 = new_n15918 ^ new_n15912;
  assign new_n16116 = new_n15892 ^ new_n15887;
  assign new_n16117 = ~new_n15891 & new_n15822;
  assign new_n16118 = ~new_n15853 & ~new_n15874;
  assign new_n16119 = new_n16118 ^ new_n16117;
  assign new_n16120 = new_n16119 ^ new_n15898;
  assign new_n16121 = new_n16120 ^ new_n16116;
  assign new_n16122 = new_n16121 ^ new_n16115;
  assign new_n16123 = new_n15725 ^ new_n15722;
  assign new_n16124 = new_n15715 ^ new_n15689;
  assign new_n16125 = ~new_n15688 & new_n15648;
  assign new_n16126 = new_n15666 & new_n15683;
  assign new_n16127 = new_n16126 ^ new_n16125;
  assign new_n16128 = new_n16127 ^ new_n15708;
  assign new_n16129 = new_n16128 ^ new_n16124;
  assign new_n16130 = new_n16129 ^ new_n16123;
  assign new_n16131 = new_n16130 ^ new_n393;
  assign new_n16132 = new_n16131 ^ new_n16122;
  assign new_n16133 = new_n16075 ^ new_n16072;
  assign new_n16134 = new_n16053 ^ new_n16048;
  assign new_n16135 = ~new_n16052 & new_n15997;
  assign new_n16136 = ~new_n16015 & ~new_n16035;
  assign new_n16137 = new_n16136 ^ new_n16135;
  assign new_n16138 = new_n16137 ^ new_n16059;
  assign new_n16139 = new_n16138 ^ new_n16134;
  assign new_n16140 = new_n16139 ^ new_n16133;
  assign new_n16141 = new_n16140 ^ new_n16132;
  assign new_n16142 = new_n16141 ^ new_n16114;
  assign new_n16143 = ~new_n15643 & ~new_n15727;
  assign new_n16144 = new_n16143 ^ new_n16126;
  assign new_n16145 = ~new_n15647 & new_n15692;
  assign new_n16146 = new_n16145 ^ new_n15726;
  assign new_n16147 = new_n16146 ^ new_n15710;
  assign new_n16148 = new_n16147 ^ new_n16144;
  assign new_n16149 = new_n16148 ^ new_n403;
  assign new_n16150 = new_n16149 ^ new_n16102;
  assign new_n16151 = ~new_n15550 & new_n16106;
  assign new_n16152 = new_n16151 ^ new_n16100;
  assign new_n16153 = ~new_n15561 & ~new_n15580;
  assign new_n16154 = new_n16153 ^ new_n15591;
  assign new_n16155 = new_n16154 ^ new_n16110;
  assign new_n16156 = new_n16155 ^ new_n16152;
  assign new_n16157 = new_n16156 ^ new_n15754;
  assign new_n16158 = new_n16157 ^ new_n16150;
  assign new_n16159 = new_n16085 ^ new_n15450;
  assign new_n16160 = ~new_n15391 & ~new_n15738;
  assign new_n16161 = new_n16160 ^ new_n15748;
  assign new_n16162 = new_n16161 ^ new_n15741;
  assign new_n16163 = new_n16162 ^ new_n16159;
  assign new_n16164 = ~new_n15992 & ~new_n16077;
  assign new_n16165 = new_n16164 ^ new_n16136;
  assign new_n16166 = ~new_n16061 & new_n15996;
  assign new_n16167 = new_n16166 ^ new_n16076;
  assign new_n16168 = new_n16167 ^ new_n16064;
  assign new_n16169 = new_n16168 ^ new_n16165;
  assign new_n16170 = ~new_n15814 & ~new_n15914;
  assign new_n16171 = new_n16170 ^ new_n16118;
  assign new_n16172 = ~new_n15900 & new_n15821;
  assign new_n16173 = new_n16172 ^ new_n15916;
  assign new_n16174 = new_n16173 ^ new_n15903;
  assign new_n16175 = new_n16174 ^ new_n16171;
  assign new_n16176 = new_n16175 ^ new_n16169;
  assign new_n16177 = new_n16176 ^ new_n16163;
  assign new_n16178 = new_n16177 ^ new_n16158;
  assign new_n16179 = new_n16178 ^ new_n16142;
  assign new_n16180 = new_n16179 ^ new_n16084;
  assign new_n16181 = ~new_n16056 & new_n15979;
  assign new_n16182 = new_n16181 ^ new_n16048;
  assign new_n16183 = new_n16166 ^ new_n16078;
  assign new_n16184 = new_n16183 ^ new_n16164;
  assign new_n16185 = new_n16184 ^ new_n16063;
  assign new_n16186 = new_n16185 ^ new_n16182;
  assign new_n16187 = ~new_n15896 & new_n15819;
  assign new_n16188 = new_n16187 ^ new_n15887;
  assign new_n16189 = new_n16172 ^ new_n15915;
  assign new_n16190 = new_n16189 ^ new_n16170;
  assign new_n16191 = new_n16190 ^ new_n15902;
  assign new_n16192 = new_n16191 ^ new_n16188;
  assign new_n16193 = new_n16192 ^ new_n16186;
  assign new_n16194 = new_n16091 ^ new_n15611;
  assign new_n16195 = new_n15526 & new_n15590;
  assign new_n16196 = new_n16195 ^ new_n16155;
  assign new_n16197 = new_n16196 ^ new_n16194;
  assign new_n16198 = new_n16197 ^ new_n16193;
  assign new_n16199 = new_n16086 ^ new_n15447;
  assign new_n16200 = new_n16160 ^ new_n15750;
  assign new_n16201 = new_n16200 ^ new_n16085;
  assign new_n16202 = new_n16201 ^ new_n15740;
  assign new_n16203 = new_n16202 ^ new_n16199;
  assign new_n16204 = ~new_n15635 & ~new_n15706;
  assign new_n16205 = new_n16204 ^ new_n15715;
  assign new_n16206 = new_n16145 ^ new_n15728;
  assign new_n16207 = new_n16206 ^ new_n16143;
  assign new_n16208 = new_n16207 ^ new_n15709;
  assign new_n16209 = new_n16208 ^ new_n16205;
  assign new_n16210 = new_n16209 ^ new_n433;
  assign new_n16211 = new_n16210 ^ new_n16203;
  assign new_n16212 = new_n16086 ^ new_n15456;
  assign new_n16213 = ~new_n15435 & new_n15367;
  assign new_n16214 = new_n16213 ^ new_n15753;
  assign new_n16215 = new_n16214 ^ new_n16212;
  assign new_n16216 = new_n16215 ^ new_n16211;
  assign new_n16217 = new_n16216 ^ new_n16198;
  assign new_n16218 = new_n16217 ^ new_n16180;
  assign new_n16219 = new_n16091 ^ new_n15602;
  assign new_n16220 = ~new_n16094 & new_n15523;
  assign new_n16221 = new_n16220 ^ new_n16108;
  assign new_n16222 = new_n16221 ^ new_n16090;
  assign new_n16223 = new_n16222 ^ new_n16096;
  assign new_n16224 = new_n16223 ^ new_n16219;
  assign new_n16225 = new_n16187 ^ new_n16170;
  assign new_n16226 = new_n16225 ^ new_n15905;
  assign new_n16227 = new_n16181 ^ new_n16164;
  assign new_n16228 = new_n16227 ^ new_n16066;
  assign new_n16229 = new_n16228 ^ new_n16226;
  assign new_n16230 = new_n16229 ^ new_n16224;
  assign new_n16231 = new_n16204 ^ new_n16143;
  assign new_n16232 = new_n16231 ^ new_n15716;
  assign new_n16233 = new_n16232 ^ new_n365;
  assign new_n16234 = new_n16233 ^ new_n16088;
  assign new_n16235 = new_n16234 ^ new_n16203;
  assign new_n16236 = new_n16235 ^ new_n16230;
  assign new_n16237 = new_n16181 ^ new_n16057;
  assign new_n16238 = new_n15977 & new_n16071;
  assign new_n16239 = new_n16238 ^ new_n16081;
  assign new_n16240 = new_n16239 ^ new_n16237;
  assign new_n16241 = new_n16187 ^ new_n15897;
  assign new_n16242 = new_n15823 & new_n15911;
  assign new_n16243 = new_n16242 ^ new_n15920;
  assign new_n16244 = new_n16243 ^ new_n16241;
  assign new_n16245 = new_n16244 ^ new_n16240;
  assign new_n16246 = new_n16245 ^ new_n16215;
  assign new_n16247 = new_n16222 ^ new_n16099;
  assign new_n16248 = new_n16201 ^ new_n15743;
  assign new_n16249 = new_n16248 ^ new_n16247;
  assign new_n16250 = new_n16204 ^ new_n15707;
  assign new_n16251 = ~new_n15721 & new_n15628;
  assign new_n16252 = new_n16251 ^ new_n15731;
  assign new_n16253 = new_n16252 ^ new_n16250;
  assign new_n16254 = new_n16253 ^ new_n444;
  assign new_n16255 = new_n16254 ^ new_n16249;
  assign new_n16256 = new_n16255 ^ new_n16246;
  assign new_n16257 = new_n16256 ^ new_n16236;
  assign new_n16258 = new_n16184 ^ new_n16065;
  assign new_n16259 = new_n16190 ^ new_n15904;
  assign new_n16260 = new_n16259 ^ new_n16258;
  assign new_n16261 = new_n16260 ^ new_n16102;
  assign new_n16262 = new_n16207 ^ new_n15714;
  assign new_n16263 = new_n16262 ^ new_n374;
  assign new_n16264 = new_n16263 ^ new_n16248;
  assign new_n16265 = new_n16090 ^ new_n15605;
  assign new_n16266 = new_n16220 ^ new_n16107;
  assign new_n16267 = new_n16266 ^ new_n16097;
  assign new_n16268 = new_n16267 ^ new_n16265;
  assign new_n16269 = new_n16268 ^ new_n16163;
  assign new_n16270 = new_n16269 ^ new_n16264;
  assign new_n16271 = new_n16270 ^ new_n16261;
  assign new_n16272 = new_n16271 ^ new_n16236;
  assign new_n16273 = new_n16272 ^ new_n16179;
  assign new_n16274 = new_n16105 ^ new_n16102;
  assign new_n16275 = new_n15919 ^ new_n15890;
  assign new_n16276 = new_n16275 ^ new_n16120;
  assign new_n16277 = new_n15730 ^ new_n15713;
  assign new_n16278 = new_n16277 ^ new_n16128;
  assign new_n16279 = new_n16278 ^ new_n413;
  assign new_n16280 = new_n16279 ^ new_n16276;
  assign new_n16281 = new_n16080 ^ new_n16051;
  assign new_n16282 = new_n16281 ^ new_n16138;
  assign new_n16283 = new_n16282 ^ new_n16280;
  assign new_n16284 = new_n16283 ^ new_n16274;
  assign new_n16285 = new_n16284 ^ new_n16273;
  assign new_n16286 = new_n16256 ^ new_n16217;
  assign new_n16287 = new_n16286 ^ new_n16284;
  assign new_n16288 = new_n16287 ^ new_n16142;
  assign new_n16289 = new_n16236 ^ new_n16084;
  assign new_n16290 = new_n16289 ^ new_n16288;
  assign new_n16291 = new_n16285 & new_n16290;
  assign new_n16292 = new_n16287 ^ new_n16271;
  assign new_n16293 = ~new_n16284 & ~new_n16292;
  assign new_n16294 = new_n16293 ^ new_n16291;
  assign new_n16295 = new_n16286 ^ new_n16273;
  assign new_n16296 = ~new_n16295 & new_n16289;
  assign new_n16297 = new_n16271 ^ new_n16256;
  assign new_n16298 = new_n16297 ^ new_n16289;
  assign new_n16299 = new_n16271 ^ new_n16084;
  assign new_n16300 = ~new_n16298 & new_n16299;
  assign new_n16301 = new_n16300 ^ new_n16296;
  assign new_n16302 = new_n16301 ^ new_n16294;
  assign new_n16303 = new_n16302 ^ new_n16257;
  assign new_n16304 = new_n16287 ^ new_n16236;
  assign new_n16305 = new_n16284 ^ new_n16218;
  assign new_n16306 = ~new_n16304 & ~new_n16305;
  assign new_n16307 = new_n16256 ^ new_n16180;
  assign new_n16308 = new_n16236 ^ new_n16142;
  assign new_n16309 = ~new_n16308 & new_n16307;
  assign new_n16310 = new_n16309 ^ new_n16306;
  assign new_n16311 = new_n16310 ^ new_n16236;
  assign new_n16312 = new_n16218 & new_n16272;
  assign new_n16313 = new_n16312 ^ new_n16296;
  assign new_n16314 = new_n16313 ^ new_n16307;
  assign new_n16315 = new_n16314 ^ new_n16311;
  assign new_n16316 = new_n16142 & new_n16287;
  assign new_n16317 = new_n16316 ^ new_n16142;
  assign new_n16318 = new_n16317 ^ new_n16309;
  assign new_n16319 = new_n16318 ^ new_n16289;
  assign new_n16320 = new_n16312 ^ new_n16300;
  assign new_n16321 = new_n16256 ^ new_n16178;
  assign new_n16322 = new_n16321 ^ new_n16320;
  assign new_n16323 = new_n16322 ^ new_n16319;
  assign new_n16324 = new_n16271 ^ new_n16142;
  assign new_n16325 = new_n16324 ^ new_n16289;
  assign new_n16326 = ~new_n16273 & ~new_n16325;
  assign new_n16327 = new_n16326 ^ new_n16217;
  assign new_n16328 = new_n16327 ^ new_n16273;
  assign new_n16329 = new_n16312 ^ new_n16291;
  assign new_n16330 = new_n16300 ^ new_n16084;
  assign new_n16331 = new_n16330 ^ new_n16329;
  assign new_n16332 = new_n16331 ^ new_n16328;
  assign new_n16333 = ~new_n16323 & new_n16332;
  assign new_n16334 = new_n16333 ^ new_n16315;
  assign new_n16335 = ~new_n16303 & new_n16334;
  assign new_n16336 = new_n16293 ^ new_n16271;
  assign new_n16337 = new_n16336 ^ new_n16327;
  assign new_n16338 = new_n16337 ^ new_n16333;
  assign new_n16339 = new_n16338 ^ new_n16314;
  assign new_n16340 = new_n16316 ^ new_n16306;
  assign new_n16341 = new_n16340 ^ new_n16301;
  assign new_n16342 = ~new_n16339 & ~new_n16341;
  assign new_n16343 = new_n16342 ^ new_n16335;
  assign new_n16344 = new_n16337 ^ new_n16311;
  assign new_n16345 = new_n16344 ^ new_n16343;
  assign new_n16346 = ~new_n16345 & new_n16218;
  assign new_n16347 = new_n16342 ^ new_n16333;
  assign new_n16348 = ~new_n16347 & new_n16315;
  assign new_n16349 = new_n16348 ^ new_n16315;
  assign new_n16350 = new_n16349 ^ new_n16323;
  assign new_n16351 = ~new_n16325 & ~new_n16350;
  assign new_n16352 = new_n16351 ^ new_n16346;
  assign new_n16353 = new_n16349 ^ new_n16342;
  assign new_n16354 = new_n16353 ^ new_n16341;
  assign new_n16355 = ~new_n16354 & new_n16290;
  assign new_n16356 = new_n16256 ^ new_n16142;
  assign new_n16357 = new_n16317 ^ new_n16291;
  assign new_n16358 = new_n16337 ^ new_n16335;
  assign new_n16359 = new_n16358 ^ new_n16314;
  assign new_n16360 = new_n16348 ^ new_n16333;
  assign new_n16361 = ~new_n16359 & new_n16360;
  assign new_n16362 = new_n16361 ^ new_n16349;
  assign new_n16363 = new_n16362 ^ new_n16357;
  assign new_n16364 = new_n16363 ^ new_n16356;
  assign new_n16365 = new_n16364 ^ new_n16271;
  assign new_n16366 = new_n16335 ^ new_n16309;
  assign new_n16367 = new_n16366 ^ new_n16327;
  assign new_n16368 = new_n16367 ^ new_n16365;
  assign new_n16369 = ~new_n16368 & new_n16299;
  assign new_n16370 = ~new_n16345 & new_n16272;
  assign new_n16371 = new_n16370 ^ new_n16369;
  assign new_n16372 = new_n16371 ^ new_n16355;
  assign new_n16373 = new_n16361 ^ new_n16303;
  assign new_n16374 = ~new_n16287 & ~new_n16373;
  assign new_n16375 = new_n16374 ^ new_n16372;
  assign new_n16376 = new_n16361 ^ new_n16335;
  assign new_n16377 = new_n16376 ^ new_n16332;
  assign new_n16378 = new_n16307 & new_n16377;
  assign new_n16379 = new_n16378 ^ new_n16375;
  assign new_n16380 = ~new_n16298 & ~new_n16368;
  assign new_n16381 = new_n16380 ^ new_n16379;
  assign new_n16382 = new_n16381 ^ new_n16352;
  assign new_n16383 = new_n16382 ^ new_n15309;
  assign new_n16384 = new_n14530 ^ new_n13669;
  assign new_n16385 = new_n12518 ^ new_n12482;
  assign new_n16386 = new_n16385 ^ new_n12547;
  assign new_n16387 = new_n16386 ^ new_n12249;
  assign new_n16388 = ~new_n12547 & ~new_n16387;
  assign new_n16389 = new_n16388 ^ new_n12249;
  assign new_n16390 = new_n12645 ^ new_n12249;
  assign new_n16391 = new_n12627 ^ new_n12566;
  assign new_n16392 = new_n16391 ^ new_n16390;
  assign new_n16393 = new_n12566 ^ new_n12249;
  assign new_n16394 = new_n12645 ^ new_n12595;
  assign new_n16395 = new_n16394 ^ new_n16393;
  assign new_n16396 = ~new_n16392 & ~new_n16395;
  assign new_n16397 = new_n16396 ^ new_n12518;
  assign new_n16398 = new_n16397 ^ new_n16389;
  assign new_n16399 = new_n16397 ^ new_n16392;
  assign new_n16400 = new_n16391 ^ new_n12595;
  assign new_n16401 = new_n16400 ^ new_n12518;
  assign new_n16402 = new_n16390 & new_n16401;
  assign new_n16403 = new_n12482 ^ new_n12249;
  assign new_n16404 = new_n16403 ^ new_n16394;
  assign new_n16405 = new_n12595 ^ new_n12249;
  assign new_n16406 = ~new_n16404 & new_n16405;
  assign new_n16407 = new_n16406 ^ new_n16402;
  assign new_n16408 = new_n16392 ^ new_n12547;
  assign new_n16409 = new_n16386 ^ new_n12566;
  assign new_n16410 = new_n16409 ^ new_n16394;
  assign new_n16411 = new_n16408 & new_n16410;
  assign new_n16412 = new_n16411 ^ new_n12595;
  assign new_n16413 = new_n16412 ^ new_n16407;
  assign new_n16414 = new_n16413 ^ new_n16399;
  assign new_n16415 = new_n12566 & new_n16386;
  assign new_n16416 = new_n16415 ^ new_n12566;
  assign new_n16417 = new_n12645 ^ new_n12566;
  assign new_n16418 = new_n16400 ^ new_n12482;
  assign new_n16419 = ~new_n16417 & new_n16418;
  assign new_n16420 = new_n16419 ^ new_n16416;
  assign new_n16421 = new_n16420 ^ new_n16394;
  assign new_n16422 = new_n12627 ^ new_n12482;
  assign new_n16423 = new_n16422 ^ new_n16407;
  assign new_n16424 = new_n16423 ^ new_n16421;
  assign new_n16425 = ~new_n16424 & new_n16414;
  assign new_n16426 = new_n16425 ^ new_n16398;
  assign new_n16427 = new_n16392 ^ new_n16385;
  assign new_n16428 = ~new_n16427 & new_n16394;
  assign new_n16429 = new_n16428 ^ new_n16402;
  assign new_n16430 = new_n16429 ^ new_n16418;
  assign new_n16431 = new_n16430 ^ new_n16426;
  assign new_n16432 = new_n16386 ^ new_n12645;
  assign new_n16433 = new_n16401 ^ new_n12547;
  assign new_n16434 = ~new_n16432 & ~new_n16433;
  assign new_n16435 = new_n16434 ^ new_n16415;
  assign new_n16436 = new_n16428 ^ new_n16406;
  assign new_n16437 = new_n16436 ^ new_n16435;
  assign new_n16438 = ~new_n16431 & ~new_n16437;
  assign new_n16439 = new_n16434 ^ new_n16419;
  assign new_n16440 = new_n16439 ^ new_n12645;
  assign new_n16441 = new_n16440 ^ new_n16430;
  assign new_n16442 = new_n16441 ^ new_n16438;
  assign new_n16443 = ~new_n16387 & new_n16442;
  assign new_n16444 = new_n12645 ^ new_n12482;
  assign new_n16445 = new_n16411 ^ new_n16388;
  assign new_n16446 = new_n16445 ^ new_n16436;
  assign new_n16447 = new_n16446 ^ new_n16444;
  assign new_n16448 = new_n16441 ^ new_n16425;
  assign new_n16449 = ~new_n16447 & new_n16448;
  assign new_n16450 = new_n16449 ^ new_n16398;
  assign new_n16451 = new_n16450 ^ new_n16430;
  assign new_n16452 = new_n16438 ^ new_n16425;
  assign new_n16453 = new_n16441 & new_n16452;
  assign new_n16454 = new_n16453 ^ new_n16448;
  assign new_n16455 = ~new_n16451 & new_n16454;
  assign new_n16456 = new_n16455 ^ new_n16449;
  assign new_n16457 = new_n16456 ^ new_n16414;
  assign new_n16458 = new_n16418 & new_n16457;
  assign new_n16459 = new_n16455 ^ new_n16447;
  assign new_n16460 = ~new_n16386 & ~new_n16459;
  assign new_n16461 = new_n16453 ^ new_n16438;
  assign new_n16462 = new_n16461 ^ new_n16437;
  assign new_n16463 = ~new_n16462 & new_n16410;
  assign new_n16464 = new_n16449 ^ new_n16438;
  assign new_n16465 = new_n16440 ^ new_n16398;
  assign new_n16466 = new_n16465 ^ new_n16464;
  assign new_n16467 = ~new_n16466 & new_n16390;
  assign new_n16468 = new_n12566 ^ new_n12482;
  assign new_n16469 = new_n16416 ^ new_n16411;
  assign new_n16470 = new_n16455 ^ new_n16453;
  assign new_n16471 = new_n16470 ^ new_n16469;
  assign new_n16472 = new_n16471 ^ new_n16468;
  assign new_n16473 = new_n16472 ^ new_n12249;
  assign new_n16474 = new_n16449 ^ new_n16419;
  assign new_n16475 = new_n16474 ^ new_n16397;
  assign new_n16476 = new_n16475 ^ new_n16473;
  assign new_n16477 = ~new_n16476 & new_n16405;
  assign new_n16478 = new_n16477 ^ new_n16467;
  assign new_n16479 = new_n16478 ^ new_n16463;
  assign new_n16480 = new_n16479 ^ new_n16460;
  assign new_n16481 = new_n16480 ^ new_n16458;
  assign new_n16482 = ~new_n16404 & ~new_n16476;
  assign new_n16483 = new_n16482 ^ new_n16481;
  assign new_n16484 = new_n16483 ^ new_n16443;
  assign new_n16485 = ~new_n16432 & ~new_n16451;
  assign new_n16486 = new_n16438 ^ new_n12645;
  assign new_n16487 = new_n16434 ^ new_n16388;
  assign new_n16488 = new_n16487 ^ new_n16472;
  assign new_n16489 = new_n16488 ^ new_n16486;
  assign new_n16490 = ~new_n16427 & new_n16489;
  assign new_n16491 = new_n16490 ^ new_n16485;
  assign new_n16492 = new_n16453 ^ new_n16424;
  assign new_n16493 = ~new_n16392 & ~new_n16492;
  assign new_n16494 = ~new_n12547 & new_n16442;
  assign new_n16495 = new_n16494 ^ new_n16493;
  assign new_n16496 = ~new_n16417 & new_n16457;
  assign new_n16497 = new_n16496 ^ new_n16495;
  assign new_n16498 = new_n16497 ^ new_n16491;
  assign new_n16499 = new_n16498 ^ new_n16484;
  assign new_n16500 = new_n16499 ^ new_n16384;
  assign new_n16501 = new_n15763 ^ new_n11514;
  assign new_n16502 = new_n12248 ^ new_n7593;
  assign new_n16503 = new_n16502 ^ new_n11330;
  assign new_n16504 = new_n16503 ^ new_n11552;
  assign new_n16505 = new_n16504 ^ new_n16501;
  assign new_n16506 = new_n12644 ^ new_n6843;
  assign new_n16507 = new_n16506 ^ new_n11456;
  assign new_n16508 = new_n15756 ^ new_n11370;
  assign new_n16509 = new_n16508 ^ new_n16507;
  assign new_n16510 = new_n16509 ^ new_n16505;
  assign new_n16511 = new_n15809 ^ new_n11449;
  assign new_n16512 = new_n12565 ^ new_n7464;
  assign new_n16513 = new_n16512 ^ new_n11541;
  assign new_n16514 = new_n16513 ^ new_n11552;
  assign new_n16515 = new_n16514 ^ new_n16511;
  assign new_n16516 = new_n12626 ^ new_n7622;
  assign new_n16517 = new_n16516 ^ new_n11486;
  assign new_n16518 = new_n16517 ^ new_n11552;
  assign new_n16519 = new_n15758 ^ new_n11572;
  assign new_n16520 = new_n16519 ^ new_n16518;
  assign new_n16521 = new_n16520 ^ new_n16515;
  assign new_n16522 = new_n16521 ^ new_n16510;
  assign new_n16523 = new_n16515 ^ new_n16505;
  assign new_n16524 = new_n12594 ^ new_n1012;
  assign new_n16525 = new_n16524 ^ new_n11494;
  assign new_n16526 = new_n15794 ^ new_n11531;
  assign new_n16527 = new_n16526 ^ new_n16525;
  assign new_n16528 = new_n16527 ^ new_n16509;
  assign new_n16529 = new_n16528 ^ new_n16523;
  assign new_n16530 = ~new_n16522 & ~new_n16529;
  assign new_n16531 = new_n12517 ^ new_n7540;
  assign new_n16532 = new_n16531 ^ new_n11412;
  assign new_n16533 = new_n15784 ^ new_n9162;
  assign new_n16534 = new_n16533 ^ new_n16532;
  assign new_n16535 = new_n16534 ^ new_n16530;
  assign new_n16536 = new_n12546 ^ new_n7648;
  assign new_n16537 = new_n16536 ^ new_n11431;
  assign new_n16538 = new_n15798 ^ new_n11552;
  assign new_n16539 = new_n16538 ^ new_n16537;
  assign new_n16540 = new_n12481 ^ new_n7574;
  assign new_n16541 = new_n16540 ^ new_n10181;
  assign new_n16542 = new_n15769 ^ new_n11474;
  assign new_n16543 = new_n16542 ^ new_n16541;
  assign new_n16544 = new_n16543 ^ new_n16534;
  assign new_n16545 = ~new_n16539 & ~new_n16544;
  assign new_n16546 = new_n16505 & new_n16539;
  assign new_n16547 = new_n16546 ^ new_n16545;
  assign new_n16548 = new_n16547 ^ new_n16535;
  assign new_n16549 = new_n16544 ^ new_n16539;
  assign new_n16550 = new_n16515 & new_n16549;
  assign new_n16551 = new_n16550 ^ new_n16515;
  assign new_n16552 = new_n16515 ^ new_n16509;
  assign new_n16553 = new_n16527 ^ new_n16521;
  assign new_n16554 = new_n16553 ^ new_n16543;
  assign new_n16555 = ~new_n16552 & new_n16554;
  assign new_n16556 = new_n16555 ^ new_n16551;
  assign new_n16557 = new_n16556 ^ new_n16528;
  assign new_n16558 = new_n16543 ^ new_n16505;
  assign new_n16559 = new_n16558 ^ new_n16528;
  assign new_n16560 = new_n16527 ^ new_n16505;
  assign new_n16561 = ~new_n16559 & new_n16560;
  assign new_n16562 = new_n16553 ^ new_n16534;
  assign new_n16563 = new_n16510 & new_n16562;
  assign new_n16564 = new_n16563 ^ new_n16561;
  assign new_n16565 = new_n16543 ^ new_n16520;
  assign new_n16566 = new_n16565 ^ new_n16564;
  assign new_n16567 = new_n16566 ^ new_n16557;
  assign new_n16568 = new_n16535 ^ new_n16522;
  assign new_n16569 = new_n16549 ^ new_n16515;
  assign new_n16570 = new_n16569 ^ new_n16528;
  assign new_n16571 = new_n16539 ^ new_n16522;
  assign new_n16572 = new_n16570 & new_n16571;
  assign new_n16573 = new_n16572 ^ new_n16563;
  assign new_n16574 = new_n16561 ^ new_n16527;
  assign new_n16575 = new_n16574 ^ new_n16573;
  assign new_n16576 = new_n16575 ^ new_n16568;
  assign new_n16577 = ~new_n16567 & new_n16576;
  assign new_n16578 = new_n16577 ^ new_n16548;
  assign new_n16579 = new_n16544 ^ new_n16522;
  assign new_n16580 = ~new_n16579 & new_n16528;
  assign new_n16581 = new_n16580 ^ new_n16563;
  assign new_n16582 = new_n16581 ^ new_n16554;
  assign new_n16583 = new_n16582 ^ new_n16578;
  assign new_n16584 = new_n16549 ^ new_n16509;
  assign new_n16585 = new_n16562 ^ new_n16539;
  assign new_n16586 = ~new_n16584 & ~new_n16585;
  assign new_n16587 = new_n16586 ^ new_n16550;
  assign new_n16588 = new_n16580 ^ new_n16561;
  assign new_n16589 = new_n16588 ^ new_n16587;
  assign new_n16590 = ~new_n16583 & ~new_n16589;
  assign new_n16591 = new_n16586 ^ new_n16555;
  assign new_n16592 = new_n16591 ^ new_n16509;
  assign new_n16593 = new_n16592 ^ new_n16582;
  assign new_n16594 = new_n16593 ^ new_n16590;
  assign new_n16595 = new_n16549 ^ new_n16505;
  assign new_n16596 = ~new_n16595 & new_n16594;
  assign new_n16597 = new_n16543 ^ new_n16509;
  assign new_n16598 = new_n16547 ^ new_n16505;
  assign new_n16599 = new_n16598 ^ new_n16572;
  assign new_n16600 = new_n16599 ^ new_n16588;
  assign new_n16601 = new_n16600 ^ new_n16597;
  assign new_n16602 = new_n16593 ^ new_n16577;
  assign new_n16603 = ~new_n16601 & new_n16602;
  assign new_n16604 = new_n16603 ^ new_n16548;
  assign new_n16605 = new_n16604 ^ new_n16582;
  assign new_n16606 = new_n16590 ^ new_n16577;
  assign new_n16607 = ~new_n16606 & new_n16593;
  assign new_n16608 = new_n16607 ^ new_n16577;
  assign new_n16609 = ~new_n16605 & new_n16608;
  assign new_n16610 = new_n16609 ^ new_n16601;
  assign new_n16611 = ~new_n16549 & ~new_n16610;
  assign new_n16612 = new_n16543 ^ new_n16515;
  assign new_n16613 = new_n16572 ^ new_n16551;
  assign new_n16614 = new_n16607 ^ new_n16593;
  assign new_n16615 = new_n16614 ^ new_n16609;
  assign new_n16616 = new_n16615 ^ new_n16613;
  assign new_n16617 = new_n16616 ^ new_n16612;
  assign new_n16618 = new_n16617 ^ new_n16505;
  assign new_n16619 = new_n16603 ^ new_n16555;
  assign new_n16620 = new_n16619 ^ new_n16535;
  assign new_n16621 = new_n16620 ^ new_n16618;
  assign new_n16622 = ~new_n16621 & new_n16560;
  assign new_n16623 = new_n16603 ^ new_n16590;
  assign new_n16624 = new_n16592 ^ new_n16548;
  assign new_n16625 = new_n16624 ^ new_n16623;
  assign new_n16626 = ~new_n16625 & new_n16510;
  assign new_n16627 = new_n16626 ^ new_n16622;
  assign new_n16628 = new_n16614 ^ new_n16590;
  assign new_n16629 = new_n16628 ^ new_n16589;
  assign new_n16630 = ~new_n16629 & new_n16570;
  assign new_n16631 = new_n16630 ^ new_n16627;
  assign new_n16632 = new_n16631 ^ new_n16611;
  assign new_n16633 = new_n16609 ^ new_n16603;
  assign new_n16634 = new_n16633 ^ new_n16576;
  assign new_n16635 = new_n16554 & new_n16634;
  assign new_n16636 = new_n16635 ^ new_n16632;
  assign new_n16637 = ~new_n16559 & ~new_n16621;
  assign new_n16638 = new_n16637 ^ new_n16636;
  assign new_n16639 = new_n16638 ^ new_n16596;
  assign new_n16640 = ~new_n16552 & new_n16634;
  assign new_n16641 = ~new_n16539 & new_n16594;
  assign new_n16642 = new_n16614 ^ new_n16567;
  assign new_n16643 = ~new_n16522 & ~new_n16642;
  assign new_n16644 = new_n16643 ^ new_n16641;
  assign new_n16645 = new_n16644 ^ new_n16640;
  assign new_n16646 = new_n16590 ^ new_n16509;
  assign new_n16647 = new_n16598 ^ new_n16586;
  assign new_n16648 = new_n16647 ^ new_n16617;
  assign new_n16649 = new_n16648 ^ new_n16646;
  assign new_n16650 = ~new_n16579 & new_n16649;
  assign new_n16651 = ~new_n16584 & ~new_n16605;
  assign new_n16652 = new_n16651 ^ new_n16650;
  assign new_n16653 = new_n16652 ^ new_n16645;
  assign new_n16654 = new_n16653 ^ new_n16639;
  assign new_n16655 = new_n16654 ^ new_n16500;
  assign new_n16656 = new_n16650 ^ new_n16640;
  assign new_n16657 = new_n16637 ^ new_n16611;
  assign new_n16658 = ~new_n16610 & new_n16569;
  assign new_n16659 = ~new_n16585 & ~new_n16605;
  assign new_n16660 = new_n16659 ^ new_n16658;
  assign new_n16661 = new_n16660 ^ new_n16627;
  assign new_n16662 = new_n16661 ^ new_n16657;
  assign new_n16663 = new_n16662 ^ new_n16656;
  assign new_n16664 = new_n14869 ^ new_n14861;
  assign new_n16665 = new_n16664 ^ new_n14880;
  assign new_n16666 = new_n16665 ^ new_n14765;
  assign new_n16667 = new_n14525 ^ new_n13640;
  assign new_n16668 = new_n16667 ^ new_n14883;
  assign new_n16669 = new_n16668 ^ new_n14895;
  assign new_n16670 = new_n16669 ^ new_n16666;
  assign new_n16671 = new_n14773 ^ new_n14650;
  assign new_n16672 = new_n14556 ^ new_n13713;
  assign new_n16673 = new_n16672 ^ new_n14861;
  assign new_n16674 = new_n16673 ^ new_n14234;
  assign new_n16675 = new_n16674 ^ new_n16671;
  assign new_n16676 = new_n16675 ^ new_n16670;
  assign new_n16677 = new_n14695 ^ new_n14511;
  assign new_n16678 = new_n14541 ^ new_n13550;
  assign new_n16679 = new_n14852 ^ new_n14845;
  assign new_n16680 = new_n16679 ^ new_n16678;
  assign new_n16681 = new_n16680 ^ new_n16677;
  assign new_n16682 = new_n16681 ^ new_n16675;
  assign new_n16683 = new_n14546 ^ new_n12868;
  assign new_n16684 = new_n16683 ^ new_n14723;
  assign new_n16685 = new_n16684 ^ new_n16664;
  assign new_n16686 = new_n14852 ^ new_n14829;
  assign new_n16687 = new_n16686 ^ new_n14815;
  assign new_n16688 = new_n16687 ^ new_n16685;
  assign new_n16689 = new_n16688 ^ new_n16675;
  assign new_n16690 = new_n14519 ^ new_n13684;
  assign new_n16691 = new_n16690 ^ new_n16664;
  assign new_n16692 = new_n16691 ^ new_n14842;
  assign new_n16693 = new_n14898 ^ new_n14815;
  assign new_n16694 = new_n16693 ^ new_n14905;
  assign new_n16695 = new_n16694 ^ new_n16692;
  assign new_n16696 = new_n16695 ^ new_n16670;
  assign new_n16697 = new_n16696 ^ new_n16689;
  assign new_n16698 = new_n14536 ^ new_n13601;
  assign new_n16699 = new_n16698 ^ new_n14780;
  assign new_n16700 = new_n16664 ^ new_n14884;
  assign new_n16701 = new_n16700 ^ new_n16699;
  assign new_n16702 = new_n16701 ^ new_n16697;
  assign new_n16703 = new_n14866 ^ new_n14742;
  assign new_n16704 = new_n14513 ^ new_n13572;
  assign new_n16705 = new_n16704 ^ new_n14234;
  assign new_n16706 = new_n16705 ^ new_n14695;
  assign new_n16707 = new_n16706 ^ new_n16703;
  assign new_n16708 = new_n16707 ^ new_n16681;
  assign new_n16709 = new_n16708 ^ new_n16701;
  assign new_n16710 = new_n16709 ^ new_n16670;
  assign new_n16711 = new_n16384 ^ new_n14905;
  assign new_n16712 = new_n14802 ^ new_n14764;
  assign new_n16713 = new_n16712 ^ new_n14824;
  assign new_n16714 = new_n16713 ^ new_n16711;
  assign new_n16715 = new_n16714 ^ new_n16675;
  assign new_n16716 = new_n16715 ^ new_n16710;
  assign new_n16717 = ~new_n16702 & ~new_n16716;
  assign new_n16718 = new_n16709 ^ new_n16688;
  assign new_n16719 = new_n16701 & new_n16718;
  assign new_n16720 = new_n16719 ^ new_n16717;
  assign new_n16721 = new_n16688 ^ new_n16681;
  assign new_n16722 = new_n16721 ^ new_n16715;
  assign new_n16723 = new_n16714 ^ new_n16688;
  assign new_n16724 = ~new_n16723 & new_n16722;
  assign new_n16725 = new_n16708 ^ new_n16697;
  assign new_n16726 = ~new_n16715 & ~new_n16725;
  assign new_n16727 = new_n16726 ^ new_n16724;
  assign new_n16728 = new_n16727 ^ new_n16720;
  assign new_n16729 = new_n16728 ^ new_n16682;
  assign new_n16730 = new_n16688 ^ new_n16670;
  assign new_n16731 = new_n16730 ^ new_n16715;
  assign new_n16732 = ~new_n16697 & ~new_n16731;
  assign new_n16733 = new_n16732 ^ new_n16707;
  assign new_n16734 = new_n16733 ^ new_n16697;
  assign new_n16735 = new_n16714 ^ new_n16696;
  assign new_n16736 = new_n16735 ^ new_n16707;
  assign new_n16737 = ~new_n16736 & new_n16689;
  assign new_n16738 = new_n16737 ^ new_n16724;
  assign new_n16739 = new_n16717 ^ new_n16714;
  assign new_n16740 = new_n16739 ^ new_n16738;
  assign new_n16741 = new_n16740 ^ new_n16734;
  assign new_n16742 = ~new_n16670 & ~new_n16709;
  assign new_n16743 = new_n16742 ^ new_n16670;
  assign new_n16744 = new_n16735 ^ new_n16681;
  assign new_n16745 = ~new_n16744 & new_n16676;
  assign new_n16746 = new_n16745 ^ new_n16743;
  assign new_n16747 = new_n16746 ^ new_n16715;
  assign new_n16748 = new_n16695 ^ new_n16681;
  assign new_n16749 = new_n16748 ^ new_n16738;
  assign new_n16750 = new_n16749 ^ new_n16747;
  assign new_n16751 = ~new_n16741 & new_n16750;
  assign new_n16752 = new_n16737 ^ new_n16726;
  assign new_n16753 = new_n16752 ^ new_n16744;
  assign new_n16754 = new_n16709 ^ new_n16675;
  assign new_n16755 = new_n16736 ^ new_n16701;
  assign new_n16756 = ~new_n16755 & new_n16754;
  assign new_n16757 = new_n16756 ^ new_n16745;
  assign new_n16758 = new_n16757 ^ new_n16675;
  assign new_n16759 = new_n16758 ^ new_n16753;
  assign new_n16760 = new_n16759 ^ new_n16751;
  assign new_n16761 = ~new_n16729 & ~new_n16760;
  assign new_n16762 = new_n16719 ^ new_n16688;
  assign new_n16763 = new_n16762 ^ new_n16733;
  assign new_n16764 = new_n16763 ^ new_n16761;
  assign new_n16765 = new_n16764 ^ new_n16753;
  assign new_n16766 = new_n16763 ^ new_n16751;
  assign new_n16767 = new_n16766 ^ new_n16753;
  assign new_n16768 = new_n16756 ^ new_n16742;
  assign new_n16769 = new_n16768 ^ new_n16727;
  assign new_n16770 = ~new_n16769 & new_n16767;
  assign new_n16771 = new_n16770 ^ new_n16751;
  assign new_n16772 = ~new_n16759 & ~new_n16771;
  assign new_n16773 = new_n16772 ^ new_n16751;
  assign new_n16774 = new_n16765 & new_n16773;
  assign new_n16775 = new_n16774 ^ new_n16761;
  assign new_n16776 = new_n16775 ^ new_n16741;
  assign new_n16777 = ~new_n16776 & new_n16676;
  assign new_n16778 = new_n16770 ^ new_n16675;
  assign new_n16779 = new_n16756 ^ new_n16719;
  assign new_n16780 = new_n16681 ^ new_n16670;
  assign new_n16781 = new_n16743 ^ new_n16717;
  assign new_n16782 = new_n16772 ^ new_n16759;
  assign new_n16783 = new_n16782 ^ new_n16774;
  assign new_n16784 = new_n16783 ^ new_n16781;
  assign new_n16785 = new_n16784 ^ new_n16780;
  assign new_n16786 = new_n16785 ^ new_n16779;
  assign new_n16787 = new_n16786 ^ new_n16778;
  assign new_n16788 = ~new_n16725 & ~new_n16787;
  assign new_n16789 = new_n16788 ^ new_n16777;
  assign new_n16790 = new_n16774 ^ new_n16729;
  assign new_n16791 = ~new_n16790 & new_n16709;
  assign new_n16792 = new_n16785 ^ new_n16688;
  assign new_n16793 = new_n16761 ^ new_n16745;
  assign new_n16794 = new_n16793 ^ new_n16733;
  assign new_n16795 = new_n16794 ^ new_n16792;
  assign new_n16796 = new_n16722 & new_n16795;
  assign new_n16797 = new_n16796 ^ new_n16791;
  assign new_n16798 = ~new_n16790 & new_n16710;
  assign new_n16799 = ~new_n16755 & new_n16765;
  assign new_n16800 = new_n16799 ^ new_n16798;
  assign new_n16801 = ~new_n16723 & new_n16795;
  assign new_n16802 = new_n16770 ^ new_n16761;
  assign new_n16803 = new_n16763 ^ new_n16758;
  assign new_n16804 = new_n16803 ^ new_n16802;
  assign new_n16805 = ~new_n16804 & new_n16689;
  assign new_n16806 = new_n16805 ^ new_n16801;
  assign new_n16807 = new_n16806 ^ new_n16800;
  assign new_n16808 = new_n16807 ^ new_n16797;
  assign new_n16809 = new_n16808 ^ new_n16789;
  assign new_n16810 = new_n16809 ^ new_n16663;
  assign new_n16811 = new_n13592 ^ new_n13516;
  assign new_n16812 = new_n14097 ^ new_n8985;
  assign new_n16813 = new_n16812 ^ new_n13718;
  assign new_n16814 = new_n16813 ^ new_n13562;
  assign new_n16815 = new_n16814 ^ new_n16811;
  assign new_n16816 = new_n13531 ^ new_n13169;
  assign new_n16817 = new_n14675 ^ new_n9024;
  assign new_n16818 = new_n16817 ^ new_n13588;
  assign new_n16819 = new_n16818 ^ new_n13497;
  assign new_n16820 = new_n16819 ^ new_n16816;
  assign new_n16821 = new_n16820 ^ new_n16815;
  assign new_n16822 = new_n13710 ^ new_n13607;
  assign new_n16823 = new_n14877 ^ new_n9001;
  assign new_n16824 = new_n16823 ^ new_n13646;
  assign new_n16825 = new_n16824 ^ new_n13614;
  assign new_n16826 = new_n16825 ^ new_n16822;
  assign new_n16827 = new_n16826 ^ new_n16821;
  assign new_n16828 = new_n14848 ^ new_n9065;
  assign new_n16829 = new_n16828 ^ new_n13710;
  assign new_n16830 = new_n16829 ^ new_n13694;
  assign new_n16831 = new_n15464 ^ new_n13461;
  assign new_n16832 = new_n16831 ^ new_n16830;
  assign new_n16833 = new_n16832 ^ new_n16827;
  assign new_n16834 = new_n13710 ^ new_n13651;
  assign new_n16835 = new_n16834 ^ new_n13621;
  assign new_n16836 = new_n14791 ^ new_n8904;
  assign new_n16837 = new_n16836 ^ new_n13678;
  assign new_n16838 = new_n16837 ^ new_n13633;
  assign new_n16839 = new_n16838 ^ new_n16835;
  assign new_n16840 = new_n16827 & new_n16839;
  assign new_n16841 = new_n16840 ^ new_n16839;
  assign new_n16842 = new_n14857 ^ new_n9044;
  assign new_n16843 = new_n16842 ^ new_n13567;
  assign new_n16844 = new_n15474 ^ new_n13454;
  assign new_n16845 = new_n16844 ^ new_n16843;
  assign new_n16846 = new_n16845 ^ new_n16839;
  assign new_n16847 = new_n13673 ^ new_n13659;
  assign new_n16848 = new_n16847 ^ new_n13700;
  assign new_n16849 = new_n14079 ^ new_n8352;
  assign new_n16850 = new_n16849 ^ new_n13634;
  assign new_n16851 = new_n16850 ^ new_n16848;
  assign new_n16852 = new_n13689 ^ new_n13468;
  assign new_n16853 = new_n16852 ^ new_n13477;
  assign new_n16854 = new_n14809 ^ new_n8931;
  assign new_n16855 = new_n16854 ^ new_n13710;
  assign new_n16856 = new_n16855 ^ new_n13664;
  assign new_n16857 = new_n16856 ^ new_n16853;
  assign new_n16858 = new_n16857 ^ new_n16839;
  assign new_n16859 = new_n16858 ^ new_n16851;
  assign new_n16860 = new_n16859 ^ new_n16820;
  assign new_n16861 = ~new_n16846 & new_n16860;
  assign new_n16862 = new_n16861 ^ new_n16841;
  assign new_n16863 = new_n16851 ^ new_n16845;
  assign new_n16864 = new_n16863 ^ new_n16862;
  assign new_n16865 = new_n16851 ^ new_n16832;
  assign new_n16866 = new_n16832 ^ new_n16820;
  assign new_n16867 = new_n16866 ^ new_n16863;
  assign new_n16868 = ~new_n16867 & new_n16865;
  assign new_n16869 = new_n16845 ^ new_n16832;
  assign new_n16870 = new_n16859 ^ new_n16815;
  assign new_n16871 = new_n16869 & new_n16870;
  assign new_n16872 = new_n16871 ^ new_n16868;
  assign new_n16873 = new_n16857 ^ new_n16820;
  assign new_n16874 = new_n16873 ^ new_n16872;
  assign new_n16875 = new_n16874 ^ new_n16864;
  assign new_n16876 = new_n16869 ^ new_n16858;
  assign new_n16877 = new_n16865 ^ new_n16846;
  assign new_n16878 = ~new_n16876 & ~new_n16877;
  assign new_n16879 = new_n16878 ^ new_n16815;
  assign new_n16880 = new_n16879 ^ new_n16876;
  assign new_n16881 = new_n16876 ^ new_n16826;
  assign new_n16882 = new_n16839 ^ new_n16827;
  assign new_n16883 = new_n16882 ^ new_n16863;
  assign new_n16884 = new_n16881 & new_n16883;
  assign new_n16885 = new_n16884 ^ new_n16871;
  assign new_n16886 = new_n16868 ^ new_n16851;
  assign new_n16887 = new_n16886 ^ new_n16885;
  assign new_n16888 = new_n16887 ^ new_n16880;
  assign new_n16889 = ~new_n16875 & new_n16888;
  assign new_n16890 = ~new_n16826 & ~new_n16833;
  assign new_n16891 = new_n16890 ^ new_n16832;
  assign new_n16892 = new_n16891 ^ new_n16879;
  assign new_n16893 = new_n16892 ^ new_n16889;
  assign new_n16894 = new_n16876 ^ new_n16821;
  assign new_n16895 = ~new_n16894 & new_n16863;
  assign new_n16896 = new_n16895 ^ new_n16871;
  assign new_n16897 = new_n16896 ^ new_n16860;
  assign new_n16898 = new_n16897 ^ new_n16893;
  assign new_n16899 = new_n16845 ^ new_n16827;
  assign new_n16900 = new_n16870 ^ new_n16826;
  assign new_n16901 = ~new_n16899 & ~new_n16900;
  assign new_n16902 = new_n16901 ^ new_n16840;
  assign new_n16903 = new_n16895 ^ new_n16868;
  assign new_n16904 = new_n16903 ^ new_n16902;
  assign new_n16905 = ~new_n16898 & ~new_n16904;
  assign new_n16906 = new_n16901 ^ new_n16861;
  assign new_n16907 = new_n16906 ^ new_n16845;
  assign new_n16908 = new_n16907 ^ new_n16897;
  assign new_n16909 = new_n16908 ^ new_n16905;
  assign new_n16910 = ~new_n16833 & new_n16909;
  assign new_n16911 = new_n16839 ^ new_n16820;
  assign new_n16912 = new_n16884 ^ new_n16841;
  assign new_n16913 = new_n16845 ^ new_n16820;
  assign new_n16914 = new_n16890 ^ new_n16884;
  assign new_n16915 = new_n16914 ^ new_n16903;
  assign new_n16916 = new_n16915 ^ new_n16913;
  assign new_n16917 = new_n16908 ^ new_n16889;
  assign new_n16918 = ~new_n16916 & new_n16917;
  assign new_n16919 = new_n16918 ^ new_n16892;
  assign new_n16920 = new_n16919 ^ new_n16897;
  assign new_n16921 = new_n16905 ^ new_n16889;
  assign new_n16922 = ~new_n16921 & new_n16908;
  assign new_n16923 = new_n16922 ^ new_n16889;
  assign new_n16924 = ~new_n16920 & new_n16923;
  assign new_n16925 = new_n16922 ^ new_n16908;
  assign new_n16926 = new_n16925 ^ new_n16924;
  assign new_n16927 = new_n16926 ^ new_n16912;
  assign new_n16928 = new_n16927 ^ new_n16911;
  assign new_n16929 = new_n16928 ^ new_n16832;
  assign new_n16930 = new_n16918 ^ new_n16861;
  assign new_n16931 = new_n16930 ^ new_n16879;
  assign new_n16932 = new_n16931 ^ new_n16929;
  assign new_n16933 = ~new_n16867 & ~new_n16932;
  assign new_n16934 = new_n16924 ^ new_n16918;
  assign new_n16935 = new_n16934 ^ new_n16888;
  assign new_n16936 = new_n16860 & new_n16935;
  assign new_n16937 = new_n16924 ^ new_n16916;
  assign new_n16938 = ~new_n16827 & ~new_n16937;
  assign new_n16939 = new_n16918 ^ new_n16905;
  assign new_n16940 = new_n16907 ^ new_n16892;
  assign new_n16941 = new_n16940 ^ new_n16939;
  assign new_n16942 = ~new_n16941 & new_n16869;
  assign new_n16943 = ~new_n16932 & new_n16865;
  assign new_n16944 = new_n16943 ^ new_n16942;
  assign new_n16945 = new_n16925 ^ new_n16905;
  assign new_n16946 = new_n16945 ^ new_n16904;
  assign new_n16947 = ~new_n16946 & new_n16883;
  assign new_n16948 = new_n16947 ^ new_n16944;
  assign new_n16949 = new_n16948 ^ new_n16938;
  assign new_n16950 = new_n16949 ^ new_n16936;
  assign new_n16951 = new_n16950 ^ new_n16933;
  assign new_n16952 = new_n16951 ^ new_n16910;
  assign new_n16953 = ~new_n16826 & new_n16909;
  assign new_n16954 = new_n16925 ^ new_n16875;
  assign new_n16955 = ~new_n16876 & ~new_n16954;
  assign new_n16956 = new_n16955 ^ new_n16953;
  assign new_n16957 = ~new_n16846 & new_n16935;
  assign new_n16958 = new_n16957 ^ new_n16956;
  assign new_n16959 = ~new_n16899 & ~new_n16920;
  assign new_n16960 = new_n16905 ^ new_n16845;
  assign new_n16961 = new_n16901 ^ new_n16890;
  assign new_n16962 = new_n16961 ^ new_n16928;
  assign new_n16963 = new_n16962 ^ new_n16960;
  assign new_n16964 = ~new_n16894 & new_n16963;
  assign new_n16965 = new_n16964 ^ new_n16959;
  assign new_n16966 = new_n16965 ^ new_n16958;
  assign new_n16967 = new_n16966 ^ new_n16952;
  assign new_n16968 = new_n13835 ^ new_n12410;
  assign new_n16969 = new_n12641 ^ new_n12638;
  assign new_n16970 = new_n16969 ^ new_n12403;
  assign new_n16971 = new_n16970 ^ new_n12621;
  assign new_n16972 = new_n16971 ^ new_n16968;
  assign new_n16973 = new_n12638 ^ new_n12504;
  assign new_n16974 = new_n16973 ^ new_n12509;
  assign new_n16975 = new_n13838 ^ new_n12144;
  assign new_n16976 = new_n16975 ^ new_n16974;
  assign new_n16977 = new_n16976 ^ new_n16972;
  assign new_n16978 = new_n16969 ^ new_n13840;
  assign new_n16979 = new_n16978 ^ new_n12540;
  assign new_n16980 = new_n12601 ^ new_n12559;
  assign new_n16981 = new_n16980 ^ new_n16979;
  assign new_n16982 = new_n16969 ^ new_n13841;
  assign new_n16983 = new_n16982 ^ new_n12590;
  assign new_n16984 = new_n12616 ^ new_n12266;
  assign new_n16985 = new_n16984 ^ new_n16983;
  assign new_n16986 = new_n16985 ^ new_n16981;
  assign new_n16987 = new_n16986 ^ new_n16977;
  assign new_n16988 = new_n16981 ^ new_n16972;
  assign new_n16989 = new_n12604 ^ new_n12585;
  assign new_n16990 = new_n16989 ^ new_n12611;
  assign new_n16991 = new_n13845 ^ new_n12560;
  assign new_n16992 = new_n16991 ^ new_n16990;
  assign new_n16993 = new_n16992 ^ new_n16976;
  assign new_n16994 = new_n16993 ^ new_n16988;
  assign new_n16995 = new_n16987 & new_n16994;
  assign new_n16996 = new_n12504 ^ new_n12428;
  assign new_n16997 = new_n16996 ^ new_n12447;
  assign new_n16998 = new_n13832 ^ new_n12636;
  assign new_n16999 = new_n16998 ^ new_n16997;
  assign new_n17000 = new_n16999 ^ new_n16995;
  assign new_n17001 = new_n12573 ^ new_n12533;
  assign new_n17002 = new_n16969 ^ new_n13830;
  assign new_n17003 = new_n17002 ^ new_n17001;
  assign new_n17004 = new_n12403 ^ new_n11845;
  assign new_n17005 = new_n17004 ^ new_n12428;
  assign new_n17006 = new_n13831 ^ new_n12500;
  assign new_n17007 = new_n17006 ^ new_n17005;
  assign new_n17008 = new_n17007 ^ new_n16999;
  assign new_n17009 = ~new_n17008 & new_n17003;
  assign new_n17010 = ~new_n17003 & new_n16972;
  assign new_n17011 = new_n17010 ^ new_n17009;
  assign new_n17012 = new_n17011 ^ new_n17000;
  assign new_n17013 = new_n17000 ^ new_n16987;
  assign new_n17014 = new_n16992 ^ new_n16986;
  assign new_n17015 = new_n17014 ^ new_n16999;
  assign new_n17016 = new_n16977 & new_n17015;
  assign new_n17017 = new_n17003 ^ new_n16987;
  assign new_n17018 = new_n17008 ^ new_n17003;
  assign new_n17019 = new_n17018 ^ new_n16981;
  assign new_n17020 = new_n17019 ^ new_n16993;
  assign new_n17021 = new_n17017 & new_n17020;
  assign new_n17022 = new_n17021 ^ new_n17016;
  assign new_n17023 = new_n17007 ^ new_n16972;
  assign new_n17024 = new_n17023 ^ new_n16993;
  assign new_n17025 = new_n16992 ^ new_n16972;
  assign new_n17026 = new_n17024 & new_n17025;
  assign new_n17027 = new_n17026 ^ new_n16992;
  assign new_n17028 = new_n17027 ^ new_n17022;
  assign new_n17029 = new_n17028 ^ new_n17013;
  assign new_n17030 = ~new_n16981 & ~new_n17018;
  assign new_n17031 = new_n17030 ^ new_n16981;
  assign new_n17032 = new_n16981 ^ new_n16976;
  assign new_n17033 = new_n17014 ^ new_n17007;
  assign new_n17034 = new_n17032 & new_n17033;
  assign new_n17035 = new_n17034 ^ new_n17031;
  assign new_n17036 = new_n17035 ^ new_n16993;
  assign new_n17037 = new_n17026 ^ new_n17016;
  assign new_n17038 = new_n17007 ^ new_n16985;
  assign new_n17039 = new_n17038 ^ new_n17037;
  assign new_n17040 = new_n17039 ^ new_n17036;
  assign new_n17041 = ~new_n17040 & new_n17029;
  assign new_n17042 = new_n17041 ^ new_n17012;
  assign new_n17043 = new_n17008 ^ new_n16987;
  assign new_n17044 = new_n16993 & new_n17043;
  assign new_n17045 = new_n17044 ^ new_n17016;
  assign new_n17046 = new_n17045 ^ new_n17033;
  assign new_n17047 = new_n17046 ^ new_n17042;
  assign new_n17048 = new_n17018 ^ new_n16976;
  assign new_n17049 = new_n17015 ^ new_n17003;
  assign new_n17050 = new_n17048 & new_n17049;
  assign new_n17051 = new_n17050 ^ new_n17030;
  assign new_n17052 = new_n17044 ^ new_n17026;
  assign new_n17053 = new_n17052 ^ new_n17051;
  assign new_n17054 = ~new_n17053 & new_n17047;
  assign new_n17055 = new_n17050 ^ new_n17034;
  assign new_n17056 = new_n17055 ^ new_n16976;
  assign new_n17057 = new_n17056 ^ new_n17046;
  assign new_n17058 = new_n17057 ^ new_n17054;
  assign new_n17059 = new_n17018 ^ new_n16972;
  assign new_n17060 = new_n17058 & new_n17059;
  assign new_n17061 = new_n17007 ^ new_n16981;
  assign new_n17062 = new_n17031 ^ new_n17021;
  assign new_n17063 = new_n17054 ^ new_n17041;
  assign new_n17064 = ~new_n17063 & new_n17057;
  assign new_n17065 = new_n17064 ^ new_n17057;
  assign new_n17066 = new_n17007 ^ new_n16976;
  assign new_n17067 = new_n17011 ^ new_n16972;
  assign new_n17068 = new_n17067 ^ new_n17021;
  assign new_n17069 = new_n17068 ^ new_n17052;
  assign new_n17070 = new_n17069 ^ new_n17066;
  assign new_n17071 = new_n17057 ^ new_n17041;
  assign new_n17072 = new_n17070 & new_n17071;
  assign new_n17073 = new_n17072 ^ new_n17012;
  assign new_n17074 = new_n17073 ^ new_n17046;
  assign new_n17075 = new_n17064 ^ new_n17041;
  assign new_n17076 = new_n17074 & new_n17075;
  assign new_n17077 = new_n17076 ^ new_n17065;
  assign new_n17078 = new_n17077 ^ new_n17062;
  assign new_n17079 = new_n17078 ^ new_n17061;
  assign new_n17080 = new_n17079 ^ new_n16972;
  assign new_n17081 = new_n17072 ^ new_n17034;
  assign new_n17082 = new_n17081 ^ new_n17000;
  assign new_n17083 = new_n17082 ^ new_n17080;
  assign new_n17084 = ~new_n17083 & new_n17024;
  assign new_n17085 = new_n17076 ^ new_n17070;
  assign new_n17086 = new_n17018 & new_n17085;
  assign new_n17087 = new_n17065 ^ new_n17054;
  assign new_n17088 = new_n17087 ^ new_n17053;
  assign new_n17089 = ~new_n17088 & new_n17020;
  assign new_n17090 = ~new_n17083 & new_n17025;
  assign new_n17091 = new_n17072 ^ new_n17054;
  assign new_n17092 = new_n17056 ^ new_n17012;
  assign new_n17093 = new_n17092 ^ new_n17091;
  assign new_n17094 = new_n16977 & new_n17093;
  assign new_n17095 = new_n17094 ^ new_n17090;
  assign new_n17096 = new_n17095 ^ new_n17089;
  assign new_n17097 = new_n17096 ^ new_n17086;
  assign new_n17098 = new_n17076 ^ new_n17072;
  assign new_n17099 = new_n17098 ^ new_n17029;
  assign new_n17100 = new_n17033 & new_n17099;
  assign new_n17101 = new_n17100 ^ new_n17097;
  assign new_n17102 = new_n17101 ^ new_n17084;
  assign new_n17103 = new_n17102 ^ new_n17060;
  assign new_n17104 = new_n17003 & new_n17058;
  assign new_n17105 = new_n17065 ^ new_n17040;
  assign new_n17106 = ~new_n17105 & new_n16987;
  assign new_n17107 = new_n17106 ^ new_n17104;
  assign new_n17108 = new_n17032 & new_n17099;
  assign new_n17109 = new_n17108 ^ new_n17107;
  assign new_n17110 = new_n17048 & new_n17074;
  assign new_n17111 = new_n17054 ^ new_n16976;
  assign new_n17112 = new_n17067 ^ new_n17050;
  assign new_n17113 = new_n17112 ^ new_n17079;
  assign new_n17114 = new_n17113 ^ new_n17111;
  assign new_n17115 = ~new_n17114 & new_n17043;
  assign new_n17116 = new_n17115 ^ new_n17110;
  assign new_n17117 = new_n17116 ^ new_n17109;
  assign new_n17118 = new_n17117 ^ new_n17103;
  assign new_n17119 = new_n17118 ^ new_n16967;
  assign new_n17120 = new_n17119 ^ new_n16810;
  assign new_n17121 = new_n17120 ^ new_n16655;
  assign new_n17122 = ~new_n16529 & ~new_n16642;
  assign new_n17123 = ~new_n16625 & new_n16562;
  assign new_n17124 = new_n17123 ^ new_n17122;
  assign new_n17125 = new_n17124 ^ new_n16638;
  assign new_n17126 = new_n16782 ^ new_n16750;
  assign new_n17127 = ~new_n16731 & ~new_n17126;
  assign new_n17128 = ~new_n16736 & ~new_n16804;
  assign new_n17129 = new_n17128 ^ new_n17127;
  assign new_n17130 = new_n16782 ^ new_n16770;
  assign new_n17131 = new_n17130 ^ new_n16769;
  assign new_n17132 = ~new_n16716 & new_n17131;
  assign new_n17133 = new_n17132 ^ new_n16806;
  assign new_n17134 = new_n17133 ^ new_n16791;
  assign new_n17135 = ~new_n16744 & ~new_n16776;
  assign new_n17136 = new_n17135 ^ new_n17134;
  assign new_n17137 = new_n17136 ^ new_n16796;
  assign new_n17138 = new_n17137 ^ new_n17129;
  assign new_n17139 = new_n17138 ^ new_n17125;
  assign new_n17140 = new_n16770 ^ new_n16759;
  assign new_n17141 = ~new_n17140 & new_n16701;
  assign new_n17142 = ~new_n16697 & ~new_n17126;
  assign new_n17143 = new_n17142 ^ new_n17141;
  assign new_n17144 = new_n17143 ^ new_n16777;
  assign new_n17145 = new_n17144 ^ new_n17135;
  assign new_n17146 = new_n17145 ^ new_n16807;
  assign new_n17147 = new_n17146 ^ new_n17139;
  assign new_n17148 = new_n17115 ^ new_n17108;
  assign new_n17149 = new_n17086 ^ new_n17084;
  assign new_n17150 = new_n17019 & new_n17085;
  assign new_n17151 = new_n17049 & new_n17074;
  assign new_n17152 = new_n17151 ^ new_n17150;
  assign new_n17153 = new_n17152 ^ new_n17095;
  assign new_n17154 = new_n17153 ^ new_n17149;
  assign new_n17155 = new_n17154 ^ new_n17148;
  assign new_n17156 = new_n17155 ^ new_n16663;
  assign new_n17157 = new_n17156 ^ new_n17147;
  assign new_n17158 = new_n16496 ^ new_n16490;
  assign new_n17159 = new_n16482 ^ new_n16460;
  assign new_n17160 = ~new_n16459 & new_n16409;
  assign new_n17161 = ~new_n16433 & ~new_n16451;
  assign new_n17162 = new_n17161 ^ new_n17160;
  assign new_n17163 = new_n17162 ^ new_n16478;
  assign new_n17164 = new_n17163 ^ new_n17159;
  assign new_n17165 = new_n17164 ^ new_n17158;
  assign new_n17166 = new_n17165 ^ new_n16667;
  assign new_n17167 = new_n16645 ^ new_n16635;
  assign new_n17168 = new_n17167 ^ new_n16661;
  assign new_n17169 = new_n17168 ^ new_n17166;
  assign new_n17170 = new_n16964 ^ new_n16957;
  assign new_n17171 = new_n16938 ^ new_n16933;
  assign new_n17172 = ~new_n16937 & new_n16882;
  assign new_n17173 = ~new_n16900 & ~new_n16920;
  assign new_n17174 = new_n17173 ^ new_n17172;
  assign new_n17175 = new_n17174 ^ new_n16944;
  assign new_n17176 = new_n17175 ^ new_n17171;
  assign new_n17177 = new_n17176 ^ new_n17170;
  assign new_n17178 = new_n17177 ^ new_n17169;
  assign new_n17179 = new_n17178 ^ new_n17157;
  assign new_n17180 = ~new_n16395 & ~new_n16492;
  assign new_n17181 = new_n17180 ^ new_n17161;
  assign new_n17182 = ~new_n16462 & new_n16408;
  assign new_n17183 = new_n17182 ^ new_n16494;
  assign new_n17184 = new_n17183 ^ new_n16480;
  assign new_n17185 = new_n17184 ^ new_n17181;
  assign new_n17186 = new_n17185 ^ new_n16690;
  assign new_n17187 = new_n17186 ^ new_n17139;
  assign new_n17188 = ~new_n17105 & new_n16994;
  assign new_n17189 = new_n17188 ^ new_n17151;
  assign new_n17190 = ~new_n17088 & new_n17017;
  assign new_n17191 = new_n17190 ^ new_n17104;
  assign new_n17192 = new_n17191 ^ new_n17097;
  assign new_n17193 = new_n17192 ^ new_n17189;
  assign new_n17194 = ~new_n16877 & ~new_n16954;
  assign new_n17195 = new_n17194 ^ new_n17173;
  assign new_n17196 = ~new_n16946 & new_n16881;
  assign new_n17197 = new_n17196 ^ new_n16953;
  assign new_n17198 = new_n17197 ^ new_n16949;
  assign new_n17199 = new_n17198 ^ new_n17195;
  assign new_n17200 = new_n17199 ^ new_n17193;
  assign new_n17201 = new_n17200 ^ new_n17187;
  assign new_n17202 = ~new_n17140 & new_n16718;
  assign new_n17203 = new_n17202 ^ new_n17137;
  assign new_n17204 = new_n16754 & new_n16765;
  assign new_n17205 = new_n17204 ^ new_n16788;
  assign new_n17206 = new_n17205 ^ new_n17144;
  assign new_n17207 = new_n17206 ^ new_n17203;
  assign new_n17208 = new_n17122 ^ new_n16659;
  assign new_n17209 = ~new_n16629 & new_n16571;
  assign new_n17210 = new_n17209 ^ new_n16641;
  assign new_n17211 = new_n17210 ^ new_n16632;
  assign new_n17212 = new_n17211 ^ new_n17208;
  assign new_n17213 = new_n17212 ^ new_n17207;
  assign new_n17214 = new_n17213 ^ new_n16654;
  assign new_n17215 = new_n17214 ^ new_n17201;
  assign new_n17216 = new_n17215 ^ new_n17179;
  assign new_n17217 = new_n17216 ^ new_n17121;
  assign new_n17218 = ~new_n16941 & new_n16870;
  assign new_n17219 = new_n17218 ^ new_n16933;
  assign new_n17220 = new_n17196 ^ new_n16955;
  assign new_n17221 = new_n17220 ^ new_n17194;
  assign new_n17222 = new_n17221 ^ new_n16948;
  assign new_n17223 = new_n17222 ^ new_n17219;
  assign new_n17224 = new_n17015 & new_n17093;
  assign new_n17225 = new_n17224 ^ new_n17084;
  assign new_n17226 = new_n17190 ^ new_n17106;
  assign new_n17227 = new_n17226 ^ new_n17188;
  assign new_n17228 = new_n17227 ^ new_n17096;
  assign new_n17229 = new_n17228 ^ new_n17225;
  assign new_n17230 = new_n17229 ^ new_n17223;
  assign new_n17231 = new_n17128 ^ new_n16805;
  assign new_n17232 = ~new_n16715 & ~new_n16787;
  assign new_n17233 = new_n17232 ^ new_n17206;
  assign new_n17234 = new_n17233 ^ new_n17231;
  assign new_n17235 = new_n17234 ^ new_n17230;
  assign new_n17236 = ~new_n16466 & new_n16401;
  assign new_n17237 = new_n17236 ^ new_n16482;
  assign new_n17238 = new_n17182 ^ new_n16493;
  assign new_n17239 = new_n17238 ^ new_n17180;
  assign new_n17240 = new_n17239 ^ new_n16479;
  assign new_n17241 = new_n17240 ^ new_n17237;
  assign new_n17242 = new_n17241 ^ new_n16704;
  assign new_n17243 = new_n17123 ^ new_n16637;
  assign new_n17244 = new_n17209 ^ new_n16643;
  assign new_n17245 = new_n17244 ^ new_n17122;
  assign new_n17246 = new_n17245 ^ new_n16631;
  assign new_n17247 = new_n17246 ^ new_n17243;
  assign new_n17248 = new_n17247 ^ new_n17242;
  assign new_n17249 = new_n17123 ^ new_n16626;
  assign new_n17250 = new_n16528 & new_n16649;
  assign new_n17251 = new_n17250 ^ new_n16653;
  assign new_n17252 = new_n17251 ^ new_n17249;
  assign new_n17253 = new_n17252 ^ new_n17248;
  assign new_n17254 = new_n17253 ^ new_n17235;
  assign new_n17255 = new_n17254 ^ new_n17217;
  assign new_n17256 = new_n17218 ^ new_n16942;
  assign new_n17257 = new_n16863 & new_n16963;
  assign new_n17258 = new_n17257 ^ new_n16966;
  assign new_n17259 = new_n17258 ^ new_n17256;
  assign new_n17260 = new_n17224 ^ new_n17094;
  assign new_n17261 = ~new_n17114 & new_n16993;
  assign new_n17262 = new_n17261 ^ new_n17117;
  assign new_n17263 = new_n17262 ^ new_n17260;
  assign new_n17264 = new_n17263 ^ new_n17259;
  assign new_n17265 = new_n17264 ^ new_n17252;
  assign new_n17266 = new_n17236 ^ new_n16467;
  assign new_n17267 = new_n16394 & new_n16489;
  assign new_n17268 = new_n17267 ^ new_n16498;
  assign new_n17269 = new_n17268 ^ new_n17266;
  assign new_n17270 = new_n17269 ^ new_n16678;
  assign new_n17271 = ~new_n16702 & new_n17131;
  assign new_n17272 = new_n17271 ^ new_n17142;
  assign new_n17273 = new_n17272 ^ new_n17127;
  assign new_n17274 = new_n17273 ^ new_n17136;
  assign new_n17275 = new_n17245 ^ new_n16636;
  assign new_n17276 = new_n17275 ^ new_n17274;
  assign new_n17277 = new_n17276 ^ new_n17270;
  assign new_n17278 = new_n17277 ^ new_n17265;
  assign new_n17279 = new_n17278 ^ new_n17217;
  assign new_n17280 = new_n17224 ^ new_n17188;
  assign new_n17281 = new_n17280 ^ new_n17102;
  assign new_n17282 = new_n17218 ^ new_n17194;
  assign new_n17283 = new_n17282 ^ new_n16951;
  assign new_n17284 = new_n17283 ^ new_n17281;
  assign new_n17285 = new_n17128 ^ new_n16796;
  assign new_n17286 = new_n17273 ^ new_n17133;
  assign new_n17287 = new_n17286 ^ new_n17285;
  assign new_n17288 = new_n17287 ^ new_n17284;
  assign new_n17289 = new_n17236 ^ new_n17180;
  assign new_n17290 = new_n17289 ^ new_n16483;
  assign new_n17291 = new_n17290 ^ new_n16672;
  assign new_n17292 = new_n17291 ^ new_n17125;
  assign new_n17293 = new_n17292 ^ new_n17247;
  assign new_n17294 = new_n17293 ^ new_n17288;
  assign new_n17295 = new_n17294 ^ new_n17179;
  assign new_n17296 = ~new_n17279 & ~new_n17295;
  assign new_n17297 = new_n16497 ^ new_n16458;
  assign new_n17298 = new_n17297 ^ new_n17163;
  assign new_n17299 = new_n17298 ^ new_n16698;
  assign new_n17300 = new_n16958 ^ new_n16936;
  assign new_n17301 = new_n17300 ^ new_n17175;
  assign new_n17302 = new_n17301 ^ new_n17299;
  assign new_n17303 = new_n17109 ^ new_n17100;
  assign new_n17304 = new_n17303 ^ new_n17153;
  assign new_n17305 = new_n17304 ^ new_n17168;
  assign new_n17306 = new_n17305 ^ new_n17139;
  assign new_n17307 = new_n17306 ^ new_n17302;
  assign new_n17308 = new_n17278 ^ new_n17254;
  assign new_n17309 = new_n17308 ^ new_n17307;
  assign new_n17310 = new_n17179 & new_n17309;
  assign new_n17311 = new_n17310 ^ new_n17179;
  assign new_n17312 = new_n17311 ^ new_n17296;
  assign new_n17313 = new_n17294 ^ new_n17121;
  assign new_n17314 = new_n17313 ^ new_n17312;
  assign new_n17315 = new_n17239 ^ new_n16481;
  assign new_n17316 = new_n17315 ^ new_n16683;
  assign new_n17317 = new_n17227 ^ new_n17101;
  assign new_n17318 = new_n17221 ^ new_n16950;
  assign new_n17319 = new_n17318 ^ new_n17317;
  assign new_n17320 = new_n17319 ^ new_n17316;
  assign new_n17321 = new_n17320 ^ new_n17139;
  assign new_n17322 = new_n17127 ^ new_n16799;
  assign new_n17323 = new_n17271 ^ new_n17141;
  assign new_n17324 = new_n17323 ^ new_n17134;
  assign new_n17325 = new_n17324 ^ new_n17322;
  assign new_n17326 = new_n17325 ^ new_n17275;
  assign new_n17327 = new_n17326 ^ new_n17212;
  assign new_n17328 = new_n17327 ^ new_n17321;
  assign new_n17329 = new_n17328 ^ new_n17294;
  assign new_n17330 = ~new_n17255 & ~new_n17329;
  assign new_n17331 = new_n17328 ^ new_n17278;
  assign new_n17332 = new_n17331 ^ new_n17313;
  assign new_n17333 = new_n17328 ^ new_n17121;
  assign new_n17334 = new_n17332 & new_n17333;
  assign new_n17335 = new_n17334 ^ new_n17330;
  assign new_n17336 = new_n17278 ^ new_n17215;
  assign new_n17337 = new_n17336 ^ new_n17335;
  assign new_n17338 = new_n17337 ^ new_n17314;
  assign new_n17339 = new_n17329 ^ new_n17216;
  assign new_n17340 = new_n17328 ^ new_n17179;
  assign new_n17341 = new_n17340 ^ new_n17313;
  assign new_n17342 = ~new_n17339 & ~new_n17341;
  assign new_n17343 = new_n17342 ^ new_n17254;
  assign new_n17344 = new_n17343 ^ new_n17339;
  assign new_n17345 = new_n17339 ^ new_n17307;
  assign new_n17346 = new_n17309 ^ new_n17179;
  assign new_n17347 = new_n17346 ^ new_n17313;
  assign new_n17348 = ~new_n17347 & new_n17345;
  assign new_n17349 = new_n17348 ^ new_n17121;
  assign new_n17350 = new_n17349 ^ new_n17335;
  assign new_n17351 = new_n17350 ^ new_n17344;
  assign new_n17352 = new_n17338 & new_n17351;
  assign new_n17353 = new_n17328 ^ new_n17309;
  assign new_n17354 = ~new_n17307 & new_n17353;
  assign new_n17355 = new_n17354 ^ new_n17328;
  assign new_n17356 = new_n17355 ^ new_n17343;
  assign new_n17357 = new_n17356 ^ new_n17352;
  assign new_n17358 = new_n17339 ^ new_n17308;
  assign new_n17359 = ~new_n17313 & ~new_n17358;
  assign new_n17360 = new_n17359 ^ new_n17330;
  assign new_n17361 = new_n17360 ^ new_n17279;
  assign new_n17362 = new_n17361 ^ new_n17357;
  assign new_n17363 = new_n17309 ^ new_n17294;
  assign new_n17364 = new_n17307 ^ new_n17255;
  assign new_n17365 = ~new_n17363 & new_n17364;
  assign new_n17366 = new_n17365 ^ new_n17310;
  assign new_n17367 = new_n17359 ^ new_n17334;
  assign new_n17368 = new_n17367 ^ new_n17366;
  assign new_n17369 = ~new_n17368 & new_n17362;
  assign new_n17370 = new_n17294 ^ new_n17278;
  assign new_n17371 = new_n17354 ^ new_n17348;
  assign new_n17372 = new_n17371 ^ new_n17367;
  assign new_n17373 = new_n17372 ^ new_n17370;
  assign new_n17374 = new_n17365 ^ new_n17296;
  assign new_n17375 = new_n17374 ^ new_n17294;
  assign new_n17376 = new_n17375 ^ new_n17361;
  assign new_n17377 = new_n17376 ^ new_n17352;
  assign new_n17378 = ~new_n17377 & new_n17373;
  assign new_n17379 = new_n17378 ^ new_n17369;
  assign new_n17380 = new_n17375 ^ new_n17356;
  assign new_n17381 = new_n17380 ^ new_n17379;
  assign new_n17382 = ~new_n17255 & ~new_n17381;
  assign new_n17383 = new_n17278 ^ new_n17179;
  assign new_n17384 = new_n17348 ^ new_n17311;
  assign new_n17385 = new_n17378 ^ new_n17356;
  assign new_n17386 = new_n17385 ^ new_n17361;
  assign new_n17387 = new_n17369 ^ new_n17352;
  assign new_n17388 = ~new_n17376 & new_n17387;
  assign new_n17389 = new_n17388 ^ new_n17377;
  assign new_n17390 = ~new_n17389 & new_n17386;
  assign new_n17391 = new_n17390 ^ new_n17388;
  assign new_n17392 = new_n17391 ^ new_n17384;
  assign new_n17393 = new_n17392 ^ new_n17383;
  assign new_n17394 = new_n17393 ^ new_n17328;
  assign new_n17395 = new_n17378 ^ new_n17296;
  assign new_n17396 = new_n17395 ^ new_n17343;
  assign new_n17397 = new_n17396 ^ new_n17394;
  assign new_n17398 = new_n17332 & new_n17397;
  assign new_n17399 = new_n17398 ^ new_n17382;
  assign new_n17400 = new_n17388 ^ new_n17369;
  assign new_n17401 = new_n17400 ^ new_n17368;
  assign new_n17402 = ~new_n17401 & new_n17345;
  assign new_n17403 = new_n17388 ^ new_n17338;
  assign new_n17404 = ~new_n17339 & new_n17403;
  assign new_n17405 = new_n17404 ^ new_n17402;
  assign new_n17406 = ~new_n17341 & new_n17403;
  assign new_n17407 = new_n17406 ^ new_n17405;
  assign new_n17408 = ~new_n17329 & ~new_n17381;
  assign new_n17409 = new_n17333 & new_n17397;
  assign new_n17410 = new_n17409 ^ new_n17408;
  assign new_n17411 = ~new_n17347 & ~new_n17401;
  assign new_n17412 = new_n17411 ^ new_n17410;
  assign new_n17413 = new_n17412 ^ new_n17407;
  assign new_n17414 = new_n17413 ^ new_n17399;
  assign new_n17415 = new_n17414 ^ new_n16383;
  assign new_n17416 = new_n14079 ^ n14;
  assign new_n17417 = new_n14848 ^ n12;
  assign new_n17418 = new_n17417 ^ new_n17416;
  assign new_n17419 = new_n14791 ^ n15;
  assign new_n17420 = new_n14857 ^ n9;
  assign new_n17421 = new_n17420 ^ new_n17419;
  assign new_n17422 = new_n17421 ^ new_n17418;
  assign new_n17423 = new_n14809 ^ n13;
  assign new_n17424 = new_n17423 ^ new_n17419;
  assign new_n17425 = new_n17424 ^ new_n17416;
  assign new_n17426 = new_n14675 ^ n11;
  assign new_n17427 = new_n17426 ^ new_n17425;
  assign new_n17428 = ~new_n17421 & new_n17427;
  assign new_n17429 = new_n14097 ^ n10;
  assign new_n17430 = new_n17429 ^ new_n17425;
  assign new_n17431 = new_n14877 ^ n16;
  assign new_n17432 = new_n17431 ^ new_n17430;
  assign new_n17433 = new_n17429 ^ new_n17426;
  assign new_n17434 = new_n17433 ^ new_n17431;
  assign new_n17435 = new_n17434 ^ new_n17420;
  assign new_n17436 = ~new_n17432 & ~new_n17435;
  assign new_n17437 = new_n17436 ^ new_n17428;
  assign new_n17438 = new_n17437 ^ new_n17420;
  assign new_n17439 = new_n17420 ^ new_n17416;
  assign new_n17440 = new_n17420 ^ new_n17417;
  assign new_n17441 = new_n17440 ^ new_n17424;
  assign new_n17442 = new_n17441 ^ new_n17433;
  assign new_n17443 = ~new_n17442 & new_n17439;
  assign new_n17444 = new_n17430 & new_n17440;
  assign new_n17445 = new_n17444 ^ new_n17443;
  assign new_n17446 = new_n17445 ^ new_n17427;
  assign new_n17447 = new_n17446 ^ new_n17438;
  assign new_n17448 = ~new_n17422 & ~new_n17441;
  assign new_n17449 = new_n17448 ^ new_n17429;
  assign new_n17450 = new_n17449 ^ new_n17441;
  assign new_n17451 = new_n17426 ^ new_n17417;
  assign new_n17452 = new_n17451 ^ new_n17439;
  assign new_n17453 = ~new_n17452 & new_n17418;
  assign new_n17454 = new_n17453 ^ new_n17444;
  assign new_n17455 = new_n17441 ^ new_n17431;
  assign new_n17456 = new_n17434 ^ new_n17419;
  assign new_n17457 = new_n17456 ^ new_n17439;
  assign new_n17458 = new_n17455 & new_n17457;
  assign new_n17459 = new_n17458 ^ new_n17416;
  assign new_n17460 = new_n17459 ^ new_n17454;
  assign new_n17461 = new_n17460 ^ new_n17450;
  assign new_n17462 = new_n17419 & new_n17434;
  assign new_n17463 = new_n17462 ^ new_n17419;
  assign new_n17464 = new_n17463 ^ new_n17428;
  assign new_n17465 = new_n17464 ^ new_n17439;
  assign new_n17466 = new_n17426 ^ new_n17423;
  assign new_n17467 = new_n17466 ^ new_n17454;
  assign new_n17468 = new_n17467 ^ new_n17465;
  assign new_n17469 = ~new_n17468 & new_n17461;
  assign new_n17470 = new_n17434 ^ new_n17417;
  assign new_n17471 = ~new_n17431 & ~new_n17470;
  assign new_n17472 = new_n17471 ^ new_n17417;
  assign new_n17473 = new_n17472 ^ new_n17449;
  assign new_n17474 = new_n17473 ^ new_n17469;
  assign new_n17475 = new_n17474 ^ new_n17446;
  assign new_n17476 = new_n17453 ^ new_n17443;
  assign new_n17477 = new_n17462 ^ new_n17436;
  assign new_n17478 = new_n17477 ^ new_n17476;
  assign new_n17479 = ~new_n17475 & ~new_n17478;
  assign new_n17480 = new_n17479 ^ new_n17469;
  assign new_n17481 = ~new_n17480 & new_n17447;
  assign new_n17482 = new_n17481 ^ new_n17447;
  assign new_n17483 = new_n17482 ^ new_n17468;
  assign new_n17484 = ~new_n17422 & ~new_n17483;
  assign new_n17485 = new_n17426 ^ new_n17420;
  assign new_n17486 = new_n17471 ^ new_n17458;
  assign new_n17487 = new_n17486 ^ new_n17476;
  assign new_n17488 = new_n17487 ^ new_n17485;
  assign new_n17489 = new_n17469 ^ new_n17447;
  assign new_n17490 = ~new_n17488 & new_n17489;
  assign new_n17491 = new_n17490 ^ new_n17473;
  assign new_n17492 = new_n17491 ^ new_n17446;
  assign new_n17493 = ~new_n17432 & ~new_n17492;
  assign new_n17494 = new_n17493 ^ new_n17484;
  assign new_n17495 = new_n17482 ^ new_n17479;
  assign new_n17496 = new_n17495 ^ new_n17478;
  assign new_n17497 = ~new_n17496 & new_n17455;
  assign new_n17498 = new_n17479 ^ new_n17447;
  assign new_n17499 = ~new_n17431 & new_n17498;
  assign new_n17500 = new_n17499 ^ new_n17497;
  assign new_n17501 = new_n17481 ^ new_n17469;
  assign new_n17502 = ~new_n17492 & new_n17501;
  assign new_n17503 = new_n17502 ^ new_n17488;
  assign new_n17504 = ~new_n17434 & ~new_n17503;
  assign new_n17505 = ~new_n17496 & new_n17457;
  assign new_n17506 = new_n17426 ^ new_n17419;
  assign new_n17507 = new_n17463 ^ new_n17458;
  assign new_n17508 = new_n17502 ^ new_n17482;
  assign new_n17509 = new_n17508 ^ new_n17507;
  assign new_n17510 = new_n17509 ^ new_n17506;
  assign new_n17511 = new_n17510 ^ new_n17417;
  assign new_n17512 = new_n17490 ^ new_n17428;
  assign new_n17513 = new_n17512 ^ new_n17449;
  assign new_n17514 = new_n17513 ^ new_n17511;
  assign new_n17515 = ~new_n17514 & new_n17418;
  assign new_n17516 = new_n17490 ^ new_n17479;
  assign new_n17517 = new_n17473 ^ new_n17438;
  assign new_n17518 = new_n17517 ^ new_n17516;
  assign new_n17519 = ~new_n17518 & new_n17440;
  assign new_n17520 = new_n17519 ^ new_n17515;
  assign new_n17521 = new_n17520 ^ new_n17505;
  assign new_n17522 = new_n17521 ^ new_n17504;
  assign new_n17523 = new_n17522 ^ new_n17500;
  assign new_n17524 = new_n17523 ^ new_n17494;
  assign new_n17525 = new_n17524 ^ new_n1175;
  assign new_n17526 = new_n17479 ^ new_n17420;
  assign new_n17527 = new_n17471 ^ new_n17436;
  assign new_n17528 = new_n17527 ^ new_n17510;
  assign new_n17529 = new_n17528 ^ new_n17526;
  assign new_n17530 = ~new_n17442 & new_n17529;
  assign new_n17531 = new_n17502 ^ new_n17490;
  assign new_n17532 = new_n17531 ^ new_n17461;
  assign new_n17533 = ~new_n17421 & new_n17532;
  assign new_n17534 = new_n17533 ^ new_n17530;
  assign new_n17535 = ~new_n17452 & ~new_n17514;
  assign new_n17536 = new_n17535 ^ new_n17504;
  assign new_n17537 = ~new_n17503 & new_n17456;
  assign new_n17538 = new_n17537 ^ new_n17493;
  assign new_n17539 = new_n17538 ^ new_n17520;
  assign new_n17540 = new_n17539 ^ new_n17536;
  assign new_n17541 = new_n17540 ^ new_n17534;
  assign new_n17542 = new_n17541 ^ new_n1183;
  assign new_n17543 = new_n17542 ^ new_n17525;
  assign new_n17544 = ~new_n17470 & new_n17498;
  assign new_n17545 = new_n17427 & new_n17532;
  assign new_n17546 = new_n17545 ^ new_n17522;
  assign new_n17547 = new_n17546 ^ new_n17535;
  assign new_n17548 = new_n17547 ^ new_n17544;
  assign new_n17549 = ~new_n17435 & ~new_n17492;
  assign new_n17550 = new_n17549 ^ new_n17530;
  assign new_n17551 = ~new_n17441 & ~new_n17483;
  assign new_n17552 = new_n17551 ^ new_n17499;
  assign new_n17553 = new_n17552 ^ new_n17533;
  assign new_n17554 = new_n17553 ^ new_n17550;
  assign new_n17555 = new_n17554 ^ new_n17548;
  assign new_n17556 = new_n17555 ^ new_n1202;
  assign new_n17557 = new_n17556 ^ new_n17543;
  assign new_n17558 = ~new_n17518 & new_n17430;
  assign new_n17559 = new_n17558 ^ new_n17535;
  assign new_n17560 = new_n17551 ^ new_n17497;
  assign new_n17561 = new_n17560 ^ new_n17484;
  assign new_n17562 = new_n17561 ^ new_n17521;
  assign new_n17563 = new_n17562 ^ new_n17559;
  assign new_n17564 = new_n17563 ^ new_n1119;
  assign new_n17565 = new_n17564 ^ new_n17557;
  assign new_n17566 = new_n17558 ^ new_n17484;
  assign new_n17567 = new_n17566 ^ new_n17547;
  assign new_n17568 = new_n17567 ^ new_n1191;
  assign new_n17569 = new_n17558 ^ new_n17519;
  assign new_n17570 = new_n17439 & new_n17529;
  assign new_n17571 = new_n17570 ^ new_n17554;
  assign new_n17572 = new_n17571 ^ new_n17569;
  assign new_n17573 = new_n17572 ^ new_n1142;
  assign new_n17574 = new_n17573 ^ new_n17568;
  assign new_n17575 = new_n17561 ^ new_n17546;
  assign new_n17576 = new_n17575 ^ new_n1164;
  assign new_n17577 = new_n17576 ^ new_n17568;
  assign new_n17578 = new_n17577 ^ new_n17543;
  assign new_n17579 = new_n17553 ^ new_n17545;
  assign new_n17580 = new_n17579 ^ new_n17539;
  assign new_n17581 = new_n17580 ^ new_n1155;
  assign new_n17582 = new_n17581 ^ new_n17578;
  assign new_n17583 = new_n17573 ^ new_n17564;
  assign new_n17584 = new_n17583 ^ new_n17581;
  assign new_n17585 = new_n17584 ^ new_n17542;
  assign new_n17586 = new_n17568 ^ new_n17556;
  assign new_n17587 = new_n17586 ^ new_n17585;
  assign new_n17588 = new_n17582 & new_n17587;
  assign new_n17589 = new_n17584 ^ new_n17576;
  assign new_n17590 = new_n17581 & new_n17589;
  assign new_n17591 = new_n17590 ^ new_n17588;
  assign new_n17592 = new_n17583 ^ new_n17578;
  assign new_n17593 = new_n17586 & new_n17592;
  assign new_n17594 = new_n17576 ^ new_n17556;
  assign new_n17595 = new_n17576 ^ new_n17573;
  assign new_n17596 = new_n17595 ^ new_n17586;
  assign new_n17597 = new_n17594 & new_n17596;
  assign new_n17598 = new_n17597 ^ new_n17593;
  assign new_n17599 = new_n17598 ^ new_n17591;
  assign new_n17600 = new_n17599 ^ new_n17574;
  assign new_n17601 = new_n17584 ^ new_n17568;
  assign new_n17602 = new_n17581 ^ new_n17565;
  assign new_n17603 = new_n17601 & new_n17602;
  assign new_n17604 = new_n17573 ^ new_n17557;
  assign new_n17605 = new_n17568 ^ new_n17542;
  assign new_n17606 = new_n17604 & new_n17605;
  assign new_n17607 = new_n17606 ^ new_n17603;
  assign new_n17608 = new_n17607 ^ new_n17568;
  assign new_n17609 = new_n17565 & new_n17577;
  assign new_n17610 = new_n17609 ^ new_n17593;
  assign new_n17611 = new_n17610 ^ new_n17604;
  assign new_n17612 = new_n17611 ^ new_n17608;
  assign new_n17613 = new_n17576 ^ new_n17542;
  assign new_n17614 = new_n17613 ^ new_n17586;
  assign new_n17615 = new_n17578 & new_n17614;
  assign new_n17616 = new_n17615 ^ new_n17564;
  assign new_n17617 = new_n17616 ^ new_n17578;
  assign new_n17618 = new_n17609 ^ new_n17597;
  assign new_n17619 = new_n17588 ^ new_n17556;
  assign new_n17620 = new_n17619 ^ new_n17618;
  assign new_n17621 = new_n17620 ^ new_n17617;
  assign new_n17622 = ~new_n17542 & ~new_n17584;
  assign new_n17623 = new_n17622 ^ new_n17542;
  assign new_n17624 = new_n17623 ^ new_n17606;
  assign new_n17625 = new_n17624 ^ new_n17586;
  assign new_n17626 = new_n17573 ^ new_n17525;
  assign new_n17627 = new_n17626 ^ new_n17618;
  assign new_n17628 = new_n17627 ^ new_n17625;
  assign new_n17629 = ~new_n17628 & new_n17621;
  assign new_n17630 = new_n17629 ^ new_n17612;
  assign new_n17631 = new_n17600 & new_n17630;
  assign new_n17632 = new_n17590 ^ new_n17576;
  assign new_n17633 = new_n17632 ^ new_n17616;
  assign new_n17634 = new_n17633 ^ new_n17629;
  assign new_n17635 = new_n17634 ^ new_n17611;
  assign new_n17636 = new_n17622 ^ new_n17603;
  assign new_n17637 = new_n17636 ^ new_n17598;
  assign new_n17638 = ~new_n17637 & new_n17635;
  assign new_n17639 = new_n17638 ^ new_n17631;
  assign new_n17640 = new_n17633 ^ new_n17608;
  assign new_n17641 = new_n17640 ^ new_n17639;
  assign new_n17642 = new_n17565 & new_n17641;
  assign new_n17643 = new_n17638 ^ new_n17629;
  assign new_n17644 = ~new_n17643 & new_n17612;
  assign new_n17645 = new_n17644 ^ new_n17612;
  assign new_n17646 = new_n17645 ^ new_n17628;
  assign new_n17647 = ~new_n17646 & new_n17614;
  assign new_n17648 = new_n17647 ^ new_n17642;
  assign new_n17649 = new_n17645 ^ new_n17638;
  assign new_n17650 = new_n17649 ^ new_n17637;
  assign new_n17651 = ~new_n17650 & new_n17587;
  assign new_n17652 = new_n17573 ^ new_n17542;
  assign new_n17653 = new_n17623 ^ new_n17588;
  assign new_n17654 = new_n17633 ^ new_n17631;
  assign new_n17655 = new_n17654 ^ new_n17611;
  assign new_n17656 = new_n17644 ^ new_n17629;
  assign new_n17657 = new_n17655 & new_n17656;
  assign new_n17658 = new_n17657 ^ new_n17645;
  assign new_n17659 = new_n17658 ^ new_n17653;
  assign new_n17660 = new_n17659 ^ new_n17652;
  assign new_n17661 = new_n17660 ^ new_n17576;
  assign new_n17662 = new_n17631 ^ new_n17606;
  assign new_n17663 = new_n17662 ^ new_n17616;
  assign new_n17664 = new_n17663 ^ new_n17661;
  assign new_n17665 = ~new_n17664 & new_n17594;
  assign new_n17666 = new_n17577 & new_n17641;
  assign new_n17667 = new_n17666 ^ new_n17665;
  assign new_n17668 = new_n17667 ^ new_n17651;
  assign new_n17669 = new_n17657 ^ new_n17600;
  assign new_n17670 = new_n17584 & new_n17669;
  assign new_n17671 = new_n17670 ^ new_n17668;
  assign new_n17672 = new_n17657 ^ new_n17631;
  assign new_n17673 = new_n17672 ^ new_n17621;
  assign new_n17674 = new_n17604 & new_n17673;
  assign new_n17675 = new_n17674 ^ new_n17671;
  assign new_n17676 = ~new_n17664 & new_n17596;
  assign new_n17677 = new_n17676 ^ new_n17675;
  assign new_n17678 = new_n17677 ^ new_n17648;
  assign new_n17679 = new_n17678 ^ new_n17291;
  assign new_n17680 = new_n17555 ^ new_n14103;
  assign new_n17681 = new_n12868 ^ new_n8532;
  assign new_n17682 = new_n17681 ^ new_n15763;
  assign new_n17683 = new_n17682 ^ new_n15786;
  assign new_n17684 = new_n11513 ^ new_n11473;
  assign new_n17685 = new_n17684 ^ new_n11486;
  assign new_n17686 = new_n17685 ^ new_n17683;
  assign new_n17687 = new_n15769 ^ new_n8060;
  assign new_n17688 = new_n13550 ^ new_n8541;
  assign new_n17689 = new_n17688 ^ new_n15760;
  assign new_n17690 = new_n17689 ^ new_n17687;
  assign new_n17691 = new_n15784 ^ new_n10181;
  assign new_n17692 = new_n13572 ^ new_n8546;
  assign new_n17693 = new_n17692 ^ new_n11369;
  assign new_n17694 = new_n17693 ^ new_n8060;
  assign new_n17695 = new_n17694 ^ new_n17691;
  assign new_n17696 = new_n17695 ^ new_n17690;
  assign new_n17697 = new_n13601 ^ new_n8552;
  assign new_n17698 = new_n17697 ^ new_n11448;
  assign new_n17699 = new_n15798 ^ new_n15786;
  assign new_n17700 = new_n17699 ^ new_n17698;
  assign new_n17701 = new_n17700 ^ new_n17696;
  assign new_n17702 = new_n17701 ^ new_n17686;
  assign new_n17703 = new_n15809 ^ new_n11431;
  assign new_n17704 = new_n17703 ^ new_n15786;
  assign new_n17705 = new_n13640 ^ new_n8563;
  assign new_n17706 = new_n17705 ^ new_n11530;
  assign new_n17707 = new_n17706 ^ new_n11448;
  assign new_n17708 = new_n17707 ^ new_n17704;
  assign new_n17709 = ~new_n17708 & new_n17701;
  assign new_n17710 = new_n17709 ^ new_n17708;
  assign new_n17711 = new_n13684 ^ new_n8580;
  assign new_n17712 = new_n17711 ^ new_n15758;
  assign new_n17713 = new_n17712 ^ new_n15786;
  assign new_n17714 = new_n11571 ^ new_n11513;
  assign new_n17715 = new_n17714 ^ new_n11494;
  assign new_n17716 = new_n17715 ^ new_n17713;
  assign new_n17717 = new_n17716 ^ new_n17708;
  assign new_n17718 = new_n15794 ^ new_n11541;
  assign new_n17719 = new_n13669 ^ new_n8588;
  assign new_n17720 = new_n17719 ^ new_n11571;
  assign new_n17721 = new_n17720 ^ new_n11530;
  assign new_n17722 = new_n17721 ^ new_n17718;
  assign new_n17723 = new_n17722 ^ new_n17717;
  assign new_n17724 = new_n17723 ^ new_n17690;
  assign new_n17725 = new_n15756 ^ new_n11412;
  assign new_n17726 = new_n13713 ^ new_n8571;
  assign new_n17727 = new_n17726 ^ new_n11551;
  assign new_n17728 = new_n17727 ^ new_n11369;
  assign new_n17729 = new_n17728 ^ new_n17725;
  assign new_n17730 = new_n17729 ^ new_n17708;
  assign new_n17731 = new_n17724 & new_n17730;
  assign new_n17732 = new_n17731 ^ new_n17710;
  assign new_n17733 = new_n17729 ^ new_n17722;
  assign new_n17734 = new_n17733 ^ new_n17732;
  assign new_n17735 = new_n17723 ^ new_n17695;
  assign new_n17736 = new_n17729 ^ new_n17686;
  assign new_n17737 = new_n17735 & new_n17736;
  assign new_n17738 = new_n17690 ^ new_n17686;
  assign new_n17739 = new_n17738 ^ new_n17733;
  assign new_n17740 = new_n17722 ^ new_n17686;
  assign new_n17741 = ~new_n17739 & new_n17740;
  assign new_n17742 = new_n17741 ^ new_n17737;
  assign new_n17743 = new_n17716 ^ new_n17690;
  assign new_n17744 = new_n17743 ^ new_n17742;
  assign new_n17745 = new_n17744 ^ new_n17734;
  assign new_n17746 = new_n17736 ^ new_n17717;
  assign new_n17747 = new_n17708 ^ new_n17686;
  assign new_n17748 = new_n17747 ^ new_n17733;
  assign new_n17749 = ~new_n17746 & new_n17748;
  assign new_n17750 = new_n17749 ^ new_n17695;
  assign new_n17751 = new_n17750 ^ new_n17746;
  assign new_n17752 = new_n17746 ^ new_n17700;
  assign new_n17753 = new_n17708 ^ new_n17701;
  assign new_n17754 = new_n17753 ^ new_n17733;
  assign new_n17755 = ~new_n17754 & new_n17752;
  assign new_n17756 = new_n17755 ^ new_n17737;
  assign new_n17757 = new_n17741 ^ new_n17722;
  assign new_n17758 = new_n17757 ^ new_n17756;
  assign new_n17759 = new_n17758 ^ new_n17751;
  assign new_n17760 = ~new_n17745 & new_n17759;
  assign new_n17761 = ~new_n17700 & ~new_n17702;
  assign new_n17762 = new_n17761 ^ new_n17686;
  assign new_n17763 = new_n17762 ^ new_n17750;
  assign new_n17764 = new_n17763 ^ new_n17760;
  assign new_n17765 = new_n17746 ^ new_n17696;
  assign new_n17766 = ~new_n17765 & new_n17733;
  assign new_n17767 = new_n17766 ^ new_n17737;
  assign new_n17768 = new_n17767 ^ new_n17724;
  assign new_n17769 = new_n17768 ^ new_n17764;
  assign new_n17770 = new_n17729 ^ new_n17701;
  assign new_n17771 = new_n17735 ^ new_n17700;
  assign new_n17772 = ~new_n17770 & ~new_n17771;
  assign new_n17773 = new_n17772 ^ new_n17709;
  assign new_n17774 = new_n17766 ^ new_n17741;
  assign new_n17775 = new_n17774 ^ new_n17773;
  assign new_n17776 = ~new_n17769 & ~new_n17775;
  assign new_n17777 = new_n17772 ^ new_n17731;
  assign new_n17778 = new_n17777 ^ new_n17729;
  assign new_n17779 = new_n17778 ^ new_n17768;
  assign new_n17780 = new_n17779 ^ new_n17776;
  assign new_n17781 = ~new_n17702 & new_n17780;
  assign new_n17782 = new_n17708 ^ new_n17690;
  assign new_n17783 = new_n17755 ^ new_n17710;
  assign new_n17784 = new_n17729 ^ new_n17690;
  assign new_n17785 = new_n17761 ^ new_n17755;
  assign new_n17786 = new_n17785 ^ new_n17774;
  assign new_n17787 = new_n17786 ^ new_n17784;
  assign new_n17788 = new_n17779 ^ new_n17760;
  assign new_n17789 = ~new_n17787 & new_n17788;
  assign new_n17790 = new_n17789 ^ new_n17763;
  assign new_n17791 = new_n17790 ^ new_n17768;
  assign new_n17792 = new_n17776 ^ new_n17760;
  assign new_n17793 = ~new_n17792 & new_n17779;
  assign new_n17794 = new_n17793 ^ new_n17760;
  assign new_n17795 = ~new_n17791 & new_n17794;
  assign new_n17796 = new_n17793 ^ new_n17779;
  assign new_n17797 = new_n17796 ^ new_n17795;
  assign new_n17798 = new_n17797 ^ new_n17783;
  assign new_n17799 = new_n17798 ^ new_n17782;
  assign new_n17800 = new_n17799 ^ new_n17686;
  assign new_n17801 = new_n17789 ^ new_n17731;
  assign new_n17802 = new_n17801 ^ new_n17750;
  assign new_n17803 = new_n17802 ^ new_n17800;
  assign new_n17804 = ~new_n17739 & ~new_n17803;
  assign new_n17805 = new_n17795 ^ new_n17787;
  assign new_n17806 = ~new_n17701 & ~new_n17805;
  assign new_n17807 = ~new_n17803 & new_n17740;
  assign new_n17808 = new_n17789 ^ new_n17776;
  assign new_n17809 = new_n17778 ^ new_n17763;
  assign new_n17810 = new_n17809 ^ new_n17808;
  assign new_n17811 = ~new_n17810 & new_n17736;
  assign new_n17812 = new_n17811 ^ new_n17807;
  assign new_n17813 = new_n17796 ^ new_n17776;
  assign new_n17814 = new_n17813 ^ new_n17775;
  assign new_n17815 = ~new_n17754 & ~new_n17814;
  assign new_n17816 = new_n17815 ^ new_n17812;
  assign new_n17817 = new_n17816 ^ new_n17806;
  assign new_n17818 = new_n17795 ^ new_n17789;
  assign new_n17819 = new_n17818 ^ new_n17759;
  assign new_n17820 = new_n17724 & new_n17819;
  assign new_n17821 = new_n17820 ^ new_n17817;
  assign new_n17822 = new_n17821 ^ new_n17804;
  assign new_n17823 = new_n17822 ^ new_n17781;
  assign new_n17824 = new_n17776 ^ new_n17729;
  assign new_n17825 = new_n17772 ^ new_n17761;
  assign new_n17826 = new_n17825 ^ new_n17799;
  assign new_n17827 = new_n17826 ^ new_n17824;
  assign new_n17828 = ~new_n17765 & new_n17827;
  assign new_n17829 = ~new_n17770 & ~new_n17791;
  assign new_n17830 = new_n17829 ^ new_n17828;
  assign new_n17831 = new_n17730 & new_n17819;
  assign new_n17832 = ~new_n17700 & new_n17780;
  assign new_n17833 = new_n17796 ^ new_n17745;
  assign new_n17834 = ~new_n17746 & ~new_n17833;
  assign new_n17835 = new_n17834 ^ new_n17832;
  assign new_n17836 = new_n17835 ^ new_n17831;
  assign new_n17837 = new_n17836 ^ new_n17830;
  assign new_n17838 = new_n17837 ^ new_n17823;
  assign new_n17839 = new_n17838 ^ new_n17680;
  assign new_n17840 = new_n15317 ^ new_n12447;
  assign new_n17841 = new_n17426 ^ new_n11990;
  assign new_n17842 = new_n17841 ^ new_n17840;
  assign new_n17843 = new_n15339 ^ new_n12509;
  assign new_n17844 = new_n17429 ^ new_n12463;
  assign new_n17845 = new_n17844 ^ new_n17843;
  assign new_n17846 = new_n17845 ^ new_n17842;
  assign new_n17847 = new_n12572 ^ new_n12540;
  assign new_n17848 = new_n17431 ^ new_n12642;
  assign new_n17849 = new_n17848 ^ new_n17847;
  assign new_n17850 = new_n17849 ^ new_n17846;
  assign new_n17851 = new_n17417 ^ new_n15331;
  assign new_n17852 = new_n17851 ^ new_n12642;
  assign new_n17853 = new_n17004 ^ new_n12409;
  assign new_n17854 = new_n17853 ^ new_n17852;
  assign new_n17855 = new_n17854 ^ new_n17850;
  assign new_n17856 = new_n17849 & new_n17855;
  assign new_n17857 = new_n17856 ^ new_n17854;
  assign new_n17858 = new_n17419 ^ new_n12642;
  assign new_n17859 = new_n15352 ^ new_n12600;
  assign new_n17860 = new_n17859 ^ new_n12560;
  assign new_n17861 = new_n17860 ^ new_n17858;
  assign new_n17862 = new_n15363 ^ new_n12258;
  assign new_n17863 = new_n17862 ^ new_n12621;
  assign new_n17864 = new_n17423 ^ new_n12642;
  assign new_n17865 = new_n17864 ^ new_n17863;
  assign new_n17866 = new_n17865 ^ new_n17861;
  assign new_n17867 = new_n17420 ^ new_n12513;
  assign new_n17868 = new_n15321 ^ new_n12641;
  assign new_n17869 = new_n17868 ^ new_n17867;
  assign new_n17870 = new_n17869 ^ new_n17854;
  assign new_n17871 = new_n17870 ^ new_n17866;
  assign new_n17872 = new_n17861 ^ new_n17854;
  assign new_n17873 = new_n15324 ^ new_n12611;
  assign new_n17874 = new_n17416 ^ new_n12590;
  assign new_n17875 = new_n17874 ^ new_n17873;
  assign new_n17876 = new_n17875 ^ new_n17869;
  assign new_n17877 = new_n17876 ^ new_n17872;
  assign new_n17878 = new_n17871 & new_n17877;
  assign new_n17879 = new_n17878 ^ new_n17845;
  assign new_n17880 = new_n17879 ^ new_n17857;
  assign new_n17881 = ~new_n17850 & ~new_n17861;
  assign new_n17882 = new_n17881 ^ new_n17861;
  assign new_n17883 = new_n17869 ^ new_n17861;
  assign new_n17884 = new_n17875 ^ new_n17866;
  assign new_n17885 = new_n17884 ^ new_n17842;
  assign new_n17886 = new_n17883 & new_n17885;
  assign new_n17887 = new_n17886 ^ new_n17882;
  assign new_n17888 = new_n17887 ^ new_n17876;
  assign new_n17889 = new_n17854 ^ new_n17842;
  assign new_n17890 = new_n17889 ^ new_n17876;
  assign new_n17891 = new_n17875 ^ new_n17854;
  assign new_n17892 = new_n17890 & new_n17891;
  assign new_n17893 = new_n17884 ^ new_n17845;
  assign new_n17894 = new_n17870 & new_n17893;
  assign new_n17895 = new_n17894 ^ new_n17892;
  assign new_n17896 = new_n17865 ^ new_n17842;
  assign new_n17897 = new_n17896 ^ new_n17895;
  assign new_n17898 = new_n17897 ^ new_n17888;
  assign new_n17899 = new_n17879 ^ new_n17871;
  assign new_n17900 = new_n17871 ^ new_n17849;
  assign new_n17901 = new_n17861 ^ new_n17850;
  assign new_n17902 = new_n17901 ^ new_n17876;
  assign new_n17903 = new_n17900 & new_n17902;
  assign new_n17904 = new_n17903 ^ new_n17895;
  assign new_n17905 = new_n17904 ^ new_n17875;
  assign new_n17906 = new_n17905 ^ new_n17899;
  assign new_n17907 = ~new_n17898 & new_n17906;
  assign new_n17908 = new_n17907 ^ new_n17880;
  assign new_n17909 = new_n17871 ^ new_n17846;
  assign new_n17910 = new_n17876 & new_n17909;
  assign new_n17911 = new_n17910 ^ new_n17894;
  assign new_n17912 = new_n17911 ^ new_n17885;
  assign new_n17913 = new_n17912 ^ new_n17908;
  assign new_n17914 = new_n17910 ^ new_n17892;
  assign new_n17915 = new_n17869 ^ new_n17850;
  assign new_n17916 = new_n17893 ^ new_n17849;
  assign new_n17917 = new_n17915 & new_n17916;
  assign new_n17918 = new_n17917 ^ new_n17881;
  assign new_n17919 = new_n17918 ^ new_n17914;
  assign new_n17920 = ~new_n17919 & new_n17913;
  assign new_n17921 = new_n17917 ^ new_n17886;
  assign new_n17922 = new_n17921 ^ new_n17869;
  assign new_n17923 = new_n17922 ^ new_n17912;
  assign new_n17924 = new_n17923 ^ new_n17920;
  assign new_n17925 = new_n17855 & new_n17924;
  assign new_n17926 = new_n17920 ^ new_n17907;
  assign new_n17927 = ~new_n17923 & ~new_n17926;
  assign new_n17928 = new_n17927 ^ new_n17920;
  assign new_n17929 = new_n17923 ^ new_n17907;
  assign new_n17930 = new_n17869 ^ new_n17842;
  assign new_n17931 = new_n17903 ^ new_n17856;
  assign new_n17932 = new_n17931 ^ new_n17914;
  assign new_n17933 = new_n17932 ^ new_n17930;
  assign new_n17934 = new_n17929 & new_n17933;
  assign new_n17935 = new_n17934 ^ new_n17880;
  assign new_n17936 = new_n17935 ^ new_n17912;
  assign new_n17937 = ~new_n17928 & new_n17936;
  assign new_n17938 = new_n17937 ^ new_n17933;
  assign new_n17939 = new_n17850 & new_n17938;
  assign new_n17940 = new_n17929 ^ new_n17928;
  assign new_n17941 = new_n17940 ^ new_n17920;
  assign new_n17942 = new_n17941 ^ new_n17919;
  assign new_n17943 = new_n17902 & new_n17942;
  assign new_n17944 = new_n17861 ^ new_n17842;
  assign new_n17945 = new_n17903 ^ new_n17882;
  assign new_n17946 = new_n17940 ^ new_n17937;
  assign new_n17947 = new_n17946 ^ new_n17945;
  assign new_n17948 = new_n17947 ^ new_n17944;
  assign new_n17949 = new_n17948 ^ new_n17854;
  assign new_n17950 = new_n17934 ^ new_n17886;
  assign new_n17951 = new_n17950 ^ new_n17879;
  assign new_n17952 = new_n17951 ^ new_n17949;
  assign new_n17953 = new_n17891 & new_n17952;
  assign new_n17954 = new_n17934 ^ new_n17920;
  assign new_n17955 = new_n17922 ^ new_n17880;
  assign new_n17956 = new_n17955 ^ new_n17954;
  assign new_n17957 = new_n17870 & new_n17956;
  assign new_n17958 = new_n17957 ^ new_n17953;
  assign new_n17959 = new_n17958 ^ new_n17943;
  assign new_n17960 = new_n17959 ^ new_n17939;
  assign new_n17961 = new_n17937 ^ new_n17934;
  assign new_n17962 = new_n17961 ^ new_n17906;
  assign new_n17963 = new_n17885 & new_n17962;
  assign new_n17964 = new_n17963 ^ new_n17960;
  assign new_n17965 = new_n17890 & new_n17952;
  assign new_n17966 = new_n17965 ^ new_n17964;
  assign new_n17967 = new_n17966 ^ new_n17925;
  assign new_n17968 = new_n17915 & new_n17936;
  assign new_n17969 = new_n17920 ^ new_n17869;
  assign new_n17970 = new_n17917 ^ new_n17856;
  assign new_n17971 = new_n17970 ^ new_n17948;
  assign new_n17972 = new_n17971 ^ new_n17969;
  assign new_n17973 = new_n17909 & new_n17972;
  assign new_n17974 = new_n17973 ^ new_n17968;
  assign new_n17975 = new_n17883 & new_n17962;
  assign new_n17976 = new_n17849 & new_n17924;
  assign new_n17977 = new_n17940 ^ new_n17898;
  assign new_n17978 = new_n17871 & new_n17977;
  assign new_n17979 = new_n17978 ^ new_n17976;
  assign new_n17980 = new_n17979 ^ new_n17975;
  assign new_n17981 = new_n17980 ^ new_n17974;
  assign new_n17982 = new_n17981 ^ new_n17967;
  assign new_n17983 = new_n11464 ^ new_n11096;
  assign new_n17984 = new_n17983 ^ new_n14870;
  assign new_n17985 = new_n17984 ^ new_n14834;
  assign new_n17986 = new_n16679 ^ new_n14716;
  assign new_n17987 = new_n17986 ^ new_n17985;
  assign new_n17988 = new_n14846 ^ new_n14742;
  assign new_n17989 = new_n11005 ^ new_n10299;
  assign new_n17990 = new_n17989 ^ new_n14695;
  assign new_n17991 = new_n17990 ^ new_n14377;
  assign new_n17992 = new_n17991 ^ new_n17988;
  assign new_n17993 = new_n14743 ^ new_n14650;
  assign new_n17994 = new_n11407 ^ new_n10687;
  assign new_n17995 = new_n17994 ^ new_n14234;
  assign new_n17996 = new_n17995 ^ new_n14865;
  assign new_n17997 = new_n17996 ^ new_n17993;
  assign new_n17998 = new_n17997 ^ new_n17992;
  assign new_n17999 = new_n11424 ^ new_n11056;
  assign new_n18000 = new_n17999 ^ new_n14880;
  assign new_n18001 = new_n15951 ^ new_n14870;
  assign new_n18002 = new_n18001 ^ new_n18000;
  assign new_n18003 = new_n18002 ^ new_n17998;
  assign new_n18004 = new_n18003 ^ new_n17987;
  assign new_n18005 = new_n16712 ^ new_n14880;
  assign new_n18006 = new_n18005 ^ new_n14870;
  assign new_n18007 = new_n11536 ^ new_n11138;
  assign new_n18008 = new_n18007 ^ new_n14782;
  assign new_n18009 = new_n18008 ^ new_n14895;
  assign new_n18010 = new_n18009 ^ new_n18006;
  assign new_n18011 = new_n18003 & new_n18010;
  assign new_n18012 = new_n18011 ^ new_n18010;
  assign new_n18013 = new_n11559 ^ new_n11181;
  assign new_n18014 = new_n18013 ^ new_n14669;
  assign new_n18015 = new_n15924 ^ new_n14869;
  assign new_n18016 = new_n18015 ^ new_n18014;
  assign new_n18017 = new_n18016 ^ new_n18010;
  assign new_n18018 = new_n14841 ^ new_n14829;
  assign new_n18019 = new_n18018 ^ new_n14815;
  assign new_n18020 = new_n11503 ^ new_n11165;
  assign new_n18021 = new_n18020 ^ new_n14870;
  assign new_n18022 = new_n18021 ^ new_n14899;
  assign new_n18023 = new_n18022 ^ new_n18019;
  assign new_n18024 = new_n18023 ^ new_n18010;
  assign new_n18025 = new_n14898 ^ new_n14820;
  assign new_n18026 = new_n18025 ^ new_n14905;
  assign new_n18027 = new_n11581 ^ new_n11210;
  assign new_n18028 = new_n18027 ^ new_n15947;
  assign new_n18029 = new_n18028 ^ new_n18026;
  assign new_n18030 = new_n18029 ^ new_n18024;
  assign new_n18031 = new_n18030 ^ new_n17992;
  assign new_n18032 = ~new_n18017 & new_n18031;
  assign new_n18033 = new_n18032 ^ new_n18012;
  assign new_n18034 = new_n18029 ^ new_n18016;
  assign new_n18035 = new_n18034 ^ new_n18033;
  assign new_n18036 = new_n18029 ^ new_n17987;
  assign new_n18037 = new_n17992 ^ new_n17987;
  assign new_n18038 = new_n18037 ^ new_n18034;
  assign new_n18039 = ~new_n18038 & new_n18036;
  assign new_n18040 = new_n18030 ^ new_n17997;
  assign new_n18041 = new_n18016 ^ new_n17987;
  assign new_n18042 = new_n18040 & new_n18041;
  assign new_n18043 = new_n18042 ^ new_n18039;
  assign new_n18044 = new_n18023 ^ new_n17992;
  assign new_n18045 = new_n18044 ^ new_n18043;
  assign new_n18046 = new_n18045 ^ new_n18035;
  assign new_n18047 = new_n18041 ^ new_n18024;
  assign new_n18048 = new_n18036 ^ new_n18017;
  assign new_n18049 = ~new_n18047 & ~new_n18048;
  assign new_n18050 = new_n18049 ^ new_n17997;
  assign new_n18051 = new_n18050 ^ new_n18047;
  assign new_n18052 = new_n18047 ^ new_n18002;
  assign new_n18053 = new_n18010 ^ new_n18003;
  assign new_n18054 = new_n18053 ^ new_n18034;
  assign new_n18055 = new_n18052 & new_n18054;
  assign new_n18056 = new_n18055 ^ new_n18042;
  assign new_n18057 = new_n18039 ^ new_n18029;
  assign new_n18058 = new_n18057 ^ new_n18056;
  assign new_n18059 = new_n18058 ^ new_n18051;
  assign new_n18060 = ~new_n18046 & new_n18059;
  assign new_n18061 = ~new_n18002 & ~new_n18004;
  assign new_n18062 = new_n18061 ^ new_n17987;
  assign new_n18063 = new_n18062 ^ new_n18050;
  assign new_n18064 = new_n18063 ^ new_n18060;
  assign new_n18065 = new_n18047 ^ new_n17998;
  assign new_n18066 = ~new_n18065 & new_n18034;
  assign new_n18067 = new_n18066 ^ new_n18042;
  assign new_n18068 = new_n18067 ^ new_n18031;
  assign new_n18069 = new_n18068 ^ new_n18064;
  assign new_n18070 = new_n18016 ^ new_n18003;
  assign new_n18071 = new_n18040 ^ new_n18002;
  assign new_n18072 = ~new_n18070 & ~new_n18071;
  assign new_n18073 = new_n18072 ^ new_n18011;
  assign new_n18074 = new_n18066 ^ new_n18039;
  assign new_n18075 = new_n18074 ^ new_n18073;
  assign new_n18076 = ~new_n18069 & ~new_n18075;
  assign new_n18077 = new_n18072 ^ new_n18032;
  assign new_n18078 = new_n18077 ^ new_n18016;
  assign new_n18079 = new_n18078 ^ new_n18068;
  assign new_n18080 = new_n18079 ^ new_n18076;
  assign new_n18081 = ~new_n18004 & new_n18080;
  assign new_n18082 = new_n18010 ^ new_n17992;
  assign new_n18083 = new_n18055 ^ new_n18012;
  assign new_n18084 = new_n18076 ^ new_n18060;
  assign new_n18085 = ~new_n18079 & ~new_n18084;
  assign new_n18086 = new_n18085 ^ new_n18076;
  assign new_n18087 = new_n18079 ^ new_n18060;
  assign new_n18088 = new_n18016 ^ new_n17992;
  assign new_n18089 = new_n18061 ^ new_n18055;
  assign new_n18090 = new_n18089 ^ new_n18074;
  assign new_n18091 = new_n18090 ^ new_n18088;
  assign new_n18092 = ~new_n18091 & new_n18087;
  assign new_n18093 = new_n18092 ^ new_n18063;
  assign new_n18094 = new_n18093 ^ new_n18068;
  assign new_n18095 = ~new_n18086 & ~new_n18094;
  assign new_n18096 = new_n18087 ^ new_n18086;
  assign new_n18097 = new_n18096 ^ new_n18095;
  assign new_n18098 = new_n18097 ^ new_n18083;
  assign new_n18099 = new_n18098 ^ new_n18082;
  assign new_n18100 = new_n18099 ^ new_n17987;
  assign new_n18101 = new_n18092 ^ new_n18032;
  assign new_n18102 = new_n18101 ^ new_n18050;
  assign new_n18103 = new_n18102 ^ new_n18100;
  assign new_n18104 = ~new_n18038 & new_n18103;
  assign new_n18105 = new_n18095 ^ new_n18092;
  assign new_n18106 = new_n18105 ^ new_n18059;
  assign new_n18107 = new_n18031 & new_n18106;
  assign new_n18108 = new_n18095 ^ new_n18091;
  assign new_n18109 = ~new_n18003 & ~new_n18108;
  assign new_n18110 = new_n18036 & new_n18103;
  assign new_n18111 = new_n18092 ^ new_n18076;
  assign new_n18112 = new_n18078 ^ new_n18063;
  assign new_n18113 = new_n18112 ^ new_n18111;
  assign new_n18114 = ~new_n18113 & new_n18041;
  assign new_n18115 = new_n18114 ^ new_n18110;
  assign new_n18116 = new_n18096 ^ new_n18076;
  assign new_n18117 = new_n18116 ^ new_n18075;
  assign new_n18118 = new_n18054 & new_n18117;
  assign new_n18119 = new_n18118 ^ new_n18115;
  assign new_n18120 = new_n18119 ^ new_n18109;
  assign new_n18121 = new_n18120 ^ new_n18107;
  assign new_n18122 = new_n18121 ^ new_n18104;
  assign new_n18123 = new_n18122 ^ new_n18081;
  assign new_n18124 = ~new_n18017 & new_n18106;
  assign new_n18125 = new_n18096 ^ new_n18046;
  assign new_n18126 = ~new_n18047 & new_n18125;
  assign new_n18127 = ~new_n18002 & new_n18080;
  assign new_n18128 = new_n18127 ^ new_n18126;
  assign new_n18129 = new_n18128 ^ new_n18124;
  assign new_n18130 = new_n18076 ^ new_n18016;
  assign new_n18131 = new_n18072 ^ new_n18061;
  assign new_n18132 = new_n18131 ^ new_n18099;
  assign new_n18133 = new_n18132 ^ new_n18130;
  assign new_n18134 = ~new_n18065 & ~new_n18133;
  assign new_n18135 = ~new_n18070 & ~new_n18094;
  assign new_n18136 = new_n18135 ^ new_n18134;
  assign new_n18137 = new_n18136 ^ new_n18129;
  assign new_n18138 = new_n18137 ^ new_n18123;
  assign new_n18139 = new_n18138 ^ new_n17982;
  assign new_n18140 = new_n17975 ^ new_n17973;
  assign new_n18141 = new_n17965 ^ new_n17939;
  assign new_n18142 = new_n17901 & new_n17938;
  assign new_n18143 = new_n17916 & new_n17936;
  assign new_n18144 = new_n18143 ^ new_n18142;
  assign new_n18145 = new_n18144 ^ new_n17958;
  assign new_n18146 = new_n18145 ^ new_n18141;
  assign new_n18147 = new_n18146 ^ new_n18140;
  assign new_n18148 = new_n15486 ^ new_n13169;
  assign new_n18149 = new_n12248 ^ new_n7966;
  assign new_n18150 = new_n18149 ^ new_n13555;
  assign new_n18151 = new_n18150 ^ new_n15490;
  assign new_n18152 = new_n18151 ^ new_n18148;
  assign new_n18153 = new_n12644 ^ new_n7938;
  assign new_n18154 = new_n18153 ^ new_n13316;
  assign new_n18155 = new_n15467 ^ new_n13710;
  assign new_n18156 = new_n18155 ^ new_n18154;
  assign new_n18157 = new_n18156 ^ new_n18152;
  assign new_n18158 = new_n15520 ^ new_n13634;
  assign new_n18159 = new_n12565 ^ new_n7788;
  assign new_n18160 = new_n18159 ^ new_n13678;
  assign new_n18161 = new_n18160 ^ new_n15490;
  assign new_n18162 = new_n18161 ^ new_n18158;
  assign new_n18163 = new_n12626 ^ new_n7823;
  assign new_n18164 = new_n18163 ^ new_n13477;
  assign new_n18165 = new_n18164 ^ new_n15490;
  assign new_n18166 = new_n15506 ^ new_n13694;
  assign new_n18167 = new_n18166 ^ new_n18165;
  assign new_n18168 = new_n18167 ^ new_n18162;
  assign new_n18169 = new_n18168 ^ new_n18157;
  assign new_n18170 = new_n12517 ^ new_n7862;
  assign new_n18171 = new_n18170 ^ new_n13718;
  assign new_n18172 = new_n15461 ^ new_n13567;
  assign new_n18173 = new_n18172 ^ new_n18171;
  assign new_n18174 = new_n12481 ^ new_n7911;
  assign new_n18175 = new_n18174 ^ new_n13588;
  assign new_n18176 = new_n15497 ^ new_n13516;
  assign new_n18177 = new_n18176 ^ new_n18175;
  assign new_n18178 = new_n18177 ^ new_n18173;
  assign new_n18179 = new_n18178 ^ new_n18169;
  assign new_n18180 = new_n12546 ^ new_n7897;
  assign new_n18181 = new_n18180 ^ new_n13646;
  assign new_n18182 = new_n15490 ^ new_n13621;
  assign new_n18183 = new_n18182 ^ new_n18181;
  assign new_n18184 = new_n18183 ^ new_n18178;
  assign new_n18185 = new_n18162 & new_n18184;
  assign new_n18186 = new_n18185 ^ new_n18162;
  assign new_n18187 = new_n12594 ^ new_n714;
  assign new_n18188 = new_n18187 ^ new_n13700;
  assign new_n18189 = new_n15476 ^ new_n13664;
  assign new_n18190 = new_n18189 ^ new_n18188;
  assign new_n18191 = new_n18190 ^ new_n18168;
  assign new_n18192 = new_n18191 ^ new_n18177;
  assign new_n18193 = new_n18162 ^ new_n18156;
  assign new_n18194 = ~new_n18193 & new_n18192;
  assign new_n18195 = new_n18194 ^ new_n18186;
  assign new_n18196 = new_n18190 ^ new_n18156;
  assign new_n18197 = new_n18196 ^ new_n18195;
  assign new_n18198 = new_n18177 ^ new_n18152;
  assign new_n18199 = new_n18198 ^ new_n18196;
  assign new_n18200 = new_n18190 ^ new_n18152;
  assign new_n18201 = ~new_n18199 & new_n18200;
  assign new_n18202 = new_n18191 ^ new_n18173;
  assign new_n18203 = new_n18157 & new_n18202;
  assign new_n18204 = new_n18203 ^ new_n18201;
  assign new_n18205 = new_n18177 ^ new_n18167;
  assign new_n18206 = new_n18205 ^ new_n18204;
  assign new_n18207 = new_n18206 ^ new_n18197;
  assign new_n18208 = new_n18162 ^ new_n18152;
  assign new_n18209 = new_n18208 ^ new_n18196;
  assign new_n18210 = ~new_n18169 & ~new_n18209;
  assign new_n18211 = new_n18210 ^ new_n18173;
  assign new_n18212 = new_n18211 ^ new_n18169;
  assign new_n18213 = new_n18183 ^ new_n18169;
  assign new_n18214 = new_n18184 ^ new_n18162;
  assign new_n18215 = new_n18214 ^ new_n18196;
  assign new_n18216 = new_n18213 & new_n18215;
  assign new_n18217 = new_n18216 ^ new_n18203;
  assign new_n18218 = new_n18201 ^ new_n18190;
  assign new_n18219 = new_n18218 ^ new_n18217;
  assign new_n18220 = new_n18219 ^ new_n18212;
  assign new_n18221 = ~new_n18207 & new_n18220;
  assign new_n18222 = new_n18184 ^ new_n18152;
  assign new_n18223 = ~new_n18183 & ~new_n18222;
  assign new_n18224 = new_n18223 ^ new_n18152;
  assign new_n18225 = new_n18224 ^ new_n18211;
  assign new_n18226 = new_n18225 ^ new_n18221;
  assign new_n18227 = ~new_n18179 & new_n18196;
  assign new_n18228 = new_n18227 ^ new_n18203;
  assign new_n18229 = new_n18228 ^ new_n18192;
  assign new_n18230 = new_n18229 ^ new_n18226;
  assign new_n18231 = new_n18227 ^ new_n18201;
  assign new_n18232 = new_n18184 ^ new_n18156;
  assign new_n18233 = new_n18202 ^ new_n18183;
  assign new_n18234 = ~new_n18232 & ~new_n18233;
  assign new_n18235 = new_n18234 ^ new_n18185;
  assign new_n18236 = new_n18235 ^ new_n18231;
  assign new_n18237 = ~new_n18230 & ~new_n18236;
  assign new_n18238 = new_n18237 ^ new_n18156;
  assign new_n18239 = new_n18234 ^ new_n18223;
  assign new_n18240 = new_n18177 ^ new_n18162;
  assign new_n18241 = new_n18216 ^ new_n18186;
  assign new_n18242 = new_n18234 ^ new_n18194;
  assign new_n18243 = new_n18242 ^ new_n18156;
  assign new_n18244 = new_n18243 ^ new_n18229;
  assign new_n18245 = new_n18244 ^ new_n18221;
  assign new_n18246 = new_n18237 ^ new_n18221;
  assign new_n18247 = ~new_n18244 & ~new_n18246;
  assign new_n18248 = new_n18247 ^ new_n18237;
  assign new_n18249 = new_n18248 ^ new_n18245;
  assign new_n18250 = new_n18177 ^ new_n18156;
  assign new_n18251 = new_n18223 ^ new_n18216;
  assign new_n18252 = new_n18251 ^ new_n18231;
  assign new_n18253 = new_n18252 ^ new_n18250;
  assign new_n18254 = ~new_n18253 & new_n18245;
  assign new_n18255 = new_n18254 ^ new_n18225;
  assign new_n18256 = new_n18255 ^ new_n18229;
  assign new_n18257 = ~new_n18248 & ~new_n18256;
  assign new_n18258 = new_n18257 ^ new_n18249;
  assign new_n18259 = new_n18258 ^ new_n18241;
  assign new_n18260 = new_n18259 ^ new_n18240;
  assign new_n18261 = new_n18260 ^ new_n18239;
  assign new_n18262 = new_n18261 ^ new_n18238;
  assign new_n18263 = ~new_n18179 & ~new_n18262;
  assign new_n18264 = new_n18257 ^ new_n18254;
  assign new_n18265 = new_n18264 ^ new_n18220;
  assign new_n18266 = ~new_n18193 & new_n18265;
  assign new_n18267 = new_n18266 ^ new_n18263;
  assign new_n18268 = new_n18257 ^ new_n18253;
  assign new_n18269 = ~new_n18184 & ~new_n18268;
  assign new_n18270 = new_n18260 ^ new_n18152;
  assign new_n18271 = new_n18254 ^ new_n18194;
  assign new_n18272 = new_n18271 ^ new_n18211;
  assign new_n18273 = new_n18272 ^ new_n18270;
  assign new_n18274 = ~new_n18199 & new_n18273;
  assign new_n18275 = new_n18274 ^ new_n18269;
  assign new_n18276 = ~new_n18268 & new_n18214;
  assign new_n18277 = ~new_n18233 & ~new_n18256;
  assign new_n18278 = new_n18277 ^ new_n18276;
  assign new_n18279 = new_n18200 & new_n18273;
  assign new_n18280 = new_n18254 ^ new_n18237;
  assign new_n18281 = new_n18243 ^ new_n18225;
  assign new_n18282 = new_n18281 ^ new_n18280;
  assign new_n18283 = ~new_n18282 & new_n18157;
  assign new_n18284 = new_n18283 ^ new_n18279;
  assign new_n18285 = new_n18284 ^ new_n18278;
  assign new_n18286 = new_n18285 ^ new_n18275;
  assign new_n18287 = new_n18286 ^ new_n18267;
  assign new_n18288 = new_n18287 ^ new_n18147;
  assign new_n18289 = new_n18288 ^ new_n18139;
  assign new_n18290 = new_n18289 ^ new_n17839;
  assign new_n18291 = new_n18134 ^ new_n18124;
  assign new_n18292 = new_n18109 ^ new_n18104;
  assign new_n18293 = ~new_n18108 & new_n18053;
  assign new_n18294 = ~new_n18071 & ~new_n18094;
  assign new_n18295 = new_n18294 ^ new_n18293;
  assign new_n18296 = new_n18295 ^ new_n18115;
  assign new_n18297 = new_n18296 ^ new_n18292;
  assign new_n18298 = new_n18297 ^ new_n18291;
  assign new_n18299 = new_n18298 ^ new_n18147;
  assign new_n18300 = new_n17980 ^ new_n17963;
  assign new_n18301 = new_n18300 ^ new_n18145;
  assign new_n18302 = new_n18244 ^ new_n18237;
  assign new_n18303 = ~new_n18183 & new_n18302;
  assign new_n18304 = new_n18249 ^ new_n18207;
  assign new_n18305 = ~new_n18169 & new_n18304;
  assign new_n18306 = new_n18305 ^ new_n18303;
  assign new_n18307 = new_n18306 ^ new_n18266;
  assign new_n18308 = new_n18192 & new_n18265;
  assign new_n18309 = new_n18308 ^ new_n18307;
  assign new_n18310 = new_n18309 ^ new_n18285;
  assign new_n18311 = new_n18310 ^ new_n18301;
  assign new_n18312 = new_n18311 ^ new_n18299;
  assign new_n18313 = new_n17541 ^ new_n14108;
  assign new_n18314 = new_n17831 ^ new_n17828;
  assign new_n18315 = new_n17806 ^ new_n17804;
  assign new_n18316 = ~new_n17753 & ~new_n17805;
  assign new_n18317 = ~new_n17771 & ~new_n17791;
  assign new_n18318 = new_n18317 ^ new_n18316;
  assign new_n18319 = new_n18318 ^ new_n17812;
  assign new_n18320 = new_n18319 ^ new_n18315;
  assign new_n18321 = new_n18320 ^ new_n18314;
  assign new_n18322 = new_n18321 ^ new_n18313;
  assign new_n18323 = ~new_n18282 & new_n18202;
  assign new_n18324 = ~new_n18209 & new_n18304;
  assign new_n18325 = new_n18324 ^ new_n18323;
  assign new_n18326 = new_n18249 ^ new_n18237;
  assign new_n18327 = new_n18326 ^ new_n18236;
  assign new_n18328 = new_n18215 & new_n18327;
  assign new_n18329 = new_n18328 ^ new_n18284;
  assign new_n18330 = new_n18329 ^ new_n18269;
  assign new_n18331 = new_n18330 ^ new_n18308;
  assign new_n18332 = new_n18331 ^ new_n18274;
  assign new_n18333 = new_n18332 ^ new_n18325;
  assign new_n18334 = new_n17893 & new_n17956;
  assign new_n18335 = new_n17877 & new_n17977;
  assign new_n18336 = new_n18335 ^ new_n18334;
  assign new_n18337 = new_n18336 ^ new_n17966;
  assign new_n18338 = new_n18337 ^ new_n18333;
  assign new_n18339 = new_n18338 ^ new_n18322;
  assign new_n18340 = new_n18339 ^ new_n18312;
  assign new_n18341 = new_n17524 ^ new_n14112;
  assign new_n18342 = ~new_n17833 & new_n17748;
  assign new_n18343 = new_n18342 ^ new_n18317;
  assign new_n18344 = ~new_n17814 & new_n17752;
  assign new_n18345 = new_n18344 ^ new_n17832;
  assign new_n18346 = new_n18345 ^ new_n17817;
  assign new_n18347 = new_n18346 ^ new_n18343;
  assign new_n18348 = new_n18347 ^ new_n18341;
  assign new_n18349 = new_n18348 ^ new_n18338;
  assign new_n18350 = ~new_n18048 & new_n18125;
  assign new_n18351 = new_n18350 ^ new_n18294;
  assign new_n18352 = new_n18052 & new_n18117;
  assign new_n18353 = new_n18352 ^ new_n18127;
  assign new_n18354 = new_n18353 ^ new_n18120;
  assign new_n18355 = new_n18354 ^ new_n18351;
  assign new_n18356 = new_n18335 ^ new_n18143;
  assign new_n18357 = new_n17900 & new_n17942;
  assign new_n18358 = new_n18357 ^ new_n17976;
  assign new_n18359 = new_n18358 ^ new_n17960;
  assign new_n18360 = new_n18359 ^ new_n18356;
  assign new_n18361 = new_n18360 ^ new_n18355;
  assign new_n18362 = ~new_n18222 & new_n18302;
  assign new_n18363 = new_n18362 ^ new_n18332;
  assign new_n18364 = ~new_n18232 & ~new_n18256;
  assign new_n18365 = new_n18364 ^ new_n18263;
  assign new_n18366 = new_n18365 ^ new_n18307;
  assign new_n18367 = new_n18366 ^ new_n18363;
  assign new_n18368 = new_n18367 ^ new_n17982;
  assign new_n18369 = new_n18368 ^ new_n18361;
  assign new_n18370 = new_n18369 ^ new_n18349;
  assign new_n18371 = new_n18370 ^ new_n18340;
  assign new_n18372 = new_n18371 ^ new_n18290;
  assign new_n18373 = new_n17563 ^ new_n14099;
  assign new_n18374 = ~new_n17810 & new_n17735;
  assign new_n18375 = new_n18374 ^ new_n17804;
  assign new_n18376 = new_n18344 ^ new_n17834;
  assign new_n18377 = new_n18376 ^ new_n18342;
  assign new_n18378 = new_n18377 ^ new_n17816;
  assign new_n18379 = new_n18378 ^ new_n18375;
  assign new_n18380 = new_n18379 ^ new_n18373;
  assign new_n18381 = ~new_n18113 & new_n18040;
  assign new_n18382 = new_n18381 ^ new_n18104;
  assign new_n18383 = new_n18352 ^ new_n18126;
  assign new_n18384 = new_n18383 ^ new_n18350;
  assign new_n18385 = new_n18384 ^ new_n18119;
  assign new_n18386 = new_n18385 ^ new_n18382;
  assign new_n18387 = new_n18334 ^ new_n17965;
  assign new_n18388 = new_n18357 ^ new_n17978;
  assign new_n18389 = new_n18388 ^ new_n18335;
  assign new_n18390 = new_n18389 ^ new_n17959;
  assign new_n18391 = new_n18390 ^ new_n18387;
  assign new_n18392 = new_n18391 ^ new_n18386;
  assign new_n18393 = new_n18323 ^ new_n18283;
  assign new_n18394 = ~new_n18262 & new_n18196;
  assign new_n18395 = new_n18394 ^ new_n18366;
  assign new_n18396 = new_n18395 ^ new_n18393;
  assign new_n18397 = new_n18334 ^ new_n17957;
  assign new_n18398 = new_n17876 & new_n17972;
  assign new_n18399 = new_n18398 ^ new_n17981;
  assign new_n18400 = new_n18399 ^ new_n18397;
  assign new_n18401 = new_n18400 ^ new_n18396;
  assign new_n18402 = new_n18401 ^ new_n18392;
  assign new_n18403 = new_n18402 ^ new_n18380;
  assign new_n18404 = new_n18403 ^ new_n18372;
  assign new_n18405 = new_n17567 ^ new_n14120;
  assign new_n18406 = new_n18374 ^ new_n18342;
  assign new_n18407 = new_n18406 ^ new_n17822;
  assign new_n18408 = new_n18407 ^ new_n18405;
  assign new_n18409 = new_n18381 ^ new_n18350;
  assign new_n18410 = new_n18409 ^ new_n18122;
  assign new_n18411 = new_n18410 ^ new_n18337;
  assign new_n18412 = new_n18323 ^ new_n18274;
  assign new_n18413 = new_n18213 & new_n18327;
  assign new_n18414 = new_n18413 ^ new_n18305;
  assign new_n18415 = new_n18414 ^ new_n18324;
  assign new_n18416 = new_n18415 ^ new_n18329;
  assign new_n18417 = new_n18416 ^ new_n18412;
  assign new_n18418 = new_n18417 ^ new_n18391;
  assign new_n18419 = new_n18418 ^ new_n18411;
  assign new_n18420 = new_n18419 ^ new_n18408;
  assign new_n18421 = new_n17572 ^ new_n14140;
  assign new_n18422 = new_n18374 ^ new_n17811;
  assign new_n18423 = new_n17733 & new_n17827;
  assign new_n18424 = new_n18423 ^ new_n17837;
  assign new_n18425 = new_n18424 ^ new_n18422;
  assign new_n18426 = new_n18425 ^ new_n18421;
  assign new_n18427 = new_n18381 ^ new_n18114;
  assign new_n18428 = ~new_n18133 & new_n18034;
  assign new_n18429 = new_n18428 ^ new_n18137;
  assign new_n18430 = new_n18429 ^ new_n18427;
  assign new_n18431 = new_n18430 ^ new_n18400;
  assign new_n18432 = new_n18389 ^ new_n17964;
  assign new_n18433 = new_n18415 ^ new_n18331;
  assign new_n18434 = new_n18433 ^ new_n18432;
  assign new_n18435 = new_n18434 ^ new_n18431;
  assign new_n18436 = new_n18435 ^ new_n18426;
  assign new_n18437 = new_n18436 ^ new_n18420;
  assign new_n18438 = new_n18384 ^ new_n18121;
  assign new_n18439 = new_n18438 ^ new_n18432;
  assign new_n18440 = new_n18324 ^ new_n18277;
  assign new_n18441 = new_n18413 ^ new_n18303;
  assign new_n18442 = new_n18441 ^ new_n18330;
  assign new_n18443 = new_n18442 ^ new_n18440;
  assign new_n18444 = new_n18443 ^ new_n18360;
  assign new_n18445 = new_n18444 ^ new_n18439;
  assign new_n18446 = new_n17575 ^ new_n14125;
  assign new_n18447 = new_n18377 ^ new_n17821;
  assign new_n18448 = new_n18447 ^ new_n18446;
  assign new_n18449 = new_n18448 ^ new_n18338;
  assign new_n18450 = new_n18449 ^ new_n18445;
  assign new_n18451 = new_n18450 ^ new_n18420;
  assign new_n18452 = new_n18451 ^ new_n18371;
  assign new_n18453 = new_n17580 ^ new_n14136;
  assign new_n18454 = new_n17836 ^ new_n17820;
  assign new_n18455 = new_n18454 ^ new_n18319;
  assign new_n18456 = new_n18455 ^ new_n18453;
  assign new_n18457 = new_n18129 ^ new_n18107;
  assign new_n18458 = new_n18457 ^ new_n18296;
  assign new_n18459 = new_n18458 ^ new_n18301;
  assign new_n18460 = new_n18459 ^ new_n18338;
  assign new_n18461 = new_n18460 ^ new_n18456;
  assign new_n18462 = new_n18461 ^ new_n18452;
  assign new_n18463 = new_n18436 ^ new_n18403;
  assign new_n18464 = new_n18463 ^ new_n18461;
  assign new_n18465 = new_n18464 ^ new_n18340;
  assign new_n18466 = new_n18420 ^ new_n18290;
  assign new_n18467 = new_n18466 ^ new_n18465;
  assign new_n18468 = new_n18462 & new_n18467;
  assign new_n18469 = new_n18464 ^ new_n18450;
  assign new_n18470 = new_n18461 & new_n18469;
  assign new_n18471 = new_n18470 ^ new_n18468;
  assign new_n18472 = new_n18463 ^ new_n18452;
  assign new_n18473 = new_n18466 & new_n18472;
  assign new_n18474 = new_n18450 ^ new_n18290;
  assign new_n18475 = new_n18450 ^ new_n18436;
  assign new_n18476 = new_n18475 ^ new_n18466;
  assign new_n18477 = new_n18474 & new_n18476;
  assign new_n18478 = new_n18477 ^ new_n18473;
  assign new_n18479 = new_n18478 ^ new_n18471;
  assign new_n18480 = new_n18479 ^ new_n18437;
  assign new_n18481 = new_n18464 ^ new_n18420;
  assign new_n18482 = new_n18461 ^ new_n18404;
  assign new_n18483 = new_n18481 & new_n18482;
  assign new_n18484 = new_n18436 ^ new_n18372;
  assign new_n18485 = new_n18420 ^ new_n18340;
  assign new_n18486 = new_n18484 & new_n18485;
  assign new_n18487 = new_n18486 ^ new_n18483;
  assign new_n18488 = new_n18487 ^ new_n18420;
  assign new_n18489 = new_n18404 & new_n18451;
  assign new_n18490 = new_n18489 ^ new_n18473;
  assign new_n18491 = new_n18490 ^ new_n18484;
  assign new_n18492 = new_n18491 ^ new_n18488;
  assign new_n18493 = ~new_n18340 & ~new_n18464;
  assign new_n18494 = new_n18493 ^ new_n18340;
  assign new_n18495 = new_n18494 ^ new_n18486;
  assign new_n18496 = new_n18495 ^ new_n18466;
  assign new_n18497 = new_n18489 ^ new_n18477;
  assign new_n18498 = new_n18436 ^ new_n18370;
  assign new_n18499 = new_n18498 ^ new_n18497;
  assign new_n18500 = new_n18499 ^ new_n18496;
  assign new_n18501 = new_n18450 ^ new_n18340;
  assign new_n18502 = new_n18501 ^ new_n18466;
  assign new_n18503 = new_n18452 & new_n18502;
  assign new_n18504 = new_n18503 ^ new_n18403;
  assign new_n18505 = new_n18504 ^ new_n18452;
  assign new_n18506 = new_n18497 ^ new_n18468;
  assign new_n18507 = new_n18506 ^ new_n18290;
  assign new_n18508 = new_n18507 ^ new_n18505;
  assign new_n18509 = ~new_n18500 & new_n18508;
  assign new_n18510 = new_n18509 ^ new_n18492;
  assign new_n18511 = new_n18480 & new_n18510;
  assign new_n18512 = new_n18470 ^ new_n18450;
  assign new_n18513 = new_n18512 ^ new_n18504;
  assign new_n18514 = new_n18513 ^ new_n18509;
  assign new_n18515 = new_n18514 ^ new_n18491;
  assign new_n18516 = new_n18493 ^ new_n18483;
  assign new_n18517 = new_n18516 ^ new_n18478;
  assign new_n18518 = ~new_n18517 & new_n18515;
  assign new_n18519 = new_n18518 ^ new_n18511;
  assign new_n18520 = new_n18513 ^ new_n18488;
  assign new_n18521 = new_n18520 ^ new_n18519;
  assign new_n18522 = new_n18404 & new_n18521;
  assign new_n18523 = new_n18518 ^ new_n18509;
  assign new_n18524 = new_n18492 & new_n18523;
  assign new_n18525 = new_n18524 ^ new_n18500;
  assign new_n18526 = ~new_n18525 & new_n18502;
  assign new_n18527 = new_n18526 ^ new_n18522;
  assign new_n18528 = new_n18436 ^ new_n18340;
  assign new_n18529 = new_n18494 ^ new_n18468;
  assign new_n18530 = new_n18513 ^ new_n18511;
  assign new_n18531 = new_n18530 ^ new_n18491;
  assign new_n18532 = new_n18524 ^ new_n18510;
  assign new_n18533 = new_n18531 & new_n18532;
  assign new_n18534 = new_n18533 ^ new_n18524;
  assign new_n18535 = new_n18534 ^ new_n18529;
  assign new_n18536 = new_n18535 ^ new_n18528;
  assign new_n18537 = new_n18536 ^ new_n18450;
  assign new_n18538 = new_n18511 ^ new_n18486;
  assign new_n18539 = new_n18538 ^ new_n18504;
  assign new_n18540 = new_n18539 ^ new_n18537;
  assign new_n18541 = ~new_n18540 & new_n18476;
  assign new_n18542 = new_n18524 ^ new_n18518;
  assign new_n18543 = new_n18542 ^ new_n18517;
  assign new_n18544 = ~new_n18543 & new_n18467;
  assign new_n18545 = ~new_n18540 & new_n18474;
  assign new_n18546 = new_n18451 & new_n18521;
  assign new_n18547 = new_n18546 ^ new_n18545;
  assign new_n18548 = new_n18547 ^ new_n18544;
  assign new_n18549 = new_n18533 ^ new_n18480;
  assign new_n18550 = new_n18464 & new_n18549;
  assign new_n18551 = new_n18550 ^ new_n18548;
  assign new_n18552 = new_n18533 ^ new_n18511;
  assign new_n18553 = new_n18552 ^ new_n18508;
  assign new_n18554 = new_n18484 & new_n18553;
  assign new_n18555 = new_n18554 ^ new_n18551;
  assign new_n18556 = new_n18555 ^ new_n18541;
  assign new_n18557 = new_n18556 ^ new_n18527;
  assign new_n18558 = new_n18557 ^ new_n17679;
  assign new_n18559 = new_n18541 ^ new_n18522;
  assign new_n18560 = ~new_n18543 & new_n18462;
  assign new_n18561 = ~new_n18525 & new_n18452;
  assign new_n18562 = new_n18561 ^ new_n18560;
  assign new_n18563 = new_n18562 ^ new_n18526;
  assign new_n18564 = new_n18563 ^ new_n18548;
  assign new_n18565 = new_n18564 ^ new_n18559;
  assign new_n18566 = new_n18565 ^ new_n18558;
  assign new_n18567 = new_n18566 ^ new_n17415;
  assign new_n18568 = new_n17376 ^ new_n17369;
  assign new_n18569 = ~new_n17307 & ~new_n18568;
  assign new_n18570 = new_n18569 ^ new_n17404;
  assign new_n18571 = new_n17390 ^ new_n17378;
  assign new_n18572 = new_n18571 ^ new_n17351;
  assign new_n18573 = ~new_n17295 & new_n18572;
  assign new_n18574 = new_n18573 ^ new_n18570;
  assign new_n18575 = ~new_n17279 & new_n18572;
  assign new_n18576 = new_n18575 ^ new_n18574;
  assign new_n18577 = new_n17364 & new_n17386;
  assign new_n18578 = new_n17390 ^ new_n17373;
  assign new_n18579 = new_n17346 & new_n18578;
  assign new_n18580 = new_n18579 ^ new_n18577;
  assign new_n18581 = new_n18580 ^ new_n17410;
  assign new_n18582 = new_n18581 ^ new_n18576;
  assign new_n18583 = new_n17406 ^ new_n17382;
  assign new_n18584 = ~new_n17309 & new_n18578;
  assign new_n18585 = new_n18584 ^ new_n17412;
  assign new_n18586 = new_n18585 ^ new_n18575;
  assign new_n18587 = new_n18586 ^ new_n17398;
  assign new_n18588 = new_n18587 ^ new_n18583;
  assign new_n18589 = new_n18588 ^ new_n18557;
  assign new_n18590 = new_n18589 ^ new_n18582;
  assign new_n18591 = new_n16342 ^ new_n16236;
  assign new_n18592 = new_n16306 ^ new_n16293;
  assign new_n18593 = new_n18592 ^ new_n16364;
  assign new_n18594 = new_n18593 ^ new_n18591;
  assign new_n18595 = ~new_n16295 & new_n18594;
  assign new_n18596 = ~new_n16308 & new_n16377;
  assign new_n18597 = new_n18596 ^ new_n18595;
  assign new_n18598 = new_n16380 ^ new_n16374;
  assign new_n18599 = ~new_n16373 & new_n16288;
  assign new_n18600 = ~new_n16305 & ~new_n16359;
  assign new_n18601 = new_n18600 ^ new_n18599;
  assign new_n18602 = new_n18601 ^ new_n16371;
  assign new_n18603 = new_n18602 ^ new_n18598;
  assign new_n18604 = new_n18603 ^ new_n18597;
  assign new_n18605 = new_n18518 ^ new_n18420;
  assign new_n18606 = new_n18483 ^ new_n18470;
  assign new_n18607 = new_n18606 ^ new_n18536;
  assign new_n18608 = new_n18607 ^ new_n18605;
  assign new_n18609 = ~new_n18608 & new_n18472;
  assign new_n18610 = new_n18485 & new_n18553;
  assign new_n18611 = new_n18610 ^ new_n18609;
  assign new_n18612 = new_n18550 ^ new_n18541;
  assign new_n18613 = new_n18465 & new_n18549;
  assign new_n18614 = new_n18482 & new_n18531;
  assign new_n18615 = new_n18614 ^ new_n18613;
  assign new_n18616 = new_n18615 ^ new_n18547;
  assign new_n18617 = new_n18616 ^ new_n18612;
  assign new_n18618 = new_n18617 ^ new_n18611;
  assign new_n18619 = new_n18618 ^ new_n18604;
  assign new_n18620 = new_n18619 ^ new_n18590;
  assign new_n18621 = new_n17638 ^ new_n17568;
  assign new_n18622 = new_n17603 ^ new_n17590;
  assign new_n18623 = new_n18622 ^ new_n17660;
  assign new_n18624 = new_n18623 ^ new_n18621;
  assign new_n18625 = ~new_n18624 & new_n17592;
  assign new_n18626 = new_n17605 & new_n17673;
  assign new_n18627 = new_n18626 ^ new_n18625;
  assign new_n18628 = new_n17676 ^ new_n17670;
  assign new_n18629 = new_n17585 & new_n17669;
  assign new_n18630 = new_n17602 & new_n17655;
  assign new_n18631 = new_n18630 ^ new_n18629;
  assign new_n18632 = new_n18631 ^ new_n17667;
  assign new_n18633 = new_n18632 ^ new_n18628;
  assign new_n18634 = new_n18633 ^ new_n18627;
  assign new_n18635 = new_n18634 ^ new_n17166;
  assign new_n18636 = new_n18518 ^ new_n18492;
  assign new_n18637 = new_n18461 & new_n18636;
  assign new_n18638 = new_n18637 ^ new_n18561;
  assign new_n18639 = new_n18638 ^ new_n18610;
  assign new_n18640 = new_n18639 ^ new_n18554;
  assign new_n18641 = new_n18640 ^ new_n18616;
  assign new_n18642 = new_n18641 ^ new_n18635;
  assign new_n18643 = new_n15269 ^ new_n15162;
  assign new_n18644 = new_n15235 ^ new_n15222;
  assign new_n18645 = new_n18644 ^ new_n15291;
  assign new_n18646 = new_n18645 ^ new_n18643;
  assign new_n18647 = ~new_n18646 & new_n15224;
  assign new_n18648 = new_n15236 & new_n15304;
  assign new_n18649 = new_n18648 ^ new_n18647;
  assign new_n18650 = new_n15307 ^ new_n15301;
  assign new_n18651 = new_n15217 & new_n15300;
  assign new_n18652 = new_n15234 & new_n15286;
  assign new_n18653 = new_n18652 ^ new_n18651;
  assign new_n18654 = new_n18653 ^ new_n15298;
  assign new_n18655 = new_n18654 ^ new_n18650;
  assign new_n18656 = new_n18655 ^ new_n18649;
  assign new_n18657 = new_n18656 ^ new_n18642;
  assign new_n18658 = new_n18657 ^ new_n18620;
  assign new_n18659 = new_n18658 ^ new_n18567;
  assign new_n18660 = new_n17638 ^ new_n17612;
  assign new_n18661 = new_n17589 & new_n18660;
  assign new_n18662 = new_n18661 ^ new_n17677;
  assign new_n18663 = new_n17601 & new_n17655;
  assign new_n18664 = new_n18663 ^ new_n18625;
  assign new_n18665 = ~new_n17646 & new_n17578;
  assign new_n18666 = new_n17581 & new_n18660;
  assign new_n18667 = new_n18666 ^ new_n18665;
  assign new_n18668 = new_n18667 ^ new_n18626;
  assign new_n18669 = new_n18668 ^ new_n18664;
  assign new_n18670 = new_n18669 ^ new_n18662;
  assign new_n18671 = new_n18670 ^ new_n16500;
  assign new_n18672 = new_n18481 & new_n18531;
  assign new_n18673 = new_n18672 ^ new_n18609;
  assign new_n18674 = new_n18673 ^ new_n18639;
  assign new_n18675 = new_n18469 & new_n18636;
  assign new_n18676 = new_n18675 ^ new_n18556;
  assign new_n18677 = new_n18676 ^ new_n18674;
  assign new_n18678 = new_n18677 ^ new_n18671;
  assign new_n18679 = new_n16342 ^ new_n16315;
  assign new_n18680 = ~new_n16292 & new_n18679;
  assign new_n18681 = new_n18680 ^ new_n16381;
  assign new_n18682 = ~new_n16304 & ~new_n16359;
  assign new_n18683 = new_n18682 ^ new_n18595;
  assign new_n18684 = ~new_n16273 & ~new_n16350;
  assign new_n18685 = ~new_n16284 & new_n18679;
  assign new_n18686 = new_n18685 ^ new_n18684;
  assign new_n18687 = new_n18686 ^ new_n18596;
  assign new_n18688 = new_n18687 ^ new_n18683;
  assign new_n18689 = new_n18688 ^ new_n18681;
  assign new_n18690 = new_n15269 ^ new_n15244;
  assign new_n18691 = new_n15221 & new_n18690;
  assign new_n18692 = new_n18691 ^ new_n15308;
  assign new_n18693 = new_n15233 & new_n15286;
  assign new_n18694 = new_n18693 ^ new_n18647;
  assign new_n18695 = ~new_n15277 & new_n15201;
  assign new_n18696 = new_n15213 & new_n18690;
  assign new_n18697 = new_n18696 ^ new_n18695;
  assign new_n18698 = new_n18697 ^ new_n18648;
  assign new_n18699 = new_n18698 ^ new_n18694;
  assign new_n18700 = new_n18699 ^ new_n18692;
  assign new_n18701 = new_n18700 ^ new_n18689;
  assign new_n18702 = new_n17369 ^ new_n17294;
  assign new_n18703 = new_n17365 ^ new_n17354;
  assign new_n18704 = new_n18703 ^ new_n17393;
  assign new_n18705 = new_n18704 ^ new_n18702;
  assign new_n18706 = ~new_n17358 & ~new_n18705;
  assign new_n18707 = new_n18706 ^ new_n18573;
  assign new_n18708 = new_n18584 ^ new_n17398;
  assign new_n18709 = new_n18708 ^ new_n18581;
  assign new_n18710 = new_n18709 ^ new_n18707;
  assign new_n18711 = new_n18710 ^ new_n18618;
  assign new_n18712 = new_n18711 ^ new_n18701;
  assign new_n18713 = new_n18712 ^ new_n18678;
  assign new_n18714 = new_n18713 ^ new_n18567;
  assign new_n18715 = new_n17666 ^ new_n17642;
  assign new_n18716 = ~new_n18624 & new_n17586;
  assign new_n18717 = new_n18716 ^ new_n18669;
  assign new_n18718 = new_n18717 ^ new_n18715;
  assign new_n18719 = new_n18718 ^ new_n17270;
  assign new_n18720 = new_n18586 ^ new_n17407;
  assign new_n18721 = new_n18563 ^ new_n18555;
  assign new_n18722 = new_n18721 ^ new_n18720;
  assign new_n18723 = new_n18722 ^ new_n18719;
  assign new_n18724 = new_n16370 ^ new_n16346;
  assign new_n18725 = new_n16289 & new_n18594;
  assign new_n18726 = new_n18725 ^ new_n18688;
  assign new_n18727 = new_n18726 ^ new_n18724;
  assign new_n18728 = new_n15297 ^ new_n15273;
  assign new_n18729 = ~new_n18646 & new_n15218;
  assign new_n18730 = new_n18729 ^ new_n18699;
  assign new_n18731 = new_n18730 ^ new_n18728;
  assign new_n18732 = new_n18731 ^ new_n18727;
  assign new_n18733 = new_n18546 ^ new_n18522;
  assign new_n18734 = ~new_n18608 & new_n18466;
  assign new_n18735 = new_n18734 ^ new_n18674;
  assign new_n18736 = new_n18735 ^ new_n18733;
  assign new_n18737 = new_n18736 ^ new_n18732;
  assign new_n18738 = new_n18737 ^ new_n18723;
  assign new_n18739 = new_n15307 ^ new_n15273;
  assign new_n18740 = ~new_n15281 & new_n15214;
  assign new_n18741 = new_n18740 ^ new_n18695;
  assign new_n18742 = new_n18741 ^ new_n15278;
  assign new_n18743 = new_n18742 ^ new_n15299;
  assign new_n18744 = new_n18743 ^ new_n18739;
  assign new_n18745 = new_n16380 ^ new_n16346;
  assign new_n18746 = ~new_n16354 & new_n16285;
  assign new_n18747 = new_n18746 ^ new_n18684;
  assign new_n18748 = new_n18747 ^ new_n16351;
  assign new_n18749 = new_n18748 ^ new_n16372;
  assign new_n18750 = new_n18749 ^ new_n18745;
  assign new_n18751 = new_n18750 ^ new_n18744;
  assign new_n18752 = new_n17408 ^ new_n17382;
  assign new_n18753 = ~new_n17313 & ~new_n18705;
  assign new_n18754 = ~new_n17363 & new_n17386;
  assign new_n18755 = new_n18754 ^ new_n18706;
  assign new_n18756 = new_n18755 ^ new_n18574;
  assign new_n18757 = new_n18756 ^ new_n18753;
  assign new_n18758 = new_n18757 ^ new_n18752;
  assign new_n18759 = new_n18758 ^ new_n18751;
  assign new_n18760 = new_n17676 ^ new_n17642;
  assign new_n18761 = ~new_n17650 & new_n17582;
  assign new_n18762 = new_n18761 ^ new_n18665;
  assign new_n18763 = new_n18762 ^ new_n17647;
  assign new_n18764 = new_n18763 ^ new_n17668;
  assign new_n18765 = new_n18764 ^ new_n18760;
  assign new_n18766 = new_n18765 ^ new_n17242;
  assign new_n18767 = new_n18766 ^ new_n18565;
  assign new_n18768 = new_n18767 ^ new_n18736;
  assign new_n18769 = new_n18768 ^ new_n18759;
  assign new_n18770 = new_n18769 ^ new_n18738;
  assign new_n18771 = new_n18763 ^ new_n17675;
  assign new_n18772 = new_n18771 ^ new_n17316;
  assign new_n18773 = new_n18748 ^ new_n16379;
  assign new_n18774 = new_n18742 ^ new_n15306;
  assign new_n18775 = new_n18774 ^ new_n18773;
  assign new_n18776 = new_n18775 ^ new_n18772;
  assign new_n18777 = new_n18776 ^ new_n18589;
  assign new_n18778 = new_n18577 ^ new_n17406;
  assign new_n18779 = new_n18569 ^ new_n17402;
  assign new_n18780 = new_n18779 ^ new_n18585;
  assign new_n18781 = new_n18780 ^ new_n18778;
  assign new_n18782 = new_n18781 ^ new_n18721;
  assign new_n18783 = new_n18614 ^ new_n18526;
  assign new_n18784 = new_n18637 ^ new_n18560;
  assign new_n18785 = new_n18784 ^ new_n18551;
  assign new_n18786 = new_n18785 ^ new_n18783;
  assign new_n18787 = new_n18786 ^ new_n18782;
  assign new_n18788 = new_n18787 ^ new_n18777;
  assign new_n18789 = new_n18788 ^ new_n18567;
  assign new_n18790 = new_n18630 ^ new_n17647;
  assign new_n18791 = new_n18761 ^ new_n18666;
  assign new_n18792 = new_n18791 ^ new_n17671;
  assign new_n18793 = new_n18792 ^ new_n18790;
  assign new_n18794 = new_n18793 ^ new_n17186;
  assign new_n18795 = new_n18794 ^ new_n18589;
  assign new_n18796 = new_n18652 ^ new_n15278;
  assign new_n18797 = new_n18740 ^ new_n18696;
  assign new_n18798 = new_n18797 ^ new_n15302;
  assign new_n18799 = new_n18798 ^ new_n18796;
  assign new_n18800 = new_n18600 ^ new_n16351;
  assign new_n18801 = new_n18746 ^ new_n18685;
  assign new_n18802 = new_n18801 ^ new_n16375;
  assign new_n18803 = new_n18802 ^ new_n18800;
  assign new_n18804 = new_n18803 ^ new_n18799;
  assign new_n18805 = new_n18804 ^ new_n18795;
  assign new_n18806 = ~new_n18568 & new_n17353;
  assign new_n18807 = new_n18806 ^ new_n18587;
  assign new_n18808 = new_n18807 ^ new_n18756;
  assign new_n18809 = new_n18808 ^ new_n18786;
  assign new_n18810 = new_n18809 ^ new_n18677;
  assign new_n18811 = new_n18810 ^ new_n18805;
  assign new_n18812 = new_n18811 ^ new_n18658;
  assign new_n18813 = new_n18812 ^ new_n18789;
  assign new_n18814 = new_n18813 ^ new_n18770;
  assign new_n18815 = ~new_n18714 & ~new_n18814;
  assign new_n18816 = new_n18812 ^ new_n18713;
  assign new_n18817 = new_n18816 ^ new_n18769;
  assign new_n18818 = ~new_n18789 & ~new_n18817;
  assign new_n18819 = new_n18818 ^ new_n18815;
  assign new_n18820 = new_n18816 ^ new_n18738;
  assign new_n18821 = new_n18820 ^ new_n18819;
  assign new_n18822 = new_n18668 ^ new_n17674;
  assign new_n18823 = new_n18822 ^ new_n18632;
  assign new_n18824 = new_n18823 ^ new_n17299;
  assign new_n18825 = new_n18698 ^ new_n15305;
  assign new_n18826 = new_n18825 ^ new_n18654;
  assign new_n18827 = new_n18826 ^ new_n18824;
  assign new_n18828 = new_n18687 ^ new_n16378;
  assign new_n18829 = new_n18828 ^ new_n18602;
  assign new_n18830 = new_n18829 ^ new_n18641;
  assign new_n18831 = new_n18830 ^ new_n18589;
  assign new_n18832 = new_n18831 ^ new_n18827;
  assign new_n18833 = new_n18832 ^ new_n18770;
  assign new_n18834 = new_n18833 ^ new_n18567;
  assign new_n18835 = new_n18832 ^ new_n18817;
  assign new_n18836 = ~new_n18834 & ~new_n18835;
  assign new_n18837 = new_n18659 & new_n18820;
  assign new_n18838 = new_n18837 ^ new_n18836;
  assign new_n18839 = new_n18838 ^ new_n18567;
  assign new_n18840 = new_n18839 ^ new_n18821;
  assign new_n18841 = new_n18833 ^ new_n18788;
  assign new_n18842 = new_n18832 & new_n18841;
  assign new_n18843 = new_n18842 ^ new_n18788;
  assign new_n18844 = new_n18788 ^ new_n18658;
  assign new_n18845 = new_n18844 ^ new_n18714;
  assign new_n18846 = new_n18813 & new_n18845;
  assign new_n18847 = new_n18846 ^ new_n18769;
  assign new_n18848 = new_n18847 ^ new_n18843;
  assign new_n18849 = new_n18847 ^ new_n18813;
  assign new_n18850 = new_n18788 ^ new_n18713;
  assign new_n18851 = new_n18788 ^ new_n18738;
  assign new_n18852 = new_n18851 ^ new_n18714;
  assign new_n18853 = new_n18850 & new_n18852;
  assign new_n18854 = new_n18853 ^ new_n18818;
  assign new_n18855 = new_n18832 ^ new_n18813;
  assign new_n18856 = new_n18833 ^ new_n18658;
  assign new_n18857 = new_n18856 ^ new_n18714;
  assign new_n18858 = new_n18855 & new_n18857;
  assign new_n18859 = new_n18858 ^ new_n18713;
  assign new_n18860 = new_n18859 ^ new_n18854;
  assign new_n18861 = new_n18860 ^ new_n18849;
  assign new_n18862 = ~new_n18658 & new_n18833;
  assign new_n18863 = new_n18862 ^ new_n18658;
  assign new_n18864 = new_n18863 ^ new_n18837;
  assign new_n18865 = new_n18864 ^ new_n18714;
  assign new_n18866 = new_n18811 ^ new_n18738;
  assign new_n18867 = new_n18866 ^ new_n18854;
  assign new_n18868 = new_n18867 ^ new_n18865;
  assign new_n18869 = ~new_n18868 & new_n18861;
  assign new_n18870 = new_n18869 ^ new_n18848;
  assign new_n18871 = new_n18870 ^ new_n18821;
  assign new_n18872 = new_n18853 ^ new_n18815;
  assign new_n18873 = new_n18862 ^ new_n18836;
  assign new_n18874 = new_n18873 ^ new_n18872;
  assign new_n18875 = ~new_n18874 & new_n18871;
  assign new_n18876 = new_n18875 ^ new_n18869;
  assign new_n18877 = ~new_n18840 & ~new_n18876;
  assign new_n18878 = new_n18877 ^ new_n18875;
  assign new_n18879 = new_n18869 ^ new_n18840;
  assign new_n18880 = new_n18738 ^ new_n18567;
  assign new_n18881 = new_n18858 ^ new_n18842;
  assign new_n18882 = new_n18881 ^ new_n18872;
  assign new_n18883 = new_n18882 ^ new_n18880;
  assign new_n18884 = new_n18879 & new_n18883;
  assign new_n18885 = new_n18884 ^ new_n18848;
  assign new_n18886 = new_n18885 ^ new_n18821;
  assign new_n18887 = ~new_n18878 & new_n18886;
  assign new_n18888 = new_n18887 ^ new_n18884;
  assign new_n18889 = new_n18888 ^ new_n18861;
  assign new_n18890 = new_n18659 & new_n18889;
  assign new_n18891 = new_n18875 ^ new_n18567;
  assign new_n18892 = new_n18842 ^ new_n18836;
  assign new_n18893 = new_n18738 ^ new_n18658;
  assign new_n18894 = new_n18863 ^ new_n18858;
  assign new_n18895 = new_n18879 ^ new_n18878;
  assign new_n18896 = new_n18895 ^ new_n18887;
  assign new_n18897 = new_n18896 ^ new_n18894;
  assign new_n18898 = new_n18897 ^ new_n18893;
  assign new_n18899 = new_n18898 ^ new_n18892;
  assign new_n18900 = new_n18899 ^ new_n18891;
  assign new_n18901 = ~new_n18814 & new_n18900;
  assign new_n18902 = new_n18901 ^ new_n18890;
  assign new_n18903 = new_n18898 ^ new_n18788;
  assign new_n18904 = new_n18884 ^ new_n18837;
  assign new_n18905 = new_n18904 ^ new_n18847;
  assign new_n18906 = new_n18905 ^ new_n18903;
  assign new_n18907 = new_n18852 & new_n18906;
  assign new_n18908 = new_n18887 ^ new_n18883;
  assign new_n18909 = ~new_n18833 & new_n18908;
  assign new_n18910 = new_n18909 ^ new_n18907;
  assign new_n18911 = ~new_n18856 & new_n18908;
  assign new_n18912 = ~new_n18835 & new_n18886;
  assign new_n18913 = new_n18912 ^ new_n18911;
  assign new_n18914 = new_n18884 ^ new_n18875;
  assign new_n18915 = new_n18848 ^ new_n18839;
  assign new_n18916 = new_n18915 ^ new_n18914;
  assign new_n18917 = ~new_n18789 & new_n18916;
  assign new_n18918 = new_n18850 & new_n18906;
  assign new_n18919 = new_n18918 ^ new_n18917;
  assign new_n18920 = new_n18919 ^ new_n18913;
  assign new_n18921 = new_n18920 ^ new_n18910;
  assign new_n18922 = new_n18921 ^ new_n18902;
  assign new_n18923 = new_n15035 ^ new_n885;
  assign new_n18924 = new_n15090 ^ new_n893;
  assign new_n18925 = new_n18924 ^ new_n18923;
  assign new_n18926 = new_n13955 ^ new_n904;
  assign new_n18927 = new_n18926 ^ new_n18925;
  assign new_n18928 = new_n15126 ^ new_n821;
  assign new_n18929 = new_n18928 ^ new_n18927;
  assign new_n18930 = new_n15206 ^ new_n857;
  assign new_n18931 = new_n15174 ^ new_n844;
  assign new_n18932 = new_n18931 ^ new_n18928;
  assign new_n18933 = new_n18932 ^ new_n18930;
  assign new_n18934 = new_n15185 ^ new_n866;
  assign new_n18935 = new_n18934 ^ new_n18933;
  assign new_n18936 = new_n18930 & new_n18935;
  assign new_n18937 = new_n18936 ^ new_n18934;
  assign new_n18938 = new_n15145 ^ new_n876;
  assign new_n18939 = new_n18938 ^ new_n18934;
  assign new_n18940 = new_n18939 ^ new_n18925;
  assign new_n18941 = new_n18934 ^ new_n18924;
  assign new_n18942 = new_n18938 ^ new_n18926;
  assign new_n18943 = new_n18942 ^ new_n18941;
  assign new_n18944 = new_n18940 & new_n18943;
  assign new_n18945 = new_n18944 ^ new_n18928;
  assign new_n18946 = new_n18945 ^ new_n18937;
  assign new_n18947 = ~new_n18924 & ~new_n18933;
  assign new_n18948 = new_n18947 ^ new_n18924;
  assign new_n18949 = new_n18931 ^ new_n18927;
  assign new_n18950 = new_n18938 ^ new_n18924;
  assign new_n18951 = new_n18949 & new_n18950;
  assign new_n18952 = new_n18951 ^ new_n18948;
  assign new_n18953 = new_n18952 ^ new_n18942;
  assign new_n18954 = new_n18929 & new_n18939;
  assign new_n18955 = new_n18934 ^ new_n18931;
  assign new_n18956 = new_n18955 ^ new_n18942;
  assign new_n18957 = new_n18934 ^ new_n18926;
  assign new_n18958 = new_n18956 & new_n18957;
  assign new_n18959 = new_n18958 ^ new_n18954;
  assign new_n18960 = new_n18931 ^ new_n18923;
  assign new_n18961 = new_n18960 ^ new_n18959;
  assign new_n18962 = new_n18961 ^ new_n18953;
  assign new_n18963 = new_n18945 ^ new_n18940;
  assign new_n18964 = new_n18940 ^ new_n18930;
  assign new_n18965 = new_n18933 ^ new_n18924;
  assign new_n18966 = new_n18965 ^ new_n18942;
  assign new_n18967 = new_n18964 & new_n18966;
  assign new_n18968 = new_n18967 ^ new_n18926;
  assign new_n18969 = new_n18968 ^ new_n18959;
  assign new_n18970 = new_n18969 ^ new_n18963;
  assign new_n18971 = ~new_n18962 & new_n18970;
  assign new_n18972 = new_n18971 ^ new_n18946;
  assign new_n18973 = new_n18940 ^ new_n18932;
  assign new_n18974 = new_n18942 & new_n18973;
  assign new_n18975 = new_n18974 ^ new_n18954;
  assign new_n18976 = new_n18975 ^ new_n18949;
  assign new_n18977 = new_n18976 ^ new_n18972;
  assign new_n18978 = new_n18938 ^ new_n18933;
  assign new_n18979 = new_n18930 ^ new_n18929;
  assign new_n18980 = new_n18978 & new_n18979;
  assign new_n18981 = new_n18980 ^ new_n18947;
  assign new_n18982 = new_n18974 ^ new_n18958;
  assign new_n18983 = new_n18982 ^ new_n18981;
  assign new_n18984 = ~new_n18983 & new_n18977;
  assign new_n18985 = new_n18938 ^ new_n18931;
  assign new_n18986 = new_n18967 ^ new_n18936;
  assign new_n18987 = new_n18986 ^ new_n18982;
  assign new_n18988 = new_n18987 ^ new_n18985;
  assign new_n18989 = new_n18980 ^ new_n18951;
  assign new_n18990 = new_n18989 ^ new_n18938;
  assign new_n18991 = new_n18990 ^ new_n18976;
  assign new_n18992 = new_n18991 ^ new_n18971;
  assign new_n18993 = new_n18988 & new_n18992;
  assign new_n18994 = new_n18993 ^ new_n18984;
  assign new_n18995 = new_n18990 ^ new_n18946;
  assign new_n18996 = new_n18995 ^ new_n18994;
  assign new_n18997 = new_n18929 & new_n18996;
  assign new_n18998 = new_n18931 ^ new_n18924;
  assign new_n18999 = new_n18967 ^ new_n18948;
  assign new_n19000 = new_n18993 ^ new_n18946;
  assign new_n19001 = new_n19000 ^ new_n18976;
  assign new_n19002 = new_n18984 ^ new_n18971;
  assign new_n19003 = new_n18991 & new_n19002;
  assign new_n19004 = new_n19003 ^ new_n18992;
  assign new_n19005 = new_n19001 & new_n19004;
  assign new_n19006 = new_n19005 ^ new_n19003;
  assign new_n19007 = new_n19006 ^ new_n18999;
  assign new_n19008 = new_n19007 ^ new_n18998;
  assign new_n19009 = new_n19008 ^ new_n18934;
  assign new_n19010 = new_n18993 ^ new_n18951;
  assign new_n19011 = new_n19010 ^ new_n18945;
  assign new_n19012 = new_n19011 ^ new_n19009;
  assign new_n19013 = ~new_n19012 & new_n18956;
  assign new_n19014 = new_n19013 ^ new_n18997;
  assign new_n19015 = new_n19003 ^ new_n18984;
  assign new_n19016 = new_n19015 ^ new_n18983;
  assign new_n19017 = ~new_n19016 & new_n18964;
  assign new_n19018 = new_n19003 ^ new_n18962;
  assign new_n19019 = ~new_n19018 & new_n18940;
  assign new_n19020 = new_n19019 ^ new_n19017;
  assign new_n19021 = ~new_n19018 & new_n18943;
  assign new_n19022 = new_n19021 ^ new_n19020;
  assign new_n19023 = ~new_n19016 & new_n18966;
  assign new_n19024 = new_n18939 & new_n18996;
  assign new_n19025 = ~new_n19012 & new_n18957;
  assign new_n19026 = new_n19025 ^ new_n19024;
  assign new_n19027 = new_n19026 ^ new_n19023;
  assign new_n19028 = new_n19027 ^ new_n19022;
  assign new_n19029 = new_n19028 ^ new_n19014;
  assign new_n19030 = new_n19029 ^ new_n16531;
  assign new_n19031 = new_n18425 ^ new_n18392;
  assign new_n19032 = new_n17241 ^ new_n10008;
  assign new_n19033 = new_n19032 ^ new_n18417;
  assign new_n19034 = new_n19033 ^ new_n18396;
  assign new_n19035 = new_n19034 ^ new_n19031;
  assign new_n19036 = new_n18321 ^ new_n18139;
  assign new_n19037 = new_n16499 ^ new_n9979;
  assign new_n19038 = new_n19037 ^ new_n18367;
  assign new_n19039 = new_n19038 ^ new_n18287;
  assign new_n19040 = new_n19039 ^ new_n19036;
  assign new_n19041 = new_n18455 ^ new_n18299;
  assign new_n19042 = new_n18407 ^ new_n18333;
  assign new_n19043 = new_n19042 ^ new_n19041;
  assign new_n19044 = new_n17165 ^ new_n9920;
  assign new_n19045 = new_n19044 ^ new_n18287;
  assign new_n19046 = new_n19045 ^ new_n18310;
  assign new_n19047 = new_n19046 ^ new_n19043;
  assign new_n19048 = new_n18443 ^ new_n18367;
  assign new_n19049 = new_n19048 ^ new_n17838;
  assign new_n19050 = new_n17185 ^ new_n9579;
  assign new_n19051 = new_n19050 ^ new_n18361;
  assign new_n19052 = new_n19051 ^ new_n19042;
  assign new_n19053 = new_n19052 ^ new_n19049;
  assign new_n19054 = new_n19053 ^ new_n19047;
  assign new_n19055 = new_n19054 ^ new_n19040;
  assign new_n19056 = new_n19055 ^ new_n19035;
  assign new_n19057 = new_n17298 ^ new_n10024;
  assign new_n19058 = new_n19057 ^ new_n18310;
  assign new_n19059 = new_n19042 ^ new_n18459;
  assign new_n19060 = new_n19059 ^ new_n19058;
  assign new_n19061 = new_n18431 ^ new_n18396;
  assign new_n19062 = new_n17269 ^ new_n10047;
  assign new_n19063 = new_n18447 ^ new_n18433;
  assign new_n19064 = new_n19063 ^ new_n19062;
  assign new_n19065 = new_n19064 ^ new_n19061;
  assign new_n19066 = new_n19065 ^ new_n19035;
  assign new_n19067 = new_n19066 ^ new_n19060;
  assign new_n19068 = new_n17315 ^ new_n10059;
  assign new_n19069 = new_n19068 ^ new_n18439;
  assign new_n19070 = new_n19069 ^ new_n19042;
  assign new_n19071 = new_n18443 ^ new_n18433;
  assign new_n19072 = new_n19071 ^ new_n18347;
  assign new_n19073 = new_n19072 ^ new_n19070;
  assign new_n19074 = new_n19073 ^ new_n19067;
  assign new_n19075 = ~new_n19060 & new_n19074;
  assign new_n19076 = new_n19075 ^ new_n19073;
  assign new_n19077 = new_n18411 ^ new_n18379;
  assign new_n19078 = new_n17290 ^ new_n10086;
  assign new_n19079 = new_n19078 ^ new_n18333;
  assign new_n19080 = new_n19079 ^ new_n18417;
  assign new_n19081 = new_n19080 ^ new_n19077;
  assign new_n19082 = new_n19081 ^ new_n19073;
  assign new_n19083 = new_n19082 ^ new_n19054;
  assign new_n19084 = new_n19081 ^ new_n19047;
  assign new_n19085 = new_n19073 ^ new_n19040;
  assign new_n19086 = new_n19085 ^ new_n19084;
  assign new_n19087 = ~new_n19083 & new_n19086;
  assign new_n19088 = new_n19087 ^ new_n19035;
  assign new_n19089 = new_n19088 ^ new_n19076;
  assign new_n19090 = ~new_n19047 & new_n19067;
  assign new_n19091 = new_n19090 ^ new_n19047;
  assign new_n19092 = new_n19065 ^ new_n19055;
  assign new_n19093 = ~new_n19092 & new_n19084;
  assign new_n19094 = new_n19093 ^ new_n19091;
  assign new_n19095 = new_n19081 ^ new_n19040;
  assign new_n19096 = new_n19095 ^ new_n19094;
  assign new_n19097 = ~new_n19056 & ~new_n19082;
  assign new_n19098 = new_n19073 ^ new_n19065;
  assign new_n19099 = new_n19098 ^ new_n19095;
  assign new_n19100 = new_n19085 & new_n19099;
  assign new_n19101 = new_n19100 ^ new_n19097;
  assign new_n19102 = new_n19065 ^ new_n19053;
  assign new_n19103 = new_n19102 ^ new_n19101;
  assign new_n19104 = new_n19103 ^ new_n19096;
  assign new_n19105 = new_n19088 ^ new_n19083;
  assign new_n19106 = new_n19083 ^ new_n19060;
  assign new_n19107 = new_n19067 ^ new_n19047;
  assign new_n19108 = new_n19107 ^ new_n19095;
  assign new_n19109 = new_n19106 & new_n19108;
  assign new_n19110 = new_n19109 ^ new_n19040;
  assign new_n19111 = new_n19110 ^ new_n19101;
  assign new_n19112 = new_n19111 ^ new_n19105;
  assign new_n19113 = new_n19104 & new_n19112;
  assign new_n19114 = new_n19113 ^ new_n19089;
  assign new_n19115 = new_n19083 ^ new_n19066;
  assign new_n19116 = ~new_n19095 & ~new_n19115;
  assign new_n19117 = new_n19116 ^ new_n19097;
  assign new_n19118 = new_n19117 ^ new_n19092;
  assign new_n19119 = new_n19118 ^ new_n19114;
  assign new_n19120 = new_n19081 ^ new_n19067;
  assign new_n19121 = new_n19060 ^ new_n19056;
  assign new_n19122 = ~new_n19120 & new_n19121;
  assign new_n19123 = new_n19122 ^ new_n19090;
  assign new_n19124 = new_n19116 ^ new_n19100;
  assign new_n19125 = new_n19124 ^ new_n19123;
  assign new_n19126 = ~new_n19125 & new_n19119;
  assign new_n19127 = new_n19081 ^ new_n19065;
  assign new_n19128 = new_n19109 ^ new_n19075;
  assign new_n19129 = new_n19128 ^ new_n19124;
  assign new_n19130 = new_n19129 ^ new_n19127;
  assign new_n19131 = new_n19122 ^ new_n19093;
  assign new_n19132 = new_n19131 ^ new_n19081;
  assign new_n19133 = new_n19132 ^ new_n19118;
  assign new_n19134 = new_n19133 ^ new_n19113;
  assign new_n19135 = ~new_n19134 & new_n19130;
  assign new_n19136 = new_n19135 ^ new_n19126;
  assign new_n19137 = new_n19132 ^ new_n19089;
  assign new_n19138 = new_n19137 ^ new_n19136;
  assign new_n19139 = ~new_n19056 & ~new_n19138;
  assign new_n19140 = new_n19065 ^ new_n19047;
  assign new_n19141 = new_n19109 ^ new_n19091;
  assign new_n19142 = new_n19135 ^ new_n19089;
  assign new_n19143 = new_n19142 ^ new_n19118;
  assign new_n19144 = new_n19126 ^ new_n19113;
  assign new_n19145 = ~new_n19133 & new_n19144;
  assign new_n19146 = new_n19145 ^ new_n19134;
  assign new_n19147 = ~new_n19146 & new_n19143;
  assign new_n19148 = new_n19147 ^ new_n19145;
  assign new_n19149 = new_n19148 ^ new_n19141;
  assign new_n19150 = new_n19149 ^ new_n19140;
  assign new_n19151 = new_n19150 ^ new_n19073;
  assign new_n19152 = new_n19135 ^ new_n19093;
  assign new_n19153 = new_n19152 ^ new_n19088;
  assign new_n19154 = new_n19153 ^ new_n19151;
  assign new_n19155 = new_n19099 & new_n19154;
  assign new_n19156 = new_n19155 ^ new_n19139;
  assign new_n19157 = new_n19145 ^ new_n19126;
  assign new_n19158 = new_n19157 ^ new_n19125;
  assign new_n19159 = ~new_n19158 & new_n19106;
  assign new_n19160 = new_n19145 ^ new_n19104;
  assign new_n19161 = ~new_n19083 & new_n19160;
  assign new_n19162 = new_n19161 ^ new_n19159;
  assign new_n19163 = new_n19086 & new_n19160;
  assign new_n19164 = new_n19163 ^ new_n19162;
  assign new_n19165 = ~new_n19158 & new_n19108;
  assign new_n19166 = ~new_n19082 & ~new_n19138;
  assign new_n19167 = new_n19085 & new_n19154;
  assign new_n19168 = new_n19167 ^ new_n19166;
  assign new_n19169 = new_n19168 ^ new_n19165;
  assign new_n19170 = new_n19169 ^ new_n19164;
  assign new_n19171 = new_n19170 ^ new_n19156;
  assign new_n19172 = new_n19171 ^ new_n19030;
  assign new_n19173 = new_n17524 ^ new_n12626;
  assign new_n19174 = new_n19173 ^ new_n1174;
  assign new_n19175 = new_n19174 ^ new_n15027;
  assign new_n19176 = new_n15159 ^ new_n15050;
  assign new_n19177 = new_n19176 ^ new_n19175;
  assign new_n19178 = new_n15066 ^ new_n12756;
  assign new_n19179 = new_n19178 ^ new_n15193;
  assign new_n19180 = new_n19179 ^ new_n19177;
  assign new_n19181 = new_n15203 ^ new_n15081;
  assign new_n19182 = new_n19181 ^ new_n15004;
  assign new_n19183 = new_n17541 ^ new_n12565;
  assign new_n19184 = new_n19183 ^ new_n1182;
  assign new_n19185 = new_n19184 ^ new_n15099;
  assign new_n19186 = new_n19185 ^ new_n19176;
  assign new_n19187 = new_n19186 ^ new_n19182;
  assign new_n19188 = new_n19187 ^ new_n19180;
  assign new_n19189 = new_n17555 ^ new_n12594;
  assign new_n19190 = new_n19189 ^ new_n1201;
  assign new_n19191 = new_n19190 ^ new_n13828;
  assign new_n19192 = new_n15076 ^ new_n15003;
  assign new_n19193 = new_n19192 ^ new_n15067;
  assign new_n19194 = new_n19193 ^ new_n19191;
  assign new_n19195 = new_n19194 ^ new_n19188;
  assign new_n19196 = new_n17563 ^ new_n12517;
  assign new_n19197 = new_n19196 ^ new_n1118;
  assign new_n19198 = new_n19197 ^ new_n15134;
  assign new_n19199 = new_n15169 ^ new_n15118;
  assign new_n19200 = new_n19199 ^ new_n15154;
  assign new_n19201 = new_n19200 ^ new_n19198;
  assign new_n19202 = new_n19201 ^ new_n19195;
  assign new_n19203 = new_n17567 ^ new_n12644;
  assign new_n19204 = new_n19203 ^ new_n1190;
  assign new_n19205 = new_n19204 ^ new_n15157;
  assign new_n19206 = new_n15153 ^ new_n15110;
  assign new_n19207 = new_n19206 ^ new_n15054;
  assign new_n19208 = new_n19207 ^ new_n19205;
  assign new_n19209 = new_n15192 ^ new_n15019;
  assign new_n19210 = new_n19209 ^ new_n15165;
  assign new_n19211 = new_n17575 ^ new_n12248;
  assign new_n19212 = new_n19211 ^ new_n1163;
  assign new_n19213 = new_n19212 ^ new_n15195;
  assign new_n19214 = new_n19213 ^ new_n19176;
  assign new_n19215 = new_n19214 ^ new_n19210;
  assign new_n19216 = new_n19215 ^ new_n19208;
  assign new_n19217 = new_n19216 ^ new_n19188;
  assign new_n19218 = new_n19215 ^ new_n19187;
  assign new_n19219 = new_n19208 ^ new_n19194;
  assign new_n19220 = new_n19219 ^ new_n19218;
  assign new_n19221 = new_n19217 & new_n19220;
  assign new_n19222 = new_n19221 ^ new_n19201;
  assign new_n19223 = new_n17580 ^ new_n12546;
  assign new_n19224 = new_n19223 ^ new_n1154;
  assign new_n19225 = new_n19224 ^ new_n15210;
  assign new_n19226 = new_n19176 ^ new_n15082;
  assign new_n19227 = new_n19226 ^ new_n19225;
  assign new_n19228 = new_n17572 ^ new_n12481;
  assign new_n19229 = new_n19228 ^ new_n1141;
  assign new_n19230 = new_n19229 ^ new_n15180;
  assign new_n19231 = new_n15197 ^ new_n15164;
  assign new_n19232 = new_n19231 ^ new_n15119;
  assign new_n19233 = new_n19232 ^ new_n19230;
  assign new_n19234 = new_n19233 ^ new_n19201;
  assign new_n19235 = ~new_n19234 & new_n19227;
  assign new_n19236 = ~new_n19227 & new_n19215;
  assign new_n19237 = new_n19236 ^ new_n19235;
  assign new_n19238 = new_n19237 ^ new_n19222;
  assign new_n19239 = new_n19234 ^ new_n19227;
  assign new_n19240 = ~new_n19187 & ~new_n19239;
  assign new_n19241 = new_n19240 ^ new_n19187;
  assign new_n19242 = new_n19233 ^ new_n19195;
  assign new_n19243 = new_n19208 ^ new_n19187;
  assign new_n19244 = new_n19242 & new_n19243;
  assign new_n19245 = new_n19244 ^ new_n19241;
  assign new_n19246 = new_n19245 ^ new_n19219;
  assign new_n19247 = new_n19202 & new_n19216;
  assign new_n19248 = new_n19233 ^ new_n19215;
  assign new_n19249 = new_n19248 ^ new_n19219;
  assign new_n19250 = new_n19215 ^ new_n19194;
  assign new_n19251 = new_n19249 & new_n19250;
  assign new_n19252 = new_n19251 ^ new_n19247;
  assign new_n19253 = new_n19233 ^ new_n19180;
  assign new_n19254 = new_n19253 ^ new_n19252;
  assign new_n19255 = new_n19254 ^ new_n19246;
  assign new_n19256 = new_n19222 ^ new_n19217;
  assign new_n19257 = new_n19239 ^ new_n19187;
  assign new_n19258 = new_n19257 ^ new_n19219;
  assign new_n19259 = new_n19227 ^ new_n19217;
  assign new_n19260 = new_n19258 & new_n19259;
  assign new_n19261 = new_n19260 ^ new_n19247;
  assign new_n19262 = new_n19251 ^ new_n19194;
  assign new_n19263 = new_n19262 ^ new_n19261;
  assign new_n19264 = new_n19263 ^ new_n19256;
  assign new_n19265 = ~new_n19255 & new_n19264;
  assign new_n19266 = new_n19265 ^ new_n19238;
  assign new_n19267 = new_n19234 ^ new_n19217;
  assign new_n19268 = new_n19219 & new_n19267;
  assign new_n19269 = new_n19268 ^ new_n19247;
  assign new_n19270 = new_n19269 ^ new_n19242;
  assign new_n19271 = new_n19270 ^ new_n19266;
  assign new_n19272 = new_n19239 ^ new_n19208;
  assign new_n19273 = new_n19227 ^ new_n19202;
  assign new_n19274 = new_n19272 & new_n19273;
  assign new_n19275 = new_n19274 ^ new_n19240;
  assign new_n19276 = new_n19268 ^ new_n19251;
  assign new_n19277 = new_n19276 ^ new_n19275;
  assign new_n19278 = ~new_n19277 & new_n19271;
  assign new_n19279 = new_n19233 ^ new_n19208;
  assign new_n19280 = new_n19237 ^ new_n19215;
  assign new_n19281 = new_n19280 ^ new_n19260;
  assign new_n19282 = new_n19281 ^ new_n19276;
  assign new_n19283 = new_n19282 ^ new_n19279;
  assign new_n19284 = new_n19274 ^ new_n19244;
  assign new_n19285 = new_n19284 ^ new_n19208;
  assign new_n19286 = new_n19285 ^ new_n19270;
  assign new_n19287 = new_n19286 ^ new_n19265;
  assign new_n19288 = new_n19283 & new_n19287;
  assign new_n19289 = new_n19288 ^ new_n19278;
  assign new_n19290 = new_n19285 ^ new_n19238;
  assign new_n19291 = new_n19290 ^ new_n19289;
  assign new_n19292 = new_n19202 & new_n19291;
  assign new_n19293 = new_n19216 & new_n19291;
  assign new_n19294 = new_n19293 ^ new_n19292;
  assign new_n19295 = new_n19278 ^ new_n19208;
  assign new_n19296 = new_n19280 ^ new_n19274;
  assign new_n19297 = new_n19233 ^ new_n19187;
  assign new_n19298 = new_n19260 ^ new_n19241;
  assign new_n19299 = new_n19288 ^ new_n19238;
  assign new_n19300 = new_n19299 ^ new_n19270;
  assign new_n19301 = new_n19278 ^ new_n19265;
  assign new_n19302 = new_n19286 & new_n19301;
  assign new_n19303 = new_n19302 ^ new_n19287;
  assign new_n19304 = new_n19300 & new_n19303;
  assign new_n19305 = new_n19304 ^ new_n19302;
  assign new_n19306 = new_n19305 ^ new_n19298;
  assign new_n19307 = new_n19306 ^ new_n19297;
  assign new_n19308 = new_n19307 ^ new_n19296;
  assign new_n19309 = new_n19308 ^ new_n19295;
  assign new_n19310 = ~new_n19309 & new_n19219;
  assign new_n19311 = new_n19304 ^ new_n19288;
  assign new_n19312 = new_n19311 ^ new_n19264;
  assign new_n19313 = new_n19243 & new_n19312;
  assign new_n19314 = new_n19302 ^ new_n19255;
  assign new_n19315 = ~new_n19314 & new_n19217;
  assign new_n19316 = new_n19286 ^ new_n19278;
  assign new_n19317 = new_n19227 & new_n19316;
  assign new_n19318 = new_n19317 ^ new_n19315;
  assign new_n19319 = new_n19318 ^ new_n19313;
  assign new_n19320 = ~new_n19309 & new_n19267;
  assign new_n19321 = new_n19272 & new_n19300;
  assign new_n19322 = new_n19321 ^ new_n19320;
  assign new_n19323 = new_n19322 ^ new_n19319;
  assign new_n19324 = new_n19323 ^ new_n19310;
  assign new_n19325 = new_n19324 ^ new_n19294;
  assign new_n19326 = new_n16156 ^ new_n15921;
  assign new_n19327 = new_n18923 ^ new_n16169;
  assign new_n19328 = new_n19327 ^ new_n19326;
  assign new_n19329 = new_n16226 ^ new_n16101;
  assign new_n19330 = new_n19329 ^ new_n16269;
  assign new_n19331 = new_n19330 ^ new_n19328;
  assign new_n19332 = new_n19329 ^ new_n15616;
  assign new_n19333 = new_n16276 ^ new_n16112;
  assign new_n19334 = new_n18924 ^ new_n16140;
  assign new_n19335 = new_n19334 ^ new_n19333;
  assign new_n19336 = new_n19335 ^ new_n19332;
  assign new_n19337 = new_n19336 ^ new_n19331;
  assign new_n19338 = new_n18926 ^ new_n16082;
  assign new_n19339 = new_n16122 ^ new_n15615;
  assign new_n19340 = new_n19339 ^ new_n16157;
  assign new_n19341 = new_n19340 ^ new_n19338;
  assign new_n19342 = new_n19341 ^ new_n19337;
  assign new_n19343 = new_n16244 ^ new_n16197;
  assign new_n19344 = new_n19343 ^ new_n16224;
  assign new_n19345 = new_n18928 ^ new_n16186;
  assign new_n19346 = new_n19345 ^ new_n16203;
  assign new_n19347 = new_n19346 ^ new_n19344;
  assign new_n19348 = new_n19347 ^ new_n19342;
  assign new_n19349 = new_n18930 ^ new_n16282;
  assign new_n19350 = new_n19329 ^ new_n16113;
  assign new_n19351 = new_n19350 ^ new_n19349;
  assign new_n19352 = new_n16268 ^ new_n16175;
  assign new_n19353 = new_n19352 ^ new_n18934;
  assign new_n19354 = new_n19353 ^ new_n19329;
  assign new_n19355 = new_n16258 ^ new_n16249;
  assign new_n19356 = new_n19355 ^ new_n19354;
  assign new_n19357 = new_n16259 ^ new_n16247;
  assign new_n19358 = new_n19357 ^ new_n16197;
  assign new_n19359 = new_n18931 ^ new_n16240;
  assign new_n19360 = new_n19359 ^ new_n16215;
  assign new_n19361 = new_n19360 ^ new_n19358;
  assign new_n19362 = new_n19361 ^ new_n19347;
  assign new_n19363 = new_n19362 ^ new_n19351;
  assign new_n19364 = new_n19363 ^ new_n19356;
  assign new_n19365 = ~new_n19351 & ~new_n19364;
  assign new_n19366 = new_n19365 ^ new_n19356;
  assign new_n19367 = new_n16224 ^ new_n16192;
  assign new_n19368 = new_n19367 ^ new_n18938;
  assign new_n19369 = new_n16228 ^ new_n16088;
  assign new_n19370 = new_n19369 ^ new_n16101;
  assign new_n19371 = new_n19370 ^ new_n19368;
  assign new_n19372 = new_n19371 ^ new_n19356;
  assign new_n19373 = new_n19372 ^ new_n19337;
  assign new_n19374 = new_n19356 ^ new_n19336;
  assign new_n19375 = new_n19371 ^ new_n19341;
  assign new_n19376 = new_n19375 ^ new_n19374;
  assign new_n19377 = ~new_n19373 & ~new_n19376;
  assign new_n19378 = new_n19377 ^ new_n19347;
  assign new_n19379 = new_n19378 ^ new_n19366;
  assign new_n19380 = new_n19336 & new_n19363;
  assign new_n19381 = new_n19380 ^ new_n19336;
  assign new_n19382 = new_n19361 ^ new_n19342;
  assign new_n19383 = new_n19371 ^ new_n19336;
  assign new_n19384 = ~new_n19383 & new_n19382;
  assign new_n19385 = new_n19384 ^ new_n19381;
  assign new_n19386 = new_n19385 ^ new_n19375;
  assign new_n19387 = new_n19348 & new_n19372;
  assign new_n19388 = new_n19361 ^ new_n19356;
  assign new_n19389 = new_n19388 ^ new_n19375;
  assign new_n19390 = new_n19356 ^ new_n19341;
  assign new_n19391 = ~new_n19389 & new_n19390;
  assign new_n19392 = new_n19391 ^ new_n19387;
  assign new_n19393 = new_n19361 ^ new_n19331;
  assign new_n19394 = new_n19393 ^ new_n19392;
  assign new_n19395 = new_n19394 ^ new_n19386;
  assign new_n19396 = new_n19378 ^ new_n19373;
  assign new_n19397 = new_n19363 ^ new_n19336;
  assign new_n19398 = new_n19397 ^ new_n19375;
  assign new_n19399 = new_n19373 ^ new_n19351;
  assign new_n19400 = new_n19398 & new_n19399;
  assign new_n19401 = new_n19400 ^ new_n19392;
  assign new_n19402 = new_n19401 ^ new_n19341;
  assign new_n19403 = new_n19402 ^ new_n19396;
  assign new_n19404 = ~new_n19395 & new_n19403;
  assign new_n19405 = new_n19404 ^ new_n19379;
  assign new_n19406 = new_n19373 ^ new_n19362;
  assign new_n19407 = ~new_n19406 & new_n19375;
  assign new_n19408 = new_n19407 ^ new_n19387;
  assign new_n19409 = new_n19408 ^ new_n19382;
  assign new_n19410 = new_n19409 ^ new_n19405;
  assign new_n19411 = new_n19371 ^ new_n19363;
  assign new_n19412 = new_n19351 ^ new_n19348;
  assign new_n19413 = ~new_n19411 & ~new_n19412;
  assign new_n19414 = new_n19413 ^ new_n19380;
  assign new_n19415 = new_n19407 ^ new_n19391;
  assign new_n19416 = new_n19415 ^ new_n19414;
  assign new_n19417 = ~new_n19410 & ~new_n19416;
  assign new_n19418 = new_n19371 ^ new_n19361;
  assign new_n19419 = new_n19400 ^ new_n19365;
  assign new_n19420 = new_n19419 ^ new_n19415;
  assign new_n19421 = new_n19420 ^ new_n19418;
  assign new_n19422 = new_n19413 ^ new_n19384;
  assign new_n19423 = new_n19422 ^ new_n19371;
  assign new_n19424 = new_n19423 ^ new_n19409;
  assign new_n19425 = new_n19424 ^ new_n19404;
  assign new_n19426 = ~new_n19421 & new_n19425;
  assign new_n19427 = new_n19426 ^ new_n19417;
  assign new_n19428 = new_n19423 ^ new_n19379;
  assign new_n19429 = new_n19428 ^ new_n19427;
  assign new_n19430 = ~new_n19429 & new_n19348;
  assign new_n19431 = ~new_n19429 & new_n19372;
  assign new_n19432 = new_n19431 ^ new_n19430;
  assign new_n19433 = new_n19417 ^ new_n19371;
  assign new_n19434 = new_n19413 ^ new_n19365;
  assign new_n19435 = new_n19361 ^ new_n19336;
  assign new_n19436 = new_n19400 ^ new_n19381;
  assign new_n19437 = new_n19426 ^ new_n19379;
  assign new_n19438 = new_n19437 ^ new_n19409;
  assign new_n19439 = new_n19417 ^ new_n19404;
  assign new_n19440 = new_n19424 & new_n19439;
  assign new_n19441 = new_n19440 ^ new_n19425;
  assign new_n19442 = ~new_n19438 & new_n19441;
  assign new_n19443 = new_n19442 ^ new_n19440;
  assign new_n19444 = new_n19443 ^ new_n19436;
  assign new_n19445 = new_n19444 ^ new_n19435;
  assign new_n19446 = new_n19445 ^ new_n19434;
  assign new_n19447 = new_n19446 ^ new_n19433;
  assign new_n19448 = new_n19375 & new_n19447;
  assign new_n19449 = ~new_n19406 & new_n19447;
  assign new_n19450 = ~new_n19411 & ~new_n19438;
  assign new_n19451 = new_n19450 ^ new_n19449;
  assign new_n19452 = new_n19442 ^ new_n19426;
  assign new_n19453 = new_n19452 ^ new_n19403;
  assign new_n19454 = ~new_n19383 & new_n19453;
  assign new_n19455 = new_n19440 ^ new_n19395;
  assign new_n19456 = ~new_n19373 & ~new_n19455;
  assign new_n19457 = new_n19424 ^ new_n19417;
  assign new_n19458 = ~new_n19351 & new_n19457;
  assign new_n19459 = new_n19458 ^ new_n19456;
  assign new_n19460 = new_n19459 ^ new_n19454;
  assign new_n19461 = new_n19460 ^ new_n19451;
  assign new_n19462 = new_n19461 ^ new_n19448;
  assign new_n19463 = new_n19462 ^ new_n19432;
  assign new_n19464 = new_n19463 ^ new_n19325;
  assign new_n19465 = new_n17263 ^ new_n17234;
  assign new_n19466 = new_n19465 ^ new_n17287;
  assign new_n19467 = new_n17994 ^ new_n16209;
  assign new_n19468 = new_n19467 ^ new_n17247;
  assign new_n19469 = new_n19468 ^ new_n17223;
  assign new_n19470 = new_n19469 ^ new_n19466;
  assign new_n19471 = new_n17207 ^ new_n16967;
  assign new_n19472 = new_n19471 ^ new_n16654;
  assign new_n19473 = new_n17155 ^ new_n16809;
  assign new_n19474 = new_n18027 ^ new_n15732;
  assign new_n19475 = new_n19474 ^ new_n19473;
  assign new_n19476 = new_n19475 ^ new_n19472;
  assign new_n19477 = new_n17325 ^ new_n17199;
  assign new_n19478 = new_n19477 ^ new_n17212;
  assign new_n19479 = new_n18020 ^ new_n16148;
  assign new_n19480 = new_n17281 ^ new_n17138;
  assign new_n19481 = new_n19480 ^ new_n19479;
  assign new_n19482 = new_n17207 ^ new_n17118;
  assign new_n19483 = new_n19482 ^ new_n19481;
  assign new_n19484 = new_n19483 ^ new_n19478;
  assign new_n19485 = new_n17146 ^ new_n16810;
  assign new_n19486 = new_n19485 ^ new_n19480;
  assign new_n19487 = new_n18007 ^ new_n16130;
  assign new_n19488 = new_n19487 ^ new_n17304;
  assign new_n19489 = new_n19488 ^ new_n17177;
  assign new_n19490 = new_n19489 ^ new_n19486;
  assign new_n19491 = new_n19490 ^ new_n19484;
  assign new_n19492 = new_n19491 ^ new_n19476;
  assign new_n19493 = new_n19492 ^ new_n19470;
  assign new_n19494 = new_n17999 ^ new_n16278;
  assign new_n19495 = new_n19494 ^ new_n17146;
  assign new_n19496 = new_n17301 ^ new_n17168;
  assign new_n19497 = new_n19496 ^ new_n19480;
  assign new_n19498 = new_n19497 ^ new_n19495;
  assign new_n19499 = new_n17317 ^ new_n17274;
  assign new_n19500 = new_n19499 ^ new_n17234;
  assign new_n19501 = new_n17989 ^ new_n16253;
  assign new_n19502 = new_n19501 ^ new_n17252;
  assign new_n19503 = new_n19502 ^ new_n17259;
  assign new_n19504 = new_n19503 ^ new_n19500;
  assign new_n19505 = new_n19504 ^ new_n19470;
  assign new_n19506 = new_n19505 ^ new_n19498;
  assign new_n19507 = new_n17983 ^ new_n16262;
  assign new_n19508 = new_n19507 ^ new_n19480;
  assign new_n19509 = new_n17325 ^ new_n17193;
  assign new_n19510 = new_n19509 ^ new_n19508;
  assign new_n19511 = new_n17318 ^ new_n17276;
  assign new_n19512 = new_n19511 ^ new_n19510;
  assign new_n19513 = new_n19512 ^ new_n19506;
  assign new_n19514 = new_n19498 & new_n19513;
  assign new_n19515 = new_n19514 ^ new_n19512;
  assign new_n19516 = new_n18013 ^ new_n16232;
  assign new_n19517 = new_n17287 ^ new_n17229;
  assign new_n19518 = new_n19517 ^ new_n19516;
  assign new_n19519 = new_n17283 ^ new_n17125;
  assign new_n19520 = new_n19519 ^ new_n17138;
  assign new_n19521 = new_n19520 ^ new_n19518;
  assign new_n19522 = new_n19521 ^ new_n19512;
  assign new_n19523 = new_n19522 ^ new_n19491;
  assign new_n19524 = new_n19521 ^ new_n19490;
  assign new_n19525 = new_n19512 ^ new_n19476;
  assign new_n19526 = new_n19525 ^ new_n19524;
  assign new_n19527 = new_n19523 & new_n19526;
  assign new_n19528 = new_n19527 ^ new_n19470;
  assign new_n19529 = new_n19528 ^ new_n19515;
  assign new_n19530 = ~new_n19490 & ~new_n19506;
  assign new_n19531 = new_n19530 ^ new_n19490;
  assign new_n19532 = new_n19504 ^ new_n19492;
  assign new_n19533 = new_n19524 & new_n19532;
  assign new_n19534 = new_n19533 ^ new_n19531;
  assign new_n19535 = new_n19521 ^ new_n19476;
  assign new_n19536 = new_n19535 ^ new_n19534;
  assign new_n19537 = new_n19493 & new_n19522;
  assign new_n19538 = new_n19512 ^ new_n19504;
  assign new_n19539 = new_n19538 ^ new_n19535;
  assign new_n19540 = new_n19525 & new_n19539;
  assign new_n19541 = new_n19540 ^ new_n19537;
  assign new_n19542 = new_n19504 ^ new_n19484;
  assign new_n19543 = new_n19542 ^ new_n19541;
  assign new_n19544 = new_n19543 ^ new_n19536;
  assign new_n19545 = new_n19528 ^ new_n19523;
  assign new_n19546 = new_n19523 ^ new_n19498;
  assign new_n19547 = new_n19506 ^ new_n19490;
  assign new_n19548 = new_n19547 ^ new_n19535;
  assign new_n19549 = new_n19546 & new_n19548;
  assign new_n19550 = new_n19549 ^ new_n19537;
  assign new_n19551 = new_n19540 ^ new_n19476;
  assign new_n19552 = new_n19551 ^ new_n19550;
  assign new_n19553 = new_n19552 ^ new_n19545;
  assign new_n19554 = ~new_n19544 & new_n19553;
  assign new_n19555 = new_n19554 ^ new_n19529;
  assign new_n19556 = new_n19523 ^ new_n19505;
  assign new_n19557 = new_n19535 & new_n19556;
  assign new_n19558 = new_n19557 ^ new_n19537;
  assign new_n19559 = new_n19558 ^ new_n19532;
  assign new_n19560 = new_n19559 ^ new_n19555;
  assign new_n19561 = new_n19521 ^ new_n19506;
  assign new_n19562 = new_n19498 ^ new_n19493;
  assign new_n19563 = new_n19561 & new_n19562;
  assign new_n19564 = new_n19563 ^ new_n19530;
  assign new_n19565 = new_n19557 ^ new_n19540;
  assign new_n19566 = new_n19565 ^ new_n19564;
  assign new_n19567 = ~new_n19566 & new_n19560;
  assign new_n19568 = new_n19521 ^ new_n19504;
  assign new_n19569 = new_n19549 ^ new_n19514;
  assign new_n19570 = new_n19569 ^ new_n19565;
  assign new_n19571 = new_n19570 ^ new_n19568;
  assign new_n19572 = new_n19563 ^ new_n19533;
  assign new_n19573 = new_n19572 ^ new_n19521;
  assign new_n19574 = new_n19573 ^ new_n19559;
  assign new_n19575 = new_n19574 ^ new_n19554;
  assign new_n19576 = new_n19571 & new_n19575;
  assign new_n19577 = new_n19576 ^ new_n19567;
  assign new_n19578 = new_n19573 ^ new_n19529;
  assign new_n19579 = new_n19578 ^ new_n19577;
  assign new_n19580 = new_n19493 & new_n19579;
  assign new_n19581 = new_n19504 ^ new_n19490;
  assign new_n19582 = new_n19549 ^ new_n19531;
  assign new_n19583 = new_n19576 ^ new_n19529;
  assign new_n19584 = new_n19583 ^ new_n19559;
  assign new_n19585 = new_n19567 ^ new_n19554;
  assign new_n19586 = new_n19574 & new_n19585;
  assign new_n19587 = new_n19586 ^ new_n19575;
  assign new_n19588 = new_n19584 & new_n19587;
  assign new_n19589 = new_n19588 ^ new_n19586;
  assign new_n19590 = new_n19589 ^ new_n19582;
  assign new_n19591 = new_n19590 ^ new_n19581;
  assign new_n19592 = new_n19591 ^ new_n19512;
  assign new_n19593 = new_n19576 ^ new_n19533;
  assign new_n19594 = new_n19593 ^ new_n19528;
  assign new_n19595 = new_n19594 ^ new_n19592;
  assign new_n19596 = ~new_n19595 & new_n19539;
  assign new_n19597 = new_n19596 ^ new_n19580;
  assign new_n19598 = new_n19586 ^ new_n19567;
  assign new_n19599 = new_n19598 ^ new_n19566;
  assign new_n19600 = ~new_n19599 & new_n19546;
  assign new_n19601 = new_n19586 ^ new_n19544;
  assign new_n19602 = ~new_n19601 & new_n19523;
  assign new_n19603 = new_n19602 ^ new_n19600;
  assign new_n19604 = ~new_n19601 & new_n19526;
  assign new_n19605 = new_n19604 ^ new_n19603;
  assign new_n19606 = ~new_n19599 & new_n19548;
  assign new_n19607 = new_n19522 & new_n19579;
  assign new_n19608 = ~new_n19595 & new_n19525;
  assign new_n19609 = new_n19608 ^ new_n19607;
  assign new_n19610 = new_n19609 ^ new_n19606;
  assign new_n19611 = new_n19610 ^ new_n19605;
  assign new_n19612 = new_n19611 ^ new_n19597;
  assign new_n19613 = new_n19445 ^ new_n19356;
  assign new_n19614 = new_n19426 ^ new_n19384;
  assign new_n19615 = new_n19614 ^ new_n19378;
  assign new_n19616 = new_n19615 ^ new_n19613;
  assign new_n19617 = ~new_n19389 & ~new_n19616;
  assign new_n19618 = new_n19617 ^ new_n19430;
  assign new_n19619 = new_n19440 ^ new_n19417;
  assign new_n19620 = new_n19619 ^ new_n19416;
  assign new_n19621 = ~new_n19620 & new_n19399;
  assign new_n19622 = new_n19621 ^ new_n19456;
  assign new_n19623 = ~new_n19376 & ~new_n19455;
  assign new_n19624 = new_n19623 ^ new_n19622;
  assign new_n19625 = ~new_n19620 & new_n19398;
  assign new_n19626 = ~new_n19616 & new_n19390;
  assign new_n19627 = new_n19626 ^ new_n19431;
  assign new_n19628 = new_n19627 ^ new_n19625;
  assign new_n19629 = new_n19628 ^ new_n19624;
  assign new_n19630 = new_n19629 ^ new_n19618;
  assign new_n19631 = new_n19630 ^ new_n19612;
  assign new_n19632 = new_n19631 ^ new_n19464;
  assign new_n19633 = new_n19632 ^ new_n19172;
  assign new_n19634 = new_n19024 ^ new_n18997;
  assign new_n19635 = new_n18984 ^ new_n18938;
  assign new_n19636 = new_n18980 ^ new_n18936;
  assign new_n19637 = new_n19636 ^ new_n19008;
  assign new_n19638 = new_n19637 ^ new_n19635;
  assign new_n19639 = ~new_n19638 & new_n18942;
  assign new_n19640 = new_n18978 & new_n19001;
  assign new_n19641 = ~new_n19638 & new_n18973;
  assign new_n19642 = new_n19641 ^ new_n19640;
  assign new_n19643 = new_n19005 ^ new_n18993;
  assign new_n19644 = new_n19643 ^ new_n18970;
  assign new_n19645 = new_n18950 & new_n19644;
  assign new_n19646 = new_n18991 ^ new_n18984;
  assign new_n19647 = new_n18930 & new_n19646;
  assign new_n19648 = new_n19647 ^ new_n19019;
  assign new_n19649 = new_n19648 ^ new_n19645;
  assign new_n19650 = new_n19649 ^ new_n19642;
  assign new_n19651 = new_n19650 ^ new_n19639;
  assign new_n19652 = new_n19651 ^ new_n19634;
  assign new_n19653 = new_n19652 ^ new_n16540;
  assign new_n19654 = new_n19166 ^ new_n19139;
  assign new_n19655 = new_n19126 ^ new_n19081;
  assign new_n19656 = new_n19122 ^ new_n19075;
  assign new_n19657 = new_n19656 ^ new_n19150;
  assign new_n19658 = new_n19657 ^ new_n19655;
  assign new_n19659 = ~new_n19095 & ~new_n19658;
  assign new_n19660 = ~new_n19120 & new_n19143;
  assign new_n19661 = ~new_n19115 & ~new_n19658;
  assign new_n19662 = new_n19661 ^ new_n19660;
  assign new_n19663 = new_n19147 ^ new_n19135;
  assign new_n19664 = new_n19663 ^ new_n19112;
  assign new_n19665 = new_n19084 & new_n19664;
  assign new_n19666 = new_n19133 ^ new_n19126;
  assign new_n19667 = ~new_n19060 & ~new_n19666;
  assign new_n19668 = new_n19667 ^ new_n19161;
  assign new_n19669 = new_n19668 ^ new_n19665;
  assign new_n19670 = new_n19669 ^ new_n19662;
  assign new_n19671 = new_n19670 ^ new_n19659;
  assign new_n19672 = new_n19671 ^ new_n19654;
  assign new_n19673 = new_n19672 ^ new_n19653;
  assign new_n19674 = new_n19302 ^ new_n19278;
  assign new_n19675 = new_n19674 ^ new_n19277;
  assign new_n19676 = ~new_n19675 & new_n19259;
  assign new_n19677 = new_n19676 ^ new_n19315;
  assign new_n19678 = ~new_n19314 & new_n19220;
  assign new_n19679 = new_n19678 ^ new_n19677;
  assign new_n19680 = new_n19307 ^ new_n19215;
  assign new_n19681 = new_n19288 ^ new_n19244;
  assign new_n19682 = new_n19681 ^ new_n19222;
  assign new_n19683 = new_n19682 ^ new_n19680;
  assign new_n19684 = ~new_n19683 & new_n19250;
  assign new_n19685 = new_n19684 ^ new_n19293;
  assign new_n19686 = ~new_n19675 & new_n19258;
  assign new_n19687 = new_n19686 ^ new_n19685;
  assign new_n19688 = new_n19304 ^ new_n19283;
  assign new_n19689 = new_n19239 & new_n19688;
  assign new_n19690 = new_n19689 ^ new_n19687;
  assign new_n19691 = new_n19242 & new_n19312;
  assign new_n19692 = new_n19691 ^ new_n19690;
  assign new_n19693 = new_n19692 ^ new_n19679;
  assign new_n19694 = new_n19442 ^ new_n19421;
  assign new_n19695 = ~new_n19363 & ~new_n19694;
  assign new_n19696 = new_n19695 ^ new_n19628;
  assign new_n19697 = new_n19382 & new_n19453;
  assign new_n19698 = new_n19697 ^ new_n19696;
  assign new_n19699 = new_n19698 ^ new_n19624;
  assign new_n19700 = new_n19699 ^ new_n19693;
  assign new_n19701 = new_n19607 ^ new_n19580;
  assign new_n19702 = new_n19567 ^ new_n19521;
  assign new_n19703 = new_n19563 ^ new_n19514;
  assign new_n19704 = new_n19703 ^ new_n19591;
  assign new_n19705 = new_n19704 ^ new_n19702;
  assign new_n19706 = ~new_n19705 & new_n19535;
  assign new_n19707 = new_n19561 & new_n19584;
  assign new_n19708 = ~new_n19705 & new_n19556;
  assign new_n19709 = new_n19708 ^ new_n19707;
  assign new_n19710 = new_n19588 ^ new_n19576;
  assign new_n19711 = new_n19710 ^ new_n19553;
  assign new_n19712 = new_n19524 & new_n19711;
  assign new_n19713 = new_n19574 ^ new_n19567;
  assign new_n19714 = new_n19498 & new_n19713;
  assign new_n19715 = new_n19714 ^ new_n19602;
  assign new_n19716 = new_n19715 ^ new_n19712;
  assign new_n19717 = new_n19716 ^ new_n19709;
  assign new_n19718 = new_n19717 ^ new_n19706;
  assign new_n19719 = new_n19718 ^ new_n19701;
  assign new_n19720 = new_n19719 ^ new_n19463;
  assign new_n19721 = new_n19720 ^ new_n19700;
  assign new_n19722 = new_n19721 ^ new_n19673;
  assign new_n19723 = new_n19722 ^ new_n19633;
  assign new_n19724 = new_n19021 ^ new_n18997;
  assign new_n19725 = new_n19005 ^ new_n18988;
  assign new_n19726 = new_n18933 & new_n19725;
  assign new_n19727 = new_n19726 ^ new_n19027;
  assign new_n19728 = new_n18949 & new_n19644;
  assign new_n19729 = new_n19728 ^ new_n19727;
  assign new_n19730 = new_n19729 ^ new_n19013;
  assign new_n19731 = new_n19730 ^ new_n19724;
  assign new_n19732 = new_n19731 ^ new_n16506;
  assign new_n19733 = new_n19163 ^ new_n19139;
  assign new_n19734 = new_n19147 ^ new_n19130;
  assign new_n19735 = ~new_n19067 & new_n19734;
  assign new_n19736 = new_n19735 ^ new_n19169;
  assign new_n19737 = ~new_n19092 & new_n19664;
  assign new_n19738 = new_n19737 ^ new_n19736;
  assign new_n19739 = new_n19738 ^ new_n19155;
  assign new_n19740 = new_n19739 ^ new_n19733;
  assign new_n19741 = new_n19740 ^ new_n19732;
  assign new_n19742 = ~new_n19683 & new_n19249;
  assign new_n19743 = new_n19742 ^ new_n19292;
  assign new_n19744 = new_n19687 ^ new_n19679;
  assign new_n19745 = new_n19744 ^ new_n19743;
  assign new_n19746 = new_n19745 ^ new_n19630;
  assign new_n19747 = new_n19604 ^ new_n19580;
  assign new_n19748 = new_n19588 ^ new_n19571;
  assign new_n19749 = new_n19506 & new_n19748;
  assign new_n19750 = new_n19749 ^ new_n19610;
  assign new_n19751 = new_n19532 & new_n19711;
  assign new_n19752 = new_n19751 ^ new_n19750;
  assign new_n19753 = new_n19752 ^ new_n19596;
  assign new_n19754 = new_n19753 ^ new_n19747;
  assign new_n19755 = new_n19623 ^ new_n19430;
  assign new_n19756 = new_n19698 ^ new_n19617;
  assign new_n19757 = new_n19756 ^ new_n19755;
  assign new_n19758 = new_n19757 ^ new_n19754;
  assign new_n19759 = new_n19758 ^ new_n19746;
  assign new_n19760 = new_n19759 ^ new_n19741;
  assign new_n19761 = new_n19273 & new_n19300;
  assign new_n19762 = new_n19761 ^ new_n19678;
  assign new_n19763 = new_n19676 ^ new_n19317;
  assign new_n19764 = new_n19763 ^ new_n19690;
  assign new_n19765 = new_n19764 ^ new_n19762;
  assign new_n19766 = ~new_n19412 & ~new_n19438;
  assign new_n19767 = new_n19766 ^ new_n19623;
  assign new_n19768 = new_n19621 ^ new_n19458;
  assign new_n19769 = new_n19768 ^ new_n19696;
  assign new_n19770 = new_n19769 ^ new_n19767;
  assign new_n19771 = new_n19770 ^ new_n19765;
  assign new_n19772 = new_n19752 ^ new_n19605;
  assign new_n19773 = new_n19772 ^ new_n19699;
  assign new_n19774 = new_n19773 ^ new_n19771;
  assign new_n19775 = new_n19729 ^ new_n19022;
  assign new_n19776 = new_n19775 ^ new_n16502;
  assign new_n19777 = new_n19738 ^ new_n19164;
  assign new_n19778 = new_n19777 ^ new_n19776;
  assign new_n19779 = new_n19678 ^ new_n19292;
  assign new_n19780 = new_n19742 ^ new_n19692;
  assign new_n19781 = new_n19780 ^ new_n19779;
  assign new_n19782 = new_n19781 ^ new_n19757;
  assign new_n19783 = new_n19782 ^ new_n19778;
  assign new_n19784 = new_n19783 ^ new_n19774;
  assign new_n19785 = new_n19784 ^ new_n19760;
  assign new_n19786 = new_n19257 & new_n19688;
  assign new_n19787 = new_n19786 ^ new_n19761;
  assign new_n19788 = new_n19787 ^ new_n19685;
  assign new_n19789 = new_n19691 ^ new_n19319;
  assign new_n19790 = new_n19789 ^ new_n19788;
  assign new_n19791 = new_n19697 ^ new_n19460;
  assign new_n19792 = ~new_n19694 & new_n19397;
  assign new_n19793 = new_n19792 ^ new_n19766;
  assign new_n19794 = new_n19793 ^ new_n19627;
  assign new_n19795 = new_n19794 ^ new_n19791;
  assign new_n19796 = new_n19795 ^ new_n19790;
  assign new_n19797 = new_n19454 ^ new_n19449;
  assign new_n19798 = new_n19695 ^ new_n19617;
  assign new_n19799 = new_n19798 ^ new_n19794;
  assign new_n19800 = new_n19799 ^ new_n19797;
  assign new_n19801 = new_n19712 ^ new_n19708;
  assign new_n19802 = new_n19749 ^ new_n19596;
  assign new_n19803 = new_n19547 & new_n19748;
  assign new_n19804 = new_n19562 & new_n19584;
  assign new_n19805 = new_n19804 ^ new_n19803;
  assign new_n19806 = new_n19805 ^ new_n19609;
  assign new_n19807 = new_n19806 ^ new_n19802;
  assign new_n19808 = new_n19807 ^ new_n19801;
  assign new_n19809 = new_n19808 ^ new_n19800;
  assign new_n19810 = new_n19809 ^ new_n19796;
  assign new_n19811 = new_n19645 ^ new_n19641;
  assign new_n19812 = new_n19726 ^ new_n19013;
  assign new_n19813 = new_n18965 & new_n19725;
  assign new_n19814 = new_n18979 & new_n19001;
  assign new_n19815 = new_n19814 ^ new_n19813;
  assign new_n19816 = new_n19815 ^ new_n19026;
  assign new_n19817 = new_n19816 ^ new_n19812;
  assign new_n19818 = new_n19817 ^ new_n19811;
  assign new_n19819 = new_n19818 ^ new_n16512;
  assign new_n19820 = new_n19665 ^ new_n19661;
  assign new_n19821 = new_n19735 ^ new_n19155;
  assign new_n19822 = ~new_n19107 & new_n19734;
  assign new_n19823 = new_n19121 & new_n19143;
  assign new_n19824 = new_n19823 ^ new_n19822;
  assign new_n19825 = new_n19824 ^ new_n19168;
  assign new_n19826 = new_n19825 ^ new_n19821;
  assign new_n19827 = new_n19826 ^ new_n19820;
  assign new_n19828 = new_n19827 ^ new_n19819;
  assign new_n19829 = new_n19828 ^ new_n19782;
  assign new_n19830 = new_n19829 ^ new_n19810;
  assign new_n19831 = new_n19814 ^ new_n19021;
  assign new_n19832 = new_n19647 ^ new_n19017;
  assign new_n19833 = new_n19832 ^ new_n19727;
  assign new_n19834 = new_n19833 ^ new_n19831;
  assign new_n19835 = new_n19834 ^ new_n16516;
  assign new_n19836 = new_n19823 ^ new_n19163;
  assign new_n19837 = new_n19667 ^ new_n19159;
  assign new_n19838 = new_n19837 ^ new_n19736;
  assign new_n19839 = new_n19838 ^ new_n19836;
  assign new_n19840 = new_n19839 ^ new_n19835;
  assign new_n19841 = new_n19840 ^ new_n19782;
  assign new_n19842 = ~new_n19364 & new_n19457;
  assign new_n19843 = new_n19842 ^ new_n19756;
  assign new_n19844 = new_n19843 ^ new_n19461;
  assign new_n19845 = new_n19239 ^ new_n19215;
  assign new_n19846 = new_n19316 & new_n19845;
  assign new_n19847 = new_n19846 ^ new_n19780;
  assign new_n19848 = new_n19847 ^ new_n19323;
  assign new_n19849 = new_n19848 ^ new_n19844;
  assign new_n19850 = new_n19804 ^ new_n19604;
  assign new_n19851 = new_n19714 ^ new_n19600;
  assign new_n19852 = new_n19851 ^ new_n19750;
  assign new_n19853 = new_n19852 ^ new_n19850;
  assign new_n19854 = new_n19853 ^ new_n19770;
  assign new_n19855 = new_n19854 ^ new_n19849;
  assign new_n19856 = new_n19855 ^ new_n19841;
  assign new_n19857 = new_n19856 ^ new_n19830;
  assign new_n19858 = new_n19857 ^ new_n19785;
  assign new_n19859 = new_n19858 ^ new_n19723;
  assign new_n19860 = new_n19728 ^ new_n19649;
  assign new_n19861 = new_n19860 ^ new_n19816;
  assign new_n19862 = new_n19861 ^ new_n16536;
  assign new_n19863 = new_n19737 ^ new_n19669;
  assign new_n19864 = new_n19863 ^ new_n19825;
  assign new_n19865 = new_n19864 ^ new_n19862;
  assign new_n19866 = new_n19751 ^ new_n19716;
  assign new_n19867 = new_n19866 ^ new_n19806;
  assign new_n19868 = new_n19867 ^ new_n19795;
  assign new_n19869 = new_n19868 ^ new_n19782;
  assign new_n19870 = new_n19869 ^ new_n19865;
  assign new_n19871 = new_n19870 ^ new_n19723;
  assign new_n19872 = new_n19871 ^ new_n19784;
  assign new_n19873 = new_n19870 & new_n19872;
  assign new_n19874 = new_n19873 ^ new_n19784;
  assign new_n19875 = new_n19830 ^ new_n19784;
  assign new_n19876 = new_n18935 & new_n19646;
  assign new_n19877 = new_n19876 ^ new_n19730;
  assign new_n19878 = new_n19877 ^ new_n19650;
  assign new_n19879 = new_n19878 ^ new_n16524;
  assign new_n19880 = ~new_n19666 & new_n19074;
  assign new_n19881 = new_n19880 ^ new_n19739;
  assign new_n19882 = new_n19881 ^ new_n19670;
  assign new_n19883 = new_n19882 ^ new_n19879;
  assign new_n19884 = new_n19320 ^ new_n19313;
  assign new_n19885 = new_n19742 ^ new_n19689;
  assign new_n19886 = new_n19885 ^ new_n19788;
  assign new_n19887 = new_n19886 ^ new_n19884;
  assign new_n19888 = new_n19887 ^ new_n19800;
  assign new_n19889 = new_n19513 & new_n19713;
  assign new_n19890 = new_n19889 ^ new_n19753;
  assign new_n19891 = new_n19890 ^ new_n19717;
  assign new_n19892 = new_n19891 ^ new_n19844;
  assign new_n19893 = new_n19892 ^ new_n19888;
  assign new_n19894 = new_n19893 ^ new_n19883;
  assign new_n19895 = new_n19894 ^ new_n19760;
  assign new_n19896 = new_n19895 ^ new_n19875;
  assign new_n19897 = new_n19858 & new_n19896;
  assign new_n19898 = new_n19897 ^ new_n19633;
  assign new_n19899 = new_n19898 ^ new_n19874;
  assign new_n19900 = new_n19898 ^ new_n19858;
  assign new_n19901 = new_n19870 ^ new_n19858;
  assign new_n19902 = new_n19871 ^ new_n19830;
  assign new_n19903 = new_n19902 ^ new_n19895;
  assign new_n19904 = new_n19901 & new_n19903;
  assign new_n19905 = new_n19894 ^ new_n19857;
  assign new_n19906 = new_n19905 ^ new_n19633;
  assign new_n19907 = new_n19785 & new_n19906;
  assign new_n19908 = new_n19907 ^ new_n19904;
  assign new_n19909 = new_n19784 ^ new_n19722;
  assign new_n19910 = new_n19909 ^ new_n19895;
  assign new_n19911 = new_n19894 ^ new_n19784;
  assign new_n19912 = new_n19910 & new_n19911;
  assign new_n19913 = new_n19912 ^ new_n19894;
  assign new_n19914 = new_n19913 ^ new_n19908;
  assign new_n19915 = new_n19914 ^ new_n19900;
  assign new_n19916 = ~new_n19830 & ~new_n19871;
  assign new_n19917 = new_n19916 ^ new_n19830;
  assign new_n19918 = new_n19905 ^ new_n19722;
  assign new_n19919 = new_n19830 ^ new_n19760;
  assign new_n19920 = new_n19918 & new_n19919;
  assign new_n19921 = new_n19920 ^ new_n19917;
  assign new_n19922 = new_n19921 ^ new_n19895;
  assign new_n19923 = new_n19912 ^ new_n19907;
  assign new_n19924 = new_n19856 ^ new_n19722;
  assign new_n19925 = new_n19924 ^ new_n19923;
  assign new_n19926 = new_n19925 ^ new_n19922;
  assign new_n19927 = ~new_n19926 & new_n19915;
  assign new_n19928 = new_n19927 ^ new_n19899;
  assign new_n19929 = new_n19859 & new_n19895;
  assign new_n19930 = new_n19929 ^ new_n19907;
  assign new_n19931 = new_n19930 ^ new_n19918;
  assign new_n19932 = new_n19931 ^ new_n19928;
  assign new_n19933 = new_n19871 ^ new_n19760;
  assign new_n19934 = new_n19906 ^ new_n19870;
  assign new_n19935 = new_n19933 & new_n19934;
  assign new_n19936 = new_n19935 ^ new_n19916;
  assign new_n19937 = new_n19929 ^ new_n19912;
  assign new_n19938 = new_n19937 ^ new_n19936;
  assign new_n19939 = ~new_n19938 & new_n19932;
  assign new_n19940 = new_n19939 ^ new_n19760;
  assign new_n19941 = new_n19935 ^ new_n19873;
  assign new_n19942 = new_n19830 ^ new_n19722;
  assign new_n19943 = new_n19917 ^ new_n19904;
  assign new_n19944 = new_n19935 ^ new_n19920;
  assign new_n19945 = new_n19944 ^ new_n19760;
  assign new_n19946 = new_n19945 ^ new_n19931;
  assign new_n19947 = new_n19939 ^ new_n19927;
  assign new_n19948 = ~new_n19946 & ~new_n19947;
  assign new_n19949 = new_n19948 ^ new_n19939;
  assign new_n19950 = new_n19946 ^ new_n19927;
  assign new_n19951 = new_n19760 ^ new_n19722;
  assign new_n19952 = new_n19904 ^ new_n19873;
  assign new_n19953 = new_n19952 ^ new_n19937;
  assign new_n19954 = new_n19953 ^ new_n19951;
  assign new_n19955 = new_n19950 & new_n19954;
  assign new_n19956 = new_n19955 ^ new_n19899;
  assign new_n19957 = new_n19956 ^ new_n19931;
  assign new_n19958 = ~new_n19949 & new_n19957;
  assign new_n19959 = new_n19950 ^ new_n19949;
  assign new_n19960 = new_n19959 ^ new_n19958;
  assign new_n19961 = new_n19960 ^ new_n19943;
  assign new_n19962 = new_n19961 ^ new_n19942;
  assign new_n19963 = new_n19962 ^ new_n19941;
  assign new_n19964 = new_n19963 ^ new_n19940;
  assign new_n19965 = new_n19859 & new_n19964;
  assign new_n19966 = new_n19958 ^ new_n19955;
  assign new_n19967 = new_n19966 ^ new_n19915;
  assign new_n19968 = new_n19919 & new_n19967;
  assign new_n19969 = new_n19968 ^ new_n19965;
  assign new_n19970 = new_n19962 ^ new_n19784;
  assign new_n19971 = new_n19955 ^ new_n19920;
  assign new_n19972 = new_n19971 ^ new_n19898;
  assign new_n19973 = new_n19972 ^ new_n19970;
  assign new_n19974 = new_n19910 & new_n19973;
  assign new_n19975 = new_n19958 ^ new_n19954;
  assign new_n19976 = new_n19871 & new_n19975;
  assign new_n19977 = new_n19976 ^ new_n19974;
  assign new_n19978 = new_n19902 & new_n19975;
  assign new_n19979 = new_n19934 & new_n19957;
  assign new_n19980 = new_n19979 ^ new_n19978;
  assign new_n19981 = new_n19955 ^ new_n19939;
  assign new_n19982 = new_n19945 ^ new_n19899;
  assign new_n19983 = new_n19982 ^ new_n19981;
  assign new_n19984 = new_n19785 & new_n19983;
  assign new_n19985 = new_n19911 & new_n19973;
  assign new_n19986 = new_n19985 ^ new_n19984;
  assign new_n19987 = new_n19986 ^ new_n19980;
  assign new_n19988 = new_n19987 ^ new_n19977;
  assign new_n19989 = new_n19988 ^ new_n19969;
  assign new_n19990 = new_n19989 ^ new_n18922;
  assign new_n19991 = new_n18875 ^ new_n18840;
  assign new_n19992 = new_n18832 & new_n19991;
  assign new_n19993 = new_n18895 ^ new_n18868;
  assign new_n19994 = new_n18813 & new_n19993;
  assign new_n19995 = new_n19994 ^ new_n19992;
  assign new_n19996 = new_n19995 ^ new_n18890;
  assign new_n19997 = new_n18820 & new_n18889;
  assign new_n19998 = new_n19997 ^ new_n19996;
  assign new_n19999 = new_n19998 ^ new_n18920;
  assign new_n20000 = new_n19999 ^ new_n19990;
  assign new_n20001 = new_n18895 ^ new_n18875;
  assign new_n20002 = new_n20001 ^ new_n18874;
  assign new_n20003 = new_n18857 & new_n20002;
  assign new_n20004 = new_n20003 ^ new_n18919;
  assign new_n20005 = new_n20004 ^ new_n18909;
  assign new_n20006 = new_n20005 ^ new_n19997;
  assign new_n20007 = new_n20006 ^ new_n18907;
  assign new_n20008 = ~new_n18817 & new_n18916;
  assign new_n20009 = new_n18845 & new_n19993;
  assign new_n20010 = new_n20009 ^ new_n20008;
  assign new_n20011 = new_n20010 ^ new_n20007;
  assign new_n20012 = new_n19206 ^ new_n15114;
  assign new_n20013 = new_n16209 ^ new_n11407;
  assign new_n20014 = new_n20013 ^ new_n432;
  assign new_n20015 = new_n20014 ^ new_n15134;
  assign new_n20016 = new_n20015 ^ new_n15180;
  assign new_n20017 = new_n20016 ^ new_n20012;
  assign new_n20018 = new_n19199 ^ new_n15180;
  assign new_n20019 = new_n16253 ^ new_n10299;
  assign new_n20020 = new_n20019 ^ new_n443;
  assign new_n20021 = new_n20020 ^ new_n15196;
  assign new_n20022 = new_n20021 ^ new_n20018;
  assign new_n20023 = new_n20022 ^ new_n20017;
  assign new_n20024 = new_n15157 ^ new_n15053;
  assign new_n20025 = new_n20024 ^ new_n15079;
  assign new_n20026 = new_n20025 ^ new_n19192;
  assign new_n20027 = new_n16130 ^ new_n11536;
  assign new_n20028 = new_n20027 ^ new_n392;
  assign new_n20029 = new_n20028 ^ new_n15099;
  assign new_n20030 = new_n20029 ^ new_n15210;
  assign new_n20031 = new_n20030 ^ new_n20026;
  assign new_n20032 = new_n15027 ^ new_n11692;
  assign new_n20033 = new_n20032 ^ new_n13828;
  assign new_n20034 = new_n16148 ^ new_n11503;
  assign new_n20035 = new_n20034 ^ new_n402;
  assign new_n20036 = new_n20035 ^ new_n20024;
  assign new_n20037 = new_n20036 ^ new_n19209;
  assign new_n20038 = new_n20037 ^ new_n20033;
  assign new_n20039 = new_n20038 ^ new_n20031;
  assign new_n20040 = new_n19176 ^ new_n15140;
  assign new_n20041 = new_n16232 ^ new_n11559;
  assign new_n20042 = new_n20041 ^ new_n364;
  assign new_n20043 = new_n20042 ^ new_n15157;
  assign new_n20044 = new_n20043 ^ new_n15134;
  assign new_n20045 = new_n20044 ^ new_n20040;
  assign new_n20046 = new_n16262 ^ new_n11464;
  assign new_n20047 = new_n20046 ^ new_n373;
  assign new_n20048 = new_n20047 ^ new_n19231;
  assign new_n20049 = new_n20048 ^ new_n20024;
  assign new_n20050 = new_n15195 ^ new_n15012;
  assign new_n20051 = new_n20050 ^ new_n15027;
  assign new_n20052 = new_n20051 ^ new_n20049;
  assign new_n20053 = new_n20052 ^ new_n20045;
  assign new_n20054 = new_n20053 ^ new_n20039;
  assign new_n20055 = new_n20054 ^ new_n20023;
  assign new_n20056 = new_n16278 ^ new_n11424;
  assign new_n20057 = new_n20056 ^ new_n412;
  assign new_n20058 = new_n20057 ^ new_n15210;
  assign new_n20059 = new_n20024 ^ new_n19181;
  assign new_n20060 = new_n20059 ^ new_n20058;
  assign new_n20061 = new_n20060 ^ new_n20023;
  assign new_n20062 = new_n20061 ^ new_n20052;
  assign new_n20063 = new_n20060 & new_n20062;
  assign new_n20064 = new_n20063 ^ new_n20052;
  assign new_n20065 = new_n19178 ^ new_n14089;
  assign new_n20066 = new_n15732 ^ new_n11581;
  assign new_n20067 = new_n20066 ^ new_n424;
  assign new_n20068 = new_n20067 ^ new_n13828;
  assign new_n20069 = new_n20068 ^ new_n15099;
  assign new_n20070 = new_n20069 ^ new_n20065;
  assign new_n20071 = new_n20070 ^ new_n20052;
  assign new_n20072 = new_n20045 ^ new_n20031;
  assign new_n20073 = new_n20072 ^ new_n20071;
  assign new_n20074 = new_n20054 & new_n20073;
  assign new_n20075 = new_n20074 ^ new_n20017;
  assign new_n20076 = new_n20075 ^ new_n20064;
  assign new_n20077 = new_n20075 ^ new_n20054;
  assign new_n20078 = new_n20060 ^ new_n20054;
  assign new_n20079 = new_n20061 ^ new_n20031;
  assign new_n20080 = new_n20070 ^ new_n20045;
  assign new_n20081 = new_n20080 ^ new_n20079;
  assign new_n20082 = new_n20078 & new_n20081;
  assign new_n20083 = new_n20070 ^ new_n20039;
  assign new_n20084 = new_n20083 ^ new_n20017;
  assign new_n20085 = new_n20053 & new_n20084;
  assign new_n20086 = new_n20085 ^ new_n20082;
  assign new_n20087 = new_n20052 ^ new_n20022;
  assign new_n20088 = new_n20087 ^ new_n20080;
  assign new_n20089 = new_n20071 & new_n20088;
  assign new_n20090 = new_n20089 ^ new_n20070;
  assign new_n20091 = new_n20090 ^ new_n20086;
  assign new_n20092 = new_n20091 ^ new_n20077;
  assign new_n20093 = ~new_n20031 & ~new_n20061;
  assign new_n20094 = new_n20093 ^ new_n20031;
  assign new_n20095 = new_n20083 ^ new_n20022;
  assign new_n20096 = new_n20072 & new_n20095;
  assign new_n20097 = new_n20096 ^ new_n20094;
  assign new_n20098 = new_n20097 ^ new_n20080;
  assign new_n20099 = new_n20089 ^ new_n20085;
  assign new_n20100 = new_n20038 ^ new_n20022;
  assign new_n20101 = new_n20100 ^ new_n20099;
  assign new_n20102 = new_n20101 ^ new_n20098;
  assign new_n20103 = ~new_n20102 & new_n20092;
  assign new_n20104 = new_n20103 ^ new_n20076;
  assign new_n20105 = new_n20055 & new_n20080;
  assign new_n20106 = new_n20105 ^ new_n20085;
  assign new_n20107 = new_n20106 ^ new_n20095;
  assign new_n20108 = new_n20107 ^ new_n20104;
  assign new_n20109 = new_n20105 ^ new_n20089;
  assign new_n20110 = new_n20061 ^ new_n20045;
  assign new_n20111 = new_n20084 ^ new_n20060;
  assign new_n20112 = new_n20110 & new_n20111;
  assign new_n20113 = new_n20112 ^ new_n20093;
  assign new_n20114 = new_n20113 ^ new_n20109;
  assign new_n20115 = ~new_n20114 & new_n20108;
  assign new_n20116 = new_n20115 ^ new_n20045;
  assign new_n20117 = new_n20112 ^ new_n20063;
  assign new_n20118 = new_n20031 ^ new_n20022;
  assign new_n20119 = new_n20094 ^ new_n20082;
  assign new_n20120 = new_n20045 ^ new_n20022;
  assign new_n20121 = new_n20082 ^ new_n20063;
  assign new_n20122 = new_n20121 ^ new_n20109;
  assign new_n20123 = new_n20122 ^ new_n20120;
  assign new_n20124 = new_n20112 ^ new_n20096;
  assign new_n20125 = new_n20124 ^ new_n20045;
  assign new_n20126 = new_n20125 ^ new_n20107;
  assign new_n20127 = new_n20126 ^ new_n20103;
  assign new_n20128 = new_n20123 & new_n20127;
  assign new_n20129 = new_n20128 ^ new_n20076;
  assign new_n20130 = new_n20129 ^ new_n20107;
  assign new_n20131 = new_n20115 ^ new_n20103;
  assign new_n20132 = ~new_n20131 & new_n20126;
  assign new_n20133 = new_n20132 ^ new_n20103;
  assign new_n20134 = new_n20130 & new_n20133;
  assign new_n20135 = new_n20132 ^ new_n20126;
  assign new_n20136 = new_n20135 ^ new_n20134;
  assign new_n20137 = new_n20136 ^ new_n20119;
  assign new_n20138 = new_n20137 ^ new_n20118;
  assign new_n20139 = new_n20138 ^ new_n20117;
  assign new_n20140 = new_n20139 ^ new_n20116;
  assign new_n20141 = ~new_n20140 & new_n20055;
  assign new_n20142 = new_n20134 ^ new_n20128;
  assign new_n20143 = new_n20142 ^ new_n20092;
  assign new_n20144 = new_n20072 & new_n20143;
  assign new_n20145 = new_n20144 ^ new_n20141;
  assign new_n20146 = new_n20138 ^ new_n20052;
  assign new_n20147 = new_n20128 ^ new_n20096;
  assign new_n20148 = new_n20147 ^ new_n20075;
  assign new_n20149 = new_n20148 ^ new_n20146;
  assign new_n20150 = ~new_n20149 & new_n20088;
  assign new_n20151 = new_n20134 ^ new_n20123;
  assign new_n20152 = new_n20061 & new_n20151;
  assign new_n20153 = new_n20152 ^ new_n20150;
  assign new_n20154 = new_n20079 & new_n20151;
  assign new_n20155 = new_n20111 & new_n20130;
  assign new_n20156 = new_n20155 ^ new_n20154;
  assign new_n20157 = new_n20128 ^ new_n20115;
  assign new_n20158 = new_n20125 ^ new_n20076;
  assign new_n20159 = new_n20158 ^ new_n20157;
  assign new_n20160 = new_n20053 & new_n20159;
  assign new_n20161 = ~new_n20149 & new_n20071;
  assign new_n20162 = new_n20161 ^ new_n20160;
  assign new_n20163 = new_n20162 ^ new_n20156;
  assign new_n20164 = new_n20163 ^ new_n20153;
  assign new_n20165 = new_n20164 ^ new_n20145;
  assign new_n20166 = new_n19367 ^ new_n16215;
  assign new_n20167 = new_n17241 ^ new_n6084;
  assign new_n20168 = new_n20167 ^ new_n16186;
  assign new_n20169 = new_n20168 ^ new_n16240;
  assign new_n20170 = new_n20169 ^ new_n20166;
  assign new_n20171 = new_n19343 ^ new_n16240;
  assign new_n20172 = new_n16258 ^ new_n16248;
  assign new_n20173 = new_n17269 ^ new_n6088;
  assign new_n20174 = new_n20173 ^ new_n20172;
  assign new_n20175 = new_n20174 ^ new_n20171;
  assign new_n20176 = new_n20175 ^ new_n20170;
  assign new_n20177 = new_n19329 ^ new_n16203;
  assign new_n20178 = new_n17290 ^ new_n6078;
  assign new_n20179 = new_n20178 ^ new_n16228;
  assign new_n20180 = new_n20179 ^ new_n16186;
  assign new_n20181 = new_n20180 ^ new_n20177;
  assign new_n20182 = new_n17315 ^ new_n6079;
  assign new_n20183 = new_n20182 ^ new_n19369;
  assign new_n20184 = new_n20183 ^ new_n19357;
  assign new_n20185 = new_n16258 ^ new_n16163;
  assign new_n20186 = new_n20185 ^ new_n16169;
  assign new_n20187 = new_n20186 ^ new_n20184;
  assign new_n20188 = new_n20187 ^ new_n20181;
  assign new_n20189 = new_n19369 ^ new_n16105;
  assign new_n20190 = new_n20189 ^ new_n19339;
  assign new_n20191 = new_n17165 ^ new_n6075;
  assign new_n20192 = new_n20191 ^ new_n16140;
  assign new_n20193 = new_n20192 ^ new_n16282;
  assign new_n20194 = new_n20193 ^ new_n20190;
  assign new_n20195 = new_n16169 ^ new_n15754;
  assign new_n20196 = new_n20195 ^ new_n16082;
  assign new_n20197 = new_n17185 ^ new_n6076;
  assign new_n20198 = new_n20197 ^ new_n19352;
  assign new_n20199 = new_n20198 ^ new_n19369;
  assign new_n20200 = new_n20199 ^ new_n20196;
  assign new_n20201 = new_n20200 ^ new_n20194;
  assign new_n20202 = new_n20201 ^ new_n20188;
  assign new_n20203 = new_n20202 ^ new_n20176;
  assign new_n20204 = new_n20194 ^ new_n20187;
  assign new_n20205 = new_n19326 ^ new_n15460;
  assign new_n20206 = new_n16499 ^ new_n6082;
  assign new_n20207 = new_n20206 ^ new_n16082;
  assign new_n20208 = new_n20207 ^ new_n16140;
  assign new_n20209 = new_n20208 ^ new_n20205;
  assign new_n20210 = new_n20209 ^ new_n20181;
  assign new_n20211 = new_n20210 ^ new_n20204;
  assign new_n20212 = new_n20202 & new_n20211;
  assign new_n20213 = new_n20212 ^ new_n20170;
  assign new_n20214 = new_n20213 ^ new_n20202;
  assign new_n20215 = new_n17298 ^ new_n6097;
  assign new_n20216 = new_n20215 ^ new_n16282;
  assign new_n20217 = new_n19369 ^ new_n19333;
  assign new_n20218 = new_n20217 ^ new_n20216;
  assign new_n20219 = new_n20218 ^ new_n20202;
  assign new_n20220 = new_n20218 ^ new_n20176;
  assign new_n20221 = new_n20220 ^ new_n20194;
  assign new_n20222 = new_n20221 ^ new_n20210;
  assign new_n20223 = ~new_n20222 & new_n20219;
  assign new_n20224 = new_n20209 ^ new_n20201;
  assign new_n20225 = new_n20224 ^ new_n20170;
  assign new_n20226 = ~new_n20188 & new_n20225;
  assign new_n20227 = new_n20226 ^ new_n20223;
  assign new_n20228 = new_n20187 ^ new_n20175;
  assign new_n20229 = new_n20228 ^ new_n20210;
  assign new_n20230 = new_n20209 ^ new_n20187;
  assign new_n20231 = ~new_n20230 & new_n20229;
  assign new_n20232 = new_n20231 ^ new_n20209;
  assign new_n20233 = new_n20232 ^ new_n20227;
  assign new_n20234 = new_n20233 ^ new_n20214;
  assign new_n20235 = ~new_n20220 & new_n20194;
  assign new_n20236 = new_n20235 ^ new_n20194;
  assign new_n20237 = new_n20224 ^ new_n20175;
  assign new_n20238 = new_n20194 ^ new_n20181;
  assign new_n20239 = ~new_n20238 & new_n20237;
  assign new_n20240 = new_n20239 ^ new_n20236;
  assign new_n20241 = new_n20240 ^ new_n20210;
  assign new_n20242 = new_n20231 ^ new_n20226;
  assign new_n20243 = new_n20200 ^ new_n20175;
  assign new_n20244 = new_n20243 ^ new_n20242;
  assign new_n20245 = new_n20244 ^ new_n20241;
  assign new_n20246 = ~new_n20234 & ~new_n20245;
  assign new_n20247 = new_n20220 ^ new_n20187;
  assign new_n20248 = ~new_n20247 & new_n20218;
  assign new_n20249 = new_n20248 ^ new_n20187;
  assign new_n20250 = new_n20249 ^ new_n20213;
  assign new_n20251 = new_n20250 ^ new_n20246;
  assign new_n20252 = new_n20203 & new_n20210;
  assign new_n20253 = new_n20252 ^ new_n20226;
  assign new_n20254 = new_n20253 ^ new_n20237;
  assign new_n20255 = new_n20254 ^ new_n20251;
  assign new_n20256 = new_n20252 ^ new_n20231;
  assign new_n20257 = new_n20220 ^ new_n20181;
  assign new_n20258 = new_n20225 ^ new_n20218;
  assign new_n20259 = new_n20257 & new_n20258;
  assign new_n20260 = new_n20259 ^ new_n20235;
  assign new_n20261 = new_n20260 ^ new_n20256;
  assign new_n20262 = ~new_n20261 & new_n20255;
  assign new_n20263 = new_n20262 ^ new_n20181;
  assign new_n20264 = new_n20259 ^ new_n20248;
  assign new_n20265 = new_n20194 ^ new_n20175;
  assign new_n20266 = new_n20236 ^ new_n20223;
  assign new_n20267 = new_n20181 ^ new_n20175;
  assign new_n20268 = new_n20248 ^ new_n20223;
  assign new_n20269 = new_n20268 ^ new_n20256;
  assign new_n20270 = new_n20269 ^ new_n20267;
  assign new_n20271 = new_n20259 ^ new_n20239;
  assign new_n20272 = new_n20271 ^ new_n20181;
  assign new_n20273 = new_n20272 ^ new_n20254;
  assign new_n20274 = new_n20273 ^ new_n20246;
  assign new_n20275 = ~new_n20270 & new_n20274;
  assign new_n20276 = new_n20275 ^ new_n20250;
  assign new_n20277 = new_n20276 ^ new_n20254;
  assign new_n20278 = new_n20262 ^ new_n20246;
  assign new_n20279 = ~new_n20278 & new_n20273;
  assign new_n20280 = new_n20279 ^ new_n20246;
  assign new_n20281 = new_n20277 & new_n20280;
  assign new_n20282 = new_n20279 ^ new_n20273;
  assign new_n20283 = new_n20282 ^ new_n20281;
  assign new_n20284 = new_n20283 ^ new_n20266;
  assign new_n20285 = new_n20284 ^ new_n20265;
  assign new_n20286 = new_n20285 ^ new_n20264;
  assign new_n20287 = new_n20286 ^ new_n20263;
  assign new_n20288 = new_n20203 & new_n20287;
  assign new_n20289 = new_n20281 ^ new_n20275;
  assign new_n20290 = new_n20289 ^ new_n20234;
  assign new_n20291 = ~new_n20238 & ~new_n20290;
  assign new_n20292 = new_n20291 ^ new_n20288;
  assign new_n20293 = new_n20285 ^ new_n20187;
  assign new_n20294 = new_n20275 ^ new_n20239;
  assign new_n20295 = new_n20294 ^ new_n20213;
  assign new_n20296 = new_n20295 ^ new_n20293;
  assign new_n20297 = new_n20229 & new_n20296;
  assign new_n20298 = new_n20281 ^ new_n20270;
  assign new_n20299 = ~new_n20298 & new_n20220;
  assign new_n20300 = new_n20299 ^ new_n20297;
  assign new_n20301 = ~new_n20221 & ~new_n20298;
  assign new_n20302 = new_n20258 & new_n20277;
  assign new_n20303 = new_n20302 ^ new_n20301;
  assign new_n20304 = ~new_n20230 & new_n20296;
  assign new_n20305 = new_n20275 ^ new_n20262;
  assign new_n20306 = new_n20272 ^ new_n20250;
  assign new_n20307 = new_n20306 ^ new_n20305;
  assign new_n20308 = ~new_n20188 & new_n20307;
  assign new_n20309 = new_n20308 ^ new_n20304;
  assign new_n20310 = new_n20309 ^ new_n20303;
  assign new_n20311 = new_n20310 ^ new_n20300;
  assign new_n20312 = new_n20311 ^ new_n20292;
  assign new_n20313 = new_n20312 ^ new_n20165;
  assign new_n20314 = new_n20182 ^ new_n20178;
  assign new_n20315 = new_n20197 ^ new_n20191;
  assign new_n20316 = new_n20315 ^ new_n20314;
  assign new_n20317 = new_n20191 ^ new_n20182;
  assign new_n20318 = new_n20206 ^ new_n20178;
  assign new_n20319 = new_n20318 ^ new_n20317;
  assign new_n20320 = ~new_n20316 & ~new_n20319;
  assign new_n20321 = new_n20320 ^ new_n20167;
  assign new_n20322 = new_n20173 ^ new_n20167;
  assign new_n20323 = ~new_n20215 & ~new_n20322;
  assign new_n20324 = ~new_n20182 & new_n20215;
  assign new_n20325 = new_n20324 ^ new_n20323;
  assign new_n20326 = new_n20325 ^ new_n20321;
  assign new_n20327 = new_n20321 ^ new_n20316;
  assign new_n20328 = new_n20206 ^ new_n20182;
  assign new_n20329 = new_n20178 ^ new_n20173;
  assign new_n20330 = new_n20329 ^ new_n20328;
  assign new_n20331 = ~new_n20328 & ~new_n20330;
  assign new_n20332 = new_n20315 ^ new_n20206;
  assign new_n20333 = new_n20332 ^ new_n20167;
  assign new_n20334 = ~new_n20314 & new_n20333;
  assign new_n20335 = new_n20334 ^ new_n20331;
  assign new_n20336 = new_n20316 ^ new_n20215;
  assign new_n20337 = new_n20322 ^ new_n20215;
  assign new_n20338 = new_n20337 ^ new_n20191;
  assign new_n20339 = new_n20338 ^ new_n20318;
  assign new_n20340 = ~new_n20339 & new_n20336;
  assign new_n20341 = new_n20340 ^ new_n20206;
  assign new_n20342 = new_n20341 ^ new_n20335;
  assign new_n20343 = new_n20342 ^ new_n20327;
  assign new_n20344 = ~new_n20191 & new_n20337;
  assign new_n20345 = new_n20344 ^ new_n20191;
  assign new_n20346 = new_n20332 ^ new_n20173;
  assign new_n20347 = new_n20191 ^ new_n20178;
  assign new_n20348 = new_n20346 & new_n20347;
  assign new_n20349 = new_n20348 ^ new_n20345;
  assign new_n20350 = new_n20349 ^ new_n20318;
  assign new_n20351 = new_n20197 ^ new_n20173;
  assign new_n20352 = new_n20351 ^ new_n20335;
  assign new_n20353 = new_n20352 ^ new_n20350;
  assign new_n20354 = ~new_n20343 & ~new_n20353;
  assign new_n20355 = new_n20354 ^ new_n20326;
  assign new_n20356 = new_n20322 ^ new_n20316;
  assign new_n20357 = ~new_n20356 & new_n20318;
  assign new_n20358 = new_n20357 ^ new_n20334;
  assign new_n20359 = new_n20358 ^ new_n20346;
  assign new_n20360 = new_n20359 ^ new_n20355;
  assign new_n20361 = new_n20357 ^ new_n20331;
  assign new_n20362 = new_n20337 ^ new_n20178;
  assign new_n20363 = new_n20333 ^ new_n20215;
  assign new_n20364 = ~new_n20362 & ~new_n20363;
  assign new_n20365 = new_n20364 ^ new_n20344;
  assign new_n20366 = new_n20365 ^ new_n20361;
  assign new_n20367 = ~new_n20366 & new_n20360;
  assign new_n20368 = new_n20364 ^ new_n20348;
  assign new_n20369 = new_n20368 ^ new_n20178;
  assign new_n20370 = new_n20369 ^ new_n20359;
  assign new_n20371 = new_n20370 ^ new_n20367;
  assign new_n20372 = new_n20337 ^ new_n20182;
  assign new_n20373 = new_n20371 & new_n20372;
  assign new_n20374 = new_n20325 ^ new_n20182;
  assign new_n20375 = new_n20374 ^ new_n20340;
  assign new_n20376 = new_n20375 ^ new_n20361;
  assign new_n20377 = new_n20376 ^ new_n20329;
  assign new_n20378 = new_n20370 ^ new_n20354;
  assign new_n20379 = ~new_n20377 & new_n20378;
  assign new_n20380 = new_n20379 ^ new_n20326;
  assign new_n20381 = new_n20380 ^ new_n20359;
  assign new_n20382 = new_n20367 ^ new_n20354;
  assign new_n20383 = ~new_n20382 & new_n20370;
  assign new_n20384 = new_n20383 ^ new_n20354;
  assign new_n20385 = new_n20381 & new_n20384;
  assign new_n20386 = new_n20385 ^ new_n20377;
  assign new_n20387 = ~new_n20337 & ~new_n20386;
  assign new_n20388 = new_n20383 ^ new_n20370;
  assign new_n20389 = new_n20388 ^ new_n20367;
  assign new_n20390 = new_n20389 ^ new_n20366;
  assign new_n20391 = ~new_n20339 & ~new_n20390;
  assign new_n20392 = new_n20191 ^ new_n20173;
  assign new_n20393 = new_n20345 ^ new_n20340;
  assign new_n20394 = new_n20388 ^ new_n20385;
  assign new_n20395 = new_n20394 ^ new_n20393;
  assign new_n20396 = new_n20395 ^ new_n20392;
  assign new_n20397 = new_n20396 ^ new_n20182;
  assign new_n20398 = new_n20379 ^ new_n20348;
  assign new_n20399 = new_n20398 ^ new_n20321;
  assign new_n20400 = new_n20399 ^ new_n20397;
  assign new_n20401 = ~new_n20328 & new_n20400;
  assign new_n20402 = new_n20379 ^ new_n20367;
  assign new_n20403 = new_n20369 ^ new_n20326;
  assign new_n20404 = new_n20403 ^ new_n20402;
  assign new_n20405 = ~new_n20314 & new_n20404;
  assign new_n20406 = new_n20405 ^ new_n20401;
  assign new_n20407 = new_n20406 ^ new_n20391;
  assign new_n20408 = new_n20407 ^ new_n20387;
  assign new_n20409 = new_n20385 ^ new_n20379;
  assign new_n20410 = new_n20409 ^ new_n20343;
  assign new_n20411 = ~new_n20410 & new_n20346;
  assign new_n20412 = new_n20411 ^ new_n20408;
  assign new_n20413 = ~new_n20330 & new_n20400;
  assign new_n20414 = new_n20413 ^ new_n20412;
  assign new_n20415 = new_n20414 ^ new_n20373;
  assign new_n20416 = new_n20367 ^ new_n20178;
  assign new_n20417 = new_n20374 ^ new_n20364;
  assign new_n20418 = new_n20417 ^ new_n20396;
  assign new_n20419 = new_n20418 ^ new_n20416;
  assign new_n20420 = ~new_n20356 & new_n20419;
  assign new_n20421 = ~new_n20362 & new_n20381;
  assign new_n20422 = new_n20421 ^ new_n20420;
  assign new_n20423 = ~new_n20410 & new_n20347;
  assign new_n20424 = ~new_n20215 & new_n20371;
  assign new_n20425 = new_n20388 ^ new_n20353;
  assign new_n20426 = ~new_n20316 & ~new_n20425;
  assign new_n20427 = new_n20426 ^ new_n20424;
  assign new_n20428 = new_n20427 ^ new_n20423;
  assign new_n20429 = new_n20428 ^ new_n20422;
  assign new_n20430 = new_n20429 ^ new_n20415;
  assign new_n20431 = new_n20430 ^ new_n8242;
  assign new_n20432 = new_n20431 ^ new_n20313;
  assign new_n20433 = new_n18439 ^ new_n18430;
  assign new_n20434 = new_n15174 ^ new_n11893;
  assign new_n20435 = new_n20434 ^ new_n18396;
  assign new_n20436 = new_n20435 ^ new_n18425;
  assign new_n20437 = new_n20436 ^ new_n20433;
  assign new_n20438 = new_n18431 ^ new_n18386;
  assign new_n20439 = new_n15126 ^ new_n11885;
  assign new_n20440 = new_n20439 ^ new_n18417;
  assign new_n20441 = new_n20440 ^ new_n18379;
  assign new_n20442 = new_n20441 ^ new_n20438;
  assign new_n20443 = new_n20442 ^ new_n20437;
  assign new_n20444 = new_n18458 ^ new_n18411;
  assign new_n20445 = new_n15206 ^ new_n11847;
  assign new_n20446 = new_n20445 ^ new_n18310;
  assign new_n20447 = new_n20446 ^ new_n18455;
  assign new_n20448 = new_n20447 ^ new_n20444;
  assign new_n20449 = new_n20448 ^ new_n20443;
  assign new_n20450 = new_n15185 ^ new_n11869;
  assign new_n20451 = new_n20450 ^ new_n18411;
  assign new_n20452 = new_n20451 ^ new_n18361;
  assign new_n20453 = new_n18447 ^ new_n18438;
  assign new_n20454 = new_n20453 ^ new_n18433;
  assign new_n20455 = new_n20454 ^ new_n20452;
  assign new_n20456 = new_n20455 ^ new_n20449;
  assign new_n20457 = new_n20448 & new_n20456;
  assign new_n20458 = new_n20457 ^ new_n20455;
  assign new_n20459 = new_n18411 ^ new_n18298;
  assign new_n20460 = new_n20459 ^ new_n18459;
  assign new_n20461 = new_n15090 ^ new_n11859;
  assign new_n20462 = new_n20461 ^ new_n18287;
  assign new_n20463 = new_n20462 ^ new_n18321;
  assign new_n20464 = new_n20463 ^ new_n20460;
  assign new_n20465 = new_n18443 ^ new_n18355;
  assign new_n20466 = new_n20465 ^ new_n18347;
  assign new_n20467 = new_n15035 ^ new_n11853;
  assign new_n20468 = new_n20467 ^ new_n18411;
  assign new_n20469 = new_n20468 ^ new_n18139;
  assign new_n20470 = new_n20469 ^ new_n20466;
  assign new_n20471 = new_n20470 ^ new_n20464;
  assign new_n20472 = new_n15145 ^ new_n11864;
  assign new_n20473 = new_n20472 ^ new_n18392;
  assign new_n20474 = new_n18410 ^ new_n18407;
  assign new_n20475 = new_n20474 ^ new_n18333;
  assign new_n20476 = new_n20475 ^ new_n20473;
  assign new_n20477 = new_n20476 ^ new_n20455;
  assign new_n20478 = new_n20477 ^ new_n20471;
  assign new_n20479 = new_n18367 ^ new_n18138;
  assign new_n20480 = new_n20479 ^ new_n17838;
  assign new_n20481 = new_n13955 ^ new_n11880;
  assign new_n20482 = new_n20481 ^ new_n18299;
  assign new_n20483 = new_n20482 ^ new_n20480;
  assign new_n20484 = new_n20483 ^ new_n20455;
  assign new_n20485 = new_n20476 ^ new_n20464;
  assign new_n20486 = new_n20485 ^ new_n20484;
  assign new_n20487 = new_n20478 & new_n20486;
  assign new_n20488 = new_n20487 ^ new_n20442;
  assign new_n20489 = new_n20488 ^ new_n20458;
  assign new_n20490 = new_n20488 ^ new_n20478;
  assign new_n20491 = new_n20478 ^ new_n20448;
  assign new_n20492 = new_n20464 ^ new_n20449;
  assign new_n20493 = new_n20483 ^ new_n20476;
  assign new_n20494 = new_n20493 ^ new_n20492;
  assign new_n20495 = new_n20491 & new_n20494;
  assign new_n20496 = new_n20483 ^ new_n20471;
  assign new_n20497 = new_n20496 ^ new_n20442;
  assign new_n20498 = new_n20477 & new_n20497;
  assign new_n20499 = new_n20498 ^ new_n20495;
  assign new_n20500 = new_n20455 ^ new_n20437;
  assign new_n20501 = new_n20500 ^ new_n20493;
  assign new_n20502 = new_n20484 & new_n20501;
  assign new_n20503 = new_n20502 ^ new_n20483;
  assign new_n20504 = new_n20503 ^ new_n20499;
  assign new_n20505 = new_n20504 ^ new_n20490;
  assign new_n20506 = ~new_n20449 & ~new_n20464;
  assign new_n20507 = new_n20506 ^ new_n20464;
  assign new_n20508 = new_n20496 ^ new_n20437;
  assign new_n20509 = new_n20485 & new_n20508;
  assign new_n20510 = new_n20509 ^ new_n20507;
  assign new_n20511 = new_n20510 ^ new_n20493;
  assign new_n20512 = new_n20502 ^ new_n20498;
  assign new_n20513 = new_n20470 ^ new_n20437;
  assign new_n20514 = new_n20513 ^ new_n20512;
  assign new_n20515 = new_n20514 ^ new_n20511;
  assign new_n20516 = ~new_n20515 & new_n20505;
  assign new_n20517 = new_n20516 ^ new_n20489;
  assign new_n20518 = new_n20478 ^ new_n20443;
  assign new_n20519 = new_n20493 & new_n20518;
  assign new_n20520 = new_n20519 ^ new_n20498;
  assign new_n20521 = new_n20520 ^ new_n20508;
  assign new_n20522 = new_n20521 ^ new_n20517;
  assign new_n20523 = new_n20476 ^ new_n20449;
  assign new_n20524 = new_n20497 ^ new_n20448;
  assign new_n20525 = new_n20523 & new_n20524;
  assign new_n20526 = new_n20525 ^ new_n20506;
  assign new_n20527 = new_n20519 ^ new_n20502;
  assign new_n20528 = new_n20527 ^ new_n20526;
  assign new_n20529 = ~new_n20528 & new_n20522;
  assign new_n20530 = new_n20525 ^ new_n20509;
  assign new_n20531 = new_n20530 ^ new_n20476;
  assign new_n20532 = new_n20531 ^ new_n20521;
  assign new_n20533 = new_n20532 ^ new_n20529;
  assign new_n20534 = new_n20456 & new_n20533;
  assign new_n20535 = new_n20464 ^ new_n20437;
  assign new_n20536 = new_n20507 ^ new_n20495;
  assign new_n20537 = new_n20476 ^ new_n20437;
  assign new_n20538 = new_n20495 ^ new_n20457;
  assign new_n20539 = new_n20538 ^ new_n20527;
  assign new_n20540 = new_n20539 ^ new_n20537;
  assign new_n20541 = new_n20532 ^ new_n20516;
  assign new_n20542 = new_n20540 & new_n20541;
  assign new_n20543 = new_n20542 ^ new_n20489;
  assign new_n20544 = new_n20543 ^ new_n20521;
  assign new_n20545 = new_n20529 ^ new_n20516;
  assign new_n20546 = ~new_n20545 & new_n20532;
  assign new_n20547 = new_n20546 ^ new_n20516;
  assign new_n20548 = new_n20544 & new_n20547;
  assign new_n20549 = new_n20546 ^ new_n20532;
  assign new_n20550 = new_n20549 ^ new_n20548;
  assign new_n20551 = new_n20550 ^ new_n20536;
  assign new_n20552 = new_n20551 ^ new_n20535;
  assign new_n20553 = new_n20552 ^ new_n20455;
  assign new_n20554 = new_n20542 ^ new_n20509;
  assign new_n20555 = new_n20554 ^ new_n20488;
  assign new_n20556 = new_n20555 ^ new_n20553;
  assign new_n20557 = ~new_n20556 & new_n20501;
  assign new_n20558 = new_n20548 ^ new_n20542;
  assign new_n20559 = new_n20558 ^ new_n20505;
  assign new_n20560 = new_n20508 & new_n20559;
  assign new_n20561 = new_n20549 ^ new_n20529;
  assign new_n20562 = new_n20561 ^ new_n20528;
  assign new_n20563 = ~new_n20562 & new_n20494;
  assign new_n20564 = new_n20542 ^ new_n20529;
  assign new_n20565 = new_n20531 ^ new_n20489;
  assign new_n20566 = new_n20565 ^ new_n20564;
  assign new_n20567 = new_n20477 & new_n20566;
  assign new_n20568 = ~new_n20556 & new_n20484;
  assign new_n20569 = new_n20568 ^ new_n20567;
  assign new_n20570 = new_n20569 ^ new_n20563;
  assign new_n20571 = new_n20548 ^ new_n20540;
  assign new_n20572 = new_n20449 & new_n20571;
  assign new_n20573 = new_n20572 ^ new_n20570;
  assign new_n20574 = new_n20573 ^ new_n20560;
  assign new_n20575 = new_n20574 ^ new_n20557;
  assign new_n20576 = new_n20575 ^ new_n20534;
  assign new_n20577 = new_n20523 & new_n20544;
  assign new_n20578 = new_n20529 ^ new_n20476;
  assign new_n20579 = new_n20525 ^ new_n20457;
  assign new_n20580 = new_n20579 ^ new_n20552;
  assign new_n20581 = new_n20580 ^ new_n20578;
  assign new_n20582 = ~new_n20581 & new_n20518;
  assign new_n20583 = new_n20582 ^ new_n20577;
  assign new_n20584 = new_n20448 & new_n20533;
  assign new_n20585 = new_n20549 ^ new_n20515;
  assign new_n20586 = ~new_n20585 & new_n20478;
  assign new_n20587 = new_n20586 ^ new_n20584;
  assign new_n20588 = new_n20485 & new_n20559;
  assign new_n20589 = new_n20588 ^ new_n20587;
  assign new_n20590 = new_n20589 ^ new_n20583;
  assign new_n20591 = new_n20590 ^ new_n20576;
  assign new_n20592 = new_n20257 & new_n20277;
  assign new_n20593 = new_n20592 ^ new_n20288;
  assign new_n20594 = new_n20282 ^ new_n20245;
  assign new_n20595 = ~new_n20594 & new_n20202;
  assign new_n20596 = new_n20273 ^ new_n20262;
  assign new_n20597 = new_n20218 & new_n20596;
  assign new_n20598 = new_n20597 ^ new_n20595;
  assign new_n20599 = new_n20598 ^ new_n20291;
  assign new_n20600 = new_n20599 ^ new_n20593;
  assign new_n20601 = ~new_n20247 & new_n20596;
  assign new_n20602 = ~new_n20290 & new_n20237;
  assign new_n20603 = new_n20282 ^ new_n20262;
  assign new_n20604 = new_n20603 ^ new_n20261;
  assign new_n20605 = ~new_n20222 & ~new_n20604;
  assign new_n20606 = new_n20605 ^ new_n20309;
  assign new_n20607 = new_n20606 ^ new_n20299;
  assign new_n20608 = new_n20607 ^ new_n20602;
  assign new_n20609 = new_n20608 ^ new_n20297;
  assign new_n20610 = new_n20609 ^ new_n20601;
  assign new_n20611 = new_n20610 ^ new_n20600;
  assign new_n20612 = new_n20611 ^ new_n20591;
  assign new_n20613 = new_n19517 ^ new_n17259;
  assign new_n20614 = new_n17563 ^ new_n15936;
  assign new_n20615 = new_n20614 ^ new_n17252;
  assign new_n20616 = new_n20615 ^ new_n17223;
  assign new_n20617 = new_n20616 ^ new_n20613;
  assign new_n20618 = new_n19465 ^ new_n17259;
  assign new_n20619 = new_n17318 ^ new_n17275;
  assign new_n20620 = new_n17572 ^ new_n15931;
  assign new_n20621 = new_n20620 ^ new_n20619;
  assign new_n20622 = new_n20621 ^ new_n20618;
  assign new_n20623 = new_n20622 ^ new_n20617;
  assign new_n20624 = new_n17580 ^ new_n15941;
  assign new_n20625 = new_n20624 ^ new_n17146;
  assign new_n20626 = new_n17304 ^ new_n17301;
  assign new_n20627 = new_n20626 ^ new_n19519;
  assign new_n20628 = new_n20627 ^ new_n20625;
  assign new_n20629 = new_n20628 ^ new_n20623;
  assign new_n20630 = new_n19480 ^ new_n17223;
  assign new_n20631 = new_n17567 ^ new_n15970;
  assign new_n20632 = new_n20631 ^ new_n17283;
  assign new_n20633 = new_n20632 ^ new_n17247;
  assign new_n20634 = new_n20633 ^ new_n20630;
  assign new_n20635 = new_n20634 ^ new_n20629;
  assign new_n20636 = new_n20634 ^ new_n20622;
  assign new_n20637 = new_n19519 ^ new_n19473;
  assign new_n20638 = new_n17541 ^ new_n15949;
  assign new_n20639 = new_n20638 ^ new_n17177;
  assign new_n20640 = new_n20639 ^ new_n19496;
  assign new_n20641 = new_n20640 ^ new_n20637;
  assign new_n20642 = new_n17199 ^ new_n16967;
  assign new_n20643 = new_n20642 ^ new_n16654;
  assign new_n20644 = new_n17524 ^ new_n15962;
  assign new_n20645 = new_n20644 ^ new_n19519;
  assign new_n20646 = new_n20645 ^ new_n19509;
  assign new_n20647 = new_n20646 ^ new_n20643;
  assign new_n20648 = new_n20647 ^ new_n20641;
  assign new_n20649 = new_n17575 ^ new_n15923;
  assign new_n20650 = new_n20649 ^ new_n19519;
  assign new_n20651 = new_n20650 ^ new_n19499;
  assign new_n20652 = new_n17318 ^ new_n17199;
  assign new_n20653 = new_n20652 ^ new_n17212;
  assign new_n20654 = new_n20653 ^ new_n20651;
  assign new_n20655 = new_n20654 ^ new_n20634;
  assign new_n20656 = new_n20655 ^ new_n20648;
  assign new_n20657 = new_n20656 ^ new_n20628;
  assign new_n20658 = new_n20641 ^ new_n20629;
  assign new_n20659 = new_n17555 ^ new_n15956;
  assign new_n20660 = new_n20659 ^ new_n16967;
  assign new_n20661 = new_n20660 ^ new_n16663;
  assign new_n20662 = new_n19482 ^ new_n17177;
  assign new_n20663 = new_n20662 ^ new_n20661;
  assign new_n20664 = new_n20663 ^ new_n20634;
  assign new_n20665 = new_n20664 ^ new_n20658;
  assign new_n20666 = new_n20657 & new_n20665;
  assign new_n20667 = new_n20654 ^ new_n20629;
  assign new_n20668 = new_n20628 & new_n20667;
  assign new_n20669 = new_n20668 ^ new_n20666;
  assign new_n20670 = new_n20654 ^ new_n20622;
  assign new_n20671 = new_n20670 ^ new_n20664;
  assign new_n20672 = new_n20663 ^ new_n20654;
  assign new_n20673 = new_n20671 & new_n20672;
  assign new_n20674 = new_n20656 ^ new_n20623;
  assign new_n20675 = new_n20664 & new_n20674;
  assign new_n20676 = new_n20675 ^ new_n20673;
  assign new_n20677 = new_n20676 ^ new_n20669;
  assign new_n20678 = new_n20677 ^ new_n20636;
  assign new_n20679 = new_n20654 ^ new_n20641;
  assign new_n20680 = new_n20679 ^ new_n20664;
  assign new_n20681 = new_n20656 & new_n20680;
  assign new_n20682 = new_n20681 ^ new_n20617;
  assign new_n20683 = new_n20682 ^ new_n20656;
  assign new_n20684 = new_n20663 ^ new_n20648;
  assign new_n20685 = new_n20684 ^ new_n20617;
  assign new_n20686 = new_n20655 & new_n20685;
  assign new_n20687 = new_n20686 ^ new_n20666;
  assign new_n20688 = new_n20673 ^ new_n20663;
  assign new_n20689 = new_n20688 ^ new_n20687;
  assign new_n20690 = new_n20689 ^ new_n20683;
  assign new_n20691 = ~new_n20629 & ~new_n20641;
  assign new_n20692 = new_n20691 ^ new_n20641;
  assign new_n20693 = new_n20641 ^ new_n20634;
  assign new_n20694 = new_n20684 ^ new_n20622;
  assign new_n20695 = new_n20693 & new_n20694;
  assign new_n20696 = new_n20695 ^ new_n20692;
  assign new_n20697 = new_n20696 ^ new_n20664;
  assign new_n20698 = new_n20686 ^ new_n20673;
  assign new_n20699 = new_n20647 ^ new_n20622;
  assign new_n20700 = new_n20699 ^ new_n20698;
  assign new_n20701 = new_n20700 ^ new_n20697;
  assign new_n20702 = ~new_n20701 & new_n20690;
  assign new_n20703 = new_n20686 ^ new_n20675;
  assign new_n20704 = new_n20703 ^ new_n20694;
  assign new_n20705 = new_n20685 ^ new_n20628;
  assign new_n20706 = new_n20635 & new_n20705;
  assign new_n20707 = new_n20706 ^ new_n20695;
  assign new_n20708 = new_n20707 ^ new_n20634;
  assign new_n20709 = new_n20708 ^ new_n20704;
  assign new_n20710 = new_n20709 ^ new_n20702;
  assign new_n20711 = new_n20678 & new_n20710;
  assign new_n20712 = new_n20668 ^ new_n20654;
  assign new_n20713 = new_n20712 ^ new_n20682;
  assign new_n20714 = new_n20713 ^ new_n20711;
  assign new_n20715 = new_n20714 ^ new_n20704;
  assign new_n20716 = new_n20635 & new_n20715;
  assign new_n20717 = new_n20713 ^ new_n20702;
  assign new_n20718 = new_n20717 ^ new_n20704;
  assign new_n20719 = new_n20706 ^ new_n20691;
  assign new_n20720 = new_n20719 ^ new_n20676;
  assign new_n20721 = ~new_n20720 & new_n20718;
  assign new_n20722 = new_n20721 ^ new_n20634;
  assign new_n20723 = new_n20706 ^ new_n20668;
  assign new_n20724 = new_n20641 ^ new_n20622;
  assign new_n20725 = new_n20692 ^ new_n20666;
  assign new_n20726 = new_n20721 ^ new_n20702;
  assign new_n20727 = ~new_n20726 & new_n20709;
  assign new_n20728 = new_n20727 ^ new_n20702;
  assign new_n20729 = new_n20715 & new_n20728;
  assign new_n20730 = new_n20727 ^ new_n20709;
  assign new_n20731 = new_n20730 ^ new_n20729;
  assign new_n20732 = new_n20731 ^ new_n20725;
  assign new_n20733 = new_n20732 ^ new_n20724;
  assign new_n20734 = new_n20733 ^ new_n20723;
  assign new_n20735 = new_n20734 ^ new_n20722;
  assign new_n20736 = ~new_n20735 & new_n20674;
  assign new_n20737 = new_n20736 ^ new_n20716;
  assign new_n20738 = new_n20721 ^ new_n20709;
  assign new_n20739 = new_n20628 & new_n20738;
  assign new_n20740 = new_n20730 ^ new_n20701;
  assign new_n20741 = ~new_n20740 & new_n20656;
  assign new_n20742 = new_n20741 ^ new_n20739;
  assign new_n20743 = new_n20729 ^ new_n20711;
  assign new_n20744 = new_n20743 ^ new_n20690;
  assign new_n20745 = new_n20693 & new_n20744;
  assign new_n20746 = new_n20745 ^ new_n20742;
  assign new_n20747 = new_n20746 ^ new_n20737;
  assign new_n20748 = new_n20667 & new_n20738;
  assign new_n20749 = new_n20733 ^ new_n20654;
  assign new_n20750 = new_n20711 ^ new_n20695;
  assign new_n20751 = new_n20750 ^ new_n20682;
  assign new_n20752 = new_n20751 ^ new_n20749;
  assign new_n20753 = ~new_n20752 & new_n20671;
  assign new_n20754 = new_n20694 & new_n20744;
  assign new_n20755 = new_n20730 ^ new_n20721;
  assign new_n20756 = new_n20755 ^ new_n20720;
  assign new_n20757 = ~new_n20756 & new_n20665;
  assign new_n20758 = ~new_n20752 & new_n20672;
  assign new_n20759 = new_n20721 ^ new_n20711;
  assign new_n20760 = new_n20713 ^ new_n20708;
  assign new_n20761 = new_n20760 ^ new_n20759;
  assign new_n20762 = new_n20655 & new_n20761;
  assign new_n20763 = new_n20762 ^ new_n20758;
  assign new_n20764 = new_n20763 ^ new_n20757;
  assign new_n20765 = new_n20729 ^ new_n20678;
  assign new_n20766 = new_n20629 & new_n20765;
  assign new_n20767 = new_n20766 ^ new_n20764;
  assign new_n20768 = new_n20767 ^ new_n20754;
  assign new_n20769 = new_n20768 ^ new_n20753;
  assign new_n20770 = new_n20769 ^ new_n20748;
  assign new_n20771 = new_n20770 ^ new_n20747;
  assign new_n20772 = new_n20771 ^ new_n20612;
  assign new_n20773 = new_n20772 ^ new_n20432;
  assign new_n20774 = new_n20225 & new_n20307;
  assign new_n20775 = ~new_n20594 & new_n20211;
  assign new_n20776 = new_n20775 ^ new_n20774;
  assign new_n20777 = new_n20776 ^ new_n20609;
  assign new_n20778 = new_n20084 & new_n20159;
  assign new_n20779 = new_n20135 ^ new_n20102;
  assign new_n20780 = ~new_n20779 & new_n20073;
  assign new_n20781 = new_n20780 ^ new_n20778;
  assign new_n20782 = new_n20095 & new_n20143;
  assign new_n20783 = new_n20135 ^ new_n20115;
  assign new_n20784 = new_n20783 ^ new_n20114;
  assign new_n20785 = ~new_n20784 & new_n20081;
  assign new_n20786 = new_n20785 ^ new_n20162;
  assign new_n20787 = new_n20786 ^ new_n20152;
  assign new_n20788 = new_n20787 ^ new_n20782;
  assign new_n20789 = new_n20788 ^ new_n20150;
  assign new_n20790 = new_n20789 ^ new_n20781;
  assign new_n20791 = new_n20790 ^ new_n20777;
  assign new_n20792 = ~new_n20363 & new_n20381;
  assign new_n20793 = ~new_n20319 & ~new_n20425;
  assign new_n20794 = new_n20793 ^ new_n20792;
  assign new_n20795 = ~new_n20390 & new_n20336;
  assign new_n20796 = new_n20795 ^ new_n20424;
  assign new_n20797 = new_n20796 ^ new_n20408;
  assign new_n20798 = new_n20797 ^ new_n20794;
  assign new_n20799 = new_n20798 ^ new_n8235;
  assign new_n20800 = new_n20799 ^ new_n20791;
  assign new_n20801 = new_n20110 & new_n20130;
  assign new_n20802 = new_n20801 ^ new_n20141;
  assign new_n20803 = ~new_n20779 & new_n20054;
  assign new_n20804 = new_n20126 ^ new_n20115;
  assign new_n20805 = new_n20060 & new_n20804;
  assign new_n20806 = new_n20805 ^ new_n20803;
  assign new_n20807 = new_n20806 ^ new_n20144;
  assign new_n20808 = new_n20807 ^ new_n20802;
  assign new_n20809 = new_n20062 & new_n20804;
  assign new_n20810 = new_n20809 ^ new_n20789;
  assign new_n20811 = new_n20810 ^ new_n20808;
  assign new_n20812 = new_n20811 ^ new_n20611;
  assign new_n20813 = new_n20812 ^ new_n20800;
  assign new_n20814 = new_n20705 & new_n20715;
  assign new_n20815 = ~new_n20740 & new_n20680;
  assign new_n20816 = new_n20815 ^ new_n20814;
  assign new_n20817 = ~new_n20756 & new_n20657;
  assign new_n20818 = new_n20817 ^ new_n20739;
  assign new_n20819 = new_n20818 ^ new_n20767;
  assign new_n20820 = new_n20819 ^ new_n20816;
  assign new_n20821 = new_n20524 & new_n20544;
  assign new_n20822 = ~new_n20585 & new_n20486;
  assign new_n20823 = new_n20822 ^ new_n20821;
  assign new_n20824 = ~new_n20562 & new_n20491;
  assign new_n20825 = new_n20824 ^ new_n20584;
  assign new_n20826 = new_n20825 ^ new_n20573;
  assign new_n20827 = new_n20826 ^ new_n20823;
  assign new_n20828 = new_n20827 ^ new_n20820;
  assign new_n20829 = new_n20775 ^ new_n20302;
  assign new_n20830 = ~new_n20604 & new_n20219;
  assign new_n20831 = new_n20830 ^ new_n20597;
  assign new_n20832 = new_n20831 ^ new_n20607;
  assign new_n20833 = new_n20832 ^ new_n20829;
  assign new_n20834 = new_n20833 ^ new_n20828;
  assign new_n20835 = new_n20834 ^ new_n20813;
  assign new_n20836 = new_n20791 ^ new_n20312;
  assign new_n20837 = new_n20602 ^ new_n20599;
  assign new_n20838 = new_n20837 ^ new_n20310;
  assign new_n20839 = new_n20807 ^ new_n20782;
  assign new_n20840 = new_n20839 ^ new_n20163;
  assign new_n20841 = new_n20840 ^ new_n20838;
  assign new_n20842 = new_n20841 ^ new_n20836;
  assign new_n20843 = new_n20588 ^ new_n20582;
  assign new_n20844 = new_n20492 & new_n20571;
  assign new_n20845 = new_n20844 ^ new_n20821;
  assign new_n20846 = new_n20845 ^ new_n20569;
  assign new_n20847 = new_n20572 ^ new_n20557;
  assign new_n20848 = new_n20847 ^ new_n20846;
  assign new_n20849 = new_n20848 ^ new_n20843;
  assign new_n20850 = new_n20423 ^ new_n20420;
  assign new_n20851 = new_n20413 ^ new_n20387;
  assign new_n20852 = ~new_n20338 & ~new_n20386;
  assign new_n20853 = new_n20852 ^ new_n20792;
  assign new_n20854 = new_n20853 ^ new_n20406;
  assign new_n20855 = new_n20854 ^ new_n20851;
  assign new_n20856 = new_n20855 ^ new_n20850;
  assign new_n20857 = new_n20856 ^ new_n8233;
  assign new_n20858 = new_n20857 ^ new_n20849;
  assign new_n20859 = new_n20745 ^ new_n20736;
  assign new_n20860 = new_n20766 ^ new_n20753;
  assign new_n20861 = new_n20658 & new_n20765;
  assign new_n20862 = new_n20861 ^ new_n20814;
  assign new_n20863 = new_n20862 ^ new_n20763;
  assign new_n20864 = new_n20863 ^ new_n20860;
  assign new_n20865 = new_n20864 ^ new_n20859;
  assign new_n20866 = new_n20865 ^ new_n20858;
  assign new_n20867 = new_n20866 ^ new_n20842;
  assign new_n20868 = new_n20867 ^ new_n20835;
  assign new_n20869 = new_n20868 ^ new_n20773;
  assign new_n20870 = new_n20497 & new_n20566;
  assign new_n20871 = new_n20870 ^ new_n20557;
  assign new_n20872 = new_n20824 ^ new_n20586;
  assign new_n20873 = new_n20872 ^ new_n20822;
  assign new_n20874 = new_n20873 ^ new_n20570;
  assign new_n20875 = new_n20874 ^ new_n20871;
  assign new_n20876 = new_n20685 & new_n20761;
  assign new_n20877 = new_n20876 ^ new_n20753;
  assign new_n20878 = new_n20817 ^ new_n20741;
  assign new_n20879 = new_n20878 ^ new_n20815;
  assign new_n20880 = new_n20879 ^ new_n20764;
  assign new_n20881 = new_n20880 ^ new_n20877;
  assign new_n20882 = new_n20881 ^ new_n20875;
  assign new_n20883 = new_n20778 ^ new_n20160;
  assign new_n20884 = ~new_n20140 & new_n20080;
  assign new_n20885 = new_n20884 ^ new_n20808;
  assign new_n20886 = new_n20885 ^ new_n20883;
  assign new_n20887 = new_n20886 ^ new_n20882;
  assign new_n20888 = new_n20774 ^ new_n20297;
  assign new_n20889 = new_n20830 ^ new_n20595;
  assign new_n20890 = new_n20889 ^ new_n20775;
  assign new_n20891 = new_n20890 ^ new_n20606;
  assign new_n20892 = new_n20891 ^ new_n20888;
  assign new_n20893 = new_n20333 & new_n20404;
  assign new_n20894 = new_n20893 ^ new_n20413;
  assign new_n20895 = new_n20795 ^ new_n20426;
  assign new_n20896 = new_n20895 ^ new_n20793;
  assign new_n20897 = new_n20896 ^ new_n20407;
  assign new_n20898 = new_n20897 ^ new_n20894;
  assign new_n20899 = new_n20898 ^ new_n8225;
  assign new_n20900 = new_n20899 ^ new_n20892;
  assign new_n20901 = new_n20774 ^ new_n20308;
  assign new_n20902 = new_n20210 & new_n20287;
  assign new_n20903 = new_n20902 ^ new_n20600;
  assign new_n20904 = new_n20903 ^ new_n20901;
  assign new_n20905 = new_n20904 ^ new_n20900;
  assign new_n20906 = new_n20905 ^ new_n20887;
  assign new_n20907 = new_n20906 ^ new_n20869;
  assign new_n20908 = new_n20870 ^ new_n20567;
  assign new_n20909 = ~new_n20581 & new_n20493;
  assign new_n20910 = new_n20909 ^ new_n20590;
  assign new_n20911 = new_n20910 ^ new_n20908;
  assign new_n20912 = new_n20876 ^ new_n20762;
  assign new_n20913 = ~new_n20735 & new_n20664;
  assign new_n20914 = new_n20913 ^ new_n20747;
  assign new_n20915 = new_n20914 ^ new_n20912;
  assign new_n20916 = new_n20915 ^ new_n20911;
  assign new_n20917 = new_n20916 ^ new_n20904;
  assign new_n20918 = ~new_n20784 & new_n20078;
  assign new_n20919 = new_n20918 ^ new_n20803;
  assign new_n20920 = new_n20919 ^ new_n20780;
  assign new_n20921 = new_n20920 ^ new_n20788;
  assign new_n20922 = new_n20890 ^ new_n20608;
  assign new_n20923 = new_n20922 ^ new_n20921;
  assign new_n20924 = new_n20893 ^ new_n20405;
  assign new_n20925 = new_n20318 & new_n20419;
  assign new_n20926 = new_n20925 ^ new_n20429;
  assign new_n20927 = new_n20926 ^ new_n20924;
  assign new_n20928 = new_n20927 ^ new_n8227;
  assign new_n20929 = new_n20928 ^ new_n20923;
  assign new_n20930 = new_n20929 ^ new_n20917;
  assign new_n20931 = new_n20930 ^ new_n20906;
  assign new_n20932 = new_n20838 ^ new_n20791;
  assign new_n20933 = new_n20589 ^ new_n20560;
  assign new_n20934 = new_n20933 ^ new_n20846;
  assign new_n20935 = new_n20428 ^ new_n20411;
  assign new_n20936 = new_n20935 ^ new_n20854;
  assign new_n20937 = new_n20936 ^ new_n8229;
  assign new_n20938 = new_n20937 ^ new_n20934;
  assign new_n20939 = new_n20754 ^ new_n20746;
  assign new_n20940 = new_n20939 ^ new_n20863;
  assign new_n20941 = new_n20940 ^ new_n20938;
  assign new_n20942 = new_n20941 ^ new_n20932;
  assign new_n20943 = new_n20942 ^ new_n20931;
  assign new_n20944 = new_n20867 & new_n20943;
  assign new_n20945 = new_n20944 ^ new_n20867;
  assign new_n20946 = new_n20930 ^ new_n20869;
  assign new_n20947 = new_n20876 ^ new_n20815;
  assign new_n20948 = new_n20947 ^ new_n20769;
  assign new_n20949 = new_n20870 ^ new_n20822;
  assign new_n20950 = new_n20949 ^ new_n20575;
  assign new_n20951 = new_n20950 ^ new_n20948;
  assign new_n20952 = new_n20778 ^ new_n20150;
  assign new_n20953 = new_n20920 ^ new_n20786;
  assign new_n20954 = new_n20953 ^ new_n20952;
  assign new_n20955 = new_n20954 ^ new_n20951;
  assign new_n20956 = new_n20893 ^ new_n20793;
  assign new_n20957 = new_n20956 ^ new_n20414;
  assign new_n20958 = new_n20957 ^ new_n8231;
  assign new_n20959 = new_n20958 ^ new_n20777;
  assign new_n20960 = new_n20959 ^ new_n20892;
  assign new_n20961 = new_n20960 ^ new_n20955;
  assign new_n20962 = new_n20961 ^ new_n20867;
  assign new_n20963 = ~new_n20962 & new_n20946;
  assign new_n20964 = new_n20963 ^ new_n20945;
  assign new_n20965 = new_n20961 ^ new_n20773;
  assign new_n20966 = new_n20965 ^ new_n20964;
  assign new_n20967 = new_n20873 ^ new_n20574;
  assign new_n20968 = new_n20879 ^ new_n20768;
  assign new_n20969 = new_n20968 ^ new_n20967;
  assign new_n20970 = new_n20969 ^ new_n20791;
  assign new_n20971 = new_n20896 ^ new_n20412;
  assign new_n20972 = new_n20971 ^ new_n8238;
  assign new_n20973 = new_n20972 ^ new_n20922;
  assign new_n20974 = new_n20780 ^ new_n20155;
  assign new_n20975 = new_n20918 ^ new_n20805;
  assign new_n20976 = new_n20975 ^ new_n20787;
  assign new_n20977 = new_n20976 ^ new_n20974;
  assign new_n20978 = new_n20977 ^ new_n20833;
  assign new_n20979 = new_n20978 ^ new_n20973;
  assign new_n20980 = new_n20979 ^ new_n20970;
  assign new_n20981 = new_n20980 ^ new_n20930;
  assign new_n20982 = new_n20981 ^ new_n20965;
  assign new_n20983 = new_n20980 ^ new_n20773;
  assign new_n20984 = ~new_n20982 & new_n20983;
  assign new_n20985 = new_n20980 ^ new_n20961;
  assign new_n20986 = new_n20907 & new_n20985;
  assign new_n20987 = new_n20986 ^ new_n20984;
  assign new_n20988 = new_n20930 ^ new_n20835;
  assign new_n20989 = new_n20988 ^ new_n20987;
  assign new_n20990 = new_n20989 ^ new_n20966;
  assign new_n20991 = new_n20985 ^ new_n20868;
  assign new_n20992 = new_n20980 ^ new_n20867;
  assign new_n20993 = new_n20992 ^ new_n20965;
  assign new_n20994 = ~new_n20991 & ~new_n20993;
  assign new_n20995 = new_n20994 ^ new_n20906;
  assign new_n20996 = new_n20995 ^ new_n20991;
  assign new_n20997 = new_n20991 ^ new_n20942;
  assign new_n20998 = new_n20943 ^ new_n20867;
  assign new_n20999 = new_n20998 ^ new_n20965;
  assign new_n21000 = new_n20997 & new_n20999;
  assign new_n21001 = new_n21000 ^ new_n20986;
  assign new_n21002 = new_n20984 ^ new_n20773;
  assign new_n21003 = new_n21002 ^ new_n21001;
  assign new_n21004 = new_n21003 ^ new_n20996;
  assign new_n21005 = ~new_n20990 & new_n21004;
  assign new_n21006 = new_n20961 ^ new_n20943;
  assign new_n21007 = new_n20942 ^ new_n20907;
  assign new_n21008 = ~new_n21006 & ~new_n21007;
  assign new_n21009 = new_n21008 ^ new_n20963;
  assign new_n21010 = new_n21009 ^ new_n20961;
  assign new_n21011 = new_n20991 ^ new_n20931;
  assign new_n21012 = ~new_n21011 & new_n20965;
  assign new_n21013 = new_n21012 ^ new_n20986;
  assign new_n21014 = new_n21013 ^ new_n20946;
  assign new_n21015 = new_n21014 ^ new_n21010;
  assign new_n21016 = new_n21015 ^ new_n21005;
  assign new_n21017 = new_n20961 ^ new_n20930;
  assign new_n21018 = new_n20980 ^ new_n20943;
  assign new_n21019 = ~new_n20942 & ~new_n21018;
  assign new_n21020 = new_n21019 ^ new_n21000;
  assign new_n21021 = new_n21012 ^ new_n20984;
  assign new_n21022 = new_n21021 ^ new_n21020;
  assign new_n21023 = new_n21022 ^ new_n21017;
  assign new_n21024 = ~new_n21023 & new_n21016;
  assign new_n21025 = new_n21019 ^ new_n20980;
  assign new_n21026 = new_n21025 ^ new_n20995;
  assign new_n21027 = new_n21026 ^ new_n21005;
  assign new_n21028 = new_n21027 ^ new_n21014;
  assign new_n21029 = new_n21008 ^ new_n20944;
  assign new_n21030 = new_n21029 ^ new_n21021;
  assign new_n21031 = ~new_n21028 & ~new_n21030;
  assign new_n21032 = new_n21031 ^ new_n21024;
  assign new_n21033 = new_n21026 ^ new_n21010;
  assign new_n21034 = new_n21033 ^ new_n21032;
  assign new_n21035 = ~new_n21034 & new_n20907;
  assign new_n21036 = new_n21031 ^ new_n21005;
  assign new_n21037 = ~new_n21015 & ~new_n21036;
  assign new_n21038 = new_n21037 ^ new_n21031;
  assign new_n21039 = new_n21038 ^ new_n21016;
  assign new_n21040 = new_n21039 ^ new_n20990;
  assign new_n21041 = ~new_n20993 & new_n21040;
  assign new_n21042 = new_n21041 ^ new_n21035;
  assign new_n21043 = new_n20930 ^ new_n20867;
  assign new_n21044 = new_n21000 ^ new_n20945;
  assign new_n21045 = new_n21026 ^ new_n21024;
  assign new_n21046 = new_n21045 ^ new_n21014;
  assign new_n21047 = ~new_n21038 & ~new_n21046;
  assign new_n21048 = new_n21047 ^ new_n21039;
  assign new_n21049 = new_n21048 ^ new_n21044;
  assign new_n21050 = new_n21049 ^ new_n21043;
  assign new_n21051 = new_n21050 ^ new_n20980;
  assign new_n21052 = new_n21024 ^ new_n20963;
  assign new_n21053 = new_n21052 ^ new_n20995;
  assign new_n21054 = new_n21053 ^ new_n21051;
  assign new_n21055 = ~new_n20982 & new_n21054;
  assign new_n21056 = new_n21047 ^ new_n21024;
  assign new_n21057 = new_n21056 ^ new_n21004;
  assign new_n21058 = new_n20946 & new_n21057;
  assign new_n21059 = new_n21047 ^ new_n21023;
  assign new_n21060 = ~new_n20943 & ~new_n21059;
  assign new_n21061 = ~new_n21034 & new_n20985;
  assign new_n21062 = new_n20983 & new_n21054;
  assign new_n21063 = new_n21062 ^ new_n21061;
  assign new_n21064 = new_n21039 ^ new_n21031;
  assign new_n21065 = new_n21064 ^ new_n21030;
  assign new_n21066 = new_n20999 & new_n21065;
  assign new_n21067 = new_n21066 ^ new_n21063;
  assign new_n21068 = new_n21067 ^ new_n21060;
  assign new_n21069 = new_n21068 ^ new_n21058;
  assign new_n21070 = new_n21069 ^ new_n21055;
  assign new_n21071 = new_n21070 ^ new_n21042;
  assign new_n21072 = new_n21071 ^ new_n20011;
  assign new_n21073 = new_n21072 ^ new_n20000;
  assign new_n21074 = new_n18765 ^ new_n8547;
  assign new_n21075 = new_n18718 ^ new_n8542;
  assign new_n21076 = new_n21075 ^ new_n21074;
  assign new_n21077 = new_n17678 ^ new_n8572;
  assign new_n21078 = new_n18771 ^ new_n8533;
  assign new_n21079 = new_n21078 ^ new_n21077;
  assign new_n21080 = new_n18634 ^ new_n8564;
  assign new_n21081 = new_n18793 ^ new_n8581;
  assign new_n21082 = new_n21081 ^ new_n21080;
  assign new_n21083 = new_n21082 ^ new_n21079;
  assign new_n21084 = new_n21083 ^ new_n21076;
  assign new_n21085 = new_n18823 ^ new_n8553;
  assign new_n21086 = new_n21085 ^ new_n21076;
  assign new_n21087 = new_n21086 ^ new_n21078;
  assign new_n21088 = ~new_n21087 & new_n21085;
  assign new_n21089 = new_n21088 ^ new_n21078;
  assign new_n21090 = new_n21080 ^ new_n21078;
  assign new_n21091 = new_n18670 ^ new_n8589;
  assign new_n21092 = new_n21091 ^ new_n21077;
  assign new_n21093 = new_n21092 ^ new_n21090;
  assign new_n21094 = ~new_n21083 & ~new_n21093;
  assign new_n21095 = new_n21094 ^ new_n21074;
  assign new_n21096 = new_n21095 ^ new_n21089;
  assign new_n21097 = new_n21095 ^ new_n21083;
  assign new_n21098 = new_n21078 ^ new_n21075;
  assign new_n21099 = new_n21098 ^ new_n21092;
  assign new_n21100 = new_n21091 ^ new_n21078;
  assign new_n21101 = ~new_n21099 & new_n21100;
  assign new_n21102 = new_n21091 ^ new_n21082;
  assign new_n21103 = new_n21102 ^ new_n21074;
  assign new_n21104 = ~new_n21103 & new_n21079;
  assign new_n21105 = new_n21104 ^ new_n21101;
  assign new_n21106 = new_n21085 ^ new_n21083;
  assign new_n21107 = new_n21086 ^ new_n21080;
  assign new_n21108 = new_n21107 ^ new_n21092;
  assign new_n21109 = ~new_n21106 & new_n21108;
  assign new_n21110 = new_n21109 ^ new_n21091;
  assign new_n21111 = new_n21110 ^ new_n21105;
  assign new_n21112 = new_n21111 ^ new_n21097;
  assign new_n21113 = new_n21080 & new_n21086;
  assign new_n21114 = new_n21113 ^ new_n21080;
  assign new_n21115 = new_n21102 ^ new_n21075;
  assign new_n21116 = new_n21080 ^ new_n21077;
  assign new_n21117 = ~new_n21116 & new_n21115;
  assign new_n21118 = new_n21117 ^ new_n21114;
  assign new_n21119 = new_n21118 ^ new_n21092;
  assign new_n21120 = new_n21081 ^ new_n21075;
  assign new_n21121 = new_n21120 ^ new_n21105;
  assign new_n21122 = new_n21121 ^ new_n21119;
  assign new_n21123 = ~new_n21112 & ~new_n21122;
  assign new_n21124 = new_n21123 ^ new_n21096;
  assign new_n21125 = new_n21084 & new_n21092;
  assign new_n21126 = new_n21125 ^ new_n21104;
  assign new_n21127 = new_n21126 ^ new_n21115;
  assign new_n21128 = new_n21127 ^ new_n21124;
  assign new_n21129 = new_n21086 ^ new_n21077;
  assign new_n21130 = new_n21103 ^ new_n21085;
  assign new_n21131 = ~new_n21129 & ~new_n21130;
  assign new_n21132 = new_n21131 ^ new_n21113;
  assign new_n21133 = new_n21125 ^ new_n21101;
  assign new_n21134 = new_n21133 ^ new_n21132;
  assign new_n21135 = ~new_n21134 & new_n21128;
  assign new_n21136 = new_n21135 ^ new_n21077;
  assign new_n21137 = new_n21131 ^ new_n21088;
  assign new_n21138 = new_n21080 ^ new_n21075;
  assign new_n21139 = new_n21114 ^ new_n21109;
  assign new_n21140 = new_n21131 ^ new_n21117;
  assign new_n21141 = new_n21140 ^ new_n21077;
  assign new_n21142 = new_n21141 ^ new_n21127;
  assign new_n21143 = new_n21135 ^ new_n21123;
  assign new_n21144 = ~new_n21142 & ~new_n21143;
  assign new_n21145 = new_n21144 ^ new_n21135;
  assign new_n21146 = new_n21142 ^ new_n21123;
  assign new_n21147 = new_n21077 ^ new_n21075;
  assign new_n21148 = new_n21109 ^ new_n21088;
  assign new_n21149 = new_n21148 ^ new_n21133;
  assign new_n21150 = new_n21149 ^ new_n21147;
  assign new_n21151 = ~new_n21150 & new_n21146;
  assign new_n21152 = new_n21151 ^ new_n21096;
  assign new_n21153 = new_n21152 ^ new_n21127;
  assign new_n21154 = ~new_n21145 & new_n21153;
  assign new_n21155 = new_n21146 ^ new_n21145;
  assign new_n21156 = new_n21155 ^ new_n21154;
  assign new_n21157 = new_n21156 ^ new_n21139;
  assign new_n21158 = new_n21157 ^ new_n21138;
  assign new_n21159 = new_n21158 ^ new_n21137;
  assign new_n21160 = new_n21159 ^ new_n21136;
  assign new_n21161 = ~new_n21160 & new_n21084;
  assign new_n21162 = new_n21154 ^ new_n21151;
  assign new_n21163 = new_n21162 ^ new_n21112;
  assign new_n21164 = ~new_n21116 & ~new_n21163;
  assign new_n21165 = new_n21164 ^ new_n21161;
  assign new_n21166 = new_n21158 ^ new_n21078;
  assign new_n21167 = new_n21151 ^ new_n21117;
  assign new_n21168 = new_n21167 ^ new_n21095;
  assign new_n21169 = new_n21168 ^ new_n21166;
  assign new_n21170 = ~new_n21099 & ~new_n21169;
  assign new_n21171 = new_n21154 ^ new_n21150;
  assign new_n21172 = ~new_n21086 & ~new_n21171;
  assign new_n21173 = new_n21172 ^ new_n21170;
  assign new_n21174 = ~new_n21171 & new_n21107;
  assign new_n21175 = ~new_n21130 & new_n21153;
  assign new_n21176 = new_n21175 ^ new_n21174;
  assign new_n21177 = new_n21151 ^ new_n21135;
  assign new_n21178 = new_n21141 ^ new_n21096;
  assign new_n21179 = new_n21178 ^ new_n21177;
  assign new_n21180 = new_n21079 & new_n21179;
  assign new_n21181 = ~new_n21169 & new_n21100;
  assign new_n21182 = new_n21181 ^ new_n21180;
  assign new_n21183 = new_n21182 ^ new_n21176;
  assign new_n21184 = new_n21183 ^ new_n21173;
  assign new_n21185 = new_n21184 ^ new_n21165;
  assign new_n21186 = new_n20856 ^ new_n19487;
  assign new_n21187 = new_n21186 ^ new_n21185;
  assign new_n21188 = ~new_n21059 & new_n20998;
  assign new_n21189 = ~new_n21007 & ~new_n21046;
  assign new_n21190 = new_n21189 ^ new_n21188;
  assign new_n21191 = new_n21190 ^ new_n21063;
  assign new_n21192 = ~new_n20962 & new_n21057;
  assign new_n21193 = ~new_n20991 & new_n21040;
  assign new_n21194 = new_n21031 ^ new_n21015;
  assign new_n21195 = ~new_n20942 & new_n21194;
  assign new_n21196 = new_n21195 ^ new_n21193;
  assign new_n21197 = new_n21196 ^ new_n21192;
  assign new_n21198 = new_n21197 ^ new_n21058;
  assign new_n21199 = new_n21198 ^ new_n21191;
  assign new_n21200 = new_n21199 ^ new_n21187;
  assign new_n21201 = new_n16149 ^ new_n16131;
  assign new_n21202 = new_n21201 ^ new_n15733;
  assign new_n21203 = new_n21202 ^ new_n16210;
  assign new_n21204 = new_n16254 ^ new_n16233;
  assign new_n21205 = new_n16263 ^ new_n16233;
  assign new_n21206 = new_n21205 ^ new_n21201;
  assign new_n21207 = new_n21206 ^ new_n16279;
  assign new_n21208 = new_n16254 ^ new_n16210;
  assign new_n21209 = new_n21208 ^ new_n16279;
  assign new_n21210 = new_n21209 ^ new_n16131;
  assign new_n21211 = new_n16233 ^ new_n15733;
  assign new_n21212 = new_n21211 ^ new_n21210;
  assign new_n21213 = new_n21207 & new_n21212;
  assign new_n21214 = new_n21209 ^ new_n16263;
  assign new_n21215 = new_n16279 & new_n21214;
  assign new_n21216 = new_n21215 ^ new_n21213;
  assign new_n21217 = new_n21208 ^ new_n21206;
  assign new_n21218 = new_n21211 & new_n21217;
  assign new_n21219 = new_n16263 ^ new_n15733;
  assign new_n21220 = new_n16263 ^ new_n16254;
  assign new_n21221 = new_n21220 ^ new_n21211;
  assign new_n21222 = new_n21219 & new_n21221;
  assign new_n21223 = new_n21222 ^ new_n21218;
  assign new_n21224 = new_n21223 ^ new_n21216;
  assign new_n21225 = new_n21224 ^ new_n21204;
  assign new_n21226 = new_n21209 ^ new_n16233;
  assign new_n21227 = new_n21203 ^ new_n16279;
  assign new_n21228 = new_n21226 & new_n21227;
  assign new_n21229 = new_n21202 ^ new_n16254;
  assign new_n21230 = new_n16233 ^ new_n16131;
  assign new_n21231 = new_n21229 & new_n21230;
  assign new_n21232 = new_n21231 ^ new_n21228;
  assign new_n21233 = new_n21232 ^ new_n16233;
  assign new_n21234 = new_n21203 & new_n21205;
  assign new_n21235 = new_n21234 ^ new_n21218;
  assign new_n21236 = new_n21235 ^ new_n21229;
  assign new_n21237 = new_n21236 ^ new_n21233;
  assign new_n21238 = new_n16263 ^ new_n16131;
  assign new_n21239 = new_n21238 ^ new_n21211;
  assign new_n21240 = new_n21206 & new_n21239;
  assign new_n21241 = new_n21240 ^ new_n16210;
  assign new_n21242 = new_n21241 ^ new_n21206;
  assign new_n21243 = new_n21234 ^ new_n21222;
  assign new_n21244 = new_n21213 ^ new_n15733;
  assign new_n21245 = new_n21244 ^ new_n21243;
  assign new_n21246 = new_n21245 ^ new_n21242;
  assign new_n21247 = ~new_n16131 & ~new_n21209;
  assign new_n21248 = new_n21247 ^ new_n16131;
  assign new_n21249 = new_n21248 ^ new_n21231;
  assign new_n21250 = new_n21249 ^ new_n21211;
  assign new_n21251 = new_n16254 ^ new_n16149;
  assign new_n21252 = new_n21251 ^ new_n21243;
  assign new_n21253 = new_n21252 ^ new_n21250;
  assign new_n21254 = ~new_n21253 & new_n21246;
  assign new_n21255 = new_n21254 ^ new_n21237;
  assign new_n21256 = new_n21225 & new_n21255;
  assign new_n21257 = new_n21215 ^ new_n16263;
  assign new_n21258 = new_n21257 ^ new_n21241;
  assign new_n21259 = new_n21258 ^ new_n21254;
  assign new_n21260 = new_n21259 ^ new_n21236;
  assign new_n21261 = new_n21247 ^ new_n21228;
  assign new_n21262 = new_n21261 ^ new_n21223;
  assign new_n21263 = ~new_n21262 & new_n21260;
  assign new_n21264 = new_n21263 ^ new_n21256;
  assign new_n21265 = new_n21258 ^ new_n21233;
  assign new_n21266 = new_n21265 ^ new_n21264;
  assign new_n21267 = new_n21203 & new_n21266;
  assign new_n21268 = new_n21263 ^ new_n21254;
  assign new_n21269 = ~new_n21268 & new_n21237;
  assign new_n21270 = new_n21269 ^ new_n21237;
  assign new_n21271 = new_n21270 ^ new_n21253;
  assign new_n21272 = ~new_n21271 & new_n21239;
  assign new_n21273 = new_n21272 ^ new_n21267;
  assign new_n21274 = new_n21258 ^ new_n21256;
  assign new_n21275 = new_n21274 ^ new_n21236;
  assign new_n21276 = new_n21269 ^ new_n21254;
  assign new_n21277 = new_n21275 & new_n21276;
  assign new_n21278 = new_n21277 ^ new_n21225;
  assign new_n21279 = new_n21209 & new_n21278;
  assign new_n21280 = new_n21270 ^ new_n21263;
  assign new_n21281 = new_n21280 ^ new_n21262;
  assign new_n21282 = ~new_n21281 & new_n21212;
  assign new_n21283 = new_n21205 & new_n21266;
  assign new_n21284 = new_n16254 ^ new_n16131;
  assign new_n21285 = new_n21248 ^ new_n21213;
  assign new_n21286 = new_n21277 ^ new_n21270;
  assign new_n21287 = new_n21286 ^ new_n21285;
  assign new_n21288 = new_n21287 ^ new_n21284;
  assign new_n21289 = new_n21288 ^ new_n16263;
  assign new_n21290 = new_n21256 ^ new_n21231;
  assign new_n21291 = new_n21290 ^ new_n21241;
  assign new_n21292 = new_n21291 ^ new_n21289;
  assign new_n21293 = ~new_n21292 & new_n21219;
  assign new_n21294 = new_n21293 ^ new_n21283;
  assign new_n21295 = new_n21294 ^ new_n21282;
  assign new_n21296 = new_n21295 ^ new_n21279;
  assign new_n21297 = new_n21277 ^ new_n21256;
  assign new_n21298 = new_n21297 ^ new_n21246;
  assign new_n21299 = new_n21229 & new_n21298;
  assign new_n21300 = new_n21299 ^ new_n21296;
  assign new_n21301 = ~new_n21292 & new_n21221;
  assign new_n21302 = new_n21301 ^ new_n21300;
  assign new_n21303 = new_n21302 ^ new_n21273;
  assign new_n21304 = new_n21303 ^ new_n15145;
  assign new_n21305 = new_n21304 ^ new_n10832;
  assign new_n21306 = new_n14901 ^ new_n13955;
  assign new_n21307 = new_n21306 ^ new_n16654;
  assign new_n21308 = new_n21307 ^ new_n17155;
  assign new_n21309 = new_n21308 ^ new_n20662;
  assign new_n21310 = new_n17284 ^ new_n17156;
  assign new_n21311 = new_n15090 ^ new_n14792;
  assign new_n21312 = new_n21311 ^ new_n16809;
  assign new_n21313 = new_n21312 ^ new_n20626;
  assign new_n21314 = new_n21313 ^ new_n21310;
  assign new_n21315 = new_n15035 ^ new_n14810;
  assign new_n21316 = new_n21315 ^ new_n17212;
  assign new_n21317 = new_n21316 ^ new_n17284;
  assign new_n21318 = new_n19509 ^ new_n17119;
  assign new_n21319 = new_n21318 ^ new_n21317;
  assign new_n21320 = new_n21319 ^ new_n21314;
  assign new_n21321 = new_n21320 ^ new_n21309;
  assign new_n21322 = new_n15126 ^ new_n14098;
  assign new_n21323 = new_n21322 ^ new_n17247;
  assign new_n21324 = new_n19517 ^ new_n17264;
  assign new_n21325 = new_n21324 ^ new_n21323;
  assign new_n21326 = new_n21325 ^ new_n21321;
  assign new_n21327 = new_n15145 ^ new_n14858;
  assign new_n21328 = new_n21327 ^ new_n17125;
  assign new_n21329 = new_n19480 ^ new_n17230;
  assign new_n21330 = new_n21329 ^ new_n21328;
  assign new_n21331 = new_n19499 ^ new_n17200;
  assign new_n21332 = new_n15185 ^ new_n14849;
  assign new_n21333 = new_n21332 ^ new_n17275;
  assign new_n21334 = new_n21333 ^ new_n17284;
  assign new_n21335 = new_n21334 ^ new_n21331;
  assign new_n21336 = new_n21335 ^ new_n21330;
  assign new_n21337 = new_n21336 ^ new_n21320;
  assign new_n21338 = new_n21330 ^ new_n21309;
  assign new_n21339 = new_n21335 ^ new_n21314;
  assign new_n21340 = new_n21339 ^ new_n21338;
  assign new_n21341 = new_n21337 & new_n21340;
  assign new_n21342 = new_n21341 ^ new_n21325;
  assign new_n21343 = new_n21342 ^ new_n21337;
  assign new_n21344 = new_n21326 & new_n21336;
  assign new_n21345 = new_n15206 ^ new_n14878;
  assign new_n21346 = new_n21345 ^ new_n17146;
  assign new_n21347 = new_n17305 ^ new_n17284;
  assign new_n21348 = new_n21347 ^ new_n21346;
  assign new_n21349 = new_n21348 ^ new_n21337;
  assign new_n21350 = new_n15174 ^ new_n14676;
  assign new_n21351 = new_n21350 ^ new_n17252;
  assign new_n21352 = new_n19465 ^ new_n17319;
  assign new_n21353 = new_n21352 ^ new_n21351;
  assign new_n21354 = new_n21353 ^ new_n21325;
  assign new_n21355 = new_n21354 ^ new_n21348;
  assign new_n21356 = new_n21355 ^ new_n21314;
  assign new_n21357 = new_n21356 ^ new_n21338;
  assign new_n21358 = new_n21349 & new_n21357;
  assign new_n21359 = new_n21358 ^ new_n21344;
  assign new_n21360 = new_n21353 ^ new_n21335;
  assign new_n21361 = new_n21360 ^ new_n21338;
  assign new_n21362 = new_n21335 ^ new_n21309;
  assign new_n21363 = new_n21361 & new_n21362;
  assign new_n21364 = new_n21363 ^ new_n21309;
  assign new_n21365 = new_n21364 ^ new_n21359;
  assign new_n21366 = new_n21365 ^ new_n21343;
  assign new_n21367 = new_n21353 ^ new_n21321;
  assign new_n21368 = new_n21330 ^ new_n21314;
  assign new_n21369 = new_n21367 & new_n21368;
  assign new_n21370 = ~new_n21314 & ~new_n21355;
  assign new_n21371 = new_n21370 ^ new_n21314;
  assign new_n21372 = new_n21371 ^ new_n21369;
  assign new_n21373 = new_n21372 ^ new_n21338;
  assign new_n21374 = new_n21363 ^ new_n21344;
  assign new_n21375 = new_n21353 ^ new_n21319;
  assign new_n21376 = new_n21375 ^ new_n21374;
  assign new_n21377 = new_n21376 ^ new_n21373;
  assign new_n21378 = ~new_n21377 & new_n21366;
  assign new_n21379 = new_n21355 ^ new_n21335;
  assign new_n21380 = new_n21348 & new_n21379;
  assign new_n21381 = new_n21380 ^ new_n21335;
  assign new_n21382 = new_n21381 ^ new_n21342;
  assign new_n21383 = new_n21382 ^ new_n21378;
  assign new_n21384 = new_n21354 ^ new_n21337;
  assign new_n21385 = new_n21338 & new_n21384;
  assign new_n21386 = new_n21385 ^ new_n21344;
  assign new_n21387 = new_n21386 ^ new_n21367;
  assign new_n21388 = new_n21387 ^ new_n21383;
  assign new_n21389 = new_n21355 ^ new_n21330;
  assign new_n21390 = new_n21348 ^ new_n21326;
  assign new_n21391 = new_n21389 & new_n21390;
  assign new_n21392 = new_n21391 ^ new_n21370;
  assign new_n21393 = new_n21385 ^ new_n21363;
  assign new_n21394 = new_n21393 ^ new_n21392;
  assign new_n21395 = ~new_n21394 & new_n21388;
  assign new_n21396 = new_n21353 ^ new_n21330;
  assign new_n21397 = new_n21380 ^ new_n21358;
  assign new_n21398 = new_n21397 ^ new_n21393;
  assign new_n21399 = new_n21398 ^ new_n21396;
  assign new_n21400 = new_n21391 ^ new_n21369;
  assign new_n21401 = new_n21400 ^ new_n21330;
  assign new_n21402 = new_n21401 ^ new_n21387;
  assign new_n21403 = new_n21402 ^ new_n21378;
  assign new_n21404 = new_n21399 & new_n21403;
  assign new_n21405 = new_n21404 ^ new_n21395;
  assign new_n21406 = new_n21401 ^ new_n21382;
  assign new_n21407 = new_n21406 ^ new_n21405;
  assign new_n21408 = new_n21326 & new_n21407;
  assign new_n21409 = new_n21353 ^ new_n21314;
  assign new_n21410 = new_n21371 ^ new_n21358;
  assign new_n21411 = new_n21404 ^ new_n21382;
  assign new_n21412 = new_n21411 ^ new_n21387;
  assign new_n21413 = new_n21395 ^ new_n21378;
  assign new_n21414 = new_n21402 & new_n21413;
  assign new_n21415 = new_n21414 ^ new_n21403;
  assign new_n21416 = new_n21412 & new_n21415;
  assign new_n21417 = new_n21416 ^ new_n21414;
  assign new_n21418 = new_n21417 ^ new_n21410;
  assign new_n21419 = new_n21418 ^ new_n21409;
  assign new_n21420 = new_n21419 ^ new_n21335;
  assign new_n21421 = new_n21404 ^ new_n21369;
  assign new_n21422 = new_n21421 ^ new_n21342;
  assign new_n21423 = new_n21422 ^ new_n21420;
  assign new_n21424 = ~new_n21423 & new_n21361;
  assign new_n21425 = new_n21424 ^ new_n21408;
  assign new_n21426 = new_n21414 ^ new_n21395;
  assign new_n21427 = new_n21426 ^ new_n21394;
  assign new_n21428 = ~new_n21427 & new_n21349;
  assign new_n21429 = new_n21414 ^ new_n21377;
  assign new_n21430 = ~new_n21429 & new_n21337;
  assign new_n21431 = new_n21430 ^ new_n21428;
  assign new_n21432 = ~new_n21429 & new_n21340;
  assign new_n21433 = new_n21432 ^ new_n21431;
  assign new_n21434 = ~new_n21427 & new_n21357;
  assign new_n21435 = new_n21336 & new_n21407;
  assign new_n21436 = ~new_n21423 & new_n21362;
  assign new_n21437 = new_n21436 ^ new_n21435;
  assign new_n21438 = new_n21437 ^ new_n21434;
  assign new_n21439 = new_n21438 ^ new_n21433;
  assign new_n21440 = new_n21439 ^ new_n21425;
  assign new_n21441 = new_n18368 ^ new_n18298;
  assign new_n21442 = new_n15732 ^ new_n13049;
  assign new_n21443 = new_n21442 ^ new_n17838;
  assign new_n21444 = new_n21443 ^ new_n18321;
  assign new_n21445 = new_n21444 ^ new_n21441;
  assign new_n21446 = new_n18347 ^ new_n18138;
  assign new_n21447 = new_n21446 ^ new_n17838;
  assign new_n21448 = new_n16148 ^ new_n13019;
  assign new_n21449 = new_n21448 ^ new_n20474;
  assign new_n21450 = new_n21449 ^ new_n18444;
  assign new_n21451 = new_n21450 ^ new_n21447;
  assign new_n21452 = new_n20474 ^ new_n18458;
  assign new_n21453 = new_n21452 ^ new_n18288;
  assign new_n21454 = new_n16130 ^ new_n13027;
  assign new_n21455 = new_n21454 ^ new_n18321;
  assign new_n21456 = new_n21455 ^ new_n18455;
  assign new_n21457 = new_n21456 ^ new_n21453;
  assign new_n21458 = new_n21457 ^ new_n21451;
  assign new_n21459 = new_n21458 ^ new_n21445;
  assign new_n21460 = new_n18430 ^ new_n18418;
  assign new_n21461 = new_n16209 ^ new_n13056;
  assign new_n21462 = new_n21461 ^ new_n18379;
  assign new_n21463 = new_n21462 ^ new_n18425;
  assign new_n21464 = new_n21463 ^ new_n21460;
  assign new_n21465 = new_n21464 ^ new_n21459;
  assign new_n21466 = new_n18386 ^ new_n18338;
  assign new_n21467 = new_n16232 ^ new_n13034;
  assign new_n21468 = new_n21467 ^ new_n18407;
  assign new_n21469 = new_n21468 ^ new_n18379;
  assign new_n21470 = new_n21469 ^ new_n21466;
  assign new_n21471 = new_n16262 ^ new_n13038;
  assign new_n21472 = new_n21471 ^ new_n18434;
  assign new_n21473 = new_n21472 ^ new_n20474;
  assign new_n21474 = new_n18447 ^ new_n18355;
  assign new_n21475 = new_n21474 ^ new_n18347;
  assign new_n21476 = new_n21475 ^ new_n21473;
  assign new_n21477 = new_n21476 ^ new_n21470;
  assign new_n21478 = new_n21477 ^ new_n21458;
  assign new_n21479 = new_n21476 ^ new_n21445;
  assign new_n21480 = new_n21470 ^ new_n21457;
  assign new_n21481 = new_n21480 ^ new_n21479;
  assign new_n21482 = new_n21478 & new_n21481;
  assign new_n21483 = new_n21482 ^ new_n21464;
  assign new_n21484 = new_n21483 ^ new_n21478;
  assign new_n21485 = new_n21465 & new_n21477;
  assign new_n21486 = new_n18425 ^ new_n18401;
  assign new_n21487 = new_n16253 ^ new_n13062;
  assign new_n21488 = new_n21487 ^ new_n20453;
  assign new_n21489 = new_n21488 ^ new_n21486;
  assign new_n21490 = new_n21489 ^ new_n21464;
  assign new_n21491 = new_n16278 ^ new_n13076;
  assign new_n21492 = new_n21491 ^ new_n18455;
  assign new_n21493 = new_n20474 ^ new_n18311;
  assign new_n21494 = new_n21493 ^ new_n21492;
  assign new_n21495 = new_n21494 ^ new_n21490;
  assign new_n21496 = new_n21495 ^ new_n21457;
  assign new_n21497 = new_n21470 ^ new_n21445;
  assign new_n21498 = new_n21497 ^ new_n21496;
  assign new_n21499 = new_n21494 ^ new_n21478;
  assign new_n21500 = new_n21498 & new_n21499;
  assign new_n21501 = new_n21500 ^ new_n21485;
  assign new_n21502 = new_n21489 ^ new_n21476;
  assign new_n21503 = new_n21502 ^ new_n21497;
  assign new_n21504 = new_n21479 & new_n21503;
  assign new_n21505 = new_n21504 ^ new_n21445;
  assign new_n21506 = new_n21505 ^ new_n21501;
  assign new_n21507 = new_n21506 ^ new_n21484;
  assign new_n21508 = new_n21489 ^ new_n21459;
  assign new_n21509 = new_n21480 & new_n21508;
  assign new_n21510 = ~new_n21457 & ~new_n21495;
  assign new_n21511 = new_n21510 ^ new_n21457;
  assign new_n21512 = new_n21511 ^ new_n21509;
  assign new_n21513 = new_n21512 ^ new_n21497;
  assign new_n21514 = new_n21504 ^ new_n21485;
  assign new_n21515 = new_n21489 ^ new_n21451;
  assign new_n21516 = new_n21515 ^ new_n21514;
  assign new_n21517 = new_n21516 ^ new_n21513;
  assign new_n21518 = ~new_n21517 & new_n21507;
  assign new_n21519 = new_n21495 ^ new_n21476;
  assign new_n21520 = new_n21494 & new_n21519;
  assign new_n21521 = new_n21520 ^ new_n21476;
  assign new_n21522 = new_n21521 ^ new_n21483;
  assign new_n21523 = new_n21522 ^ new_n21518;
  assign new_n21524 = new_n21490 ^ new_n21478;
  assign new_n21525 = new_n21497 & new_n21524;
  assign new_n21526 = new_n21525 ^ new_n21485;
  assign new_n21527 = new_n21526 ^ new_n21508;
  assign new_n21528 = new_n21527 ^ new_n21523;
  assign new_n21529 = new_n21494 ^ new_n21465;
  assign new_n21530 = new_n21495 ^ new_n21470;
  assign new_n21531 = new_n21529 & new_n21530;
  assign new_n21532 = new_n21531 ^ new_n21510;
  assign new_n21533 = new_n21525 ^ new_n21504;
  assign new_n21534 = new_n21533 ^ new_n21532;
  assign new_n21535 = ~new_n21534 & new_n21528;
  assign new_n21536 = new_n21489 ^ new_n21470;
  assign new_n21537 = new_n21520 ^ new_n21500;
  assign new_n21538 = new_n21537 ^ new_n21533;
  assign new_n21539 = new_n21538 ^ new_n21536;
  assign new_n21540 = new_n21531 ^ new_n21509;
  assign new_n21541 = new_n21540 ^ new_n21470;
  assign new_n21542 = new_n21541 ^ new_n21527;
  assign new_n21543 = new_n21542 ^ new_n21518;
  assign new_n21544 = new_n21539 & new_n21543;
  assign new_n21545 = new_n21544 ^ new_n21535;
  assign new_n21546 = new_n21541 ^ new_n21522;
  assign new_n21547 = new_n21546 ^ new_n21545;
  assign new_n21548 = new_n21465 & new_n21547;
  assign new_n21549 = new_n21489 ^ new_n21457;
  assign new_n21550 = new_n21511 ^ new_n21500;
  assign new_n21551 = new_n21544 ^ new_n21522;
  assign new_n21552 = new_n21551 ^ new_n21527;
  assign new_n21553 = new_n21535 ^ new_n21518;
  assign new_n21554 = new_n21542 & new_n21553;
  assign new_n21555 = new_n21554 ^ new_n21543;
  assign new_n21556 = new_n21552 & new_n21555;
  assign new_n21557 = new_n21556 ^ new_n21554;
  assign new_n21558 = new_n21557 ^ new_n21550;
  assign new_n21559 = new_n21558 ^ new_n21549;
  assign new_n21560 = new_n21559 ^ new_n21476;
  assign new_n21561 = new_n21544 ^ new_n21509;
  assign new_n21562 = new_n21561 ^ new_n21483;
  assign new_n21563 = new_n21562 ^ new_n21560;
  assign new_n21564 = ~new_n21563 & new_n21503;
  assign new_n21565 = new_n21564 ^ new_n21548;
  assign new_n21566 = new_n21554 ^ new_n21535;
  assign new_n21567 = new_n21566 ^ new_n21534;
  assign new_n21568 = ~new_n21567 & new_n21499;
  assign new_n21569 = new_n21554 ^ new_n21517;
  assign new_n21570 = ~new_n21569 & new_n21478;
  assign new_n21571 = new_n21570 ^ new_n21568;
  assign new_n21572 = ~new_n21569 & new_n21481;
  assign new_n21573 = new_n21572 ^ new_n21571;
  assign new_n21574 = ~new_n21567 & new_n21498;
  assign new_n21575 = ~new_n21563 & new_n21479;
  assign new_n21576 = new_n21477 & new_n21547;
  assign new_n21577 = new_n21576 ^ new_n21575;
  assign new_n21578 = new_n21577 ^ new_n21574;
  assign new_n21579 = new_n21578 ^ new_n21573;
  assign new_n21580 = new_n21579 ^ new_n21565;
  assign new_n21581 = new_n21580 ^ new_n21440;
  assign new_n21582 = new_n21581 ^ new_n21305;
  assign new_n21583 = new_n15076 ^ new_n15067;
  assign new_n21584 = new_n16499 ^ new_n13669;
  assign new_n21585 = new_n21584 ^ new_n3529;
  assign new_n21586 = new_n21585 ^ new_n12756;
  assign new_n21587 = new_n21586 ^ new_n15099;
  assign new_n21588 = new_n21587 ^ new_n21583;
  assign new_n21589 = new_n17185 ^ new_n13684;
  assign new_n21590 = new_n21589 ^ new_n3594;
  assign new_n21591 = new_n21590 ^ new_n15193;
  assign new_n21592 = new_n21591 ^ new_n15160;
  assign new_n21593 = new_n15019 ^ new_n12756;
  assign new_n21594 = new_n21593 ^ new_n13828;
  assign new_n21595 = new_n21594 ^ new_n21592;
  assign new_n21596 = new_n15203 ^ new_n15004;
  assign new_n21597 = new_n21596 ^ new_n15160;
  assign new_n21598 = new_n17165 ^ new_n13640;
  assign new_n21599 = new_n21598 ^ new_n3421;
  assign new_n21600 = new_n21599 ^ new_n15210;
  assign new_n21601 = new_n21600 ^ new_n15076;
  assign new_n21602 = new_n21601 ^ new_n21597;
  assign new_n21603 = new_n21602 ^ new_n21595;
  assign new_n21604 = new_n21603 ^ new_n21588;
  assign new_n21605 = new_n15169 ^ new_n15154;
  assign new_n21606 = new_n17241 ^ new_n13572;
  assign new_n21607 = new_n21606 ^ new_n3621;
  assign new_n21608 = new_n21607 ^ new_n15180;
  assign new_n21609 = new_n21608 ^ new_n15110;
  assign new_n21610 = new_n21609 ^ new_n21605;
  assign new_n21611 = new_n21610 ^ new_n21604;
  assign new_n21612 = new_n15110 ^ new_n15054;
  assign new_n21613 = new_n17290 ^ new_n13713;
  assign new_n21614 = new_n21613 ^ new_n3474;
  assign new_n21615 = new_n21614 ^ new_n15159;
  assign new_n21616 = new_n21615 ^ new_n15134;
  assign new_n21617 = new_n21616 ^ new_n21612;
  assign new_n21618 = new_n15169 ^ new_n15119;
  assign new_n21619 = new_n17269 ^ new_n13550;
  assign new_n21620 = new_n21619 ^ new_n3646;
  assign new_n21621 = new_n15197 ^ new_n15195;
  assign new_n21622 = new_n21621 ^ new_n21620;
  assign new_n21623 = new_n21622 ^ new_n21618;
  assign new_n21624 = new_n21623 ^ new_n21610;
  assign new_n21625 = new_n17298 ^ new_n13601;
  assign new_n21626 = new_n21625 ^ new_n3661;
  assign new_n21627 = new_n21626 ^ new_n15203;
  assign new_n21628 = new_n15160 ^ new_n15082;
  assign new_n21629 = new_n21628 ^ new_n21627;
  assign new_n21630 = new_n21629 ^ new_n21624;
  assign new_n21631 = new_n21630 ^ new_n21617;
  assign new_n21632 = new_n21629 ^ new_n21611;
  assign new_n21633 = ~new_n21631 & new_n21632;
  assign new_n21634 = new_n21623 ^ new_n21604;
  assign new_n21635 = new_n21617 ^ new_n21602;
  assign new_n21636 = ~new_n21634 & new_n21635;
  assign new_n21637 = new_n21636 ^ new_n21633;
  assign new_n21638 = new_n21637 ^ new_n21617;
  assign new_n21639 = new_n21617 ^ new_n21588;
  assign new_n21640 = new_n17315 ^ new_n12868;
  assign new_n21641 = new_n21640 ^ new_n3553;
  assign new_n21642 = new_n21641 ^ new_n15165;
  assign new_n21643 = new_n21642 ^ new_n15160;
  assign new_n21644 = new_n15197 ^ new_n15019;
  assign new_n21645 = new_n21644 ^ new_n15027;
  assign new_n21646 = new_n21645 ^ new_n21643;
  assign new_n21647 = new_n21646 ^ new_n21617;
  assign new_n21648 = new_n21647 ^ new_n21603;
  assign new_n21649 = new_n21648 ^ new_n21624;
  assign new_n21650 = new_n21639 & new_n21649;
  assign new_n21651 = ~new_n21611 & ~new_n21647;
  assign new_n21652 = new_n21651 ^ new_n21650;
  assign new_n21653 = new_n21652 ^ new_n21634;
  assign new_n21654 = new_n21653 ^ new_n21638;
  assign new_n21655 = new_n21646 ^ new_n21602;
  assign new_n21656 = new_n21655 ^ new_n21639;
  assign new_n21657 = ~new_n21656 & new_n21648;
  assign new_n21658 = new_n21657 ^ new_n21610;
  assign new_n21659 = new_n21658 ^ new_n21648;
  assign new_n21660 = new_n21648 ^ new_n21629;
  assign new_n21661 = new_n21630 ^ new_n21602;
  assign new_n21662 = new_n21661 ^ new_n21639;
  assign new_n21663 = ~new_n21660 & ~new_n21662;
  assign new_n21664 = new_n21663 ^ new_n21651;
  assign new_n21665 = new_n21646 ^ new_n21588;
  assign new_n21666 = new_n21646 ^ new_n21623;
  assign new_n21667 = new_n21666 ^ new_n21639;
  assign new_n21668 = ~new_n21665 & ~new_n21667;
  assign new_n21669 = new_n21668 ^ new_n21588;
  assign new_n21670 = new_n21669 ^ new_n21664;
  assign new_n21671 = new_n21670 ^ new_n21659;
  assign new_n21672 = ~new_n21602 & new_n21630;
  assign new_n21673 = new_n21672 ^ new_n21602;
  assign new_n21674 = new_n21673 ^ new_n21636;
  assign new_n21675 = new_n21674 ^ new_n21639;
  assign new_n21676 = new_n21668 ^ new_n21651;
  assign new_n21677 = new_n21623 ^ new_n21595;
  assign new_n21678 = new_n21677 ^ new_n21676;
  assign new_n21679 = new_n21678 ^ new_n21675;
  assign new_n21680 = new_n21671 & new_n21679;
  assign new_n21681 = new_n21680 ^ new_n21654;
  assign new_n21682 = new_n21623 ^ new_n21617;
  assign new_n21683 = new_n21646 ^ new_n21630;
  assign new_n21684 = ~new_n21629 & new_n21683;
  assign new_n21685 = new_n21684 ^ new_n21663;
  assign new_n21686 = new_n21668 ^ new_n21650;
  assign new_n21687 = new_n21686 ^ new_n21685;
  assign new_n21688 = new_n21687 ^ new_n21682;
  assign new_n21689 = ~new_n21681 & new_n21688;
  assign new_n21690 = new_n21684 ^ new_n21646;
  assign new_n21691 = new_n21690 ^ new_n21658;
  assign new_n21692 = new_n21691 ^ new_n21680;
  assign new_n21693 = new_n21692 ^ new_n21653;
  assign new_n21694 = new_n21672 ^ new_n21633;
  assign new_n21695 = new_n21694 ^ new_n21686;
  assign new_n21696 = ~new_n21695 & new_n21693;
  assign new_n21697 = new_n21696 ^ new_n21689;
  assign new_n21698 = new_n21691 ^ new_n21638;
  assign new_n21699 = new_n21698 ^ new_n21697;
  assign new_n21700 = ~new_n21611 & ~new_n21699;
  assign new_n21701 = new_n21696 ^ new_n21680;
  assign new_n21702 = ~new_n21701 & new_n21654;
  assign new_n21703 = new_n21702 ^ new_n21696;
  assign new_n21704 = new_n21703 ^ new_n21681;
  assign new_n21705 = new_n21704 ^ new_n21679;
  assign new_n21706 = ~new_n21656 & new_n21705;
  assign new_n21707 = new_n21706 ^ new_n21700;
  assign new_n21708 = new_n21691 ^ new_n21689;
  assign new_n21709 = new_n21708 ^ new_n21653;
  assign new_n21710 = ~new_n21703 & new_n21709;
  assign new_n21711 = new_n21710 ^ new_n21688;
  assign new_n21712 = ~new_n21630 & new_n21711;
  assign new_n21713 = new_n21704 ^ new_n21696;
  assign new_n21714 = new_n21713 ^ new_n21695;
  assign new_n21715 = ~new_n21662 & ~new_n21714;
  assign new_n21716 = ~new_n21647 & ~new_n21699;
  assign new_n21717 = new_n21623 ^ new_n21602;
  assign new_n21718 = new_n21673 ^ new_n21663;
  assign new_n21719 = new_n21710 ^ new_n21704;
  assign new_n21720 = new_n21719 ^ new_n21718;
  assign new_n21721 = new_n21720 ^ new_n21717;
  assign new_n21722 = new_n21721 ^ new_n21646;
  assign new_n21723 = new_n21689 ^ new_n21636;
  assign new_n21724 = new_n21723 ^ new_n21658;
  assign new_n21725 = new_n21724 ^ new_n21722;
  assign new_n21726 = ~new_n21665 & new_n21725;
  assign new_n21727 = new_n21726 ^ new_n21716;
  assign new_n21728 = new_n21727 ^ new_n21715;
  assign new_n21729 = new_n21728 ^ new_n21712;
  assign new_n21730 = new_n21710 ^ new_n21689;
  assign new_n21731 = new_n21730 ^ new_n21671;
  assign new_n21732 = ~new_n21634 & new_n21731;
  assign new_n21733 = new_n21732 ^ new_n21729;
  assign new_n21734 = ~new_n21667 & new_n21725;
  assign new_n21735 = new_n21734 ^ new_n21733;
  assign new_n21736 = new_n21735 ^ new_n21707;
  assign new_n21737 = new_n21572 ^ new_n21548;
  assign new_n21738 = new_n21556 ^ new_n21539;
  assign new_n21739 = new_n21495 & new_n21738;
  assign new_n21740 = new_n21739 ^ new_n21578;
  assign new_n21741 = new_n21556 ^ new_n21544;
  assign new_n21742 = new_n21741 ^ new_n21507;
  assign new_n21743 = new_n21508 & new_n21742;
  assign new_n21744 = new_n21743 ^ new_n21740;
  assign new_n21745 = new_n21744 ^ new_n21564;
  assign new_n21746 = new_n21745 ^ new_n21737;
  assign new_n21747 = new_n21746 ^ new_n21736;
  assign new_n21748 = new_n16157 ^ new_n16140;
  assign new_n21749 = new_n17556 ^ new_n15921;
  assign new_n21750 = new_n21749 ^ new_n16122;
  assign new_n21751 = new_n21750 ^ new_n21748;
  assign new_n21752 = new_n16175 ^ new_n15921;
  assign new_n21753 = new_n21752 ^ new_n16082;
  assign new_n21754 = new_n17525 ^ new_n16229;
  assign new_n21755 = new_n21754 ^ new_n16269;
  assign new_n21756 = new_n21755 ^ new_n21753;
  assign new_n21757 = new_n16282 ^ new_n16229;
  assign new_n21758 = new_n21757 ^ new_n15616;
  assign new_n21759 = new_n17542 ^ new_n16122;
  assign new_n21760 = new_n21759 ^ new_n16276;
  assign new_n21761 = new_n21760 ^ new_n21758;
  assign new_n21762 = new_n21761 ^ new_n21756;
  assign new_n21763 = new_n21762 ^ new_n21751;
  assign new_n21764 = new_n17564 ^ new_n16203;
  assign new_n21765 = new_n19367 ^ new_n16245;
  assign new_n21766 = new_n21765 ^ new_n21764;
  assign new_n21767 = new_n21766 ^ new_n21763;
  assign new_n21768 = new_n17568 ^ new_n16088;
  assign new_n21769 = new_n19329 ^ new_n16193;
  assign new_n21770 = new_n21769 ^ new_n21768;
  assign new_n21771 = new_n17573 ^ new_n16215;
  assign new_n21772 = new_n19343 ^ new_n16260;
  assign new_n21773 = new_n21772 ^ new_n21771;
  assign new_n21774 = new_n21773 ^ new_n21766;
  assign new_n21775 = new_n17581 ^ new_n16276;
  assign new_n21776 = new_n16229 ^ new_n16113;
  assign new_n21777 = new_n21776 ^ new_n21775;
  assign new_n21778 = new_n21777 ^ new_n21774;
  assign new_n21779 = new_n21778 ^ new_n21770;
  assign new_n21780 = new_n21777 ^ new_n21767;
  assign new_n21781 = ~new_n21779 & ~new_n21780;
  assign new_n21782 = new_n21770 ^ new_n21761;
  assign new_n21783 = new_n21773 ^ new_n21763;
  assign new_n21784 = ~new_n21782 & new_n21783;
  assign new_n21785 = new_n21784 ^ new_n21781;
  assign new_n21786 = new_n21785 ^ new_n21770;
  assign new_n21787 = new_n21770 ^ new_n21751;
  assign new_n21788 = new_n17576 ^ new_n16229;
  assign new_n21789 = new_n21788 ^ new_n19357;
  assign new_n21790 = new_n16248 ^ new_n16176;
  assign new_n21791 = new_n21790 ^ new_n21789;
  assign new_n21792 = new_n21791 ^ new_n21770;
  assign new_n21793 = new_n21792 ^ new_n21762;
  assign new_n21794 = new_n21793 ^ new_n21774;
  assign new_n21795 = ~new_n21794 & new_n21787;
  assign new_n21796 = new_n21767 & new_n21792;
  assign new_n21797 = new_n21796 ^ new_n21795;
  assign new_n21798 = new_n21797 ^ new_n21783;
  assign new_n21799 = new_n21798 ^ new_n21786;
  assign new_n21800 = new_n21791 ^ new_n21751;
  assign new_n21801 = new_n21800 ^ new_n21782;
  assign new_n21802 = ~new_n21793 & ~new_n21801;
  assign new_n21803 = new_n21802 ^ new_n21766;
  assign new_n21804 = new_n21803 ^ new_n21793;
  assign new_n21805 = new_n21793 ^ new_n21777;
  assign new_n21806 = new_n21778 ^ new_n21761;
  assign new_n21807 = new_n21806 ^ new_n21787;
  assign new_n21808 = new_n21805 & new_n21807;
  assign new_n21809 = new_n21808 ^ new_n21796;
  assign new_n21810 = new_n21791 ^ new_n21773;
  assign new_n21811 = new_n21810 ^ new_n21787;
  assign new_n21812 = ~new_n21811 & new_n21800;
  assign new_n21813 = new_n21812 ^ new_n21751;
  assign new_n21814 = new_n21813 ^ new_n21809;
  assign new_n21815 = new_n21814 ^ new_n21804;
  assign new_n21816 = new_n21761 & new_n21778;
  assign new_n21817 = new_n21816 ^ new_n21761;
  assign new_n21818 = new_n21817 ^ new_n21784;
  assign new_n21819 = new_n21818 ^ new_n21787;
  assign new_n21820 = new_n21812 ^ new_n21796;
  assign new_n21821 = new_n21773 ^ new_n21756;
  assign new_n21822 = new_n21821 ^ new_n21820;
  assign new_n21823 = new_n21822 ^ new_n21819;
  assign new_n21824 = ~new_n21823 & new_n21815;
  assign new_n21825 = new_n21824 ^ new_n21799;
  assign new_n21826 = new_n21773 ^ new_n21770;
  assign new_n21827 = new_n21791 ^ new_n21778;
  assign new_n21828 = ~new_n21777 & ~new_n21827;
  assign new_n21829 = new_n21828 ^ new_n21808;
  assign new_n21830 = new_n21812 ^ new_n21795;
  assign new_n21831 = new_n21830 ^ new_n21829;
  assign new_n21832 = new_n21831 ^ new_n21826;
  assign new_n21833 = ~new_n21832 & new_n21825;
  assign new_n21834 = new_n21828 ^ new_n21791;
  assign new_n21835 = new_n21834 ^ new_n21803;
  assign new_n21836 = new_n21835 ^ new_n21824;
  assign new_n21837 = new_n21836 ^ new_n21798;
  assign new_n21838 = new_n21816 ^ new_n21781;
  assign new_n21839 = new_n21838 ^ new_n21830;
  assign new_n21840 = ~new_n21837 & ~new_n21839;
  assign new_n21841 = new_n21840 ^ new_n21833;
  assign new_n21842 = new_n21835 ^ new_n21786;
  assign new_n21843 = new_n21842 ^ new_n21841;
  assign new_n21844 = ~new_n21843 & new_n21767;
  assign new_n21845 = new_n21840 ^ new_n21824;
  assign new_n21846 = ~new_n21799 & ~new_n21845;
  assign new_n21847 = new_n21846 ^ new_n21840;
  assign new_n21848 = new_n21847 ^ new_n21825;
  assign new_n21849 = new_n21848 ^ new_n21823;
  assign new_n21850 = ~new_n21801 & new_n21849;
  assign new_n21851 = new_n21850 ^ new_n21844;
  assign new_n21852 = new_n21835 ^ new_n21833;
  assign new_n21853 = new_n21852 ^ new_n21798;
  assign new_n21854 = ~new_n21847 & ~new_n21853;
  assign new_n21855 = new_n21854 ^ new_n21832;
  assign new_n21856 = ~new_n21778 & ~new_n21855;
  assign new_n21857 = new_n21848 ^ new_n21840;
  assign new_n21858 = new_n21857 ^ new_n21839;
  assign new_n21859 = new_n21807 & new_n21858;
  assign new_n21860 = ~new_n21843 & new_n21792;
  assign new_n21861 = new_n21773 ^ new_n21761;
  assign new_n21862 = new_n21817 ^ new_n21808;
  assign new_n21863 = new_n21854 ^ new_n21848;
  assign new_n21864 = new_n21863 ^ new_n21862;
  assign new_n21865 = new_n21864 ^ new_n21861;
  assign new_n21866 = new_n21865 ^ new_n21791;
  assign new_n21867 = new_n21833 ^ new_n21784;
  assign new_n21868 = new_n21867 ^ new_n21803;
  assign new_n21869 = new_n21868 ^ new_n21866;
  assign new_n21870 = new_n21800 & new_n21869;
  assign new_n21871 = new_n21870 ^ new_n21860;
  assign new_n21872 = new_n21871 ^ new_n21859;
  assign new_n21873 = new_n21872 ^ new_n21856;
  assign new_n21874 = new_n21854 ^ new_n21833;
  assign new_n21875 = new_n21874 ^ new_n21815;
  assign new_n21876 = new_n21783 & new_n21875;
  assign new_n21877 = new_n21876 ^ new_n21873;
  assign new_n21878 = ~new_n21811 & new_n21869;
  assign new_n21879 = new_n21878 ^ new_n21877;
  assign new_n21880 = new_n21879 ^ new_n21851;
  assign new_n21881 = new_n21880 ^ new_n21747;
  assign new_n21882 = new_n21881 ^ new_n21582;
  assign new_n21883 = new_n21840 ^ new_n21770;
  assign new_n21884 = new_n21828 ^ new_n21781;
  assign new_n21885 = new_n21884 ^ new_n21865;
  assign new_n21886 = new_n21885 ^ new_n21883;
  assign new_n21887 = ~new_n21794 & ~new_n21886;
  assign new_n21888 = ~new_n21782 & new_n21875;
  assign new_n21889 = new_n21888 ^ new_n21887;
  assign new_n21890 = new_n21878 ^ new_n21856;
  assign new_n21891 = ~new_n21855 & new_n21806;
  assign new_n21892 = ~new_n21780 & ~new_n21853;
  assign new_n21893 = new_n21892 ^ new_n21891;
  assign new_n21894 = new_n21893 ^ new_n21871;
  assign new_n21895 = new_n21894 ^ new_n21890;
  assign new_n21896 = new_n21895 ^ new_n21889;
  assign new_n21897 = new_n21432 ^ new_n21408;
  assign new_n21898 = new_n21416 ^ new_n21404;
  assign new_n21899 = new_n21898 ^ new_n21366;
  assign new_n21900 = new_n21367 & new_n21899;
  assign new_n21901 = new_n21416 ^ new_n21399;
  assign new_n21902 = new_n21355 & new_n21901;
  assign new_n21903 = new_n21902 ^ new_n21438;
  assign new_n21904 = new_n21903 ^ new_n21900;
  assign new_n21905 = new_n21904 ^ new_n21424;
  assign new_n21906 = new_n21905 ^ new_n21897;
  assign new_n21907 = new_n21906 ^ new_n21746;
  assign new_n21908 = new_n21907 ^ new_n21896;
  assign new_n21909 = new_n21356 & new_n21901;
  assign new_n21910 = new_n21390 & new_n21412;
  assign new_n21911 = new_n21910 ^ new_n21909;
  assign new_n21912 = new_n21911 ^ new_n21437;
  assign new_n21913 = new_n21368 & new_n21899;
  assign new_n21914 = new_n21402 ^ new_n21395;
  assign new_n21915 = new_n21348 & new_n21914;
  assign new_n21916 = new_n21915 ^ new_n21430;
  assign new_n21917 = new_n21916 ^ new_n21913;
  assign new_n21918 = new_n21917 ^ new_n21900;
  assign new_n21919 = new_n21918 ^ new_n21912;
  assign new_n21920 = new_n21480 & new_n21742;
  assign new_n21921 = new_n21542 ^ new_n21535;
  assign new_n21922 = new_n21494 & new_n21921;
  assign new_n21923 = new_n21922 ^ new_n21570;
  assign new_n21924 = new_n21923 ^ new_n21920;
  assign new_n21925 = new_n21924 ^ new_n21743;
  assign new_n21926 = new_n21496 & new_n21738;
  assign new_n21927 = new_n21529 & new_n21552;
  assign new_n21928 = new_n21927 ^ new_n21926;
  assign new_n21929 = new_n21928 ^ new_n21577;
  assign new_n21930 = new_n21929 ^ new_n21925;
  assign new_n21931 = new_n21930 ^ new_n21919;
  assign new_n21932 = new_n21931 ^ new_n21908;
  assign new_n21933 = new_n21535 ^ new_n21470;
  assign new_n21934 = new_n21531 ^ new_n21520;
  assign new_n21935 = new_n21934 ^ new_n21559;
  assign new_n21936 = new_n21935 ^ new_n21933;
  assign new_n21937 = ~new_n21936 & new_n21524;
  assign new_n21938 = new_n21937 ^ new_n21920;
  assign new_n21939 = new_n21739 ^ new_n21564;
  assign new_n21940 = new_n21939 ^ new_n21929;
  assign new_n21941 = new_n21940 ^ new_n21938;
  assign new_n21942 = new_n21263 ^ new_n16233;
  assign new_n21943 = new_n21228 ^ new_n21215;
  assign new_n21944 = new_n21943 ^ new_n21288;
  assign new_n21945 = new_n21944 ^ new_n21942;
  assign new_n21946 = ~new_n21945 & new_n21217;
  assign new_n21947 = new_n21230 & new_n21298;
  assign new_n21948 = new_n21947 ^ new_n21946;
  assign new_n21949 = new_n21301 ^ new_n21279;
  assign new_n21950 = new_n21210 & new_n21278;
  assign new_n21951 = new_n21227 & new_n21275;
  assign new_n21952 = new_n21951 ^ new_n21950;
  assign new_n21953 = new_n21952 ^ new_n21294;
  assign new_n21954 = new_n21953 ^ new_n21949;
  assign new_n21955 = new_n21954 ^ new_n21948;
  assign new_n21956 = new_n21955 ^ new_n15090;
  assign new_n21957 = new_n21956 ^ new_n10840;
  assign new_n21958 = new_n21696 ^ new_n21617;
  assign new_n21959 = new_n21684 ^ new_n21633;
  assign new_n21960 = new_n21959 ^ new_n21721;
  assign new_n21961 = new_n21960 ^ new_n21958;
  assign new_n21962 = ~new_n21961 & new_n21649;
  assign new_n21963 = new_n21635 & new_n21731;
  assign new_n21964 = new_n21963 ^ new_n21962;
  assign new_n21965 = new_n21734 ^ new_n21712;
  assign new_n21966 = ~new_n21661 & new_n21711;
  assign new_n21967 = new_n21632 & new_n21709;
  assign new_n21968 = new_n21967 ^ new_n21966;
  assign new_n21969 = new_n21968 ^ new_n21727;
  assign new_n21970 = new_n21969 ^ new_n21965;
  assign new_n21971 = new_n21970 ^ new_n21964;
  assign new_n21972 = new_n21971 ^ new_n21957;
  assign new_n21973 = new_n21972 ^ new_n21941;
  assign new_n21974 = new_n21973 ^ new_n21932;
  assign new_n21975 = new_n21974 ^ new_n21882;
  assign new_n21976 = new_n21840 ^ new_n21799;
  assign new_n21977 = ~new_n21827 & new_n21976;
  assign new_n21978 = new_n21977 ^ new_n21879;
  assign new_n21979 = ~new_n21779 & ~new_n21853;
  assign new_n21980 = new_n21979 ^ new_n21887;
  assign new_n21981 = ~new_n21793 & new_n21849;
  assign new_n21982 = ~new_n21777 & new_n21976;
  assign new_n21983 = new_n21982 ^ new_n21981;
  assign new_n21984 = new_n21983 ^ new_n21888;
  assign new_n21985 = new_n21984 ^ new_n21980;
  assign new_n21986 = new_n21985 ^ new_n21978;
  assign new_n21987 = new_n21530 & new_n21552;
  assign new_n21988 = new_n21987 ^ new_n21937;
  assign new_n21989 = new_n21988 ^ new_n21924;
  assign new_n21990 = new_n21519 & new_n21921;
  assign new_n21991 = new_n21990 ^ new_n21745;
  assign new_n21992 = new_n21991 ^ new_n21989;
  assign new_n21993 = new_n21992 ^ new_n21986;
  assign new_n21994 = new_n21696 ^ new_n21654;
  assign new_n21995 = ~new_n21994 & new_n21683;
  assign new_n21996 = new_n21995 ^ new_n21735;
  assign new_n21997 = ~new_n21631 & new_n21709;
  assign new_n21998 = new_n21997 ^ new_n21962;
  assign new_n21999 = new_n21648 & new_n21705;
  assign new_n22000 = ~new_n21629 & ~new_n21994;
  assign new_n22001 = new_n22000 ^ new_n21999;
  assign new_n22002 = new_n22001 ^ new_n21963;
  assign new_n22003 = new_n22002 ^ new_n21998;
  assign new_n22004 = new_n22003 ^ new_n21996;
  assign new_n22005 = new_n22004 ^ new_n21993;
  assign new_n22006 = new_n21263 ^ new_n21237;
  assign new_n22007 = new_n21214 & new_n22006;
  assign new_n22008 = new_n22007 ^ new_n21302;
  assign new_n22009 = new_n21226 & new_n21275;
  assign new_n22010 = new_n22009 ^ new_n21946;
  assign new_n22011 = ~new_n21271 & new_n21206;
  assign new_n22012 = new_n16279 & new_n22006;
  assign new_n22013 = new_n22012 ^ new_n22011;
  assign new_n22014 = new_n22013 ^ new_n21947;
  assign new_n22015 = new_n22014 ^ new_n22010;
  assign new_n22016 = new_n22015 ^ new_n22008;
  assign new_n22017 = new_n22016 ^ new_n13955;
  assign new_n22018 = new_n22017 ^ new_n10829;
  assign new_n22019 = new_n21395 ^ new_n21330;
  assign new_n22020 = new_n21391 ^ new_n21380;
  assign new_n22021 = new_n22020 ^ new_n21419;
  assign new_n22022 = new_n22021 ^ new_n22019;
  assign new_n22023 = ~new_n22022 & new_n21384;
  assign new_n22024 = new_n22023 ^ new_n21913;
  assign new_n22025 = new_n21902 ^ new_n21424;
  assign new_n22026 = new_n22025 ^ new_n21912;
  assign new_n22027 = new_n22026 ^ new_n22024;
  assign new_n22028 = new_n22027 ^ new_n21941;
  assign new_n22029 = new_n22028 ^ new_n22018;
  assign new_n22030 = new_n22029 ^ new_n22005;
  assign new_n22031 = new_n22030 ^ new_n21882;
  assign new_n22032 = new_n21878 ^ new_n21844;
  assign new_n22033 = new_n21805 & new_n21858;
  assign new_n22034 = new_n22033 ^ new_n21981;
  assign new_n22035 = new_n22034 ^ new_n21850;
  assign new_n22036 = new_n22035 ^ new_n21872;
  assign new_n22037 = new_n22036 ^ new_n22032;
  assign new_n22038 = new_n21435 ^ new_n21408;
  assign new_n22039 = ~new_n22022 & new_n21338;
  assign new_n22040 = new_n21389 & new_n21412;
  assign new_n22041 = new_n22040 ^ new_n22023;
  assign new_n22042 = new_n22041 ^ new_n21917;
  assign new_n22043 = new_n22042 ^ new_n22039;
  assign new_n22044 = new_n22043 ^ new_n22038;
  assign new_n22045 = new_n21576 ^ new_n21548;
  assign new_n22046 = ~new_n21936 & new_n21497;
  assign new_n22047 = new_n22046 ^ new_n21989;
  assign new_n22048 = new_n22047 ^ new_n22045;
  assign new_n22049 = new_n22048 ^ new_n22044;
  assign new_n22050 = new_n22049 ^ new_n22037;
  assign new_n22051 = new_n21301 ^ new_n21267;
  assign new_n22052 = ~new_n21281 & new_n21207;
  assign new_n22053 = new_n22052 ^ new_n22011;
  assign new_n22054 = new_n22053 ^ new_n21272;
  assign new_n22055 = new_n22054 ^ new_n21295;
  assign new_n22056 = new_n22055 ^ new_n22051;
  assign new_n22057 = new_n22056 ^ new_n15126;
  assign new_n22058 = new_n22057 ^ new_n10846;
  assign new_n22059 = new_n21734 ^ new_n21700;
  assign new_n22060 = ~new_n21660 & ~new_n21714;
  assign new_n22061 = new_n22060 ^ new_n21999;
  assign new_n22062 = new_n22061 ^ new_n21706;
  assign new_n22063 = new_n22062 ^ new_n21728;
  assign new_n22064 = new_n22063 ^ new_n22059;
  assign new_n22065 = new_n22064 ^ new_n22058;
  assign new_n22066 = new_n22065 ^ new_n21580;
  assign new_n22067 = new_n22066 ^ new_n22050;
  assign new_n22068 = new_n21860 ^ new_n21844;
  assign new_n22069 = ~new_n21886 & new_n21787;
  assign new_n22070 = new_n22069 ^ new_n21985;
  assign new_n22071 = new_n22070 ^ new_n22068;
  assign new_n22072 = new_n21904 ^ new_n21433;
  assign new_n22073 = new_n21744 ^ new_n21573;
  assign new_n22074 = new_n22073 ^ new_n22072;
  assign new_n22075 = new_n22074 ^ new_n22071;
  assign new_n22076 = new_n21283 ^ new_n21267;
  assign new_n22077 = ~new_n21945 & new_n21211;
  assign new_n22078 = new_n22077 ^ new_n22015;
  assign new_n22079 = new_n22078 ^ new_n22076;
  assign new_n22080 = new_n22079 ^ new_n15174;
  assign new_n22081 = new_n22080 ^ new_n10817;
  assign new_n22082 = new_n21716 ^ new_n21700;
  assign new_n22083 = ~new_n21961 & new_n21639;
  assign new_n22084 = new_n22083 ^ new_n22003;
  assign new_n22085 = new_n22084 ^ new_n22082;
  assign new_n22086 = new_n22085 ^ new_n22081;
  assign new_n22087 = new_n22086 ^ new_n22048;
  assign new_n22088 = new_n22087 ^ new_n22075;
  assign new_n22089 = new_n22088 ^ new_n22067;
  assign new_n22090 = new_n22054 ^ new_n21300;
  assign new_n22091 = new_n22090 ^ new_n15185;
  assign new_n22092 = new_n22091 ^ new_n10821;
  assign new_n22093 = new_n22092 ^ new_n21907;
  assign new_n22094 = new_n21910 ^ new_n21432;
  assign new_n22095 = new_n21915 ^ new_n21428;
  assign new_n22096 = new_n22095 ^ new_n21903;
  assign new_n22097 = new_n22096 ^ new_n22094;
  assign new_n22098 = new_n21927 ^ new_n21572;
  assign new_n22099 = new_n21922 ^ new_n21568;
  assign new_n22100 = new_n22099 ^ new_n21740;
  assign new_n22101 = new_n22100 ^ new_n22098;
  assign new_n22102 = new_n22101 ^ new_n22097;
  assign new_n22103 = new_n22102 ^ new_n22093;
  assign new_n22104 = new_n22062 ^ new_n21733;
  assign new_n22105 = new_n22104 ^ new_n22073;
  assign new_n22106 = new_n22035 ^ new_n21877;
  assign new_n22107 = new_n22106 ^ new_n22105;
  assign new_n22108 = new_n22107 ^ new_n22103;
  assign new_n22109 = new_n22108 ^ new_n21882;
  assign new_n22110 = new_n21892 ^ new_n21850;
  assign new_n22111 = new_n22033 ^ new_n21982;
  assign new_n22112 = new_n22111 ^ new_n21873;
  assign new_n22113 = new_n22112 ^ new_n22110;
  assign new_n22114 = new_n22113 ^ new_n22101;
  assign new_n22115 = new_n21967 ^ new_n21706;
  assign new_n22116 = new_n22060 ^ new_n22000;
  assign new_n22117 = new_n22116 ^ new_n21729;
  assign new_n22118 = new_n22117 ^ new_n22115;
  assign new_n22119 = new_n22118 ^ new_n22114;
  assign new_n22120 = new_n21951 ^ new_n21272;
  assign new_n22121 = new_n22052 ^ new_n22012;
  assign new_n22122 = new_n22121 ^ new_n21296;
  assign new_n22123 = new_n22122 ^ new_n22120;
  assign new_n22124 = new_n22123 ^ new_n15035;
  assign new_n22125 = new_n22124 ^ new_n10861;
  assign new_n22126 = new_n22125 ^ new_n21907;
  assign new_n22127 = new_n21379 & new_n21914;
  assign new_n22128 = new_n22127 ^ new_n21905;
  assign new_n22129 = new_n22128 ^ new_n22042;
  assign new_n22130 = new_n22129 ^ new_n21992;
  assign new_n22131 = new_n22130 ^ new_n22126;
  assign new_n22132 = new_n22131 ^ new_n22119;
  assign new_n22133 = new_n22132 ^ new_n21974;
  assign new_n22134 = new_n22133 ^ new_n22109;
  assign new_n22135 = new_n22134 ^ new_n22089;
  assign new_n22136 = ~new_n22135 & new_n22031;
  assign new_n22137 = new_n22133 ^ new_n22030;
  assign new_n22138 = new_n22137 ^ new_n22067;
  assign new_n22139 = new_n22109 & new_n22138;
  assign new_n22140 = new_n22139 ^ new_n22136;
  assign new_n22141 = new_n22137 ^ new_n22088;
  assign new_n22142 = new_n22141 ^ new_n22140;
  assign new_n22143 = new_n21984 ^ new_n21876;
  assign new_n22144 = new_n22143 ^ new_n21894;
  assign new_n22145 = new_n22144 ^ new_n21907;
  assign new_n22146 = new_n22014 ^ new_n21299;
  assign new_n22147 = new_n22146 ^ new_n21953;
  assign new_n22148 = new_n22147 ^ new_n15206;
  assign new_n22149 = new_n22148 ^ new_n10852;
  assign new_n22150 = new_n22002 ^ new_n21732;
  assign new_n22151 = new_n22150 ^ new_n21969;
  assign new_n22152 = new_n22151 ^ new_n22149;
  assign new_n22153 = new_n22152 ^ new_n21930;
  assign new_n22154 = new_n22153 ^ new_n22145;
  assign new_n22155 = new_n22154 ^ new_n22089;
  assign new_n22156 = new_n22155 ^ new_n21882;
  assign new_n22157 = new_n22154 ^ new_n22138;
  assign new_n22158 = ~new_n22156 & ~new_n22157;
  assign new_n22159 = ~new_n21975 & new_n22141;
  assign new_n22160 = new_n22159 ^ new_n22158;
  assign new_n22161 = new_n22160 ^ new_n21882;
  assign new_n22162 = new_n22161 ^ new_n22142;
  assign new_n22163 = new_n22155 ^ new_n22108;
  assign new_n22164 = ~new_n22154 & ~new_n22163;
  assign new_n22165 = new_n22164 ^ new_n22108;
  assign new_n22166 = new_n22108 ^ new_n22030;
  assign new_n22167 = new_n22166 ^ new_n21975;
  assign new_n22168 = ~new_n22134 & ~new_n22167;
  assign new_n22169 = new_n22168 ^ new_n22067;
  assign new_n22170 = new_n22169 ^ new_n22165;
  assign new_n22171 = new_n21974 & new_n22155;
  assign new_n22172 = new_n22171 ^ new_n21974;
  assign new_n22173 = new_n22172 ^ new_n22159;
  assign new_n22174 = new_n22173 ^ new_n22031;
  assign new_n22175 = new_n22108 ^ new_n22088;
  assign new_n22176 = new_n22175 ^ new_n22031;
  assign new_n22177 = ~new_n22176 & new_n22166;
  assign new_n22178 = new_n22177 ^ new_n22139;
  assign new_n22179 = new_n22132 ^ new_n22088;
  assign new_n22180 = new_n22179 ^ new_n22178;
  assign new_n22181 = new_n22180 ^ new_n22174;
  assign new_n22182 = new_n22169 ^ new_n22134;
  assign new_n22183 = new_n22154 ^ new_n22134;
  assign new_n22184 = new_n22155 ^ new_n21974;
  assign new_n22185 = new_n22184 ^ new_n22031;
  assign new_n22186 = new_n22183 & new_n22185;
  assign new_n22187 = new_n22186 ^ new_n22139;
  assign new_n22188 = new_n22177 ^ new_n22030;
  assign new_n22189 = new_n22188 ^ new_n22187;
  assign new_n22190 = new_n22189 ^ new_n22182;
  assign new_n22191 = ~new_n22181 & new_n22190;
  assign new_n22192 = new_n22191 ^ new_n22170;
  assign new_n22193 = new_n22192 ^ new_n22142;
  assign new_n22194 = new_n22177 ^ new_n22136;
  assign new_n22195 = new_n22171 ^ new_n22158;
  assign new_n22196 = new_n22195 ^ new_n22194;
  assign new_n22197 = ~new_n22193 & ~new_n22196;
  assign new_n22198 = new_n22197 ^ new_n22191;
  assign new_n22199 = ~new_n22162 & ~new_n22198;
  assign new_n22200 = new_n22199 ^ new_n22197;
  assign new_n22201 = new_n22191 ^ new_n22162;
  assign new_n22202 = new_n22088 ^ new_n21882;
  assign new_n22203 = new_n22186 ^ new_n22164;
  assign new_n22204 = new_n22203 ^ new_n22194;
  assign new_n22205 = new_n22204 ^ new_n22202;
  assign new_n22206 = ~new_n22205 & new_n22201;
  assign new_n22207 = new_n22206 ^ new_n22170;
  assign new_n22208 = new_n22207 ^ new_n22142;
  assign new_n22209 = ~new_n22200 & ~new_n22208;
  assign new_n22210 = new_n22209 ^ new_n22206;
  assign new_n22211 = new_n22210 ^ new_n22190;
  assign new_n22212 = ~new_n21975 & new_n22211;
  assign new_n22213 = new_n22197 ^ new_n21882;
  assign new_n22214 = new_n22164 ^ new_n22158;
  assign new_n22215 = new_n22088 ^ new_n21974;
  assign new_n22216 = new_n22186 ^ new_n22172;
  assign new_n22217 = new_n22201 ^ new_n22200;
  assign new_n22218 = new_n22217 ^ new_n22209;
  assign new_n22219 = new_n22218 ^ new_n22216;
  assign new_n22220 = new_n22219 ^ new_n22215;
  assign new_n22221 = new_n22220 ^ new_n22214;
  assign new_n22222 = new_n22221 ^ new_n22213;
  assign new_n22223 = ~new_n22135 & ~new_n22222;
  assign new_n22224 = new_n22223 ^ new_n22212;
  assign new_n22225 = new_n22220 ^ new_n22108;
  assign new_n22226 = new_n22206 ^ new_n22159;
  assign new_n22227 = new_n22226 ^ new_n22169;
  assign new_n22228 = new_n22227 ^ new_n22225;
  assign new_n22229 = ~new_n22176 & new_n22228;
  assign new_n22230 = new_n22209 ^ new_n22205;
  assign new_n22231 = ~new_n22155 & ~new_n22230;
  assign new_n22232 = new_n22231 ^ new_n22229;
  assign new_n22233 = ~new_n22230 & new_n22184;
  assign new_n22234 = ~new_n22157 & ~new_n22208;
  assign new_n22235 = new_n22234 ^ new_n22233;
  assign new_n22236 = new_n22166 & new_n22228;
  assign new_n22237 = new_n22206 ^ new_n22197;
  assign new_n22238 = new_n22170 ^ new_n22161;
  assign new_n22239 = new_n22238 ^ new_n22237;
  assign new_n22240 = ~new_n22239 & new_n22109;
  assign new_n22241 = new_n22240 ^ new_n22236;
  assign new_n22242 = new_n22241 ^ new_n22235;
  assign new_n22243 = new_n22242 ^ new_n22232;
  assign new_n22244 = new_n22243 ^ new_n22224;
  assign new_n22245 = new_n22244 ^ new_n21200;
  assign new_n22246 = new_n22245 ^ new_n21073;
  assign new_n22247 = new_n21155 ^ new_n21135;
  assign new_n22248 = new_n22247 ^ new_n21134;
  assign new_n22249 = new_n21108 & new_n22248;
  assign new_n22250 = new_n22249 ^ new_n21182;
  assign new_n22251 = new_n22250 ^ new_n21172;
  assign new_n22252 = ~new_n21163 & new_n21115;
  assign new_n22253 = new_n22252 ^ new_n22251;
  assign new_n22254 = new_n22253 ^ new_n21170;
  assign new_n22255 = ~new_n21103 & new_n21179;
  assign new_n22256 = new_n21155 ^ new_n21122;
  assign new_n22257 = ~new_n21093 & new_n22256;
  assign new_n22258 = new_n22257 ^ new_n22255;
  assign new_n22259 = new_n22258 ^ new_n22254;
  assign new_n22260 = new_n20957 ^ new_n19516;
  assign new_n22261 = new_n22260 ^ new_n22259;
  assign new_n22262 = new_n20008 ^ new_n18907;
  assign new_n22263 = new_n18855 & new_n20002;
  assign new_n22264 = new_n22263 ^ new_n19994;
  assign new_n22265 = new_n22264 ^ new_n20009;
  assign new_n22266 = new_n22265 ^ new_n20004;
  assign new_n22267 = new_n22266 ^ new_n22262;
  assign new_n22268 = new_n21055 ^ new_n21035;
  assign new_n22269 = new_n20997 & new_n21065;
  assign new_n22270 = new_n22269 ^ new_n21193;
  assign new_n22271 = new_n22270 ^ new_n21041;
  assign new_n22272 = new_n22271 ^ new_n21067;
  assign new_n22273 = new_n22272 ^ new_n22268;
  assign new_n22274 = new_n22273 ^ new_n22267;
  assign new_n22275 = new_n22274 ^ new_n22261;
  assign new_n22276 = new_n19959 ^ new_n19939;
  assign new_n22277 = new_n22276 ^ new_n19938;
  assign new_n22278 = new_n19903 & new_n22277;
  assign new_n22279 = new_n22278 ^ new_n19986;
  assign new_n22280 = new_n22279 ^ new_n19976;
  assign new_n22281 = new_n19918 & new_n19967;
  assign new_n22282 = new_n22281 ^ new_n22280;
  assign new_n22283 = new_n22282 ^ new_n19974;
  assign new_n22284 = new_n19906 & new_n19983;
  assign new_n22285 = new_n19959 ^ new_n19926;
  assign new_n22286 = new_n19896 & new_n22285;
  assign new_n22287 = new_n22286 ^ new_n22284;
  assign new_n22288 = new_n22287 ^ new_n22283;
  assign new_n22289 = new_n22141 & new_n22211;
  assign new_n22290 = new_n22217 ^ new_n22197;
  assign new_n22291 = new_n22290 ^ new_n22196;
  assign new_n22292 = new_n22185 & new_n22291;
  assign new_n22293 = new_n22292 ^ new_n22241;
  assign new_n22294 = new_n22293 ^ new_n22231;
  assign new_n22295 = new_n22294 ^ new_n22289;
  assign new_n22296 = new_n22295 ^ new_n22229;
  assign new_n22297 = ~new_n22239 & new_n22138;
  assign new_n22298 = new_n22217 ^ new_n22181;
  assign new_n22299 = ~new_n22167 & new_n22298;
  assign new_n22300 = new_n22299 ^ new_n22297;
  assign new_n22301 = new_n22300 ^ new_n22296;
  assign new_n22302 = new_n22301 ^ new_n22288;
  assign new_n22303 = new_n22302 ^ new_n20011;
  assign new_n22304 = new_n22303 ^ new_n22275;
  assign new_n22305 = new_n22304 ^ new_n22246;
  assign new_n22306 = new_n22271 ^ new_n21069;
  assign new_n22307 = new_n22265 ^ new_n20006;
  assign new_n22308 = new_n22307 ^ new_n22306;
  assign new_n22309 = new_n20008 ^ new_n18917;
  assign new_n22310 = ~new_n18714 & new_n18900;
  assign new_n22311 = ~new_n18834 & new_n18886;
  assign new_n22312 = new_n22311 ^ new_n18901;
  assign new_n22313 = new_n22312 ^ new_n19996;
  assign new_n22314 = new_n22313 ^ new_n22310;
  assign new_n22315 = new_n22314 ^ new_n22309;
  assign new_n22316 = new_n22315 ^ new_n22308;
  assign new_n22317 = new_n22255 ^ new_n21180;
  assign new_n22318 = ~new_n21129 & new_n21153;
  assign new_n22319 = new_n22318 ^ new_n21161;
  assign new_n22320 = new_n21142 ^ new_n21135;
  assign new_n22321 = new_n21085 & new_n22320;
  assign new_n22322 = ~new_n21083 & new_n22256;
  assign new_n22323 = new_n22322 ^ new_n22321;
  assign new_n22324 = new_n22323 ^ new_n21164;
  assign new_n22325 = new_n22324 ^ new_n22319;
  assign new_n22326 = ~new_n21160 & new_n21092;
  assign new_n22327 = new_n22326 ^ new_n22325;
  assign new_n22328 = new_n22327 ^ new_n22317;
  assign new_n22329 = new_n20927 ^ new_n19501;
  assign new_n22330 = new_n22329 ^ new_n22328;
  assign new_n22331 = new_n22284 ^ new_n19984;
  assign new_n22332 = new_n19933 & new_n19957;
  assign new_n22333 = new_n22332 ^ new_n19965;
  assign new_n22334 = new_n19946 ^ new_n19939;
  assign new_n22335 = new_n19870 & new_n22334;
  assign new_n22336 = new_n19858 & new_n22285;
  assign new_n22337 = new_n22336 ^ new_n22335;
  assign new_n22338 = new_n22337 ^ new_n19968;
  assign new_n22339 = new_n22338 ^ new_n22333;
  assign new_n22340 = new_n19895 & new_n19964;
  assign new_n22341 = new_n22340 ^ new_n22339;
  assign new_n22342 = new_n22341 ^ new_n22331;
  assign new_n22343 = new_n22342 ^ new_n22330;
  assign new_n22344 = new_n22297 ^ new_n22240;
  assign new_n22345 = ~new_n22156 & ~new_n22208;
  assign new_n22346 = new_n22345 ^ new_n22223;
  assign new_n22347 = new_n22197 ^ new_n22162;
  assign new_n22348 = ~new_n22154 & new_n22347;
  assign new_n22349 = ~new_n22134 & new_n22298;
  assign new_n22350 = new_n22349 ^ new_n22348;
  assign new_n22351 = new_n22350 ^ new_n22212;
  assign new_n22352 = new_n22351 ^ new_n22346;
  assign new_n22353 = ~new_n22222 & new_n22031;
  assign new_n22354 = new_n22353 ^ new_n22352;
  assign new_n22355 = new_n22354 ^ new_n22344;
  assign new_n22356 = new_n22355 ^ new_n22343;
  assign new_n22357 = new_n22356 ^ new_n22316;
  assign new_n22358 = new_n22357 ^ new_n22304;
  assign new_n22359 = new_n22324 ^ new_n22252;
  assign new_n22360 = new_n22359 ^ new_n21183;
  assign new_n22361 = new_n20936 ^ new_n19494;
  assign new_n22362 = new_n22361 ^ new_n22360;
  assign new_n22363 = new_n22362 ^ new_n19999;
  assign new_n22364 = new_n22351 ^ new_n22289;
  assign new_n22365 = new_n22364 ^ new_n22242;
  assign new_n22366 = new_n22338 ^ new_n22281;
  assign new_n22367 = new_n22366 ^ new_n19987;
  assign new_n22368 = new_n22367 ^ new_n22365;
  assign new_n22369 = new_n22368 ^ new_n21072;
  assign new_n22370 = new_n22369 ^ new_n22363;
  assign new_n22371 = new_n22299 ^ new_n22234;
  assign new_n22372 = new_n22183 & new_n22291;
  assign new_n22373 = new_n22372 ^ new_n22348;
  assign new_n22374 = new_n22373 ^ new_n22294;
  assign new_n22375 = new_n22374 ^ new_n22371;
  assign new_n22376 = new_n20009 ^ new_n18912;
  assign new_n22377 = new_n22263 ^ new_n19992;
  assign new_n22378 = new_n22377 ^ new_n20005;
  assign new_n22379 = new_n22378 ^ new_n22376;
  assign new_n22380 = new_n22379 ^ new_n22375;
  assign new_n22381 = new_n22286 ^ new_n19979;
  assign new_n22382 = new_n19901 & new_n22277;
  assign new_n22383 = new_n22382 ^ new_n22335;
  assign new_n22384 = new_n22383 ^ new_n22280;
  assign new_n22385 = new_n22384 ^ new_n22381;
  assign new_n22386 = new_n22385 ^ new_n22380;
  assign new_n22387 = new_n22257 ^ new_n21175;
  assign new_n22388 = ~new_n21106 & new_n22248;
  assign new_n22389 = new_n22388 ^ new_n22321;
  assign new_n22390 = new_n22389 ^ new_n22251;
  assign new_n22391 = new_n22390 ^ new_n22387;
  assign new_n22392 = new_n20798 ^ new_n19479;
  assign new_n22393 = new_n22392 ^ new_n22391;
  assign new_n22394 = new_n22393 ^ new_n21072;
  assign new_n22395 = new_n18841 & new_n19991;
  assign new_n22396 = new_n22395 ^ new_n20007;
  assign new_n22397 = new_n22396 ^ new_n22313;
  assign new_n22398 = new_n21031 ^ new_n20961;
  assign new_n22399 = new_n21019 ^ new_n21008;
  assign new_n22400 = new_n22399 ^ new_n21050;
  assign new_n22401 = new_n22400 ^ new_n22398;
  assign new_n22402 = ~new_n21011 & ~new_n22401;
  assign new_n22403 = ~new_n21006 & ~new_n21046;
  assign new_n22404 = new_n22403 ^ new_n22402;
  assign new_n22405 = new_n22404 ^ new_n21197;
  assign new_n22406 = ~new_n21018 & new_n21194;
  assign new_n22407 = new_n22406 ^ new_n21070;
  assign new_n22408 = new_n22407 ^ new_n22405;
  assign new_n22409 = new_n22408 ^ new_n22397;
  assign new_n22410 = new_n22409 ^ new_n22394;
  assign new_n22411 = new_n22410 ^ new_n22386;
  assign new_n22412 = new_n22411 ^ new_n22246;
  assign new_n22413 = new_n22388 ^ new_n22322;
  assign new_n22414 = new_n22413 ^ new_n22257;
  assign new_n22415 = new_n22414 ^ new_n22253;
  assign new_n22416 = new_n20971 ^ new_n19507;
  assign new_n22417 = new_n22416 ^ new_n22415;
  assign new_n22418 = new_n22417 ^ new_n21072;
  assign new_n22419 = new_n21189 ^ new_n21041;
  assign new_n22420 = new_n22269 ^ new_n21195;
  assign new_n22421 = new_n22420 ^ new_n21068;
  assign new_n22422 = new_n22421 ^ new_n22419;
  assign new_n22423 = new_n22422 ^ new_n22379;
  assign new_n22424 = new_n22423 ^ new_n22418;
  assign new_n22425 = new_n22382 ^ new_n22336;
  assign new_n22426 = new_n22425 ^ new_n22286;
  assign new_n22427 = new_n22426 ^ new_n22282;
  assign new_n22428 = new_n22427 ^ new_n22307;
  assign new_n22429 = new_n22372 ^ new_n22349;
  assign new_n22430 = new_n22429 ^ new_n22299;
  assign new_n22431 = new_n22430 ^ new_n22295;
  assign new_n22432 = new_n22431 ^ new_n22428;
  assign new_n22433 = new_n22432 ^ new_n22424;
  assign new_n22434 = new_n22433 ^ new_n22304;
  assign new_n22435 = new_n22434 ^ new_n22412;
  assign new_n22436 = new_n22435 ^ new_n22370;
  assign new_n22437 = new_n21061 ^ new_n21035;
  assign new_n22438 = ~new_n22401 & new_n20965;
  assign new_n22439 = new_n22438 ^ new_n22405;
  assign new_n22440 = new_n22439 ^ new_n22437;
  assign new_n22441 = new_n22440 ^ new_n22315;
  assign new_n22442 = new_n22441 ^ new_n22267;
  assign new_n22443 = new_n22255 ^ new_n21170;
  assign new_n22444 = new_n22414 ^ new_n22250;
  assign new_n22445 = new_n22444 ^ new_n22443;
  assign new_n22446 = new_n20898 ^ new_n19467;
  assign new_n22447 = new_n22446 ^ new_n22445;
  assign new_n22448 = new_n22284 ^ new_n19974;
  assign new_n22449 = new_n22426 ^ new_n22279;
  assign new_n22450 = new_n22449 ^ new_n22448;
  assign new_n22451 = new_n22450 ^ new_n22447;
  assign new_n22452 = new_n22297 ^ new_n22229;
  assign new_n22453 = new_n22430 ^ new_n22293;
  assign new_n22454 = new_n22453 ^ new_n22452;
  assign new_n22455 = new_n22454 ^ new_n22451;
  assign new_n22456 = new_n22455 ^ new_n22442;
  assign new_n22457 = new_n22456 ^ new_n22357;
  assign new_n22458 = new_n22457 ^ new_n22370;
  assign new_n22459 = new_n22458 ^ new_n22246;
  assign new_n22460 = ~new_n22163 & new_n22347;
  assign new_n22461 = new_n22460 ^ new_n22296;
  assign new_n22462 = new_n22461 ^ new_n22352;
  assign new_n22463 = new_n22462 ^ new_n22397;
  assign new_n22464 = new_n19872 & new_n22334;
  assign new_n22465 = new_n22464 ^ new_n22283;
  assign new_n22466 = new_n22465 ^ new_n22339;
  assign new_n22467 = new_n22466 ^ new_n22463;
  assign new_n22468 = ~new_n21087 & new_n22320;
  assign new_n22469 = new_n22468 ^ new_n22254;
  assign new_n22470 = new_n22469 ^ new_n22325;
  assign new_n22471 = new_n20430 ^ new_n19474;
  assign new_n22472 = new_n22471 ^ new_n22470;
  assign new_n22473 = new_n22402 ^ new_n21192;
  assign new_n22474 = new_n21060 ^ new_n21055;
  assign new_n22475 = new_n22474 ^ new_n21191;
  assign new_n22476 = new_n22475 ^ new_n22473;
  assign new_n22477 = new_n22476 ^ new_n18922;
  assign new_n22478 = new_n22477 ^ new_n22472;
  assign new_n22479 = new_n22478 ^ new_n22467;
  assign new_n22480 = new_n22479 ^ new_n22304;
  assign new_n22481 = new_n22480 ^ new_n22459;
  assign new_n22482 = new_n22436 & new_n22481;
  assign new_n22483 = new_n22458 ^ new_n22433;
  assign new_n22484 = new_n22370 & new_n22483;
  assign new_n22485 = new_n22484 ^ new_n22482;
  assign new_n22486 = new_n22479 ^ new_n22433;
  assign new_n22487 = new_n22433 ^ new_n22357;
  assign new_n22488 = new_n22487 ^ new_n22480;
  assign new_n22489 = new_n22486 & new_n22488;
  assign new_n22490 = new_n22457 ^ new_n22435;
  assign new_n22491 = new_n22480 & new_n22490;
  assign new_n22492 = new_n22491 ^ new_n22489;
  assign new_n22493 = new_n22492 ^ new_n22485;
  assign new_n22494 = new_n22493 ^ new_n22358;
  assign new_n22495 = ~new_n22246 & ~new_n22458;
  assign new_n22496 = new_n22495 ^ new_n22246;
  assign new_n22497 = new_n22479 ^ new_n22412;
  assign new_n22498 = new_n22497 ^ new_n22357;
  assign new_n22499 = new_n22305 & new_n22498;
  assign new_n22500 = new_n22499 ^ new_n22496;
  assign new_n22501 = new_n22500 ^ new_n22480;
  assign new_n22502 = new_n22497 ^ new_n22456;
  assign new_n22503 = new_n22434 & new_n22502;
  assign new_n22504 = new_n22503 ^ new_n22489;
  assign new_n22505 = new_n22411 ^ new_n22357;
  assign new_n22506 = new_n22505 ^ new_n22504;
  assign new_n22507 = new_n22506 ^ new_n22501;
  assign new_n22508 = new_n22486 ^ new_n22305;
  assign new_n22509 = new_n22435 & new_n22508;
  assign new_n22510 = new_n22509 ^ new_n22456;
  assign new_n22511 = new_n22510 ^ new_n22435;
  assign new_n22512 = new_n22503 ^ new_n22482;
  assign new_n22513 = new_n22489 ^ new_n22479;
  assign new_n22514 = new_n22513 ^ new_n22512;
  assign new_n22515 = new_n22514 ^ new_n22511;
  assign new_n22516 = ~new_n22507 & new_n22515;
  assign new_n22517 = new_n22503 ^ new_n22491;
  assign new_n22518 = new_n22517 ^ new_n22498;
  assign new_n22519 = new_n22458 ^ new_n22304;
  assign new_n22520 = new_n22502 ^ new_n22370;
  assign new_n22521 = new_n22519 & new_n22520;
  assign new_n22522 = new_n22521 ^ new_n22499;
  assign new_n22523 = new_n22522 ^ new_n22304;
  assign new_n22524 = new_n22523 ^ new_n22518;
  assign new_n22525 = new_n22524 ^ new_n22516;
  assign new_n22526 = new_n22494 & new_n22525;
  assign new_n22527 = new_n22484 ^ new_n22433;
  assign new_n22528 = new_n22527 ^ new_n22510;
  assign new_n22529 = new_n22528 ^ new_n22526;
  assign new_n22530 = new_n22529 ^ new_n22518;
  assign new_n22531 = new_n22528 ^ new_n22516;
  assign new_n22532 = new_n22531 ^ new_n22518;
  assign new_n22533 = new_n22521 ^ new_n22495;
  assign new_n22534 = new_n22533 ^ new_n22492;
  assign new_n22535 = ~new_n22534 & new_n22532;
  assign new_n22536 = new_n22535 ^ new_n22516;
  assign new_n22537 = ~new_n22536 & new_n22524;
  assign new_n22538 = new_n22537 ^ new_n22516;
  assign new_n22539 = new_n22530 & new_n22538;
  assign new_n22540 = new_n22539 ^ new_n22526;
  assign new_n22541 = new_n22540 ^ new_n22515;
  assign new_n22542 = new_n22305 & new_n22541;
  assign new_n22543 = new_n22535 ^ new_n22304;
  assign new_n22544 = new_n22521 ^ new_n22484;
  assign new_n22545 = new_n22357 ^ new_n22246;
  assign new_n22546 = new_n22496 ^ new_n22482;
  assign new_n22547 = new_n22537 ^ new_n22524;
  assign new_n22548 = new_n22547 ^ new_n22539;
  assign new_n22549 = new_n22548 ^ new_n22546;
  assign new_n22550 = new_n22549 ^ new_n22545;
  assign new_n22551 = new_n22550 ^ new_n22544;
  assign new_n22552 = new_n22551 ^ new_n22543;
  assign new_n22553 = ~new_n22552 & new_n22490;
  assign new_n22554 = new_n22553 ^ new_n22542;
  assign new_n22555 = new_n22550 ^ new_n22433;
  assign new_n22556 = new_n22526 ^ new_n22499;
  assign new_n22557 = new_n22556 ^ new_n22510;
  assign new_n22558 = new_n22557 ^ new_n22555;
  assign new_n22559 = ~new_n22558 & new_n22488;
  assign new_n22560 = new_n22539 ^ new_n22494;
  assign new_n22561 = new_n22458 & new_n22560;
  assign new_n22562 = new_n22561 ^ new_n22559;
  assign new_n22563 = new_n22459 & new_n22560;
  assign new_n22564 = new_n22520 & new_n22530;
  assign new_n22565 = new_n22564 ^ new_n22563;
  assign new_n22566 = new_n22535 ^ new_n22526;
  assign new_n22567 = new_n22528 ^ new_n22523;
  assign new_n22568 = new_n22567 ^ new_n22566;
  assign new_n22569 = new_n22434 & new_n22568;
  assign new_n22570 = ~new_n22558 & new_n22486;
  assign new_n22571 = new_n22570 ^ new_n22569;
  assign new_n22572 = new_n22571 ^ new_n22565;
  assign new_n22573 = new_n22572 ^ new_n22562;
  assign new_n22574 = new_n22573 ^ new_n22554;
  assign new_n22575 = new_n22123 ^ new_n598;
  assign new_n22576 = new_n21955 ^ new_n592;
  assign new_n22577 = new_n22576 ^ new_n22575;
  assign new_n22578 = new_n22016 ^ new_n606;
  assign new_n22579 = new_n22578 ^ new_n22577;
  assign new_n22580 = new_n22056 ^ new_n567;
  assign new_n22581 = new_n22580 ^ new_n22579;
  assign new_n22582 = new_n22147 ^ new_n576;
  assign new_n22583 = new_n22079 ^ new_n561;
  assign new_n22584 = new_n22583 ^ new_n22580;
  assign new_n22585 = new_n22584 ^ new_n22582;
  assign new_n22586 = new_n22090 ^ new_n541;
  assign new_n22587 = new_n22586 ^ new_n22585;
  assign new_n22588 = new_n22582 & new_n22587;
  assign new_n22589 = new_n22588 ^ new_n22586;
  assign new_n22590 = new_n21303 ^ new_n585;
  assign new_n22591 = new_n22590 ^ new_n22586;
  assign new_n22592 = new_n22591 ^ new_n22577;
  assign new_n22593 = new_n22586 ^ new_n22576;
  assign new_n22594 = new_n22590 ^ new_n22578;
  assign new_n22595 = new_n22594 ^ new_n22593;
  assign new_n22596 = new_n22592 & new_n22595;
  assign new_n22597 = new_n22596 ^ new_n22580;
  assign new_n22598 = new_n22597 ^ new_n22589;
  assign new_n22599 = ~new_n22576 & ~new_n22585;
  assign new_n22600 = new_n22599 ^ new_n22576;
  assign new_n22601 = new_n22583 ^ new_n22579;
  assign new_n22602 = new_n22590 ^ new_n22576;
  assign new_n22603 = new_n22601 & new_n22602;
  assign new_n22604 = new_n22603 ^ new_n22600;
  assign new_n22605 = new_n22604 ^ new_n22594;
  assign new_n22606 = new_n22581 & new_n22591;
  assign new_n22607 = new_n22586 ^ new_n22583;
  assign new_n22608 = new_n22607 ^ new_n22594;
  assign new_n22609 = new_n22586 ^ new_n22578;
  assign new_n22610 = new_n22608 & new_n22609;
  assign new_n22611 = new_n22610 ^ new_n22606;
  assign new_n22612 = new_n22583 ^ new_n22575;
  assign new_n22613 = new_n22612 ^ new_n22611;
  assign new_n22614 = new_n22613 ^ new_n22605;
  assign new_n22615 = new_n22597 ^ new_n22592;
  assign new_n22616 = new_n22585 ^ new_n22576;
  assign new_n22617 = new_n22616 ^ new_n22594;
  assign new_n22618 = new_n22592 ^ new_n22582;
  assign new_n22619 = new_n22617 & new_n22618;
  assign new_n22620 = new_n22619 ^ new_n22578;
  assign new_n22621 = new_n22620 ^ new_n22611;
  assign new_n22622 = new_n22621 ^ new_n22615;
  assign new_n22623 = ~new_n22614 & new_n22622;
  assign new_n22624 = new_n22623 ^ new_n22598;
  assign new_n22625 = new_n22592 ^ new_n22584;
  assign new_n22626 = new_n22594 & new_n22625;
  assign new_n22627 = new_n22626 ^ new_n22606;
  assign new_n22628 = new_n22627 ^ new_n22601;
  assign new_n22629 = new_n22628 ^ new_n22624;
  assign new_n22630 = new_n22590 ^ new_n22585;
  assign new_n22631 = new_n22582 ^ new_n22581;
  assign new_n22632 = new_n22630 & new_n22631;
  assign new_n22633 = new_n22632 ^ new_n22599;
  assign new_n22634 = new_n22626 ^ new_n22610;
  assign new_n22635 = new_n22634 ^ new_n22633;
  assign new_n22636 = ~new_n22635 & new_n22629;
  assign new_n22637 = new_n22590 ^ new_n22583;
  assign new_n22638 = new_n22619 ^ new_n22588;
  assign new_n22639 = new_n22638 ^ new_n22634;
  assign new_n22640 = new_n22639 ^ new_n22637;
  assign new_n22641 = new_n22632 ^ new_n22603;
  assign new_n22642 = new_n22641 ^ new_n22590;
  assign new_n22643 = new_n22642 ^ new_n22628;
  assign new_n22644 = new_n22643 ^ new_n22623;
  assign new_n22645 = new_n22640 & new_n22644;
  assign new_n22646 = new_n22645 ^ new_n22636;
  assign new_n22647 = new_n22642 ^ new_n22598;
  assign new_n22648 = new_n22647 ^ new_n22646;
  assign new_n22649 = new_n22581 & new_n22648;
  assign new_n22650 = new_n22591 & new_n22648;
  assign new_n22651 = new_n22650 ^ new_n22649;
  assign new_n22652 = new_n22645 ^ new_n22598;
  assign new_n22653 = new_n22652 ^ new_n22628;
  assign new_n22654 = new_n22630 & new_n22653;
  assign new_n22655 = new_n22636 ^ new_n22590;
  assign new_n22656 = new_n22632 ^ new_n22588;
  assign new_n22657 = new_n22583 ^ new_n22576;
  assign new_n22658 = new_n22619 ^ new_n22600;
  assign new_n22659 = new_n22636 ^ new_n22623;
  assign new_n22660 = new_n22643 & new_n22659;
  assign new_n22661 = new_n22660 ^ new_n22644;
  assign new_n22662 = new_n22653 & new_n22661;
  assign new_n22663 = new_n22662 ^ new_n22660;
  assign new_n22664 = new_n22663 ^ new_n22658;
  assign new_n22665 = new_n22664 ^ new_n22657;
  assign new_n22666 = new_n22665 ^ new_n22656;
  assign new_n22667 = new_n22666 ^ new_n22655;
  assign new_n22668 = ~new_n22667 & new_n22625;
  assign new_n22669 = new_n22668 ^ new_n22654;
  assign new_n22670 = new_n22660 ^ new_n22614;
  assign new_n22671 = ~new_n22670 & new_n22592;
  assign new_n22672 = new_n22643 ^ new_n22636;
  assign new_n22673 = new_n22582 & new_n22672;
  assign new_n22674 = new_n22673 ^ new_n22671;
  assign new_n22675 = new_n22662 ^ new_n22645;
  assign new_n22676 = new_n22675 ^ new_n22622;
  assign new_n22677 = new_n22602 & new_n22676;
  assign new_n22678 = new_n22677 ^ new_n22674;
  assign new_n22679 = new_n22678 ^ new_n22669;
  assign new_n22680 = ~new_n22667 & new_n22594;
  assign new_n22681 = new_n22680 ^ new_n22679;
  assign new_n22682 = new_n22681 ^ new_n22651;
  assign new_n22683 = new_n22682 ^ new_n19652;
  assign new_n22684 = new_n22683 ^ new_n7912;
  assign new_n22685 = new_n22130 ^ new_n21896;
  assign new_n22686 = new_n18670 ^ new_n16499;
  assign new_n22687 = new_n22686 ^ new_n4753;
  assign new_n22688 = new_n22687 ^ new_n21986;
  assign new_n22689 = new_n22688 ^ new_n21971;
  assign new_n22690 = new_n22689 ^ new_n22685;
  assign new_n22691 = new_n22113 ^ new_n21986;
  assign new_n22692 = new_n22691 ^ new_n22004;
  assign new_n22693 = new_n18793 ^ new_n17185;
  assign new_n22694 = new_n22693 ^ new_n4777;
  assign new_n22695 = new_n22694 ^ new_n22102;
  assign new_n22696 = new_n21880 ^ new_n21736;
  assign new_n22697 = new_n22696 ^ new_n22695;
  assign new_n22698 = new_n22697 ^ new_n22692;
  assign new_n22699 = new_n22144 ^ new_n22028;
  assign new_n22700 = new_n22699 ^ new_n22696;
  assign new_n22701 = new_n18634 ^ new_n17165;
  assign new_n22702 = new_n22701 ^ new_n4704;
  assign new_n22703 = new_n22702 ^ new_n22151;
  assign new_n22704 = new_n22703 ^ new_n21896;
  assign new_n22705 = new_n22704 ^ new_n22700;
  assign new_n22706 = new_n22705 ^ new_n22698;
  assign new_n22707 = new_n22706 ^ new_n22690;
  assign new_n22708 = new_n22071 ^ new_n21581;
  assign new_n22709 = new_n18765 ^ new_n17241;
  assign new_n22710 = new_n22709 ^ new_n4634;
  assign new_n22711 = new_n22710 ^ new_n22085;
  assign new_n22712 = new_n22711 ^ new_n22037;
  assign new_n22713 = new_n22712 ^ new_n22708;
  assign new_n22714 = new_n22713 ^ new_n22707;
  assign new_n22715 = new_n18823 ^ new_n17298;
  assign new_n22716 = new_n22715 ^ new_n4664;
  assign new_n22717 = new_n22716 ^ new_n22144;
  assign new_n22718 = new_n22696 ^ new_n21931;
  assign new_n22719 = new_n22718 ^ new_n22717;
  assign new_n22720 = new_n18771 ^ new_n17315;
  assign new_n22721 = new_n22720 ^ new_n1403;
  assign new_n22722 = new_n22721 ^ new_n22074;
  assign new_n22723 = new_n22722 ^ new_n22696;
  assign new_n22724 = new_n22113 ^ new_n22106;
  assign new_n22725 = new_n22724 ^ new_n22118;
  assign new_n22726 = new_n22725 ^ new_n22723;
  assign new_n22727 = new_n18718 ^ new_n17269;
  assign new_n22728 = new_n22727 ^ new_n4616;
  assign new_n22729 = new_n22106 ^ new_n22104;
  assign new_n22730 = new_n22729 ^ new_n22728;
  assign new_n22731 = new_n22071 ^ new_n22049;
  assign new_n22732 = new_n22731 ^ new_n22730;
  assign new_n22733 = new_n22732 ^ new_n22713;
  assign new_n22734 = new_n22733 ^ new_n22719;
  assign new_n22735 = new_n22734 ^ new_n22726;
  assign new_n22736 = new_n22719 & new_n22735;
  assign new_n22737 = new_n22736 ^ new_n22726;
  assign new_n22738 = new_n22037 ^ new_n21907;
  assign new_n22739 = new_n17678 ^ new_n17290;
  assign new_n22740 = new_n22739 ^ new_n4732;
  assign new_n22741 = new_n22740 ^ new_n21880;
  assign new_n22742 = new_n22741 ^ new_n22064;
  assign new_n22743 = new_n22742 ^ new_n22738;
  assign new_n22744 = new_n22743 ^ new_n22726;
  assign new_n22745 = new_n22744 ^ new_n22706;
  assign new_n22746 = new_n22726 ^ new_n22705;
  assign new_n22747 = new_n22743 ^ new_n22690;
  assign new_n22748 = new_n22747 ^ new_n22746;
  assign new_n22749 = ~new_n22745 & ~new_n22748;
  assign new_n22750 = new_n22749 ^ new_n22713;
  assign new_n22751 = new_n22750 ^ new_n22737;
  assign new_n22752 = ~new_n22705 & new_n22734;
  assign new_n22753 = new_n22752 ^ new_n22705;
  assign new_n22754 = new_n22743 ^ new_n22705;
  assign new_n22755 = new_n22732 ^ new_n22707;
  assign new_n22756 = new_n22754 & new_n22755;
  assign new_n22757 = new_n22756 ^ new_n22753;
  assign new_n22758 = new_n22757 ^ new_n22747;
  assign new_n22759 = ~new_n22714 & ~new_n22744;
  assign new_n22760 = new_n22732 ^ new_n22726;
  assign new_n22761 = new_n22760 ^ new_n22747;
  assign new_n22762 = new_n22726 ^ new_n22690;
  assign new_n22763 = ~new_n22761 & ~new_n22762;
  assign new_n22764 = new_n22763 ^ new_n22759;
  assign new_n22765 = new_n22732 ^ new_n22698;
  assign new_n22766 = new_n22765 ^ new_n22764;
  assign new_n22767 = new_n22766 ^ new_n22758;
  assign new_n22768 = new_n22750 ^ new_n22745;
  assign new_n22769 = new_n22745 ^ new_n22719;
  assign new_n22770 = new_n22734 ^ new_n22705;
  assign new_n22771 = new_n22770 ^ new_n22747;
  assign new_n22772 = ~new_n22769 & ~new_n22771;
  assign new_n22773 = new_n22772 ^ new_n22764;
  assign new_n22774 = new_n22773 ^ new_n22690;
  assign new_n22775 = new_n22774 ^ new_n22768;
  assign new_n22776 = ~new_n22767 & new_n22775;
  assign new_n22777 = new_n22776 ^ new_n22751;
  assign new_n22778 = new_n22745 ^ new_n22733;
  assign new_n22779 = new_n22747 & new_n22778;
  assign new_n22780 = new_n22779 ^ new_n22759;
  assign new_n22781 = new_n22780 ^ new_n22755;
  assign new_n22782 = new_n22781 ^ new_n22777;
  assign new_n22783 = new_n22743 ^ new_n22734;
  assign new_n22784 = new_n22719 ^ new_n22714;
  assign new_n22785 = ~new_n22783 & ~new_n22784;
  assign new_n22786 = new_n22785 ^ new_n22752;
  assign new_n22787 = new_n22779 ^ new_n22763;
  assign new_n22788 = new_n22787 ^ new_n22786;
  assign new_n22789 = ~new_n22788 & new_n22782;
  assign new_n22790 = new_n22743 ^ new_n22732;
  assign new_n22791 = new_n22772 ^ new_n22736;
  assign new_n22792 = new_n22791 ^ new_n22787;
  assign new_n22793 = new_n22792 ^ new_n22790;
  assign new_n22794 = new_n22785 ^ new_n22756;
  assign new_n22795 = new_n22794 ^ new_n22743;
  assign new_n22796 = new_n22795 ^ new_n22781;
  assign new_n22797 = new_n22796 ^ new_n22776;
  assign new_n22798 = new_n22793 & new_n22797;
  assign new_n22799 = new_n22798 ^ new_n22789;
  assign new_n22800 = new_n22795 ^ new_n22751;
  assign new_n22801 = new_n22800 ^ new_n22799;
  assign new_n22802 = ~new_n22714 & new_n22801;
  assign new_n22803 = ~new_n22744 & new_n22801;
  assign new_n22804 = new_n22803 ^ new_n22802;
  assign new_n22805 = new_n22789 ^ new_n22743;
  assign new_n22806 = new_n22785 ^ new_n22736;
  assign new_n22807 = new_n22732 ^ new_n22705;
  assign new_n22808 = new_n22772 ^ new_n22753;
  assign new_n22809 = new_n22798 ^ new_n22751;
  assign new_n22810 = new_n22809 ^ new_n22781;
  assign new_n22811 = new_n22789 ^ new_n22776;
  assign new_n22812 = new_n22796 & new_n22811;
  assign new_n22813 = new_n22812 ^ new_n22797;
  assign new_n22814 = new_n22810 & new_n22813;
  assign new_n22815 = new_n22814 ^ new_n22812;
  assign new_n22816 = new_n22815 ^ new_n22808;
  assign new_n22817 = new_n22816 ^ new_n22807;
  assign new_n22818 = new_n22817 ^ new_n22806;
  assign new_n22819 = new_n22818 ^ new_n22805;
  assign new_n22820 = ~new_n22819 & new_n22747;
  assign new_n22821 = ~new_n22783 & new_n22810;
  assign new_n22822 = ~new_n22819 & new_n22778;
  assign new_n22823 = new_n22822 ^ new_n22821;
  assign new_n22824 = new_n22812 ^ new_n22767;
  assign new_n22825 = ~new_n22745 & ~new_n22824;
  assign new_n22826 = new_n22796 ^ new_n22789;
  assign new_n22827 = new_n22719 & new_n22826;
  assign new_n22828 = new_n22827 ^ new_n22825;
  assign new_n22829 = new_n22814 ^ new_n22798;
  assign new_n22830 = new_n22829 ^ new_n22775;
  assign new_n22831 = new_n22754 & new_n22830;
  assign new_n22832 = new_n22831 ^ new_n22828;
  assign new_n22833 = new_n22832 ^ new_n22823;
  assign new_n22834 = new_n22833 ^ new_n22820;
  assign new_n22835 = new_n22834 ^ new_n22804;
  assign new_n22836 = new_n22835 ^ new_n22684;
  assign new_n22837 = new_n19731 ^ new_n6844;
  assign new_n22838 = new_n22837 ^ new_n20777;
  assign new_n22839 = new_n20950 ^ new_n20790;
  assign new_n22840 = new_n22839 ^ new_n20882;
  assign new_n22841 = new_n22840 ^ new_n22838;
  assign new_n22842 = new_n19775 ^ new_n7594;
  assign new_n22843 = new_n22842 ^ new_n20951;
  assign new_n22844 = new_n20967 ^ new_n20921;
  assign new_n22845 = new_n22844 ^ new_n22843;
  assign new_n22846 = new_n20922 ^ new_n20828;
  assign new_n22847 = new_n22846 ^ new_n22845;
  assign new_n22848 = new_n22847 ^ new_n22841;
  assign new_n22849 = new_n20951 ^ new_n20940;
  assign new_n22850 = new_n22849 ^ new_n20313;
  assign new_n22851 = new_n19818 ^ new_n7465;
  assign new_n22852 = new_n22851 ^ new_n20849;
  assign new_n22853 = new_n22852 ^ new_n20934;
  assign new_n22854 = new_n22853 ^ new_n22850;
  assign new_n22855 = new_n20827 ^ new_n20591;
  assign new_n22856 = new_n22855 ^ new_n20771;
  assign new_n22857 = new_n19834 ^ new_n7623;
  assign new_n22858 = new_n22857 ^ new_n20951;
  assign new_n22859 = new_n22858 ^ new_n20978;
  assign new_n22860 = new_n22859 ^ new_n22856;
  assign new_n22861 = new_n22860 ^ new_n22854;
  assign new_n22862 = new_n22861 ^ new_n22848;
  assign new_n22863 = new_n19861 ^ new_n7649;
  assign new_n22864 = new_n22863 ^ new_n20934;
  assign new_n22865 = new_n20951 ^ new_n20841;
  assign new_n22866 = new_n22865 ^ new_n22864;
  assign new_n22867 = new_n22866 ^ new_n22862;
  assign new_n22868 = new_n20865 ^ new_n20812;
  assign new_n22869 = new_n19878 ^ new_n7523;
  assign new_n22870 = new_n22869 ^ new_n20591;
  assign new_n22871 = new_n22870 ^ new_n20849;
  assign new_n22872 = new_n22871 ^ new_n22868;
  assign new_n22873 = new_n22872 ^ new_n22861;
  assign new_n22874 = new_n19029 ^ new_n7541;
  assign new_n22875 = new_n22874 ^ new_n20892;
  assign new_n22876 = new_n20954 ^ new_n20875;
  assign new_n22877 = new_n22876 ^ new_n20916;
  assign new_n22878 = new_n22877 ^ new_n22875;
  assign new_n22879 = new_n22878 ^ new_n22873;
  assign new_n22880 = new_n22848 & new_n22879;
  assign new_n22881 = new_n22872 ^ new_n22841;
  assign new_n22882 = new_n19652 ^ new_n7575;
  assign new_n22883 = new_n22882 ^ new_n20904;
  assign new_n22884 = new_n20911 ^ new_n20886;
  assign new_n22885 = new_n22884 ^ new_n20969;
  assign new_n22886 = new_n22885 ^ new_n22883;
  assign new_n22887 = new_n22886 ^ new_n22878;
  assign new_n22888 = new_n22887 ^ new_n22862;
  assign new_n22889 = ~new_n22888 & new_n22881;
  assign new_n22890 = new_n22889 ^ new_n22880;
  assign new_n22891 = new_n22886 ^ new_n22873;
  assign new_n22892 = new_n22891 ^ new_n22890;
  assign new_n22893 = new_n22879 ^ new_n22866;
  assign new_n22894 = new_n22887 ^ new_n22866;
  assign new_n22895 = new_n22894 ^ new_n22841;
  assign new_n22896 = ~new_n22893 & ~new_n22895;
  assign new_n22897 = new_n22854 ^ new_n22841;
  assign new_n22898 = ~new_n22897 & new_n22891;
  assign new_n22899 = new_n22898 ^ new_n22896;
  assign new_n22900 = new_n22899 ^ new_n22841;
  assign new_n22901 = new_n22900 ^ new_n22892;
  assign new_n22902 = new_n22872 ^ new_n22847;
  assign new_n22903 = new_n22902 ^ new_n22897;
  assign new_n22904 = ~new_n22862 & ~new_n22903;
  assign new_n22905 = new_n22904 ^ new_n22878;
  assign new_n22906 = ~new_n22866 & ~new_n22887;
  assign new_n22907 = new_n22847 & new_n22866;
  assign new_n22908 = new_n22907 ^ new_n22906;
  assign new_n22909 = new_n22908 ^ new_n22905;
  assign new_n22910 = new_n22854 & new_n22894;
  assign new_n22911 = new_n22910 ^ new_n22854;
  assign new_n22912 = new_n22911 ^ new_n22898;
  assign new_n22913 = new_n22912 ^ new_n22881;
  assign new_n22914 = new_n22886 ^ new_n22847;
  assign new_n22915 = new_n22914 ^ new_n22881;
  assign new_n22916 = ~new_n22915 & new_n22902;
  assign new_n22917 = new_n22916 ^ new_n22880;
  assign new_n22918 = new_n22886 ^ new_n22860;
  assign new_n22919 = new_n22918 ^ new_n22917;
  assign new_n22920 = new_n22919 ^ new_n22913;
  assign new_n22921 = new_n22905 ^ new_n22862;
  assign new_n22922 = new_n22894 ^ new_n22854;
  assign new_n22923 = new_n22922 ^ new_n22881;
  assign new_n22924 = new_n22867 & new_n22923;
  assign new_n22925 = new_n22924 ^ new_n22917;
  assign new_n22926 = new_n22925 ^ new_n22872;
  assign new_n22927 = new_n22926 ^ new_n22921;
  assign new_n22928 = ~new_n22920 & new_n22927;
  assign new_n22929 = new_n22928 ^ new_n22909;
  assign new_n22930 = new_n22929 ^ new_n22892;
  assign new_n22931 = new_n22910 ^ new_n22896;
  assign new_n22932 = new_n22916 ^ new_n22889;
  assign new_n22933 = new_n22932 ^ new_n22931;
  assign new_n22934 = ~new_n22930 & ~new_n22933;
  assign new_n22935 = new_n22934 ^ new_n22928;
  assign new_n22936 = new_n22901 & new_n22935;
  assign new_n22937 = new_n22936 ^ new_n22934;
  assign new_n22938 = new_n22937 ^ new_n22933;
  assign new_n22939 = ~new_n22938 & new_n22867;
  assign new_n22940 = new_n22936 ^ new_n22920;
  assign new_n22941 = ~new_n22862 & ~new_n22940;
  assign new_n22942 = new_n22941 ^ new_n22939;
  assign new_n22943 = ~new_n22903 & ~new_n22940;
  assign new_n22944 = new_n22943 ^ new_n22942;
  assign new_n22945 = new_n22886 ^ new_n22841;
  assign new_n22946 = new_n22908 ^ new_n22847;
  assign new_n22947 = new_n22946 ^ new_n22924;
  assign new_n22948 = new_n22947 ^ new_n22932;
  assign new_n22949 = new_n22948 ^ new_n22945;
  assign new_n22950 = new_n22928 ^ new_n22901;
  assign new_n22951 = ~new_n22949 & new_n22950;
  assign new_n22952 = new_n22951 ^ new_n22909;
  assign new_n22953 = new_n22952 ^ new_n22892;
  assign new_n22954 = new_n22950 ^ new_n22936;
  assign new_n22955 = ~new_n22953 & new_n22954;
  assign new_n22956 = new_n22955 ^ new_n22949;
  assign new_n22957 = ~new_n22894 & ~new_n22956;
  assign new_n22958 = ~new_n22938 & new_n22923;
  assign new_n22959 = new_n22886 ^ new_n22854;
  assign new_n22960 = new_n22924 ^ new_n22911;
  assign new_n22961 = new_n22955 ^ new_n22936;
  assign new_n22962 = new_n22961 ^ new_n22960;
  assign new_n22963 = new_n22962 ^ new_n22959;
  assign new_n22964 = new_n22963 ^ new_n22847;
  assign new_n22965 = new_n22951 ^ new_n22898;
  assign new_n22966 = new_n22965 ^ new_n22905;
  assign new_n22967 = new_n22966 ^ new_n22964;
  assign new_n22968 = ~new_n22967 & new_n22902;
  assign new_n22969 = new_n22951 ^ new_n22934;
  assign new_n22970 = new_n22909 ^ new_n22900;
  assign new_n22971 = new_n22970 ^ new_n22969;
  assign new_n22972 = ~new_n22971 & new_n22848;
  assign new_n22973 = new_n22972 ^ new_n22968;
  assign new_n22974 = new_n22973 ^ new_n22958;
  assign new_n22975 = new_n22974 ^ new_n22957;
  assign new_n22976 = new_n22955 ^ new_n22951;
  assign new_n22977 = new_n22976 ^ new_n22927;
  assign new_n22978 = new_n22891 & new_n22977;
  assign new_n22979 = new_n22978 ^ new_n22975;
  assign new_n22980 = new_n22979 ^ new_n22944;
  assign new_n22981 = new_n21327 ^ new_n21303;
  assign new_n22982 = new_n22981 ^ new_n18557;
  assign new_n22983 = new_n18588 ^ new_n16382;
  assign new_n22984 = new_n22983 ^ new_n18751;
  assign new_n22985 = new_n22984 ^ new_n22982;
  assign new_n22986 = new_n18773 ^ new_n18720;
  assign new_n22987 = new_n22986 ^ new_n18804;
  assign new_n22988 = new_n22090 ^ new_n21332;
  assign new_n22989 = new_n22988 ^ new_n18721;
  assign new_n22990 = new_n22989 ^ new_n16383;
  assign new_n22991 = new_n22990 ^ new_n22987;
  assign new_n22992 = new_n22991 ^ new_n22985;
  assign new_n22993 = new_n22123 ^ new_n21315;
  assign new_n22994 = new_n22993 ^ new_n18786;
  assign new_n22995 = new_n22994 ^ new_n16383;
  assign new_n22996 = new_n18803 ^ new_n18781;
  assign new_n22997 = new_n22996 ^ new_n18701;
  assign new_n22998 = new_n22997 ^ new_n22995;
  assign new_n22999 = new_n18619 ^ new_n16383;
  assign new_n23000 = new_n21955 ^ new_n21311;
  assign new_n23001 = new_n23000 ^ new_n18710;
  assign new_n23002 = new_n18829 ^ new_n18826;
  assign new_n23003 = new_n23002 ^ new_n23001;
  assign new_n23004 = new_n23003 ^ new_n22999;
  assign new_n23005 = new_n23004 ^ new_n22998;
  assign new_n23006 = new_n23005 ^ new_n22992;
  assign new_n23007 = new_n22147 ^ new_n21345;
  assign new_n23008 = new_n23007 ^ new_n18582;
  assign new_n23009 = new_n18830 ^ new_n16383;
  assign new_n23010 = new_n23009 ^ new_n23008;
  assign new_n23011 = new_n23010 ^ new_n23006;
  assign new_n23012 = new_n22016 ^ new_n21306;
  assign new_n23013 = new_n23012 ^ new_n18677;
  assign new_n23014 = new_n23013 ^ new_n18604;
  assign new_n23015 = new_n18808 ^ new_n18689;
  assign new_n23016 = new_n23015 ^ new_n18656;
  assign new_n23017 = new_n23016 ^ new_n23014;
  assign new_n23018 = new_n23017 ^ new_n23005;
  assign new_n23019 = new_n22056 ^ new_n21322;
  assign new_n23020 = new_n23019 ^ new_n18565;
  assign new_n23021 = new_n18750 ^ new_n17414;
  assign new_n23022 = new_n23021 ^ new_n18732;
  assign new_n23023 = new_n23022 ^ new_n23020;
  assign new_n23024 = new_n23023 ^ new_n23018;
  assign new_n23025 = new_n22992 & new_n23024;
  assign new_n23026 = new_n23017 ^ new_n22985;
  assign new_n23027 = new_n22079 ^ new_n21350;
  assign new_n23028 = new_n23027 ^ new_n18736;
  assign new_n23029 = new_n18758 ^ new_n18727;
  assign new_n23030 = new_n23029 ^ new_n18775;
  assign new_n23031 = new_n23030 ^ new_n23028;
  assign new_n23032 = new_n23031 ^ new_n23023;
  assign new_n23033 = new_n23032 ^ new_n23006;
  assign new_n23034 = ~new_n23033 & new_n23026;
  assign new_n23035 = new_n23034 ^ new_n23025;
  assign new_n23036 = new_n23031 ^ new_n23018;
  assign new_n23037 = new_n23036 ^ new_n23035;
  assign new_n23038 = new_n23024 ^ new_n23010;
  assign new_n23039 = new_n23032 ^ new_n23010;
  assign new_n23040 = new_n23039 ^ new_n22985;
  assign new_n23041 = ~new_n23038 & ~new_n23040;
  assign new_n23042 = new_n23004 ^ new_n22985;
  assign new_n23043 = ~new_n23042 & new_n23036;
  assign new_n23044 = new_n23043 ^ new_n23041;
  assign new_n23045 = new_n23044 ^ new_n22985;
  assign new_n23046 = new_n23045 ^ new_n23037;
  assign new_n23047 = new_n23004 ^ new_n22991;
  assign new_n23048 = new_n23047 ^ new_n23026;
  assign new_n23049 = ~new_n23006 & ~new_n23048;
  assign new_n23050 = new_n23049 ^ new_n23023;
  assign new_n23051 = ~new_n23010 & ~new_n23032;
  assign new_n23052 = new_n22991 & new_n23010;
  assign new_n23053 = new_n23052 ^ new_n23051;
  assign new_n23054 = new_n23053 ^ new_n23050;
  assign new_n23055 = new_n23004 & new_n23039;
  assign new_n23056 = new_n23055 ^ new_n23004;
  assign new_n23057 = new_n23056 ^ new_n23043;
  assign new_n23058 = new_n23057 ^ new_n23026;
  assign new_n23059 = new_n23031 ^ new_n22991;
  assign new_n23060 = new_n23059 ^ new_n23026;
  assign new_n23061 = new_n23017 ^ new_n22991;
  assign new_n23062 = ~new_n23060 & new_n23061;
  assign new_n23063 = new_n23062 ^ new_n23025;
  assign new_n23064 = new_n23031 ^ new_n22998;
  assign new_n23065 = new_n23064 ^ new_n23063;
  assign new_n23066 = new_n23065 ^ new_n23058;
  assign new_n23067 = new_n23050 ^ new_n23006;
  assign new_n23068 = new_n23039 ^ new_n23004;
  assign new_n23069 = new_n23068 ^ new_n23026;
  assign new_n23070 = new_n23011 & new_n23069;
  assign new_n23071 = new_n23070 ^ new_n23025;
  assign new_n23072 = new_n23062 ^ new_n23017;
  assign new_n23073 = new_n23072 ^ new_n23071;
  assign new_n23074 = new_n23073 ^ new_n23067;
  assign new_n23075 = ~new_n23066 & new_n23074;
  assign new_n23076 = new_n23075 ^ new_n23054;
  assign new_n23077 = new_n23076 ^ new_n23037;
  assign new_n23078 = new_n23055 ^ new_n23041;
  assign new_n23079 = new_n23062 ^ new_n23034;
  assign new_n23080 = new_n23079 ^ new_n23078;
  assign new_n23081 = ~new_n23077 & ~new_n23080;
  assign new_n23082 = new_n23081 ^ new_n23075;
  assign new_n23083 = new_n23046 & new_n23082;
  assign new_n23084 = new_n23083 ^ new_n23081;
  assign new_n23085 = new_n23084 ^ new_n23080;
  assign new_n23086 = ~new_n23085 & new_n23011;
  assign new_n23087 = new_n23083 ^ new_n23066;
  assign new_n23088 = ~new_n23006 & ~new_n23087;
  assign new_n23089 = new_n23088 ^ new_n23086;
  assign new_n23090 = ~new_n23048 & ~new_n23087;
  assign new_n23091 = new_n23090 ^ new_n23089;
  assign new_n23092 = new_n23031 ^ new_n22985;
  assign new_n23093 = new_n23053 ^ new_n22991;
  assign new_n23094 = new_n23093 ^ new_n23070;
  assign new_n23095 = new_n23094 ^ new_n23079;
  assign new_n23096 = new_n23095 ^ new_n23092;
  assign new_n23097 = new_n23075 ^ new_n23046;
  assign new_n23098 = ~new_n23096 & new_n23097;
  assign new_n23099 = new_n23098 ^ new_n23054;
  assign new_n23100 = new_n23099 ^ new_n23037;
  assign new_n23101 = new_n23097 ^ new_n23083;
  assign new_n23102 = ~new_n23100 & new_n23101;
  assign new_n23103 = new_n23102 ^ new_n23096;
  assign new_n23104 = ~new_n23039 & ~new_n23103;
  assign new_n23105 = ~new_n23085 & new_n23069;
  assign new_n23106 = new_n23031 ^ new_n23004;
  assign new_n23107 = new_n23070 ^ new_n23056;
  assign new_n23108 = new_n23102 ^ new_n23083;
  assign new_n23109 = new_n23108 ^ new_n23107;
  assign new_n23110 = new_n23109 ^ new_n23106;
  assign new_n23111 = new_n23110 ^ new_n22991;
  assign new_n23112 = new_n23098 ^ new_n23043;
  assign new_n23113 = new_n23112 ^ new_n23050;
  assign new_n23114 = new_n23113 ^ new_n23111;
  assign new_n23115 = ~new_n23114 & new_n23061;
  assign new_n23116 = new_n23098 ^ new_n23081;
  assign new_n23117 = new_n23054 ^ new_n23045;
  assign new_n23118 = new_n23117 ^ new_n23116;
  assign new_n23119 = ~new_n23118 & new_n22992;
  assign new_n23120 = new_n23119 ^ new_n23115;
  assign new_n23121 = new_n23120 ^ new_n23105;
  assign new_n23122 = new_n23121 ^ new_n23104;
  assign new_n23123 = new_n23102 ^ new_n23098;
  assign new_n23124 = new_n23123 ^ new_n23074;
  assign new_n23125 = new_n23036 & new_n23124;
  assign new_n23126 = new_n23125 ^ new_n23122;
  assign new_n23127 = new_n23126 ^ new_n23091;
  assign new_n23128 = new_n23127 ^ new_n22980;
  assign new_n23129 = new_n19891 ^ new_n19839;
  assign new_n23130 = new_n23129 ^ new_n19882;
  assign new_n23131 = new_n20798 ^ new_n11504;
  assign new_n23132 = new_n19754 ^ new_n19740;
  assign new_n23133 = new_n23132 ^ new_n23131;
  assign new_n23134 = new_n23133 ^ new_n19771;
  assign new_n23135 = new_n23134 ^ new_n23130;
  assign new_n23136 = new_n23132 ^ new_n19867;
  assign new_n23137 = new_n23136 ^ new_n19888;
  assign new_n23138 = new_n20856 ^ new_n11537;
  assign new_n23139 = new_n23138 ^ new_n19827;
  assign new_n23140 = new_n23139 ^ new_n19864;
  assign new_n23141 = new_n23140 ^ new_n23137;
  assign new_n23142 = new_n23141 ^ new_n23135;
  assign new_n23143 = new_n19849 ^ new_n19808;
  assign new_n23144 = new_n20430 ^ new_n11582;
  assign new_n23145 = new_n23144 ^ new_n19882;
  assign new_n23146 = new_n23145 ^ new_n19827;
  assign new_n23147 = new_n23146 ^ new_n23143;
  assign new_n23148 = new_n23147 ^ new_n23142;
  assign new_n23149 = new_n19746 ^ new_n19719;
  assign new_n23150 = new_n20898 ^ new_n11408;
  assign new_n23151 = new_n23150 ^ new_n19171;
  assign new_n23152 = new_n23151 ^ new_n19672;
  assign new_n23153 = new_n23152 ^ new_n23149;
  assign new_n23154 = new_n23153 ^ new_n23148;
  assign new_n23155 = new_n19782 ^ new_n19612;
  assign new_n23156 = new_n20957 ^ new_n11560;
  assign new_n23157 = new_n23156 ^ new_n19740;
  assign new_n23158 = new_n23157 ^ new_n19171;
  assign new_n23159 = new_n23158 ^ new_n23155;
  assign new_n23160 = new_n20971 ^ new_n11465;
  assign new_n23161 = new_n23160 ^ new_n19700;
  assign new_n23162 = new_n23161 ^ new_n23132;
  assign new_n23163 = new_n19853 ^ new_n19777;
  assign new_n23164 = new_n23163 ^ new_n19839;
  assign new_n23165 = new_n23164 ^ new_n23162;
  assign new_n23166 = new_n23165 ^ new_n23159;
  assign new_n23167 = new_n23166 ^ new_n23142;
  assign new_n23168 = new_n23159 ^ new_n23141;
  assign new_n23169 = new_n23165 ^ new_n23147;
  assign new_n23170 = new_n23169 ^ new_n23168;
  assign new_n23171 = new_n23167 & new_n23170;
  assign new_n23172 = new_n23171 ^ new_n23153;
  assign new_n23173 = new_n20936 ^ new_n11425;
  assign new_n23174 = new_n23173 ^ new_n19864;
  assign new_n23175 = new_n23132 ^ new_n19796;
  assign new_n23176 = new_n23175 ^ new_n23174;
  assign new_n23177 = new_n19672 ^ new_n19464;
  assign new_n23178 = new_n20927 ^ new_n10300;
  assign new_n23179 = new_n19777 ^ new_n19772;
  assign new_n23180 = new_n23179 ^ new_n23178;
  assign new_n23181 = new_n23180 ^ new_n23177;
  assign new_n23182 = new_n23181 ^ new_n23153;
  assign new_n23183 = ~new_n23182 & new_n23176;
  assign new_n23184 = ~new_n23176 & new_n23165;
  assign new_n23185 = new_n23184 ^ new_n23183;
  assign new_n23186 = new_n23185 ^ new_n23172;
  assign new_n23187 = new_n23182 ^ new_n23176;
  assign new_n23188 = ~new_n23141 & ~new_n23187;
  assign new_n23189 = new_n23188 ^ new_n23141;
  assign new_n23190 = new_n23181 ^ new_n23148;
  assign new_n23191 = new_n23168 & new_n23190;
  assign new_n23192 = new_n23191 ^ new_n23189;
  assign new_n23193 = new_n23159 ^ new_n23147;
  assign new_n23194 = new_n23193 ^ new_n23192;
  assign new_n23195 = new_n23154 & new_n23166;
  assign new_n23196 = new_n23181 ^ new_n23165;
  assign new_n23197 = new_n23196 ^ new_n23193;
  assign new_n23198 = new_n23169 & new_n23197;
  assign new_n23199 = new_n23198 ^ new_n23195;
  assign new_n23200 = new_n23181 ^ new_n23135;
  assign new_n23201 = new_n23200 ^ new_n23199;
  assign new_n23202 = new_n23201 ^ new_n23194;
  assign new_n23203 = new_n23172 ^ new_n23167;
  assign new_n23204 = new_n23187 ^ new_n23141;
  assign new_n23205 = new_n23204 ^ new_n23193;
  assign new_n23206 = new_n23176 ^ new_n23167;
  assign new_n23207 = new_n23205 & new_n23206;
  assign new_n23208 = new_n23207 ^ new_n23195;
  assign new_n23209 = new_n23198 ^ new_n23147;
  assign new_n23210 = new_n23209 ^ new_n23208;
  assign new_n23211 = new_n23210 ^ new_n23203;
  assign new_n23212 = ~new_n23202 & new_n23211;
  assign new_n23213 = new_n23212 ^ new_n23186;
  assign new_n23214 = new_n23182 ^ new_n23167;
  assign new_n23215 = new_n23193 & new_n23214;
  assign new_n23216 = new_n23215 ^ new_n23195;
  assign new_n23217 = new_n23216 ^ new_n23190;
  assign new_n23218 = new_n23217 ^ new_n23213;
  assign new_n23219 = new_n23187 ^ new_n23159;
  assign new_n23220 = new_n23176 ^ new_n23154;
  assign new_n23221 = new_n23219 & new_n23220;
  assign new_n23222 = new_n23221 ^ new_n23188;
  assign new_n23223 = new_n23215 ^ new_n23198;
  assign new_n23224 = new_n23223 ^ new_n23222;
  assign new_n23225 = ~new_n23224 & new_n23218;
  assign new_n23226 = new_n23181 ^ new_n23159;
  assign new_n23227 = new_n23185 ^ new_n23165;
  assign new_n23228 = new_n23227 ^ new_n23207;
  assign new_n23229 = new_n23228 ^ new_n23223;
  assign new_n23230 = new_n23229 ^ new_n23226;
  assign new_n23231 = new_n23221 ^ new_n23191;
  assign new_n23232 = new_n23231 ^ new_n23159;
  assign new_n23233 = new_n23232 ^ new_n23217;
  assign new_n23234 = new_n23233 ^ new_n23212;
  assign new_n23235 = new_n23230 & new_n23234;
  assign new_n23236 = new_n23235 ^ new_n23225;
  assign new_n23237 = new_n23232 ^ new_n23186;
  assign new_n23238 = new_n23237 ^ new_n23236;
  assign new_n23239 = new_n23154 & new_n23238;
  assign new_n23240 = new_n23166 & new_n23238;
  assign new_n23241 = new_n23240 ^ new_n23239;
  assign new_n23242 = new_n23225 ^ new_n23159;
  assign new_n23243 = new_n23227 ^ new_n23221;
  assign new_n23244 = new_n23181 ^ new_n23141;
  assign new_n23245 = new_n23207 ^ new_n23189;
  assign new_n23246 = new_n23235 ^ new_n23186;
  assign new_n23247 = new_n23246 ^ new_n23217;
  assign new_n23248 = new_n23225 ^ new_n23212;
  assign new_n23249 = new_n23233 & new_n23248;
  assign new_n23250 = new_n23249 ^ new_n23234;
  assign new_n23251 = new_n23247 & new_n23250;
  assign new_n23252 = new_n23251 ^ new_n23249;
  assign new_n23253 = new_n23252 ^ new_n23245;
  assign new_n23254 = new_n23253 ^ new_n23244;
  assign new_n23255 = new_n23254 ^ new_n23243;
  assign new_n23256 = new_n23255 ^ new_n23242;
  assign new_n23257 = ~new_n23256 & new_n23193;
  assign new_n23258 = new_n23219 & new_n23247;
  assign new_n23259 = ~new_n23256 & new_n23214;
  assign new_n23260 = new_n23259 ^ new_n23258;
  assign new_n23261 = new_n23249 ^ new_n23202;
  assign new_n23262 = ~new_n23261 & new_n23167;
  assign new_n23263 = new_n23233 ^ new_n23225;
  assign new_n23264 = new_n23176 & new_n23263;
  assign new_n23265 = new_n23264 ^ new_n23262;
  assign new_n23266 = new_n23251 ^ new_n23235;
  assign new_n23267 = new_n23266 ^ new_n23211;
  assign new_n23268 = new_n23168 & new_n23267;
  assign new_n23269 = new_n23268 ^ new_n23265;
  assign new_n23270 = new_n23269 ^ new_n23260;
  assign new_n23271 = new_n23270 ^ new_n23257;
  assign new_n23272 = new_n23271 ^ new_n23241;
  assign new_n23273 = ~new_n23118 & new_n23024;
  assign new_n23274 = new_n23273 ^ new_n23119;
  assign new_n23275 = new_n23081 ^ new_n22985;
  assign new_n23276 = new_n23093 ^ new_n23041;
  assign new_n23277 = new_n23276 ^ new_n23110;
  assign new_n23278 = new_n23277 ^ new_n23275;
  assign new_n23279 = new_n23026 & new_n23278;
  assign new_n23280 = ~new_n23040 & ~new_n23100;
  assign new_n23281 = ~new_n23033 & new_n23278;
  assign new_n23282 = new_n23281 ^ new_n23280;
  assign new_n23283 = new_n23081 ^ new_n23046;
  assign new_n23284 = ~new_n23010 & new_n23283;
  assign new_n23285 = new_n23284 ^ new_n23088;
  assign new_n23286 = ~new_n23042 & new_n23124;
  assign new_n23287 = new_n23286 ^ new_n23285;
  assign new_n23288 = new_n23287 ^ new_n23282;
  assign new_n23289 = new_n23288 ^ new_n23279;
  assign new_n23290 = new_n23289 ^ new_n23274;
  assign new_n23291 = new_n23290 ^ new_n23272;
  assign new_n23292 = new_n23291 ^ new_n23128;
  assign new_n23293 = new_n23292 ^ new_n22836;
  assign new_n23294 = new_n22665 ^ new_n22586;
  assign new_n23295 = new_n22645 ^ new_n22603;
  assign new_n23296 = new_n23295 ^ new_n22597;
  assign new_n23297 = new_n23296 ^ new_n23294;
  assign new_n23298 = ~new_n23297 & new_n22608;
  assign new_n23299 = new_n23298 ^ new_n22649;
  assign new_n23300 = new_n22660 ^ new_n22636;
  assign new_n23301 = new_n23300 ^ new_n22635;
  assign new_n23302 = ~new_n23301 & new_n22618;
  assign new_n23303 = new_n23302 ^ new_n22671;
  assign new_n23304 = ~new_n22670 & new_n22595;
  assign new_n23305 = new_n23304 ^ new_n23303;
  assign new_n23306 = ~new_n23301 & new_n22617;
  assign new_n23307 = ~new_n23297 & new_n22609;
  assign new_n23308 = new_n23307 ^ new_n22650;
  assign new_n23309 = new_n23308 ^ new_n23306;
  assign new_n23310 = new_n23309 ^ new_n23305;
  assign new_n23311 = new_n23310 ^ new_n23299;
  assign new_n23312 = new_n23311 ^ new_n19029;
  assign new_n23313 = new_n23312 ^ new_n7863;
  assign new_n23314 = new_n22817 ^ new_n22726;
  assign new_n23315 = new_n22798 ^ new_n22756;
  assign new_n23316 = new_n23315 ^ new_n22750;
  assign new_n23317 = new_n23316 ^ new_n23314;
  assign new_n23318 = ~new_n22761 & ~new_n23317;
  assign new_n23319 = new_n23318 ^ new_n22802;
  assign new_n23320 = new_n22812 ^ new_n22789;
  assign new_n23321 = new_n23320 ^ new_n22788;
  assign new_n23322 = ~new_n22769 & ~new_n23321;
  assign new_n23323 = new_n23322 ^ new_n22825;
  assign new_n23324 = ~new_n22748 & ~new_n22824;
  assign new_n23325 = new_n23324 ^ new_n23323;
  assign new_n23326 = ~new_n22771 & ~new_n23321;
  assign new_n23327 = ~new_n22762 & ~new_n23317;
  assign new_n23328 = new_n23327 ^ new_n22803;
  assign new_n23329 = new_n23328 ^ new_n23326;
  assign new_n23330 = new_n23329 ^ new_n23325;
  assign new_n23331 = new_n23330 ^ new_n23319;
  assign new_n23332 = new_n23331 ^ new_n23313;
  assign new_n23333 = ~new_n22971 & new_n22879;
  assign new_n23334 = new_n23333 ^ new_n22972;
  assign new_n23335 = new_n22934 ^ new_n22841;
  assign new_n23336 = new_n22946 ^ new_n22896;
  assign new_n23337 = new_n23336 ^ new_n22963;
  assign new_n23338 = new_n23337 ^ new_n23335;
  assign new_n23339 = new_n22881 & new_n23338;
  assign new_n23340 = ~new_n22888 & new_n23338;
  assign new_n23341 = ~new_n22895 & ~new_n22953;
  assign new_n23342 = new_n23341 ^ new_n23340;
  assign new_n23343 = ~new_n22897 & new_n22977;
  assign new_n23344 = new_n22934 ^ new_n22901;
  assign new_n23345 = ~new_n22866 & new_n23344;
  assign new_n23346 = new_n23345 ^ new_n22941;
  assign new_n23347 = new_n23346 ^ new_n23343;
  assign new_n23348 = new_n23347 ^ new_n23342;
  assign new_n23349 = new_n23348 ^ new_n23339;
  assign new_n23350 = new_n23349 ^ new_n23334;
  assign new_n23351 = new_n23350 ^ new_n23290;
  assign new_n23352 = new_n23254 ^ new_n23165;
  assign new_n23353 = new_n23235 ^ new_n23191;
  assign new_n23354 = new_n23353 ^ new_n23172;
  assign new_n23355 = new_n23354 ^ new_n23352;
  assign new_n23356 = ~new_n23355 & new_n23197;
  assign new_n23357 = new_n23356 ^ new_n23239;
  assign new_n23358 = new_n23249 ^ new_n23225;
  assign new_n23359 = new_n23358 ^ new_n23224;
  assign new_n23360 = ~new_n23359 & new_n23206;
  assign new_n23361 = new_n23360 ^ new_n23262;
  assign new_n23362 = ~new_n23261 & new_n23170;
  assign new_n23363 = new_n23362 ^ new_n23361;
  assign new_n23364 = ~new_n23359 & new_n23205;
  assign new_n23365 = ~new_n23355 & new_n23169;
  assign new_n23366 = new_n23365 ^ new_n23240;
  assign new_n23367 = new_n23366 ^ new_n23364;
  assign new_n23368 = new_n23367 ^ new_n23363;
  assign new_n23369 = new_n23368 ^ new_n23357;
  assign new_n23370 = ~new_n23060 & ~new_n23114;
  assign new_n23371 = new_n23370 ^ new_n23273;
  assign new_n23372 = new_n23121 ^ new_n23091;
  assign new_n23373 = new_n23372 ^ new_n23371;
  assign new_n23374 = new_n23373 ^ new_n23369;
  assign new_n23375 = new_n23374 ^ new_n23351;
  assign new_n23376 = new_n23375 ^ new_n23332;
  assign new_n23377 = new_n23376 ^ new_n23293;
  assign new_n23378 = new_n22601 & new_n22676;
  assign new_n23379 = new_n23378 ^ new_n22678;
  assign new_n23380 = new_n22662 ^ new_n22640;
  assign new_n23381 = new_n22616 & new_n23380;
  assign new_n23382 = new_n22631 & new_n22653;
  assign new_n23383 = new_n23382 ^ new_n23381;
  assign new_n23384 = new_n23383 ^ new_n23308;
  assign new_n23385 = new_n23384 ^ new_n23379;
  assign new_n23386 = new_n23385 ^ new_n19861;
  assign new_n23387 = new_n23386 ^ new_n7898;
  assign new_n23388 = new_n22755 & new_n22830;
  assign new_n23389 = new_n23388 ^ new_n22832;
  assign new_n23390 = new_n22814 ^ new_n22793;
  assign new_n23391 = ~new_n22770 & new_n23390;
  assign new_n23392 = ~new_n22784 & new_n22810;
  assign new_n23393 = new_n23392 ^ new_n23391;
  assign new_n23394 = new_n23393 ^ new_n23328;
  assign new_n23395 = new_n23394 ^ new_n23389;
  assign new_n23396 = new_n23395 ^ new_n23387;
  assign new_n23397 = new_n23190 & new_n23267;
  assign new_n23398 = new_n23397 ^ new_n23269;
  assign new_n23399 = new_n23251 ^ new_n23230;
  assign new_n23400 = new_n23204 & new_n23399;
  assign new_n23401 = new_n23220 & new_n23247;
  assign new_n23402 = new_n23401 ^ new_n23400;
  assign new_n23403 = new_n23402 ^ new_n23366;
  assign new_n23404 = new_n23403 ^ new_n23398;
  assign new_n23405 = new_n23287 ^ new_n23125;
  assign new_n23406 = ~new_n23038 & ~new_n23100;
  assign new_n23407 = ~new_n23103 & new_n23068;
  assign new_n23408 = new_n23407 ^ new_n23406;
  assign new_n23409 = new_n23408 ^ new_n23120;
  assign new_n23410 = new_n23409 ^ new_n23405;
  assign new_n23411 = new_n23410 ^ new_n23404;
  assign new_n23412 = new_n23273 ^ new_n23090;
  assign new_n23413 = new_n23370 ^ new_n23126;
  assign new_n23414 = new_n23413 ^ new_n23412;
  assign new_n23415 = new_n23333 ^ new_n22943;
  assign new_n23416 = ~new_n22915 & ~new_n22967;
  assign new_n23417 = new_n23416 ^ new_n22979;
  assign new_n23418 = new_n23417 ^ new_n23415;
  assign new_n23419 = new_n23418 ^ new_n23414;
  assign new_n23420 = new_n23419 ^ new_n23411;
  assign new_n23421 = new_n23420 ^ new_n23396;
  assign new_n23422 = new_n23421 ^ new_n23377;
  assign new_n23423 = ~new_n22893 & ~new_n22953;
  assign new_n23424 = new_n23423 ^ new_n22943;
  assign new_n23425 = new_n23345 ^ new_n22939;
  assign new_n23426 = new_n23425 ^ new_n22975;
  assign new_n23427 = new_n23426 ^ new_n23424;
  assign new_n23428 = new_n23406 ^ new_n23090;
  assign new_n23429 = new_n23284 ^ new_n23086;
  assign new_n23430 = new_n23429 ^ new_n23122;
  assign new_n23431 = new_n23430 ^ new_n23428;
  assign new_n23432 = new_n23431 ^ new_n23427;
  assign new_n23433 = new_n23187 & new_n23399;
  assign new_n23434 = new_n23433 ^ new_n23367;
  assign new_n23435 = new_n23434 ^ new_n23397;
  assign new_n23436 = new_n23435 ^ new_n23363;
  assign new_n23437 = new_n23436 ^ new_n23127;
  assign new_n23438 = new_n23437 ^ new_n23432;
  assign new_n23439 = new_n22585 & new_n23380;
  assign new_n23440 = new_n23439 ^ new_n23309;
  assign new_n23441 = new_n23440 ^ new_n23378;
  assign new_n23442 = new_n23441 ^ new_n23305;
  assign new_n23443 = new_n23442 ^ new_n19775;
  assign new_n23444 = new_n23443 ^ new_n7967;
  assign new_n23445 = ~new_n22734 & new_n23390;
  assign new_n23446 = new_n23445 ^ new_n23329;
  assign new_n23447 = new_n23446 ^ new_n23388;
  assign new_n23448 = new_n23447 ^ new_n23325;
  assign new_n23449 = new_n23448 ^ new_n23444;
  assign new_n23450 = new_n23449 ^ new_n23419;
  assign new_n23451 = new_n23450 ^ new_n23438;
  assign new_n23452 = new_n23451 ^ new_n23422;
  assign new_n23453 = ~new_n23421 & ~new_n23452;
  assign new_n23454 = new_n23453 ^ new_n23451;
  assign new_n23455 = new_n23304 ^ new_n22649;
  assign new_n23456 = new_n23441 ^ new_n23298;
  assign new_n23457 = new_n23456 ^ new_n23455;
  assign new_n23458 = new_n23457 ^ new_n19731;
  assign new_n23459 = new_n23458 ^ new_n7939;
  assign new_n23460 = new_n23324 ^ new_n22802;
  assign new_n23461 = new_n23447 ^ new_n23318;
  assign new_n23462 = new_n23461 ^ new_n23460;
  assign new_n23463 = new_n23462 ^ new_n23459;
  assign new_n23464 = new_n23416 ^ new_n23333;
  assign new_n23465 = new_n22974 ^ new_n22944;
  assign new_n23466 = new_n23465 ^ new_n23464;
  assign new_n23467 = new_n23466 ^ new_n23373;
  assign new_n23468 = new_n23362 ^ new_n23239;
  assign new_n23469 = new_n23435 ^ new_n23356;
  assign new_n23470 = new_n23469 ^ new_n23468;
  assign new_n23471 = new_n23470 ^ new_n23414;
  assign new_n23472 = new_n23471 ^ new_n23467;
  assign new_n23473 = new_n23472 ^ new_n23463;
  assign new_n23474 = new_n23473 ^ new_n23451;
  assign new_n23475 = new_n23382 ^ new_n23304;
  assign new_n23476 = new_n23302 ^ new_n22673;
  assign new_n23477 = new_n23476 ^ new_n23440;
  assign new_n23478 = new_n23477 ^ new_n23475;
  assign new_n23479 = new_n23478 ^ new_n19834;
  assign new_n23480 = new_n23479 ^ new_n7824;
  assign new_n23481 = new_n23392 ^ new_n23324;
  assign new_n23482 = new_n23322 ^ new_n22827;
  assign new_n23483 = new_n23482 ^ new_n23446;
  assign new_n23484 = new_n23483 ^ new_n23481;
  assign new_n23485 = new_n23484 ^ new_n23480;
  assign new_n23486 = new_n23485 ^ new_n23419;
  assign new_n23487 = new_n22894 ^ new_n22847;
  assign new_n23488 = ~new_n23487 & new_n23344;
  assign new_n23489 = new_n23488 ^ new_n23417;
  assign new_n23490 = new_n23489 ^ new_n23348;
  assign new_n23491 = new_n23039 ^ new_n22991;
  assign new_n23492 = ~new_n23491 & new_n23283;
  assign new_n23493 = new_n23492 ^ new_n23413;
  assign new_n23494 = new_n23493 ^ new_n23288;
  assign new_n23495 = new_n23494 ^ new_n23490;
  assign new_n23496 = new_n23401 ^ new_n23362;
  assign new_n23497 = new_n23360 ^ new_n23264;
  assign new_n23498 = new_n23497 ^ new_n23434;
  assign new_n23499 = new_n23498 ^ new_n23496;
  assign new_n23500 = new_n23499 ^ new_n23431;
  assign new_n23501 = new_n23500 ^ new_n23495;
  assign new_n23502 = new_n23501 ^ new_n23486;
  assign new_n23503 = ~new_n22956 & new_n22922;
  assign new_n23504 = new_n23503 ^ new_n23423;
  assign new_n23505 = new_n23504 ^ new_n22973;
  assign new_n23506 = new_n23347 ^ new_n22978;
  assign new_n23507 = new_n23506 ^ new_n23505;
  assign new_n23508 = new_n23507 ^ new_n23410;
  assign new_n23509 = new_n23286 ^ new_n23281;
  assign new_n23510 = new_n23370 ^ new_n23104;
  assign new_n23511 = new_n23510 ^ new_n23409;
  assign new_n23512 = new_n23511 ^ new_n23509;
  assign new_n23513 = new_n23268 ^ new_n23259;
  assign new_n23514 = new_n23433 ^ new_n23356;
  assign new_n23515 = new_n23514 ^ new_n23403;
  assign new_n23516 = new_n23515 ^ new_n23513;
  assign new_n23517 = new_n23516 ^ new_n23512;
  assign new_n23518 = new_n23517 ^ new_n23508;
  assign new_n23519 = new_n22677 ^ new_n22668;
  assign new_n23520 = new_n23439 ^ new_n23298;
  assign new_n23521 = new_n23520 ^ new_n23384;
  assign new_n23522 = new_n23521 ^ new_n23519;
  assign new_n23523 = new_n23522 ^ new_n19818;
  assign new_n23524 = new_n23523 ^ new_n7789;
  assign new_n23525 = new_n22831 ^ new_n22822;
  assign new_n23526 = new_n23445 ^ new_n23318;
  assign new_n23527 = new_n23526 ^ new_n23394;
  assign new_n23528 = new_n23527 ^ new_n23525;
  assign new_n23529 = new_n23528 ^ new_n23524;
  assign new_n23530 = new_n23529 ^ new_n23419;
  assign new_n23531 = new_n23530 ^ new_n23518;
  assign new_n23532 = new_n23531 ^ new_n23502;
  assign new_n23533 = new_n23532 ^ new_n23474;
  assign new_n23534 = new_n23531 ^ new_n23451;
  assign new_n23535 = new_n22587 & new_n22672;
  assign new_n23536 = new_n23535 ^ new_n23456;
  assign new_n23537 = new_n23536 ^ new_n22679;
  assign new_n23538 = new_n23537 ^ new_n19878;
  assign new_n23539 = new_n23538 ^ new_n1013;
  assign new_n23540 = new_n22735 & new_n22826;
  assign new_n23541 = new_n23540 ^ new_n23461;
  assign new_n23542 = new_n23541 ^ new_n22833;
  assign new_n23543 = new_n23542 ^ new_n23539;
  assign new_n23544 = new_n23343 ^ new_n23340;
  assign new_n23545 = new_n23416 ^ new_n22957;
  assign new_n23546 = new_n23545 ^ new_n23505;
  assign new_n23547 = new_n23546 ^ new_n23544;
  assign new_n23548 = new_n23547 ^ new_n23512;
  assign new_n23549 = new_n23187 ^ new_n23165;
  assign new_n23550 = new_n23263 & new_n23549;
  assign new_n23551 = new_n23550 ^ new_n23469;
  assign new_n23552 = new_n23551 ^ new_n23270;
  assign new_n23553 = new_n23552 ^ new_n23494;
  assign new_n23554 = new_n23553 ^ new_n23548;
  assign new_n23555 = new_n23554 ^ new_n23543;
  assign new_n23556 = new_n23555 ^ new_n23473;
  assign new_n23557 = new_n23556 ^ new_n23534;
  assign new_n23558 = ~new_n23533 & ~new_n23557;
  assign new_n23559 = new_n23558 ^ new_n23376;
  assign new_n23560 = new_n23559 ^ new_n23454;
  assign new_n23561 = new_n23559 ^ new_n23533;
  assign new_n23562 = new_n23533 ^ new_n23421;
  assign new_n23563 = new_n23531 ^ new_n23422;
  assign new_n23564 = new_n23563 ^ new_n23556;
  assign new_n23565 = new_n23562 & new_n23564;
  assign new_n23566 = new_n23555 ^ new_n23532;
  assign new_n23567 = new_n23566 ^ new_n23376;
  assign new_n23568 = new_n23474 & new_n23567;
  assign new_n23569 = new_n23568 ^ new_n23565;
  assign new_n23570 = new_n23451 ^ new_n23293;
  assign new_n23571 = new_n23570 ^ new_n23556;
  assign new_n23572 = new_n23555 ^ new_n23451;
  assign new_n23573 = ~new_n23571 & new_n23572;
  assign new_n23574 = new_n23573 ^ new_n23555;
  assign new_n23575 = new_n23574 ^ new_n23569;
  assign new_n23576 = new_n23575 ^ new_n23561;
  assign new_n23577 = new_n23422 & new_n23531;
  assign new_n23578 = new_n23577 ^ new_n23531;
  assign new_n23579 = new_n23566 ^ new_n23293;
  assign new_n23580 = new_n23531 ^ new_n23473;
  assign new_n23581 = ~new_n23580 & new_n23579;
  assign new_n23582 = new_n23581 ^ new_n23578;
  assign new_n23583 = new_n23582 ^ new_n23556;
  assign new_n23584 = new_n23573 ^ new_n23568;
  assign new_n23585 = new_n23502 ^ new_n23293;
  assign new_n23586 = new_n23585 ^ new_n23584;
  assign new_n23587 = new_n23586 ^ new_n23583;
  assign new_n23588 = ~new_n23587 & new_n23576;
  assign new_n23589 = new_n23588 ^ new_n23560;
  assign new_n23590 = new_n23533 ^ new_n23377;
  assign new_n23591 = ~new_n23590 & new_n23556;
  assign new_n23592 = new_n23591 ^ new_n23568;
  assign new_n23593 = new_n23592 ^ new_n23579;
  assign new_n23594 = new_n23593 ^ new_n23589;
  assign new_n23595 = new_n23473 ^ new_n23422;
  assign new_n23596 = new_n23567 ^ new_n23421;
  assign new_n23597 = ~new_n23595 & ~new_n23596;
  assign new_n23598 = new_n23597 ^ new_n23577;
  assign new_n23599 = new_n23591 ^ new_n23573;
  assign new_n23600 = new_n23599 ^ new_n23598;
  assign new_n23601 = ~new_n23594 & ~new_n23600;
  assign new_n23602 = new_n23597 ^ new_n23581;
  assign new_n23603 = new_n23602 ^ new_n23473;
  assign new_n23604 = new_n23603 ^ new_n23593;
  assign new_n23605 = new_n23604 ^ new_n23601;
  assign new_n23606 = ~new_n23452 & new_n23605;
  assign new_n23607 = new_n23531 ^ new_n23293;
  assign new_n23608 = new_n23578 ^ new_n23565;
  assign new_n23609 = new_n23601 ^ new_n23588;
  assign new_n23610 = ~new_n23604 & ~new_n23609;
  assign new_n23611 = new_n23610 ^ new_n23601;
  assign new_n23612 = new_n23604 ^ new_n23588;
  assign new_n23613 = new_n23473 ^ new_n23293;
  assign new_n23614 = new_n23565 ^ new_n23453;
  assign new_n23615 = new_n23614 ^ new_n23599;
  assign new_n23616 = new_n23615 ^ new_n23613;
  assign new_n23617 = ~new_n23616 & new_n23612;
  assign new_n23618 = new_n23617 ^ new_n23560;
  assign new_n23619 = new_n23618 ^ new_n23593;
  assign new_n23620 = ~new_n23611 & ~new_n23619;
  assign new_n23621 = new_n23612 ^ new_n23611;
  assign new_n23622 = new_n23621 ^ new_n23620;
  assign new_n23623 = new_n23622 ^ new_n23608;
  assign new_n23624 = new_n23623 ^ new_n23607;
  assign new_n23625 = new_n23624 ^ new_n23451;
  assign new_n23626 = new_n23617 ^ new_n23581;
  assign new_n23627 = new_n23626 ^ new_n23559;
  assign new_n23628 = new_n23627 ^ new_n23625;
  assign new_n23629 = ~new_n23571 & new_n23628;
  assign new_n23630 = new_n23620 ^ new_n23617;
  assign new_n23631 = new_n23630 ^ new_n23576;
  assign new_n23632 = new_n23579 & new_n23631;
  assign new_n23633 = new_n23621 ^ new_n23601;
  assign new_n23634 = new_n23633 ^ new_n23600;
  assign new_n23635 = new_n23564 & new_n23634;
  assign new_n23636 = new_n23572 & new_n23628;
  assign new_n23637 = new_n23617 ^ new_n23601;
  assign new_n23638 = new_n23603 ^ new_n23560;
  assign new_n23639 = new_n23638 ^ new_n23637;
  assign new_n23640 = ~new_n23639 & new_n23474;
  assign new_n23641 = new_n23640 ^ new_n23636;
  assign new_n23642 = new_n23641 ^ new_n23635;
  assign new_n23643 = new_n23620 ^ new_n23616;
  assign new_n23644 = ~new_n23422 & ~new_n23643;
  assign new_n23645 = new_n23644 ^ new_n23642;
  assign new_n23646 = new_n23645 ^ new_n23632;
  assign new_n23647 = new_n23646 ^ new_n23629;
  assign new_n23648 = new_n23647 ^ new_n23606;
  assign new_n23649 = ~new_n23595 & ~new_n23619;
  assign new_n23650 = new_n23601 ^ new_n23473;
  assign new_n23651 = new_n23597 ^ new_n23453;
  assign new_n23652 = new_n23651 ^ new_n23624;
  assign new_n23653 = new_n23652 ^ new_n23650;
  assign new_n23654 = ~new_n23590 & ~new_n23653;
  assign new_n23655 = new_n23654 ^ new_n23649;
  assign new_n23656 = ~new_n23421 & new_n23605;
  assign new_n23657 = new_n23621 ^ new_n23587;
  assign new_n23658 = ~new_n23533 & new_n23657;
  assign new_n23659 = new_n23658 ^ new_n23656;
  assign new_n23660 = ~new_n23580 & new_n23631;
  assign new_n23661 = new_n23660 ^ new_n23659;
  assign new_n23662 = new_n23661 ^ new_n23655;
  assign new_n23663 = new_n23662 ^ new_n23648;
  assign new_n23664 = new_n19808 ^ new_n19758;
  assign new_n23665 = new_n23664 ^ new_n19868;
  assign new_n23666 = new_n21955 ^ new_n15800;
  assign new_n23667 = new_n23666 ^ new_n19887;
  assign new_n23668 = new_n23667 ^ new_n19827;
  assign new_n23669 = new_n23668 ^ new_n23665;
  assign new_n23670 = new_n19853 ^ new_n19765;
  assign new_n23671 = new_n23670 ^ new_n19839;
  assign new_n23672 = new_n22123 ^ new_n15792;
  assign new_n23673 = new_n23672 ^ new_n19758;
  assign new_n23674 = new_n23673 ^ new_n19892;
  assign new_n23675 = new_n23674 ^ new_n23671;
  assign new_n23676 = new_n23675 ^ new_n23669;
  assign new_n23677 = new_n21303 ^ new_n15783;
  assign new_n23678 = new_n23677 ^ new_n19631;
  assign new_n23679 = new_n23132 ^ new_n19781;
  assign new_n23680 = new_n23679 ^ new_n23678;
  assign new_n23681 = new_n22090 ^ new_n15755;
  assign new_n23682 = new_n23681 ^ new_n19758;
  assign new_n23683 = new_n23682 ^ new_n19854;
  assign new_n23684 = new_n23179 ^ new_n19693;
  assign new_n23685 = new_n23684 ^ new_n23683;
  assign new_n23686 = new_n23685 ^ new_n23680;
  assign new_n23687 = new_n23686 ^ new_n23676;
  assign new_n23688 = new_n19867 ^ new_n19758;
  assign new_n23689 = new_n22147 ^ new_n15777;
  assign new_n23690 = new_n23689 ^ new_n19790;
  assign new_n23691 = new_n23690 ^ new_n19864;
  assign new_n23692 = new_n23691 ^ new_n23688;
  assign new_n23693 = new_n23692 ^ new_n23687;
  assign new_n23694 = new_n19720 ^ new_n19612;
  assign new_n23695 = new_n22056 ^ new_n15771;
  assign new_n23696 = new_n23695 ^ new_n19745;
  assign new_n23697 = new_n23696 ^ new_n19171;
  assign new_n23698 = new_n23697 ^ new_n23694;
  assign new_n23699 = new_n19891 ^ new_n19848;
  assign new_n23700 = new_n23699 ^ new_n19882;
  assign new_n23701 = new_n22016 ^ new_n15808;
  assign new_n23702 = new_n23701 ^ new_n19809;
  assign new_n23703 = new_n23702 ^ new_n23700;
  assign new_n23704 = new_n23703 ^ new_n23676;
  assign new_n23705 = new_n23704 ^ new_n23698;
  assign new_n23706 = new_n23705 ^ new_n23692;
  assign new_n23707 = new_n19773 ^ new_n19719;
  assign new_n23708 = new_n22079 ^ new_n15765;
  assign new_n23709 = new_n23708 ^ new_n19325;
  assign new_n23710 = new_n23709 ^ new_n19672;
  assign new_n23711 = new_n23710 ^ new_n23707;
  assign new_n23712 = new_n23711 ^ new_n23698;
  assign new_n23713 = new_n23712 ^ new_n23692;
  assign new_n23714 = new_n23713 ^ new_n23680;
  assign new_n23715 = new_n23706 & new_n23714;
  assign new_n23716 = new_n23711 ^ new_n23704;
  assign new_n23717 = new_n23680 ^ new_n23669;
  assign new_n23718 = new_n23716 & new_n23717;
  assign new_n23719 = new_n23718 ^ new_n23715;
  assign new_n23720 = new_n23719 ^ new_n23680;
  assign new_n23721 = new_n23703 ^ new_n23680;
  assign new_n23722 = new_n23712 ^ new_n23687;
  assign new_n23723 = new_n23721 & new_n23722;
  assign new_n23724 = new_n23686 & new_n23705;
  assign new_n23725 = new_n23724 ^ new_n23723;
  assign new_n23726 = new_n23725 ^ new_n23716;
  assign new_n23727 = new_n23726 ^ new_n23720;
  assign new_n23728 = new_n23713 ^ new_n23685;
  assign new_n23729 = new_n23692 & new_n23728;
  assign new_n23730 = new_n23729 ^ new_n23685;
  assign new_n23731 = new_n23703 ^ new_n23685;
  assign new_n23732 = new_n23731 ^ new_n23717;
  assign new_n23733 = new_n23687 & new_n23732;
  assign new_n23734 = new_n23733 ^ new_n23698;
  assign new_n23735 = new_n23734 ^ new_n23730;
  assign new_n23736 = ~new_n23669 & ~new_n23713;
  assign new_n23737 = new_n23736 ^ new_n23669;
  assign new_n23738 = new_n23737 ^ new_n23718;
  assign new_n23739 = new_n23738 ^ new_n23721;
  assign new_n23740 = new_n23711 ^ new_n23685;
  assign new_n23741 = new_n23740 ^ new_n23721;
  assign new_n23742 = new_n23731 & new_n23741;
  assign new_n23743 = new_n23742 ^ new_n23724;
  assign new_n23744 = new_n23711 ^ new_n23675;
  assign new_n23745 = new_n23744 ^ new_n23743;
  assign new_n23746 = new_n23745 ^ new_n23739;
  assign new_n23747 = new_n23734 ^ new_n23687;
  assign new_n23748 = new_n23713 ^ new_n23669;
  assign new_n23749 = new_n23748 ^ new_n23721;
  assign new_n23750 = new_n23693 & new_n23749;
  assign new_n23751 = new_n23750 ^ new_n23743;
  assign new_n23752 = new_n23751 ^ new_n23703;
  assign new_n23753 = new_n23752 ^ new_n23747;
  assign new_n23754 = ~new_n23746 & new_n23753;
  assign new_n23755 = new_n23754 ^ new_n23735;
  assign new_n23756 = new_n23755 ^ new_n23726;
  assign new_n23757 = new_n23742 ^ new_n23723;
  assign new_n23758 = new_n23736 ^ new_n23715;
  assign new_n23759 = new_n23758 ^ new_n23757;
  assign new_n23760 = ~new_n23759 & new_n23756;
  assign new_n23761 = new_n23760 ^ new_n23754;
  assign new_n23762 = ~new_n23727 & ~new_n23761;
  assign new_n23763 = new_n23762 ^ new_n23760;
  assign new_n23764 = new_n23754 ^ new_n23727;
  assign new_n23765 = new_n23764 ^ new_n23763;
  assign new_n23766 = new_n23765 ^ new_n23760;
  assign new_n23767 = new_n23766 ^ new_n23759;
  assign new_n23768 = new_n23693 & new_n23767;
  assign new_n23769 = new_n23765 ^ new_n23746;
  assign new_n23770 = new_n23687 & new_n23769;
  assign new_n23771 = new_n23770 ^ new_n23768;
  assign new_n23772 = new_n23732 & new_n23769;
  assign new_n23773 = new_n23772 ^ new_n23771;
  assign new_n23774 = new_n23711 ^ new_n23680;
  assign new_n23775 = new_n23750 ^ new_n23729;
  assign new_n23776 = new_n23775 ^ new_n23757;
  assign new_n23777 = new_n23776 ^ new_n23774;
  assign new_n23778 = new_n23764 & new_n23777;
  assign new_n23779 = new_n23778 ^ new_n23735;
  assign new_n23780 = new_n23779 ^ new_n23726;
  assign new_n23781 = ~new_n23763 & new_n23780;
  assign new_n23782 = new_n23781 ^ new_n23777;
  assign new_n23783 = new_n23713 & new_n23782;
  assign new_n23784 = new_n23749 & new_n23767;
  assign new_n23785 = new_n23711 ^ new_n23669;
  assign new_n23786 = new_n23750 ^ new_n23737;
  assign new_n23787 = new_n23781 ^ new_n23765;
  assign new_n23788 = new_n23787 ^ new_n23786;
  assign new_n23789 = new_n23788 ^ new_n23785;
  assign new_n23790 = new_n23789 ^ new_n23685;
  assign new_n23791 = new_n23778 ^ new_n23718;
  assign new_n23792 = new_n23791 ^ new_n23734;
  assign new_n23793 = new_n23792 ^ new_n23790;
  assign new_n23794 = new_n23731 & new_n23793;
  assign new_n23795 = new_n23778 ^ new_n23760;
  assign new_n23796 = new_n23735 ^ new_n23720;
  assign new_n23797 = new_n23796 ^ new_n23795;
  assign new_n23798 = new_n23686 & new_n23797;
  assign new_n23799 = new_n23798 ^ new_n23794;
  assign new_n23800 = new_n23799 ^ new_n23784;
  assign new_n23801 = new_n23800 ^ new_n23783;
  assign new_n23802 = new_n23781 ^ new_n23778;
  assign new_n23803 = new_n23802 ^ new_n23753;
  assign new_n23804 = new_n23716 & new_n23803;
  assign new_n23805 = new_n23804 ^ new_n23801;
  assign new_n23806 = new_n23805 ^ new_n23773;
  assign new_n23807 = new_n21930 ^ new_n21747;
  assign new_n23808 = new_n22027 ^ new_n21896;
  assign new_n23809 = new_n23808 ^ new_n23807;
  assign new_n23810 = new_n20856 ^ new_n16130;
  assign new_n23811 = new_n23810 ^ new_n8394;
  assign new_n23812 = new_n23811 ^ new_n21971;
  assign new_n23813 = new_n23812 ^ new_n22151;
  assign new_n23814 = new_n23813 ^ new_n23809;
  assign new_n23815 = new_n22118 ^ new_n21992;
  assign new_n23816 = new_n23815 ^ new_n22004;
  assign new_n23817 = new_n20798 ^ new_n16148;
  assign new_n23818 = new_n23817 ^ new_n8402;
  assign new_n23819 = new_n23818 ^ new_n21747;
  assign new_n23820 = new_n22113 ^ new_n22097;
  assign new_n23821 = new_n23820 ^ new_n23819;
  assign new_n23822 = new_n23821 ^ new_n23816;
  assign new_n23823 = new_n23822 ^ new_n23814;
  assign new_n23824 = new_n21906 ^ new_n21880;
  assign new_n23825 = new_n23824 ^ new_n21580;
  assign new_n23826 = new_n20957 ^ new_n16232;
  assign new_n23827 = new_n23826 ^ new_n8411;
  assign new_n23828 = new_n23827 ^ new_n21736;
  assign new_n23829 = new_n23828 ^ new_n22064;
  assign new_n23830 = new_n23829 ^ new_n23825;
  assign new_n23831 = new_n20971 ^ new_n16262;
  assign new_n23832 = new_n23831 ^ new_n8380;
  assign new_n23833 = new_n22106 ^ new_n22072;
  assign new_n23834 = new_n23833 ^ new_n23832;
  assign new_n23835 = new_n23834 ^ new_n21747;
  assign new_n23836 = new_n22104 ^ new_n22101;
  assign new_n23837 = new_n23836 ^ new_n22118;
  assign new_n23838 = new_n23837 ^ new_n23835;
  assign new_n23839 = new_n23838 ^ new_n23830;
  assign new_n23840 = new_n23839 ^ new_n23823;
  assign new_n23841 = new_n20936 ^ new_n16278;
  assign new_n23842 = new_n23841 ^ new_n8371;
  assign new_n23843 = new_n23842 ^ new_n22151;
  assign new_n23844 = new_n22144 ^ new_n21919;
  assign new_n23845 = new_n23844 ^ new_n21747;
  assign new_n23846 = new_n23845 ^ new_n23843;
  assign new_n23847 = new_n23846 ^ new_n23840;
  assign new_n23848 = new_n22129 ^ new_n21986;
  assign new_n23849 = new_n23848 ^ new_n21941;
  assign new_n23850 = new_n20430 ^ new_n15732;
  assign new_n23851 = new_n23850 ^ new_n8421;
  assign new_n23852 = new_n23851 ^ new_n22004;
  assign new_n23853 = new_n23852 ^ new_n21971;
  assign new_n23854 = new_n23853 ^ new_n23849;
  assign new_n23855 = new_n23854 ^ new_n23823;
  assign new_n23856 = new_n22037 ^ new_n21440;
  assign new_n23857 = new_n23856 ^ new_n22048;
  assign new_n23858 = new_n20898 ^ new_n16209;
  assign new_n23859 = new_n23858 ^ new_n8358;
  assign new_n23860 = new_n23859 ^ new_n22064;
  assign new_n23861 = new_n23860 ^ new_n22085;
  assign new_n23862 = new_n23861 ^ new_n23857;
  assign new_n23863 = new_n23862 ^ new_n23855;
  assign new_n23864 = new_n23863 ^ new_n23846;
  assign new_n23865 = new_n22071 ^ new_n22044;
  assign new_n23866 = new_n23865 ^ new_n22085;
  assign new_n23867 = new_n20927 ^ new_n16253;
  assign new_n23868 = new_n23867 ^ new_n8365;
  assign new_n23869 = new_n23868 ^ new_n22105;
  assign new_n23870 = new_n23869 ^ new_n23866;
  assign new_n23871 = new_n23870 ^ new_n23862;
  assign new_n23872 = new_n23871 ^ new_n23846;
  assign new_n23873 = new_n23872 ^ new_n23830;
  assign new_n23874 = ~new_n23864 & ~new_n23873;
  assign new_n23875 = new_n23830 ^ new_n23814;
  assign new_n23876 = new_n23870 ^ new_n23855;
  assign new_n23877 = ~new_n23875 & new_n23876;
  assign new_n23878 = new_n23877 ^ new_n23874;
  assign new_n23879 = new_n23878 ^ new_n23830;
  assign new_n23880 = new_n23854 ^ new_n23830;
  assign new_n23881 = new_n23871 ^ new_n23840;
  assign new_n23882 = ~new_n23881 & new_n23880;
  assign new_n23883 = new_n23839 & new_n23863;
  assign new_n23884 = new_n23883 ^ new_n23882;
  assign new_n23885 = new_n23884 ^ new_n23876;
  assign new_n23886 = new_n23885 ^ new_n23879;
  assign new_n23887 = new_n23814 & new_n23872;
  assign new_n23888 = new_n23887 ^ new_n23814;
  assign new_n23889 = new_n23888 ^ new_n23877;
  assign new_n23890 = new_n23889 ^ new_n23880;
  assign new_n23891 = new_n23854 ^ new_n23838;
  assign new_n23892 = new_n23870 ^ new_n23838;
  assign new_n23893 = new_n23892 ^ new_n23880;
  assign new_n23894 = ~new_n23893 & new_n23891;
  assign new_n23895 = new_n23894 ^ new_n23883;
  assign new_n23896 = new_n23870 ^ new_n23822;
  assign new_n23897 = new_n23896 ^ new_n23895;
  assign new_n23898 = new_n23897 ^ new_n23890;
  assign new_n23899 = new_n23891 ^ new_n23875;
  assign new_n23900 = ~new_n23840 & ~new_n23899;
  assign new_n23901 = new_n23900 ^ new_n23862;
  assign new_n23902 = new_n23901 ^ new_n23840;
  assign new_n23903 = new_n23872 ^ new_n23814;
  assign new_n23904 = new_n23903 ^ new_n23880;
  assign new_n23905 = new_n23847 & new_n23904;
  assign new_n23906 = new_n23905 ^ new_n23883;
  assign new_n23907 = new_n23894 ^ new_n23854;
  assign new_n23908 = new_n23907 ^ new_n23906;
  assign new_n23909 = new_n23908 ^ new_n23902;
  assign new_n23910 = ~new_n23898 & new_n23909;
  assign new_n23911 = new_n23872 ^ new_n23838;
  assign new_n23912 = ~new_n23846 & ~new_n23911;
  assign new_n23913 = new_n23912 ^ new_n23838;
  assign new_n23914 = new_n23913 ^ new_n23901;
  assign new_n23915 = new_n23914 ^ new_n23910;
  assign new_n23916 = new_n23915 ^ new_n23885;
  assign new_n23917 = new_n23894 ^ new_n23882;
  assign new_n23918 = new_n23887 ^ new_n23874;
  assign new_n23919 = new_n23918 ^ new_n23917;
  assign new_n23920 = ~new_n23916 & ~new_n23919;
  assign new_n23921 = new_n23920 ^ new_n23910;
  assign new_n23922 = ~new_n23921 & new_n23886;
  assign new_n23923 = new_n23922 ^ new_n23886;
  assign new_n23924 = new_n23923 ^ new_n23920;
  assign new_n23925 = new_n23924 ^ new_n23919;
  assign new_n23926 = ~new_n23925 & new_n23847;
  assign new_n23927 = new_n23923 ^ new_n23898;
  assign new_n23928 = ~new_n23840 & ~new_n23927;
  assign new_n23929 = new_n23928 ^ new_n23926;
  assign new_n23930 = ~new_n23899 & ~new_n23927;
  assign new_n23931 = new_n23930 ^ new_n23929;
  assign new_n23932 = ~new_n23925 & new_n23904;
  assign new_n23933 = new_n23870 ^ new_n23814;
  assign new_n23934 = new_n23905 ^ new_n23888;
  assign new_n23935 = new_n23870 ^ new_n23830;
  assign new_n23936 = new_n23912 ^ new_n23905;
  assign new_n23937 = new_n23936 ^ new_n23917;
  assign new_n23938 = new_n23937 ^ new_n23935;
  assign new_n23939 = new_n23910 ^ new_n23886;
  assign new_n23940 = ~new_n23938 & new_n23939;
  assign new_n23941 = new_n23940 ^ new_n23914;
  assign new_n23942 = new_n23941 ^ new_n23885;
  assign new_n23943 = new_n23922 ^ new_n23910;
  assign new_n23944 = ~new_n23942 & new_n23943;
  assign new_n23945 = new_n23944 ^ new_n23923;
  assign new_n23946 = new_n23945 ^ new_n23934;
  assign new_n23947 = new_n23946 ^ new_n23933;
  assign new_n23948 = new_n23947 ^ new_n23838;
  assign new_n23949 = new_n23940 ^ new_n23877;
  assign new_n23950 = new_n23949 ^ new_n23901;
  assign new_n23951 = new_n23950 ^ new_n23948;
  assign new_n23952 = ~new_n23951 & new_n23891;
  assign new_n23953 = new_n23940 ^ new_n23920;
  assign new_n23954 = new_n23914 ^ new_n23879;
  assign new_n23955 = new_n23954 ^ new_n23953;
  assign new_n23956 = ~new_n23955 & new_n23839;
  assign new_n23957 = new_n23956 ^ new_n23952;
  assign new_n23958 = new_n23957 ^ new_n23932;
  assign new_n23959 = new_n23944 ^ new_n23938;
  assign new_n23960 = ~new_n23872 & ~new_n23959;
  assign new_n23961 = new_n23960 ^ new_n23958;
  assign new_n23962 = new_n23944 ^ new_n23940;
  assign new_n23963 = new_n23962 ^ new_n23909;
  assign new_n23964 = new_n23876 & new_n23963;
  assign new_n23965 = new_n23964 ^ new_n23961;
  assign new_n23966 = new_n23965 ^ new_n23931;
  assign new_n23967 = new_n23966 ^ new_n23806;
  assign new_n23968 = ~new_n23955 & new_n23863;
  assign new_n23969 = new_n23968 ^ new_n23956;
  assign new_n23970 = new_n23920 ^ new_n23830;
  assign new_n23971 = new_n23912 ^ new_n23874;
  assign new_n23972 = new_n23971 ^ new_n23947;
  assign new_n23973 = new_n23972 ^ new_n23970;
  assign new_n23974 = new_n23880 & new_n23973;
  assign new_n23975 = ~new_n23873 & ~new_n23942;
  assign new_n23976 = ~new_n23881 & new_n23973;
  assign new_n23977 = new_n23976 ^ new_n23975;
  assign new_n23978 = ~new_n23875 & new_n23963;
  assign new_n23979 = new_n23920 ^ new_n23886;
  assign new_n23980 = ~new_n23846 & new_n23979;
  assign new_n23981 = new_n23980 ^ new_n23928;
  assign new_n23982 = new_n23981 ^ new_n23978;
  assign new_n23983 = new_n23982 ^ new_n23977;
  assign new_n23984 = new_n23983 ^ new_n23974;
  assign new_n23985 = new_n23984 ^ new_n23969;
  assign new_n23986 = new_n23985 ^ new_n23967;
  assign new_n23987 = new_n20659 ^ new_n19878;
  assign new_n23988 = new_n23987 ^ new_n18700;
  assign new_n23989 = new_n23988 ^ new_n18618;
  assign new_n23990 = new_n23989 ^ new_n23016;
  assign new_n23991 = new_n18557 ^ new_n15309;
  assign new_n23992 = new_n18710 ^ new_n18604;
  assign new_n23993 = new_n23992 ^ new_n23991;
  assign new_n23994 = new_n20638 ^ new_n19818;
  assign new_n23995 = new_n23994 ^ new_n18656;
  assign new_n23996 = new_n18826 ^ new_n18641;
  assign new_n23997 = new_n23996 ^ new_n23995;
  assign new_n23998 = new_n23997 ^ new_n23993;
  assign new_n23999 = new_n18799 ^ new_n18700;
  assign new_n24000 = new_n23999 ^ new_n18677;
  assign new_n24001 = new_n20644 ^ new_n19834;
  assign new_n24002 = new_n24001 ^ new_n23991;
  assign new_n24003 = new_n24002 ^ new_n22996;
  assign new_n24004 = new_n24003 ^ new_n24000;
  assign new_n24005 = new_n24004 ^ new_n23998;
  assign new_n24006 = new_n24005 ^ new_n23990;
  assign new_n24007 = new_n23021 ^ new_n18731;
  assign new_n24008 = new_n20614 ^ new_n19029;
  assign new_n24009 = new_n24008 ^ new_n18736;
  assign new_n24010 = new_n24009 ^ new_n18744;
  assign new_n24011 = new_n24010 ^ new_n24007;
  assign new_n24012 = new_n24011 ^ new_n24006;
  assign new_n24013 = new_n22983 ^ new_n18744;
  assign new_n24014 = new_n20631 ^ new_n19731;
  assign new_n24015 = new_n24014 ^ new_n15309;
  assign new_n24016 = new_n24015 ^ new_n18565;
  assign new_n24017 = new_n24016 ^ new_n24013;
  assign new_n24018 = new_n20649 ^ new_n19775;
  assign new_n24019 = new_n24018 ^ new_n23991;
  assign new_n24020 = new_n24019 ^ new_n22986;
  assign new_n24021 = new_n18799 ^ new_n18774;
  assign new_n24022 = new_n24021 ^ new_n18786;
  assign new_n24023 = new_n24022 ^ new_n24020;
  assign new_n24024 = new_n24023 ^ new_n24017;
  assign new_n24025 = new_n24024 ^ new_n24005;
  assign new_n24026 = new_n24023 ^ new_n23998;
  assign new_n24027 = new_n24017 ^ new_n23990;
  assign new_n24028 = new_n24027 ^ new_n24026;
  assign new_n24029 = ~new_n24025 & ~new_n24028;
  assign new_n24030 = new_n24029 ^ new_n24011;
  assign new_n24031 = new_n20624 ^ new_n19861;
  assign new_n24032 = new_n24031 ^ new_n18582;
  assign new_n24033 = new_n23991 ^ new_n23002;
  assign new_n24034 = new_n24033 ^ new_n24032;
  assign new_n24035 = new_n23029 ^ new_n18731;
  assign new_n24036 = new_n20620 ^ new_n19652;
  assign new_n24037 = new_n18774 ^ new_n18721;
  assign new_n24038 = new_n24037 ^ new_n24036;
  assign new_n24039 = new_n24038 ^ new_n24035;
  assign new_n24040 = new_n24039 ^ new_n24011;
  assign new_n24041 = ~new_n24034 & ~new_n24040;
  assign new_n24042 = new_n24023 & new_n24034;
  assign new_n24043 = new_n24042 ^ new_n24041;
  assign new_n24044 = new_n24043 ^ new_n24030;
  assign new_n24045 = new_n24040 ^ new_n24034;
  assign new_n24046 = new_n23998 & new_n24045;
  assign new_n24047 = new_n24046 ^ new_n23998;
  assign new_n24048 = new_n24039 ^ new_n24006;
  assign new_n24049 = new_n24017 ^ new_n23998;
  assign new_n24050 = ~new_n24049 & new_n24048;
  assign new_n24051 = new_n24050 ^ new_n24047;
  assign new_n24052 = new_n24051 ^ new_n24027;
  assign new_n24053 = new_n24012 & new_n24024;
  assign new_n24054 = new_n24039 ^ new_n24023;
  assign new_n24055 = new_n24054 ^ new_n24027;
  assign new_n24056 = new_n24023 ^ new_n23990;
  assign new_n24057 = ~new_n24055 & new_n24056;
  assign new_n24058 = new_n24057 ^ new_n24053;
  assign new_n24059 = new_n24039 ^ new_n24004;
  assign new_n24060 = new_n24059 ^ new_n24058;
  assign new_n24061 = new_n24060 ^ new_n24052;
  assign new_n24062 = new_n24030 ^ new_n24025;
  assign new_n24063 = new_n24034 ^ new_n24025;
  assign new_n24064 = new_n24045 ^ new_n23998;
  assign new_n24065 = new_n24064 ^ new_n24027;
  assign new_n24066 = new_n24063 & new_n24065;
  assign new_n24067 = new_n24066 ^ new_n24058;
  assign new_n24068 = new_n24067 ^ new_n23990;
  assign new_n24069 = new_n24068 ^ new_n24062;
  assign new_n24070 = ~new_n24061 & new_n24069;
  assign new_n24071 = new_n24070 ^ new_n24044;
  assign new_n24072 = new_n24040 ^ new_n24025;
  assign new_n24073 = ~new_n24072 & new_n24027;
  assign new_n24074 = new_n24073 ^ new_n24053;
  assign new_n24075 = new_n24074 ^ new_n24048;
  assign new_n24076 = new_n24075 ^ new_n24071;
  assign new_n24077 = new_n24045 ^ new_n24017;
  assign new_n24078 = new_n24034 ^ new_n24012;
  assign new_n24079 = ~new_n24077 & ~new_n24078;
  assign new_n24080 = new_n24079 ^ new_n24046;
  assign new_n24081 = new_n24073 ^ new_n24057;
  assign new_n24082 = new_n24081 ^ new_n24080;
  assign new_n24083 = ~new_n24076 & ~new_n24082;
  assign new_n24084 = new_n24039 ^ new_n24017;
  assign new_n24085 = new_n24043 ^ new_n24023;
  assign new_n24086 = new_n24085 ^ new_n24066;
  assign new_n24087 = new_n24086 ^ new_n24081;
  assign new_n24088 = new_n24087 ^ new_n24084;
  assign new_n24089 = new_n24079 ^ new_n24050;
  assign new_n24090 = new_n24089 ^ new_n24017;
  assign new_n24091 = new_n24090 ^ new_n24075;
  assign new_n24092 = new_n24091 ^ new_n24070;
  assign new_n24093 = ~new_n24088 & new_n24092;
  assign new_n24094 = new_n24093 ^ new_n24083;
  assign new_n24095 = new_n24090 ^ new_n24044;
  assign new_n24096 = new_n24095 ^ new_n24094;
  assign new_n24097 = ~new_n24096 & new_n24012;
  assign new_n24098 = ~new_n24096 & new_n24024;
  assign new_n24099 = new_n24098 ^ new_n24097;
  assign new_n24100 = new_n24093 ^ new_n24044;
  assign new_n24101 = new_n24100 ^ new_n24075;
  assign new_n24102 = ~new_n24077 & ~new_n24101;
  assign new_n24103 = new_n24083 ^ new_n24017;
  assign new_n24104 = new_n24085 ^ new_n24079;
  assign new_n24105 = new_n24039 ^ new_n23998;
  assign new_n24106 = new_n24066 ^ new_n24047;
  assign new_n24107 = new_n24083 ^ new_n24070;
  assign new_n24108 = new_n24091 & new_n24107;
  assign new_n24109 = new_n24108 ^ new_n24092;
  assign new_n24110 = ~new_n24101 & new_n24109;
  assign new_n24111 = new_n24110 ^ new_n24108;
  assign new_n24112 = new_n24111 ^ new_n24106;
  assign new_n24113 = new_n24112 ^ new_n24105;
  assign new_n24114 = new_n24113 ^ new_n24104;
  assign new_n24115 = new_n24114 ^ new_n24103;
  assign new_n24116 = ~new_n24072 & new_n24115;
  assign new_n24117 = new_n24116 ^ new_n24102;
  assign new_n24118 = new_n24108 ^ new_n24061;
  assign new_n24119 = ~new_n24025 & ~new_n24118;
  assign new_n24120 = new_n24091 ^ new_n24083;
  assign new_n24121 = ~new_n24034 & new_n24120;
  assign new_n24122 = new_n24121 ^ new_n24119;
  assign new_n24123 = new_n24110 ^ new_n24093;
  assign new_n24124 = new_n24123 ^ new_n24069;
  assign new_n24125 = ~new_n24049 & new_n24124;
  assign new_n24126 = new_n24125 ^ new_n24122;
  assign new_n24127 = new_n24126 ^ new_n24117;
  assign new_n24128 = new_n24027 & new_n24115;
  assign new_n24129 = new_n24128 ^ new_n24127;
  assign new_n24130 = new_n24129 ^ new_n24099;
  assign new_n24131 = new_n20857 ^ new_n20799;
  assign new_n24132 = new_n24131 ^ new_n20431;
  assign new_n24133 = new_n24132 ^ new_n20899;
  assign new_n24134 = new_n20928 ^ new_n20899;
  assign new_n24135 = new_n24134 ^ new_n20937;
  assign new_n24136 = new_n24135 ^ new_n20972;
  assign new_n24137 = new_n20937 & new_n24136;
  assign new_n24138 = new_n24137 ^ new_n20972;
  assign new_n24139 = new_n20972 ^ new_n20958;
  assign new_n24140 = new_n24139 ^ new_n24131;
  assign new_n24141 = new_n20972 ^ new_n20857;
  assign new_n24142 = new_n20958 ^ new_n20431;
  assign new_n24143 = new_n24142 ^ new_n24141;
  assign new_n24144 = new_n24140 & new_n24143;
  assign new_n24145 = new_n24144 ^ new_n20899;
  assign new_n24146 = new_n24145 ^ new_n24138;
  assign new_n24147 = new_n24145 ^ new_n24140;
  assign new_n24148 = new_n24133 & new_n24139;
  assign new_n24149 = new_n20972 ^ new_n20928;
  assign new_n24150 = new_n24149 ^ new_n24142;
  assign new_n24151 = new_n20972 ^ new_n20431;
  assign new_n24152 = new_n24150 & new_n24151;
  assign new_n24153 = new_n24152 ^ new_n24148;
  assign new_n24154 = new_n24140 ^ new_n20937;
  assign new_n24155 = new_n24135 ^ new_n20857;
  assign new_n24156 = new_n24155 ^ new_n24142;
  assign new_n24157 = new_n24154 & new_n24156;
  assign new_n24158 = new_n24157 ^ new_n20431;
  assign new_n24159 = new_n24158 ^ new_n24153;
  assign new_n24160 = new_n24159 ^ new_n24147;
  assign new_n24161 = ~new_n20857 & ~new_n24135;
  assign new_n24162 = new_n24161 ^ new_n20857;
  assign new_n24163 = new_n24132 ^ new_n20928;
  assign new_n24164 = new_n20958 ^ new_n20857;
  assign new_n24165 = new_n24163 & new_n24164;
  assign new_n24166 = new_n24165 ^ new_n24162;
  assign new_n24167 = new_n24166 ^ new_n24142;
  assign new_n24168 = new_n20928 ^ new_n20799;
  assign new_n24169 = new_n24168 ^ new_n24153;
  assign new_n24170 = new_n24169 ^ new_n24167;
  assign new_n24171 = ~new_n24170 & new_n24160;
  assign new_n24172 = new_n24171 ^ new_n24146;
  assign new_n24173 = new_n24140 ^ new_n24134;
  assign new_n24174 = new_n24142 & new_n24173;
  assign new_n24175 = new_n24174 ^ new_n24148;
  assign new_n24176 = new_n24175 ^ new_n24163;
  assign new_n24177 = new_n24176 ^ new_n24172;
  assign new_n24178 = new_n24135 ^ new_n20958;
  assign new_n24179 = new_n24133 ^ new_n20937;
  assign new_n24180 = new_n24178 & new_n24179;
  assign new_n24181 = new_n24180 ^ new_n24161;
  assign new_n24182 = new_n24174 ^ new_n24152;
  assign new_n24183 = new_n24182 ^ new_n24181;
  assign new_n24184 = ~new_n24183 & new_n24177;
  assign new_n24185 = new_n20958 ^ new_n20928;
  assign new_n24186 = new_n24157 ^ new_n24137;
  assign new_n24187 = new_n24186 ^ new_n24182;
  assign new_n24188 = new_n24187 ^ new_n24185;
  assign new_n24189 = new_n24180 ^ new_n24165;
  assign new_n24190 = new_n24189 ^ new_n20958;
  assign new_n24191 = new_n24190 ^ new_n24176;
  assign new_n24192 = new_n24191 ^ new_n24171;
  assign new_n24193 = new_n24188 & new_n24192;
  assign new_n24194 = new_n24193 ^ new_n24184;
  assign new_n24195 = new_n24190 ^ new_n24146;
  assign new_n24196 = new_n24195 ^ new_n24194;
  assign new_n24197 = new_n24133 & new_n24196;
  assign new_n24198 = new_n24139 & new_n24196;
  assign new_n24199 = new_n24198 ^ new_n24197;
  assign new_n24200 = new_n24184 ^ new_n20958;
  assign new_n24201 = new_n24180 ^ new_n24137;
  assign new_n24202 = new_n20928 ^ new_n20857;
  assign new_n24203 = new_n24162 ^ new_n24157;
  assign new_n24204 = new_n24193 ^ new_n24146;
  assign new_n24205 = new_n24204 ^ new_n24176;
  assign new_n24206 = new_n24184 ^ new_n24171;
  assign new_n24207 = new_n24191 & new_n24206;
  assign new_n24208 = new_n24207 ^ new_n24192;
  assign new_n24209 = new_n24205 & new_n24208;
  assign new_n24210 = new_n24209 ^ new_n24207;
  assign new_n24211 = new_n24210 ^ new_n24203;
  assign new_n24212 = new_n24211 ^ new_n24202;
  assign new_n24213 = new_n24212 ^ new_n24201;
  assign new_n24214 = new_n24213 ^ new_n24200;
  assign new_n24215 = ~new_n24214 & new_n24142;
  assign new_n24216 = new_n24178 & new_n24205;
  assign new_n24217 = ~new_n24214 & new_n24173;
  assign new_n24218 = new_n24217 ^ new_n24216;
  assign new_n24219 = new_n24191 ^ new_n24184;
  assign new_n24220 = new_n20937 & new_n24219;
  assign new_n24221 = new_n24207 ^ new_n24170;
  assign new_n24222 = ~new_n24221 & new_n24140;
  assign new_n24223 = new_n24222 ^ new_n24220;
  assign new_n24224 = new_n24209 ^ new_n24193;
  assign new_n24225 = new_n24224 ^ new_n24160;
  assign new_n24226 = new_n24164 & new_n24225;
  assign new_n24227 = new_n24226 ^ new_n24223;
  assign new_n24228 = new_n24227 ^ new_n24218;
  assign new_n24229 = new_n24228 ^ new_n24215;
  assign new_n24230 = new_n24229 ^ new_n24199;
  assign new_n24231 = new_n24230 ^ new_n9025;
  assign new_n24232 = new_n24231 ^ new_n24130;
  assign new_n24233 = new_n20820 ^ new_n20611;
  assign new_n24234 = new_n24233 ^ new_n20771;
  assign new_n24235 = new_n20977 ^ new_n20827;
  assign new_n24236 = new_n24235 ^ new_n21081;
  assign new_n24237 = new_n20948 ^ new_n20777;
  assign new_n24238 = new_n24237 ^ new_n24236;
  assign new_n24239 = new_n24238 ^ new_n24234;
  assign new_n24240 = new_n20811 ^ new_n20591;
  assign new_n24241 = new_n24240 ^ new_n20312;
  assign new_n24242 = new_n21091 ^ new_n20771;
  assign new_n24243 = new_n24242 ^ new_n20865;
  assign new_n24244 = new_n24243 ^ new_n24241;
  assign new_n24245 = new_n24244 ^ new_n24239;
  assign new_n24246 = new_n24237 ^ new_n20838;
  assign new_n24247 = new_n20849 ^ new_n20165;
  assign new_n24248 = new_n24247 ^ new_n24246;
  assign new_n24249 = new_n21080 ^ new_n20865;
  assign new_n24250 = new_n24249 ^ new_n20940;
  assign new_n24251 = new_n24250 ^ new_n24248;
  assign new_n24252 = new_n24251 ^ new_n24245;
  assign new_n24253 = new_n22876 ^ new_n20904;
  assign new_n24254 = new_n21074 ^ new_n20881;
  assign new_n24255 = new_n24254 ^ new_n20915;
  assign new_n24256 = new_n24255 ^ new_n24253;
  assign new_n24257 = new_n24256 ^ new_n24252;
  assign new_n24258 = new_n22839 ^ new_n20892;
  assign new_n24259 = new_n21077 ^ new_n20948;
  assign new_n24260 = new_n24259 ^ new_n20881;
  assign new_n24261 = new_n24260 ^ new_n24258;
  assign new_n24262 = new_n24237 ^ new_n21078;
  assign new_n24263 = new_n24262 ^ new_n22844;
  assign new_n24264 = new_n20968 ^ new_n20833;
  assign new_n24265 = new_n24264 ^ new_n20820;
  assign new_n24266 = new_n24265 ^ new_n24263;
  assign new_n24267 = new_n24266 ^ new_n24261;
  assign new_n24268 = new_n24251 ^ new_n24239;
  assign new_n24269 = new_n24268 ^ new_n24267;
  assign new_n24270 = new_n24266 ^ new_n24251;
  assign new_n24271 = new_n24261 ^ new_n24244;
  assign new_n24272 = new_n24271 ^ new_n24270;
  assign new_n24273 = new_n24269 & new_n24272;
  assign new_n24274 = new_n24273 ^ new_n24256;
  assign new_n24275 = new_n21085 ^ new_n20940;
  assign new_n24276 = new_n20934 ^ new_n20840;
  assign new_n24277 = new_n24276 ^ new_n24237;
  assign new_n24278 = new_n24277 ^ new_n24275;
  assign new_n24279 = new_n20968 ^ new_n20922;
  assign new_n24280 = new_n24279 ^ new_n21075;
  assign new_n24281 = new_n22884 ^ new_n20915;
  assign new_n24282 = new_n24281 ^ new_n24280;
  assign new_n24283 = new_n24282 ^ new_n24256;
  assign new_n24284 = ~new_n24278 & new_n24283;
  assign new_n24285 = new_n24266 & new_n24278;
  assign new_n24286 = new_n24285 ^ new_n24284;
  assign new_n24287 = new_n24286 ^ new_n24274;
  assign new_n24288 = new_n24283 ^ new_n24278;
  assign new_n24289 = ~new_n24251 & ~new_n24288;
  assign new_n24290 = new_n24289 ^ new_n24251;
  assign new_n24291 = new_n24282 ^ new_n24252;
  assign new_n24292 = new_n24261 ^ new_n24251;
  assign new_n24293 = new_n24291 & new_n24292;
  assign new_n24294 = new_n24293 ^ new_n24290;
  assign new_n24295 = new_n24294 ^ new_n24271;
  assign new_n24296 = ~new_n24257 & new_n24267;
  assign new_n24297 = new_n24282 ^ new_n24266;
  assign new_n24298 = new_n24297 ^ new_n24271;
  assign new_n24299 = new_n24266 ^ new_n24244;
  assign new_n24300 = new_n24298 & new_n24299;
  assign new_n24301 = new_n24300 ^ new_n24296;
  assign new_n24302 = new_n24282 ^ new_n24239;
  assign new_n24303 = new_n24302 ^ new_n24301;
  assign new_n24304 = new_n24303 ^ new_n24295;
  assign new_n24305 = new_n24274 ^ new_n24269;
  assign new_n24306 = new_n24288 ^ new_n24251;
  assign new_n24307 = new_n24306 ^ new_n24271;
  assign new_n24308 = new_n24278 ^ new_n24269;
  assign new_n24309 = ~new_n24308 & new_n24307;
  assign new_n24310 = new_n24309 ^ new_n24296;
  assign new_n24311 = new_n24300 ^ new_n24244;
  assign new_n24312 = new_n24311 ^ new_n24310;
  assign new_n24313 = new_n24312 ^ new_n24305;
  assign new_n24314 = ~new_n24304 & ~new_n24313;
  assign new_n24315 = new_n24314 ^ new_n24287;
  assign new_n24316 = new_n24283 ^ new_n24269;
  assign new_n24317 = ~new_n24316 & new_n24271;
  assign new_n24318 = new_n24317 ^ new_n24296;
  assign new_n24319 = new_n24318 ^ new_n24291;
  assign new_n24320 = new_n24319 ^ new_n24315;
  assign new_n24321 = new_n24288 ^ new_n24261;
  assign new_n24322 = new_n24278 ^ new_n24257;
  assign new_n24323 = new_n24321 & new_n24322;
  assign new_n24324 = new_n24323 ^ new_n24289;
  assign new_n24325 = new_n24317 ^ new_n24300;
  assign new_n24326 = new_n24325 ^ new_n24324;
  assign new_n24327 = ~new_n24320 & ~new_n24326;
  assign new_n24328 = new_n24282 ^ new_n24261;
  assign new_n24329 = new_n24286 ^ new_n24266;
  assign new_n24330 = new_n24329 ^ new_n24309;
  assign new_n24331 = new_n24330 ^ new_n24325;
  assign new_n24332 = new_n24331 ^ new_n24328;
  assign new_n24333 = new_n24323 ^ new_n24293;
  assign new_n24334 = new_n24333 ^ new_n24261;
  assign new_n24335 = new_n24334 ^ new_n24319;
  assign new_n24336 = new_n24335 ^ new_n24314;
  assign new_n24337 = new_n24332 & new_n24336;
  assign new_n24338 = new_n24337 ^ new_n24327;
  assign new_n24339 = new_n24334 ^ new_n24287;
  assign new_n24340 = new_n24339 ^ new_n24338;
  assign new_n24341 = ~new_n24257 & ~new_n24340;
  assign new_n24342 = ~new_n24340 & new_n24267;
  assign new_n24343 = new_n24342 ^ new_n24341;
  assign new_n24344 = new_n24337 ^ new_n24287;
  assign new_n24345 = new_n24344 ^ new_n24319;
  assign new_n24346 = ~new_n24345 & new_n24321;
  assign new_n24347 = new_n24327 ^ new_n24261;
  assign new_n24348 = new_n24329 ^ new_n24323;
  assign new_n24349 = new_n24282 ^ new_n24251;
  assign new_n24350 = new_n24309 ^ new_n24290;
  assign new_n24351 = new_n24327 ^ new_n24314;
  assign new_n24352 = new_n24335 & new_n24351;
  assign new_n24353 = new_n24352 ^ new_n24336;
  assign new_n24354 = ~new_n24345 & new_n24353;
  assign new_n24355 = new_n24354 ^ new_n24352;
  assign new_n24356 = new_n24355 ^ new_n24350;
  assign new_n24357 = new_n24356 ^ new_n24349;
  assign new_n24358 = new_n24357 ^ new_n24348;
  assign new_n24359 = new_n24358 ^ new_n24347;
  assign new_n24360 = ~new_n24316 & ~new_n24359;
  assign new_n24361 = new_n24360 ^ new_n24346;
  assign new_n24362 = new_n24352 ^ new_n24304;
  assign new_n24363 = ~new_n24362 & new_n24269;
  assign new_n24364 = new_n24335 ^ new_n24327;
  assign new_n24365 = ~new_n24278 & new_n24364;
  assign new_n24366 = new_n24365 ^ new_n24363;
  assign new_n24367 = new_n24354 ^ new_n24337;
  assign new_n24368 = new_n24367 ^ new_n24313;
  assign new_n24369 = ~new_n24368 & new_n24292;
  assign new_n24370 = new_n24369 ^ new_n24366;
  assign new_n24371 = new_n24370 ^ new_n24361;
  assign new_n24372 = ~new_n24359 & new_n24271;
  assign new_n24373 = new_n24372 ^ new_n24371;
  assign new_n24374 = new_n24373 ^ new_n24343;
  assign new_n24375 = new_n24374 ^ new_n24232;
  assign new_n24376 = new_n24375 ^ new_n23986;
  assign new_n24377 = new_n23705 & new_n23797;
  assign new_n24378 = new_n24377 ^ new_n23798;
  assign new_n24379 = new_n23760 ^ new_n23680;
  assign new_n24380 = new_n23729 ^ new_n23715;
  assign new_n24381 = new_n24380 ^ new_n23789;
  assign new_n24382 = new_n24381 ^ new_n24379;
  assign new_n24383 = new_n23721 & new_n24382;
  assign new_n24384 = new_n23722 & new_n24382;
  assign new_n24385 = new_n23714 & new_n23780;
  assign new_n24386 = new_n24385 ^ new_n24384;
  assign new_n24387 = new_n23717 & new_n23803;
  assign new_n24388 = new_n23760 ^ new_n23727;
  assign new_n24389 = new_n23692 & new_n24388;
  assign new_n24390 = new_n24389 ^ new_n23770;
  assign new_n24391 = new_n24390 ^ new_n24387;
  assign new_n24392 = new_n24391 ^ new_n24386;
  assign new_n24393 = new_n24392 ^ new_n24383;
  assign new_n24394 = new_n24393 ^ new_n24378;
  assign new_n24395 = new_n24394 ^ new_n23985;
  assign new_n24396 = ~new_n23893 & ~new_n23951;
  assign new_n24397 = new_n24396 ^ new_n23968;
  assign new_n24398 = new_n23958 ^ new_n23931;
  assign new_n24399 = new_n24398 ^ new_n24397;
  assign new_n24400 = new_n24399 ^ new_n24395;
  assign new_n24401 = new_n24113 ^ new_n24023;
  assign new_n24402 = new_n24093 ^ new_n24050;
  assign new_n24403 = new_n24402 ^ new_n24030;
  assign new_n24404 = new_n24403 ^ new_n24401;
  assign new_n24405 = ~new_n24055 & ~new_n24404;
  assign new_n24406 = new_n24405 ^ new_n24097;
  assign new_n24407 = new_n24108 ^ new_n24083;
  assign new_n24408 = new_n24407 ^ new_n24082;
  assign new_n24409 = ~new_n24408 & new_n24063;
  assign new_n24410 = new_n24409 ^ new_n24119;
  assign new_n24411 = ~new_n24028 & ~new_n24118;
  assign new_n24412 = new_n24411 ^ new_n24410;
  assign new_n24413 = ~new_n24408 & new_n24065;
  assign new_n24414 = ~new_n24404 & new_n24056;
  assign new_n24415 = new_n24414 ^ new_n24098;
  assign new_n24416 = new_n24415 ^ new_n24413;
  assign new_n24417 = new_n24416 ^ new_n24412;
  assign new_n24418 = new_n24417 ^ new_n24406;
  assign new_n24419 = new_n24212 ^ new_n20972;
  assign new_n24420 = new_n24193 ^ new_n24165;
  assign new_n24421 = new_n24420 ^ new_n24145;
  assign new_n24422 = new_n24421 ^ new_n24419;
  assign new_n24423 = ~new_n24422 & new_n24150;
  assign new_n24424 = new_n24423 ^ new_n24197;
  assign new_n24425 = new_n24207 ^ new_n24184;
  assign new_n24426 = new_n24425 ^ new_n24183;
  assign new_n24427 = ~new_n24426 & new_n24154;
  assign new_n24428 = new_n24427 ^ new_n24222;
  assign new_n24429 = ~new_n24221 & new_n24143;
  assign new_n24430 = new_n24429 ^ new_n24428;
  assign new_n24431 = ~new_n24426 & new_n24156;
  assign new_n24432 = ~new_n24422 & new_n24151;
  assign new_n24433 = new_n24432 ^ new_n24198;
  assign new_n24434 = new_n24433 ^ new_n24431;
  assign new_n24435 = new_n24434 ^ new_n24430;
  assign new_n24436 = new_n24435 ^ new_n24424;
  assign new_n24437 = new_n24436 ^ new_n8986;
  assign new_n24438 = new_n24437 ^ new_n24418;
  assign new_n24439 = new_n24357 ^ new_n24266;
  assign new_n24440 = new_n24337 ^ new_n24293;
  assign new_n24441 = new_n24440 ^ new_n24274;
  assign new_n24442 = new_n24441 ^ new_n24439;
  assign new_n24443 = new_n24298 & new_n24442;
  assign new_n24444 = new_n24443 ^ new_n24341;
  assign new_n24445 = new_n24352 ^ new_n24327;
  assign new_n24446 = new_n24445 ^ new_n24326;
  assign new_n24447 = ~new_n24308 & ~new_n24446;
  assign new_n24448 = new_n24447 ^ new_n24363;
  assign new_n24449 = ~new_n24362 & new_n24272;
  assign new_n24450 = new_n24449 ^ new_n24448;
  assign new_n24451 = ~new_n24446 & new_n24307;
  assign new_n24452 = new_n24299 & new_n24442;
  assign new_n24453 = new_n24452 ^ new_n24342;
  assign new_n24454 = new_n24453 ^ new_n24451;
  assign new_n24455 = new_n24454 ^ new_n24450;
  assign new_n24456 = new_n24455 ^ new_n24444;
  assign new_n24457 = new_n24456 ^ new_n24438;
  assign new_n24458 = new_n24457 ^ new_n24400;
  assign new_n24459 = new_n24458 ^ new_n24376;
  assign new_n24460 = new_n24048 & new_n24124;
  assign new_n24461 = new_n24460 ^ new_n24126;
  assign new_n24462 = new_n24110 ^ new_n24088;
  assign new_n24463 = ~new_n24462 & new_n24064;
  assign new_n24464 = ~new_n24078 & ~new_n24101;
  assign new_n24465 = new_n24464 ^ new_n24463;
  assign new_n24466 = new_n24465 ^ new_n24415;
  assign new_n24467 = new_n24466 ^ new_n24461;
  assign new_n24468 = new_n24163 & new_n24225;
  assign new_n24469 = new_n24468 ^ new_n24227;
  assign new_n24470 = new_n24209 ^ new_n24188;
  assign new_n24471 = new_n24155 & new_n24470;
  assign new_n24472 = new_n24179 & new_n24205;
  assign new_n24473 = new_n24472 ^ new_n24471;
  assign new_n24474 = new_n24473 ^ new_n24433;
  assign new_n24475 = new_n24474 ^ new_n24469;
  assign new_n24476 = new_n24475 ^ new_n9002;
  assign new_n24477 = new_n24476 ^ new_n24467;
  assign new_n24478 = ~new_n24368 & new_n24291;
  assign new_n24479 = new_n24478 ^ new_n24370;
  assign new_n24480 = new_n24354 ^ new_n24332;
  assign new_n24481 = new_n24306 & new_n24480;
  assign new_n24482 = ~new_n24345 & new_n24322;
  assign new_n24483 = new_n24482 ^ new_n24481;
  assign new_n24484 = new_n24483 ^ new_n24453;
  assign new_n24485 = new_n24484 ^ new_n24479;
  assign new_n24486 = ~new_n23864 & ~new_n23942;
  assign new_n24487 = ~new_n23959 & new_n23903;
  assign new_n24488 = new_n24487 ^ new_n24486;
  assign new_n24489 = new_n24488 ^ new_n23957;
  assign new_n24490 = new_n23982 ^ new_n23964;
  assign new_n24491 = new_n24490 ^ new_n24489;
  assign new_n24492 = new_n24491 ^ new_n24485;
  assign new_n24493 = new_n23968 ^ new_n23930;
  assign new_n24494 = new_n24396 ^ new_n23965;
  assign new_n24495 = new_n24494 ^ new_n24493;
  assign new_n24496 = new_n24377 ^ new_n23772;
  assign new_n24497 = new_n23741 & new_n23793;
  assign new_n24498 = new_n24497 ^ new_n23805;
  assign new_n24499 = new_n24498 ^ new_n24496;
  assign new_n24500 = new_n24499 ^ new_n24495;
  assign new_n24501 = new_n24500 ^ new_n24492;
  assign new_n24502 = new_n24501 ^ new_n24477;
  assign new_n24503 = new_n24502 ^ new_n24459;
  assign new_n24504 = new_n23706 & new_n23780;
  assign new_n24505 = new_n24504 ^ new_n23772;
  assign new_n24506 = new_n24389 ^ new_n23768;
  assign new_n24507 = new_n24506 ^ new_n23801;
  assign new_n24508 = new_n24507 ^ new_n24505;
  assign new_n24509 = new_n24486 ^ new_n23930;
  assign new_n24510 = new_n23980 ^ new_n23926;
  assign new_n24511 = new_n24510 ^ new_n23961;
  assign new_n24512 = new_n24511 ^ new_n24509;
  assign new_n24513 = new_n24512 ^ new_n24508;
  assign new_n24514 = new_n24135 & new_n24470;
  assign new_n24515 = new_n24514 ^ new_n24434;
  assign new_n24516 = new_n24515 ^ new_n24468;
  assign new_n24517 = new_n24516 ^ new_n24430;
  assign new_n24518 = new_n24517 ^ new_n9066;
  assign new_n24519 = new_n24518 ^ new_n24513;
  assign new_n24520 = new_n24519 ^ new_n24500;
  assign new_n24521 = new_n24288 & new_n24480;
  assign new_n24522 = new_n24521 ^ new_n24454;
  assign new_n24523 = new_n24522 ^ new_n24478;
  assign new_n24524 = new_n24523 ^ new_n24450;
  assign new_n24525 = new_n24524 ^ new_n23966;
  assign new_n24526 = ~new_n24045 & ~new_n24462;
  assign new_n24527 = new_n24526 ^ new_n24416;
  assign new_n24528 = new_n24527 ^ new_n24460;
  assign new_n24529 = new_n24528 ^ new_n24412;
  assign new_n24530 = new_n24529 ^ new_n24525;
  assign new_n24531 = new_n24530 ^ new_n24520;
  assign new_n24532 = new_n24531 ^ new_n24503;
  assign new_n24533 = ~new_n24502 & ~new_n24532;
  assign new_n24534 = new_n24533 ^ new_n24531;
  assign new_n24535 = new_n24497 ^ new_n24377;
  assign new_n24536 = new_n23800 ^ new_n23773;
  assign new_n24537 = new_n24536 ^ new_n24535;
  assign new_n24538 = new_n24537 ^ new_n24399;
  assign new_n24539 = new_n24429 ^ new_n24197;
  assign new_n24540 = new_n24516 ^ new_n24423;
  assign new_n24541 = new_n24540 ^ new_n24539;
  assign new_n24542 = new_n24541 ^ new_n9045;
  assign new_n24543 = new_n24542 ^ new_n24538;
  assign new_n24544 = new_n24449 ^ new_n24341;
  assign new_n24545 = new_n24523 ^ new_n24443;
  assign new_n24546 = new_n24545 ^ new_n24544;
  assign new_n24547 = new_n24546 ^ new_n24495;
  assign new_n24548 = new_n24411 ^ new_n24097;
  assign new_n24549 = new_n24528 ^ new_n24405;
  assign new_n24550 = new_n24549 ^ new_n24548;
  assign new_n24551 = new_n24550 ^ new_n24547;
  assign new_n24552 = new_n24551 ^ new_n24543;
  assign new_n24553 = new_n24552 ^ new_n24531;
  assign new_n24554 = new_n24464 ^ new_n24411;
  assign new_n24555 = new_n24409 ^ new_n24121;
  assign new_n24556 = new_n24555 ^ new_n24527;
  assign new_n24557 = new_n24556 ^ new_n24554;
  assign new_n24558 = new_n24472 ^ new_n24429;
  assign new_n24559 = new_n24427 ^ new_n24220;
  assign new_n24560 = new_n24559 ^ new_n24515;
  assign new_n24561 = new_n24560 ^ new_n24558;
  assign new_n24562 = new_n24561 ^ new_n8932;
  assign new_n24563 = new_n24562 ^ new_n24557;
  assign new_n24564 = new_n23728 & new_n24388;
  assign new_n24565 = new_n24564 ^ new_n24498;
  assign new_n24566 = new_n24565 ^ new_n24392;
  assign new_n24567 = ~new_n23911 & new_n23979;
  assign new_n24568 = new_n24567 ^ new_n24494;
  assign new_n24569 = new_n24568 ^ new_n23983;
  assign new_n24570 = new_n24569 ^ new_n24566;
  assign new_n24571 = new_n24570 ^ new_n24563;
  assign new_n24572 = new_n24482 ^ new_n24449;
  assign new_n24573 = new_n24447 ^ new_n24365;
  assign new_n24574 = new_n24573 ^ new_n24522;
  assign new_n24575 = new_n24574 ^ new_n24572;
  assign new_n24576 = new_n24575 ^ new_n24512;
  assign new_n24577 = new_n24576 ^ new_n24500;
  assign new_n24578 = new_n24577 ^ new_n24571;
  assign new_n24579 = new_n23978 ^ new_n23976;
  assign new_n24580 = new_n24396 ^ new_n23960;
  assign new_n24581 = new_n24580 ^ new_n24489;
  assign new_n24582 = new_n24581 ^ new_n24579;
  assign new_n24583 = new_n24369 ^ new_n24360;
  assign new_n24584 = new_n24521 ^ new_n24443;
  assign new_n24585 = new_n24584 ^ new_n24484;
  assign new_n24586 = new_n24585 ^ new_n24583;
  assign new_n24587 = new_n24586 ^ new_n24582;
  assign new_n24588 = new_n24587 ^ new_n24500;
  assign new_n24589 = new_n24125 ^ new_n24116;
  assign new_n24590 = new_n24526 ^ new_n24405;
  assign new_n24591 = new_n24590 ^ new_n24466;
  assign new_n24592 = new_n24591 ^ new_n24589;
  assign new_n24593 = new_n24226 ^ new_n24217;
  assign new_n24594 = new_n24514 ^ new_n24423;
  assign new_n24595 = new_n24594 ^ new_n24474;
  assign new_n24596 = new_n24595 ^ new_n24593;
  assign new_n24597 = new_n24596 ^ new_n8905;
  assign new_n24598 = new_n24597 ^ new_n24592;
  assign new_n24599 = new_n23748 & new_n23782;
  assign new_n24600 = new_n24599 ^ new_n24504;
  assign new_n24601 = new_n24600 ^ new_n23799;
  assign new_n24602 = new_n24391 ^ new_n23804;
  assign new_n24603 = new_n24602 ^ new_n24601;
  assign new_n24604 = new_n24603 ^ new_n24491;
  assign new_n24605 = new_n24604 ^ new_n24598;
  assign new_n24606 = new_n24605 ^ new_n24588;
  assign new_n24607 = new_n24606 ^ new_n24578;
  assign new_n24608 = new_n24607 ^ new_n24553;
  assign new_n24609 = new_n24606 ^ new_n24531;
  assign new_n24610 = new_n24045 ^ new_n24023;
  assign new_n24611 = ~new_n24610 & new_n24120;
  assign new_n24612 = new_n24611 ^ new_n24549;
  assign new_n24613 = new_n24612 ^ new_n24127;
  assign new_n24614 = new_n24136 & new_n24219;
  assign new_n24615 = new_n24614 ^ new_n24540;
  assign new_n24616 = new_n24615 ^ new_n24228;
  assign new_n24617 = new_n24616 ^ new_n8353;
  assign new_n24618 = new_n24617 ^ new_n24613;
  assign new_n24619 = new_n24387 ^ new_n24384;
  assign new_n24620 = new_n24497 ^ new_n23783;
  assign new_n24621 = new_n24620 ^ new_n24601;
  assign new_n24622 = new_n24621 ^ new_n24619;
  assign new_n24623 = new_n24622 ^ new_n24582;
  assign new_n24624 = new_n24288 ^ new_n24266;
  assign new_n24625 = new_n24364 & new_n24624;
  assign new_n24626 = new_n24625 ^ new_n24545;
  assign new_n24627 = new_n24626 ^ new_n24371;
  assign new_n24628 = new_n24627 ^ new_n24569;
  assign new_n24629 = new_n24628 ^ new_n24623;
  assign new_n24630 = new_n24629 ^ new_n24618;
  assign new_n24631 = new_n24630 ^ new_n24552;
  assign new_n24632 = new_n24631 ^ new_n24609;
  assign new_n24633 = ~new_n24608 & ~new_n24632;
  assign new_n24634 = new_n24633 ^ new_n24458;
  assign new_n24635 = new_n24634 ^ new_n24534;
  assign new_n24636 = new_n24634 ^ new_n24608;
  assign new_n24637 = new_n24608 ^ new_n24502;
  assign new_n24638 = new_n24606 ^ new_n24503;
  assign new_n24639 = new_n24638 ^ new_n24631;
  assign new_n24640 = new_n24637 & new_n24639;
  assign new_n24641 = new_n24630 ^ new_n24607;
  assign new_n24642 = new_n24641 ^ new_n24458;
  assign new_n24643 = new_n24553 & new_n24642;
  assign new_n24644 = new_n24643 ^ new_n24640;
  assign new_n24645 = new_n24531 ^ new_n24376;
  assign new_n24646 = new_n24645 ^ new_n24631;
  assign new_n24647 = new_n24630 ^ new_n24531;
  assign new_n24648 = ~new_n24646 & new_n24647;
  assign new_n24649 = new_n24648 ^ new_n24630;
  assign new_n24650 = new_n24649 ^ new_n24644;
  assign new_n24651 = new_n24650 ^ new_n24636;
  assign new_n24652 = new_n24503 & new_n24606;
  assign new_n24653 = new_n24652 ^ new_n24606;
  assign new_n24654 = new_n24641 ^ new_n24376;
  assign new_n24655 = new_n24606 ^ new_n24552;
  assign new_n24656 = ~new_n24655 & new_n24654;
  assign new_n24657 = new_n24656 ^ new_n24653;
  assign new_n24658 = new_n24657 ^ new_n24631;
  assign new_n24659 = new_n24648 ^ new_n24643;
  assign new_n24660 = new_n24578 ^ new_n24376;
  assign new_n24661 = new_n24660 ^ new_n24659;
  assign new_n24662 = new_n24661 ^ new_n24658;
  assign new_n24663 = ~new_n24662 & new_n24651;
  assign new_n24664 = new_n24663 ^ new_n24635;
  assign new_n24665 = new_n24608 ^ new_n24459;
  assign new_n24666 = ~new_n24665 & new_n24631;
  assign new_n24667 = new_n24666 ^ new_n24643;
  assign new_n24668 = new_n24667 ^ new_n24654;
  assign new_n24669 = new_n24668 ^ new_n24664;
  assign new_n24670 = new_n24552 ^ new_n24503;
  assign new_n24671 = new_n24642 ^ new_n24502;
  assign new_n24672 = ~new_n24670 & ~new_n24671;
  assign new_n24673 = new_n24672 ^ new_n24652;
  assign new_n24674 = new_n24666 ^ new_n24648;
  assign new_n24675 = new_n24674 ^ new_n24673;
  assign new_n24676 = ~new_n24669 & ~new_n24675;
  assign new_n24677 = new_n24672 ^ new_n24656;
  assign new_n24678 = new_n24677 ^ new_n24552;
  assign new_n24679 = new_n24678 ^ new_n24668;
  assign new_n24680 = new_n24679 ^ new_n24676;
  assign new_n24681 = ~new_n24532 & new_n24680;
  assign new_n24682 = new_n24606 ^ new_n24376;
  assign new_n24683 = new_n24653 ^ new_n24640;
  assign new_n24684 = new_n24676 ^ new_n24663;
  assign new_n24685 = ~new_n24679 & ~new_n24684;
  assign new_n24686 = new_n24685 ^ new_n24676;
  assign new_n24687 = new_n24679 ^ new_n24663;
  assign new_n24688 = new_n24552 ^ new_n24376;
  assign new_n24689 = new_n24640 ^ new_n24533;
  assign new_n24690 = new_n24689 ^ new_n24674;
  assign new_n24691 = new_n24690 ^ new_n24688;
  assign new_n24692 = ~new_n24691 & new_n24687;
  assign new_n24693 = new_n24692 ^ new_n24635;
  assign new_n24694 = new_n24693 ^ new_n24668;
  assign new_n24695 = ~new_n24686 & ~new_n24694;
  assign new_n24696 = new_n24687 ^ new_n24686;
  assign new_n24697 = new_n24696 ^ new_n24695;
  assign new_n24698 = new_n24697 ^ new_n24683;
  assign new_n24699 = new_n24698 ^ new_n24682;
  assign new_n24700 = new_n24699 ^ new_n24531;
  assign new_n24701 = new_n24692 ^ new_n24656;
  assign new_n24702 = new_n24701 ^ new_n24634;
  assign new_n24703 = new_n24702 ^ new_n24700;
  assign new_n24704 = ~new_n24646 & new_n24703;
  assign new_n24705 = new_n24695 ^ new_n24692;
  assign new_n24706 = new_n24705 ^ new_n24651;
  assign new_n24707 = new_n24654 & new_n24706;
  assign new_n24708 = new_n24696 ^ new_n24676;
  assign new_n24709 = new_n24708 ^ new_n24675;
  assign new_n24710 = new_n24639 & new_n24709;
  assign new_n24711 = new_n24647 & new_n24703;
  assign new_n24712 = new_n24692 ^ new_n24676;
  assign new_n24713 = new_n24678 ^ new_n24635;
  assign new_n24714 = new_n24713 ^ new_n24712;
  assign new_n24715 = ~new_n24714 & new_n24553;
  assign new_n24716 = new_n24715 ^ new_n24711;
  assign new_n24717 = new_n24716 ^ new_n24710;
  assign new_n24718 = new_n24695 ^ new_n24691;
  assign new_n24719 = ~new_n24503 & ~new_n24718;
  assign new_n24720 = new_n24719 ^ new_n24717;
  assign new_n24721 = new_n24720 ^ new_n24707;
  assign new_n24722 = new_n24721 ^ new_n24704;
  assign new_n24723 = new_n24722 ^ new_n24681;
  assign new_n24724 = ~new_n24670 & ~new_n24694;
  assign new_n24725 = new_n24676 ^ new_n24552;
  assign new_n24726 = new_n24672 ^ new_n24533;
  assign new_n24727 = new_n24726 ^ new_n24699;
  assign new_n24728 = new_n24727 ^ new_n24725;
  assign new_n24729 = ~new_n24665 & ~new_n24728;
  assign new_n24730 = new_n24729 ^ new_n24724;
  assign new_n24731 = ~new_n24502 & new_n24680;
  assign new_n24732 = new_n24696 ^ new_n24662;
  assign new_n24733 = ~new_n24608 & new_n24732;
  assign new_n24734 = new_n24733 ^ new_n24731;
  assign new_n24735 = ~new_n24655 & new_n24706;
  assign new_n24736 = new_n24735 ^ new_n24734;
  assign new_n24737 = new_n24736 ^ new_n24730;
  assign new_n24738 = new_n24737 ^ new_n24723;
  assign new_n24739 = new_n24738 ^ new_n23663;
  assign new_n24740 = new_n24739 ^ new_n22574;
  assign new_n24741 = new_n22857 ^ new_n22851;
  assign new_n24742 = new_n24741 ^ new_n22869;
  assign new_n24743 = new_n24742 ^ new_n22874;
  assign new_n24744 = new_n22842 ^ new_n22837;
  assign new_n24745 = new_n24744 ^ new_n24741;
  assign new_n24746 = new_n22851 ^ new_n22842;
  assign new_n24747 = new_n22869 ^ new_n22837;
  assign new_n24748 = new_n24747 ^ new_n24746;
  assign new_n24749 = new_n24745 & new_n24748;
  assign new_n24750 = new_n24749 ^ new_n22874;
  assign new_n24751 = new_n22882 ^ new_n22874;
  assign new_n24752 = ~new_n24751 & new_n22863;
  assign new_n24753 = ~new_n22863 & new_n22842;
  assign new_n24754 = new_n24753 ^ new_n24752;
  assign new_n24755 = new_n24754 ^ new_n24750;
  assign new_n24756 = new_n24751 ^ new_n22863;
  assign new_n24757 = ~new_n22851 & ~new_n24756;
  assign new_n24758 = new_n24757 ^ new_n22851;
  assign new_n24759 = new_n24742 ^ new_n22882;
  assign new_n24760 = new_n22851 ^ new_n22837;
  assign new_n24761 = new_n24759 & new_n24760;
  assign new_n24762 = new_n24761 ^ new_n24758;
  assign new_n24763 = new_n24762 ^ new_n24747;
  assign new_n24764 = new_n24743 & new_n24744;
  assign new_n24765 = new_n22882 ^ new_n22842;
  assign new_n24766 = new_n24765 ^ new_n24747;
  assign new_n24767 = new_n22869 ^ new_n22842;
  assign new_n24768 = new_n24766 & new_n24767;
  assign new_n24769 = new_n24768 ^ new_n24764;
  assign new_n24770 = new_n22882 ^ new_n22857;
  assign new_n24771 = new_n24770 ^ new_n24769;
  assign new_n24772 = new_n24771 ^ new_n24763;
  assign new_n24773 = new_n24750 ^ new_n24745;
  assign new_n24774 = new_n24745 ^ new_n22863;
  assign new_n24775 = new_n24756 ^ new_n22851;
  assign new_n24776 = new_n24775 ^ new_n24747;
  assign new_n24777 = new_n24774 & new_n24776;
  assign new_n24778 = new_n24777 ^ new_n22869;
  assign new_n24779 = new_n24778 ^ new_n24769;
  assign new_n24780 = new_n24779 ^ new_n24773;
  assign new_n24781 = ~new_n24772 & new_n24780;
  assign new_n24782 = new_n24781 ^ new_n24755;
  assign new_n24783 = new_n24751 ^ new_n24745;
  assign new_n24784 = new_n24747 & new_n24783;
  assign new_n24785 = new_n24784 ^ new_n24764;
  assign new_n24786 = new_n24785 ^ new_n24759;
  assign new_n24787 = new_n24786 ^ new_n24782;
  assign new_n24788 = new_n24743 ^ new_n22863;
  assign new_n24789 = new_n24756 ^ new_n22837;
  assign new_n24790 = new_n24788 & new_n24789;
  assign new_n24791 = new_n24790 ^ new_n24757;
  assign new_n24792 = new_n24784 ^ new_n24768;
  assign new_n24793 = new_n24792 ^ new_n24791;
  assign new_n24794 = ~new_n24793 & new_n24787;
  assign new_n24795 = new_n22882 ^ new_n22837;
  assign new_n24796 = new_n24754 ^ new_n22842;
  assign new_n24797 = new_n24796 ^ new_n24777;
  assign new_n24798 = new_n24797 ^ new_n24792;
  assign new_n24799 = new_n24798 ^ new_n24795;
  assign new_n24800 = new_n24790 ^ new_n24761;
  assign new_n24801 = new_n24800 ^ new_n22837;
  assign new_n24802 = new_n24801 ^ new_n24786;
  assign new_n24803 = new_n24802 ^ new_n24781;
  assign new_n24804 = new_n24799 & new_n24803;
  assign new_n24805 = new_n24804 ^ new_n24794;
  assign new_n24806 = new_n24801 ^ new_n24755;
  assign new_n24807 = new_n24806 ^ new_n24805;
  assign new_n24808 = new_n24743 & new_n24807;
  assign new_n24809 = new_n22882 ^ new_n22851;
  assign new_n24810 = new_n24777 ^ new_n24758;
  assign new_n24811 = new_n24804 ^ new_n24755;
  assign new_n24812 = new_n24811 ^ new_n24786;
  assign new_n24813 = new_n24794 ^ new_n24781;
  assign new_n24814 = new_n24802 & new_n24813;
  assign new_n24815 = new_n24814 ^ new_n24803;
  assign new_n24816 = new_n24812 & new_n24815;
  assign new_n24817 = new_n24816 ^ new_n24814;
  assign new_n24818 = new_n24817 ^ new_n24810;
  assign new_n24819 = new_n24818 ^ new_n24809;
  assign new_n24820 = new_n24819 ^ new_n22842;
  assign new_n24821 = new_n24804 ^ new_n24761;
  assign new_n24822 = new_n24821 ^ new_n24750;
  assign new_n24823 = new_n24822 ^ new_n24820;
  assign new_n24824 = ~new_n24823 & new_n24766;
  assign new_n24825 = new_n24824 ^ new_n24808;
  assign new_n24826 = new_n24814 ^ new_n24794;
  assign new_n24827 = new_n24826 ^ new_n24793;
  assign new_n24828 = ~new_n24827 & new_n24774;
  assign new_n24829 = new_n24814 ^ new_n24772;
  assign new_n24830 = ~new_n24829 & new_n24745;
  assign new_n24831 = new_n24830 ^ new_n24828;
  assign new_n24832 = ~new_n24829 & new_n24748;
  assign new_n24833 = new_n24832 ^ new_n24831;
  assign new_n24834 = ~new_n24827 & new_n24776;
  assign new_n24835 = ~new_n24823 & new_n24767;
  assign new_n24836 = new_n24744 & new_n24807;
  assign new_n24837 = new_n24836 ^ new_n24835;
  assign new_n24838 = new_n24837 ^ new_n24834;
  assign new_n24839 = new_n24838 ^ new_n24833;
  assign new_n24840 = new_n24839 ^ new_n24825;
  assign new_n24841 = new_n24840 ^ new_n10193;
  assign new_n24842 = new_n24836 ^ new_n24808;
  assign new_n24843 = new_n24794 ^ new_n22837;
  assign new_n24844 = new_n24796 ^ new_n24790;
  assign new_n24845 = new_n24844 ^ new_n24819;
  assign new_n24846 = new_n24845 ^ new_n24843;
  assign new_n24847 = ~new_n24846 & new_n24747;
  assign new_n24848 = new_n24789 & new_n24812;
  assign new_n24849 = ~new_n24846 & new_n24783;
  assign new_n24850 = new_n24849 ^ new_n24848;
  assign new_n24851 = new_n24802 ^ new_n24794;
  assign new_n24852 = new_n22863 & new_n24851;
  assign new_n24853 = new_n24852 ^ new_n24830;
  assign new_n24854 = new_n24816 ^ new_n24804;
  assign new_n24855 = new_n24854 ^ new_n24780;
  assign new_n24856 = new_n24760 & new_n24855;
  assign new_n24857 = new_n24856 ^ new_n24853;
  assign new_n24858 = new_n24857 ^ new_n24850;
  assign new_n24859 = new_n24858 ^ new_n24847;
  assign new_n24860 = new_n24859 ^ new_n24842;
  assign new_n24861 = new_n24860 ^ new_n10191;
  assign new_n24862 = new_n24861 ^ new_n24841;
  assign new_n24863 = new_n24759 & new_n24855;
  assign new_n24864 = new_n24863 ^ new_n24857;
  assign new_n24865 = new_n24816 ^ new_n24799;
  assign new_n24866 = new_n24775 & new_n24865;
  assign new_n24867 = new_n24788 & new_n24812;
  assign new_n24868 = new_n24867 ^ new_n24866;
  assign new_n24869 = new_n24868 ^ new_n24837;
  assign new_n24870 = new_n24869 ^ new_n24864;
  assign new_n24871 = new_n24870 ^ new_n10189;
  assign new_n24872 = new_n24871 ^ new_n24862;
  assign new_n24873 = new_n24756 & new_n24865;
  assign new_n24874 = new_n24873 ^ new_n24838;
  assign new_n24875 = new_n24874 ^ new_n24863;
  assign new_n24876 = new_n24875 ^ new_n24833;
  assign new_n24877 = new_n24876 ^ new_n10186;
  assign new_n24878 = new_n24877 ^ new_n24872;
  assign new_n24879 = ~new_n24878 & new_n24871;
  assign new_n24880 = new_n24879 ^ new_n24877;
  assign new_n24881 = new_n24867 ^ new_n24832;
  assign new_n24882 = new_n24852 ^ new_n24828;
  assign new_n24883 = new_n24882 ^ new_n24874;
  assign new_n24884 = new_n24883 ^ new_n24881;
  assign new_n24885 = new_n24884 ^ new_n10208;
  assign new_n24886 = new_n24856 ^ new_n24849;
  assign new_n24887 = new_n24873 ^ new_n24824;
  assign new_n24888 = new_n24887 ^ new_n24869;
  assign new_n24889 = new_n24888 ^ new_n24886;
  assign new_n24890 = new_n24889 ^ new_n10201;
  assign new_n24891 = new_n24890 ^ new_n24885;
  assign new_n24892 = new_n24832 ^ new_n24808;
  assign new_n24893 = new_n24875 ^ new_n24824;
  assign new_n24894 = new_n24893 ^ new_n24892;
  assign new_n24895 = new_n24894 ^ new_n10184;
  assign new_n24896 = new_n24895 ^ new_n24877;
  assign new_n24897 = new_n24896 ^ new_n24891;
  assign new_n24898 = new_n24890 ^ new_n24877;
  assign new_n24899 = new_n24756 ^ new_n22842;
  assign new_n24900 = new_n24851 & new_n24899;
  assign new_n24901 = new_n24900 ^ new_n24893;
  assign new_n24902 = new_n24901 ^ new_n24858;
  assign new_n24903 = new_n24902 ^ new_n10204;
  assign new_n24904 = new_n24903 ^ new_n24895;
  assign new_n24905 = new_n24904 ^ new_n24898;
  assign new_n24906 = ~new_n24905 & new_n24897;
  assign new_n24907 = new_n24906 ^ new_n24841;
  assign new_n24908 = new_n24907 ^ new_n24880;
  assign new_n24909 = ~new_n24890 & new_n24872;
  assign new_n24910 = new_n24909 ^ new_n24890;
  assign new_n24911 = new_n24903 ^ new_n24891;
  assign new_n24912 = new_n24911 ^ new_n24861;
  assign new_n24913 = new_n24895 ^ new_n24890;
  assign new_n24914 = ~new_n24912 & new_n24913;
  assign new_n24915 = new_n24914 ^ new_n24910;
  assign new_n24916 = new_n24915 ^ new_n24904;
  assign new_n24917 = new_n24903 ^ new_n24877;
  assign new_n24918 = new_n24895 ^ new_n24861;
  assign new_n24919 = new_n24918 ^ new_n24917;
  assign new_n24920 = ~new_n24917 & ~new_n24919;
  assign new_n24921 = new_n24911 ^ new_n24841;
  assign new_n24922 = new_n24896 & new_n24921;
  assign new_n24923 = new_n24922 ^ new_n24920;
  assign new_n24924 = new_n24885 ^ new_n24861;
  assign new_n24925 = new_n24924 ^ new_n24923;
  assign new_n24926 = new_n24925 ^ new_n24916;
  assign new_n24927 = new_n24907 ^ new_n24897;
  assign new_n24928 = new_n24897 ^ new_n24871;
  assign new_n24929 = new_n24890 ^ new_n24872;
  assign new_n24930 = new_n24929 ^ new_n24904;
  assign new_n24931 = new_n24928 & new_n24930;
  assign new_n24932 = new_n24931 ^ new_n24922;
  assign new_n24933 = new_n24920 ^ new_n24903;
  assign new_n24934 = new_n24933 ^ new_n24932;
  assign new_n24935 = new_n24934 ^ new_n24927;
  assign new_n24936 = new_n24926 & new_n24935;
  assign new_n24937 = new_n24936 ^ new_n24908;
  assign new_n24938 = new_n24897 ^ new_n24862;
  assign new_n24939 = ~new_n24904 & ~new_n24938;
  assign new_n24940 = new_n24939 ^ new_n24922;
  assign new_n24941 = new_n24940 ^ new_n24912;
  assign new_n24942 = new_n24941 ^ new_n24937;
  assign new_n24943 = new_n24895 ^ new_n24872;
  assign new_n24944 = new_n24921 ^ new_n24871;
  assign new_n24945 = ~new_n24943 & new_n24944;
  assign new_n24946 = new_n24945 ^ new_n24909;
  assign new_n24947 = new_n24939 ^ new_n24920;
  assign new_n24948 = new_n24947 ^ new_n24946;
  assign new_n24949 = ~new_n24948 & new_n24942;
  assign new_n24950 = new_n24945 ^ new_n24914;
  assign new_n24951 = new_n24950 ^ new_n24895;
  assign new_n24952 = new_n24951 ^ new_n24941;
  assign new_n24953 = new_n24952 ^ new_n24949;
  assign new_n24954 = ~new_n24878 & ~new_n24953;
  assign new_n24955 = new_n24890 ^ new_n24861;
  assign new_n24956 = new_n24931 ^ new_n24910;
  assign new_n24957 = new_n24949 ^ new_n24936;
  assign new_n24958 = ~new_n24957 & new_n24952;
  assign new_n24959 = new_n24958 ^ new_n24949;
  assign new_n24960 = new_n24952 ^ new_n24936;
  assign new_n24961 = new_n24931 ^ new_n24879;
  assign new_n24962 = new_n24961 ^ new_n24947;
  assign new_n24963 = new_n24962 ^ new_n24918;
  assign new_n24964 = ~new_n24960 & new_n24963;
  assign new_n24965 = new_n24964 ^ new_n24908;
  assign new_n24966 = new_n24965 ^ new_n24941;
  assign new_n24967 = ~new_n24959 & new_n24966;
  assign new_n24968 = new_n24960 ^ new_n24959;
  assign new_n24969 = new_n24968 ^ new_n24967;
  assign new_n24970 = new_n24969 ^ new_n24956;
  assign new_n24971 = new_n24970 ^ new_n24955;
  assign new_n24972 = new_n24971 ^ new_n24877;
  assign new_n24973 = new_n24964 ^ new_n24914;
  assign new_n24974 = new_n24973 ^ new_n24907;
  assign new_n24975 = new_n24974 ^ new_n24972;
  assign new_n24976 = ~new_n24919 & new_n24975;
  assign new_n24977 = new_n24967 ^ new_n24964;
  assign new_n24978 = new_n24977 ^ new_n24935;
  assign new_n24979 = ~new_n24912 & new_n24978;
  assign new_n24980 = new_n24968 ^ new_n24949;
  assign new_n24981 = new_n24980 ^ new_n24948;
  assign new_n24982 = ~new_n24981 & new_n24930;
  assign new_n24983 = new_n24964 ^ new_n24949;
  assign new_n24984 = new_n24951 ^ new_n24908;
  assign new_n24985 = new_n24984 ^ new_n24983;
  assign new_n24986 = ~new_n24985 & new_n24896;
  assign new_n24987 = ~new_n24917 & new_n24975;
  assign new_n24988 = new_n24987 ^ new_n24986;
  assign new_n24989 = new_n24988 ^ new_n24982;
  assign new_n24990 = new_n24967 ^ new_n24963;
  assign new_n24991 = ~new_n24872 & new_n24990;
  assign new_n24992 = new_n24991 ^ new_n24989;
  assign new_n24993 = new_n24992 ^ new_n24979;
  assign new_n24994 = new_n24993 ^ new_n24976;
  assign new_n24995 = new_n24994 ^ new_n24954;
  assign new_n24996 = ~new_n24943 & new_n24966;
  assign new_n24997 = new_n24949 ^ new_n24895;
  assign new_n24998 = new_n24945 ^ new_n24879;
  assign new_n24999 = new_n24998 ^ new_n24971;
  assign new_n25000 = new_n24999 ^ new_n24997;
  assign new_n25001 = ~new_n24938 & ~new_n25000;
  assign new_n25002 = new_n25001 ^ new_n24996;
  assign new_n25003 = ~new_n24953 & new_n24871;
  assign new_n25004 = new_n24968 ^ new_n24926;
  assign new_n25005 = new_n24897 & new_n25004;
  assign new_n25006 = new_n25005 ^ new_n25003;
  assign new_n25007 = new_n24913 & new_n24978;
  assign new_n25008 = new_n25007 ^ new_n25006;
  assign new_n25009 = new_n25008 ^ new_n25002;
  assign new_n25010 = new_n25009 ^ new_n24995;
  assign new_n25011 = new_n25010 ^ new_n23144;
  assign new_n25012 = new_n24840 ^ new_n19032;
  assign new_n25013 = new_n19029 ^ new_n17563;
  assign new_n25014 = new_n25013 ^ new_n9179;
  assign new_n25015 = new_n25014 ^ new_n22064;
  assign new_n25016 = new_n23865 ^ new_n21581;
  assign new_n25017 = new_n25016 ^ new_n25015;
  assign new_n25018 = new_n19834 ^ new_n17524;
  assign new_n25019 = new_n25018 ^ new_n9172;
  assign new_n25020 = new_n25019 ^ new_n22118;
  assign new_n25021 = new_n25020 ^ new_n23824;
  assign new_n25022 = new_n23848 ^ new_n22102;
  assign new_n25023 = new_n25022 ^ new_n25021;
  assign new_n25024 = new_n23844 ^ new_n22028;
  assign new_n25025 = new_n19818 ^ new_n17541;
  assign new_n25026 = new_n25025 ^ new_n9168;
  assign new_n25027 = new_n25026 ^ new_n21971;
  assign new_n25028 = new_n25027 ^ new_n23824;
  assign new_n25029 = new_n25028 ^ new_n25024;
  assign new_n25030 = new_n25029 ^ new_n25023;
  assign new_n25031 = new_n19878 ^ new_n17555;
  assign new_n25032 = new_n25031 ^ new_n9163;
  assign new_n25033 = new_n25032 ^ new_n22004;
  assign new_n25034 = new_n23808 ^ new_n22130;
  assign new_n25035 = new_n25034 ^ new_n25033;
  assign new_n25036 = new_n25035 ^ new_n25030;
  assign new_n25037 = new_n25036 ^ new_n25017;
  assign new_n25038 = new_n19861 ^ new_n17580;
  assign new_n25039 = new_n25038 ^ new_n9184;
  assign new_n25040 = new_n25039 ^ new_n22151;
  assign new_n25041 = new_n23824 ^ new_n21931;
  assign new_n25042 = new_n25041 ^ new_n25040;
  assign new_n25043 = new_n23820 ^ new_n22074;
  assign new_n25044 = new_n19775 ^ new_n17575;
  assign new_n25045 = new_n25044 ^ new_n9190;
  assign new_n25046 = new_n25045 ^ new_n22104;
  assign new_n25047 = new_n25046 ^ new_n23824;
  assign new_n25048 = new_n25047 ^ new_n25043;
  assign new_n25049 = new_n19652 ^ new_n17572;
  assign new_n25050 = new_n25049 ^ new_n9207;
  assign new_n25051 = new_n25050 ^ new_n22085;
  assign new_n25052 = new_n23833 ^ new_n22049;
  assign new_n25053 = new_n25052 ^ new_n25051;
  assign new_n25054 = new_n25053 ^ new_n25017;
  assign new_n25055 = new_n25054 ^ new_n25042;
  assign new_n25056 = new_n25055 ^ new_n25048;
  assign new_n25057 = ~new_n25042 & ~new_n25056;
  assign new_n25058 = new_n25057 ^ new_n25048;
  assign new_n25059 = new_n19731 ^ new_n17567;
  assign new_n25060 = new_n25059 ^ new_n9194;
  assign new_n25061 = new_n25060 ^ new_n21736;
  assign new_n25062 = new_n23856 ^ new_n21907;
  assign new_n25063 = new_n25062 ^ new_n25061;
  assign new_n25064 = new_n25063 ^ new_n25048;
  assign new_n25065 = new_n25064 ^ new_n25030;
  assign new_n25066 = new_n25048 ^ new_n25029;
  assign new_n25067 = new_n25063 ^ new_n25035;
  assign new_n25068 = new_n25067 ^ new_n25066;
  assign new_n25069 = ~new_n25065 & ~new_n25068;
  assign new_n25070 = new_n25069 ^ new_n25017;
  assign new_n25071 = new_n25070 ^ new_n25058;
  assign new_n25072 = new_n25070 ^ new_n25065;
  assign new_n25073 = new_n25037 & new_n25064;
  assign new_n25074 = new_n25055 ^ new_n25029;
  assign new_n25075 = new_n25074 ^ new_n25067;
  assign new_n25076 = new_n25065 ^ new_n25042;
  assign new_n25077 = new_n25075 & new_n25076;
  assign new_n25078 = new_n25077 ^ new_n25073;
  assign new_n25079 = new_n25053 ^ new_n25048;
  assign new_n25080 = new_n25079 ^ new_n25067;
  assign new_n25081 = new_n25048 ^ new_n25035;
  assign new_n25082 = ~new_n25080 & new_n25081;
  assign new_n25083 = new_n25082 ^ new_n25035;
  assign new_n25084 = new_n25083 ^ new_n25078;
  assign new_n25085 = new_n25084 ^ new_n25072;
  assign new_n25086 = new_n25029 & new_n25055;
  assign new_n25087 = new_n25086 ^ new_n25029;
  assign new_n25088 = new_n25053 ^ new_n25036;
  assign new_n25089 = new_n25063 ^ new_n25029;
  assign new_n25090 = ~new_n25089 & new_n25088;
  assign new_n25091 = new_n25090 ^ new_n25087;
  assign new_n25092 = new_n25091 ^ new_n25067;
  assign new_n25093 = new_n25082 ^ new_n25073;
  assign new_n25094 = new_n25053 ^ new_n25023;
  assign new_n25095 = new_n25094 ^ new_n25093;
  assign new_n25096 = new_n25095 ^ new_n25092;
  assign new_n25097 = ~new_n25096 & new_n25085;
  assign new_n25098 = new_n25097 ^ new_n25071;
  assign new_n25099 = new_n25065 ^ new_n25054;
  assign new_n25100 = ~new_n25099 & new_n25067;
  assign new_n25101 = new_n25100 ^ new_n25073;
  assign new_n25102 = new_n25101 ^ new_n25088;
  assign new_n25103 = new_n25102 ^ new_n25098;
  assign new_n25104 = new_n25063 ^ new_n25055;
  assign new_n25105 = new_n25042 ^ new_n25037;
  assign new_n25106 = ~new_n25104 & ~new_n25105;
  assign new_n25107 = new_n25106 ^ new_n25086;
  assign new_n25108 = new_n25100 ^ new_n25082;
  assign new_n25109 = new_n25108 ^ new_n25107;
  assign new_n25110 = ~new_n25103 & ~new_n25109;
  assign new_n25111 = new_n25063 ^ new_n25053;
  assign new_n25112 = new_n25077 ^ new_n25057;
  assign new_n25113 = new_n25112 ^ new_n25108;
  assign new_n25114 = new_n25113 ^ new_n25111;
  assign new_n25115 = new_n25106 ^ new_n25090;
  assign new_n25116 = new_n25115 ^ new_n25063;
  assign new_n25117 = new_n25116 ^ new_n25102;
  assign new_n25118 = new_n25117 ^ new_n25097;
  assign new_n25119 = ~new_n25114 & new_n25118;
  assign new_n25120 = new_n25119 ^ new_n25110;
  assign new_n25121 = new_n25116 ^ new_n25071;
  assign new_n25122 = new_n25121 ^ new_n25120;
  assign new_n25123 = ~new_n25122 & new_n25037;
  assign new_n25124 = new_n25053 ^ new_n25029;
  assign new_n25125 = new_n25087 ^ new_n25077;
  assign new_n25126 = new_n25119 ^ new_n25071;
  assign new_n25127 = new_n25126 ^ new_n25102;
  assign new_n25128 = new_n25110 ^ new_n25097;
  assign new_n25129 = new_n25117 & new_n25128;
  assign new_n25130 = new_n25129 ^ new_n25118;
  assign new_n25131 = ~new_n25127 & new_n25130;
  assign new_n25132 = new_n25131 ^ new_n25129;
  assign new_n25133 = new_n25132 ^ new_n25125;
  assign new_n25134 = new_n25133 ^ new_n25124;
  assign new_n25135 = new_n25134 ^ new_n25048;
  assign new_n25136 = new_n25119 ^ new_n25090;
  assign new_n25137 = new_n25136 ^ new_n25070;
  assign new_n25138 = new_n25137 ^ new_n25135;
  assign new_n25139 = ~new_n25080 & ~new_n25138;
  assign new_n25140 = new_n25139 ^ new_n25123;
  assign new_n25141 = new_n25129 ^ new_n25110;
  assign new_n25142 = new_n25141 ^ new_n25109;
  assign new_n25143 = ~new_n25142 & new_n25076;
  assign new_n25144 = new_n25129 ^ new_n25096;
  assign new_n25145 = ~new_n25065 & ~new_n25144;
  assign new_n25146 = new_n25145 ^ new_n25143;
  assign new_n25147 = ~new_n25068 & ~new_n25144;
  assign new_n25148 = new_n25147 ^ new_n25146;
  assign new_n25149 = ~new_n25142 & new_n25075;
  assign new_n25150 = ~new_n25122 & new_n25064;
  assign new_n25151 = ~new_n25138 & new_n25081;
  assign new_n25152 = new_n25151 ^ new_n25150;
  assign new_n25153 = new_n25152 ^ new_n25149;
  assign new_n25154 = new_n25153 ^ new_n25148;
  assign new_n25155 = new_n25154 ^ new_n25140;
  assign new_n25156 = new_n25155 ^ new_n25012;
  assign new_n25157 = new_n25150 ^ new_n25123;
  assign new_n25158 = new_n25110 ^ new_n25063;
  assign new_n25159 = new_n25106 ^ new_n25057;
  assign new_n25160 = new_n25159 ^ new_n25134;
  assign new_n25161 = new_n25160 ^ new_n25158;
  assign new_n25162 = new_n25067 & new_n25161;
  assign new_n25163 = ~new_n25099 & new_n25161;
  assign new_n25164 = ~new_n25104 & ~new_n25127;
  assign new_n25165 = new_n25164 ^ new_n25163;
  assign new_n25166 = new_n25131 ^ new_n25119;
  assign new_n25167 = new_n25166 ^ new_n25085;
  assign new_n25168 = ~new_n25089 & new_n25167;
  assign new_n25169 = new_n25117 ^ new_n25110;
  assign new_n25170 = ~new_n25042 & new_n25169;
  assign new_n25171 = new_n25170 ^ new_n25145;
  assign new_n25172 = new_n25171 ^ new_n25168;
  assign new_n25173 = new_n25172 ^ new_n25165;
  assign new_n25174 = new_n25173 ^ new_n25162;
  assign new_n25175 = new_n25174 ^ new_n25157;
  assign new_n25176 = new_n25175 ^ new_n25156;
  assign new_n25177 = new_n23029 ^ new_n17414;
  assign new_n25178 = new_n22446 ^ new_n18565;
  assign new_n25179 = new_n25178 ^ new_n18744;
  assign new_n25180 = new_n25179 ^ new_n25177;
  assign new_n25181 = new_n18808 ^ new_n18700;
  assign new_n25182 = new_n25181 ^ new_n18677;
  assign new_n25183 = new_n23992 ^ new_n22471;
  assign new_n25184 = new_n25183 ^ new_n25182;
  assign new_n25185 = new_n18711 ^ new_n18582;
  assign new_n25186 = new_n25185 ^ new_n22983;
  assign new_n25187 = new_n21186 ^ new_n18829;
  assign new_n25188 = new_n25187 ^ new_n18656;
  assign new_n25189 = new_n25188 ^ new_n25186;
  assign new_n25190 = new_n18799 ^ new_n18781;
  assign new_n25191 = new_n25190 ^ new_n18786;
  assign new_n25192 = new_n22983 ^ new_n22392;
  assign new_n25193 = new_n25192 ^ new_n23015;
  assign new_n25194 = new_n25193 ^ new_n25191;
  assign new_n25195 = new_n25194 ^ new_n25189;
  assign new_n25196 = new_n25195 ^ new_n25184;
  assign new_n25197 = new_n25196 ^ new_n25180;
  assign new_n25198 = new_n22361 ^ new_n18582;
  assign new_n25199 = new_n23996 ^ new_n22983;
  assign new_n25200 = new_n25199 ^ new_n25198;
  assign new_n25201 = new_n22986 ^ new_n18758;
  assign new_n25202 = new_n22329 ^ new_n18736;
  assign new_n25203 = new_n25202 ^ new_n18731;
  assign new_n25204 = new_n25203 ^ new_n25201;
  assign new_n25205 = new_n25204 ^ new_n25180;
  assign new_n25206 = new_n25205 ^ new_n25200;
  assign new_n25207 = new_n22983 ^ new_n22416;
  assign new_n25208 = new_n25207 ^ new_n22996;
  assign new_n25209 = new_n18774 ^ new_n18722;
  assign new_n25210 = new_n25209 ^ new_n25208;
  assign new_n25211 = new_n25210 ^ new_n25206;
  assign new_n25212 = ~new_n25200 & ~new_n25211;
  assign new_n25213 = new_n25212 ^ new_n25210;
  assign new_n25214 = new_n23021 ^ new_n22260;
  assign new_n25215 = new_n18589 ^ new_n15309;
  assign new_n25216 = new_n25215 ^ new_n25214;
  assign new_n25217 = new_n25216 ^ new_n25210;
  assign new_n25218 = new_n25217 ^ new_n25195;
  assign new_n25219 = new_n25216 ^ new_n25189;
  assign new_n25220 = new_n25210 ^ new_n25184;
  assign new_n25221 = new_n25220 ^ new_n25219;
  assign new_n25222 = ~new_n25218 & ~new_n25221;
  assign new_n25223 = new_n25222 ^ new_n25180;
  assign new_n25224 = new_n25223 ^ new_n25213;
  assign new_n25225 = new_n25223 ^ new_n25218;
  assign new_n25226 = new_n25197 & new_n25217;
  assign new_n25227 = new_n25218 ^ new_n25200;
  assign new_n25228 = new_n25206 ^ new_n25189;
  assign new_n25229 = new_n25216 ^ new_n25184;
  assign new_n25230 = new_n25229 ^ new_n25228;
  assign new_n25231 = new_n25227 & new_n25230;
  assign new_n25232 = new_n25231 ^ new_n25226;
  assign new_n25233 = new_n25210 ^ new_n25204;
  assign new_n25234 = new_n25233 ^ new_n25229;
  assign new_n25235 = ~new_n25234 & new_n25220;
  assign new_n25236 = new_n25235 ^ new_n25184;
  assign new_n25237 = new_n25236 ^ new_n25232;
  assign new_n25238 = new_n25237 ^ new_n25225;
  assign new_n25239 = new_n25189 & new_n25206;
  assign new_n25240 = new_n25239 ^ new_n25189;
  assign new_n25241 = new_n25204 ^ new_n25196;
  assign new_n25242 = ~new_n25219 & new_n25241;
  assign new_n25243 = new_n25242 ^ new_n25240;
  assign new_n25244 = new_n25243 ^ new_n25229;
  assign new_n25245 = new_n25235 ^ new_n25226;
  assign new_n25246 = new_n25204 ^ new_n25194;
  assign new_n25247 = new_n25246 ^ new_n25245;
  assign new_n25248 = new_n25247 ^ new_n25244;
  assign new_n25249 = ~new_n25248 & new_n25238;
  assign new_n25250 = new_n25249 ^ new_n25224;
  assign new_n25251 = new_n25218 ^ new_n25205;
  assign new_n25252 = ~new_n25251 & new_n25229;
  assign new_n25253 = new_n25252 ^ new_n25226;
  assign new_n25254 = new_n25253 ^ new_n25241;
  assign new_n25255 = new_n25254 ^ new_n25250;
  assign new_n25256 = new_n25216 ^ new_n25206;
  assign new_n25257 = new_n25200 ^ new_n25197;
  assign new_n25258 = ~new_n25256 & ~new_n25257;
  assign new_n25259 = new_n25258 ^ new_n25239;
  assign new_n25260 = new_n25252 ^ new_n25235;
  assign new_n25261 = new_n25260 ^ new_n25259;
  assign new_n25262 = ~new_n25255 & ~new_n25261;
  assign new_n25263 = new_n25216 ^ new_n25204;
  assign new_n25264 = new_n25231 ^ new_n25212;
  assign new_n25265 = new_n25264 ^ new_n25260;
  assign new_n25266 = new_n25265 ^ new_n25263;
  assign new_n25267 = new_n25258 ^ new_n25242;
  assign new_n25268 = new_n25267 ^ new_n25216;
  assign new_n25269 = new_n25268 ^ new_n25254;
  assign new_n25270 = new_n25269 ^ new_n25249;
  assign new_n25271 = ~new_n25266 & new_n25270;
  assign new_n25272 = new_n25271 ^ new_n25262;
  assign new_n25273 = new_n25268 ^ new_n25224;
  assign new_n25274 = new_n25273 ^ new_n25272;
  assign new_n25275 = ~new_n25274 & new_n25197;
  assign new_n25276 = new_n25204 ^ new_n25189;
  assign new_n25277 = new_n25240 ^ new_n25231;
  assign new_n25278 = new_n25271 ^ new_n25224;
  assign new_n25279 = new_n25278 ^ new_n25254;
  assign new_n25280 = new_n25262 ^ new_n25249;
  assign new_n25281 = new_n25269 & new_n25280;
  assign new_n25282 = new_n25281 ^ new_n25270;
  assign new_n25283 = ~new_n25279 & new_n25282;
  assign new_n25284 = new_n25283 ^ new_n25281;
  assign new_n25285 = new_n25284 ^ new_n25277;
  assign new_n25286 = new_n25285 ^ new_n25276;
  assign new_n25287 = new_n25286 ^ new_n25210;
  assign new_n25288 = new_n25271 ^ new_n25242;
  assign new_n25289 = new_n25288 ^ new_n25223;
  assign new_n25290 = new_n25289 ^ new_n25287;
  assign new_n25291 = ~new_n25234 & ~new_n25290;
  assign new_n25292 = new_n25291 ^ new_n25275;
  assign new_n25293 = new_n25281 ^ new_n25262;
  assign new_n25294 = new_n25293 ^ new_n25261;
  assign new_n25295 = ~new_n25294 & new_n25227;
  assign new_n25296 = new_n25281 ^ new_n25248;
  assign new_n25297 = ~new_n25218 & ~new_n25296;
  assign new_n25298 = new_n25297 ^ new_n25295;
  assign new_n25299 = ~new_n25221 & ~new_n25296;
  assign new_n25300 = new_n25299 ^ new_n25298;
  assign new_n25301 = ~new_n25294 & new_n25230;
  assign new_n25302 = ~new_n25290 & new_n25220;
  assign new_n25303 = ~new_n25274 & new_n25217;
  assign new_n25304 = new_n25303 ^ new_n25302;
  assign new_n25305 = new_n25304 ^ new_n25301;
  assign new_n25306 = new_n25305 ^ new_n25300;
  assign new_n25307 = new_n25306 ^ new_n25292;
  assign new_n25308 = new_n22884 ^ new_n20954;
  assign new_n25309 = new_n22580 ^ new_n20881;
  assign new_n25310 = new_n25309 ^ new_n20892;
  assign new_n25311 = new_n25310 ^ new_n25308;
  assign new_n25312 = new_n22578 ^ new_n20771;
  assign new_n25313 = new_n24247 ^ new_n20812;
  assign new_n25314 = new_n25313 ^ new_n25312;
  assign new_n25315 = new_n22575 ^ new_n20820;
  assign new_n25316 = new_n25315 ^ new_n24240;
  assign new_n25317 = new_n22839 ^ new_n20978;
  assign new_n25318 = new_n25317 ^ new_n25316;
  assign new_n25319 = new_n22839 ^ new_n20313;
  assign new_n25320 = new_n22576 ^ new_n20865;
  assign new_n25321 = new_n25320 ^ new_n24276;
  assign new_n25322 = new_n25321 ^ new_n25319;
  assign new_n25323 = new_n25322 ^ new_n25318;
  assign new_n25324 = new_n25323 ^ new_n25314;
  assign new_n25325 = new_n25324 ^ new_n25311;
  assign new_n25326 = new_n22582 ^ new_n20940;
  assign new_n25327 = new_n22839 ^ new_n20841;
  assign new_n25328 = new_n25327 ^ new_n25326;
  assign new_n25329 = new_n22844 ^ new_n20886;
  assign new_n25330 = new_n22583 ^ new_n20915;
  assign new_n25331 = new_n25330 ^ new_n20904;
  assign new_n25332 = new_n25331 ^ new_n25329;
  assign new_n25333 = new_n25332 ^ new_n25311;
  assign new_n25334 = new_n25333 ^ new_n25328;
  assign new_n25335 = new_n24235 ^ new_n22586;
  assign new_n25336 = new_n25335 ^ new_n22839;
  assign new_n25337 = new_n20968 ^ new_n20923;
  assign new_n25338 = new_n25337 ^ new_n25336;
  assign new_n25339 = new_n25338 ^ new_n25334;
  assign new_n25340 = ~new_n25328 & ~new_n25339;
  assign new_n25341 = new_n25340 ^ new_n25338;
  assign new_n25342 = new_n22876 ^ new_n22590;
  assign new_n25343 = new_n24237 ^ new_n20790;
  assign new_n25344 = new_n25343 ^ new_n25342;
  assign new_n25345 = new_n25344 ^ new_n25338;
  assign new_n25346 = new_n25345 ^ new_n25323;
  assign new_n25347 = new_n25338 ^ new_n25322;
  assign new_n25348 = new_n25344 ^ new_n25314;
  assign new_n25349 = new_n25348 ^ new_n25347;
  assign new_n25350 = ~new_n25346 & ~new_n25349;
  assign new_n25351 = new_n25350 ^ new_n25311;
  assign new_n25352 = new_n25351 ^ new_n25341;
  assign new_n25353 = new_n25351 ^ new_n25346;
  assign new_n25354 = new_n25325 & new_n25345;
  assign new_n25355 = new_n25346 ^ new_n25328;
  assign new_n25356 = new_n25334 ^ new_n25322;
  assign new_n25357 = new_n25356 ^ new_n25348;
  assign new_n25358 = new_n25355 & new_n25357;
  assign new_n25359 = new_n25358 ^ new_n25354;
  assign new_n25360 = new_n25338 ^ new_n25314;
  assign new_n25361 = new_n25338 ^ new_n25332;
  assign new_n25362 = new_n25361 ^ new_n25348;
  assign new_n25363 = ~new_n25362 & new_n25360;
  assign new_n25364 = new_n25363 ^ new_n25314;
  assign new_n25365 = new_n25364 ^ new_n25359;
  assign new_n25366 = new_n25365 ^ new_n25353;
  assign new_n25367 = new_n25322 & new_n25334;
  assign new_n25368 = new_n25367 ^ new_n25322;
  assign new_n25369 = new_n25332 ^ new_n25324;
  assign new_n25370 = new_n25344 ^ new_n25322;
  assign new_n25371 = ~new_n25370 & new_n25369;
  assign new_n25372 = new_n25371 ^ new_n25368;
  assign new_n25373 = new_n25372 ^ new_n25348;
  assign new_n25374 = new_n25363 ^ new_n25354;
  assign new_n25375 = new_n25332 ^ new_n25318;
  assign new_n25376 = new_n25375 ^ new_n25374;
  assign new_n25377 = new_n25376 ^ new_n25373;
  assign new_n25378 = ~new_n25377 & new_n25366;
  assign new_n25379 = new_n25378 ^ new_n25352;
  assign new_n25380 = new_n25346 ^ new_n25333;
  assign new_n25381 = ~new_n25380 & new_n25348;
  assign new_n25382 = new_n25381 ^ new_n25354;
  assign new_n25383 = new_n25382 ^ new_n25369;
  assign new_n25384 = new_n25383 ^ new_n25379;
  assign new_n25385 = new_n25344 ^ new_n25334;
  assign new_n25386 = new_n25328 ^ new_n25325;
  assign new_n25387 = ~new_n25385 & ~new_n25386;
  assign new_n25388 = new_n25387 ^ new_n25367;
  assign new_n25389 = new_n25381 ^ new_n25363;
  assign new_n25390 = new_n25389 ^ new_n25388;
  assign new_n25391 = ~new_n25384 & ~new_n25390;
  assign new_n25392 = new_n25344 ^ new_n25332;
  assign new_n25393 = new_n25358 ^ new_n25340;
  assign new_n25394 = new_n25393 ^ new_n25389;
  assign new_n25395 = new_n25394 ^ new_n25392;
  assign new_n25396 = new_n25387 ^ new_n25371;
  assign new_n25397 = new_n25396 ^ new_n25344;
  assign new_n25398 = new_n25397 ^ new_n25383;
  assign new_n25399 = new_n25398 ^ new_n25378;
  assign new_n25400 = ~new_n25395 & new_n25399;
  assign new_n25401 = new_n25400 ^ new_n25391;
  assign new_n25402 = new_n25397 ^ new_n25352;
  assign new_n25403 = new_n25402 ^ new_n25401;
  assign new_n25404 = ~new_n25403 & new_n25325;
  assign new_n25405 = new_n25332 ^ new_n25322;
  assign new_n25406 = new_n25368 ^ new_n25358;
  assign new_n25407 = new_n25400 ^ new_n25352;
  assign new_n25408 = new_n25407 ^ new_n25383;
  assign new_n25409 = new_n25391 ^ new_n25378;
  assign new_n25410 = new_n25398 & new_n25409;
  assign new_n25411 = new_n25410 ^ new_n25399;
  assign new_n25412 = ~new_n25408 & new_n25411;
  assign new_n25413 = new_n25412 ^ new_n25410;
  assign new_n25414 = new_n25413 ^ new_n25406;
  assign new_n25415 = new_n25414 ^ new_n25405;
  assign new_n25416 = new_n25415 ^ new_n25338;
  assign new_n25417 = new_n25400 ^ new_n25371;
  assign new_n25418 = new_n25417 ^ new_n25351;
  assign new_n25419 = new_n25418 ^ new_n25416;
  assign new_n25420 = ~new_n25362 & ~new_n25419;
  assign new_n25421 = new_n25420 ^ new_n25404;
  assign new_n25422 = new_n25410 ^ new_n25391;
  assign new_n25423 = new_n25422 ^ new_n25390;
  assign new_n25424 = ~new_n25423 & new_n25355;
  assign new_n25425 = new_n25410 ^ new_n25377;
  assign new_n25426 = ~new_n25346 & ~new_n25425;
  assign new_n25427 = new_n25426 ^ new_n25424;
  assign new_n25428 = ~new_n25349 & ~new_n25425;
  assign new_n25429 = new_n25428 ^ new_n25427;
  assign new_n25430 = ~new_n25423 & new_n25357;
  assign new_n25431 = ~new_n25403 & new_n25345;
  assign new_n25432 = ~new_n25419 & new_n25360;
  assign new_n25433 = new_n25432 ^ new_n25431;
  assign new_n25434 = new_n25433 ^ new_n25430;
  assign new_n25435 = new_n25434 ^ new_n25429;
  assign new_n25436 = new_n25435 ^ new_n25421;
  assign new_n25437 = new_n25436 ^ new_n25307;
  assign new_n25438 = new_n18793 ^ new_n17711;
  assign new_n25439 = new_n25438 ^ new_n19854;
  assign new_n25440 = new_n19781 ^ new_n19740;
  assign new_n25441 = new_n25440 ^ new_n25439;
  assign new_n25442 = new_n19848 ^ new_n19765;
  assign new_n25443 = new_n25442 ^ new_n19882;
  assign new_n25444 = new_n25443 ^ new_n25441;
  assign new_n25445 = new_n19864 ^ new_n19809;
  assign new_n25446 = new_n25445 ^ new_n25440;
  assign new_n25447 = new_n18634 ^ new_n17705;
  assign new_n25448 = new_n25447 ^ new_n19887;
  assign new_n25449 = new_n25448 ^ new_n19790;
  assign new_n25450 = new_n25449 ^ new_n25446;
  assign new_n25451 = new_n25450 ^ new_n25444;
  assign new_n25452 = new_n19892 ^ new_n19827;
  assign new_n25453 = new_n18670 ^ new_n17719;
  assign new_n25454 = new_n25453 ^ new_n19848;
  assign new_n25455 = new_n25454 ^ new_n19887;
  assign new_n25456 = new_n25455 ^ new_n25452;
  assign new_n25457 = new_n25456 ^ new_n25451;
  assign new_n25458 = new_n19672 ^ new_n19631;
  assign new_n25459 = new_n18765 ^ new_n17692;
  assign new_n25460 = new_n25459 ^ new_n19745;
  assign new_n25461 = new_n25460 ^ new_n19325;
  assign new_n25462 = new_n25461 ^ new_n25458;
  assign new_n25463 = new_n25462 ^ new_n25457;
  assign new_n25464 = new_n19758 ^ new_n19171;
  assign new_n25465 = new_n17726 ^ new_n17678;
  assign new_n25466 = new_n25465 ^ new_n19781;
  assign new_n25467 = new_n25466 ^ new_n19745;
  assign new_n25468 = new_n25467 ^ new_n25464;
  assign new_n25469 = new_n18771 ^ new_n17681;
  assign new_n25470 = new_n25469 ^ new_n19773;
  assign new_n25471 = new_n25470 ^ new_n25440;
  assign new_n25472 = new_n19765 ^ new_n19693;
  assign new_n25473 = new_n25472 ^ new_n19839;
  assign new_n25474 = new_n25473 ^ new_n25471;
  assign new_n25475 = new_n25474 ^ new_n25468;
  assign new_n25476 = new_n25475 ^ new_n25451;
  assign new_n25477 = new_n25474 ^ new_n25450;
  assign new_n25478 = new_n25468 ^ new_n25456;
  assign new_n25479 = new_n25478 ^ new_n25477;
  assign new_n25480 = ~new_n25479 & new_n25476;
  assign new_n25481 = new_n25480 ^ new_n25462;
  assign new_n25482 = new_n18823 ^ new_n17697;
  assign new_n25483 = new_n25482 ^ new_n19790;
  assign new_n25484 = new_n25440 ^ new_n19868;
  assign new_n25485 = new_n25484 ^ new_n25483;
  assign new_n25486 = new_n18718 ^ new_n17688;
  assign new_n25487 = new_n19777 ^ new_n19693;
  assign new_n25488 = new_n25487 ^ new_n25486;
  assign new_n25489 = new_n19720 ^ new_n19325;
  assign new_n25490 = new_n25489 ^ new_n25488;
  assign new_n25491 = new_n25490 ^ new_n25462;
  assign new_n25492 = new_n25485 & new_n25491;
  assign new_n25493 = ~new_n25485 & new_n25474;
  assign new_n25494 = new_n25493 ^ new_n25492;
  assign new_n25495 = new_n25494 ^ new_n25481;
  assign new_n25496 = new_n25481 ^ new_n25476;
  assign new_n25497 = new_n25463 & new_n25475;
  assign new_n25498 = new_n25491 ^ new_n25485;
  assign new_n25499 = new_n25498 ^ new_n25450;
  assign new_n25500 = new_n25499 ^ new_n25478;
  assign new_n25501 = new_n25485 ^ new_n25476;
  assign new_n25502 = new_n25500 & new_n25501;
  assign new_n25503 = new_n25502 ^ new_n25497;
  assign new_n25504 = new_n25490 ^ new_n25474;
  assign new_n25505 = new_n25504 ^ new_n25478;
  assign new_n25506 = new_n25474 ^ new_n25456;
  assign new_n25507 = ~new_n25505 & new_n25506;
  assign new_n25508 = new_n25507 ^ new_n25456;
  assign new_n25509 = new_n25508 ^ new_n25503;
  assign new_n25510 = new_n25509 ^ new_n25496;
  assign new_n25511 = new_n25450 & new_n25498;
  assign new_n25512 = new_n25511 ^ new_n25450;
  assign new_n25513 = new_n25468 ^ new_n25450;
  assign new_n25514 = new_n25490 ^ new_n25457;
  assign new_n25515 = ~new_n25513 & ~new_n25514;
  assign new_n25516 = new_n25515 ^ new_n25512;
  assign new_n25517 = new_n25516 ^ new_n25478;
  assign new_n25518 = new_n25507 ^ new_n25497;
  assign new_n25519 = new_n25490 ^ new_n25444;
  assign new_n25520 = new_n25519 ^ new_n25518;
  assign new_n25521 = new_n25520 ^ new_n25517;
  assign new_n25522 = new_n25510 & new_n25521;
  assign new_n25523 = new_n25522 ^ new_n25495;
  assign new_n25524 = new_n25491 ^ new_n25476;
  assign new_n25525 = ~new_n25524 & new_n25478;
  assign new_n25526 = new_n25525 ^ new_n25497;
  assign new_n25527 = new_n25526 ^ new_n25514;
  assign new_n25528 = new_n25527 ^ new_n25523;
  assign new_n25529 = new_n25498 ^ new_n25468;
  assign new_n25530 = new_n25485 ^ new_n25463;
  assign new_n25531 = ~new_n25529 & new_n25530;
  assign new_n25532 = new_n25531 ^ new_n25511;
  assign new_n25533 = new_n25525 ^ new_n25507;
  assign new_n25534 = new_n25533 ^ new_n25532;
  assign new_n25535 = ~new_n25528 & ~new_n25534;
  assign new_n25536 = new_n25490 ^ new_n25468;
  assign new_n25537 = new_n25494 ^ new_n25474;
  assign new_n25538 = new_n25537 ^ new_n25502;
  assign new_n25539 = new_n25538 ^ new_n25533;
  assign new_n25540 = new_n25539 ^ new_n25536;
  assign new_n25541 = new_n25531 ^ new_n25515;
  assign new_n25542 = new_n25541 ^ new_n25468;
  assign new_n25543 = new_n25542 ^ new_n25527;
  assign new_n25544 = new_n25543 ^ new_n25522;
  assign new_n25545 = ~new_n25540 & ~new_n25544;
  assign new_n25546 = new_n25545 ^ new_n25535;
  assign new_n25547 = new_n25542 ^ new_n25495;
  assign new_n25548 = new_n25547 ^ new_n25546;
  assign new_n25549 = new_n25463 & new_n25548;
  assign new_n25550 = new_n25475 & new_n25548;
  assign new_n25551 = new_n25550 ^ new_n25549;
  assign new_n25552 = new_n25535 ^ new_n25468;
  assign new_n25553 = new_n25537 ^ new_n25531;
  assign new_n25554 = new_n25490 ^ new_n25450;
  assign new_n25555 = new_n25512 ^ new_n25502;
  assign new_n25556 = new_n25545 ^ new_n25495;
  assign new_n25557 = new_n25556 ^ new_n25527;
  assign new_n25558 = new_n25535 ^ new_n25522;
  assign new_n25559 = ~new_n25543 & new_n25558;
  assign new_n25560 = new_n25559 ^ new_n25544;
  assign new_n25561 = ~new_n25557 & ~new_n25560;
  assign new_n25562 = new_n25561 ^ new_n25559;
  assign new_n25563 = new_n25562 ^ new_n25555;
  assign new_n25564 = new_n25563 ^ new_n25554;
  assign new_n25565 = new_n25564 ^ new_n25553;
  assign new_n25566 = new_n25565 ^ new_n25552;
  assign new_n25567 = new_n25478 & new_n25566;
  assign new_n25568 = new_n25561 ^ new_n25545;
  assign new_n25569 = new_n25568 ^ new_n25510;
  assign new_n25570 = ~new_n25513 & new_n25569;
  assign new_n25571 = new_n25559 ^ new_n25521;
  assign new_n25572 = new_n25476 & new_n25571;
  assign new_n25573 = new_n25543 ^ new_n25535;
  assign new_n25574 = ~new_n25573 & new_n25485;
  assign new_n25575 = new_n25574 ^ new_n25572;
  assign new_n25576 = new_n25575 ^ new_n25570;
  assign new_n25577 = ~new_n25524 & new_n25566;
  assign new_n25578 = ~new_n25529 & ~new_n25557;
  assign new_n25579 = new_n25578 ^ new_n25577;
  assign new_n25580 = new_n25579 ^ new_n25576;
  assign new_n25581 = new_n25580 ^ new_n25567;
  assign new_n25582 = new_n25581 ^ new_n25551;
  assign new_n25583 = new_n25582 ^ new_n25437;
  assign new_n25584 = new_n25583 ^ new_n25176;
  assign new_n25585 = new_n25431 ^ new_n25404;
  assign new_n25586 = new_n25391 ^ new_n25344;
  assign new_n25587 = new_n25387 ^ new_n25340;
  assign new_n25588 = new_n25587 ^ new_n25415;
  assign new_n25589 = new_n25588 ^ new_n25586;
  assign new_n25590 = new_n25348 & new_n25589;
  assign new_n25591 = ~new_n25385 & ~new_n25408;
  assign new_n25592 = ~new_n25380 & new_n25589;
  assign new_n25593 = new_n25592 ^ new_n25591;
  assign new_n25594 = new_n25412 ^ new_n25400;
  assign new_n25595 = new_n25594 ^ new_n25366;
  assign new_n25596 = ~new_n25370 & new_n25595;
  assign new_n25597 = new_n25398 ^ new_n25391;
  assign new_n25598 = ~new_n25328 & new_n25597;
  assign new_n25599 = new_n25598 ^ new_n25426;
  assign new_n25600 = new_n25599 ^ new_n25596;
  assign new_n25601 = new_n25600 ^ new_n25593;
  assign new_n25602 = new_n25601 ^ new_n25590;
  assign new_n25603 = new_n25602 ^ new_n25585;
  assign new_n25604 = new_n25303 ^ new_n25275;
  assign new_n25605 = new_n25262 ^ new_n25216;
  assign new_n25606 = new_n25258 ^ new_n25212;
  assign new_n25607 = new_n25606 ^ new_n25286;
  assign new_n25608 = new_n25607 ^ new_n25605;
  assign new_n25609 = new_n25229 & new_n25608;
  assign new_n25610 = ~new_n25256 & ~new_n25279;
  assign new_n25611 = ~new_n25251 & new_n25608;
  assign new_n25612 = new_n25611 ^ new_n25610;
  assign new_n25613 = new_n25283 ^ new_n25271;
  assign new_n25614 = new_n25613 ^ new_n25238;
  assign new_n25615 = ~new_n25219 & new_n25614;
  assign new_n25616 = new_n25269 ^ new_n25262;
  assign new_n25617 = ~new_n25200 & new_n25616;
  assign new_n25618 = new_n25617 ^ new_n25297;
  assign new_n25619 = new_n25618 ^ new_n25615;
  assign new_n25620 = new_n25619 ^ new_n25612;
  assign new_n25621 = new_n25620 ^ new_n25609;
  assign new_n25622 = new_n25621 ^ new_n25604;
  assign new_n25623 = new_n25622 ^ new_n25603;
  assign new_n25624 = new_n25623 ^ new_n25175;
  assign new_n25625 = new_n24860 ^ new_n19062;
  assign new_n25626 = new_n25559 ^ new_n25535;
  assign new_n25627 = new_n25626 ^ new_n25534;
  assign new_n25628 = ~new_n25627 & new_n25501;
  assign new_n25629 = new_n25628 ^ new_n25572;
  assign new_n25630 = ~new_n25479 & new_n25571;
  assign new_n25631 = new_n25630 ^ new_n25629;
  assign new_n25632 = ~new_n25514 & new_n25569;
  assign new_n25633 = ~new_n25627 & new_n25500;
  assign new_n25634 = new_n25564 ^ new_n25474;
  assign new_n25635 = new_n25545 ^ new_n25515;
  assign new_n25636 = new_n25635 ^ new_n25481;
  assign new_n25637 = new_n25636 ^ new_n25634;
  assign new_n25638 = new_n25506 & new_n25637;
  assign new_n25639 = new_n25638 ^ new_n25550;
  assign new_n25640 = new_n25639 ^ new_n25633;
  assign new_n25641 = new_n25561 ^ new_n25540;
  assign new_n25642 = ~new_n25498 & ~new_n25641;
  assign new_n25643 = new_n25642 ^ new_n25640;
  assign new_n25644 = new_n25643 ^ new_n25632;
  assign new_n25645 = new_n25644 ^ new_n25631;
  assign new_n25646 = new_n25131 ^ new_n25114;
  assign new_n25647 = ~new_n25055 & ~new_n25646;
  assign new_n25648 = new_n25647 ^ new_n25153;
  assign new_n25649 = new_n25088 & new_n25167;
  assign new_n25650 = new_n25649 ^ new_n25648;
  assign new_n25651 = new_n25650 ^ new_n25148;
  assign new_n25652 = new_n25651 ^ new_n25645;
  assign new_n25653 = new_n25652 ^ new_n25625;
  assign new_n25654 = new_n25653 ^ new_n25624;
  assign new_n25655 = new_n25654 ^ new_n25584;
  assign new_n25656 = new_n25428 ^ new_n25404;
  assign new_n25657 = new_n25412 ^ new_n25395;
  assign new_n25658 = ~new_n25334 & ~new_n25657;
  assign new_n25659 = new_n25658 ^ new_n25434;
  assign new_n25660 = new_n25369 & new_n25595;
  assign new_n25661 = new_n25660 ^ new_n25659;
  assign new_n25662 = new_n25661 ^ new_n25420;
  assign new_n25663 = new_n25662 ^ new_n25656;
  assign new_n25664 = new_n25299 ^ new_n25275;
  assign new_n25665 = new_n25283 ^ new_n25266;
  assign new_n25666 = ~new_n25206 & ~new_n25665;
  assign new_n25667 = new_n25666 ^ new_n25305;
  assign new_n25668 = new_n25241 & new_n25614;
  assign new_n25669 = new_n25668 ^ new_n25667;
  assign new_n25670 = new_n25669 ^ new_n25291;
  assign new_n25671 = new_n25670 ^ new_n25664;
  assign new_n25672 = new_n25671 ^ new_n25663;
  assign new_n25673 = ~new_n25505 & new_n25637;
  assign new_n25674 = new_n25673 ^ new_n25549;
  assign new_n25675 = new_n25640 ^ new_n25631;
  assign new_n25676 = new_n25675 ^ new_n25674;
  assign new_n25677 = new_n25676 ^ new_n25672;
  assign new_n25678 = new_n24894 ^ new_n19078;
  assign new_n25679 = new_n25147 ^ new_n25123;
  assign new_n25680 = new_n25650 ^ new_n25139;
  assign new_n25681 = new_n25680 ^ new_n25679;
  assign new_n25682 = new_n25681 ^ new_n25678;
  assign new_n25683 = new_n25682 ^ new_n25155;
  assign new_n25684 = new_n25683 ^ new_n25677;
  assign new_n25685 = new_n24876 ^ new_n19068;
  assign new_n25686 = new_n25661 ^ new_n25429;
  assign new_n25687 = new_n25669 ^ new_n25300;
  assign new_n25688 = new_n25687 ^ new_n25686;
  assign new_n25689 = new_n25688 ^ new_n25685;
  assign new_n25690 = new_n25630 ^ new_n25549;
  assign new_n25691 = new_n25673 ^ new_n25644;
  assign new_n25692 = new_n25691 ^ new_n25690;
  assign new_n25693 = new_n25692 ^ new_n25681;
  assign new_n25694 = new_n25693 ^ new_n25689;
  assign new_n25695 = ~new_n25105 & ~new_n25127;
  assign new_n25696 = new_n25695 ^ new_n25147;
  assign new_n25697 = new_n25170 ^ new_n25143;
  assign new_n25698 = new_n25697 ^ new_n25648;
  assign new_n25699 = new_n25698 ^ new_n25696;
  assign new_n25700 = new_n25699 ^ new_n25651;
  assign new_n25701 = ~new_n25557 & new_n25530;
  assign new_n25702 = new_n25701 ^ new_n25630;
  assign new_n25703 = new_n25628 ^ new_n25574;
  assign new_n25704 = new_n25703 ^ new_n25643;
  assign new_n25705 = new_n25704 ^ new_n25702;
  assign new_n25706 = new_n25705 ^ new_n25700;
  assign new_n25707 = new_n25706 ^ new_n25694;
  assign new_n25708 = new_n25707 ^ new_n25684;
  assign new_n25709 = new_n25615 ^ new_n25611;
  assign new_n25710 = new_n25666 ^ new_n25291;
  assign new_n25711 = ~new_n25665 & new_n25228;
  assign new_n25712 = ~new_n25257 & ~new_n25279;
  assign new_n25713 = new_n25712 ^ new_n25711;
  assign new_n25714 = new_n25713 ^ new_n25304;
  assign new_n25715 = new_n25714 ^ new_n25710;
  assign new_n25716 = new_n25715 ^ new_n25709;
  assign new_n25717 = new_n25596 ^ new_n25592;
  assign new_n25718 = new_n25658 ^ new_n25420;
  assign new_n25719 = ~new_n25657 & new_n25356;
  assign new_n25720 = ~new_n25386 & ~new_n25408;
  assign new_n25721 = new_n25720 ^ new_n25719;
  assign new_n25722 = new_n25721 ^ new_n25433;
  assign new_n25723 = new_n25722 ^ new_n25718;
  assign new_n25724 = new_n25723 ^ new_n25717;
  assign new_n25725 = new_n25724 ^ new_n25716;
  assign new_n25726 = ~new_n25641 & new_n25499;
  assign new_n25727 = new_n25726 ^ new_n25701;
  assign new_n25728 = new_n25727 ^ new_n25639;
  assign new_n25729 = new_n25632 ^ new_n25576;
  assign new_n25730 = new_n25729 ^ new_n25728;
  assign new_n25731 = new_n25730 ^ new_n25725;
  assign new_n25732 = new_n25731 ^ new_n25693;
  assign new_n25733 = new_n25168 ^ new_n25163;
  assign new_n25734 = new_n25647 ^ new_n25139;
  assign new_n25735 = ~new_n25646 & new_n25074;
  assign new_n25736 = new_n25735 ^ new_n25695;
  assign new_n25737 = new_n25736 ^ new_n25152;
  assign new_n25738 = new_n25737 ^ new_n25734;
  assign new_n25739 = new_n25738 ^ new_n25733;
  assign new_n25740 = new_n24889 ^ new_n19044;
  assign new_n25741 = new_n25740 ^ new_n25739;
  assign new_n25742 = new_n25649 ^ new_n25172;
  assign new_n25743 = new_n25742 ^ new_n25737;
  assign new_n25744 = new_n25743 ^ new_n25741;
  assign new_n25745 = new_n25744 ^ new_n25732;
  assign new_n25746 = ~new_n25056 & new_n25169;
  assign new_n25747 = new_n25746 ^ new_n25680;
  assign new_n25748 = new_n25747 ^ new_n25173;
  assign new_n25749 = new_n25748 ^ new_n25699;
  assign new_n25750 = new_n25498 ^ new_n25474;
  assign new_n25751 = ~new_n25573 & ~new_n25750;
  assign new_n25752 = new_n25751 ^ new_n25691;
  assign new_n25753 = new_n25752 ^ new_n25580;
  assign new_n25754 = new_n25753 ^ new_n25749;
  assign new_n25755 = new_n24884 ^ new_n19050;
  assign new_n25756 = new_n25720 ^ new_n25428;
  assign new_n25757 = new_n25598 ^ new_n25424;
  assign new_n25758 = new_n25757 ^ new_n25659;
  assign new_n25759 = new_n25758 ^ new_n25756;
  assign new_n25760 = new_n25712 ^ new_n25299;
  assign new_n25761 = new_n25617 ^ new_n25295;
  assign new_n25762 = new_n25761 ^ new_n25667;
  assign new_n25763 = new_n25762 ^ new_n25760;
  assign new_n25764 = new_n25763 ^ new_n25759;
  assign new_n25765 = new_n25764 ^ new_n25755;
  assign new_n25766 = new_n25765 ^ new_n25693;
  assign new_n25767 = new_n25766 ^ new_n25754;
  assign new_n25768 = new_n25767 ^ new_n25745;
  assign new_n25769 = new_n25768 ^ new_n25708;
  assign new_n25770 = new_n25769 ^ new_n25655;
  assign new_n25771 = new_n24870 ^ new_n19057;
  assign new_n25772 = new_n25771 ^ new_n25743;
  assign new_n25773 = new_n25668 ^ new_n25619;
  assign new_n25774 = new_n25773 ^ new_n25714;
  assign new_n25775 = new_n25660 ^ new_n25600;
  assign new_n25776 = new_n25775 ^ new_n25722;
  assign new_n25777 = new_n25776 ^ new_n25774;
  assign new_n25778 = new_n25777 ^ new_n25693;
  assign new_n25779 = new_n25778 ^ new_n25772;
  assign new_n25780 = new_n25779 ^ new_n25655;
  assign new_n25781 = new_n25780 ^ new_n25707;
  assign new_n25782 = new_n25779 & new_n25781;
  assign new_n25783 = new_n25782 ^ new_n25707;
  assign new_n25784 = ~new_n25339 & new_n25597;
  assign new_n25785 = new_n25784 ^ new_n25662;
  assign new_n25786 = new_n25785 ^ new_n25601;
  assign new_n25787 = ~new_n25211 & new_n25616;
  assign new_n25788 = new_n25787 ^ new_n25670;
  assign new_n25789 = new_n25788 ^ new_n25620;
  assign new_n25790 = new_n25789 ^ new_n25786;
  assign new_n25791 = new_n25577 ^ new_n25570;
  assign new_n25792 = new_n25673 ^ new_n25642;
  assign new_n25793 = new_n25792 ^ new_n25728;
  assign new_n25794 = new_n25793 ^ new_n25791;
  assign new_n25795 = new_n25794 ^ new_n25790;
  assign new_n25796 = new_n24902 ^ new_n19037;
  assign new_n25797 = new_n25796 ^ new_n25748;
  assign new_n25798 = new_n25797 ^ new_n25739;
  assign new_n25799 = new_n25798 ^ new_n25795;
  assign new_n25800 = new_n25799 ^ new_n25707;
  assign new_n25801 = new_n25745 ^ new_n25684;
  assign new_n25802 = new_n25801 ^ new_n25800;
  assign new_n25803 = ~new_n25802 & new_n25769;
  assign new_n25804 = new_n25803 ^ new_n25584;
  assign new_n25805 = new_n25804 ^ new_n25783;
  assign new_n25806 = new_n25745 & new_n25780;
  assign new_n25807 = new_n25806 ^ new_n25745;
  assign new_n25808 = new_n25799 ^ new_n25768;
  assign new_n25809 = new_n25808 ^ new_n25654;
  assign new_n25810 = ~new_n25801 & ~new_n25809;
  assign new_n25811 = new_n25810 ^ new_n25807;
  assign new_n25812 = new_n25799 ^ new_n25684;
  assign new_n25813 = new_n25812 ^ new_n25811;
  assign new_n25814 = new_n25707 ^ new_n25654;
  assign new_n25815 = new_n25814 ^ new_n25812;
  assign new_n25816 = ~new_n25815 & new_n25800;
  assign new_n25817 = new_n25808 ^ new_n25584;
  assign new_n25818 = ~new_n25708 & new_n25817;
  assign new_n25819 = new_n25818 ^ new_n25816;
  assign new_n25820 = new_n25767 ^ new_n25654;
  assign new_n25821 = new_n25820 ^ new_n25819;
  assign new_n25822 = new_n25821 ^ new_n25813;
  assign new_n25823 = new_n25804 ^ new_n25769;
  assign new_n25824 = new_n25779 ^ new_n25769;
  assign new_n25825 = new_n25780 ^ new_n25745;
  assign new_n25826 = new_n25825 ^ new_n25812;
  assign new_n25827 = ~new_n25826 & new_n25824;
  assign new_n25828 = new_n25827 ^ new_n25799;
  assign new_n25829 = new_n25828 ^ new_n25819;
  assign new_n25830 = new_n25829 ^ new_n25823;
  assign new_n25831 = ~new_n25830 & new_n25822;
  assign new_n25832 = new_n25831 ^ new_n25805;
  assign new_n25833 = ~new_n25770 & ~new_n25812;
  assign new_n25834 = new_n25833 ^ new_n25818;
  assign new_n25835 = new_n25834 ^ new_n25809;
  assign new_n25836 = new_n25835 ^ new_n25832;
  assign new_n25837 = new_n25780 ^ new_n25684;
  assign new_n25838 = new_n25817 ^ new_n25779;
  assign new_n25839 = ~new_n25837 & new_n25838;
  assign new_n25840 = new_n25839 ^ new_n25806;
  assign new_n25841 = new_n25833 ^ new_n25816;
  assign new_n25842 = new_n25841 ^ new_n25840;
  assign new_n25843 = ~new_n25842 & new_n25836;
  assign new_n25844 = new_n25843 ^ new_n25684;
  assign new_n25845 = new_n25839 ^ new_n25782;
  assign new_n25846 = new_n25745 ^ new_n25654;
  assign new_n25847 = new_n25827 ^ new_n25807;
  assign new_n25848 = new_n25684 ^ new_n25654;
  assign new_n25849 = new_n25827 ^ new_n25782;
  assign new_n25850 = new_n25849 ^ new_n25841;
  assign new_n25851 = new_n25850 ^ new_n25848;
  assign new_n25852 = new_n25839 ^ new_n25810;
  assign new_n25853 = new_n25852 ^ new_n25684;
  assign new_n25854 = new_n25853 ^ new_n25835;
  assign new_n25855 = new_n25854 ^ new_n25831;
  assign new_n25856 = ~new_n25851 & ~new_n25855;
  assign new_n25857 = new_n25856 ^ new_n25805;
  assign new_n25858 = new_n25857 ^ new_n25835;
  assign new_n25859 = new_n25843 ^ new_n25831;
  assign new_n25860 = ~new_n25854 & ~new_n25859;
  assign new_n25861 = new_n25860 ^ new_n25831;
  assign new_n25862 = new_n25858 & new_n25861;
  assign new_n25863 = new_n25860 ^ new_n25854;
  assign new_n25864 = new_n25863 ^ new_n25862;
  assign new_n25865 = new_n25864 ^ new_n25847;
  assign new_n25866 = new_n25865 ^ new_n25846;
  assign new_n25867 = new_n25866 ^ new_n25845;
  assign new_n25868 = new_n25867 ^ new_n25844;
  assign new_n25869 = ~new_n25770 & ~new_n25868;
  assign new_n25870 = ~new_n25837 & new_n25858;
  assign new_n25871 = new_n25870 ^ new_n25869;
  assign new_n25872 = new_n25862 ^ new_n25856;
  assign new_n25873 = new_n25872 ^ new_n25830;
  assign new_n25874 = ~new_n25801 & ~new_n25873;
  assign new_n25875 = new_n25854 ^ new_n25843;
  assign new_n25876 = ~new_n25875 & new_n25779;
  assign new_n25877 = new_n25863 ^ new_n25822;
  assign new_n25878 = ~new_n25877 & new_n25769;
  assign new_n25879 = new_n25878 ^ new_n25876;
  assign new_n25880 = new_n25879 ^ new_n25874;
  assign new_n25881 = new_n25880 ^ new_n25871;
  assign new_n25882 = ~new_n25875 & new_n25781;
  assign new_n25883 = new_n25866 ^ new_n25707;
  assign new_n25884 = new_n25856 ^ new_n25810;
  assign new_n25885 = new_n25884 ^ new_n25804;
  assign new_n25886 = new_n25885 ^ new_n25883;
  assign new_n25887 = ~new_n25815 & new_n25886;
  assign new_n25888 = new_n25863 ^ new_n25843;
  assign new_n25889 = new_n25888 ^ new_n25842;
  assign new_n25890 = ~new_n25826 & new_n25889;
  assign new_n25891 = new_n25856 ^ new_n25843;
  assign new_n25892 = new_n25853 ^ new_n25805;
  assign new_n25893 = new_n25892 ^ new_n25891;
  assign new_n25894 = ~new_n25708 & ~new_n25893;
  assign new_n25895 = new_n25800 & new_n25886;
  assign new_n25896 = new_n25895 ^ new_n25894;
  assign new_n25897 = new_n25896 ^ new_n25890;
  assign new_n25898 = new_n25862 ^ new_n25851;
  assign new_n25899 = ~new_n25780 & ~new_n25898;
  assign new_n25900 = new_n25899 ^ new_n25897;
  assign new_n25901 = ~new_n25809 & ~new_n25873;
  assign new_n25902 = new_n25901 ^ new_n25900;
  assign new_n25903 = new_n25902 ^ new_n25887;
  assign new_n25904 = new_n25903 ^ new_n25882;
  assign new_n25905 = new_n25904 ^ new_n25881;
  assign new_n25906 = new_n25905 ^ new_n25011;
  assign new_n25907 = new_n25874 ^ new_n25869;
  assign new_n25908 = new_n25899 ^ new_n25887;
  assign new_n25909 = ~new_n25898 & new_n25825;
  assign new_n25910 = new_n25838 & new_n25858;
  assign new_n25911 = new_n25910 ^ new_n25909;
  assign new_n25912 = new_n25911 ^ new_n25896;
  assign new_n25913 = new_n25912 ^ new_n25908;
  assign new_n25914 = new_n25913 ^ new_n25907;
  assign new_n25915 = new_n25914 ^ new_n25906;
  assign new_n25916 = new_n25915 ^ new_n24740;
  assign new_n25917 = new_n22547 ^ new_n22507;
  assign new_n25918 = ~new_n25917 & new_n22435;
  assign new_n25919 = new_n22535 ^ new_n22524;
  assign new_n25920 = new_n22370 & new_n25919;
  assign new_n25921 = new_n25920 ^ new_n25918;
  assign new_n25922 = new_n25921 ^ new_n22542;
  assign new_n25923 = new_n22498 & new_n22541;
  assign new_n25924 = new_n25923 ^ new_n25922;
  assign new_n25925 = new_n25924 ^ new_n22572;
  assign new_n25926 = ~new_n25893 & new_n25817;
  assign new_n25927 = ~new_n25802 & ~new_n25877;
  assign new_n25928 = new_n25927 ^ new_n25926;
  assign new_n25929 = new_n25928 ^ new_n25903;
  assign new_n25930 = new_n22547 ^ new_n22535;
  assign new_n25931 = new_n25930 ^ new_n22534;
  assign new_n25932 = ~new_n25931 & new_n22481;
  assign new_n25933 = new_n25932 ^ new_n22571;
  assign new_n25934 = new_n25933 ^ new_n22561;
  assign new_n25935 = new_n25934 ^ new_n25923;
  assign new_n25936 = new_n25935 ^ new_n22559;
  assign new_n25937 = new_n22502 & new_n22568;
  assign new_n25938 = ~new_n25917 & new_n22508;
  assign new_n25939 = new_n25938 ^ new_n25937;
  assign new_n25940 = new_n25939 ^ new_n25936;
  assign new_n25941 = new_n25940 ^ new_n25929;
  assign new_n25942 = new_n25941 ^ new_n25925;
  assign new_n25943 = new_n24735 ^ new_n24729;
  assign new_n25944 = new_n24719 ^ new_n24704;
  assign new_n25945 = ~new_n24718 & new_n24638;
  assign new_n25946 = ~new_n24671 & ~new_n24694;
  assign new_n25947 = new_n25946 ^ new_n25945;
  assign new_n25948 = new_n25947 ^ new_n24716;
  assign new_n25949 = new_n25948 ^ new_n25944;
  assign new_n25950 = new_n25949 ^ new_n25943;
  assign new_n25951 = new_n23660 ^ new_n23654;
  assign new_n25952 = new_n23644 ^ new_n23629;
  assign new_n25953 = ~new_n23643 & new_n23563;
  assign new_n25954 = ~new_n23596 & ~new_n23619;
  assign new_n25955 = new_n25954 ^ new_n25953;
  assign new_n25956 = new_n25955 ^ new_n23641;
  assign new_n25957 = new_n25956 ^ new_n25952;
  assign new_n25958 = new_n25957 ^ new_n25951;
  assign new_n25959 = new_n25958 ^ new_n25950;
  assign new_n25960 = new_n25959 ^ new_n25942;
  assign new_n25961 = new_n25007 ^ new_n25001;
  assign new_n25962 = ~new_n24929 & new_n24990;
  assign new_n25963 = new_n24944 & new_n24966;
  assign new_n25964 = new_n25963 ^ new_n25962;
  assign new_n25965 = new_n25964 ^ new_n24988;
  assign new_n25966 = new_n24991 ^ new_n24976;
  assign new_n25967 = new_n25966 ^ new_n25965;
  assign new_n25968 = new_n25967 ^ new_n25961;
  assign new_n25969 = new_n25968 ^ new_n23138;
  assign new_n25970 = new_n25969 ^ new_n25914;
  assign new_n25971 = new_n25901 ^ new_n25880;
  assign new_n25972 = new_n25971 ^ new_n25912;
  assign new_n25973 = new_n25972 ^ new_n25970;
  assign new_n25974 = new_n25973 ^ new_n25960;
  assign new_n25975 = new_n22519 & new_n22530;
  assign new_n25976 = new_n25975 ^ new_n22553;
  assign new_n25977 = new_n25976 ^ new_n25922;
  assign new_n25978 = new_n22483 & new_n25919;
  assign new_n25979 = new_n25978 ^ new_n25936;
  assign new_n25980 = new_n25979 ^ new_n25977;
  assign new_n25981 = new_n25927 ^ new_n25910;
  assign new_n25982 = new_n25824 & new_n25889;
  assign new_n25983 = new_n25982 ^ new_n25876;
  assign new_n25984 = new_n25983 ^ new_n25900;
  assign new_n25985 = new_n25984 ^ new_n25981;
  assign new_n25986 = new_n25985 ^ new_n25980;
  assign new_n25987 = new_n25986 ^ new_n25905;
  assign new_n25988 = ~new_n23557 & new_n23657;
  assign new_n25989 = new_n25988 ^ new_n25954;
  assign new_n25990 = new_n23562 & new_n23634;
  assign new_n25991 = new_n25990 ^ new_n23656;
  assign new_n25992 = new_n25991 ^ new_n23645;
  assign new_n25993 = new_n25992 ^ new_n25989;
  assign new_n25994 = ~new_n24632 & new_n24732;
  assign new_n25995 = new_n25994 ^ new_n25946;
  assign new_n25996 = new_n24637 & new_n24709;
  assign new_n25997 = new_n25996 ^ new_n24731;
  assign new_n25998 = new_n25997 ^ new_n24720;
  assign new_n25999 = new_n25998 ^ new_n25995;
  assign new_n26000 = new_n25999 ^ new_n25993;
  assign new_n26001 = ~new_n24905 & new_n25004;
  assign new_n26002 = new_n26001 ^ new_n25963;
  assign new_n26003 = ~new_n24981 & new_n24928;
  assign new_n26004 = new_n26003 ^ new_n25003;
  assign new_n26005 = new_n26004 ^ new_n24992;
  assign new_n26006 = new_n26005 ^ new_n26002;
  assign new_n26007 = new_n26006 ^ new_n23131;
  assign new_n26008 = new_n26007 ^ new_n25941;
  assign new_n26009 = new_n26008 ^ new_n26000;
  assign new_n26010 = new_n26009 ^ new_n25987;
  assign new_n26011 = new_n26010 ^ new_n25974;
  assign new_n26012 = new_n26011 ^ new_n25916;
  assign new_n26013 = new_n25937 ^ new_n22569;
  assign new_n26014 = ~new_n22552 & new_n22480;
  assign new_n26015 = new_n26014 ^ new_n25977;
  assign new_n26016 = new_n26015 ^ new_n26013;
  assign new_n26017 = ~new_n24714 & new_n24642;
  assign new_n26018 = new_n26017 ^ new_n24704;
  assign new_n26019 = new_n25996 ^ new_n24733;
  assign new_n26020 = new_n26019 ^ new_n25994;
  assign new_n26021 = new_n26020 ^ new_n24717;
  assign new_n26022 = new_n26021 ^ new_n26018;
  assign new_n26023 = ~new_n23639 & new_n23567;
  assign new_n26024 = new_n26023 ^ new_n23629;
  assign new_n26025 = new_n25990 ^ new_n23658;
  assign new_n26026 = new_n26025 ^ new_n25988;
  assign new_n26027 = new_n26026 ^ new_n23642;
  assign new_n26028 = new_n26027 ^ new_n26024;
  assign new_n26029 = new_n26028 ^ new_n26022;
  assign new_n26030 = new_n26029 ^ new_n26016;
  assign new_n26031 = ~new_n24985 & new_n24921;
  assign new_n26032 = new_n26031 ^ new_n24976;
  assign new_n26033 = new_n26003 ^ new_n25005;
  assign new_n26034 = new_n26033 ^ new_n26001;
  assign new_n26035 = new_n26034 ^ new_n24989;
  assign new_n26036 = new_n26035 ^ new_n26032;
  assign new_n26037 = new_n26036 ^ new_n23150;
  assign new_n26038 = new_n25926 ^ new_n25887;
  assign new_n26039 = new_n25982 ^ new_n25878;
  assign new_n26040 = new_n26039 ^ new_n25927;
  assign new_n26041 = new_n26040 ^ new_n25897;
  assign new_n26042 = new_n26041 ^ new_n26038;
  assign new_n26043 = new_n26042 ^ new_n26037;
  assign new_n26044 = new_n25926 ^ new_n25894;
  assign new_n26045 = ~new_n25812 & ~new_n25868;
  assign new_n26046 = new_n26045 ^ new_n25881;
  assign new_n26047 = new_n26046 ^ new_n26044;
  assign new_n26048 = new_n26047 ^ new_n26043;
  assign new_n26049 = new_n26048 ^ new_n26030;
  assign new_n26050 = new_n26049 ^ new_n26012;
  assign new_n26051 = new_n26017 ^ new_n24715;
  assign new_n26052 = ~new_n24728 & new_n24631;
  assign new_n26053 = new_n26052 ^ new_n24737;
  assign new_n26054 = new_n26053 ^ new_n26051;
  assign new_n26055 = new_n26023 ^ new_n23640;
  assign new_n26056 = ~new_n23653 & new_n23556;
  assign new_n26057 = new_n26056 ^ new_n23662;
  assign new_n26058 = new_n26057 ^ new_n26055;
  assign new_n26059 = new_n26058 ^ new_n26054;
  assign new_n26060 = new_n26059 ^ new_n26047;
  assign new_n26061 = new_n26031 ^ new_n24986;
  assign new_n26062 = ~new_n24904 & ~new_n25000;
  assign new_n26063 = new_n26062 ^ new_n25009;
  assign new_n26064 = new_n26063 ^ new_n26061;
  assign new_n26065 = new_n26064 ^ new_n23178;
  assign new_n26066 = ~new_n25931 & new_n22436;
  assign new_n26067 = new_n26066 ^ new_n25918;
  assign new_n26068 = new_n26067 ^ new_n25938;
  assign new_n26069 = new_n26068 ^ new_n25935;
  assign new_n26070 = new_n26040 ^ new_n25902;
  assign new_n26071 = new_n26070 ^ new_n26069;
  assign new_n26072 = new_n26071 ^ new_n26065;
  assign new_n26073 = new_n26072 ^ new_n26060;
  assign new_n26074 = new_n26073 ^ new_n26049;
  assign new_n26075 = new_n25008 ^ new_n24979;
  assign new_n26076 = new_n26075 ^ new_n25965;
  assign new_n26077 = new_n26076 ^ new_n23173;
  assign new_n26078 = new_n26077 ^ new_n25972;
  assign new_n26079 = new_n24736 ^ new_n24707;
  assign new_n26080 = new_n26079 ^ new_n25948;
  assign new_n26081 = new_n23661 ^ new_n23632;
  assign new_n26082 = new_n26081 ^ new_n25956;
  assign new_n26083 = new_n26082 ^ new_n26080;
  assign new_n26084 = new_n26083 ^ new_n25941;
  assign new_n26085 = new_n26084 ^ new_n26078;
  assign new_n26086 = new_n26085 ^ new_n26074;
  assign new_n26087 = new_n25974 & new_n26086;
  assign new_n26088 = new_n26087 ^ new_n25974;
  assign new_n26089 = new_n26073 ^ new_n26012;
  assign new_n26090 = new_n25937 ^ new_n22559;
  assign new_n26091 = new_n26068 ^ new_n25933;
  assign new_n26092 = new_n26091 ^ new_n26090;
  assign new_n26093 = new_n26023 ^ new_n25988;
  assign new_n26094 = new_n26093 ^ new_n23647;
  assign new_n26095 = new_n26017 ^ new_n25994;
  assign new_n26096 = new_n26095 ^ new_n24722;
  assign new_n26097 = new_n26096 ^ new_n26094;
  assign new_n26098 = new_n26097 ^ new_n26092;
  assign new_n26099 = new_n26031 ^ new_n26001;
  assign new_n26100 = new_n26099 ^ new_n24994;
  assign new_n26101 = new_n26100 ^ new_n23156;
  assign new_n26102 = new_n26101 ^ new_n25929;
  assign new_n26103 = new_n26102 ^ new_n26042;
  assign new_n26104 = new_n26103 ^ new_n26098;
  assign new_n26105 = new_n26104 ^ new_n25974;
  assign new_n26106 = ~new_n26105 & new_n26089;
  assign new_n26107 = new_n26106 ^ new_n26088;
  assign new_n26108 = new_n26104 ^ new_n25916;
  assign new_n26109 = new_n26108 ^ new_n26107;
  assign new_n26110 = new_n26034 ^ new_n24993;
  assign new_n26111 = new_n26110 ^ new_n23160;
  assign new_n26112 = new_n26026 ^ new_n23646;
  assign new_n26113 = new_n26020 ^ new_n24721;
  assign new_n26114 = new_n26113 ^ new_n26112;
  assign new_n26115 = new_n26114 ^ new_n26111;
  assign new_n26116 = new_n26115 ^ new_n25941;
  assign new_n26117 = new_n25938 ^ new_n22564;
  assign new_n26118 = new_n26066 ^ new_n25920;
  assign new_n26119 = new_n26118 ^ new_n25934;
  assign new_n26120 = new_n26119 ^ new_n26117;
  assign new_n26121 = new_n26120 ^ new_n26070;
  assign new_n26122 = new_n26121 ^ new_n25985;
  assign new_n26123 = new_n26122 ^ new_n26116;
  assign new_n26124 = new_n26123 ^ new_n25916;
  assign new_n26125 = new_n26123 ^ new_n26073;
  assign new_n26126 = new_n26125 ^ new_n26108;
  assign new_n26127 = ~new_n26126 & new_n26124;
  assign new_n26128 = new_n26123 ^ new_n26104;
  assign new_n26129 = new_n26050 & new_n26128;
  assign new_n26130 = new_n26129 ^ new_n26127;
  assign new_n26131 = new_n26073 ^ new_n26010;
  assign new_n26132 = new_n26131 ^ new_n26130;
  assign new_n26133 = new_n26132 ^ new_n26109;
  assign new_n26134 = new_n26128 ^ new_n26011;
  assign new_n26135 = new_n26124 ^ new_n26105;
  assign new_n26136 = ~new_n26134 & ~new_n26135;
  assign new_n26137 = new_n26136 ^ new_n26049;
  assign new_n26138 = new_n26137 ^ new_n26134;
  assign new_n26139 = new_n26134 ^ new_n26085;
  assign new_n26140 = new_n26086 ^ new_n25974;
  assign new_n26141 = new_n26140 ^ new_n26108;
  assign new_n26142 = new_n26139 & new_n26141;
  assign new_n26143 = new_n26142 ^ new_n26130;
  assign new_n26144 = new_n26143 ^ new_n25916;
  assign new_n26145 = new_n26144 ^ new_n26138;
  assign new_n26146 = ~new_n26133 & new_n26145;
  assign new_n26147 = new_n26134 ^ new_n26074;
  assign new_n26148 = ~new_n26147 & new_n26108;
  assign new_n26149 = new_n26148 ^ new_n26129;
  assign new_n26150 = new_n26149 ^ new_n26089;
  assign new_n26151 = new_n26104 ^ new_n26086;
  assign new_n26152 = new_n26085 ^ new_n26050;
  assign new_n26153 = ~new_n26151 & ~new_n26152;
  assign new_n26154 = new_n26153 ^ new_n26106;
  assign new_n26155 = new_n26154 ^ new_n26104;
  assign new_n26156 = new_n26155 ^ new_n26150;
  assign new_n26157 = new_n26156 ^ new_n26146;
  assign new_n26158 = new_n26104 ^ new_n26073;
  assign new_n26159 = new_n26123 ^ new_n26086;
  assign new_n26160 = ~new_n26085 & ~new_n26159;
  assign new_n26161 = new_n26160 ^ new_n26142;
  assign new_n26162 = new_n26148 ^ new_n26127;
  assign new_n26163 = new_n26162 ^ new_n26161;
  assign new_n26164 = new_n26163 ^ new_n26158;
  assign new_n26165 = ~new_n26164 & new_n26157;
  assign new_n26166 = new_n26160 ^ new_n26123;
  assign new_n26167 = new_n26166 ^ new_n26137;
  assign new_n26168 = new_n26167 ^ new_n26146;
  assign new_n26169 = new_n26168 ^ new_n26150;
  assign new_n26170 = new_n26153 ^ new_n26087;
  assign new_n26171 = new_n26170 ^ new_n26162;
  assign new_n26172 = ~new_n26169 & ~new_n26171;
  assign new_n26173 = new_n26172 ^ new_n26165;
  assign new_n26174 = new_n26167 ^ new_n26155;
  assign new_n26175 = new_n26174 ^ new_n26173;
  assign new_n26176 = ~new_n26175 & new_n26050;
  assign new_n26177 = ~new_n26175 & new_n26128;
  assign new_n26178 = new_n26177 ^ new_n26176;
  assign new_n26179 = new_n26172 ^ new_n26104;
  assign new_n26180 = new_n26160 ^ new_n26153;
  assign new_n26181 = new_n26073 ^ new_n25974;
  assign new_n26182 = new_n26142 ^ new_n26088;
  assign new_n26183 = new_n26167 ^ new_n26165;
  assign new_n26184 = new_n26183 ^ new_n26150;
  assign new_n26185 = new_n26172 ^ new_n26146;
  assign new_n26186 = ~new_n26185 & new_n26156;
  assign new_n26187 = new_n26186 ^ new_n26146;
  assign new_n26188 = ~new_n26184 & new_n26187;
  assign new_n26189 = new_n26186 ^ new_n26156;
  assign new_n26190 = new_n26189 ^ new_n26188;
  assign new_n26191 = new_n26190 ^ new_n26182;
  assign new_n26192 = new_n26191 ^ new_n26181;
  assign new_n26193 = new_n26192 ^ new_n26180;
  assign new_n26194 = new_n26193 ^ new_n26179;
  assign new_n26195 = new_n26108 & new_n26194;
  assign new_n26196 = ~new_n26151 & ~new_n26184;
  assign new_n26197 = ~new_n26147 & new_n26194;
  assign new_n26198 = new_n26197 ^ new_n26196;
  assign new_n26199 = new_n26188 ^ new_n26165;
  assign new_n26200 = new_n26199 ^ new_n26145;
  assign new_n26201 = ~new_n26105 & new_n26200;
  assign new_n26202 = new_n26172 ^ new_n26156;
  assign new_n26203 = ~new_n26085 & new_n26202;
  assign new_n26204 = new_n26189 ^ new_n26133;
  assign new_n26205 = ~new_n26134 & ~new_n26204;
  assign new_n26206 = new_n26205 ^ new_n26203;
  assign new_n26207 = new_n26206 ^ new_n26201;
  assign new_n26208 = new_n26207 ^ new_n26198;
  assign new_n26209 = new_n26208 ^ new_n26195;
  assign new_n26210 = new_n26209 ^ new_n26178;
  assign new_n26211 = new_n23987 ^ new_n23537;
  assign new_n26212 = new_n26211 ^ new_n22462;
  assign new_n26213 = new_n26212 ^ new_n19989;
  assign new_n26214 = new_n22409 ^ new_n22244;
  assign new_n26215 = new_n26214 ^ new_n26213;
  assign new_n26216 = new_n22477 ^ new_n22302;
  assign new_n26217 = new_n23994 ^ new_n23522;
  assign new_n26218 = new_n26217 ^ new_n22244;
  assign new_n26219 = new_n26218 ^ new_n22368;
  assign new_n26220 = new_n26219 ^ new_n26216;
  assign new_n26221 = new_n22462 ^ new_n22375;
  assign new_n26222 = new_n26221 ^ new_n22466;
  assign new_n26223 = new_n24001 ^ new_n23478;
  assign new_n26224 = new_n26223 ^ new_n22302;
  assign new_n26225 = new_n26224 ^ new_n22423;
  assign new_n26226 = new_n26225 ^ new_n26222;
  assign new_n26227 = new_n26226 ^ new_n26220;
  assign new_n26228 = new_n26227 ^ new_n26215;
  assign new_n26229 = new_n22355 ^ new_n22274;
  assign new_n26230 = new_n24008 ^ new_n23311;
  assign new_n26231 = new_n26230 ^ new_n22342;
  assign new_n26232 = new_n26231 ^ new_n22454;
  assign new_n26233 = new_n26232 ^ new_n26229;
  assign new_n26234 = new_n26233 ^ new_n26228;
  assign new_n26235 = new_n22454 ^ new_n21072;
  assign new_n26236 = new_n24014 ^ new_n23457;
  assign new_n26237 = new_n26236 ^ new_n22301;
  assign new_n26238 = new_n26237 ^ new_n22450;
  assign new_n26239 = new_n26238 ^ new_n26235;
  assign new_n26240 = new_n26239 ^ new_n26215;
  assign new_n26241 = new_n22441 ^ new_n22355;
  assign new_n26242 = new_n24036 ^ new_n22682;
  assign new_n26243 = new_n22431 ^ new_n22427;
  assign new_n26244 = new_n26243 ^ new_n26242;
  assign new_n26245 = new_n26244 ^ new_n26241;
  assign new_n26246 = new_n26245 ^ new_n26233;
  assign new_n26247 = new_n24018 ^ new_n23442;
  assign new_n26248 = new_n26247 ^ new_n22302;
  assign new_n26249 = new_n26248 ^ new_n22308;
  assign new_n26250 = new_n22431 ^ new_n22375;
  assign new_n26251 = new_n26250 ^ new_n22385;
  assign new_n26252 = new_n26251 ^ new_n26249;
  assign new_n26253 = new_n26252 ^ new_n26239;
  assign new_n26254 = new_n26253 ^ new_n26227;
  assign new_n26255 = new_n26254 ^ new_n26246;
  assign new_n26256 = new_n26240 & new_n26255;
  assign new_n26257 = new_n26234 & new_n26253;
  assign new_n26258 = new_n26257 ^ new_n26256;
  assign new_n26259 = new_n26245 ^ new_n26228;
  assign new_n26260 = new_n26259 ^ new_n26258;
  assign new_n26261 = new_n24031 ^ new_n23385;
  assign new_n26262 = new_n26261 ^ new_n19999;
  assign new_n26263 = new_n22365 ^ new_n21199;
  assign new_n26264 = new_n26263 ^ new_n22302;
  assign new_n26265 = new_n26264 ^ new_n26262;
  assign new_n26266 = new_n26265 ^ new_n26246;
  assign new_n26267 = new_n26266 ^ new_n26239;
  assign new_n26268 = new_n26265 ^ new_n26234;
  assign new_n26269 = new_n26267 & new_n26268;
  assign new_n26270 = new_n26239 ^ new_n26220;
  assign new_n26271 = new_n26259 & new_n26270;
  assign new_n26272 = new_n26271 ^ new_n26269;
  assign new_n26273 = new_n26272 ^ new_n26239;
  assign new_n26274 = new_n26273 ^ new_n26260;
  assign new_n26275 = ~new_n26220 & ~new_n26266;
  assign new_n26276 = new_n26275 ^ new_n26220;
  assign new_n26277 = new_n26276 ^ new_n26271;
  assign new_n26278 = new_n26277 ^ new_n26240;
  assign new_n26279 = new_n26252 ^ new_n26215;
  assign new_n26280 = new_n26252 ^ new_n26245;
  assign new_n26281 = new_n26280 ^ new_n26240;
  assign new_n26282 = new_n26279 & new_n26281;
  assign new_n26283 = new_n26282 ^ new_n26257;
  assign new_n26284 = new_n26245 ^ new_n26226;
  assign new_n26285 = new_n26284 ^ new_n26283;
  assign new_n26286 = new_n26285 ^ new_n26278;
  assign new_n26287 = new_n26252 ^ new_n26220;
  assign new_n26288 = new_n26287 ^ new_n26240;
  assign new_n26289 = new_n26254 & new_n26288;
  assign new_n26290 = new_n26289 ^ new_n26233;
  assign new_n26291 = new_n26290 ^ new_n26254;
  assign new_n26292 = new_n26265 ^ new_n26254;
  assign new_n26293 = new_n26266 ^ new_n26220;
  assign new_n26294 = new_n26293 ^ new_n26240;
  assign new_n26295 = new_n26292 & new_n26294;
  assign new_n26296 = new_n26295 ^ new_n26283;
  assign new_n26297 = new_n26296 ^ new_n26215;
  assign new_n26298 = new_n26297 ^ new_n26291;
  assign new_n26299 = ~new_n26286 & new_n26298;
  assign new_n26300 = new_n26299 ^ new_n26274;
  assign new_n26301 = new_n26245 ^ new_n26239;
  assign new_n26302 = new_n26266 ^ new_n26252;
  assign new_n26303 = new_n26265 & new_n26302;
  assign new_n26304 = new_n26303 ^ new_n26295;
  assign new_n26305 = new_n26282 ^ new_n26256;
  assign new_n26306 = new_n26305 ^ new_n26304;
  assign new_n26307 = new_n26306 ^ new_n26301;
  assign new_n26308 = new_n26300 & new_n26307;
  assign new_n26309 = new_n26303 ^ new_n26252;
  assign new_n26310 = new_n26309 ^ new_n26290;
  assign new_n26311 = new_n26310 ^ new_n26299;
  assign new_n26312 = new_n26311 ^ new_n26260;
  assign new_n26313 = new_n26275 ^ new_n26269;
  assign new_n26314 = new_n26313 ^ new_n26305;
  assign new_n26315 = ~new_n26314 & new_n26312;
  assign new_n26316 = new_n26315 ^ new_n26308;
  assign new_n26317 = new_n26310 ^ new_n26273;
  assign new_n26318 = new_n26317 ^ new_n26316;
  assign new_n26319 = new_n26234 & new_n26318;
  assign new_n26320 = new_n26315 ^ new_n26299;
  assign new_n26321 = ~new_n26274 & ~new_n26320;
  assign new_n26322 = new_n26321 ^ new_n26315;
  assign new_n26323 = new_n26322 ^ new_n26300;
  assign new_n26324 = new_n26323 ^ new_n26286;
  assign new_n26325 = new_n26288 & new_n26324;
  assign new_n26326 = new_n26325 ^ new_n26319;
  assign new_n26327 = new_n26310 ^ new_n26308;
  assign new_n26328 = new_n26327 ^ new_n26260;
  assign new_n26329 = ~new_n26322 & new_n26328;
  assign new_n26330 = new_n26329 ^ new_n26308;
  assign new_n26331 = new_n26330 ^ new_n26298;
  assign new_n26332 = new_n26259 & new_n26331;
  assign new_n26333 = new_n26329 ^ new_n26307;
  assign new_n26334 = new_n26266 & new_n26333;
  assign new_n26335 = new_n26253 & new_n26318;
  assign new_n26336 = new_n26245 ^ new_n26220;
  assign new_n26337 = new_n26295 ^ new_n26276;
  assign new_n26338 = new_n26329 ^ new_n26323;
  assign new_n26339 = new_n26338 ^ new_n26337;
  assign new_n26340 = new_n26339 ^ new_n26336;
  assign new_n26341 = new_n26340 ^ new_n26252;
  assign new_n26342 = new_n26308 ^ new_n26271;
  assign new_n26343 = new_n26342 ^ new_n26290;
  assign new_n26344 = new_n26343 ^ new_n26341;
  assign new_n26345 = new_n26279 & new_n26344;
  assign new_n26346 = new_n26345 ^ new_n26335;
  assign new_n26347 = new_n26323 ^ new_n26315;
  assign new_n26348 = new_n26347 ^ new_n26314;
  assign new_n26349 = new_n26294 & new_n26348;
  assign new_n26350 = new_n26349 ^ new_n26346;
  assign new_n26351 = new_n26350 ^ new_n26334;
  assign new_n26352 = new_n26351 ^ new_n26332;
  assign new_n26353 = new_n26281 & new_n26344;
  assign new_n26354 = new_n26353 ^ new_n26352;
  assign new_n26355 = new_n26354 ^ new_n26326;
  assign new_n26356 = new_n25688 ^ new_n25622;
  assign new_n26357 = new_n24230 ^ new_n20434;
  assign new_n26358 = new_n26357 ^ new_n25175;
  assign new_n26359 = new_n26358 ^ new_n25582;
  assign new_n26360 = new_n26359 ^ new_n26356;
  assign new_n26361 = new_n25716 ^ new_n25672;
  assign new_n26362 = new_n26361 ^ new_n25777;
  assign new_n26363 = new_n24596 ^ new_n20461;
  assign new_n26364 = new_n26363 ^ new_n25739;
  assign new_n26365 = new_n26364 ^ new_n25794;
  assign new_n26366 = new_n26365 ^ new_n26362;
  assign new_n26367 = new_n25763 ^ new_n25699;
  assign new_n26368 = new_n26367 ^ new_n25705;
  assign new_n26369 = new_n24561 ^ new_n20467;
  assign new_n26370 = new_n26369 ^ new_n25672;
  assign new_n26371 = new_n26370 ^ new_n25790;
  assign new_n26372 = new_n26371 ^ new_n26368;
  assign new_n26373 = new_n26372 ^ new_n26366;
  assign new_n26374 = new_n25789 ^ new_n25748;
  assign new_n26375 = new_n26374 ^ new_n25753;
  assign new_n26376 = new_n24616 ^ new_n20481;
  assign new_n26377 = new_n26376 ^ new_n25725;
  assign new_n26378 = new_n26377 ^ new_n26375;
  assign new_n26379 = new_n26378 ^ new_n26373;
  assign new_n26380 = new_n26379 ^ new_n26360;
  assign new_n26381 = new_n24541 ^ new_n20472;
  assign new_n26382 = new_n26381 ^ new_n25437;
  assign new_n26383 = new_n25692 ^ new_n25671;
  assign new_n26384 = new_n26383 ^ new_n25681;
  assign new_n26385 = new_n26384 ^ new_n26382;
  assign new_n26386 = new_n26385 ^ new_n26360;
  assign new_n26387 = new_n26385 ^ new_n26378;
  assign new_n26388 = new_n24517 ^ new_n20450;
  assign new_n26389 = new_n26388 ^ new_n25672;
  assign new_n26390 = new_n26389 ^ new_n25764;
  assign new_n26391 = new_n25687 ^ new_n25645;
  assign new_n26392 = new_n26391 ^ new_n25651;
  assign new_n26393 = new_n26392 ^ new_n26390;
  assign new_n26394 = new_n26393 ^ new_n26385;
  assign new_n26395 = new_n26394 ^ new_n26373;
  assign new_n26396 = new_n25623 ^ new_n25307;
  assign new_n26397 = new_n24436 ^ new_n20439;
  assign new_n26398 = new_n26397 ^ new_n25155;
  assign new_n26399 = new_n26398 ^ new_n25676;
  assign new_n26400 = new_n26399 ^ new_n26396;
  assign new_n26401 = new_n26400 ^ new_n26360;
  assign new_n26402 = new_n26401 ^ new_n26395;
  assign new_n26403 = ~new_n26402 & new_n26387;
  assign new_n26404 = new_n26393 ^ new_n26378;
  assign new_n26405 = new_n26393 ^ new_n26360;
  assign new_n26406 = new_n26405 ^ new_n26387;
  assign new_n26407 = ~new_n26406 & new_n26404;
  assign new_n26408 = new_n26407 ^ new_n26403;
  assign new_n26409 = new_n25774 ^ new_n25672;
  assign new_n26410 = new_n24475 ^ new_n20445;
  assign new_n26411 = new_n26410 ^ new_n25743;
  assign new_n26412 = new_n26411 ^ new_n25730;
  assign new_n26413 = new_n26412 ^ new_n26409;
  assign new_n26414 = new_n26413 ^ new_n26401;
  assign new_n26415 = new_n26414 ^ new_n26366;
  assign new_n26416 = new_n26415 ^ new_n26387;
  assign new_n26417 = new_n26413 ^ new_n26395;
  assign new_n26418 = new_n26416 & new_n26417;
  assign new_n26419 = new_n26414 ^ new_n26393;
  assign new_n26420 = ~new_n26413 & ~new_n26419;
  assign new_n26421 = new_n26420 ^ new_n26418;
  assign new_n26422 = new_n26421 ^ new_n26408;
  assign new_n26423 = new_n26422 ^ new_n26386;
  assign new_n26424 = new_n26400 ^ new_n26379;
  assign new_n26425 = new_n26394 & new_n26424;
  assign new_n26426 = new_n26425 ^ new_n26403;
  assign new_n26427 = new_n26426 ^ new_n26380;
  assign new_n26428 = new_n26385 ^ new_n26366;
  assign new_n26429 = ~new_n26428 & new_n26380;
  assign new_n26430 = new_n26414 ^ new_n26385;
  assign new_n26431 = new_n26424 ^ new_n26413;
  assign new_n26432 = ~new_n26430 & ~new_n26431;
  assign new_n26433 = new_n26432 ^ new_n26429;
  assign new_n26434 = new_n26433 ^ new_n26385;
  assign new_n26435 = new_n26434 ^ new_n26427;
  assign new_n26436 = new_n26366 & new_n26414;
  assign new_n26437 = new_n26436 ^ new_n26366;
  assign new_n26438 = new_n26437 ^ new_n26429;
  assign new_n26439 = new_n26438 ^ new_n26387;
  assign new_n26440 = new_n26425 ^ new_n26407;
  assign new_n26441 = new_n26372 ^ new_n26360;
  assign new_n26442 = new_n26441 ^ new_n26440;
  assign new_n26443 = new_n26442 ^ new_n26439;
  assign new_n26444 = new_n26428 ^ new_n26404;
  assign new_n26445 = ~new_n26395 & ~new_n26444;
  assign new_n26446 = new_n26445 ^ new_n26400;
  assign new_n26447 = new_n26446 ^ new_n26395;
  assign new_n26448 = new_n26440 ^ new_n26418;
  assign new_n26449 = new_n26448 ^ new_n26378;
  assign new_n26450 = new_n26449 ^ new_n26447;
  assign new_n26451 = ~new_n26443 & new_n26450;
  assign new_n26452 = new_n26451 ^ new_n26435;
  assign new_n26453 = ~new_n26423 & new_n26452;
  assign new_n26454 = new_n26420 ^ new_n26393;
  assign new_n26455 = new_n26454 ^ new_n26446;
  assign new_n26456 = new_n26455 ^ new_n26453;
  assign new_n26457 = new_n26456 ^ new_n26427;
  assign new_n26458 = new_n26455 ^ new_n26451;
  assign new_n26459 = new_n26458 ^ new_n26427;
  assign new_n26460 = new_n26436 ^ new_n26432;
  assign new_n26461 = new_n26460 ^ new_n26408;
  assign new_n26462 = ~new_n26459 & ~new_n26461;
  assign new_n26463 = new_n26462 ^ new_n26451;
  assign new_n26464 = ~new_n26463 & new_n26435;
  assign new_n26465 = new_n26464 ^ new_n26451;
  assign new_n26466 = ~new_n26457 & new_n26465;
  assign new_n26467 = new_n26466 ^ new_n26453;
  assign new_n26468 = new_n26467 ^ new_n26450;
  assign new_n26469 = new_n26380 & new_n26468;
  assign new_n26470 = new_n26466 ^ new_n26423;
  assign new_n26471 = ~new_n26414 & ~new_n26470;
  assign new_n26472 = new_n26464 ^ new_n26435;
  assign new_n26473 = new_n26472 ^ new_n26462;
  assign new_n26474 = new_n26473 ^ new_n26461;
  assign new_n26475 = ~new_n26474 & new_n26416;
  assign new_n26476 = new_n26366 ^ new_n26360;
  assign new_n26477 = new_n26437 ^ new_n26418;
  assign new_n26478 = new_n26472 ^ new_n26466;
  assign new_n26479 = new_n26478 ^ new_n26477;
  assign new_n26480 = new_n26479 ^ new_n26476;
  assign new_n26481 = new_n26480 ^ new_n26393;
  assign new_n26482 = new_n26453 ^ new_n26429;
  assign new_n26483 = new_n26482 ^ new_n26446;
  assign new_n26484 = new_n26483 ^ new_n26481;
  assign new_n26485 = ~new_n26484 & new_n26404;
  assign new_n26486 = new_n26462 ^ new_n26453;
  assign new_n26487 = new_n26455 ^ new_n26434;
  assign new_n26488 = new_n26487 ^ new_n26486;
  assign new_n26489 = ~new_n26488 & new_n26394;
  assign new_n26490 = new_n26489 ^ new_n26485;
  assign new_n26491 = new_n26490 ^ new_n26475;
  assign new_n26492 = new_n26491 ^ new_n26471;
  assign new_n26493 = new_n26492 ^ new_n26469;
  assign new_n26494 = ~new_n26406 & ~new_n26484;
  assign new_n26495 = new_n26494 ^ new_n26493;
  assign new_n26496 = new_n26472 ^ new_n26443;
  assign new_n26497 = ~new_n26444 & ~new_n26496;
  assign new_n26498 = ~new_n26488 & new_n26424;
  assign new_n26499 = new_n26498 ^ new_n26497;
  assign new_n26500 = new_n26499 ^ new_n26495;
  assign new_n26501 = new_n26500 ^ new_n26355;
  assign new_n26502 = new_n24542 ^ new_n24518;
  assign new_n26503 = new_n24597 ^ new_n24562;
  assign new_n26504 = new_n26503 ^ new_n26502;
  assign new_n26505 = new_n26504 ^ new_n24476;
  assign new_n26506 = new_n26503 ^ new_n24617;
  assign new_n26507 = new_n26506 ^ new_n24437;
  assign new_n26508 = new_n26502 & new_n26507;
  assign new_n26509 = new_n24617 ^ new_n24542;
  assign new_n26510 = new_n24437 ^ new_n24231;
  assign new_n26511 = new_n26510 ^ new_n26504;
  assign new_n26512 = new_n26509 & new_n26511;
  assign new_n26513 = new_n26512 ^ new_n26508;
  assign new_n26514 = new_n26506 ^ new_n24231;
  assign new_n26515 = new_n26514 ^ new_n26513;
  assign new_n26516 = new_n24597 ^ new_n24542;
  assign new_n26517 = new_n26514 & new_n26516;
  assign new_n26518 = new_n26510 ^ new_n24476;
  assign new_n26519 = new_n26518 ^ new_n24542;
  assign new_n26520 = new_n26507 ^ new_n24476;
  assign new_n26521 = new_n26519 & new_n26520;
  assign new_n26522 = new_n26521 ^ new_n26517;
  assign new_n26523 = new_n26522 ^ new_n24542;
  assign new_n26524 = new_n26523 ^ new_n26515;
  assign new_n26525 = ~new_n24597 & ~new_n26518;
  assign new_n26526 = new_n26525 ^ new_n24597;
  assign new_n26527 = new_n26526 ^ new_n26517;
  assign new_n26528 = new_n26527 ^ new_n26509;
  assign new_n26529 = new_n24518 ^ new_n24231;
  assign new_n26530 = new_n26529 ^ new_n26509;
  assign new_n26531 = new_n24617 ^ new_n24518;
  assign new_n26532 = new_n26530 & new_n26531;
  assign new_n26533 = new_n26532 ^ new_n26508;
  assign new_n26534 = new_n24562 ^ new_n24231;
  assign new_n26535 = new_n26534 ^ new_n26533;
  assign new_n26536 = new_n26535 ^ new_n26528;
  assign new_n26537 = new_n24597 ^ new_n24518;
  assign new_n26538 = new_n26537 ^ new_n26509;
  assign new_n26539 = new_n26504 & new_n26538;
  assign new_n26540 = new_n26539 ^ new_n24437;
  assign new_n26541 = new_n26540 ^ new_n26504;
  assign new_n26542 = new_n26518 ^ new_n24597;
  assign new_n26543 = new_n26542 ^ new_n26509;
  assign new_n26544 = new_n26505 & new_n26543;
  assign new_n26545 = new_n26544 ^ new_n24617;
  assign new_n26546 = new_n26545 ^ new_n26533;
  assign new_n26547 = new_n26546 ^ new_n26541;
  assign new_n26548 = ~new_n26536 & new_n26547;
  assign new_n26549 = new_n26518 ^ new_n24518;
  assign new_n26550 = new_n24476 & new_n26549;
  assign new_n26551 = new_n26550 ^ new_n24518;
  assign new_n26552 = new_n26551 ^ new_n26540;
  assign new_n26553 = new_n26552 ^ new_n26548;
  assign new_n26554 = new_n26553 ^ new_n26515;
  assign new_n26555 = new_n26525 ^ new_n26521;
  assign new_n26556 = new_n26532 ^ new_n26512;
  assign new_n26557 = new_n26556 ^ new_n26555;
  assign new_n26558 = ~new_n26557 & new_n26554;
  assign new_n26559 = new_n26558 ^ new_n26548;
  assign new_n26560 = ~new_n26559 & new_n26524;
  assign new_n26561 = new_n26560 ^ new_n26524;
  assign new_n26562 = new_n26561 ^ new_n26558;
  assign new_n26563 = new_n26562 ^ new_n26557;
  assign new_n26564 = ~new_n26563 & new_n26505;
  assign new_n26565 = new_n26561 ^ new_n26536;
  assign new_n26566 = ~new_n26565 & new_n26504;
  assign new_n26567 = new_n26566 ^ new_n26564;
  assign new_n26568 = ~new_n26565 & new_n26538;
  assign new_n26569 = new_n26568 ^ new_n26567;
  assign new_n26570 = new_n24542 ^ new_n24231;
  assign new_n26571 = new_n26550 ^ new_n26544;
  assign new_n26572 = new_n26571 ^ new_n26556;
  assign new_n26573 = new_n26572 ^ new_n26570;
  assign new_n26574 = new_n26548 ^ new_n26524;
  assign new_n26575 = new_n26573 & new_n26574;
  assign new_n26576 = new_n26575 ^ new_n26552;
  assign new_n26577 = new_n26576 ^ new_n26515;
  assign new_n26578 = new_n26560 ^ new_n26548;
  assign new_n26579 = new_n26577 & new_n26578;
  assign new_n26580 = new_n26579 ^ new_n26573;
  assign new_n26581 = new_n26518 & new_n26580;
  assign new_n26582 = new_n26575 ^ new_n26558;
  assign new_n26583 = new_n26552 ^ new_n26523;
  assign new_n26584 = new_n26583 ^ new_n26582;
  assign new_n26585 = new_n26502 & new_n26584;
  assign new_n26586 = new_n24597 ^ new_n24231;
  assign new_n26587 = new_n26544 ^ new_n26526;
  assign new_n26588 = new_n26579 ^ new_n26561;
  assign new_n26589 = new_n26588 ^ new_n26587;
  assign new_n26590 = new_n26589 ^ new_n26586;
  assign new_n26591 = new_n26590 ^ new_n24518;
  assign new_n26592 = new_n26575 ^ new_n26517;
  assign new_n26593 = new_n26592 ^ new_n26540;
  assign new_n26594 = new_n26593 ^ new_n26591;
  assign new_n26595 = ~new_n26594 & new_n26531;
  assign new_n26596 = new_n26595 ^ new_n26585;
  assign new_n26597 = ~new_n26563 & new_n26543;
  assign new_n26598 = new_n26597 ^ new_n26596;
  assign new_n26599 = new_n26598 ^ new_n26581;
  assign new_n26600 = new_n26579 ^ new_n26575;
  assign new_n26601 = new_n26600 ^ new_n26547;
  assign new_n26602 = new_n26514 & new_n26601;
  assign new_n26603 = new_n26602 ^ new_n26599;
  assign new_n26604 = new_n26603 ^ new_n26569;
  assign new_n26605 = new_n26604 ^ new_n12249;
  assign new_n26606 = new_n26605 ^ new_n26501;
  assign new_n26607 = new_n23419 ^ new_n23369;
  assign new_n26608 = new_n22259 ^ new_n20957;
  assign new_n26609 = new_n26608 ^ new_n11703;
  assign new_n26610 = new_n26609 ^ new_n23462;
  assign new_n26611 = new_n26610 ^ new_n23331;
  assign new_n26612 = new_n26611 ^ new_n26607;
  assign new_n26613 = new_n22415 ^ new_n20971;
  assign new_n26614 = new_n26613 ^ new_n11694;
  assign new_n26615 = new_n26614 ^ new_n23128;
  assign new_n26616 = new_n23470 ^ new_n23462;
  assign new_n26617 = new_n26616 ^ new_n26615;
  assign new_n26618 = new_n23499 ^ new_n23448;
  assign new_n26619 = new_n26618 ^ new_n23484;
  assign new_n26620 = new_n26619 ^ new_n26617;
  assign new_n26621 = new_n26620 ^ new_n26612;
  assign new_n26622 = new_n23552 ^ new_n23484;
  assign new_n26623 = new_n26622 ^ new_n23542;
  assign new_n26624 = new_n22391 ^ new_n20798;
  assign new_n26625 = new_n26624 ^ new_n11718;
  assign new_n26626 = new_n26625 ^ new_n26616;
  assign new_n26627 = new_n26626 ^ new_n23432;
  assign new_n26628 = new_n26627 ^ new_n26623;
  assign new_n26629 = new_n26616 ^ new_n23404;
  assign new_n26630 = new_n26629 ^ new_n23548;
  assign new_n26631 = new_n21185 ^ new_n20856;
  assign new_n26632 = new_n26631 ^ new_n11711;
  assign new_n26633 = new_n26632 ^ new_n23528;
  assign new_n26634 = new_n26633 ^ new_n23395;
  assign new_n26635 = new_n26634 ^ new_n26630;
  assign new_n26636 = new_n26635 ^ new_n26628;
  assign new_n26637 = new_n26636 ^ new_n26621;
  assign new_n26638 = new_n22360 ^ new_n20936;
  assign new_n26639 = new_n26638 ^ new_n11755;
  assign new_n26640 = new_n26639 ^ new_n23395;
  assign new_n26641 = new_n26616 ^ new_n23508;
  assign new_n26642 = new_n26641 ^ new_n26640;
  assign new_n26643 = new_n26642 ^ new_n26637;
  assign new_n26644 = new_n23516 ^ new_n23495;
  assign new_n26645 = new_n22470 ^ new_n20430;
  assign new_n26646 = new_n26645 ^ new_n11726;
  assign new_n26647 = new_n26646 ^ new_n23542;
  assign new_n26648 = new_n26647 ^ new_n23528;
  assign new_n26649 = new_n26648 ^ new_n26644;
  assign new_n26650 = new_n26649 ^ new_n26636;
  assign new_n26651 = new_n23467 ^ new_n23272;
  assign new_n26652 = new_n22445 ^ new_n20898;
  assign new_n26653 = new_n26652 ^ new_n11739;
  assign new_n26654 = new_n26653 ^ new_n23331;
  assign new_n26655 = new_n26654 ^ new_n22835;
  assign new_n26656 = new_n26655 ^ new_n26651;
  assign new_n26657 = new_n26656 ^ new_n26650;
  assign new_n26658 = new_n26621 & new_n26657;
  assign new_n26659 = new_n26649 ^ new_n26612;
  assign new_n26660 = new_n23351 ^ new_n22835;
  assign new_n26661 = new_n22328 ^ new_n20927;
  assign new_n26662 = new_n26661 ^ new_n11733;
  assign new_n26663 = new_n23448 ^ new_n23436;
  assign new_n26664 = new_n26663 ^ new_n26662;
  assign new_n26665 = new_n26664 ^ new_n26660;
  assign new_n26666 = new_n26665 ^ new_n26656;
  assign new_n26667 = new_n26666 ^ new_n26637;
  assign new_n26668 = ~new_n26667 & new_n26659;
  assign new_n26669 = new_n26668 ^ new_n26658;
  assign new_n26670 = new_n26665 ^ new_n26650;
  assign new_n26671 = new_n26670 ^ new_n26669;
  assign new_n26672 = new_n26635 ^ new_n26612;
  assign new_n26673 = ~new_n26672 & new_n26670;
  assign new_n26674 = new_n26666 ^ new_n26642;
  assign new_n26675 = new_n26674 ^ new_n26612;
  assign new_n26676 = new_n26657 ^ new_n26642;
  assign new_n26677 = ~new_n26675 & ~new_n26676;
  assign new_n26678 = new_n26677 ^ new_n26673;
  assign new_n26679 = new_n26678 ^ new_n26612;
  assign new_n26680 = new_n26679 ^ new_n26671;
  assign new_n26681 = new_n26635 & new_n26674;
  assign new_n26682 = new_n26681 ^ new_n26635;
  assign new_n26683 = new_n26682 ^ new_n26673;
  assign new_n26684 = new_n26683 ^ new_n26659;
  assign new_n26685 = new_n26649 ^ new_n26620;
  assign new_n26686 = new_n26665 ^ new_n26620;
  assign new_n26687 = new_n26686 ^ new_n26659;
  assign new_n26688 = ~new_n26687 & new_n26685;
  assign new_n26689 = new_n26688 ^ new_n26658;
  assign new_n26690 = new_n26665 ^ new_n26628;
  assign new_n26691 = new_n26690 ^ new_n26689;
  assign new_n26692 = new_n26691 ^ new_n26684;
  assign new_n26693 = new_n26685 ^ new_n26672;
  assign new_n26694 = ~new_n26637 & ~new_n26693;
  assign new_n26695 = new_n26694 ^ new_n26656;
  assign new_n26696 = new_n26695 ^ new_n26637;
  assign new_n26697 = new_n26674 ^ new_n26635;
  assign new_n26698 = new_n26697 ^ new_n26659;
  assign new_n26699 = new_n26643 & new_n26698;
  assign new_n26700 = new_n26699 ^ new_n26658;
  assign new_n26701 = new_n26688 ^ new_n26649;
  assign new_n26702 = new_n26701 ^ new_n26700;
  assign new_n26703 = new_n26702 ^ new_n26696;
  assign new_n26704 = ~new_n26692 & new_n26703;
  assign new_n26705 = new_n26674 ^ new_n26620;
  assign new_n26706 = ~new_n26642 & ~new_n26705;
  assign new_n26707 = new_n26706 ^ new_n26620;
  assign new_n26708 = new_n26707 ^ new_n26695;
  assign new_n26709 = new_n26708 ^ new_n26704;
  assign new_n26710 = new_n26709 ^ new_n26671;
  assign new_n26711 = new_n26681 ^ new_n26677;
  assign new_n26712 = new_n26688 ^ new_n26668;
  assign new_n26713 = new_n26712 ^ new_n26711;
  assign new_n26714 = ~new_n26710 & ~new_n26713;
  assign new_n26715 = new_n26714 ^ new_n26704;
  assign new_n26716 = ~new_n26715 & new_n26680;
  assign new_n26717 = new_n26716 ^ new_n26680;
  assign new_n26718 = new_n26717 ^ new_n26714;
  assign new_n26719 = new_n26718 ^ new_n26713;
  assign new_n26720 = ~new_n26719 & new_n26643;
  assign new_n26721 = new_n26717 ^ new_n26692;
  assign new_n26722 = ~new_n26637 & ~new_n26721;
  assign new_n26723 = new_n26722 ^ new_n26720;
  assign new_n26724 = ~new_n26693 & ~new_n26721;
  assign new_n26725 = new_n26724 ^ new_n26723;
  assign new_n26726 = new_n26665 ^ new_n26612;
  assign new_n26727 = new_n26706 ^ new_n26699;
  assign new_n26728 = new_n26727 ^ new_n26712;
  assign new_n26729 = new_n26728 ^ new_n26726;
  assign new_n26730 = new_n26704 ^ new_n26680;
  assign new_n26731 = ~new_n26729 & new_n26730;
  assign new_n26732 = new_n26731 ^ new_n26708;
  assign new_n26733 = new_n26732 ^ new_n26671;
  assign new_n26734 = new_n26716 ^ new_n26704;
  assign new_n26735 = ~new_n26733 & new_n26734;
  assign new_n26736 = new_n26735 ^ new_n26729;
  assign new_n26737 = ~new_n26674 & ~new_n26736;
  assign new_n26738 = new_n26731 ^ new_n26714;
  assign new_n26739 = new_n26708 ^ new_n26679;
  assign new_n26740 = new_n26739 ^ new_n26738;
  assign new_n26741 = ~new_n26740 & new_n26621;
  assign new_n26742 = new_n26665 ^ new_n26635;
  assign new_n26743 = new_n26699 ^ new_n26682;
  assign new_n26744 = new_n26735 ^ new_n26717;
  assign new_n26745 = new_n26744 ^ new_n26743;
  assign new_n26746 = new_n26745 ^ new_n26742;
  assign new_n26747 = new_n26746 ^ new_n26620;
  assign new_n26748 = new_n26731 ^ new_n26673;
  assign new_n26749 = new_n26748 ^ new_n26695;
  assign new_n26750 = new_n26749 ^ new_n26747;
  assign new_n26751 = ~new_n26750 & new_n26685;
  assign new_n26752 = new_n26751 ^ new_n26741;
  assign new_n26753 = ~new_n26719 & new_n26698;
  assign new_n26754 = new_n26753 ^ new_n26752;
  assign new_n26755 = new_n26754 ^ new_n26737;
  assign new_n26756 = new_n26735 ^ new_n26731;
  assign new_n26757 = new_n26756 ^ new_n26703;
  assign new_n26758 = new_n26670 & new_n26757;
  assign new_n26759 = new_n26758 ^ new_n26755;
  assign new_n26760 = new_n26759 ^ new_n26725;
  assign new_n26761 = ~new_n26395 & ~new_n26496;
  assign new_n26762 = ~new_n26474 & new_n26417;
  assign new_n26763 = new_n26762 ^ new_n26761;
  assign new_n26764 = new_n26763 ^ new_n26497;
  assign new_n26765 = new_n26764 ^ new_n26493;
  assign new_n26766 = new_n26765 ^ new_n26760;
  assign new_n26767 = new_n26766 ^ new_n26606;
  assign new_n26768 = new_n24500 ^ new_n24456;
  assign new_n26769 = new_n24895 ^ new_n24550;
  assign new_n26770 = new_n26769 ^ new_n24418;
  assign new_n26771 = new_n26770 ^ new_n26768;
  assign new_n26772 = new_n24550 ^ new_n24546;
  assign new_n26773 = new_n26772 ^ new_n24877;
  assign new_n26774 = new_n26773 ^ new_n23967;
  assign new_n26775 = new_n24575 ^ new_n24529;
  assign new_n26776 = new_n26775 ^ new_n24557;
  assign new_n26777 = new_n26776 ^ new_n26774;
  assign new_n26778 = new_n26777 ^ new_n26771;
  assign new_n26779 = new_n24627 ^ new_n24557;
  assign new_n26780 = new_n26779 ^ new_n24613;
  assign new_n26781 = new_n24885 ^ new_n24513;
  assign new_n26782 = new_n26781 ^ new_n26772;
  assign new_n26783 = new_n26782 ^ new_n26780;
  assign new_n26784 = new_n26772 ^ new_n24485;
  assign new_n26785 = new_n26784 ^ new_n24623;
  assign new_n26786 = new_n24890 ^ new_n24592;
  assign new_n26787 = new_n26786 ^ new_n24467;
  assign new_n26788 = new_n26787 ^ new_n26785;
  assign new_n26789 = new_n26788 ^ new_n26783;
  assign new_n26790 = new_n26789 ^ new_n26778;
  assign new_n26791 = new_n24871 ^ new_n24467;
  assign new_n26792 = new_n26772 ^ new_n24604;
  assign new_n26793 = new_n26792 ^ new_n26791;
  assign new_n26794 = new_n26793 ^ new_n26790;
  assign new_n26795 = new_n24395 ^ new_n24130;
  assign new_n26796 = new_n24529 ^ new_n24524;
  assign new_n26797 = new_n26796 ^ new_n24861;
  assign new_n26798 = new_n26797 ^ new_n26795;
  assign new_n26799 = new_n24841 ^ new_n24418;
  assign new_n26800 = new_n26799 ^ new_n24130;
  assign new_n26801 = new_n24538 ^ new_n24374;
  assign new_n26802 = new_n26801 ^ new_n26800;
  assign new_n26803 = new_n26802 ^ new_n26798;
  assign new_n26804 = new_n26803 ^ new_n26793;
  assign new_n26805 = ~new_n26804 & new_n26788;
  assign new_n26806 = new_n26805 ^ new_n26788;
  assign new_n26807 = new_n24586 ^ new_n24570;
  assign new_n26808 = new_n24903 ^ new_n24613;
  assign new_n26809 = new_n26808 ^ new_n24592;
  assign new_n26810 = new_n26809 ^ new_n26807;
  assign new_n26811 = new_n26810 ^ new_n26789;
  assign new_n26812 = new_n26811 ^ new_n26798;
  assign new_n26813 = new_n26788 ^ new_n26771;
  assign new_n26814 = ~new_n26812 & ~new_n26813;
  assign new_n26815 = new_n26814 ^ new_n26806;
  assign new_n26816 = new_n26810 ^ new_n26771;
  assign new_n26817 = new_n26816 ^ new_n26815;
  assign new_n26818 = new_n26798 ^ new_n26777;
  assign new_n26819 = new_n26818 ^ new_n26816;
  assign new_n26820 = new_n26810 ^ new_n26777;
  assign new_n26821 = ~new_n26820 & new_n26819;
  assign new_n26822 = new_n26811 ^ new_n26802;
  assign new_n26823 = new_n26778 & new_n26822;
  assign new_n26824 = new_n26823 ^ new_n26821;
  assign new_n26825 = new_n26798 ^ new_n26783;
  assign new_n26826 = new_n26825 ^ new_n26824;
  assign new_n26827 = new_n26826 ^ new_n26817;
  assign new_n26828 = new_n26788 ^ new_n26777;
  assign new_n26829 = new_n26828 ^ new_n26816;
  assign new_n26830 = ~new_n26790 & new_n26829;
  assign new_n26831 = new_n26830 ^ new_n26802;
  assign new_n26832 = new_n26831 ^ new_n26790;
  assign new_n26833 = new_n26804 ^ new_n26788;
  assign new_n26834 = new_n26833 ^ new_n26816;
  assign new_n26835 = new_n26794 & new_n26834;
  assign new_n26836 = new_n26835 ^ new_n26810;
  assign new_n26837 = new_n26836 ^ new_n26824;
  assign new_n26838 = new_n26837 ^ new_n26832;
  assign new_n26839 = new_n26827 & new_n26838;
  assign new_n26840 = new_n26803 ^ new_n26790;
  assign new_n26841 = ~new_n26816 & new_n26840;
  assign new_n26842 = new_n26841 ^ new_n26823;
  assign new_n26843 = new_n26842 ^ new_n26812;
  assign new_n26844 = new_n26804 ^ new_n26771;
  assign new_n26845 = new_n26822 ^ new_n26793;
  assign new_n26846 = ~new_n26845 & new_n26844;
  assign new_n26847 = new_n26846 ^ new_n26814;
  assign new_n26848 = new_n26847 ^ new_n26771;
  assign new_n26849 = new_n26848 ^ new_n26843;
  assign new_n26850 = new_n26849 ^ new_n26839;
  assign new_n26851 = new_n26804 ^ new_n26777;
  assign new_n26852 = ~new_n26793 & new_n26851;
  assign new_n26853 = new_n26852 ^ new_n26777;
  assign new_n26854 = new_n26853 ^ new_n26831;
  assign new_n26855 = new_n26854 ^ new_n26839;
  assign new_n26856 = new_n26855 ^ new_n26843;
  assign new_n26857 = new_n26846 ^ new_n26805;
  assign new_n26858 = new_n26841 ^ new_n26821;
  assign new_n26859 = new_n26858 ^ new_n26857;
  assign new_n26860 = ~new_n26856 & ~new_n26859;
  assign new_n26861 = new_n26860 ^ new_n26839;
  assign new_n26862 = ~new_n26861 & new_n26849;
  assign new_n26863 = new_n26862 ^ new_n26860;
  assign new_n26864 = new_n26863 ^ new_n26850;
  assign new_n26865 = new_n26864 ^ new_n26860;
  assign new_n26866 = new_n26865 ^ new_n26859;
  assign new_n26867 = ~new_n26866 & new_n26794;
  assign new_n26868 = new_n26864 ^ new_n26827;
  assign new_n26869 = ~new_n26790 & new_n26868;
  assign new_n26870 = new_n26869 ^ new_n26867;
  assign new_n26871 = new_n26829 & new_n26868;
  assign new_n26872 = new_n26871 ^ new_n26870;
  assign new_n26873 = new_n26798 ^ new_n26771;
  assign new_n26874 = new_n26852 ^ new_n26835;
  assign new_n26875 = new_n26874 ^ new_n26858;
  assign new_n26876 = new_n26875 ^ new_n26873;
  assign new_n26877 = ~new_n26850 & ~new_n26876;
  assign new_n26878 = new_n26877 ^ new_n26854;
  assign new_n26879 = new_n26878 ^ new_n26843;
  assign new_n26880 = ~new_n26863 & ~new_n26879;
  assign new_n26881 = new_n26880 ^ new_n26876;
  assign new_n26882 = ~new_n26881 & new_n26804;
  assign new_n26883 = new_n26877 ^ new_n26860;
  assign new_n26884 = new_n26854 ^ new_n26848;
  assign new_n26885 = new_n26884 ^ new_n26883;
  assign new_n26886 = new_n26778 & new_n26885;
  assign new_n26887 = new_n26798 ^ new_n26788;
  assign new_n26888 = new_n26835 ^ new_n26806;
  assign new_n26889 = new_n26880 ^ new_n26864;
  assign new_n26890 = new_n26889 ^ new_n26888;
  assign new_n26891 = new_n26890 ^ new_n26887;
  assign new_n26892 = new_n26891 ^ new_n26777;
  assign new_n26893 = new_n26877 ^ new_n26814;
  assign new_n26894 = new_n26893 ^ new_n26831;
  assign new_n26895 = new_n26894 ^ new_n26892;
  assign new_n26896 = ~new_n26820 & new_n26895;
  assign new_n26897 = new_n26896 ^ new_n26886;
  assign new_n26898 = ~new_n26866 & new_n26834;
  assign new_n26899 = new_n26898 ^ new_n26897;
  assign new_n26900 = new_n26899 ^ new_n26882;
  assign new_n26901 = new_n26880 ^ new_n26877;
  assign new_n26902 = new_n26901 ^ new_n26838;
  assign new_n26903 = ~new_n26812 & new_n26902;
  assign new_n26904 = new_n26903 ^ new_n26900;
  assign new_n26905 = new_n26904 ^ new_n26872;
  assign new_n26906 = new_n26268 & new_n26328;
  assign new_n26907 = new_n26906 ^ new_n26325;
  assign new_n26908 = new_n26315 ^ new_n26274;
  assign new_n26909 = new_n26265 & new_n26908;
  assign new_n26910 = new_n26292 & new_n26348;
  assign new_n26911 = new_n26910 ^ new_n26909;
  assign new_n26912 = new_n26911 ^ new_n26351;
  assign new_n26913 = new_n26912 ^ new_n26907;
  assign new_n26914 = ~new_n26431 & ~new_n26457;
  assign new_n26915 = new_n26914 ^ new_n26497;
  assign new_n26916 = new_n26462 ^ new_n26435;
  assign new_n26917 = ~new_n26413 & new_n26916;
  assign new_n26918 = new_n26917 ^ new_n26762;
  assign new_n26919 = new_n26918 ^ new_n26492;
  assign new_n26920 = new_n26919 ^ new_n26915;
  assign new_n26921 = new_n26920 ^ new_n26913;
  assign new_n26922 = new_n26921 ^ new_n26905;
  assign new_n26923 = new_n26922 ^ new_n26767;
  assign new_n26924 = new_n26822 & new_n26885;
  assign new_n26925 = new_n26924 ^ new_n26886;
  assign new_n26926 = new_n26860 ^ new_n26771;
  assign new_n26927 = new_n26852 ^ new_n26846;
  assign new_n26928 = new_n26927 ^ new_n26891;
  assign new_n26929 = new_n26928 ^ new_n26926;
  assign new_n26930 = ~new_n26816 & new_n26929;
  assign new_n26931 = ~new_n26813 & new_n26902;
  assign new_n26932 = new_n26860 ^ new_n26849;
  assign new_n26933 = ~new_n26793 & ~new_n26932;
  assign new_n26934 = new_n26933 ^ new_n26869;
  assign new_n26935 = new_n26934 ^ new_n26931;
  assign new_n26936 = new_n26840 & new_n26929;
  assign new_n26937 = ~new_n26879 & new_n26844;
  assign new_n26938 = new_n26937 ^ new_n26936;
  assign new_n26939 = new_n26938 ^ new_n26935;
  assign new_n26940 = new_n26939 ^ new_n26930;
  assign new_n26941 = new_n26940 ^ new_n26925;
  assign new_n26942 = new_n26507 & new_n26584;
  assign new_n26943 = new_n26942 ^ new_n26585;
  assign new_n26944 = new_n26558 ^ new_n24542;
  assign new_n26945 = new_n26550 ^ new_n26521;
  assign new_n26946 = new_n26945 ^ new_n26590;
  assign new_n26947 = new_n26946 ^ new_n26944;
  assign new_n26948 = ~new_n26947 & new_n26509;
  assign new_n26949 = new_n26516 & new_n26601;
  assign new_n26950 = new_n26558 ^ new_n26524;
  assign new_n26951 = new_n24476 & new_n26950;
  assign new_n26952 = new_n26951 ^ new_n26566;
  assign new_n26953 = new_n26952 ^ new_n26949;
  assign new_n26954 = ~new_n26947 & new_n26511;
  assign new_n26955 = new_n26519 & new_n26577;
  assign new_n26956 = new_n26955 ^ new_n26954;
  assign new_n26957 = new_n26956 ^ new_n26953;
  assign new_n26958 = new_n26957 ^ new_n26948;
  assign new_n26959 = new_n26958 ^ new_n26943;
  assign new_n26960 = new_n26959 ^ new_n12482;
  assign new_n26961 = new_n26960 ^ new_n26941;
  assign new_n26962 = new_n26254 & new_n26324;
  assign new_n26963 = new_n26962 ^ new_n26910;
  assign new_n26964 = new_n26963 ^ new_n26325;
  assign new_n26965 = new_n26964 ^ new_n26352;
  assign new_n26966 = new_n26965 ^ new_n26765;
  assign new_n26967 = ~new_n26740 & new_n26657;
  assign new_n26968 = new_n26967 ^ new_n26741;
  assign new_n26969 = new_n26714 ^ new_n26612;
  assign new_n26970 = new_n26706 ^ new_n26677;
  assign new_n26971 = new_n26970 ^ new_n26746;
  assign new_n26972 = new_n26971 ^ new_n26969;
  assign new_n26973 = new_n26659 & new_n26972;
  assign new_n26974 = ~new_n26672 & new_n26757;
  assign new_n26975 = new_n26714 ^ new_n26680;
  assign new_n26976 = ~new_n26642 & new_n26975;
  assign new_n26977 = new_n26976 ^ new_n26722;
  assign new_n26978 = new_n26977 ^ new_n26974;
  assign new_n26979 = ~new_n26667 & new_n26972;
  assign new_n26980 = ~new_n26675 & ~new_n26733;
  assign new_n26981 = new_n26980 ^ new_n26979;
  assign new_n26982 = new_n26981 ^ new_n26978;
  assign new_n26983 = new_n26982 ^ new_n26973;
  assign new_n26984 = new_n26983 ^ new_n26968;
  assign new_n26985 = new_n26498 ^ new_n26489;
  assign new_n26986 = new_n26462 ^ new_n26385;
  assign new_n26987 = new_n26432 ^ new_n26420;
  assign new_n26988 = new_n26987 ^ new_n26480;
  assign new_n26989 = new_n26988 ^ new_n26986;
  assign new_n26990 = new_n26387 & new_n26989;
  assign new_n26991 = new_n26917 ^ new_n26761;
  assign new_n26992 = ~new_n26428 & new_n26468;
  assign new_n26993 = new_n26992 ^ new_n26991;
  assign new_n26994 = ~new_n26430 & ~new_n26457;
  assign new_n26995 = ~new_n26402 & new_n26989;
  assign new_n26996 = new_n26995 ^ new_n26994;
  assign new_n26997 = new_n26996 ^ new_n26993;
  assign new_n26998 = new_n26997 ^ new_n26990;
  assign new_n26999 = new_n26998 ^ new_n26985;
  assign new_n27000 = new_n26999 ^ new_n26984;
  assign new_n27001 = new_n27000 ^ new_n26966;
  assign new_n27002 = new_n27001 ^ new_n26961;
  assign new_n27003 = new_n27002 ^ new_n26923;
  assign new_n27004 = new_n26270 & new_n26331;
  assign new_n27005 = new_n26315 ^ new_n26239;
  assign new_n27006 = new_n26303 ^ new_n26269;
  assign new_n27007 = new_n27006 ^ new_n26340;
  assign new_n27008 = new_n27007 ^ new_n27005;
  assign new_n27009 = new_n26255 & new_n27008;
  assign new_n27010 = new_n27009 ^ new_n27004;
  assign new_n27011 = new_n26353 ^ new_n26334;
  assign new_n27012 = new_n26293 & new_n26333;
  assign new_n27013 = new_n27012 ^ new_n26906;
  assign new_n27014 = new_n27013 ^ new_n26346;
  assign new_n27015 = new_n27014 ^ new_n27011;
  assign new_n27016 = new_n27015 ^ new_n27010;
  assign new_n27017 = ~new_n26705 & new_n26975;
  assign new_n27018 = ~new_n26687 & ~new_n26750;
  assign new_n27019 = new_n27018 ^ new_n26759;
  assign new_n27020 = new_n27019 ^ new_n27017;
  assign new_n27021 = new_n27020 ^ new_n26982;
  assign new_n27022 = ~new_n26932 & new_n26851;
  assign new_n27023 = new_n26819 & new_n26895;
  assign new_n27024 = new_n27023 ^ new_n26904;
  assign new_n27025 = new_n27024 ^ new_n27022;
  assign new_n27026 = new_n27025 ^ new_n26939;
  assign new_n27027 = new_n27026 ^ new_n27021;
  assign new_n27028 = new_n27027 ^ new_n27016;
  assign new_n27029 = ~new_n26419 & new_n26916;
  assign new_n27030 = new_n27029 ^ new_n26495;
  assign new_n27031 = new_n27030 ^ new_n26997;
  assign new_n27032 = new_n26549 & new_n26950;
  assign new_n27033 = ~new_n26594 & new_n26530;
  assign new_n27034 = new_n27033 ^ new_n26603;
  assign new_n27035 = new_n27034 ^ new_n27032;
  assign new_n27036 = new_n27035 ^ new_n26957;
  assign new_n27037 = new_n27036 ^ new_n12595;
  assign new_n27038 = new_n27037 ^ new_n27031;
  assign new_n27039 = new_n26995 ^ new_n26992;
  assign new_n27040 = new_n26494 ^ new_n26471;
  assign new_n27041 = ~new_n26470 & new_n26415;
  assign new_n27042 = new_n27041 ^ new_n26914;
  assign new_n27043 = new_n27042 ^ new_n26490;
  assign new_n27044 = new_n27043 ^ new_n27040;
  assign new_n27045 = new_n27044 ^ new_n27039;
  assign new_n27046 = new_n27045 ^ new_n27038;
  assign new_n27047 = new_n27046 ^ new_n27028;
  assign new_n27048 = new_n26924 ^ new_n26871;
  assign new_n27049 = new_n27048 ^ new_n27024;
  assign new_n27050 = new_n26942 ^ new_n26568;
  assign new_n27051 = new_n27050 ^ new_n27034;
  assign new_n27052 = new_n27051 ^ new_n12645;
  assign new_n27053 = new_n27052 ^ new_n27049;
  assign new_n27054 = new_n26498 ^ new_n26494;
  assign new_n27055 = new_n26764 ^ new_n26491;
  assign new_n27056 = new_n27055 ^ new_n27054;
  assign new_n27057 = new_n26353 ^ new_n26319;
  assign new_n27058 = new_n26964 ^ new_n26350;
  assign new_n27059 = new_n27058 ^ new_n27057;
  assign new_n27060 = new_n27059 ^ new_n27056;
  assign new_n27061 = new_n26967 ^ new_n26724;
  assign new_n27062 = new_n27061 ^ new_n27019;
  assign new_n27063 = new_n27062 ^ new_n26500;
  assign new_n27064 = new_n27063 ^ new_n27060;
  assign new_n27065 = new_n27064 ^ new_n27053;
  assign new_n27066 = new_n27065 ^ new_n27047;
  assign new_n27067 = new_n27066 ^ new_n27003;
  assign new_n27068 = new_n26962 ^ new_n26909;
  assign new_n27069 = new_n27068 ^ new_n27004;
  assign new_n27070 = new_n27069 ^ new_n26332;
  assign new_n27071 = new_n27070 ^ new_n27014;
  assign new_n27072 = new_n27071 ^ new_n26501;
  assign new_n27073 = new_n26979 ^ new_n26974;
  assign new_n27074 = new_n27018 ^ new_n26737;
  assign new_n27075 = ~new_n26676 & ~new_n26733;
  assign new_n27076 = ~new_n26736 & new_n26697;
  assign new_n27077 = new_n27076 ^ new_n27075;
  assign new_n27078 = new_n27077 ^ new_n26752;
  assign new_n27079 = new_n27078 ^ new_n27074;
  assign new_n27080 = new_n27079 ^ new_n27073;
  assign new_n27081 = new_n26936 ^ new_n26931;
  assign new_n27082 = new_n27023 ^ new_n26882;
  assign new_n27083 = ~new_n26845 & ~new_n26879;
  assign new_n27084 = ~new_n26833 & ~new_n26881;
  assign new_n27085 = new_n27084 ^ new_n27083;
  assign new_n27086 = new_n27085 ^ new_n26897;
  assign new_n27087 = new_n27086 ^ new_n27082;
  assign new_n27088 = new_n27087 ^ new_n27081;
  assign new_n27089 = new_n27088 ^ new_n27080;
  assign new_n27090 = new_n27089 ^ new_n27072;
  assign new_n27091 = new_n26954 ^ new_n26949;
  assign new_n27092 = new_n27033 ^ new_n26581;
  assign new_n27093 = new_n26520 & new_n26577;
  assign new_n27094 = new_n26542 & new_n26580;
  assign new_n27095 = new_n27094 ^ new_n27093;
  assign new_n27096 = new_n27095 ^ new_n26596;
  assign new_n27097 = new_n27096 ^ new_n27092;
  assign new_n27098 = new_n27097 ^ new_n27091;
  assign new_n27099 = new_n27098 ^ new_n12566;
  assign new_n27100 = new_n27099 ^ new_n27045;
  assign new_n27101 = new_n26993 ^ new_n26469;
  assign new_n27102 = new_n27101 ^ new_n27043;
  assign new_n27103 = new_n27102 ^ new_n27100;
  assign new_n27104 = new_n27103 ^ new_n27090;
  assign new_n27105 = new_n27104 ^ new_n27002;
  assign new_n27106 = new_n27023 ^ new_n26924;
  assign new_n27107 = new_n26899 ^ new_n26872;
  assign new_n27108 = new_n27107 ^ new_n27106;
  assign new_n27109 = new_n27033 ^ new_n26942;
  assign new_n27110 = new_n26598 ^ new_n26569;
  assign new_n27111 = new_n27110 ^ new_n27109;
  assign new_n27112 = new_n27111 ^ new_n12518;
  assign new_n27113 = new_n27112 ^ new_n27108;
  assign new_n27114 = new_n26335 ^ new_n26319;
  assign new_n27115 = new_n26267 & new_n26328;
  assign new_n27116 = new_n27115 ^ new_n27009;
  assign new_n27117 = new_n27116 ^ new_n27069;
  assign new_n27118 = new_n26240 & new_n27008;
  assign new_n27119 = new_n27118 ^ new_n27117;
  assign new_n27120 = new_n27119 ^ new_n27114;
  assign new_n27121 = new_n27120 ^ new_n26999;
  assign new_n27122 = new_n27018 ^ new_n26967;
  assign new_n27123 = new_n26754 ^ new_n26725;
  assign new_n27124 = new_n27123 ^ new_n27122;
  assign new_n27125 = new_n27124 ^ new_n27056;
  assign new_n27126 = new_n27125 ^ new_n27121;
  assign new_n27127 = new_n27126 ^ new_n27113;
  assign new_n27128 = new_n27127 ^ new_n27002;
  assign new_n27129 = new_n26953 ^ new_n26602;
  assign new_n27130 = new_n27129 ^ new_n27096;
  assign new_n27131 = new_n27130 ^ new_n12547;
  assign new_n27132 = new_n27131 ^ new_n27102;
  assign new_n27133 = new_n26978 ^ new_n26758;
  assign new_n27134 = new_n27133 ^ new_n27078;
  assign new_n27135 = new_n26935 ^ new_n26903;
  assign new_n27136 = new_n27135 ^ new_n27086;
  assign new_n27137 = new_n27136 ^ new_n27134;
  assign new_n27138 = new_n27137 ^ new_n26501;
  assign new_n27139 = new_n27138 ^ new_n27132;
  assign new_n27140 = new_n27139 ^ new_n27128;
  assign new_n27141 = new_n27104 & new_n27140;
  assign new_n27142 = new_n27141 ^ new_n27104;
  assign new_n27143 = new_n27140 ^ new_n27104;
  assign new_n27144 = new_n27143 ^ new_n27066;
  assign new_n27145 = new_n27065 ^ new_n26923;
  assign new_n27146 = new_n26302 & new_n26908;
  assign new_n27147 = new_n27146 ^ new_n26354;
  assign new_n27148 = new_n27147 ^ new_n27117;
  assign new_n27149 = new_n27031 ^ new_n26920;
  assign new_n27150 = new_n27149 ^ new_n27148;
  assign new_n27151 = new_n27075 ^ new_n26724;
  assign new_n27152 = new_n26976 ^ new_n26720;
  assign new_n27153 = new_n27152 ^ new_n26755;
  assign new_n27154 = new_n27153 ^ new_n27151;
  assign new_n27155 = new_n27083 ^ new_n26871;
  assign new_n27156 = new_n26933 ^ new_n26867;
  assign new_n27157 = new_n27156 ^ new_n26900;
  assign new_n27158 = new_n27157 ^ new_n27155;
  assign new_n27159 = new_n27158 ^ new_n27154;
  assign new_n27160 = new_n27093 ^ new_n26568;
  assign new_n27161 = new_n26951 ^ new_n26564;
  assign new_n27162 = new_n27161 ^ new_n26599;
  assign new_n27163 = new_n27162 ^ new_n27160;
  assign new_n27164 = new_n27163 ^ new_n12627;
  assign new_n27165 = new_n27164 ^ new_n26501;
  assign new_n27166 = new_n27165 ^ new_n27159;
  assign new_n27167 = new_n27166 ^ new_n27150;
  assign new_n27168 = new_n27167 ^ new_n27104;
  assign new_n27169 = new_n27168 ^ new_n27145;
  assign new_n27170 = new_n27169 ^ new_n27139;
  assign new_n27171 = new_n27144 & new_n27170;
  assign new_n27172 = new_n27171 ^ new_n27142;
  assign new_n27173 = new_n27104 ^ new_n27065;
  assign new_n27174 = new_n27047 ^ new_n26923;
  assign new_n27175 = new_n27174 ^ new_n27173;
  assign new_n27176 = ~new_n27169 & ~new_n27175;
  assign new_n27177 = new_n27176 ^ new_n27127;
  assign new_n27178 = ~new_n27128 & ~new_n27139;
  assign new_n27179 = new_n26923 & new_n27139;
  assign new_n27180 = new_n27179 ^ new_n27178;
  assign new_n27181 = new_n27180 ^ new_n27177;
  assign new_n27182 = new_n27065 ^ new_n27002;
  assign new_n27183 = new_n27169 ^ new_n27128;
  assign new_n27184 = ~new_n27183 & new_n27066;
  assign new_n27185 = ~new_n27067 & new_n27174;
  assign new_n27186 = new_n27185 ^ new_n27184;
  assign new_n27187 = new_n27180 ^ new_n26923;
  assign new_n27188 = new_n27187 ^ new_n27171;
  assign new_n27189 = new_n27188 ^ new_n27186;
  assign new_n27190 = new_n27189 ^ new_n27182;
  assign new_n27191 = new_n27168 ^ new_n27047;
  assign new_n27192 = new_n27191 ^ new_n27127;
  assign new_n27193 = new_n27145 & new_n27192;
  assign new_n27194 = new_n27193 ^ new_n27184;
  assign new_n27195 = new_n27191 ^ new_n27002;
  assign new_n27196 = new_n27195 ^ new_n27194;
  assign new_n27197 = ~new_n27173 & new_n27195;
  assign new_n27198 = new_n27140 ^ new_n27065;
  assign new_n27199 = new_n27192 ^ new_n27139;
  assign new_n27200 = ~new_n27198 & ~new_n27199;
  assign new_n27201 = new_n27200 ^ new_n27197;
  assign new_n27202 = new_n27201 ^ new_n27065;
  assign new_n27203 = new_n27202 ^ new_n27196;
  assign new_n27204 = new_n27197 ^ new_n27142;
  assign new_n27205 = new_n27204 ^ new_n27066;
  assign new_n27206 = new_n27193 ^ new_n27185;
  assign new_n27207 = new_n27167 ^ new_n27002;
  assign new_n27208 = new_n27207 ^ new_n27206;
  assign new_n27209 = new_n27208 ^ new_n27205;
  assign new_n27210 = new_n27177 ^ new_n27169;
  assign new_n27211 = new_n27206 ^ new_n27171;
  assign new_n27212 = new_n27211 ^ new_n27047;
  assign new_n27213 = new_n27212 ^ new_n27210;
  assign new_n27214 = ~new_n27209 & new_n27213;
  assign new_n27215 = new_n27214 ^ new_n27203;
  assign new_n27216 = ~new_n27190 & new_n27215;
  assign new_n27217 = new_n27216 ^ new_n27181;
  assign new_n27218 = new_n27217 ^ new_n27196;
  assign new_n27219 = new_n27214 ^ new_n27181;
  assign new_n27220 = new_n27219 ^ new_n27196;
  assign new_n27221 = new_n27200 ^ new_n27141;
  assign new_n27222 = new_n27221 ^ new_n27186;
  assign new_n27223 = ~new_n27220 & ~new_n27222;
  assign new_n27224 = new_n27223 ^ new_n27214;
  assign new_n27225 = new_n27203 & new_n27224;
  assign new_n27226 = new_n27225 ^ new_n27215;
  assign new_n27227 = ~new_n27218 & new_n27226;
  assign new_n27228 = new_n27227 ^ new_n27225;
  assign new_n27229 = new_n27228 ^ new_n27172;
  assign new_n27230 = new_n27229 ^ new_n27105;
  assign new_n27231 = new_n27230 ^ new_n26923;
  assign new_n27232 = new_n27216 ^ new_n27197;
  assign new_n27233 = new_n27232 ^ new_n27177;
  assign new_n27234 = new_n27233 ^ new_n27231;
  assign new_n27235 = ~new_n27067 & ~new_n27234;
  assign new_n27236 = new_n27223 ^ new_n27216;
  assign new_n27237 = new_n27202 ^ new_n27181;
  assign new_n27238 = new_n27237 ^ new_n27236;
  assign new_n27239 = ~new_n27238 & new_n27192;
  assign new_n27240 = new_n27239 ^ new_n27235;
  assign new_n27241 = new_n27225 ^ new_n27223;
  assign new_n27242 = new_n27241 ^ new_n27222;
  assign new_n27243 = ~new_n27242 & new_n27170;
  assign new_n27244 = new_n27225 ^ new_n27209;
  assign new_n27245 = ~new_n27169 & ~new_n27244;
  assign new_n27246 = new_n27245 ^ new_n27243;
  assign new_n27247 = ~new_n27175 & ~new_n27244;
  assign new_n27248 = new_n27247 ^ new_n27246;
  assign new_n27249 = ~new_n27242 & new_n27144;
  assign new_n27250 = ~new_n27234 & new_n27174;
  assign new_n27251 = ~new_n27238 & new_n27145;
  assign new_n27252 = new_n27251 ^ new_n27250;
  assign new_n27253 = new_n27252 ^ new_n27249;
  assign new_n27254 = new_n27253 ^ new_n27248;
  assign new_n27255 = new_n27254 ^ new_n27240;
  assign new_n27256 = new_n22301 ^ new_n21071;
  assign new_n27257 = new_n27256 ^ new_n22267;
  assign new_n27258 = new_n24894 ^ new_n17679;
  assign new_n27259 = new_n27258 ^ new_n22288;
  assign new_n27260 = new_n27259 ^ new_n22450;
  assign new_n27261 = new_n27260 ^ new_n27257;
  assign new_n27262 = new_n24876 ^ new_n18772;
  assign new_n27263 = new_n22431 ^ new_n22306;
  assign new_n27264 = new_n27263 ^ new_n27262;
  assign new_n27265 = new_n22288 ^ new_n20011;
  assign new_n27266 = new_n27265 ^ new_n27264;
  assign new_n27267 = new_n22427 ^ new_n22379;
  assign new_n27268 = new_n27267 ^ new_n22385;
  assign new_n27269 = new_n27268 ^ new_n27266;
  assign new_n27270 = new_n27269 ^ new_n27261;
  assign new_n27271 = new_n24884 ^ new_n18794;
  assign new_n27272 = new_n27271 ^ new_n27265;
  assign new_n27273 = new_n22422 ^ new_n22375;
  assign new_n27274 = new_n27273 ^ new_n27272;
  assign new_n27275 = new_n22397 ^ new_n22385;
  assign new_n27276 = new_n27275 ^ new_n22466;
  assign new_n27277 = new_n27276 ^ new_n27274;
  assign new_n27278 = new_n27265 ^ new_n19999;
  assign new_n27279 = new_n22476 ^ new_n19989;
  assign new_n27280 = new_n27279 ^ new_n27278;
  assign new_n27281 = new_n24889 ^ new_n18635;
  assign new_n27282 = new_n27281 ^ new_n22367;
  assign new_n27283 = new_n27282 ^ new_n22244;
  assign new_n27284 = new_n27283 ^ new_n27280;
  assign new_n27285 = new_n27284 ^ new_n27277;
  assign new_n27286 = new_n27285 ^ new_n27270;
  assign new_n27287 = new_n24870 ^ new_n18824;
  assign new_n27288 = new_n27287 ^ new_n22365;
  assign new_n27289 = new_n22367 ^ new_n21199;
  assign new_n27290 = new_n27289 ^ new_n27265;
  assign new_n27291 = new_n27290 ^ new_n27288;
  assign new_n27292 = new_n27291 ^ new_n27286;
  assign new_n27293 = new_n24902 ^ new_n18671;
  assign new_n27294 = new_n27293 ^ new_n22466;
  assign new_n27295 = new_n22462 ^ new_n22408;
  assign new_n27296 = new_n27295 ^ new_n19990;
  assign new_n27297 = new_n27296 ^ new_n27294;
  assign new_n27298 = new_n27297 ^ new_n27285;
  assign new_n27299 = new_n24840 ^ new_n18766;
  assign new_n27300 = new_n27299 ^ new_n22450;
  assign new_n27301 = new_n27300 ^ new_n22342;
  assign new_n27302 = new_n22454 ^ new_n22273;
  assign new_n27303 = new_n27302 ^ new_n22315;
  assign new_n27304 = new_n27303 ^ new_n27301;
  assign new_n27305 = new_n27304 ^ new_n27298;
  assign new_n27306 = ~new_n27270 & new_n27305;
  assign new_n27307 = new_n27297 ^ new_n27261;
  assign new_n27308 = new_n24860 ^ new_n18719;
  assign new_n27309 = new_n27308 ^ new_n22428;
  assign new_n27310 = new_n22440 ^ new_n22355;
  assign new_n27311 = new_n27310 ^ new_n22342;
  assign new_n27312 = new_n27311 ^ new_n27309;
  assign new_n27313 = new_n27312 ^ new_n27304;
  assign new_n27314 = new_n27313 ^ new_n27286;
  assign new_n27315 = ~new_n27307 & ~new_n27314;
  assign new_n27316 = new_n27315 ^ new_n27306;
  assign new_n27317 = new_n27312 ^ new_n27298;
  assign new_n27318 = new_n27317 ^ new_n27316;
  assign new_n27319 = new_n27284 ^ new_n27261;
  assign new_n27320 = ~new_n27319 & new_n27317;
  assign new_n27321 = new_n27313 ^ new_n27291;
  assign new_n27322 = new_n27321 ^ new_n27261;
  assign new_n27323 = new_n27305 ^ new_n27291;
  assign new_n27324 = ~new_n27322 & ~new_n27323;
  assign new_n27325 = new_n27324 ^ new_n27320;
  assign new_n27326 = new_n27325 ^ new_n27261;
  assign new_n27327 = new_n27326 ^ new_n27318;
  assign new_n27328 = new_n27284 & new_n27321;
  assign new_n27329 = new_n27328 ^ new_n27284;
  assign new_n27330 = new_n27329 ^ new_n27320;
  assign new_n27331 = new_n27330 ^ new_n27307;
  assign new_n27332 = new_n27312 ^ new_n27269;
  assign new_n27333 = new_n27332 ^ new_n27307;
  assign new_n27334 = new_n27297 ^ new_n27269;
  assign new_n27335 = ~new_n27333 & new_n27334;
  assign new_n27336 = new_n27335 ^ new_n27306;
  assign new_n27337 = new_n27312 ^ new_n27277;
  assign new_n27338 = new_n27337 ^ new_n27336;
  assign new_n27339 = new_n27338 ^ new_n27331;
  assign new_n27340 = new_n27284 ^ new_n27269;
  assign new_n27341 = new_n27340 ^ new_n27307;
  assign new_n27342 = ~new_n27286 & ~new_n27341;
  assign new_n27343 = new_n27342 ^ new_n27304;
  assign new_n27344 = new_n27343 ^ new_n27286;
  assign new_n27345 = new_n27321 ^ new_n27284;
  assign new_n27346 = new_n27345 ^ new_n27307;
  assign new_n27347 = ~new_n27346 & new_n27292;
  assign new_n27348 = new_n27347 ^ new_n27297;
  assign new_n27349 = new_n27348 ^ new_n27336;
  assign new_n27350 = new_n27349 ^ new_n27344;
  assign new_n27351 = ~new_n27339 & ~new_n27350;
  assign new_n27352 = new_n27321 ^ new_n27269;
  assign new_n27353 = ~new_n27291 & new_n27352;
  assign new_n27354 = new_n27353 ^ new_n27269;
  assign new_n27355 = new_n27354 ^ new_n27343;
  assign new_n27356 = new_n27355 ^ new_n27351;
  assign new_n27357 = new_n27356 ^ new_n27318;
  assign new_n27358 = new_n27328 ^ new_n27324;
  assign new_n27359 = new_n27335 ^ new_n27315;
  assign new_n27360 = new_n27359 ^ new_n27358;
  assign new_n27361 = ~new_n27360 & new_n27357;
  assign new_n27362 = new_n27361 ^ new_n27351;
  assign new_n27363 = ~new_n27362 & new_n27327;
  assign new_n27364 = new_n27363 ^ new_n27327;
  assign new_n27365 = new_n27364 ^ new_n27361;
  assign new_n27366 = new_n27365 ^ new_n27360;
  assign new_n27367 = ~new_n27366 & new_n27292;
  assign new_n27368 = new_n27364 ^ new_n27339;
  assign new_n27369 = ~new_n27286 & ~new_n27368;
  assign new_n27370 = new_n27369 ^ new_n27367;
  assign new_n27371 = ~new_n27341 & ~new_n27368;
  assign new_n27372 = new_n27371 ^ new_n27370;
  assign new_n27373 = new_n27312 ^ new_n27261;
  assign new_n27374 = new_n27353 ^ new_n27347;
  assign new_n27375 = new_n27374 ^ new_n27359;
  assign new_n27376 = new_n27375 ^ new_n27373;
  assign new_n27377 = new_n27351 ^ new_n27327;
  assign new_n27378 = ~new_n27376 & new_n27377;
  assign new_n27379 = new_n27378 ^ new_n27355;
  assign new_n27380 = new_n27379 ^ new_n27318;
  assign new_n27381 = new_n27363 ^ new_n27351;
  assign new_n27382 = new_n27380 & new_n27381;
  assign new_n27383 = new_n27382 ^ new_n27376;
  assign new_n27384 = ~new_n27321 & ~new_n27383;
  assign new_n27385 = new_n27378 ^ new_n27361;
  assign new_n27386 = new_n27355 ^ new_n27326;
  assign new_n27387 = new_n27386 ^ new_n27385;
  assign new_n27388 = ~new_n27270 & new_n27387;
  assign new_n27389 = new_n27312 ^ new_n27284;
  assign new_n27390 = new_n27347 ^ new_n27329;
  assign new_n27391 = new_n27382 ^ new_n27364;
  assign new_n27392 = new_n27391 ^ new_n27390;
  assign new_n27393 = new_n27392 ^ new_n27389;
  assign new_n27394 = new_n27393 ^ new_n27269;
  assign new_n27395 = new_n27378 ^ new_n27320;
  assign new_n27396 = new_n27395 ^ new_n27343;
  assign new_n27397 = new_n27396 ^ new_n27394;
  assign new_n27398 = new_n27334 & new_n27397;
  assign new_n27399 = new_n27398 ^ new_n27388;
  assign new_n27400 = ~new_n27346 & ~new_n27366;
  assign new_n27401 = new_n27400 ^ new_n27399;
  assign new_n27402 = new_n27401 ^ new_n27384;
  assign new_n27403 = new_n27382 ^ new_n27378;
  assign new_n27404 = new_n27403 ^ new_n27350;
  assign new_n27405 = ~new_n27404 & new_n27317;
  assign new_n27406 = new_n27405 ^ new_n27402;
  assign new_n27407 = new_n27406 ^ new_n27372;
  assign new_n27408 = new_n24550 ^ new_n24499;
  assign new_n27409 = new_n27408 ^ new_n24399;
  assign new_n27410 = new_n22259 ^ new_n13967;
  assign new_n27411 = new_n27410 ^ new_n24546;
  assign new_n27412 = new_n27411 ^ new_n24456;
  assign new_n27413 = new_n27412 ^ new_n27409;
  assign new_n27414 = new_n24529 ^ new_n23806;
  assign new_n27415 = new_n27414 ^ new_n24547;
  assign new_n27416 = new_n22415 ^ new_n13961;
  assign new_n27417 = new_n27416 ^ new_n24524;
  assign new_n27418 = new_n27417 ^ new_n24576;
  assign new_n27419 = new_n27418 ^ new_n27415;
  assign new_n27420 = new_n27419 ^ new_n27413;
  assign new_n27421 = new_n24586 ^ new_n24547;
  assign new_n27422 = new_n27421 ^ new_n24492;
  assign new_n27423 = new_n21185 ^ new_n13965;
  assign new_n27424 = new_n27423 ^ new_n24622;
  assign new_n27425 = new_n27424 ^ new_n24592;
  assign new_n27426 = new_n27425 ^ new_n27422;
  assign new_n27427 = new_n22391 ^ new_n13972;
  assign new_n27428 = new_n27427 ^ new_n24547;
  assign new_n27429 = new_n27428 ^ new_n24628;
  assign new_n27430 = new_n24557 ^ new_n24508;
  assign new_n27431 = new_n27430 ^ new_n24575;
  assign new_n27432 = new_n27431 ^ new_n27429;
  assign new_n27433 = new_n27432 ^ new_n27426;
  assign new_n27434 = new_n27433 ^ new_n27420;
  assign new_n27435 = new_n24537 ^ new_n24418;
  assign new_n27436 = new_n27435 ^ new_n23985;
  assign new_n27437 = new_n22445 ^ new_n13956;
  assign new_n27438 = new_n27437 ^ new_n24456;
  assign new_n27439 = new_n27438 ^ new_n24374;
  assign new_n27440 = new_n27439 ^ new_n27436;
  assign new_n27441 = new_n22470 ^ new_n13968;
  assign new_n27442 = new_n27441 ^ new_n24587;
  assign new_n27443 = new_n24627 ^ new_n24566;
  assign new_n27444 = new_n27443 ^ new_n24613;
  assign new_n27445 = new_n27444 ^ new_n27442;
  assign new_n27446 = new_n27445 ^ new_n27433;
  assign new_n27447 = new_n27446 ^ new_n27440;
  assign new_n27448 = new_n27420 & new_n27447;
  assign new_n27449 = new_n27445 ^ new_n27413;
  assign new_n27450 = new_n24394 ^ new_n24130;
  assign new_n27451 = new_n27450 ^ new_n24374;
  assign new_n27452 = new_n22328 ^ new_n13957;
  assign new_n27453 = new_n27452 ^ new_n24525;
  assign new_n27454 = new_n27453 ^ new_n27451;
  assign new_n27455 = new_n27454 ^ new_n27440;
  assign new_n27456 = new_n27455 ^ new_n27434;
  assign new_n27457 = ~new_n27456 & new_n27449;
  assign new_n27458 = new_n27457 ^ new_n27448;
  assign new_n27459 = new_n27454 ^ new_n27446;
  assign new_n27460 = new_n27459 ^ new_n27458;
  assign new_n27461 = new_n27426 ^ new_n27413;
  assign new_n27462 = ~new_n27461 & new_n27459;
  assign new_n27463 = new_n24547 ^ new_n24485;
  assign new_n27464 = new_n22360 ^ new_n13959;
  assign new_n27465 = new_n27464 ^ new_n24603;
  assign new_n27466 = new_n27465 ^ new_n24467;
  assign new_n27467 = new_n27466 ^ new_n27463;
  assign new_n27468 = new_n27467 ^ new_n27455;
  assign new_n27469 = new_n27468 ^ new_n27413;
  assign new_n27470 = new_n27467 ^ new_n27447;
  assign new_n27471 = ~new_n27469 & ~new_n27470;
  assign new_n27472 = new_n27471 ^ new_n27462;
  assign new_n27473 = new_n27472 ^ new_n27413;
  assign new_n27474 = new_n27473 ^ new_n27460;
  assign new_n27475 = new_n27426 & new_n27468;
  assign new_n27476 = new_n27475 ^ new_n27426;
  assign new_n27477 = new_n27476 ^ new_n27462;
  assign new_n27478 = new_n27477 ^ new_n27449;
  assign new_n27479 = new_n27454 ^ new_n27419;
  assign new_n27480 = new_n27479 ^ new_n27449;
  assign new_n27481 = new_n27445 ^ new_n27419;
  assign new_n27482 = ~new_n27480 & new_n27481;
  assign new_n27483 = new_n27482 ^ new_n27448;
  assign new_n27484 = new_n27454 ^ new_n27432;
  assign new_n27485 = new_n27484 ^ new_n27483;
  assign new_n27486 = new_n27485 ^ new_n27478;
  assign new_n27487 = new_n27426 ^ new_n27419;
  assign new_n27488 = new_n27487 ^ new_n27449;
  assign new_n27489 = ~new_n27434 & ~new_n27488;
  assign new_n27490 = new_n27489 ^ new_n27440;
  assign new_n27491 = new_n27490 ^ new_n27434;
  assign new_n27492 = new_n27468 ^ new_n27426;
  assign new_n27493 = new_n27492 ^ new_n27449;
  assign new_n27494 = new_n27467 ^ new_n27434;
  assign new_n27495 = new_n27493 & new_n27494;
  assign new_n27496 = new_n27495 ^ new_n27483;
  assign new_n27497 = new_n27496 ^ new_n27445;
  assign new_n27498 = new_n27497 ^ new_n27491;
  assign new_n27499 = ~new_n27486 & new_n27498;
  assign new_n27500 = new_n27468 ^ new_n27419;
  assign new_n27501 = ~new_n27467 & ~new_n27500;
  assign new_n27502 = new_n27501 ^ new_n27419;
  assign new_n27503 = new_n27502 ^ new_n27490;
  assign new_n27504 = new_n27503 ^ new_n27499;
  assign new_n27505 = new_n27504 ^ new_n27460;
  assign new_n27506 = new_n27475 ^ new_n27471;
  assign new_n27507 = new_n27482 ^ new_n27457;
  assign new_n27508 = new_n27507 ^ new_n27506;
  assign new_n27509 = ~new_n27505 & ~new_n27508;
  assign new_n27510 = new_n27509 ^ new_n27499;
  assign new_n27511 = ~new_n27510 & new_n27474;
  assign new_n27512 = new_n27511 ^ new_n27474;
  assign new_n27513 = new_n27512 ^ new_n27486;
  assign new_n27514 = ~new_n27434 & ~new_n27513;
  assign new_n27515 = new_n27512 ^ new_n27509;
  assign new_n27516 = new_n27515 ^ new_n27508;
  assign new_n27517 = ~new_n27516 & new_n27494;
  assign new_n27518 = new_n27517 ^ new_n27514;
  assign new_n27519 = ~new_n27488 & ~new_n27513;
  assign new_n27520 = new_n27519 ^ new_n27518;
  assign new_n27521 = new_n27454 ^ new_n27413;
  assign new_n27522 = new_n27501 ^ new_n27495;
  assign new_n27523 = new_n27522 ^ new_n27507;
  assign new_n27524 = new_n27523 ^ new_n27521;
  assign new_n27525 = new_n27499 ^ new_n27474;
  assign new_n27526 = ~new_n27524 & new_n27525;
  assign new_n27527 = new_n27526 ^ new_n27503;
  assign new_n27528 = new_n27527 ^ new_n27460;
  assign new_n27529 = new_n27511 ^ new_n27499;
  assign new_n27530 = ~new_n27528 & new_n27529;
  assign new_n27531 = new_n27530 ^ new_n27526;
  assign new_n27532 = new_n27531 ^ new_n27498;
  assign new_n27533 = new_n27459 & new_n27532;
  assign new_n27534 = new_n27530 ^ new_n27524;
  assign new_n27535 = ~new_n27468 & ~new_n27534;
  assign new_n27536 = new_n27454 ^ new_n27426;
  assign new_n27537 = new_n27495 ^ new_n27476;
  assign new_n27538 = new_n27530 ^ new_n27512;
  assign new_n27539 = new_n27538 ^ new_n27537;
  assign new_n27540 = new_n27539 ^ new_n27536;
  assign new_n27541 = new_n27540 ^ new_n27419;
  assign new_n27542 = new_n27526 ^ new_n27462;
  assign new_n27543 = new_n27542 ^ new_n27490;
  assign new_n27544 = new_n27543 ^ new_n27541;
  assign new_n27545 = ~new_n27544 & new_n27481;
  assign new_n27546 = new_n27526 ^ new_n27509;
  assign new_n27547 = new_n27503 ^ new_n27473;
  assign new_n27548 = new_n27547 ^ new_n27546;
  assign new_n27549 = ~new_n27548 & new_n27420;
  assign new_n27550 = new_n27549 ^ new_n27545;
  assign new_n27551 = ~new_n27516 & new_n27493;
  assign new_n27552 = new_n27551 ^ new_n27550;
  assign new_n27553 = new_n27552 ^ new_n27535;
  assign new_n27554 = new_n27553 ^ new_n27533;
  assign new_n27555 = new_n27554 ^ new_n27520;
  assign new_n27556 = new_n27555 ^ new_n27407;
  assign new_n27557 = new_n23507 ^ new_n23471;
  assign new_n27558 = new_n24475 ^ new_n22147;
  assign new_n27559 = new_n27558 ^ new_n14268;
  assign new_n27560 = new_n27559 ^ new_n23395;
  assign new_n27561 = new_n27560 ^ new_n23404;
  assign new_n27562 = new_n27561 ^ new_n27557;
  assign new_n27563 = new_n23466 ^ new_n23291;
  assign new_n27564 = new_n24436 ^ new_n22056;
  assign new_n27565 = new_n27564 ^ new_n14256;
  assign new_n27566 = new_n27565 ^ new_n23331;
  assign new_n27567 = new_n27566 ^ new_n23369;
  assign new_n27568 = new_n27567 ^ new_n27563;
  assign new_n27569 = new_n23552 ^ new_n23490;
  assign new_n27570 = new_n27569 ^ new_n23542;
  assign new_n27571 = new_n24616 ^ new_n22016;
  assign new_n27572 = new_n27571 ^ new_n14238;
  assign new_n27573 = new_n27572 ^ new_n23517;
  assign new_n27574 = new_n27573 ^ new_n27570;
  assign new_n27575 = new_n23547 ^ new_n23471;
  assign new_n27576 = new_n27575 ^ new_n23411;
  assign new_n27577 = new_n24596 ^ new_n21955;
  assign new_n27578 = new_n27577 ^ new_n14249;
  assign new_n27579 = new_n27578 ^ new_n23528;
  assign new_n27580 = new_n27579 ^ new_n23516;
  assign new_n27581 = new_n27580 ^ new_n27576;
  assign new_n27582 = new_n23499 ^ new_n23427;
  assign new_n27583 = new_n27582 ^ new_n23484;
  assign new_n27584 = new_n24561 ^ new_n22123;
  assign new_n27585 = new_n27584 ^ new_n14243;
  assign new_n27586 = new_n27585 ^ new_n23471;
  assign new_n27587 = new_n27586 ^ new_n23553;
  assign new_n27588 = new_n27587 ^ new_n27583;
  assign new_n27589 = new_n27588 ^ new_n27581;
  assign new_n27590 = new_n27589 ^ new_n27574;
  assign new_n27591 = new_n27590 ^ new_n27568;
  assign new_n27592 = new_n27591 ^ new_n27562;
  assign new_n27593 = new_n24541 ^ new_n21303;
  assign new_n27594 = new_n27593 ^ new_n14275;
  assign new_n27595 = new_n27594 ^ new_n23374;
  assign new_n27596 = new_n26616 ^ new_n23418;
  assign new_n27597 = new_n27596 ^ new_n27595;
  assign new_n27598 = new_n27597 ^ new_n27574;
  assign new_n27599 = new_n23437 ^ new_n23350;
  assign new_n27600 = new_n24230 ^ new_n22079;
  assign new_n27601 = new_n27600 ^ new_n14262;
  assign new_n27602 = new_n27601 ^ new_n22835;
  assign new_n27603 = new_n27602 ^ new_n23272;
  assign new_n27604 = new_n27603 ^ new_n27599;
  assign new_n27605 = new_n27604 ^ new_n27568;
  assign new_n27606 = new_n24517 ^ new_n22090;
  assign new_n27607 = new_n27606 ^ new_n14285;
  assign new_n27608 = new_n27607 ^ new_n23471;
  assign new_n27609 = new_n27608 ^ new_n23500;
  assign new_n27610 = new_n23448 ^ new_n22980;
  assign new_n27611 = new_n27610 ^ new_n23436;
  assign new_n27612 = new_n27611 ^ new_n27609;
  assign new_n27613 = new_n27612 ^ new_n27597;
  assign new_n27614 = new_n27613 ^ new_n27589;
  assign new_n27615 = new_n27614 ^ new_n27605;
  assign new_n27616 = ~new_n27615 & new_n27598;
  assign new_n27617 = new_n27591 & new_n27613;
  assign new_n27618 = new_n27617 ^ new_n27616;
  assign new_n27619 = new_n27604 ^ new_n27590;
  assign new_n27620 = new_n27619 ^ new_n27618;
  assign new_n27621 = new_n27605 ^ new_n27562;
  assign new_n27622 = new_n27621 ^ new_n27597;
  assign new_n27623 = ~new_n27592 & ~new_n27622;
  assign new_n27624 = new_n27597 ^ new_n27581;
  assign new_n27625 = ~new_n27624 & new_n27619;
  assign new_n27626 = new_n27625 ^ new_n27623;
  assign new_n27627 = new_n27626 ^ new_n27597;
  assign new_n27628 = new_n27627 ^ new_n27620;
  assign new_n27629 = new_n27581 & new_n27621;
  assign new_n27630 = new_n27629 ^ new_n27581;
  assign new_n27631 = new_n27630 ^ new_n27625;
  assign new_n27632 = new_n27631 ^ new_n27598;
  assign new_n27633 = new_n27612 ^ new_n27574;
  assign new_n27634 = new_n27612 ^ new_n27604;
  assign new_n27635 = new_n27634 ^ new_n27598;
  assign new_n27636 = ~new_n27635 & new_n27633;
  assign new_n27637 = new_n27636 ^ new_n27617;
  assign new_n27638 = new_n27604 ^ new_n27588;
  assign new_n27639 = new_n27638 ^ new_n27637;
  assign new_n27640 = new_n27639 ^ new_n27632;
  assign new_n27641 = new_n27633 ^ new_n27624;
  assign new_n27642 = ~new_n27614 & ~new_n27641;
  assign new_n27643 = new_n27642 ^ new_n27568;
  assign new_n27644 = new_n27643 ^ new_n27614;
  assign new_n27645 = new_n27614 ^ new_n27562;
  assign new_n27646 = new_n27621 ^ new_n27581;
  assign new_n27647 = new_n27646 ^ new_n27598;
  assign new_n27648 = new_n27645 & new_n27647;
  assign new_n27649 = new_n27648 ^ new_n27637;
  assign new_n27650 = new_n27649 ^ new_n27574;
  assign new_n27651 = new_n27650 ^ new_n27644;
  assign new_n27652 = ~new_n27640 & new_n27651;
  assign new_n27653 = new_n27652 ^ new_n27628;
  assign new_n27654 = new_n27604 ^ new_n27597;
  assign new_n27655 = new_n27621 ^ new_n27612;
  assign new_n27656 = ~new_n27562 & ~new_n27655;
  assign new_n27657 = new_n27656 ^ new_n27648;
  assign new_n27658 = new_n27636 ^ new_n27616;
  assign new_n27659 = new_n27658 ^ new_n27657;
  assign new_n27660 = new_n27659 ^ new_n27654;
  assign new_n27661 = ~new_n27660 & new_n27653;
  assign new_n27662 = new_n27656 ^ new_n27612;
  assign new_n27663 = new_n27662 ^ new_n27643;
  assign new_n27664 = new_n27663 ^ new_n27661;
  assign new_n27665 = new_n27664 ^ new_n27620;
  assign new_n27666 = ~new_n27592 & ~new_n27665;
  assign new_n27667 = new_n27663 ^ new_n27652;
  assign new_n27668 = new_n27667 ^ new_n27620;
  assign new_n27669 = new_n27629 ^ new_n27623;
  assign new_n27670 = new_n27669 ^ new_n27658;
  assign new_n27671 = ~new_n27668 & ~new_n27670;
  assign new_n27672 = new_n27671 ^ new_n27652;
  assign new_n27673 = ~new_n27628 & ~new_n27672;
  assign new_n27674 = new_n27673 ^ new_n27671;
  assign new_n27675 = new_n27674 ^ new_n27653;
  assign new_n27676 = new_n27675 ^ new_n27640;
  assign new_n27677 = ~new_n27641 & new_n27676;
  assign new_n27678 = new_n27677 ^ new_n27666;
  assign new_n27679 = new_n27671 ^ new_n27628;
  assign new_n27680 = ~new_n27562 & new_n27679;
  assign new_n27681 = new_n27675 ^ new_n27671;
  assign new_n27682 = new_n27681 ^ new_n27670;
  assign new_n27683 = new_n27645 & new_n27682;
  assign new_n27684 = new_n27683 ^ new_n27680;
  assign new_n27685 = ~new_n27665 & ~new_n27674;
  assign new_n27686 = new_n27685 ^ new_n27660;
  assign new_n27687 = ~new_n27621 & ~new_n27686;
  assign new_n27688 = new_n27671 ^ new_n27661;
  assign new_n27689 = new_n27663 ^ new_n27627;
  assign new_n27690 = new_n27689 ^ new_n27688;
  assign new_n27691 = ~new_n27690 & new_n27613;
  assign new_n27692 = new_n27604 ^ new_n27581;
  assign new_n27693 = new_n27648 ^ new_n27630;
  assign new_n27694 = new_n27685 ^ new_n27675;
  assign new_n27695 = new_n27694 ^ new_n27693;
  assign new_n27696 = new_n27695 ^ new_n27692;
  assign new_n27697 = new_n27696 ^ new_n27612;
  assign new_n27698 = new_n27661 ^ new_n27625;
  assign new_n27699 = new_n27698 ^ new_n27643;
  assign new_n27700 = new_n27699 ^ new_n27697;
  assign new_n27701 = new_n27633 & new_n27700;
  assign new_n27702 = new_n27701 ^ new_n27691;
  assign new_n27703 = new_n27647 & new_n27682;
  assign new_n27704 = new_n27703 ^ new_n27702;
  assign new_n27705 = new_n27704 ^ new_n27687;
  assign new_n27706 = new_n27705 ^ new_n27684;
  assign new_n27707 = new_n27706 ^ new_n27678;
  assign new_n27708 = ~new_n27470 & ~new_n27528;
  assign new_n27709 = new_n27708 ^ new_n27519;
  assign new_n27710 = new_n27509 ^ new_n27474;
  assign new_n27711 = ~new_n27467 & new_n27710;
  assign new_n27712 = new_n27711 ^ new_n27517;
  assign new_n27713 = new_n27712 ^ new_n27553;
  assign new_n27714 = new_n27713 ^ new_n27709;
  assign new_n27715 = new_n27714 ^ new_n27707;
  assign new_n27716 = new_n27715 ^ new_n27556;
  assign new_n27717 = new_n23457 ^ new_n18405;
  assign new_n27718 = new_n27717 ^ new_n25692;
  assign new_n27719 = new_n25436 ^ new_n25155;
  assign new_n27720 = new_n27719 ^ new_n25672;
  assign new_n27721 = new_n27720 ^ new_n27718;
  assign new_n27722 = new_n25759 ^ new_n25699;
  assign new_n27723 = new_n27722 ^ new_n25688;
  assign new_n27724 = new_n23442 ^ new_n18446;
  assign new_n27725 = new_n27724 ^ new_n25645;
  assign new_n27726 = new_n25681 ^ new_n25663;
  assign new_n27727 = new_n27726 ^ new_n27725;
  assign new_n27728 = new_n27727 ^ new_n27723;
  assign new_n27729 = new_n27728 ^ new_n27721;
  assign new_n27730 = new_n23478 ^ new_n18341;
  assign new_n27731 = new_n27730 ^ new_n25705;
  assign new_n27732 = new_n27731 ^ new_n27726;
  assign new_n27733 = new_n25786 ^ new_n25748;
  assign new_n27734 = new_n27733 ^ new_n25764;
  assign new_n27735 = new_n27734 ^ new_n27732;
  assign new_n27736 = new_n25776 ^ new_n25743;
  assign new_n27737 = new_n27736 ^ new_n25725;
  assign new_n27738 = new_n23522 ^ new_n18313;
  assign new_n27739 = new_n27738 ^ new_n25794;
  assign new_n27740 = new_n27739 ^ new_n27726;
  assign new_n27741 = new_n27740 ^ new_n27737;
  assign new_n27742 = new_n27741 ^ new_n27735;
  assign new_n27743 = new_n27742 ^ new_n27729;
  assign new_n27744 = new_n23385 ^ new_n18453;
  assign new_n27745 = new_n27744 ^ new_n25730;
  assign new_n27746 = new_n27726 ^ new_n25777;
  assign new_n27747 = new_n27746 ^ new_n27745;
  assign new_n27748 = new_n27747 ^ new_n27743;
  assign new_n27749 = new_n23537 ^ new_n17680;
  assign new_n27750 = new_n27749 ^ new_n25753;
  assign new_n27751 = new_n25739 ^ new_n25724;
  assign new_n27752 = new_n27751 ^ new_n25790;
  assign new_n27753 = new_n27752 ^ new_n27750;
  assign new_n27754 = new_n27753 ^ new_n27742;
  assign new_n27755 = new_n23311 ^ new_n18373;
  assign new_n27756 = new_n27755 ^ new_n25676;
  assign new_n27757 = new_n25603 ^ new_n25175;
  assign new_n27758 = new_n27757 ^ new_n25437;
  assign new_n27759 = new_n27758 ^ new_n27756;
  assign new_n27760 = new_n27759 ^ new_n27754;
  assign new_n27761 = new_n27729 & new_n27760;
  assign new_n27762 = new_n27753 ^ new_n27721;
  assign new_n27763 = new_n22682 ^ new_n18421;
  assign new_n27764 = new_n27763 ^ new_n25582;
  assign new_n27765 = new_n25686 ^ new_n25651;
  assign new_n27766 = new_n27765 ^ new_n25623;
  assign new_n27767 = new_n27766 ^ new_n27764;
  assign new_n27768 = new_n27767 ^ new_n27759;
  assign new_n27769 = new_n27768 ^ new_n27743;
  assign new_n27770 = ~new_n27769 & new_n27762;
  assign new_n27771 = new_n27770 ^ new_n27761;
  assign new_n27772 = new_n27767 ^ new_n27754;
  assign new_n27773 = new_n27772 ^ new_n27771;
  assign new_n27774 = new_n27741 ^ new_n27721;
  assign new_n27775 = ~new_n27774 & new_n27772;
  assign new_n27776 = new_n27768 ^ new_n27747;
  assign new_n27777 = new_n27776 ^ new_n27721;
  assign new_n27778 = new_n27760 ^ new_n27747;
  assign new_n27779 = ~new_n27777 & ~new_n27778;
  assign new_n27780 = new_n27779 ^ new_n27775;
  assign new_n27781 = new_n27780 ^ new_n27721;
  assign new_n27782 = new_n27781 ^ new_n27773;
  assign new_n27783 = new_n27741 & new_n27776;
  assign new_n27784 = new_n27783 ^ new_n27741;
  assign new_n27785 = new_n27784 ^ new_n27775;
  assign new_n27786 = new_n27785 ^ new_n27762;
  assign new_n27787 = new_n27767 ^ new_n27728;
  assign new_n27788 = new_n27787 ^ new_n27762;
  assign new_n27789 = new_n27753 ^ new_n27728;
  assign new_n27790 = ~new_n27788 & new_n27789;
  assign new_n27791 = new_n27790 ^ new_n27761;
  assign new_n27792 = new_n27767 ^ new_n27735;
  assign new_n27793 = new_n27792 ^ new_n27791;
  assign new_n27794 = new_n27793 ^ new_n27786;
  assign new_n27795 = new_n27741 ^ new_n27728;
  assign new_n27796 = new_n27795 ^ new_n27762;
  assign new_n27797 = ~new_n27743 & ~new_n27796;
  assign new_n27798 = new_n27797 ^ new_n27759;
  assign new_n27799 = new_n27798 ^ new_n27743;
  assign new_n27800 = new_n27776 ^ new_n27741;
  assign new_n27801 = new_n27800 ^ new_n27762;
  assign new_n27802 = new_n27748 & new_n27801;
  assign new_n27803 = new_n27802 ^ new_n27761;
  assign new_n27804 = new_n27790 ^ new_n27753;
  assign new_n27805 = new_n27804 ^ new_n27803;
  assign new_n27806 = new_n27805 ^ new_n27799;
  assign new_n27807 = ~new_n27794 & new_n27806;
  assign new_n27808 = new_n27776 ^ new_n27728;
  assign new_n27809 = ~new_n27747 & ~new_n27808;
  assign new_n27810 = new_n27809 ^ new_n27728;
  assign new_n27811 = new_n27810 ^ new_n27798;
  assign new_n27812 = new_n27811 ^ new_n27807;
  assign new_n27813 = new_n27812 ^ new_n27773;
  assign new_n27814 = new_n27783 ^ new_n27779;
  assign new_n27815 = new_n27790 ^ new_n27770;
  assign new_n27816 = new_n27815 ^ new_n27814;
  assign new_n27817 = ~new_n27813 & ~new_n27816;
  assign new_n27818 = new_n27817 ^ new_n27807;
  assign new_n27819 = ~new_n27818 & new_n27782;
  assign new_n27820 = new_n27819 ^ new_n27782;
  assign new_n27821 = new_n27820 ^ new_n27817;
  assign new_n27822 = new_n27821 ^ new_n27816;
  assign new_n27823 = ~new_n27822 & new_n27748;
  assign new_n27824 = new_n27820 ^ new_n27794;
  assign new_n27825 = ~new_n27743 & ~new_n27824;
  assign new_n27826 = new_n27825 ^ new_n27823;
  assign new_n27827 = ~new_n27796 & ~new_n27824;
  assign new_n27828 = new_n27827 ^ new_n27826;
  assign new_n27829 = new_n27767 ^ new_n27721;
  assign new_n27830 = new_n27809 ^ new_n27802;
  assign new_n27831 = new_n27830 ^ new_n27815;
  assign new_n27832 = new_n27831 ^ new_n27829;
  assign new_n27833 = new_n27807 ^ new_n27782;
  assign new_n27834 = ~new_n27832 & new_n27833;
  assign new_n27835 = new_n27834 ^ new_n27811;
  assign new_n27836 = new_n27835 ^ new_n27773;
  assign new_n27837 = new_n27819 ^ new_n27807;
  assign new_n27838 = ~new_n27836 & new_n27837;
  assign new_n27839 = new_n27838 ^ new_n27832;
  assign new_n27840 = ~new_n27776 & ~new_n27839;
  assign new_n27841 = new_n27834 ^ new_n27817;
  assign new_n27842 = new_n27811 ^ new_n27781;
  assign new_n27843 = new_n27842 ^ new_n27841;
  assign new_n27844 = ~new_n27843 & new_n27729;
  assign new_n27845 = new_n27767 ^ new_n27741;
  assign new_n27846 = new_n27802 ^ new_n27784;
  assign new_n27847 = new_n27838 ^ new_n27820;
  assign new_n27848 = new_n27847 ^ new_n27846;
  assign new_n27849 = new_n27848 ^ new_n27845;
  assign new_n27850 = new_n27849 ^ new_n27728;
  assign new_n27851 = new_n27834 ^ new_n27775;
  assign new_n27852 = new_n27851 ^ new_n27798;
  assign new_n27853 = new_n27852 ^ new_n27850;
  assign new_n27854 = ~new_n27853 & new_n27789;
  assign new_n27855 = new_n27854 ^ new_n27844;
  assign new_n27856 = ~new_n27822 & new_n27801;
  assign new_n27857 = new_n27856 ^ new_n27855;
  assign new_n27858 = new_n27857 ^ new_n27840;
  assign new_n27859 = new_n27838 ^ new_n27834;
  assign new_n27860 = new_n27859 ^ new_n27806;
  assign new_n27861 = new_n27772 & new_n27860;
  assign new_n27862 = new_n27861 ^ new_n27858;
  assign new_n27863 = new_n27862 ^ new_n27828;
  assign new_n27864 = new_n27416 ^ new_n27410;
  assign new_n27865 = new_n27427 ^ new_n27423;
  assign new_n27866 = new_n27865 ^ new_n27864;
  assign new_n27867 = new_n27866 ^ new_n27464;
  assign new_n27868 = new_n27865 ^ new_n27441;
  assign new_n27869 = new_n27868 ^ new_n27437;
  assign new_n27870 = new_n27864 & new_n27869;
  assign new_n27871 = new_n27441 ^ new_n27410;
  assign new_n27872 = new_n27452 ^ new_n27437;
  assign new_n27873 = new_n27872 ^ new_n27866;
  assign new_n27874 = new_n27871 & new_n27873;
  assign new_n27875 = new_n27874 ^ new_n27870;
  assign new_n27876 = new_n27868 ^ new_n27452;
  assign new_n27877 = new_n27876 ^ new_n27875;
  assign new_n27878 = new_n27423 ^ new_n27410;
  assign new_n27879 = new_n27876 & new_n27878;
  assign new_n27880 = new_n27872 ^ new_n27464;
  assign new_n27881 = new_n27880 ^ new_n27410;
  assign new_n27882 = new_n27869 ^ new_n27464;
  assign new_n27883 = new_n27881 & new_n27882;
  assign new_n27884 = new_n27883 ^ new_n27879;
  assign new_n27885 = new_n27884 ^ new_n27410;
  assign new_n27886 = new_n27885 ^ new_n27877;
  assign new_n27887 = ~new_n27423 & ~new_n27880;
  assign new_n27888 = new_n27887 ^ new_n27423;
  assign new_n27889 = new_n27888 ^ new_n27879;
  assign new_n27890 = new_n27889 ^ new_n27871;
  assign new_n27891 = new_n27452 ^ new_n27416;
  assign new_n27892 = new_n27891 ^ new_n27871;
  assign new_n27893 = new_n27441 ^ new_n27416;
  assign new_n27894 = new_n27892 & new_n27893;
  assign new_n27895 = new_n27894 ^ new_n27870;
  assign new_n27896 = new_n27452 ^ new_n27427;
  assign new_n27897 = new_n27896 ^ new_n27895;
  assign new_n27898 = new_n27897 ^ new_n27890;
  assign new_n27899 = new_n27423 ^ new_n27416;
  assign new_n27900 = new_n27899 ^ new_n27871;
  assign new_n27901 = new_n27866 & new_n27900;
  assign new_n27902 = new_n27901 ^ new_n27437;
  assign new_n27903 = new_n27902 ^ new_n27866;
  assign new_n27904 = new_n27880 ^ new_n27423;
  assign new_n27905 = new_n27904 ^ new_n27871;
  assign new_n27906 = new_n27867 & new_n27905;
  assign new_n27907 = new_n27906 ^ new_n27441;
  assign new_n27908 = new_n27907 ^ new_n27895;
  assign new_n27909 = new_n27908 ^ new_n27903;
  assign new_n27910 = ~new_n27898 & new_n27909;
  assign new_n27911 = new_n27880 ^ new_n27416;
  assign new_n27912 = new_n27464 & new_n27911;
  assign new_n27913 = new_n27912 ^ new_n27416;
  assign new_n27914 = new_n27913 ^ new_n27902;
  assign new_n27915 = new_n27914 ^ new_n27910;
  assign new_n27916 = new_n27915 ^ new_n27877;
  assign new_n27917 = new_n27887 ^ new_n27883;
  assign new_n27918 = new_n27894 ^ new_n27874;
  assign new_n27919 = new_n27918 ^ new_n27917;
  assign new_n27920 = ~new_n27919 & new_n27916;
  assign new_n27921 = new_n27920 ^ new_n27910;
  assign new_n27922 = ~new_n27921 & new_n27886;
  assign new_n27923 = new_n27922 ^ new_n27886;
  assign new_n27924 = new_n27923 ^ new_n27920;
  assign new_n27925 = new_n27924 ^ new_n27919;
  assign new_n27926 = ~new_n27925 & new_n27867;
  assign new_n27927 = new_n27923 ^ new_n27898;
  assign new_n27928 = ~new_n27927 & new_n27866;
  assign new_n27929 = new_n27928 ^ new_n27926;
  assign new_n27930 = ~new_n27927 & new_n27900;
  assign new_n27931 = new_n27930 ^ new_n27929;
  assign new_n27932 = new_n27452 ^ new_n27410;
  assign new_n27933 = new_n27912 ^ new_n27906;
  assign new_n27934 = new_n27933 ^ new_n27918;
  assign new_n27935 = new_n27934 ^ new_n27932;
  assign new_n27936 = new_n27910 ^ new_n27886;
  assign new_n27937 = new_n27935 & new_n27936;
  assign new_n27938 = new_n27937 ^ new_n27914;
  assign new_n27939 = new_n27938 ^ new_n27877;
  assign new_n27940 = new_n27922 ^ new_n27910;
  assign new_n27941 = new_n27939 & new_n27940;
  assign new_n27942 = new_n27941 ^ new_n27935;
  assign new_n27943 = new_n27880 & new_n27942;
  assign new_n27944 = new_n27937 ^ new_n27920;
  assign new_n27945 = new_n27914 ^ new_n27885;
  assign new_n27946 = new_n27945 ^ new_n27944;
  assign new_n27947 = new_n27864 & new_n27946;
  assign new_n27948 = new_n27452 ^ new_n27423;
  assign new_n27949 = new_n27906 ^ new_n27888;
  assign new_n27950 = new_n27941 ^ new_n27923;
  assign new_n27951 = new_n27950 ^ new_n27949;
  assign new_n27952 = new_n27951 ^ new_n27948;
  assign new_n27953 = new_n27952 ^ new_n27416;
  assign new_n27954 = new_n27937 ^ new_n27879;
  assign new_n27955 = new_n27954 ^ new_n27902;
  assign new_n27956 = new_n27955 ^ new_n27953;
  assign new_n27957 = ~new_n27956 & new_n27893;
  assign new_n27958 = new_n27957 ^ new_n27947;
  assign new_n27959 = ~new_n27925 & new_n27905;
  assign new_n27960 = new_n27959 ^ new_n27958;
  assign new_n27961 = new_n27960 ^ new_n27943;
  assign new_n27962 = new_n27941 ^ new_n27937;
  assign new_n27963 = new_n27962 ^ new_n27909;
  assign new_n27964 = new_n27876 & new_n27963;
  assign new_n27965 = new_n27964 ^ new_n27961;
  assign new_n27966 = new_n27965 ^ new_n27931;
  assign new_n27967 = new_n24517 ^ new_n22988;
  assign new_n27968 = new_n27967 ^ new_n27966;
  assign new_n27969 = new_n27968 ^ new_n27863;
  assign new_n27970 = ~new_n27690 & new_n27591;
  assign new_n27971 = new_n27970 ^ new_n27677;
  assign new_n27972 = new_n27685 ^ new_n27661;
  assign new_n27973 = new_n27972 ^ new_n27651;
  assign new_n27974 = new_n27619 & new_n27973;
  assign new_n27975 = new_n27974 ^ new_n27705;
  assign new_n27976 = ~new_n27635 & new_n27700;
  assign new_n27977 = new_n27976 ^ new_n27975;
  assign new_n27978 = new_n27977 ^ new_n27971;
  assign new_n27979 = ~new_n27480 & ~new_n27544;
  assign new_n27980 = new_n27979 ^ new_n27554;
  assign new_n27981 = ~new_n27548 & new_n27447;
  assign new_n27982 = new_n27981 ^ new_n27519;
  assign new_n27983 = new_n27982 ^ new_n27980;
  assign new_n27984 = new_n27983 ^ new_n27978;
  assign new_n27985 = new_n27984 ^ new_n27969;
  assign new_n27986 = new_n27985 ^ new_n27716;
  assign new_n27987 = ~new_n27843 & new_n27760;
  assign new_n27988 = new_n27987 ^ new_n27844;
  assign new_n27989 = new_n27817 ^ new_n27721;
  assign new_n27990 = new_n27809 ^ new_n27779;
  assign new_n27991 = new_n27990 ^ new_n27849;
  assign new_n27992 = new_n27991 ^ new_n27989;
  assign new_n27993 = new_n27762 & new_n27992;
  assign new_n27994 = ~new_n27774 & new_n27860;
  assign new_n27995 = new_n27817 ^ new_n27782;
  assign new_n27996 = ~new_n27747 & new_n27995;
  assign new_n27997 = new_n27996 ^ new_n27825;
  assign new_n27998 = new_n27997 ^ new_n27994;
  assign new_n27999 = ~new_n27769 & new_n27992;
  assign new_n28000 = ~new_n27777 & ~new_n27836;
  assign new_n28001 = new_n28000 ^ new_n27999;
  assign new_n28002 = new_n28001 ^ new_n27998;
  assign new_n28003 = new_n28002 ^ new_n27993;
  assign new_n28004 = new_n28003 ^ new_n27988;
  assign new_n28005 = new_n27869 & new_n27946;
  assign new_n28006 = new_n28005 ^ new_n27947;
  assign new_n28007 = new_n27920 ^ new_n27410;
  assign new_n28008 = new_n27912 ^ new_n27883;
  assign new_n28009 = new_n28008 ^ new_n27952;
  assign new_n28010 = new_n28009 ^ new_n28007;
  assign new_n28011 = ~new_n28010 & new_n27871;
  assign new_n28012 = new_n27878 & new_n27963;
  assign new_n28013 = new_n27920 ^ new_n27886;
  assign new_n28014 = new_n27464 & new_n28013;
  assign new_n28015 = new_n28014 ^ new_n27928;
  assign new_n28016 = new_n28015 ^ new_n28012;
  assign new_n28017 = ~new_n28010 & new_n27873;
  assign new_n28018 = new_n27881 & new_n27939;
  assign new_n28019 = new_n28018 ^ new_n28017;
  assign new_n28020 = new_n28019 ^ new_n28016;
  assign new_n28021 = new_n28020 ^ new_n28011;
  assign new_n28022 = new_n28021 ^ new_n28006;
  assign new_n28023 = new_n24230 ^ new_n23027;
  assign new_n28024 = new_n28023 ^ new_n28022;
  assign new_n28025 = new_n28024 ^ new_n28004;
  assign new_n28026 = ~new_n27614 & new_n27676;
  assign new_n28027 = new_n28026 ^ new_n27683;
  assign new_n28028 = new_n28027 ^ new_n27677;
  assign new_n28029 = new_n28028 ^ new_n27975;
  assign new_n28030 = new_n28029 ^ new_n27555;
  assign new_n28031 = new_n27305 & new_n27387;
  assign new_n28032 = new_n28031 ^ new_n27388;
  assign new_n28033 = new_n27361 ^ new_n27261;
  assign new_n28034 = new_n27353 ^ new_n27324;
  assign new_n28035 = new_n28034 ^ new_n27393;
  assign new_n28036 = new_n28035 ^ new_n28033;
  assign new_n28037 = ~new_n27307 & new_n28036;
  assign new_n28038 = ~new_n27319 & ~new_n27404;
  assign new_n28039 = new_n27361 ^ new_n27327;
  assign new_n28040 = ~new_n27291 & new_n28039;
  assign new_n28041 = new_n28040 ^ new_n27369;
  assign new_n28042 = new_n28041 ^ new_n28038;
  assign new_n28043 = ~new_n27314 & new_n28036;
  assign new_n28044 = ~new_n27322 & new_n27380;
  assign new_n28045 = new_n28044 ^ new_n28043;
  assign new_n28046 = new_n28045 ^ new_n28042;
  assign new_n28047 = new_n28046 ^ new_n28037;
  assign new_n28048 = new_n28047 ^ new_n28032;
  assign new_n28049 = new_n27981 ^ new_n27549;
  assign new_n28050 = new_n27509 ^ new_n27413;
  assign new_n28051 = new_n27501 ^ new_n27471;
  assign new_n28052 = new_n28051 ^ new_n27540;
  assign new_n28053 = new_n28052 ^ new_n28050;
  assign new_n28054 = new_n27449 & new_n28053;
  assign new_n28055 = new_n27711 ^ new_n27514;
  assign new_n28056 = ~new_n27461 & new_n27532;
  assign new_n28057 = new_n28056 ^ new_n28055;
  assign new_n28058 = ~new_n27469 & ~new_n27528;
  assign new_n28059 = ~new_n27456 & new_n28053;
  assign new_n28060 = new_n28059 ^ new_n28058;
  assign new_n28061 = new_n28060 ^ new_n28057;
  assign new_n28062 = new_n28061 ^ new_n28054;
  assign new_n28063 = new_n28062 ^ new_n28049;
  assign new_n28064 = new_n28063 ^ new_n28048;
  assign new_n28065 = new_n28064 ^ new_n28030;
  assign new_n28066 = new_n28065 ^ new_n28025;
  assign new_n28067 = new_n28066 ^ new_n27986;
  assign new_n28068 = ~new_n27624 & new_n27973;
  assign new_n28069 = new_n27671 ^ new_n27597;
  assign new_n28070 = new_n27656 ^ new_n27623;
  assign new_n28071 = new_n28070 ^ new_n27696;
  assign new_n28072 = new_n28071 ^ new_n28069;
  assign new_n28073 = ~new_n27615 & ~new_n28072;
  assign new_n28074 = new_n28073 ^ new_n28068;
  assign new_n28075 = new_n27976 ^ new_n27687;
  assign new_n28076 = ~new_n27686 & new_n27646;
  assign new_n28077 = new_n28076 ^ new_n27666;
  assign new_n28078 = new_n28077 ^ new_n27702;
  assign new_n28079 = new_n28078 ^ new_n28075;
  assign new_n28080 = new_n28079 ^ new_n28074;
  assign new_n28081 = new_n27352 & new_n28039;
  assign new_n28082 = ~new_n27333 & new_n27397;
  assign new_n28083 = new_n28082 ^ new_n27406;
  assign new_n28084 = new_n28083 ^ new_n28081;
  assign new_n28085 = new_n28084 ^ new_n28046;
  assign new_n28086 = ~new_n27500 & new_n27710;
  assign new_n28087 = new_n28086 ^ new_n27980;
  assign new_n28088 = new_n28087 ^ new_n28061;
  assign new_n28089 = new_n28088 ^ new_n28085;
  assign new_n28090 = new_n28089 ^ new_n28080;
  assign new_n28091 = ~new_n27808 & new_n27995;
  assign new_n28092 = ~new_n27788 & ~new_n27853;
  assign new_n28093 = new_n28092 ^ new_n27862;
  assign new_n28094 = new_n28093 ^ new_n28091;
  assign new_n28095 = new_n28094 ^ new_n28002;
  assign new_n28096 = new_n27911 & new_n28013;
  assign new_n28097 = ~new_n27956 & new_n27892;
  assign new_n28098 = new_n28097 ^ new_n27965;
  assign new_n28099 = new_n28098 ^ new_n28096;
  assign new_n28100 = new_n28099 ^ new_n28020;
  assign new_n28101 = new_n24616 ^ new_n23012;
  assign new_n28102 = new_n28101 ^ new_n28100;
  assign new_n28103 = new_n28102 ^ new_n28095;
  assign new_n28104 = new_n28059 ^ new_n28056;
  assign new_n28105 = new_n27979 ^ new_n27535;
  assign new_n28106 = ~new_n27534 & new_n27492;
  assign new_n28107 = new_n28106 ^ new_n27708;
  assign new_n28108 = new_n28107 ^ new_n27550;
  assign new_n28109 = new_n28108 ^ new_n28105;
  assign new_n28110 = new_n28109 ^ new_n28104;
  assign new_n28111 = new_n28110 ^ new_n28103;
  assign new_n28112 = new_n28111 ^ new_n28090;
  assign new_n28113 = new_n27987 ^ new_n27827;
  assign new_n28114 = new_n28113 ^ new_n28093;
  assign new_n28115 = new_n28005 ^ new_n27930;
  assign new_n28116 = new_n28115 ^ new_n28098;
  assign new_n28117 = new_n24541 ^ new_n22981;
  assign new_n28118 = new_n28117 ^ new_n28116;
  assign new_n28119 = new_n28118 ^ new_n28114;
  assign new_n28120 = new_n27981 ^ new_n27979;
  assign new_n28121 = new_n27552 ^ new_n27520;
  assign new_n28122 = new_n28121 ^ new_n28120;
  assign new_n28123 = new_n27976 ^ new_n27970;
  assign new_n28124 = new_n28028 ^ new_n27704;
  assign new_n28125 = new_n28124 ^ new_n28123;
  assign new_n28126 = new_n28125 ^ new_n28122;
  assign new_n28127 = new_n28031 ^ new_n27371;
  assign new_n28128 = new_n28127 ^ new_n28083;
  assign new_n28129 = new_n28128 ^ new_n27983;
  assign new_n28130 = new_n28129 ^ new_n28126;
  assign new_n28131 = new_n28130 ^ new_n28119;
  assign new_n28132 = new_n28131 ^ new_n28112;
  assign new_n28133 = new_n28132 ^ new_n28067;
  assign new_n28134 = new_n27999 ^ new_n27994;
  assign new_n28135 = new_n28092 ^ new_n27840;
  assign new_n28136 = ~new_n27778 & ~new_n27836;
  assign new_n28137 = ~new_n27839 & new_n27800;
  assign new_n28138 = new_n28137 ^ new_n28136;
  assign new_n28139 = new_n28138 ^ new_n27855;
  assign new_n28140 = new_n28139 ^ new_n28135;
  assign new_n28141 = new_n28140 ^ new_n28134;
  assign new_n28142 = new_n28141 ^ new_n28110;
  assign new_n28143 = new_n28142 ^ new_n27984;
  assign new_n28144 = new_n28026 ^ new_n27680;
  assign new_n28145 = new_n28144 ^ new_n28068;
  assign new_n28146 = new_n28145 ^ new_n27974;
  assign new_n28147 = new_n28146 ^ new_n28078;
  assign new_n28148 = new_n28057 ^ new_n27533;
  assign new_n28149 = new_n28148 ^ new_n28108;
  assign new_n28150 = new_n28149 ^ new_n28147;
  assign new_n28151 = new_n28017 ^ new_n28012;
  assign new_n28152 = new_n28097 ^ new_n27943;
  assign new_n28153 = new_n27882 & new_n27939;
  assign new_n28154 = new_n27904 & new_n27942;
  assign new_n28155 = new_n28154 ^ new_n28153;
  assign new_n28156 = new_n28155 ^ new_n27958;
  assign new_n28157 = new_n28156 ^ new_n28152;
  assign new_n28158 = new_n28157 ^ new_n28151;
  assign new_n28159 = new_n24596 ^ new_n23000;
  assign new_n28160 = new_n28159 ^ new_n28158;
  assign new_n28161 = new_n28043 ^ new_n28038;
  assign new_n28162 = new_n28082 ^ new_n27384;
  assign new_n28163 = ~new_n27323 & new_n27380;
  assign new_n28164 = ~new_n27383 & new_n27345;
  assign new_n28165 = new_n28164 ^ new_n28163;
  assign new_n28166 = new_n28165 ^ new_n27399;
  assign new_n28167 = new_n28166 ^ new_n28162;
  assign new_n28168 = new_n28167 ^ new_n28161;
  assign new_n28169 = new_n28168 ^ new_n28160;
  assign new_n28170 = new_n28169 ^ new_n28150;
  assign new_n28171 = new_n28170 ^ new_n28143;
  assign new_n28172 = new_n28171 ^ new_n28066;
  assign new_n28173 = new_n28092 ^ new_n27987;
  assign new_n28174 = new_n27857 ^ new_n27828;
  assign new_n28175 = new_n28174 ^ new_n28173;
  assign new_n28176 = new_n28097 ^ new_n28005;
  assign new_n28177 = new_n27960 ^ new_n27931;
  assign new_n28178 = new_n28177 ^ new_n28176;
  assign new_n28179 = new_n24436 ^ new_n23019;
  assign new_n28180 = new_n28179 ^ new_n28178;
  assign new_n28181 = new_n28180 ^ new_n28175;
  assign new_n28182 = new_n27970 ^ new_n27691;
  assign new_n28183 = ~new_n27622 & ~new_n27665;
  assign new_n28184 = new_n28183 ^ new_n28073;
  assign new_n28185 = new_n28184 ^ new_n28145;
  assign new_n28186 = ~new_n28072 & new_n27598;
  assign new_n28187 = new_n28186 ^ new_n28185;
  assign new_n28188 = new_n28187 ^ new_n28182;
  assign new_n28189 = new_n28188 ^ new_n28063;
  assign new_n28190 = new_n28082 ^ new_n28031;
  assign new_n28191 = new_n27401 ^ new_n27372;
  assign new_n28192 = new_n28191 ^ new_n28190;
  assign new_n28193 = new_n28192 ^ new_n28122;
  assign new_n28194 = new_n28193 ^ new_n28189;
  assign new_n28195 = new_n28194 ^ new_n28181;
  assign new_n28196 = new_n28195 ^ new_n28066;
  assign new_n28197 = new_n28042 ^ new_n27405;
  assign new_n28198 = new_n28197 ^ new_n28166;
  assign new_n28199 = new_n28016 ^ new_n27964;
  assign new_n28200 = new_n28199 ^ new_n28156;
  assign new_n28201 = new_n24475 ^ new_n23007;
  assign new_n28202 = new_n28201 ^ new_n28200;
  assign new_n28203 = new_n28202 ^ new_n28198;
  assign new_n28204 = new_n27998 ^ new_n27861;
  assign new_n28205 = new_n28204 ^ new_n28139;
  assign new_n28206 = new_n28205 ^ new_n28149;
  assign new_n28207 = new_n28206 ^ new_n27984;
  assign new_n28208 = new_n28207 ^ new_n28203;
  assign new_n28209 = new_n28208 ^ new_n28196;
  assign new_n28210 = new_n28171 & new_n28209;
  assign new_n28211 = new_n28210 ^ new_n28171;
  assign new_n28212 = new_n28209 ^ new_n28171;
  assign new_n28213 = new_n28212 ^ new_n28132;
  assign new_n28214 = new_n28131 ^ new_n27986;
  assign new_n28215 = new_n28136 ^ new_n27827;
  assign new_n28216 = new_n27996 ^ new_n27823;
  assign new_n28217 = new_n28216 ^ new_n27858;
  assign new_n28218 = new_n28217 ^ new_n28215;
  assign new_n28219 = new_n28153 ^ new_n27930;
  assign new_n28220 = new_n28014 ^ new_n27926;
  assign new_n28221 = new_n28220 ^ new_n27961;
  assign new_n28222 = new_n28221 ^ new_n28219;
  assign new_n28223 = new_n24561 ^ new_n22993;
  assign new_n28224 = new_n28223 ^ new_n28222;
  assign new_n28225 = new_n28224 ^ new_n28218;
  assign new_n28226 = new_n28225 ^ new_n27984;
  assign new_n28227 = ~new_n27655 & new_n27679;
  assign new_n28228 = new_n28227 ^ new_n27977;
  assign new_n28229 = new_n28228 ^ new_n28185;
  assign new_n28230 = new_n28229 ^ new_n28088;
  assign new_n28231 = new_n28163 ^ new_n27371;
  assign new_n28232 = new_n28040 ^ new_n27367;
  assign new_n28233 = new_n28232 ^ new_n27402;
  assign new_n28234 = new_n28233 ^ new_n28231;
  assign new_n28235 = new_n28234 ^ new_n27714;
  assign new_n28236 = new_n28235 ^ new_n28230;
  assign new_n28237 = new_n28236 ^ new_n28226;
  assign new_n28238 = new_n28237 ^ new_n28171;
  assign new_n28239 = new_n28238 ^ new_n28214;
  assign new_n28240 = new_n28239 ^ new_n28208;
  assign new_n28241 = new_n28213 & new_n28240;
  assign new_n28242 = new_n28241 ^ new_n28211;
  assign new_n28243 = new_n28171 ^ new_n27986;
  assign new_n28244 = new_n28243 ^ new_n28132;
  assign new_n28245 = ~new_n28239 & ~new_n28244;
  assign new_n28246 = new_n28245 ^ new_n28195;
  assign new_n28247 = ~new_n28196 & ~new_n28208;
  assign new_n28248 = new_n27986 & new_n28208;
  assign new_n28249 = new_n28248 ^ new_n28247;
  assign new_n28250 = new_n28249 ^ new_n28246;
  assign new_n28251 = new_n28131 ^ new_n28066;
  assign new_n28252 = new_n28239 ^ new_n28196;
  assign new_n28253 = ~new_n28252 & new_n28132;
  assign new_n28254 = new_n28112 ^ new_n27986;
  assign new_n28255 = ~new_n28133 & new_n28254;
  assign new_n28256 = new_n28255 ^ new_n28253;
  assign new_n28257 = new_n28249 ^ new_n27986;
  assign new_n28258 = new_n28257 ^ new_n28241;
  assign new_n28259 = new_n28258 ^ new_n28256;
  assign new_n28260 = new_n28259 ^ new_n28251;
  assign new_n28261 = new_n28238 ^ new_n28112;
  assign new_n28262 = new_n28261 ^ new_n28195;
  assign new_n28263 = new_n28214 & new_n28262;
  assign new_n28264 = new_n28263 ^ new_n28253;
  assign new_n28265 = new_n28261 ^ new_n28066;
  assign new_n28266 = new_n28265 ^ new_n28264;
  assign new_n28267 = new_n28171 ^ new_n28131;
  assign new_n28268 = ~new_n28267 & new_n28265;
  assign new_n28269 = new_n28209 ^ new_n28131;
  assign new_n28270 = new_n28262 ^ new_n28208;
  assign new_n28271 = ~new_n28269 & ~new_n28270;
  assign new_n28272 = new_n28271 ^ new_n28268;
  assign new_n28273 = new_n28272 ^ new_n28131;
  assign new_n28274 = new_n28273 ^ new_n28266;
  assign new_n28275 = new_n28268 ^ new_n28211;
  assign new_n28276 = new_n28275 ^ new_n28132;
  assign new_n28277 = new_n28263 ^ new_n28255;
  assign new_n28278 = new_n28237 ^ new_n28066;
  assign new_n28279 = new_n28278 ^ new_n28277;
  assign new_n28280 = new_n28279 ^ new_n28276;
  assign new_n28281 = new_n28246 ^ new_n28239;
  assign new_n28282 = new_n28277 ^ new_n28241;
  assign new_n28283 = new_n28282 ^ new_n28112;
  assign new_n28284 = new_n28283 ^ new_n28281;
  assign new_n28285 = ~new_n28280 & new_n28284;
  assign new_n28286 = new_n28285 ^ new_n28274;
  assign new_n28287 = ~new_n28260 & new_n28286;
  assign new_n28288 = new_n28287 ^ new_n28250;
  assign new_n28289 = new_n28288 ^ new_n28266;
  assign new_n28290 = new_n28285 ^ new_n28250;
  assign new_n28291 = new_n28290 ^ new_n28266;
  assign new_n28292 = new_n28271 ^ new_n28210;
  assign new_n28293 = new_n28292 ^ new_n28256;
  assign new_n28294 = ~new_n28291 & ~new_n28293;
  assign new_n28295 = new_n28294 ^ new_n28285;
  assign new_n28296 = new_n28274 & new_n28295;
  assign new_n28297 = new_n28296 ^ new_n28286;
  assign new_n28298 = ~new_n28289 & new_n28297;
  assign new_n28299 = new_n28298 ^ new_n28296;
  assign new_n28300 = new_n28299 ^ new_n28242;
  assign new_n28301 = new_n28300 ^ new_n28172;
  assign new_n28302 = new_n28301 ^ new_n27986;
  assign new_n28303 = new_n28287 ^ new_n28268;
  assign new_n28304 = new_n28303 ^ new_n28246;
  assign new_n28305 = new_n28304 ^ new_n28302;
  assign new_n28306 = ~new_n28133 & ~new_n28305;
  assign new_n28307 = new_n28294 ^ new_n28287;
  assign new_n28308 = new_n28273 ^ new_n28250;
  assign new_n28309 = new_n28308 ^ new_n28307;
  assign new_n28310 = ~new_n28309 & new_n28262;
  assign new_n28311 = new_n28310 ^ new_n28306;
  assign new_n28312 = new_n28296 ^ new_n28294;
  assign new_n28313 = new_n28312 ^ new_n28293;
  assign new_n28314 = ~new_n28313 & new_n28240;
  assign new_n28315 = new_n28296 ^ new_n28280;
  assign new_n28316 = ~new_n28239 & ~new_n28315;
  assign new_n28317 = new_n28316 ^ new_n28314;
  assign new_n28318 = ~new_n28244 & ~new_n28315;
  assign new_n28319 = new_n28318 ^ new_n28317;
  assign new_n28320 = ~new_n28313 & new_n28213;
  assign new_n28321 = ~new_n28305 & new_n28254;
  assign new_n28322 = ~new_n28309 & new_n28214;
  assign new_n28323 = new_n28322 ^ new_n28321;
  assign new_n28324 = new_n28323 ^ new_n28320;
  assign new_n28325 = new_n28324 ^ new_n28319;
  assign new_n28326 = new_n28325 ^ new_n28311;
  assign new_n28327 = new_n28326 ^ new_n27255;
  assign new_n28328 = new_n28327 ^ new_n26210;
  assign new_n28329 = new_n23522 ^ new_n12759;
  assign new_n28330 = new_n23478 ^ new_n12758;
  assign new_n28331 = new_n28330 ^ new_n28329;
  assign new_n28332 = new_n23457 ^ new_n12761;
  assign new_n28333 = new_n23442 ^ new_n12762;
  assign new_n28334 = new_n28333 ^ new_n28332;
  assign new_n28335 = new_n28334 ^ new_n28331;
  assign new_n28336 = new_n23311 ^ new_n12768;
  assign new_n28337 = new_n22682 ^ new_n12767;
  assign new_n28338 = new_n28337 ^ new_n28336;
  assign new_n28339 = new_n23385 ^ new_n12780;
  assign new_n28340 = new_n28339 ^ new_n28338;
  assign new_n28341 = new_n28340 ^ new_n28332;
  assign new_n28342 = new_n23537 ^ new_n12765;
  assign new_n28343 = new_n28342 ^ new_n28331;
  assign new_n28344 = new_n28343 ^ new_n28336;
  assign new_n28345 = new_n28344 ^ new_n28339;
  assign new_n28346 = new_n28341 & new_n28345;
  assign new_n28347 = new_n28343 ^ new_n28337;
  assign new_n28348 = new_n28332 ^ new_n28329;
  assign new_n28349 = new_n28347 & new_n28348;
  assign new_n28350 = new_n28349 ^ new_n28346;
  assign new_n28351 = new_n28350 ^ new_n28332;
  assign new_n28352 = new_n28342 ^ new_n28332;
  assign new_n28353 = new_n28338 ^ new_n28335;
  assign new_n28354 = new_n28352 & new_n28353;
  assign new_n28355 = new_n28334 & new_n28344;
  assign new_n28356 = new_n28355 ^ new_n28354;
  assign new_n28357 = new_n28356 ^ new_n28347;
  assign new_n28358 = new_n28357 ^ new_n28351;
  assign new_n28359 = ~new_n28329 & ~new_n28340;
  assign new_n28360 = new_n28359 ^ new_n28329;
  assign new_n28361 = new_n28360 ^ new_n28349;
  assign new_n28362 = new_n28361 ^ new_n28352;
  assign new_n28363 = new_n28337 ^ new_n28333;
  assign new_n28364 = new_n28363 ^ new_n28352;
  assign new_n28365 = new_n28342 ^ new_n28333;
  assign new_n28366 = new_n28364 & new_n28365;
  assign new_n28367 = new_n28366 ^ new_n28355;
  assign new_n28368 = new_n28337 ^ new_n28330;
  assign new_n28369 = new_n28368 ^ new_n28367;
  assign new_n28370 = new_n28369 ^ new_n28362;
  assign new_n28371 = new_n28333 ^ new_n28329;
  assign new_n28372 = new_n28371 ^ new_n28352;
  assign new_n28373 = new_n28335 & new_n28372;
  assign new_n28374 = new_n28373 ^ new_n28336;
  assign new_n28375 = new_n28374 ^ new_n28335;
  assign new_n28376 = new_n28339 ^ new_n28335;
  assign new_n28377 = new_n28340 ^ new_n28329;
  assign new_n28378 = new_n28377 ^ new_n28352;
  assign new_n28379 = new_n28376 & new_n28378;
  assign new_n28380 = new_n28379 ^ new_n28342;
  assign new_n28381 = new_n28380 ^ new_n28367;
  assign new_n28382 = new_n28381 ^ new_n28375;
  assign new_n28383 = ~new_n28370 & new_n28382;
  assign new_n28384 = new_n28340 ^ new_n28333;
  assign new_n28385 = new_n28339 & new_n28384;
  assign new_n28386 = new_n28385 ^ new_n28333;
  assign new_n28387 = new_n28386 ^ new_n28374;
  assign new_n28388 = new_n28387 ^ new_n28383;
  assign new_n28389 = new_n28388 ^ new_n28357;
  assign new_n28390 = new_n28366 ^ new_n28354;
  assign new_n28391 = new_n28359 ^ new_n28346;
  assign new_n28392 = new_n28391 ^ new_n28390;
  assign new_n28393 = ~new_n28392 & new_n28389;
  assign new_n28394 = new_n28393 ^ new_n28383;
  assign new_n28395 = ~new_n28394 & new_n28358;
  assign new_n28396 = new_n28395 ^ new_n28358;
  assign new_n28397 = new_n28396 ^ new_n28370;
  assign new_n28398 = ~new_n28397 & new_n28335;
  assign new_n28399 = new_n28396 ^ new_n28393;
  assign new_n28400 = new_n28399 ^ new_n28392;
  assign new_n28401 = ~new_n28400 & new_n28376;
  assign new_n28402 = new_n28401 ^ new_n28398;
  assign new_n28403 = ~new_n28397 & new_n28372;
  assign new_n28404 = new_n28403 ^ new_n28402;
  assign new_n28405 = new_n28337 ^ new_n28332;
  assign new_n28406 = new_n28385 ^ new_n28379;
  assign new_n28407 = new_n28406 ^ new_n28390;
  assign new_n28408 = new_n28407 ^ new_n28405;
  assign new_n28409 = new_n28383 ^ new_n28358;
  assign new_n28410 = new_n28408 & new_n28409;
  assign new_n28411 = new_n28410 ^ new_n28387;
  assign new_n28412 = new_n28411 ^ new_n28357;
  assign new_n28413 = new_n28395 ^ new_n28383;
  assign new_n28414 = new_n28412 & new_n28413;
  assign new_n28415 = new_n28414 ^ new_n28410;
  assign new_n28416 = new_n28415 ^ new_n28382;
  assign new_n28417 = new_n28347 & new_n28416;
  assign new_n28418 = new_n28414 ^ new_n28408;
  assign new_n28419 = new_n28340 & new_n28418;
  assign new_n28420 = ~new_n28400 & new_n28378;
  assign new_n28421 = new_n28410 ^ new_n28393;
  assign new_n28422 = new_n28387 ^ new_n28351;
  assign new_n28423 = new_n28422 ^ new_n28421;
  assign new_n28424 = new_n28334 & new_n28423;
  assign new_n28425 = new_n28337 ^ new_n28329;
  assign new_n28426 = new_n28379 ^ new_n28360;
  assign new_n28427 = new_n28414 ^ new_n28396;
  assign new_n28428 = new_n28427 ^ new_n28426;
  assign new_n28429 = new_n28428 ^ new_n28425;
  assign new_n28430 = new_n28429 ^ new_n28333;
  assign new_n28431 = new_n28410 ^ new_n28349;
  assign new_n28432 = new_n28431 ^ new_n28374;
  assign new_n28433 = new_n28432 ^ new_n28430;
  assign new_n28434 = ~new_n28433 & new_n28365;
  assign new_n28435 = new_n28434 ^ new_n28424;
  assign new_n28436 = new_n28435 ^ new_n28420;
  assign new_n28437 = new_n28436 ^ new_n28419;
  assign new_n28438 = new_n28437 ^ new_n28417;
  assign new_n28439 = new_n28438 ^ new_n28404;
  assign new_n28440 = new_n28439 ^ new_n15343;
  assign new_n28441 = new_n28344 & new_n28423;
  assign new_n28442 = new_n28441 ^ new_n28424;
  assign new_n28443 = new_n28393 ^ new_n28332;
  assign new_n28444 = new_n28385 ^ new_n28346;
  assign new_n28445 = new_n28444 ^ new_n28429;
  assign new_n28446 = new_n28445 ^ new_n28443;
  assign new_n28447 = ~new_n28446 & new_n28352;
  assign new_n28448 = new_n28341 & new_n28412;
  assign new_n28449 = ~new_n28446 & new_n28353;
  assign new_n28450 = new_n28449 ^ new_n28448;
  assign new_n28451 = new_n28393 ^ new_n28358;
  assign new_n28452 = new_n28339 & new_n28451;
  assign new_n28453 = new_n28452 ^ new_n28398;
  assign new_n28454 = new_n28348 & new_n28416;
  assign new_n28455 = new_n28454 ^ new_n28453;
  assign new_n28456 = new_n28455 ^ new_n28450;
  assign new_n28457 = new_n28456 ^ new_n28447;
  assign new_n28458 = new_n28457 ^ new_n28442;
  assign new_n28459 = new_n28458 ^ new_n15312;
  assign new_n28460 = new_n28459 ^ new_n28440;
  assign new_n28461 = new_n28384 & new_n28451;
  assign new_n28462 = ~new_n28433 & new_n28364;
  assign new_n28463 = new_n28462 ^ new_n28438;
  assign new_n28464 = new_n28463 ^ new_n28461;
  assign new_n28465 = new_n28464 ^ new_n28456;
  assign new_n28466 = new_n28465 ^ new_n15364;
  assign new_n28467 = new_n28441 ^ new_n28403;
  assign new_n28468 = new_n28467 ^ new_n28463;
  assign new_n28469 = new_n28468 ^ new_n15337;
  assign new_n28470 = new_n28469 ^ new_n28466;
  assign new_n28471 = new_n28470 ^ new_n28460;
  assign new_n28472 = new_n28454 ^ new_n28449;
  assign new_n28473 = new_n28462 ^ new_n28419;
  assign new_n28474 = new_n28377 & new_n28418;
  assign new_n28475 = new_n28345 & new_n28412;
  assign new_n28476 = new_n28475 ^ new_n28474;
  assign new_n28477 = new_n28476 ^ new_n28435;
  assign new_n28478 = new_n28477 ^ new_n28473;
  assign new_n28479 = new_n28478 ^ new_n28472;
  assign new_n28480 = new_n28479 ^ new_n15322;
  assign new_n28481 = new_n28480 ^ new_n28459;
  assign new_n28482 = new_n28462 ^ new_n28441;
  assign new_n28483 = new_n28436 ^ new_n28404;
  assign new_n28484 = new_n28483 ^ new_n28482;
  assign new_n28485 = new_n28484 ^ new_n15315;
  assign new_n28486 = new_n28485 ^ new_n28459;
  assign new_n28487 = new_n28455 ^ new_n28417;
  assign new_n28488 = new_n28487 ^ new_n28477;
  assign new_n28489 = new_n28488 ^ new_n15353;
  assign new_n28490 = new_n28489 ^ new_n28486;
  assign new_n28491 = ~new_n28480 & ~new_n28490;
  assign new_n28492 = new_n28491 ^ new_n28480;
  assign new_n28493 = new_n28490 ^ new_n28480;
  assign new_n28494 = new_n28493 ^ new_n28470;
  assign new_n28495 = new_n28469 ^ new_n28440;
  assign new_n28496 = new_n28475 ^ new_n28403;
  assign new_n28497 = new_n28452 ^ new_n28401;
  assign new_n28498 = new_n28497 ^ new_n28437;
  assign new_n28499 = new_n28498 ^ new_n28496;
  assign new_n28500 = new_n28499 ^ new_n15329;
  assign new_n28501 = new_n28500 ^ new_n28480;
  assign new_n28502 = new_n28501 ^ new_n28495;
  assign new_n28503 = new_n28502 ^ new_n28489;
  assign new_n28504 = ~new_n28494 & new_n28503;
  assign new_n28505 = new_n28504 ^ new_n28492;
  assign new_n28506 = new_n28480 ^ new_n28440;
  assign new_n28507 = new_n28506 ^ new_n28470;
  assign new_n28508 = ~new_n28507 & new_n28502;
  assign new_n28509 = new_n28508 ^ new_n28485;
  assign new_n28510 = ~new_n28486 & new_n28489;
  assign new_n28511 = ~new_n28489 & new_n28440;
  assign new_n28512 = new_n28511 ^ new_n28510;
  assign new_n28513 = new_n28512 ^ new_n28509;
  assign new_n28514 = new_n28469 ^ new_n28459;
  assign new_n28515 = new_n28502 ^ new_n28486;
  assign new_n28516 = ~new_n28470 & new_n28515;
  assign new_n28517 = new_n28466 ^ new_n28440;
  assign new_n28518 = ~new_n28471 & new_n28517;
  assign new_n28519 = new_n28518 ^ new_n28516;
  assign new_n28520 = new_n28512 ^ new_n28440;
  assign new_n28521 = new_n28520 ^ new_n28504;
  assign new_n28522 = new_n28521 ^ new_n28519;
  assign new_n28523 = new_n28522 ^ new_n28514;
  assign new_n28524 = new_n28501 ^ new_n28466;
  assign new_n28525 = new_n28524 ^ new_n28485;
  assign new_n28526 = ~new_n28495 & ~new_n28525;
  assign new_n28527 = new_n28526 ^ new_n28516;
  assign new_n28528 = new_n28524 ^ new_n28459;
  assign new_n28529 = new_n28528 ^ new_n28527;
  assign new_n28530 = new_n28480 ^ new_n28469;
  assign new_n28531 = ~new_n28528 & ~new_n28530;
  assign new_n28532 = new_n28490 ^ new_n28469;
  assign new_n28533 = new_n28525 ^ new_n28489;
  assign new_n28534 = ~new_n28532 & ~new_n28533;
  assign new_n28535 = new_n28534 ^ new_n28531;
  assign new_n28536 = new_n28535 ^ new_n28469;
  assign new_n28537 = new_n28536 ^ new_n28529;
  assign new_n28538 = new_n28531 ^ new_n28492;
  assign new_n28539 = new_n28538 ^ new_n28470;
  assign new_n28540 = new_n28526 ^ new_n28518;
  assign new_n28541 = new_n28500 ^ new_n28459;
  assign new_n28542 = new_n28541 ^ new_n28540;
  assign new_n28543 = new_n28542 ^ new_n28539;
  assign new_n28544 = new_n28509 ^ new_n28502;
  assign new_n28545 = new_n28526 ^ new_n28504;
  assign new_n28546 = new_n28518 ^ new_n28466;
  assign new_n28547 = new_n28546 ^ new_n28545;
  assign new_n28548 = new_n28547 ^ new_n28544;
  assign new_n28549 = ~new_n28543 & new_n28548;
  assign new_n28550 = new_n28549 ^ new_n28537;
  assign new_n28551 = ~new_n28523 & new_n28550;
  assign new_n28552 = new_n28551 ^ new_n28513;
  assign new_n28553 = new_n28552 ^ new_n28529;
  assign new_n28554 = new_n28549 ^ new_n28513;
  assign new_n28555 = new_n28554 ^ new_n28529;
  assign new_n28556 = new_n28534 ^ new_n28491;
  assign new_n28557 = new_n28556 ^ new_n28519;
  assign new_n28558 = ~new_n28555 & ~new_n28557;
  assign new_n28559 = new_n28558 ^ new_n28549;
  assign new_n28560 = new_n28537 & new_n28559;
  assign new_n28561 = new_n28560 ^ new_n28550;
  assign new_n28562 = ~new_n28553 & new_n28561;
  assign new_n28563 = new_n28562 ^ new_n28560;
  assign new_n28564 = new_n28563 ^ new_n28505;
  assign new_n28565 = new_n28564 ^ new_n28481;
  assign new_n28566 = new_n28565 ^ new_n28440;
  assign new_n28567 = new_n28551 ^ new_n28531;
  assign new_n28568 = new_n28567 ^ new_n28509;
  assign new_n28569 = new_n28568 ^ new_n28566;
  assign new_n28570 = ~new_n28471 & ~new_n28569;
  assign new_n28571 = new_n28558 ^ new_n28551;
  assign new_n28572 = new_n28536 ^ new_n28513;
  assign new_n28573 = new_n28572 ^ new_n28571;
  assign new_n28574 = ~new_n28525 & ~new_n28573;
  assign new_n28575 = new_n28574 ^ new_n28570;
  assign new_n28576 = new_n28560 ^ new_n28558;
  assign new_n28577 = new_n28576 ^ new_n28557;
  assign new_n28578 = ~new_n28577 & new_n28503;
  assign new_n28579 = new_n28560 ^ new_n28543;
  assign new_n28580 = ~new_n28579 & new_n28502;
  assign new_n28581 = new_n28580 ^ new_n28578;
  assign new_n28582 = ~new_n28507 & ~new_n28579;
  assign new_n28583 = new_n28582 ^ new_n28581;
  assign new_n28584 = ~new_n28494 & ~new_n28577;
  assign new_n28585 = ~new_n28569 & new_n28517;
  assign new_n28586 = ~new_n28495 & ~new_n28573;
  assign new_n28587 = new_n28586 ^ new_n28585;
  assign new_n28588 = new_n28587 ^ new_n28584;
  assign new_n28589 = new_n28588 ^ new_n28583;
  assign new_n28590 = new_n28589 ^ new_n28575;
  assign new_n28591 = new_n28590 ^ new_n26036;
  assign new_n28592 = new_n28591 ^ new_n20014;
  assign new_n28593 = new_n28439 ^ new_n24876;
  assign new_n28594 = new_n28593 ^ new_n12869;
  assign new_n28595 = new_n27279 ^ new_n27256;
  assign new_n28596 = new_n28159 ^ new_n18922;
  assign new_n28597 = new_n28596 ^ new_n26263;
  assign new_n28598 = new_n28597 ^ new_n28595;
  assign new_n28599 = new_n28223 ^ new_n22385;
  assign new_n28600 = new_n28599 ^ new_n27256;
  assign new_n28601 = new_n27295 ^ new_n22423;
  assign new_n28602 = new_n28601 ^ new_n28600;
  assign new_n28603 = new_n28602 ^ new_n28598;
  assign new_n28604 = new_n28117 ^ new_n22288;
  assign new_n28605 = new_n27302 ^ new_n21072;
  assign new_n28606 = new_n28605 ^ new_n28604;
  assign new_n28607 = new_n27273 ^ new_n22308;
  assign new_n28608 = new_n27967 ^ new_n22427;
  assign new_n28609 = new_n28608 ^ new_n27256;
  assign new_n28610 = new_n28609 ^ new_n28607;
  assign new_n28611 = new_n28610 ^ new_n28606;
  assign new_n28612 = new_n28611 ^ new_n28603;
  assign new_n28613 = new_n28179 ^ new_n22450;
  assign new_n28614 = new_n27310 ^ new_n22274;
  assign new_n28615 = new_n28614 ^ new_n28613;
  assign new_n28616 = new_n28023 ^ new_n22342;
  assign new_n28617 = new_n27263 ^ new_n22441;
  assign new_n28618 = new_n28617 ^ new_n28616;
  assign new_n28619 = new_n28618 ^ new_n28615;
  assign new_n28620 = new_n28201 ^ new_n19999;
  assign new_n28621 = new_n27289 ^ new_n27256;
  assign new_n28622 = new_n28621 ^ new_n28620;
  assign new_n28623 = new_n28622 ^ new_n28619;
  assign new_n28624 = new_n28623 ^ new_n28606;
  assign new_n28625 = new_n28101 ^ new_n22466;
  assign new_n28626 = new_n28625 ^ new_n22476;
  assign new_n28627 = new_n28626 ^ new_n26214;
  assign new_n28628 = new_n28627 ^ new_n28603;
  assign new_n28629 = new_n28628 ^ new_n28615;
  assign new_n28630 = new_n28629 ^ new_n28622;
  assign new_n28631 = new_n28624 & new_n28630;
  assign new_n28632 = new_n28628 ^ new_n28618;
  assign new_n28633 = new_n28606 ^ new_n28598;
  assign new_n28634 = new_n28632 & new_n28633;
  assign new_n28635 = new_n28634 ^ new_n28631;
  assign new_n28636 = new_n28635 ^ new_n28606;
  assign new_n28637 = new_n28627 ^ new_n28606;
  assign new_n28638 = new_n28619 ^ new_n28612;
  assign new_n28639 = new_n28637 & new_n28638;
  assign new_n28640 = new_n28611 & new_n28629;
  assign new_n28641 = new_n28640 ^ new_n28639;
  assign new_n28642 = new_n28641 ^ new_n28632;
  assign new_n28643 = new_n28642 ^ new_n28636;
  assign new_n28644 = new_n28623 ^ new_n28610;
  assign new_n28645 = new_n28622 & new_n28644;
  assign new_n28646 = new_n28645 ^ new_n28610;
  assign new_n28647 = new_n28610 ^ new_n28598;
  assign new_n28648 = new_n28647 ^ new_n28637;
  assign new_n28649 = new_n28612 & new_n28648;
  assign new_n28650 = new_n28649 ^ new_n28615;
  assign new_n28651 = new_n28650 ^ new_n28646;
  assign new_n28652 = ~new_n28598 & ~new_n28623;
  assign new_n28653 = new_n28652 ^ new_n28598;
  assign new_n28654 = new_n28653 ^ new_n28634;
  assign new_n28655 = new_n28654 ^ new_n28637;
  assign new_n28656 = new_n28618 ^ new_n28610;
  assign new_n28657 = new_n28656 ^ new_n28637;
  assign new_n28658 = new_n28627 ^ new_n28610;
  assign new_n28659 = new_n28657 & new_n28658;
  assign new_n28660 = new_n28659 ^ new_n28640;
  assign new_n28661 = new_n28618 ^ new_n28602;
  assign new_n28662 = new_n28661 ^ new_n28660;
  assign new_n28663 = new_n28662 ^ new_n28655;
  assign new_n28664 = new_n28650 ^ new_n28612;
  assign new_n28665 = new_n28622 ^ new_n28612;
  assign new_n28666 = new_n28623 ^ new_n28598;
  assign new_n28667 = new_n28666 ^ new_n28637;
  assign new_n28668 = new_n28665 & new_n28667;
  assign new_n28669 = new_n28668 ^ new_n28640;
  assign new_n28670 = new_n28659 ^ new_n28627;
  assign new_n28671 = new_n28670 ^ new_n28669;
  assign new_n28672 = new_n28671 ^ new_n28664;
  assign new_n28673 = ~new_n28663 & new_n28672;
  assign new_n28674 = new_n28673 ^ new_n28651;
  assign new_n28675 = new_n28674 ^ new_n28642;
  assign new_n28676 = new_n28652 ^ new_n28631;
  assign new_n28677 = new_n28659 ^ new_n28639;
  assign new_n28678 = new_n28677 ^ new_n28676;
  assign new_n28679 = ~new_n28678 & new_n28675;
  assign new_n28680 = new_n28679 ^ new_n28673;
  assign new_n28681 = ~new_n28643 & ~new_n28680;
  assign new_n28682 = new_n28681 ^ new_n28679;
  assign new_n28683 = new_n28673 ^ new_n28643;
  assign new_n28684 = new_n28683 ^ new_n28682;
  assign new_n28685 = new_n28684 ^ new_n28663;
  assign new_n28686 = new_n28612 & new_n28685;
  assign new_n28687 = new_n28684 ^ new_n28679;
  assign new_n28688 = new_n28687 ^ new_n28678;
  assign new_n28689 = new_n28665 & new_n28688;
  assign new_n28690 = new_n28689 ^ new_n28686;
  assign new_n28691 = new_n28648 & new_n28685;
  assign new_n28692 = new_n28691 ^ new_n28690;
  assign new_n28693 = new_n28618 ^ new_n28606;
  assign new_n28694 = new_n28668 ^ new_n28645;
  assign new_n28695 = new_n28694 ^ new_n28677;
  assign new_n28696 = new_n28695 ^ new_n28693;
  assign new_n28697 = new_n28683 & new_n28696;
  assign new_n28698 = new_n28697 ^ new_n28651;
  assign new_n28699 = new_n28698 ^ new_n28642;
  assign new_n28700 = ~new_n28682 & new_n28699;
  assign new_n28701 = new_n28700 ^ new_n28697;
  assign new_n28702 = new_n28701 ^ new_n28672;
  assign new_n28703 = new_n28632 & new_n28702;
  assign new_n28704 = new_n28700 ^ new_n28696;
  assign new_n28705 = new_n28623 & new_n28704;
  assign new_n28706 = new_n28667 & new_n28688;
  assign new_n28707 = new_n28618 ^ new_n28598;
  assign new_n28708 = new_n28668 ^ new_n28653;
  assign new_n28709 = new_n28700 ^ new_n28684;
  assign new_n28710 = new_n28709 ^ new_n28708;
  assign new_n28711 = new_n28710 ^ new_n28707;
  assign new_n28712 = new_n28711 ^ new_n28610;
  assign new_n28713 = new_n28697 ^ new_n28634;
  assign new_n28714 = new_n28713 ^ new_n28650;
  assign new_n28715 = new_n28714 ^ new_n28712;
  assign new_n28716 = new_n28658 & new_n28715;
  assign new_n28717 = new_n28697 ^ new_n28679;
  assign new_n28718 = new_n28651 ^ new_n28636;
  assign new_n28719 = new_n28718 ^ new_n28717;
  assign new_n28720 = new_n28611 & new_n28719;
  assign new_n28721 = new_n28720 ^ new_n28716;
  assign new_n28722 = new_n28721 ^ new_n28706;
  assign new_n28723 = new_n28722 ^ new_n28705;
  assign new_n28724 = new_n28723 ^ new_n28703;
  assign new_n28725 = new_n28724 ^ new_n28692;
  assign new_n28726 = new_n26383 ^ new_n25774;
  assign new_n28727 = new_n28726 ^ new_n27751;
  assign new_n28728 = new_n21454 ^ new_n21185;
  assign new_n28729 = new_n28728 ^ new_n25794;
  assign new_n28730 = new_n28729 ^ new_n25730;
  assign new_n28731 = new_n28730 ^ new_n28727;
  assign new_n28732 = new_n25789 ^ new_n25705;
  assign new_n28733 = new_n28732 ^ new_n25753;
  assign new_n28734 = new_n22391 ^ new_n21448;
  assign new_n28735 = new_n28734 ^ new_n26383;
  assign new_n28736 = new_n28735 ^ new_n27722;
  assign new_n28737 = new_n28736 ^ new_n28733;
  assign new_n28738 = new_n28737 ^ new_n28731;
  assign new_n28739 = new_n27726 ^ new_n25307;
  assign new_n28740 = new_n22259 ^ new_n21467;
  assign new_n28741 = new_n28740 ^ new_n25692;
  assign new_n28742 = new_n28741 ^ new_n25676;
  assign new_n28743 = new_n28742 ^ new_n28739;
  assign new_n28744 = new_n22415 ^ new_n21471;
  assign new_n28745 = new_n28744 ^ new_n27765;
  assign new_n28746 = new_n28745 ^ new_n26383;
  assign new_n28747 = new_n25763 ^ new_n25645;
  assign new_n28748 = new_n28747 ^ new_n25705;
  assign new_n28749 = new_n28748 ^ new_n28746;
  assign new_n28750 = new_n28749 ^ new_n28743;
  assign new_n28751 = new_n28750 ^ new_n28738;
  assign new_n28752 = new_n27719 ^ new_n25622;
  assign new_n28753 = new_n22445 ^ new_n21461;
  assign new_n28754 = new_n28753 ^ new_n25676;
  assign new_n28755 = new_n28754 ^ new_n25582;
  assign new_n28756 = new_n28755 ^ new_n28752;
  assign new_n28757 = new_n27757 ^ new_n25582;
  assign new_n28758 = new_n22328 ^ new_n21487;
  assign new_n28759 = new_n28758 ^ new_n26391;
  assign new_n28760 = new_n28759 ^ new_n28757;
  assign new_n28761 = new_n28760 ^ new_n28756;
  assign new_n28762 = new_n22360 ^ new_n21491;
  assign new_n28763 = new_n28762 ^ new_n25730;
  assign new_n28764 = new_n27736 ^ new_n26383;
  assign new_n28765 = new_n28764 ^ new_n28763;
  assign new_n28766 = new_n28765 ^ new_n28761;
  assign new_n28767 = new_n28766 ^ new_n28743;
  assign new_n28768 = new_n27733 ^ new_n25716;
  assign new_n28769 = new_n22470 ^ new_n21442;
  assign new_n28770 = new_n28769 ^ new_n25753;
  assign new_n28771 = new_n28770 ^ new_n25794;
  assign new_n28772 = new_n28771 ^ new_n28768;
  assign new_n28773 = new_n28772 ^ new_n28738;
  assign new_n28774 = new_n28773 ^ new_n28756;
  assign new_n28775 = new_n28774 ^ new_n28765;
  assign new_n28776 = ~new_n28767 & ~new_n28775;
  assign new_n28777 = new_n28743 ^ new_n28731;
  assign new_n28778 = new_n28773 ^ new_n28760;
  assign new_n28779 = ~new_n28777 & new_n28778;
  assign new_n28780 = new_n28779 ^ new_n28776;
  assign new_n28781 = new_n28780 ^ new_n28743;
  assign new_n28782 = new_n28772 ^ new_n28743;
  assign new_n28783 = new_n28761 ^ new_n28751;
  assign new_n28784 = ~new_n28783 & new_n28782;
  assign new_n28785 = new_n28750 & new_n28774;
  assign new_n28786 = new_n28785 ^ new_n28784;
  assign new_n28787 = new_n28786 ^ new_n28778;
  assign new_n28788 = new_n28787 ^ new_n28781;
  assign new_n28789 = new_n28766 ^ new_n28749;
  assign new_n28790 = ~new_n28765 & ~new_n28789;
  assign new_n28791 = new_n28790 ^ new_n28749;
  assign new_n28792 = new_n28772 ^ new_n28749;
  assign new_n28793 = new_n28792 ^ new_n28777;
  assign new_n28794 = ~new_n28751 & ~new_n28793;
  assign new_n28795 = new_n28794 ^ new_n28756;
  assign new_n28796 = new_n28795 ^ new_n28791;
  assign new_n28797 = new_n28731 & new_n28766;
  assign new_n28798 = new_n28797 ^ new_n28731;
  assign new_n28799 = new_n28798 ^ new_n28779;
  assign new_n28800 = new_n28799 ^ new_n28782;
  assign new_n28801 = new_n28760 ^ new_n28749;
  assign new_n28802 = new_n28801 ^ new_n28782;
  assign new_n28803 = ~new_n28802 & new_n28792;
  assign new_n28804 = new_n28803 ^ new_n28785;
  assign new_n28805 = new_n28760 ^ new_n28737;
  assign new_n28806 = new_n28805 ^ new_n28804;
  assign new_n28807 = new_n28806 ^ new_n28800;
  assign new_n28808 = new_n28795 ^ new_n28751;
  assign new_n28809 = new_n28765 ^ new_n28751;
  assign new_n28810 = new_n28766 ^ new_n28731;
  assign new_n28811 = new_n28810 ^ new_n28782;
  assign new_n28812 = new_n28809 & new_n28811;
  assign new_n28813 = new_n28812 ^ new_n28785;
  assign new_n28814 = new_n28803 ^ new_n28772;
  assign new_n28815 = new_n28814 ^ new_n28813;
  assign new_n28816 = new_n28815 ^ new_n28808;
  assign new_n28817 = ~new_n28807 & new_n28816;
  assign new_n28818 = new_n28817 ^ new_n28796;
  assign new_n28819 = new_n28818 ^ new_n28787;
  assign new_n28820 = new_n28797 ^ new_n28776;
  assign new_n28821 = new_n28803 ^ new_n28784;
  assign new_n28822 = new_n28821 ^ new_n28820;
  assign new_n28823 = ~new_n28819 & ~new_n28822;
  assign new_n28824 = new_n28823 ^ new_n28817;
  assign new_n28825 = ~new_n28788 & ~new_n28824;
  assign new_n28826 = new_n28825 ^ new_n28823;
  assign new_n28827 = new_n28817 ^ new_n28788;
  assign new_n28828 = new_n28827 ^ new_n28826;
  assign new_n28829 = new_n28828 ^ new_n28807;
  assign new_n28830 = ~new_n28751 & new_n28829;
  assign new_n28831 = new_n28828 ^ new_n28823;
  assign new_n28832 = new_n28831 ^ new_n28822;
  assign new_n28833 = new_n28809 & new_n28832;
  assign new_n28834 = new_n28833 ^ new_n28830;
  assign new_n28835 = ~new_n28793 & new_n28829;
  assign new_n28836 = new_n28835 ^ new_n28834;
  assign new_n28837 = new_n28760 ^ new_n28743;
  assign new_n28838 = new_n28812 ^ new_n28790;
  assign new_n28839 = new_n28838 ^ new_n28821;
  assign new_n28840 = new_n28839 ^ new_n28837;
  assign new_n28841 = ~new_n28840 & new_n28827;
  assign new_n28842 = new_n28841 ^ new_n28796;
  assign new_n28843 = new_n28842 ^ new_n28787;
  assign new_n28844 = ~new_n28826 & ~new_n28843;
  assign new_n28845 = new_n28844 ^ new_n28841;
  assign new_n28846 = new_n28845 ^ new_n28816;
  assign new_n28847 = new_n28778 & new_n28846;
  assign new_n28848 = new_n28844 ^ new_n28840;
  assign new_n28849 = ~new_n28766 & ~new_n28848;
  assign new_n28850 = new_n28811 & new_n28832;
  assign new_n28851 = new_n28760 ^ new_n28731;
  assign new_n28852 = new_n28812 ^ new_n28798;
  assign new_n28853 = new_n28844 ^ new_n28828;
  assign new_n28854 = new_n28853 ^ new_n28852;
  assign new_n28855 = new_n28854 ^ new_n28851;
  assign new_n28856 = new_n28855 ^ new_n28749;
  assign new_n28857 = new_n28841 ^ new_n28779;
  assign new_n28858 = new_n28857 ^ new_n28795;
  assign new_n28859 = new_n28858 ^ new_n28856;
  assign new_n28860 = new_n28792 & new_n28859;
  assign new_n28861 = new_n28841 ^ new_n28823;
  assign new_n28862 = new_n28796 ^ new_n28781;
  assign new_n28863 = new_n28862 ^ new_n28861;
  assign new_n28864 = ~new_n28863 & new_n28750;
  assign new_n28865 = new_n28864 ^ new_n28860;
  assign new_n28866 = new_n28865 ^ new_n28850;
  assign new_n28867 = new_n28866 ^ new_n28849;
  assign new_n28868 = new_n28867 ^ new_n28847;
  assign new_n28869 = new_n28868 ^ new_n28836;
  assign new_n28870 = new_n28869 ^ new_n28725;
  assign new_n28871 = new_n28870 ^ new_n28594;
  assign new_n28872 = new_n24628 ^ new_n24592;
  assign new_n28873 = new_n28342 ^ new_n24566;
  assign new_n28874 = new_n28873 ^ new_n24622;
  assign new_n28875 = new_n28874 ^ new_n28872;
  assign new_n28876 = new_n27408 ^ new_n24467;
  assign new_n28877 = new_n28876 ^ new_n24587;
  assign new_n28878 = new_n28329 ^ new_n24622;
  assign new_n28879 = new_n28878 ^ new_n24603;
  assign new_n28880 = new_n28879 ^ new_n28877;
  assign new_n28881 = new_n24566 ^ new_n24508;
  assign new_n28882 = new_n28881 ^ new_n24613;
  assign new_n28883 = new_n28330 ^ new_n27408;
  assign new_n28884 = new_n28883 ^ new_n24576;
  assign new_n28885 = new_n28884 ^ new_n28882;
  assign new_n28886 = new_n28885 ^ new_n28880;
  assign new_n28887 = new_n28886 ^ new_n28875;
  assign new_n28888 = new_n28336 ^ new_n24456;
  assign new_n28889 = new_n27450 ^ new_n24538;
  assign new_n28890 = new_n28889 ^ new_n28888;
  assign new_n28891 = new_n28890 ^ new_n28887;
  assign new_n28892 = new_n28332 ^ new_n24546;
  assign new_n28893 = new_n27435 ^ new_n24500;
  assign new_n28894 = new_n28893 ^ new_n28892;
  assign new_n28895 = new_n28337 ^ new_n24374;
  assign new_n28896 = new_n27414 ^ new_n24395;
  assign new_n28897 = new_n28896 ^ new_n28895;
  assign new_n28898 = new_n28897 ^ new_n28894;
  assign new_n28899 = new_n28333 ^ new_n27408;
  assign new_n28900 = new_n28899 ^ new_n23967;
  assign new_n28901 = new_n27430 ^ new_n24524;
  assign new_n28902 = new_n28901 ^ new_n28900;
  assign new_n28903 = new_n28902 ^ new_n28894;
  assign new_n28904 = new_n28903 ^ new_n28886;
  assign new_n28905 = new_n28339 ^ new_n24603;
  assign new_n28906 = new_n27408 ^ new_n24492;
  assign new_n28907 = new_n28906 ^ new_n28905;
  assign new_n28908 = new_n28907 ^ new_n28904;
  assign new_n28909 = new_n28897 ^ new_n28890;
  assign new_n28910 = new_n28909 ^ new_n28907;
  assign new_n28911 = new_n28910 ^ new_n28880;
  assign new_n28912 = new_n28894 ^ new_n28875;
  assign new_n28913 = new_n28912 ^ new_n28911;
  assign new_n28914 = new_n28908 & new_n28913;
  assign new_n28915 = new_n28910 ^ new_n28902;
  assign new_n28916 = ~new_n28907 & ~new_n28915;
  assign new_n28917 = new_n28916 ^ new_n28914;
  assign new_n28918 = new_n28909 ^ new_n28904;
  assign new_n28919 = ~new_n28918 & new_n28912;
  assign new_n28920 = new_n28902 ^ new_n28875;
  assign new_n28921 = new_n28902 ^ new_n28897;
  assign new_n28922 = new_n28921 ^ new_n28912;
  assign new_n28923 = ~new_n28922 & new_n28920;
  assign new_n28924 = new_n28923 ^ new_n28919;
  assign new_n28925 = new_n28924 ^ new_n28917;
  assign new_n28926 = new_n28925 ^ new_n28898;
  assign new_n28927 = new_n28910 ^ new_n28894;
  assign new_n28928 = new_n28907 ^ new_n28891;
  assign new_n28929 = ~new_n28927 & ~new_n28928;
  assign new_n28930 = new_n28894 ^ new_n28880;
  assign new_n28931 = new_n28897 ^ new_n28887;
  assign new_n28932 = ~new_n28930 & new_n28931;
  assign new_n28933 = new_n28932 ^ new_n28929;
  assign new_n28934 = new_n28933 ^ new_n28894;
  assign new_n28935 = new_n28891 & new_n28903;
  assign new_n28936 = new_n28935 ^ new_n28919;
  assign new_n28937 = new_n28936 ^ new_n28931;
  assign new_n28938 = new_n28937 ^ new_n28934;
  assign new_n28939 = new_n28880 & new_n28910;
  assign new_n28940 = new_n28939 ^ new_n28880;
  assign new_n28941 = new_n28940 ^ new_n28932;
  assign new_n28942 = new_n28941 ^ new_n28912;
  assign new_n28943 = new_n28935 ^ new_n28923;
  assign new_n28944 = new_n28897 ^ new_n28885;
  assign new_n28945 = new_n28944 ^ new_n28943;
  assign new_n28946 = new_n28945 ^ new_n28942;
  assign new_n28947 = new_n28930 ^ new_n28920;
  assign new_n28948 = ~new_n28904 & ~new_n28947;
  assign new_n28949 = new_n28948 ^ new_n28890;
  assign new_n28950 = new_n28949 ^ new_n28904;
  assign new_n28951 = new_n28943 ^ new_n28914;
  assign new_n28952 = new_n28951 ^ new_n28875;
  assign new_n28953 = new_n28952 ^ new_n28950;
  assign new_n28954 = ~new_n28946 & new_n28953;
  assign new_n28955 = new_n28954 ^ new_n28938;
  assign new_n28956 = ~new_n28926 & new_n28955;
  assign new_n28957 = new_n28916 ^ new_n28902;
  assign new_n28958 = new_n28957 ^ new_n28949;
  assign new_n28959 = new_n28958 ^ new_n28954;
  assign new_n28960 = new_n28959 ^ new_n28937;
  assign new_n28961 = new_n28939 ^ new_n28929;
  assign new_n28962 = new_n28961 ^ new_n28924;
  assign new_n28963 = ~new_n28960 & ~new_n28962;
  assign new_n28964 = new_n28963 ^ new_n28956;
  assign new_n28965 = new_n28958 ^ new_n28934;
  assign new_n28966 = new_n28965 ^ new_n28964;
  assign new_n28967 = ~new_n28966 & new_n28891;
  assign new_n28968 = new_n28963 ^ new_n28954;
  assign new_n28969 = new_n28938 & new_n28968;
  assign new_n28970 = new_n28969 ^ new_n28946;
  assign new_n28971 = ~new_n28947 & ~new_n28970;
  assign new_n28972 = new_n28971 ^ new_n28967;
  assign new_n28973 = new_n28897 ^ new_n28880;
  assign new_n28974 = new_n28940 ^ new_n28914;
  assign new_n28975 = new_n28958 ^ new_n28956;
  assign new_n28976 = new_n28975 ^ new_n28937;
  assign new_n28977 = new_n28969 ^ new_n28955;
  assign new_n28978 = ~new_n28976 & new_n28977;
  assign new_n28979 = new_n28978 ^ new_n28969;
  assign new_n28980 = new_n28979 ^ new_n28974;
  assign new_n28981 = new_n28980 ^ new_n28973;
  assign new_n28982 = new_n28981 ^ new_n28902;
  assign new_n28983 = new_n28956 ^ new_n28932;
  assign new_n28984 = new_n28983 ^ new_n28949;
  assign new_n28985 = new_n28984 ^ new_n28982;
  assign new_n28986 = ~new_n28922 & ~new_n28985;
  assign new_n28987 = new_n28978 ^ new_n28956;
  assign new_n28988 = new_n28987 ^ new_n28953;
  assign new_n28989 = new_n28931 & new_n28988;
  assign new_n28990 = new_n28978 ^ new_n28926;
  assign new_n28991 = ~new_n28910 & ~new_n28990;
  assign new_n28992 = new_n28969 ^ new_n28963;
  assign new_n28993 = new_n28992 ^ new_n28962;
  assign new_n28994 = ~new_n28993 & new_n28913;
  assign new_n28995 = ~new_n28985 & new_n28920;
  assign new_n28996 = ~new_n28966 & new_n28903;
  assign new_n28997 = new_n28996 ^ new_n28995;
  assign new_n28998 = new_n28997 ^ new_n28994;
  assign new_n28999 = new_n28998 ^ new_n28991;
  assign new_n29000 = new_n28999 ^ new_n28989;
  assign new_n29001 = new_n29000 ^ new_n28986;
  assign new_n29002 = new_n29001 ^ new_n28972;
  assign new_n29003 = new_n23553 ^ new_n23547;
  assign new_n29004 = new_n24902 ^ new_n18670;
  assign new_n29005 = new_n29004 ^ new_n13172;
  assign new_n29006 = new_n29005 ^ new_n23490;
  assign new_n29007 = new_n29006 ^ new_n23528;
  assign new_n29008 = new_n29007 ^ new_n29003;
  assign new_n29009 = new_n23517 ^ new_n23507;
  assign new_n29010 = new_n23462 ^ new_n23418;
  assign new_n29011 = new_n29010 ^ new_n29009;
  assign new_n29012 = new_n24889 ^ new_n18634;
  assign new_n29013 = new_n29012 ^ new_n13185;
  assign new_n29014 = new_n29013 ^ new_n23395;
  assign new_n29015 = new_n29014 ^ new_n23547;
  assign new_n29016 = new_n29015 ^ new_n29011;
  assign new_n29017 = new_n23490 ^ new_n23427;
  assign new_n29018 = new_n29017 ^ new_n23542;
  assign new_n29019 = new_n24884 ^ new_n18793;
  assign new_n29020 = new_n29019 ^ new_n13216;
  assign new_n29021 = new_n29020 ^ new_n23500;
  assign new_n29022 = new_n29021 ^ new_n29010;
  assign new_n29023 = new_n29022 ^ new_n29018;
  assign new_n29024 = new_n29023 ^ new_n29016;
  assign new_n29025 = new_n29024 ^ new_n29008;
  assign new_n29026 = new_n24840 ^ new_n18765;
  assign new_n29027 = new_n29026 ^ new_n13207;
  assign new_n29028 = new_n29027 ^ new_n22835;
  assign new_n29029 = new_n29028 ^ new_n23466;
  assign new_n29030 = new_n23374 ^ new_n23350;
  assign new_n29031 = new_n29030 ^ new_n29029;
  assign new_n29032 = new_n29031 ^ new_n29025;
  assign new_n29033 = new_n23471 ^ new_n23466;
  assign new_n29034 = new_n24894 ^ new_n17678;
  assign new_n29035 = new_n29034 ^ new_n13177;
  assign new_n29036 = new_n29035 ^ new_n23418;
  assign new_n29037 = new_n29036 ^ new_n23331;
  assign new_n29038 = new_n29037 ^ new_n29033;
  assign new_n29039 = new_n24860 ^ new_n18718;
  assign new_n29040 = new_n29039 ^ new_n13202;
  assign new_n29041 = new_n29040 ^ new_n27610;
  assign new_n29042 = new_n23350 ^ new_n23291;
  assign new_n29043 = new_n29042 ^ new_n29041;
  assign new_n29044 = new_n29043 ^ new_n29038;
  assign new_n29045 = new_n24876 ^ new_n18771;
  assign new_n29046 = new_n29045 ^ new_n13189;
  assign new_n29047 = new_n29046 ^ new_n23437;
  assign new_n29048 = new_n29047 ^ new_n29010;
  assign new_n29049 = new_n23427 ^ new_n22980;
  assign new_n29050 = new_n29049 ^ new_n23484;
  assign new_n29051 = new_n29050 ^ new_n29048;
  assign new_n29052 = new_n29051 ^ new_n29038;
  assign new_n29053 = new_n29052 ^ new_n29024;
  assign new_n29054 = new_n24870 ^ new_n18823;
  assign new_n29055 = new_n29054 ^ new_n13197;
  assign new_n29056 = new_n29055 ^ new_n23507;
  assign new_n29057 = new_n29010 ^ new_n23411;
  assign new_n29058 = new_n29057 ^ new_n29056;
  assign new_n29059 = new_n29058 ^ new_n29053;
  assign new_n29060 = new_n29043 ^ new_n29031;
  assign new_n29061 = new_n29060 ^ new_n29058;
  assign new_n29062 = new_n29061 ^ new_n29016;
  assign new_n29063 = new_n29038 ^ new_n29008;
  assign new_n29064 = new_n29063 ^ new_n29062;
  assign new_n29065 = ~new_n29059 & new_n29064;
  assign new_n29066 = new_n29061 ^ new_n29051;
  assign new_n29067 = ~new_n29058 & ~new_n29066;
  assign new_n29068 = new_n29067 ^ new_n29065;
  assign new_n29069 = new_n29060 ^ new_n29053;
  assign new_n29070 = ~new_n29063 & new_n29069;
  assign new_n29071 = new_n29051 ^ new_n29008;
  assign new_n29072 = new_n29051 ^ new_n29043;
  assign new_n29073 = new_n29072 ^ new_n29063;
  assign new_n29074 = ~new_n29071 & ~new_n29073;
  assign new_n29075 = new_n29074 ^ new_n29070;
  assign new_n29076 = new_n29075 ^ new_n29068;
  assign new_n29077 = new_n29076 ^ new_n29044;
  assign new_n29078 = new_n29061 ^ new_n29038;
  assign new_n29079 = new_n29058 ^ new_n29032;
  assign new_n29080 = ~new_n29078 & new_n29079;
  assign new_n29081 = new_n29043 ^ new_n29025;
  assign new_n29082 = new_n29038 ^ new_n29016;
  assign new_n29083 = ~new_n29081 & new_n29082;
  assign new_n29084 = new_n29083 ^ new_n29080;
  assign new_n29085 = new_n29084 ^ new_n29038;
  assign new_n29086 = ~new_n29032 & new_n29052;
  assign new_n29087 = new_n29086 ^ new_n29070;
  assign new_n29088 = new_n29087 ^ new_n29081;
  assign new_n29089 = new_n29088 ^ new_n29085;
  assign new_n29090 = ~new_n29016 & new_n29061;
  assign new_n29091 = new_n29090 ^ new_n29016;
  assign new_n29092 = new_n29091 ^ new_n29083;
  assign new_n29093 = new_n29092 ^ new_n29063;
  assign new_n29094 = new_n29086 ^ new_n29074;
  assign new_n29095 = new_n29043 ^ new_n29023;
  assign new_n29096 = new_n29095 ^ new_n29094;
  assign new_n29097 = new_n29096 ^ new_n29093;
  assign new_n29098 = new_n29051 ^ new_n29016;
  assign new_n29099 = new_n29098 ^ new_n29063;
  assign new_n29100 = ~new_n29099 & new_n29053;
  assign new_n29101 = new_n29100 ^ new_n29031;
  assign new_n29102 = new_n29101 ^ new_n29053;
  assign new_n29103 = new_n29065 ^ new_n29008;
  assign new_n29104 = new_n29103 ^ new_n29094;
  assign new_n29105 = new_n29104 ^ new_n29102;
  assign new_n29106 = ~new_n29105 & new_n29097;
  assign new_n29107 = new_n29106 ^ new_n29089;
  assign new_n29108 = ~new_n29107 & new_n29077;
  assign new_n29109 = new_n29067 ^ new_n29051;
  assign new_n29110 = new_n29109 ^ new_n29101;
  assign new_n29111 = new_n29110 ^ new_n29106;
  assign new_n29112 = new_n29111 ^ new_n29088;
  assign new_n29113 = new_n29090 ^ new_n29080;
  assign new_n29114 = new_n29113 ^ new_n29075;
  assign new_n29115 = ~new_n29112 & ~new_n29114;
  assign new_n29116 = new_n29115 ^ new_n29108;
  assign new_n29117 = new_n29110 ^ new_n29085;
  assign new_n29118 = new_n29117 ^ new_n29116;
  assign new_n29119 = ~new_n29032 & new_n29118;
  assign new_n29120 = new_n29115 ^ new_n29106;
  assign new_n29121 = ~new_n29089 & new_n29120;
  assign new_n29122 = new_n29121 ^ new_n29097;
  assign new_n29123 = ~new_n29099 & new_n29122;
  assign new_n29124 = new_n29123 ^ new_n29119;
  assign new_n29125 = new_n29043 ^ new_n29016;
  assign new_n29126 = new_n29091 ^ new_n29065;
  assign new_n29127 = new_n29110 ^ new_n29108;
  assign new_n29128 = new_n29127 ^ new_n29088;
  assign new_n29129 = new_n29121 ^ new_n29107;
  assign new_n29130 = ~new_n29128 & ~new_n29129;
  assign new_n29131 = new_n29130 ^ new_n29121;
  assign new_n29132 = new_n29131 ^ new_n29126;
  assign new_n29133 = new_n29132 ^ new_n29125;
  assign new_n29134 = new_n29133 ^ new_n29051;
  assign new_n29135 = new_n29108 ^ new_n29083;
  assign new_n29136 = new_n29135 ^ new_n29101;
  assign new_n29137 = new_n29136 ^ new_n29134;
  assign new_n29138 = ~new_n29073 & ~new_n29137;
  assign new_n29139 = new_n29130 ^ new_n29108;
  assign new_n29140 = new_n29139 ^ new_n29105;
  assign new_n29141 = ~new_n29081 & ~new_n29140;
  assign new_n29142 = new_n29130 ^ new_n29077;
  assign new_n29143 = ~new_n29061 & new_n29142;
  assign new_n29144 = new_n29121 ^ new_n29115;
  assign new_n29145 = new_n29144 ^ new_n29114;
  assign new_n29146 = ~new_n29145 & new_n29064;
  assign new_n29147 = new_n29052 & new_n29118;
  assign new_n29148 = ~new_n29071 & ~new_n29137;
  assign new_n29149 = new_n29148 ^ new_n29147;
  assign new_n29150 = new_n29149 ^ new_n29146;
  assign new_n29151 = new_n29150 ^ new_n29143;
  assign new_n29152 = new_n29151 ^ new_n29141;
  assign new_n29153 = new_n29152 ^ new_n29138;
  assign new_n29154 = new_n29153 ^ new_n29124;
  assign new_n29155 = new_n29154 ^ new_n29002;
  assign new_n29156 = new_n29155 ^ new_n28871;
  assign new_n29157 = ~new_n29128 & new_n29079;
  assign new_n29158 = new_n29157 ^ new_n29123;
  assign new_n29159 = ~new_n29059 & ~new_n29145;
  assign new_n29160 = new_n29115 ^ new_n29089;
  assign new_n29161 = ~new_n29058 & ~new_n29160;
  assign new_n29162 = new_n29161 ^ new_n29159;
  assign new_n29163 = new_n29162 ^ new_n29151;
  assign new_n29164 = new_n29163 ^ new_n29158;
  assign new_n29165 = ~new_n28993 & new_n28908;
  assign new_n29166 = ~new_n28904 & ~new_n28970;
  assign new_n29167 = new_n29166 ^ new_n29165;
  assign new_n29168 = new_n29167 ^ new_n28971;
  assign new_n29169 = new_n29168 ^ new_n29000;
  assign new_n29170 = ~new_n28928 & ~new_n28976;
  assign new_n29171 = new_n29170 ^ new_n28971;
  assign new_n29172 = new_n28963 ^ new_n28938;
  assign new_n29173 = ~new_n28907 & new_n29172;
  assign new_n29174 = new_n29173 ^ new_n29165;
  assign new_n29175 = new_n29174 ^ new_n28999;
  assign new_n29176 = new_n29175 ^ new_n29171;
  assign new_n29177 = new_n29176 ^ new_n29169;
  assign new_n29178 = new_n29177 ^ new_n29164;
  assign new_n29179 = new_n29178 ^ new_n29156;
  assign new_n29180 = new_n28996 ^ new_n28967;
  assign new_n29181 = new_n28963 ^ new_n28894;
  assign new_n29182 = new_n28929 ^ new_n28916;
  assign new_n29183 = new_n29182 ^ new_n28981;
  assign new_n29184 = new_n29183 ^ new_n29181;
  assign new_n29185 = new_n28912 & new_n29184;
  assign new_n29186 = ~new_n28918 & new_n29184;
  assign new_n29187 = ~new_n28927 & ~new_n28976;
  assign new_n29188 = new_n29187 ^ new_n29186;
  assign new_n29189 = ~new_n28930 & new_n28988;
  assign new_n29190 = new_n29173 ^ new_n29166;
  assign new_n29191 = new_n29190 ^ new_n29189;
  assign new_n29192 = new_n29191 ^ new_n29188;
  assign new_n29193 = new_n29192 ^ new_n29185;
  assign new_n29194 = new_n29193 ^ new_n29180;
  assign new_n29195 = new_n28629 & new_n28719;
  assign new_n29196 = new_n29195 ^ new_n28720;
  assign new_n29197 = new_n28679 ^ new_n28606;
  assign new_n29198 = new_n28645 ^ new_n28631;
  assign new_n29199 = new_n29198 ^ new_n28711;
  assign new_n29200 = new_n29199 ^ new_n29197;
  assign new_n29201 = new_n28637 & new_n29200;
  assign new_n29202 = new_n28624 & new_n28699;
  assign new_n29203 = new_n28638 & new_n29200;
  assign new_n29204 = new_n29203 ^ new_n29202;
  assign new_n29205 = new_n28679 ^ new_n28643;
  assign new_n29206 = new_n28622 & new_n29205;
  assign new_n29207 = new_n29206 ^ new_n28686;
  assign new_n29208 = new_n28633 & new_n28702;
  assign new_n29209 = new_n29208 ^ new_n29207;
  assign new_n29210 = new_n29209 ^ new_n29204;
  assign new_n29211 = new_n29210 ^ new_n29201;
  assign new_n29212 = new_n29211 ^ new_n29196;
  assign new_n29213 = ~new_n28863 & new_n28774;
  assign new_n29214 = new_n29213 ^ new_n28864;
  assign new_n29215 = new_n28823 ^ new_n28743;
  assign new_n29216 = new_n28790 ^ new_n28776;
  assign new_n29217 = new_n29216 ^ new_n28855;
  assign new_n29218 = new_n29217 ^ new_n29215;
  assign new_n29219 = ~new_n29218 & new_n28782;
  assign new_n29220 = ~new_n28767 & ~new_n28843;
  assign new_n29221 = ~new_n28783 & ~new_n29218;
  assign new_n29222 = new_n29221 ^ new_n29220;
  assign new_n29223 = new_n28823 ^ new_n28788;
  assign new_n29224 = ~new_n28765 & new_n29223;
  assign new_n29225 = new_n29224 ^ new_n28830;
  assign new_n29226 = ~new_n28777 & new_n28846;
  assign new_n29227 = new_n29226 ^ new_n29225;
  assign new_n29228 = new_n29227 ^ new_n29222;
  assign new_n29229 = new_n29228 ^ new_n29219;
  assign new_n29230 = new_n29229 ^ new_n29214;
  assign new_n29231 = new_n29230 ^ new_n29212;
  assign new_n29232 = new_n29231 ^ new_n29194;
  assign new_n29233 = new_n28458 ^ new_n24860;
  assign new_n29234 = new_n29233 ^ new_n13551;
  assign new_n29235 = new_n29053 & new_n29122;
  assign new_n29236 = new_n29235 ^ new_n29159;
  assign new_n29237 = new_n29236 ^ new_n29123;
  assign new_n29238 = new_n29237 ^ new_n29152;
  assign new_n29239 = new_n29238 ^ new_n29169;
  assign new_n29240 = new_n29239 ^ new_n29234;
  assign new_n29241 = new_n29240 ^ new_n29232;
  assign new_n29242 = new_n29241 ^ new_n29179;
  assign new_n29243 = new_n29195 ^ new_n28691;
  assign new_n29244 = new_n28657 & new_n28715;
  assign new_n29245 = new_n29244 ^ new_n28724;
  assign new_n29246 = new_n29245 ^ new_n29243;
  assign new_n29247 = new_n29213 ^ new_n28835;
  assign new_n29248 = ~new_n28802 & new_n28859;
  assign new_n29249 = new_n29248 ^ new_n28868;
  assign new_n29250 = new_n29249 ^ new_n29247;
  assign new_n29251 = new_n29250 ^ new_n29246;
  assign new_n29252 = new_n28986 ^ new_n28967;
  assign new_n29253 = new_n29168 ^ new_n28998;
  assign new_n29254 = new_n29253 ^ new_n29252;
  assign new_n29255 = new_n29254 ^ new_n29251;
  assign new_n29256 = new_n29138 ^ new_n29119;
  assign new_n29257 = new_n29237 ^ new_n29150;
  assign new_n29258 = new_n29257 ^ new_n29256;
  assign new_n29259 = new_n28468 ^ new_n24894;
  assign new_n29260 = new_n29259 ^ new_n13714;
  assign new_n29261 = new_n29260 ^ new_n29002;
  assign new_n29262 = new_n29261 ^ new_n29258;
  assign new_n29263 = new_n29262 ^ new_n29255;
  assign new_n29264 = new_n28644 & new_n29205;
  assign new_n29265 = new_n29264 ^ new_n29245;
  assign new_n29266 = new_n29265 ^ new_n29210;
  assign new_n29267 = ~new_n28789 & new_n29223;
  assign new_n29268 = new_n29267 ^ new_n29249;
  assign new_n29269 = new_n29268 ^ new_n29228;
  assign new_n29270 = new_n29269 ^ new_n29266;
  assign new_n29271 = new_n29189 ^ new_n29186;
  assign new_n29272 = ~new_n28990 & new_n28911;
  assign new_n29273 = new_n29272 ^ new_n29170;
  assign new_n29274 = new_n29273 ^ new_n28997;
  assign new_n29275 = new_n28991 ^ new_n28986;
  assign new_n29276 = new_n29275 ^ new_n29274;
  assign new_n29277 = new_n29276 ^ new_n29271;
  assign new_n29278 = new_n29277 ^ new_n29270;
  assign new_n29279 = ~new_n29140 & new_n29082;
  assign new_n29280 = new_n29115 ^ new_n29038;
  assign new_n29281 = new_n29080 ^ new_n29067;
  assign new_n29282 = new_n29281 ^ new_n29133;
  assign new_n29283 = new_n29282 ^ new_n29280;
  assign new_n29284 = ~new_n29283 & new_n29069;
  assign new_n29285 = new_n29284 ^ new_n29279;
  assign new_n29286 = new_n29143 ^ new_n29138;
  assign new_n29287 = ~new_n29062 & new_n29142;
  assign new_n29288 = new_n29287 ^ new_n29157;
  assign new_n29289 = new_n29288 ^ new_n29149;
  assign new_n29290 = new_n29289 ^ new_n29286;
  assign new_n29291 = new_n29290 ^ new_n29285;
  assign new_n29292 = new_n28465 ^ new_n24902;
  assign new_n29293 = new_n29292 ^ new_n13670;
  assign new_n29294 = ~new_n28915 & new_n29172;
  assign new_n29295 = new_n29294 ^ new_n29001;
  assign new_n29296 = new_n29295 ^ new_n29192;
  assign new_n29297 = new_n29296 ^ new_n29293;
  assign new_n29298 = new_n29297 ^ new_n29291;
  assign new_n29299 = new_n29298 ^ new_n29278;
  assign new_n29300 = new_n29299 ^ new_n29263;
  assign new_n29301 = new_n29300 ^ new_n29242;
  assign new_n29302 = new_n29208 ^ new_n29203;
  assign new_n29303 = new_n29244 ^ new_n28705;
  assign new_n29304 = new_n28666 & new_n28704;
  assign new_n29305 = new_n28630 & new_n28699;
  assign new_n29306 = new_n29305 ^ new_n29304;
  assign new_n29307 = new_n29306 ^ new_n28721;
  assign new_n29308 = new_n29307 ^ new_n29303;
  assign new_n29309 = new_n29308 ^ new_n29302;
  assign new_n29310 = new_n29226 ^ new_n29221;
  assign new_n29311 = new_n29248 ^ new_n28849;
  assign new_n29312 = ~new_n28848 & new_n28810;
  assign new_n29313 = ~new_n28775 & ~new_n28843;
  assign new_n29314 = new_n29313 ^ new_n29312;
  assign new_n29315 = new_n29314 ^ new_n28865;
  assign new_n29316 = new_n29315 ^ new_n29311;
  assign new_n29317 = new_n29316 ^ new_n29310;
  assign new_n29318 = new_n29317 ^ new_n29309;
  assign new_n29319 = new_n29191 ^ new_n28989;
  assign new_n29320 = new_n29319 ^ new_n29274;
  assign new_n29321 = new_n29320 ^ new_n29318;
  assign new_n29322 = new_n29321 ^ new_n29155;
  assign new_n29323 = new_n28479 ^ new_n24889;
  assign new_n29324 = new_n29323 ^ new_n13641;
  assign new_n29325 = new_n29235 ^ new_n29161;
  assign new_n29326 = new_n29325 ^ new_n29279;
  assign new_n29327 = new_n29326 ^ new_n29141;
  assign new_n29328 = new_n29327 ^ new_n29289;
  assign new_n29329 = new_n29328 ^ new_n29324;
  assign new_n29330 = new_n29329 ^ new_n29277;
  assign new_n29331 = new_n29330 ^ new_n29322;
  assign new_n29332 = new_n29331 ^ new_n29241;
  assign new_n29333 = new_n28484 ^ new_n24840;
  assign new_n29334 = new_n29333 ^ new_n13573;
  assign new_n29335 = new_n29147 ^ new_n29119;
  assign new_n29336 = ~new_n29063 & ~new_n29283;
  assign new_n29337 = ~new_n29078 & ~new_n29128;
  assign new_n29338 = new_n29337 ^ new_n29284;
  assign new_n29339 = new_n29338 ^ new_n29326;
  assign new_n29340 = new_n29339 ^ new_n29336;
  assign new_n29341 = new_n29340 ^ new_n29335;
  assign new_n29342 = new_n29341 ^ new_n29334;
  assign new_n29343 = new_n29342 ^ new_n29254;
  assign new_n29344 = new_n29244 ^ new_n29195;
  assign new_n29345 = new_n28722 ^ new_n28692;
  assign new_n29346 = new_n29345 ^ new_n29344;
  assign new_n29347 = new_n29248 ^ new_n29213;
  assign new_n29348 = new_n28866 ^ new_n28836;
  assign new_n29349 = new_n29348 ^ new_n29347;
  assign new_n29350 = new_n29349 ^ new_n29346;
  assign new_n29351 = new_n29350 ^ new_n29194;
  assign new_n29352 = new_n29351 ^ new_n29343;
  assign new_n29353 = new_n29352 ^ new_n29241;
  assign new_n29354 = new_n28488 ^ new_n24870;
  assign new_n29355 = new_n29354 ^ new_n13602;
  assign new_n29356 = new_n29355 ^ new_n29320;
  assign new_n29357 = new_n29209 ^ new_n28703;
  assign new_n29358 = new_n29357 ^ new_n29307;
  assign new_n29359 = new_n29227 ^ new_n28847;
  assign new_n29360 = new_n29359 ^ new_n29315;
  assign new_n29361 = new_n29360 ^ new_n29358;
  assign new_n29362 = new_n29361 ^ new_n29155;
  assign new_n29363 = new_n29362 ^ new_n29356;
  assign new_n29364 = new_n29363 ^ new_n29353;
  assign new_n29365 = ~new_n29364 & new_n29331;
  assign new_n29366 = new_n29365 ^ new_n29331;
  assign new_n29367 = new_n29364 ^ new_n29331;
  assign new_n29368 = new_n29367 ^ new_n29300;
  assign new_n29369 = new_n29263 ^ new_n29179;
  assign new_n29370 = new_n28499 ^ new_n24884;
  assign new_n29371 = new_n29370 ^ new_n13685;
  assign new_n29372 = new_n29305 ^ new_n28691;
  assign new_n29373 = new_n29206 ^ new_n28689;
  assign new_n29374 = new_n29373 ^ new_n28723;
  assign new_n29375 = new_n29374 ^ new_n29372;
  assign new_n29376 = new_n29313 ^ new_n28835;
  assign new_n29377 = new_n29224 ^ new_n28833;
  assign new_n29378 = new_n29377 ^ new_n28867;
  assign new_n29379 = new_n29378 ^ new_n29376;
  assign new_n29380 = new_n29379 ^ new_n29375;
  assign new_n29381 = new_n29380 ^ new_n29371;
  assign new_n29382 = new_n29381 ^ new_n29155;
  assign new_n29383 = ~new_n29066 & ~new_n29160;
  assign new_n29384 = new_n29383 ^ new_n29153;
  assign new_n29385 = new_n29384 ^ new_n29339;
  assign new_n29386 = new_n29296 ^ new_n29176;
  assign new_n29387 = new_n29386 ^ new_n29385;
  assign new_n29388 = new_n29387 ^ new_n29382;
  assign new_n29389 = new_n29388 ^ new_n29331;
  assign new_n29390 = new_n29389 ^ new_n29369;
  assign new_n29391 = new_n29390 ^ new_n29363;
  assign new_n29392 = ~new_n29368 & new_n29391;
  assign new_n29393 = new_n29392 ^ new_n29366;
  assign new_n29394 = new_n29331 ^ new_n29179;
  assign new_n29395 = new_n29394 ^ new_n29300;
  assign new_n29396 = ~new_n29390 & ~new_n29395;
  assign new_n29397 = new_n29396 ^ new_n29352;
  assign new_n29398 = ~new_n29363 & new_n29353;
  assign new_n29399 = new_n29179 & new_n29363;
  assign new_n29400 = new_n29399 ^ new_n29398;
  assign new_n29401 = new_n29400 ^ new_n29397;
  assign new_n29402 = new_n29263 ^ new_n29241;
  assign new_n29403 = new_n29390 ^ new_n29353;
  assign new_n29404 = new_n29300 & new_n29403;
  assign new_n29405 = new_n29299 ^ new_n29179;
  assign new_n29406 = ~new_n29301 & ~new_n29405;
  assign new_n29407 = new_n29406 ^ new_n29404;
  assign new_n29408 = new_n29400 ^ new_n29179;
  assign new_n29409 = new_n29408 ^ new_n29392;
  assign new_n29410 = new_n29409 ^ new_n29407;
  assign new_n29411 = new_n29410 ^ new_n29402;
  assign new_n29412 = new_n29389 ^ new_n29299;
  assign new_n29413 = new_n29412 ^ new_n29352;
  assign new_n29414 = ~new_n29369 & ~new_n29413;
  assign new_n29415 = new_n29414 ^ new_n29404;
  assign new_n29416 = new_n29412 ^ new_n29241;
  assign new_n29417 = new_n29416 ^ new_n29415;
  assign new_n29418 = new_n29364 ^ new_n29263;
  assign new_n29419 = new_n29413 ^ new_n29363;
  assign new_n29420 = ~new_n29418 & new_n29419;
  assign new_n29421 = new_n29331 ^ new_n29263;
  assign new_n29422 = new_n29416 & new_n29421;
  assign new_n29423 = new_n29422 ^ new_n29420;
  assign new_n29424 = new_n29423 ^ new_n29263;
  assign new_n29425 = new_n29424 ^ new_n29417;
  assign new_n29426 = new_n29422 ^ new_n29366;
  assign new_n29427 = new_n29426 ^ new_n29300;
  assign new_n29428 = new_n29414 ^ new_n29406;
  assign new_n29429 = new_n29388 ^ new_n29241;
  assign new_n29430 = new_n29429 ^ new_n29428;
  assign new_n29431 = new_n29430 ^ new_n29427;
  assign new_n29432 = new_n29397 ^ new_n29390;
  assign new_n29433 = new_n29392 ^ new_n29299;
  assign new_n29434 = new_n29433 ^ new_n29428;
  assign new_n29435 = new_n29434 ^ new_n29432;
  assign new_n29436 = new_n29431 & new_n29435;
  assign new_n29437 = new_n29436 ^ new_n29425;
  assign new_n29438 = ~new_n29437 & new_n29411;
  assign new_n29439 = new_n29438 ^ new_n29401;
  assign new_n29440 = new_n29439 ^ new_n29417;
  assign new_n29441 = new_n29436 ^ new_n29401;
  assign new_n29442 = new_n29441 ^ new_n29417;
  assign new_n29443 = new_n29420 ^ new_n29365;
  assign new_n29444 = new_n29443 ^ new_n29407;
  assign new_n29445 = ~new_n29444 & new_n29442;
  assign new_n29446 = new_n29445 ^ new_n29436;
  assign new_n29447 = ~new_n29425 & new_n29446;
  assign new_n29448 = new_n29447 ^ new_n29437;
  assign new_n29449 = ~new_n29448 & new_n29440;
  assign new_n29450 = new_n29449 ^ new_n29447;
  assign new_n29451 = new_n29450 ^ new_n29393;
  assign new_n29452 = new_n29451 ^ new_n29332;
  assign new_n29453 = new_n29452 ^ new_n29179;
  assign new_n29454 = new_n29438 ^ new_n29422;
  assign new_n29455 = new_n29454 ^ new_n29397;
  assign new_n29456 = new_n29455 ^ new_n29453;
  assign new_n29457 = ~new_n29301 & new_n29456;
  assign new_n29458 = new_n29445 ^ new_n29438;
  assign new_n29459 = new_n29424 ^ new_n29401;
  assign new_n29460 = new_n29459 ^ new_n29458;
  assign new_n29461 = ~new_n29413 & ~new_n29460;
  assign new_n29462 = new_n29461 ^ new_n29457;
  assign new_n29463 = new_n29447 ^ new_n29445;
  assign new_n29464 = new_n29463 ^ new_n29444;
  assign new_n29465 = ~new_n29464 & new_n29391;
  assign new_n29466 = new_n29447 ^ new_n29431;
  assign new_n29467 = ~new_n29390 & new_n29466;
  assign new_n29468 = new_n29467 ^ new_n29465;
  assign new_n29469 = ~new_n29395 & new_n29466;
  assign new_n29470 = new_n29469 ^ new_n29468;
  assign new_n29471 = ~new_n29368 & ~new_n29464;
  assign new_n29472 = ~new_n29369 & ~new_n29460;
  assign new_n29473 = ~new_n29405 & new_n29456;
  assign new_n29474 = new_n29473 ^ new_n29472;
  assign new_n29475 = new_n29474 ^ new_n29471;
  assign new_n29476 = new_n29475 ^ new_n29470;
  assign new_n29477 = new_n29476 ^ new_n29462;
  assign new_n29478 = new_n29477 ^ new_n28592;
  assign new_n29479 = new_n29472 ^ new_n29461;
  assign new_n29480 = new_n29445 ^ new_n29263;
  assign new_n29481 = new_n29420 ^ new_n29408;
  assign new_n29482 = new_n29481 ^ new_n29452;
  assign new_n29483 = new_n29482 ^ new_n29480;
  assign new_n29484 = ~new_n29483 & new_n29300;
  assign new_n29485 = ~new_n29418 & new_n29440;
  assign new_n29486 = ~new_n29483 & new_n29403;
  assign new_n29487 = new_n29486 ^ new_n29485;
  assign new_n29488 = new_n29445 ^ new_n29425;
  assign new_n29489 = ~new_n29363 & ~new_n29488;
  assign new_n29490 = new_n29489 ^ new_n29467;
  assign new_n29491 = new_n29449 ^ new_n29438;
  assign new_n29492 = new_n29491 ^ new_n29435;
  assign new_n29493 = new_n29421 & new_n29492;
  assign new_n29494 = new_n29493 ^ new_n29490;
  assign new_n29495 = new_n29494 ^ new_n29487;
  assign new_n29496 = new_n29495 ^ new_n29484;
  assign new_n29497 = new_n29496 ^ new_n29479;
  assign new_n29498 = new_n29497 ^ new_n29478;
  assign new_n29499 = new_n29498 ^ new_n28328;
  assign new_n29500 = new_n26201 ^ new_n26197;
  assign new_n29501 = new_n26192 ^ new_n26123;
  assign new_n29502 = new_n26165 ^ new_n26106;
  assign new_n29503 = new_n29502 ^ new_n26137;
  assign new_n29504 = new_n29503 ^ new_n29501;
  assign new_n29505 = ~new_n26126 & ~new_n29504;
  assign new_n29506 = new_n26188 ^ new_n26164;
  assign new_n29507 = ~new_n26086 & ~new_n29506;
  assign new_n29508 = new_n29507 ^ new_n29505;
  assign new_n29509 = ~new_n26152 & ~new_n26184;
  assign new_n29510 = ~new_n29506 & new_n26140;
  assign new_n29511 = new_n29510 ^ new_n29509;
  assign new_n29512 = ~new_n29504 & new_n26124;
  assign new_n29513 = new_n29512 ^ new_n26177;
  assign new_n29514 = new_n29513 ^ new_n29511;
  assign new_n29515 = new_n29514 ^ new_n29508;
  assign new_n29516 = new_n29515 ^ new_n29500;
  assign new_n29517 = new_n27223 ^ new_n27203;
  assign new_n29518 = new_n27140 ^ new_n26923;
  assign new_n29519 = ~new_n29518 & new_n29517;
  assign new_n29520 = new_n27227 ^ new_n27216;
  assign new_n29521 = new_n29520 ^ new_n27213;
  assign new_n29522 = new_n27195 & new_n29521;
  assign new_n29523 = new_n27227 ^ new_n27190;
  assign new_n29524 = ~new_n27140 & ~new_n29523;
  assign new_n29525 = new_n29524 ^ new_n27253;
  assign new_n29526 = new_n29525 ^ new_n29522;
  assign new_n29527 = new_n29526 ^ new_n27235;
  assign new_n29528 = new_n29527 ^ new_n29519;
  assign new_n29529 = ~new_n27139 & new_n29517;
  assign new_n29530 = new_n29529 ^ new_n27245;
  assign new_n29531 = ~new_n27173 & new_n29521;
  assign new_n29532 = new_n29531 ^ new_n29530;
  assign new_n29533 = ~new_n27198 & ~new_n27218;
  assign new_n29534 = new_n27223 ^ new_n27065;
  assign new_n29535 = new_n27200 ^ new_n27187;
  assign new_n29536 = new_n29535 ^ new_n27230;
  assign new_n29537 = new_n29536 ^ new_n29534;
  assign new_n29538 = ~new_n27183 & new_n29537;
  assign new_n29539 = new_n29538 ^ new_n29533;
  assign new_n29540 = new_n29539 ^ new_n29532;
  assign new_n29541 = new_n29540 ^ new_n29528;
  assign new_n29542 = new_n28294 ^ new_n28274;
  assign new_n29543 = new_n28209 ^ new_n27986;
  assign new_n29544 = ~new_n29543 & new_n29542;
  assign new_n29545 = new_n28298 ^ new_n28287;
  assign new_n29546 = new_n29545 ^ new_n28284;
  assign new_n29547 = new_n28265 & new_n29546;
  assign new_n29548 = new_n28298 ^ new_n28260;
  assign new_n29549 = ~new_n28209 & ~new_n29548;
  assign new_n29550 = new_n29549 ^ new_n28324;
  assign new_n29551 = new_n29550 ^ new_n29547;
  assign new_n29552 = new_n29551 ^ new_n28306;
  assign new_n29553 = new_n29552 ^ new_n29544;
  assign new_n29554 = ~new_n28208 & new_n29542;
  assign new_n29555 = new_n29554 ^ new_n28316;
  assign new_n29556 = ~new_n28267 & new_n29546;
  assign new_n29557 = new_n29556 ^ new_n29555;
  assign new_n29558 = ~new_n28269 & ~new_n28289;
  assign new_n29559 = new_n28294 ^ new_n28131;
  assign new_n29560 = new_n28271 ^ new_n28257;
  assign new_n29561 = new_n29560 ^ new_n28301;
  assign new_n29562 = new_n29561 ^ new_n29559;
  assign new_n29563 = ~new_n28252 & new_n29562;
  assign new_n29564 = new_n29563 ^ new_n29558;
  assign new_n29565 = new_n29564 ^ new_n29557;
  assign new_n29566 = new_n29565 ^ new_n29553;
  assign new_n29567 = new_n29566 ^ new_n29541;
  assign new_n29568 = new_n29567 ^ new_n29516;
  assign new_n29569 = new_n28558 ^ new_n28537;
  assign new_n29570 = new_n28490 ^ new_n28440;
  assign new_n29571 = new_n29569 & new_n29570;
  assign new_n29572 = new_n28562 ^ new_n28551;
  assign new_n29573 = new_n29572 ^ new_n28548;
  assign new_n29574 = ~new_n28528 & new_n29573;
  assign new_n29575 = new_n28562 ^ new_n28523;
  assign new_n29576 = ~new_n29575 & new_n28490;
  assign new_n29577 = new_n29576 ^ new_n28588;
  assign new_n29578 = new_n29577 ^ new_n29574;
  assign new_n29579 = new_n29578 ^ new_n28570;
  assign new_n29580 = new_n29579 ^ new_n29571;
  assign new_n29581 = new_n28489 & new_n29569;
  assign new_n29582 = new_n29581 ^ new_n28580;
  assign new_n29583 = ~new_n28530 & new_n29573;
  assign new_n29584 = new_n29583 ^ new_n29582;
  assign new_n29585 = ~new_n28532 & ~new_n28553;
  assign new_n29586 = new_n28558 ^ new_n28469;
  assign new_n29587 = new_n28534 ^ new_n28520;
  assign new_n29588 = new_n29587 ^ new_n28565;
  assign new_n29589 = new_n29588 ^ new_n29586;
  assign new_n29590 = new_n28515 & new_n29589;
  assign new_n29591 = new_n29590 ^ new_n29585;
  assign new_n29592 = new_n29591 ^ new_n29584;
  assign new_n29593 = new_n29592 ^ new_n29580;
  assign new_n29594 = new_n29593 ^ new_n25010;
  assign new_n29595 = new_n29594 ^ new_n20067;
  assign new_n29596 = new_n29364 ^ new_n29179;
  assign new_n29597 = ~new_n29488 & new_n29596;
  assign new_n29598 = new_n29449 ^ new_n29411;
  assign new_n29599 = new_n29364 & new_n29598;
  assign new_n29600 = new_n29599 ^ new_n29475;
  assign new_n29601 = new_n29416 & new_n29492;
  assign new_n29602 = new_n29601 ^ new_n29600;
  assign new_n29603 = new_n29602 ^ new_n29457;
  assign new_n29604 = new_n29603 ^ new_n29597;
  assign new_n29605 = new_n29604 ^ new_n29495;
  assign new_n29606 = new_n29605 ^ new_n29595;
  assign new_n29607 = new_n29493 ^ new_n29486;
  assign new_n29608 = new_n29419 & new_n29440;
  assign new_n29609 = ~new_n29367 & new_n29598;
  assign new_n29610 = new_n29609 ^ new_n29608;
  assign new_n29611 = new_n29610 ^ new_n29474;
  assign new_n29612 = new_n29599 ^ new_n29457;
  assign new_n29613 = new_n29612 ^ new_n29611;
  assign new_n29614 = new_n29613 ^ new_n29607;
  assign new_n29615 = new_n29614 ^ new_n29606;
  assign new_n29616 = new_n29615 ^ new_n29568;
  assign new_n29617 = ~new_n26159 & new_n26202;
  assign new_n29618 = new_n26189 ^ new_n26172;
  assign new_n29619 = new_n29618 ^ new_n26171;
  assign new_n29620 = ~new_n29619 & new_n26141;
  assign new_n29621 = new_n29620 ^ new_n29513;
  assign new_n29622 = new_n29621 ^ new_n29507;
  assign new_n29623 = new_n26089 & new_n26200;
  assign new_n29624 = new_n29623 ^ new_n29622;
  assign new_n29625 = new_n29624 ^ new_n29505;
  assign new_n29626 = new_n29625 ^ new_n29617;
  assign new_n29627 = new_n29626 ^ new_n26208;
  assign new_n29628 = new_n29608 ^ new_n29469;
  assign new_n29629 = new_n29489 ^ new_n29465;
  assign new_n29630 = new_n29629 ^ new_n29600;
  assign new_n29631 = new_n29630 ^ new_n29628;
  assign new_n29632 = new_n29631 ^ new_n29627;
  assign new_n29633 = new_n29632 ^ new_n29605;
  assign new_n29634 = ~new_n27199 & ~new_n27218;
  assign new_n29635 = new_n29634 ^ new_n27247;
  assign new_n29636 = new_n29529 ^ new_n27243;
  assign new_n29637 = new_n29636 ^ new_n29525;
  assign new_n29638 = new_n29637 ^ new_n29635;
  assign new_n29639 = ~new_n28270 & ~new_n28289;
  assign new_n29640 = new_n29639 ^ new_n28318;
  assign new_n29641 = new_n29554 ^ new_n28314;
  assign new_n29642 = new_n29641 ^ new_n29550;
  assign new_n29643 = new_n29642 ^ new_n29640;
  assign new_n29644 = new_n29643 ^ new_n29638;
  assign new_n29645 = ~new_n28533 & ~new_n28553;
  assign new_n29646 = new_n29645 ^ new_n28582;
  assign new_n29647 = new_n29581 ^ new_n28578;
  assign new_n29648 = new_n29647 ^ new_n29577;
  assign new_n29649 = new_n29648 ^ new_n29646;
  assign new_n29650 = new_n29649 ^ new_n26006;
  assign new_n29651 = new_n29650 ^ new_n20035;
  assign new_n29652 = new_n29469 ^ new_n29461;
  assign new_n29653 = new_n29652 ^ new_n29603;
  assign new_n29654 = ~new_n26135 & ~new_n26204;
  assign new_n29655 = new_n29654 ^ new_n26176;
  assign new_n29656 = new_n29655 ^ new_n29625;
  assign new_n29657 = new_n29656 ^ new_n29653;
  assign new_n29658 = new_n29657 ^ new_n29651;
  assign new_n29659 = new_n29658 ^ new_n29644;
  assign new_n29660 = new_n29659 ^ new_n29633;
  assign new_n29661 = new_n29623 ^ new_n26207;
  assign new_n29662 = new_n29661 ^ new_n29514;
  assign new_n29663 = new_n29662 ^ new_n29657;
  assign new_n29664 = new_n29538 ^ new_n29531;
  assign new_n29665 = ~new_n29523 & new_n27143;
  assign new_n29666 = new_n29665 ^ new_n29634;
  assign new_n29667 = new_n29666 ^ new_n27252;
  assign new_n29668 = new_n29524 ^ new_n27235;
  assign new_n29669 = new_n29668 ^ new_n29667;
  assign new_n29670 = new_n29669 ^ new_n29664;
  assign new_n29671 = new_n29563 ^ new_n29556;
  assign new_n29672 = ~new_n29548 & new_n28212;
  assign new_n29673 = new_n29672 ^ new_n29639;
  assign new_n29674 = new_n29673 ^ new_n28323;
  assign new_n29675 = new_n29549 ^ new_n28306;
  assign new_n29676 = new_n29675 ^ new_n29674;
  assign new_n29677 = new_n29676 ^ new_n29671;
  assign new_n29678 = new_n29677 ^ new_n29670;
  assign new_n29679 = new_n29678 ^ new_n29663;
  assign new_n29680 = new_n29601 ^ new_n29494;
  assign new_n29681 = new_n29680 ^ new_n29611;
  assign new_n29682 = new_n29590 ^ new_n29583;
  assign new_n29683 = ~new_n29575 & new_n28493;
  assign new_n29684 = new_n29683 ^ new_n29645;
  assign new_n29685 = new_n29684 ^ new_n28587;
  assign new_n29686 = new_n29576 ^ new_n28570;
  assign new_n29687 = new_n29686 ^ new_n29685;
  assign new_n29688 = new_n29687 ^ new_n29682;
  assign new_n29689 = new_n29688 ^ new_n25968;
  assign new_n29690 = new_n29689 ^ new_n20028;
  assign new_n29691 = new_n29690 ^ new_n29614;
  assign new_n29692 = new_n29691 ^ new_n29681;
  assign new_n29693 = new_n29692 ^ new_n29679;
  assign new_n29694 = new_n29693 ^ new_n29660;
  assign new_n29695 = new_n29694 ^ new_n29616;
  assign new_n29696 = new_n29695 ^ new_n29499;
  assign new_n29697 = new_n29584 ^ new_n29574;
  assign new_n29698 = new_n29697 ^ new_n29685;
  assign new_n29699 = new_n29698 ^ new_n26076;
  assign new_n29700 = new_n29699 ^ new_n20057;
  assign new_n29701 = new_n29700 ^ new_n29681;
  assign new_n29702 = new_n29532 ^ new_n29522;
  assign new_n29703 = new_n29702 ^ new_n29667;
  assign new_n29704 = new_n29557 ^ new_n29547;
  assign new_n29705 = new_n29704 ^ new_n29674;
  assign new_n29706 = new_n29705 ^ new_n29703;
  assign new_n29707 = new_n29706 ^ new_n29657;
  assign new_n29708 = new_n29707 ^ new_n29701;
  assign new_n29709 = new_n29578 ^ new_n28583;
  assign new_n29710 = new_n29709 ^ new_n26110;
  assign new_n29711 = new_n29710 ^ new_n20047;
  assign new_n29712 = new_n29526 ^ new_n27248;
  assign new_n29713 = new_n29551 ^ new_n28319;
  assign new_n29714 = new_n29713 ^ new_n29712;
  assign new_n29715 = new_n29714 ^ new_n29711;
  assign new_n29716 = new_n29715 ^ new_n29657;
  assign new_n29717 = new_n29654 ^ new_n29509;
  assign new_n29718 = ~new_n29619 & new_n26139;
  assign new_n29719 = new_n29718 ^ new_n26203;
  assign new_n29720 = new_n29719 ^ new_n29622;
  assign new_n29721 = new_n29720 ^ new_n29717;
  assign new_n29722 = new_n29602 ^ new_n29470;
  assign new_n29723 = new_n29722 ^ new_n29721;
  assign new_n29724 = new_n29723 ^ new_n29631;
  assign new_n29725 = new_n29724 ^ new_n29716;
  assign new_n29726 = new_n27251 ^ new_n27239;
  assign new_n29727 = new_n27066 & new_n29537;
  assign new_n29728 = new_n29727 ^ new_n29540;
  assign new_n29729 = new_n29728 ^ new_n29726;
  assign new_n29730 = new_n28322 ^ new_n28310;
  assign new_n29731 = new_n28132 & new_n29562;
  assign new_n29732 = new_n29731 ^ new_n29565;
  assign new_n29733 = new_n29732 ^ new_n29730;
  assign new_n29734 = new_n29733 ^ new_n29729;
  assign new_n29735 = new_n29734 ^ new_n29497;
  assign new_n29736 = new_n28586 ^ new_n28574;
  assign new_n29737 = ~new_n28470 & new_n29589;
  assign new_n29738 = new_n29737 ^ new_n29592;
  assign new_n29739 = new_n29738 ^ new_n29736;
  assign new_n29740 = new_n29739 ^ new_n26064;
  assign new_n29741 = new_n29740 ^ new_n20020;
  assign new_n29742 = new_n29718 ^ new_n26205;
  assign new_n29743 = new_n29742 ^ new_n29654;
  assign new_n29744 = new_n29743 ^ new_n29624;
  assign new_n29745 = new_n29744 ^ new_n29722;
  assign new_n29746 = new_n29745 ^ new_n29741;
  assign new_n29747 = new_n29746 ^ new_n29735;
  assign new_n29748 = new_n29747 ^ new_n29499;
  assign new_n29749 = new_n29748 ^ new_n29708;
  assign new_n29750 = new_n29749 ^ new_n29725;
  assign new_n29751 = new_n29708 & new_n29750;
  assign new_n29752 = new_n29751 ^ new_n29725;
  assign new_n29753 = new_n29505 ^ new_n26176;
  assign new_n29754 = new_n29743 ^ new_n29621;
  assign new_n29755 = new_n29754 ^ new_n29753;
  assign new_n29756 = new_n27247 ^ new_n27239;
  assign new_n29757 = new_n29756 ^ new_n29527;
  assign new_n29758 = new_n28318 ^ new_n28310;
  assign new_n29759 = new_n29758 ^ new_n29552;
  assign new_n29760 = new_n29759 ^ new_n29757;
  assign new_n29761 = new_n29760 ^ new_n29755;
  assign new_n29762 = new_n28582 ^ new_n28574;
  assign new_n29763 = new_n29762 ^ new_n29579;
  assign new_n29764 = new_n29763 ^ new_n26100;
  assign new_n29765 = new_n29764 ^ new_n20042;
  assign new_n29766 = new_n29765 ^ new_n29653;
  assign new_n29767 = new_n29766 ^ new_n29477;
  assign new_n29768 = new_n29767 ^ new_n29761;
  assign new_n29769 = new_n29768 ^ new_n29725;
  assign new_n29770 = new_n29769 ^ new_n29694;
  assign new_n29771 = new_n29768 ^ new_n29693;
  assign new_n29772 = new_n29725 ^ new_n29616;
  assign new_n29773 = new_n29772 ^ new_n29771;
  assign new_n29774 = new_n29770 & new_n29773;
  assign new_n29775 = new_n29774 ^ new_n29499;
  assign new_n29776 = new_n29775 ^ new_n29752;
  assign new_n29777 = ~new_n29693 & ~new_n29749;
  assign new_n29778 = new_n29777 ^ new_n29693;
  assign new_n29779 = new_n29747 ^ new_n29695;
  assign new_n29780 = new_n29771 & new_n29779;
  assign new_n29781 = new_n29780 ^ new_n29778;
  assign new_n29782 = new_n29768 ^ new_n29616;
  assign new_n29783 = new_n29782 ^ new_n29781;
  assign new_n29784 = new_n29696 & new_n29769;
  assign new_n29785 = new_n29747 ^ new_n29725;
  assign new_n29786 = new_n29785 ^ new_n29782;
  assign new_n29787 = new_n29772 & new_n29786;
  assign new_n29788 = new_n29787 ^ new_n29784;
  assign new_n29789 = new_n29747 ^ new_n29660;
  assign new_n29790 = new_n29789 ^ new_n29788;
  assign new_n29791 = new_n29790 ^ new_n29783;
  assign new_n29792 = new_n29775 ^ new_n29770;
  assign new_n29793 = new_n29749 ^ new_n29693;
  assign new_n29794 = new_n29793 ^ new_n29782;
  assign new_n29795 = new_n29770 ^ new_n29708;
  assign new_n29796 = new_n29794 & new_n29795;
  assign new_n29797 = new_n29796 ^ new_n29784;
  assign new_n29798 = new_n29787 ^ new_n29616;
  assign new_n29799 = new_n29798 ^ new_n29797;
  assign new_n29800 = new_n29799 ^ new_n29792;
  assign new_n29801 = ~new_n29791 & new_n29800;
  assign new_n29802 = new_n29801 ^ new_n29776;
  assign new_n29803 = new_n29770 ^ new_n29748;
  assign new_n29804 = new_n29782 & new_n29803;
  assign new_n29805 = new_n29804 ^ new_n29784;
  assign new_n29806 = new_n29805 ^ new_n29779;
  assign new_n29807 = new_n29806 ^ new_n29802;
  assign new_n29808 = new_n29768 ^ new_n29749;
  assign new_n29809 = new_n29708 ^ new_n29696;
  assign new_n29810 = new_n29808 & new_n29809;
  assign new_n29811 = new_n29810 ^ new_n29777;
  assign new_n29812 = new_n29804 ^ new_n29787;
  assign new_n29813 = new_n29812 ^ new_n29811;
  assign new_n29814 = ~new_n29813 & new_n29807;
  assign new_n29815 = new_n29768 ^ new_n29747;
  assign new_n29816 = new_n29796 ^ new_n29751;
  assign new_n29817 = new_n29816 ^ new_n29812;
  assign new_n29818 = new_n29817 ^ new_n29815;
  assign new_n29819 = new_n29810 ^ new_n29780;
  assign new_n29820 = new_n29819 ^ new_n29768;
  assign new_n29821 = new_n29820 ^ new_n29806;
  assign new_n29822 = new_n29821 ^ new_n29801;
  assign new_n29823 = new_n29818 & new_n29822;
  assign new_n29824 = new_n29823 ^ new_n29814;
  assign new_n29825 = new_n29820 ^ new_n29776;
  assign new_n29826 = new_n29825 ^ new_n29824;
  assign new_n29827 = new_n29696 & new_n29826;
  assign new_n29828 = new_n29814 ^ new_n29801;
  assign new_n29829 = new_n29821 & new_n29828;
  assign new_n29830 = new_n29829 ^ new_n29791;
  assign new_n29831 = ~new_n29830 & new_n29773;
  assign new_n29832 = new_n29831 ^ new_n29827;
  assign new_n29833 = new_n29747 ^ new_n29693;
  assign new_n29834 = new_n29796 ^ new_n29778;
  assign new_n29835 = new_n29823 ^ new_n29776;
  assign new_n29836 = new_n29835 ^ new_n29806;
  assign new_n29837 = new_n29829 ^ new_n29822;
  assign new_n29838 = new_n29836 & new_n29837;
  assign new_n29839 = new_n29838 ^ new_n29829;
  assign new_n29840 = new_n29839 ^ new_n29834;
  assign new_n29841 = new_n29840 ^ new_n29833;
  assign new_n29842 = new_n29841 ^ new_n29725;
  assign new_n29843 = new_n29823 ^ new_n29780;
  assign new_n29844 = new_n29843 ^ new_n29775;
  assign new_n29845 = new_n29844 ^ new_n29842;
  assign new_n29846 = ~new_n29845 & new_n29786;
  assign new_n29847 = new_n29838 ^ new_n29818;
  assign new_n29848 = new_n29749 & new_n29847;
  assign new_n29849 = new_n29829 ^ new_n29814;
  assign new_n29850 = new_n29849 ^ new_n29813;
  assign new_n29851 = ~new_n29850 & new_n29794;
  assign new_n29852 = ~new_n29845 & new_n29772;
  assign new_n29853 = new_n29769 & new_n29826;
  assign new_n29854 = new_n29853 ^ new_n29852;
  assign new_n29855 = new_n29854 ^ new_n29851;
  assign new_n29856 = new_n29855 ^ new_n29848;
  assign new_n29857 = new_n29838 ^ new_n29823;
  assign new_n29858 = new_n29857 ^ new_n29800;
  assign new_n29859 = new_n29779 & new_n29858;
  assign new_n29860 = new_n29859 ^ new_n29856;
  assign new_n29861 = new_n29860 ^ new_n29846;
  assign new_n29862 = new_n29861 ^ new_n29832;
  assign new_n29863 = new_n26960 ^ new_n26605;
  assign new_n29864 = new_n27052 ^ new_n27037;
  assign new_n29865 = new_n29864 ^ new_n29863;
  assign new_n29866 = new_n27099 ^ new_n26960;
  assign new_n29867 = new_n27112 ^ new_n26960;
  assign new_n29868 = new_n29867 ^ new_n27131;
  assign new_n29869 = ~new_n27099 & ~new_n29868;
  assign new_n29870 = new_n29869 ^ new_n27099;
  assign new_n29871 = new_n29868 ^ new_n27099;
  assign new_n29872 = new_n29871 ^ new_n29864;
  assign new_n29873 = new_n27052 ^ new_n26605;
  assign new_n29874 = new_n27164 ^ new_n27099;
  assign new_n29875 = new_n29874 ^ new_n29873;
  assign new_n29876 = new_n29875 ^ new_n27131;
  assign new_n29877 = new_n29872 & new_n29876;
  assign new_n29878 = new_n29877 ^ new_n29870;
  assign new_n29879 = new_n27099 ^ new_n26605;
  assign new_n29880 = new_n29879 ^ new_n29864;
  assign new_n29881 = new_n29875 & new_n29880;
  assign new_n29882 = new_n29881 ^ new_n27112;
  assign new_n29883 = ~new_n29867 & new_n27131;
  assign new_n29884 = ~new_n27131 & new_n26605;
  assign new_n29885 = new_n29884 ^ new_n29883;
  assign new_n29886 = new_n29885 ^ new_n29882;
  assign new_n29887 = new_n27052 ^ new_n26960;
  assign new_n29888 = new_n29875 ^ new_n29867;
  assign new_n29889 = new_n29864 & new_n29888;
  assign new_n29890 = new_n27037 ^ new_n26605;
  assign new_n29891 = new_n29865 & new_n29890;
  assign new_n29892 = new_n29891 ^ new_n29889;
  assign new_n29893 = new_n29885 ^ new_n26605;
  assign new_n29894 = new_n29893 ^ new_n29877;
  assign new_n29895 = new_n29894 ^ new_n29892;
  assign new_n29896 = new_n29895 ^ new_n29887;
  assign new_n29897 = new_n29874 ^ new_n27037;
  assign new_n29898 = new_n29897 ^ new_n27112;
  assign new_n29899 = new_n29873 & new_n29898;
  assign new_n29900 = new_n29899 ^ new_n29889;
  assign new_n29901 = new_n29897 ^ new_n26960;
  assign new_n29902 = new_n29901 ^ new_n29900;
  assign new_n29903 = new_n27099 ^ new_n27052;
  assign new_n29904 = new_n29901 & new_n29903;
  assign new_n29905 = new_n29868 ^ new_n27052;
  assign new_n29906 = new_n29898 ^ new_n27131;
  assign new_n29907 = new_n29905 & new_n29906;
  assign new_n29908 = new_n29907 ^ new_n29904;
  assign new_n29909 = new_n29908 ^ new_n27052;
  assign new_n29910 = new_n29909 ^ new_n29902;
  assign new_n29911 = new_n29904 ^ new_n29870;
  assign new_n29912 = new_n29911 ^ new_n29864;
  assign new_n29913 = new_n29899 ^ new_n29891;
  assign new_n29914 = new_n27164 ^ new_n26960;
  assign new_n29915 = new_n29914 ^ new_n29913;
  assign new_n29916 = new_n29915 ^ new_n29912;
  assign new_n29917 = new_n29882 ^ new_n29875;
  assign new_n29918 = new_n29899 ^ new_n29877;
  assign new_n29919 = new_n29891 ^ new_n27037;
  assign new_n29920 = new_n29919 ^ new_n29918;
  assign new_n29921 = new_n29920 ^ new_n29917;
  assign new_n29922 = ~new_n29916 & new_n29921;
  assign new_n29923 = new_n29922 ^ new_n29910;
  assign new_n29924 = new_n29896 & new_n29923;
  assign new_n29925 = new_n29924 ^ new_n29886;
  assign new_n29926 = new_n29925 ^ new_n29902;
  assign new_n29927 = new_n29922 ^ new_n29886;
  assign new_n29928 = new_n29927 ^ new_n29902;
  assign new_n29929 = new_n29907 ^ new_n29869;
  assign new_n29930 = new_n29929 ^ new_n29892;
  assign new_n29931 = ~new_n29930 & new_n29928;
  assign new_n29932 = new_n29931 ^ new_n29922;
  assign new_n29933 = new_n29910 & new_n29932;
  assign new_n29934 = new_n29933 ^ new_n29923;
  assign new_n29935 = new_n29926 & new_n29934;
  assign new_n29936 = new_n29935 ^ new_n29933;
  assign new_n29937 = new_n29936 ^ new_n29878;
  assign new_n29938 = new_n29937 ^ new_n29866;
  assign new_n29939 = new_n29938 ^ new_n26605;
  assign new_n29940 = new_n29924 ^ new_n29904;
  assign new_n29941 = new_n29940 ^ new_n29882;
  assign new_n29942 = new_n29941 ^ new_n29939;
  assign new_n29943 = ~new_n29942 & new_n29865;
  assign new_n29944 = new_n29931 ^ new_n29924;
  assign new_n29945 = new_n29909 ^ new_n29886;
  assign new_n29946 = new_n29945 ^ new_n29944;
  assign new_n29947 = new_n29898 & new_n29946;
  assign new_n29948 = new_n29947 ^ new_n29943;
  assign new_n29949 = new_n29933 ^ new_n29931;
  assign new_n29950 = new_n29949 ^ new_n29930;
  assign new_n29951 = ~new_n29950 & new_n29876;
  assign new_n29952 = new_n29933 ^ new_n29916;
  assign new_n29953 = ~new_n29952 & new_n29875;
  assign new_n29954 = new_n29953 ^ new_n29951;
  assign new_n29955 = ~new_n29952 & new_n29880;
  assign new_n29956 = new_n29955 ^ new_n29954;
  assign new_n29957 = ~new_n29950 & new_n29872;
  assign new_n29958 = ~new_n29942 & new_n29890;
  assign new_n29959 = new_n29873 & new_n29946;
  assign new_n29960 = new_n29959 ^ new_n29958;
  assign new_n29961 = new_n29960 ^ new_n29957;
  assign new_n29962 = new_n29961 ^ new_n29956;
  assign new_n29963 = new_n29962 ^ new_n29948;
  assign new_n29964 = new_n29963 ^ new_n20167;
  assign new_n29965 = new_n29931 ^ new_n29910;
  assign new_n29966 = new_n29868 ^ new_n26605;
  assign new_n29967 = new_n29965 & new_n29966;
  assign new_n29968 = new_n29935 ^ new_n29924;
  assign new_n29969 = new_n29968 ^ new_n29921;
  assign new_n29970 = new_n29901 & new_n29969;
  assign new_n29971 = new_n29935 ^ new_n29896;
  assign new_n29972 = new_n29868 & new_n29971;
  assign new_n29973 = new_n29972 ^ new_n29961;
  assign new_n29974 = new_n29973 ^ new_n29970;
  assign new_n29975 = new_n29974 ^ new_n29943;
  assign new_n29976 = new_n29975 ^ new_n29967;
  assign new_n29977 = new_n27131 & new_n29965;
  assign new_n29978 = new_n29977 ^ new_n29953;
  assign new_n29979 = new_n29903 & new_n29969;
  assign new_n29980 = new_n29979 ^ new_n29978;
  assign new_n29981 = new_n29905 & new_n29926;
  assign new_n29982 = new_n29931 ^ new_n27052;
  assign new_n29983 = new_n29907 ^ new_n29893;
  assign new_n29984 = new_n29983 ^ new_n29938;
  assign new_n29985 = new_n29984 ^ new_n29982;
  assign new_n29986 = ~new_n29985 & new_n29888;
  assign new_n29987 = new_n29986 ^ new_n29981;
  assign new_n29988 = new_n29987 ^ new_n29980;
  assign new_n29989 = new_n29988 ^ new_n29976;
  assign new_n29990 = new_n29989 ^ new_n20206;
  assign new_n29991 = new_n29906 & new_n29926;
  assign new_n29992 = new_n29991 ^ new_n29955;
  assign new_n29993 = new_n29977 ^ new_n29951;
  assign new_n29994 = new_n29993 ^ new_n29973;
  assign new_n29995 = new_n29994 ^ new_n29992;
  assign new_n29996 = new_n29995 ^ new_n20197;
  assign new_n29997 = new_n29986 ^ new_n29979;
  assign new_n29998 = new_n29871 & new_n29971;
  assign new_n29999 = new_n29998 ^ new_n29991;
  assign new_n30000 = new_n29999 ^ new_n29960;
  assign new_n30001 = new_n29972 ^ new_n29943;
  assign new_n30002 = new_n30001 ^ new_n30000;
  assign new_n30003 = new_n30002 ^ new_n29997;
  assign new_n30004 = new_n30003 ^ new_n20191;
  assign new_n30005 = new_n30004 ^ new_n29996;
  assign new_n30006 = new_n30005 ^ new_n29990;
  assign new_n30007 = new_n30006 ^ new_n29964;
  assign new_n30008 = new_n29980 ^ new_n29970;
  assign new_n30009 = new_n30008 ^ new_n30000;
  assign new_n30010 = new_n30009 ^ new_n20215;
  assign new_n30011 = new_n29974 ^ new_n29956;
  assign new_n30012 = new_n30011 ^ new_n20182;
  assign new_n30013 = new_n29959 ^ new_n29947;
  assign new_n30014 = ~new_n29985 & new_n29864;
  assign new_n30015 = new_n30014 ^ new_n29988;
  assign new_n30016 = new_n30015 ^ new_n30013;
  assign new_n30017 = new_n30016 ^ new_n20173;
  assign new_n30018 = new_n30017 ^ new_n29964;
  assign new_n30019 = new_n30018 ^ new_n30010;
  assign new_n30020 = new_n30019 ^ new_n30012;
  assign new_n30021 = ~new_n30010 & ~new_n30020;
  assign new_n30022 = new_n30021 ^ new_n30012;
  assign new_n30023 = new_n29955 ^ new_n29947;
  assign new_n30024 = new_n30023 ^ new_n29975;
  assign new_n30025 = new_n30024 ^ new_n20178;
  assign new_n30026 = new_n30025 ^ new_n30012;
  assign new_n30027 = new_n30026 ^ new_n30005;
  assign new_n30028 = new_n30012 ^ new_n30004;
  assign new_n30029 = new_n30025 ^ new_n29990;
  assign new_n30030 = new_n30029 ^ new_n30028;
  assign new_n30031 = ~new_n30027 & new_n30030;
  assign new_n30032 = new_n30031 ^ new_n29964;
  assign new_n30033 = new_n30032 ^ new_n30022;
  assign new_n30034 = ~new_n30004 & new_n30019;
  assign new_n30035 = new_n30034 ^ new_n30004;
  assign new_n30036 = new_n30017 ^ new_n30006;
  assign new_n30037 = new_n30025 ^ new_n30004;
  assign new_n30038 = new_n30036 & new_n30037;
  assign new_n30039 = new_n30038 ^ new_n30035;
  assign new_n30040 = new_n30039 ^ new_n30029;
  assign new_n30041 = new_n30007 & new_n30026;
  assign new_n30042 = new_n30017 ^ new_n30012;
  assign new_n30043 = new_n30042 ^ new_n30029;
  assign new_n30044 = new_n30012 ^ new_n29990;
  assign new_n30045 = ~new_n30043 & new_n30044;
  assign new_n30046 = new_n30045 ^ new_n30041;
  assign new_n30047 = new_n30017 ^ new_n29996;
  assign new_n30048 = new_n30047 ^ new_n30046;
  assign new_n30049 = new_n30048 ^ new_n30040;
  assign new_n30050 = new_n30032 ^ new_n30027;
  assign new_n30051 = new_n30019 ^ new_n30004;
  assign new_n30052 = new_n30051 ^ new_n30029;
  assign new_n30053 = new_n30027 ^ new_n30010;
  assign new_n30054 = ~new_n30052 & new_n30053;
  assign new_n30055 = new_n30054 ^ new_n29990;
  assign new_n30056 = new_n30055 ^ new_n30046;
  assign new_n30057 = new_n30056 ^ new_n30050;
  assign new_n30058 = ~new_n30049 & new_n30057;
  assign new_n30059 = new_n30058 ^ new_n30033;
  assign new_n30060 = new_n30027 ^ new_n30018;
  assign new_n30061 = ~new_n30060 & new_n30029;
  assign new_n30062 = new_n30061 ^ new_n30041;
  assign new_n30063 = new_n30062 ^ new_n30036;
  assign new_n30064 = new_n30063 ^ new_n30059;
  assign new_n30065 = new_n30025 ^ new_n30019;
  assign new_n30066 = new_n30010 ^ new_n30007;
  assign new_n30067 = ~new_n30065 & ~new_n30066;
  assign new_n30068 = new_n30067 ^ new_n30034;
  assign new_n30069 = new_n30061 ^ new_n30045;
  assign new_n30070 = new_n30069 ^ new_n30068;
  assign new_n30071 = ~new_n30064 & ~new_n30070;
  assign new_n30072 = new_n30025 ^ new_n30017;
  assign new_n30073 = new_n30054 ^ new_n30021;
  assign new_n30074 = new_n30073 ^ new_n30069;
  assign new_n30075 = new_n30074 ^ new_n30072;
  assign new_n30076 = new_n30067 ^ new_n30038;
  assign new_n30077 = new_n30076 ^ new_n30025;
  assign new_n30078 = new_n30077 ^ new_n30063;
  assign new_n30079 = new_n30078 ^ new_n30058;
  assign new_n30080 = ~new_n30075 & new_n30079;
  assign new_n30081 = new_n30080 ^ new_n30071;
  assign new_n30082 = new_n30077 ^ new_n30033;
  assign new_n30083 = new_n30082 ^ new_n30081;
  assign new_n30084 = ~new_n30083 & new_n30007;
  assign new_n30085 = new_n30071 ^ new_n30058;
  assign new_n30086 = new_n30078 & new_n30085;
  assign new_n30087 = new_n30086 ^ new_n30049;
  assign new_n30088 = ~new_n30087 & new_n30030;
  assign new_n30089 = new_n30088 ^ new_n30084;
  assign new_n30090 = new_n30017 ^ new_n30004;
  assign new_n30091 = new_n30054 ^ new_n30035;
  assign new_n30092 = new_n30080 ^ new_n30033;
  assign new_n30093 = new_n30092 ^ new_n30063;
  assign new_n30094 = new_n30086 ^ new_n30079;
  assign new_n30095 = ~new_n30093 & new_n30094;
  assign new_n30096 = new_n30095 ^ new_n30086;
  assign new_n30097 = new_n30096 ^ new_n30091;
  assign new_n30098 = new_n30097 ^ new_n30090;
  assign new_n30099 = new_n30098 ^ new_n30012;
  assign new_n30100 = new_n30080 ^ new_n30038;
  assign new_n30101 = new_n30100 ^ new_n30032;
  assign new_n30102 = new_n30101 ^ new_n30099;
  assign new_n30103 = ~new_n30043 & ~new_n30102;
  assign new_n30104 = new_n30095 ^ new_n30075;
  assign new_n30105 = ~new_n30019 & ~new_n30104;
  assign new_n30106 = new_n30086 ^ new_n30071;
  assign new_n30107 = new_n30106 ^ new_n30070;
  assign new_n30108 = ~new_n30052 & ~new_n30107;
  assign new_n30109 = ~new_n30102 & new_n30044;
  assign new_n30110 = ~new_n30083 & new_n30026;
  assign new_n30111 = new_n30110 ^ new_n30109;
  assign new_n30112 = new_n30111 ^ new_n30108;
  assign new_n30113 = new_n30112 ^ new_n30105;
  assign new_n30114 = new_n30095 ^ new_n30080;
  assign new_n30115 = new_n30114 ^ new_n30057;
  assign new_n30116 = new_n30036 & new_n30115;
  assign new_n30117 = new_n30116 ^ new_n30113;
  assign new_n30118 = new_n30117 ^ new_n30103;
  assign new_n30119 = new_n30118 ^ new_n30089;
  assign new_n30120 = new_n30119 ^ new_n20958;
  assign new_n30121 = new_n30120 ^ new_n29862;
  assign new_n30122 = new_n30103 ^ new_n30084;
  assign new_n30123 = ~new_n30027 & ~new_n30087;
  assign new_n30124 = ~new_n30107 & new_n30053;
  assign new_n30125 = new_n30124 ^ new_n30123;
  assign new_n30126 = new_n30125 ^ new_n30088;
  assign new_n30127 = new_n30126 ^ new_n30112;
  assign new_n30128 = new_n30127 ^ new_n30122;
  assign new_n30129 = new_n30128 ^ new_n20899;
  assign new_n30130 = new_n29846 ^ new_n29827;
  assign new_n30131 = ~new_n29830 & new_n29770;
  assign new_n30132 = ~new_n29850 & new_n29795;
  assign new_n30133 = new_n30132 ^ new_n30131;
  assign new_n30134 = new_n30133 ^ new_n29831;
  assign new_n30135 = new_n30134 ^ new_n29855;
  assign new_n30136 = new_n30135 ^ new_n30130;
  assign new_n30137 = new_n30136 ^ new_n30129;
  assign new_n30138 = new_n30110 ^ new_n30084;
  assign new_n30139 = new_n30071 ^ new_n30025;
  assign new_n30140 = new_n30067 ^ new_n30021;
  assign new_n30141 = new_n30140 ^ new_n30098;
  assign new_n30142 = new_n30141 ^ new_n30139;
  assign new_n30143 = new_n30029 & new_n30142;
  assign new_n30144 = new_n30037 & new_n30115;
  assign new_n30145 = new_n30078 ^ new_n30071;
  assign new_n30146 = ~new_n30010 & new_n30145;
  assign new_n30147 = new_n30146 ^ new_n30123;
  assign new_n30148 = new_n30147 ^ new_n30144;
  assign new_n30149 = ~new_n30060 & new_n30142;
  assign new_n30150 = ~new_n30065 & ~new_n30093;
  assign new_n30151 = new_n30150 ^ new_n30149;
  assign new_n30152 = new_n30151 ^ new_n30148;
  assign new_n30153 = new_n30152 ^ new_n30143;
  assign new_n30154 = new_n30153 ^ new_n30138;
  assign new_n30155 = new_n30154 ^ new_n20928;
  assign new_n30156 = new_n29853 ^ new_n29827;
  assign new_n30157 = new_n29814 ^ new_n29768;
  assign new_n30158 = new_n29810 ^ new_n29751;
  assign new_n30159 = new_n30158 ^ new_n29841;
  assign new_n30160 = new_n30159 ^ new_n30157;
  assign new_n30161 = ~new_n30160 & new_n29782;
  assign new_n30162 = new_n29771 & new_n29858;
  assign new_n30163 = new_n29821 ^ new_n29814;
  assign new_n30164 = new_n29708 & new_n30163;
  assign new_n30165 = new_n30164 ^ new_n30131;
  assign new_n30166 = new_n30165 ^ new_n30162;
  assign new_n30167 = ~new_n30160 & new_n29803;
  assign new_n30168 = new_n29808 & new_n29836;
  assign new_n30169 = new_n30168 ^ new_n30167;
  assign new_n30170 = new_n30169 ^ new_n30166;
  assign new_n30171 = new_n30170 ^ new_n30161;
  assign new_n30172 = new_n30171 ^ new_n30156;
  assign new_n30173 = new_n30172 ^ new_n30155;
  assign new_n30174 = new_n30134 ^ new_n29860;
  assign new_n30175 = new_n30126 ^ new_n30117;
  assign new_n30176 = new_n30175 ^ new_n20972;
  assign new_n30177 = new_n30176 ^ new_n30174;
  assign new_n30178 = new_n29809 & new_n29836;
  assign new_n30179 = new_n30178 ^ new_n29831;
  assign new_n30180 = new_n30164 ^ new_n30132;
  assign new_n30181 = new_n30180 ^ new_n29856;
  assign new_n30182 = new_n30181 ^ new_n30179;
  assign new_n30183 = ~new_n30066 & ~new_n30093;
  assign new_n30184 = new_n30183 ^ new_n30088;
  assign new_n30185 = new_n30146 ^ new_n30124;
  assign new_n30186 = new_n30185 ^ new_n30113;
  assign new_n30187 = new_n30186 ^ new_n30184;
  assign new_n30188 = new_n30187 ^ new_n20799;
  assign new_n30189 = new_n30188 ^ new_n30182;
  assign new_n30190 = new_n29750 & new_n30163;
  assign new_n30191 = new_n30190 ^ new_n29861;
  assign new_n30192 = new_n30191 ^ new_n30170;
  assign new_n30193 = ~new_n30020 & new_n30145;
  assign new_n30194 = new_n30193 ^ new_n30118;
  assign new_n30195 = new_n30194 ^ new_n30152;
  assign new_n30196 = new_n30195 ^ new_n20431;
  assign new_n30197 = new_n30196 ^ new_n30192;
  assign new_n30198 = new_n30149 ^ new_n30144;
  assign new_n30199 = ~new_n30051 & ~new_n30104;
  assign new_n30200 = new_n30199 ^ new_n30183;
  assign new_n30201 = new_n30200 ^ new_n30111;
  assign new_n30202 = new_n30105 ^ new_n30103;
  assign new_n30203 = new_n30202 ^ new_n30201;
  assign new_n30204 = new_n30203 ^ new_n30198;
  assign new_n30205 = new_n30204 ^ new_n20857;
  assign new_n30206 = new_n30167 ^ new_n30162;
  assign new_n30207 = new_n29793 & new_n29847;
  assign new_n30208 = new_n30207 ^ new_n30178;
  assign new_n30209 = new_n30208 ^ new_n29854;
  assign new_n30210 = new_n29848 ^ new_n29846;
  assign new_n30211 = new_n30210 ^ new_n30209;
  assign new_n30212 = new_n30211 ^ new_n30206;
  assign new_n30213 = new_n30212 ^ new_n30205;
  assign new_n30214 = new_n30148 ^ new_n30116;
  assign new_n30215 = new_n30214 ^ new_n30201;
  assign new_n30216 = new_n30215 ^ new_n20937;
  assign new_n30217 = new_n30166 ^ new_n29859;
  assign new_n30218 = new_n30217 ^ new_n30209;
  assign new_n30219 = new_n30218 ^ new_n30216;
  assign new_n30220 = new_n28100 ^ new_n17416;
  assign new_n30221 = new_n30220 ^ new_n27148;
  assign new_n30222 = new_n27080 ^ new_n27045;
  assign new_n30223 = new_n30222 ^ new_n27027;
  assign new_n30224 = new_n30223 ^ new_n30221;
  assign new_n30225 = new_n27089 ^ new_n27063;
  assign new_n30226 = new_n27134 ^ new_n27102;
  assign new_n30227 = new_n28158 ^ new_n17419;
  assign new_n30228 = new_n30227 ^ new_n27016;
  assign new_n30229 = new_n30228 ^ new_n30226;
  assign new_n30230 = new_n30229 ^ new_n30225;
  assign new_n30231 = new_n27031 ^ new_n27021;
  assign new_n30232 = new_n28222 ^ new_n17423;
  assign new_n30233 = new_n30232 ^ new_n26913;
  assign new_n30234 = new_n30233 ^ new_n30231;
  assign new_n30235 = new_n27159 ^ new_n27063;
  assign new_n30236 = new_n30235 ^ new_n30234;
  assign new_n30237 = new_n30236 ^ new_n30230;
  assign new_n30238 = new_n30237 ^ new_n30224;
  assign new_n30239 = new_n27124 ^ new_n27000;
  assign new_n30240 = new_n28178 ^ new_n17429;
  assign new_n30241 = new_n30240 ^ new_n27059;
  assign new_n30242 = new_n30241 ^ new_n27108;
  assign new_n30243 = new_n30242 ^ new_n30239;
  assign new_n30244 = new_n30243 ^ new_n30238;
  assign new_n30245 = new_n26984 ^ new_n26766;
  assign new_n30246 = new_n28022 ^ new_n17426;
  assign new_n30247 = new_n30246 ^ new_n27120;
  assign new_n30248 = new_n30247 ^ new_n26941;
  assign new_n30249 = new_n30248 ^ new_n30245;
  assign new_n30250 = new_n30249 ^ new_n30243;
  assign new_n30251 = new_n28200 ^ new_n17431;
  assign new_n30252 = new_n30251 ^ new_n27071;
  assign new_n30253 = new_n27137 ^ new_n27063;
  assign new_n30254 = new_n30253 ^ new_n30252;
  assign new_n30255 = new_n30254 ^ new_n30250;
  assign new_n30256 = new_n30230 & new_n30255;
  assign new_n30257 = new_n30256 ^ new_n30230;
  assign new_n30258 = new_n30249 ^ new_n30238;
  assign new_n30259 = new_n28116 ^ new_n17420;
  assign new_n30260 = new_n30259 ^ new_n27125;
  assign new_n30261 = new_n27062 ^ new_n27049;
  assign new_n30262 = new_n30261 ^ new_n26355;
  assign new_n30263 = new_n30262 ^ new_n30260;
  assign new_n30264 = new_n30263 ^ new_n30230;
  assign new_n30265 = ~new_n30264 & new_n30258;
  assign new_n30266 = new_n30265 ^ new_n30257;
  assign new_n30267 = new_n30263 ^ new_n30224;
  assign new_n30268 = new_n30267 ^ new_n30266;
  assign new_n30269 = new_n27154 ^ new_n26920;
  assign new_n30270 = new_n27966 ^ new_n17417;
  assign new_n30271 = new_n30270 ^ new_n30269;
  assign new_n30272 = new_n30271 ^ new_n27063;
  assign new_n30273 = new_n26905 ^ new_n26760;
  assign new_n30274 = new_n30273 ^ new_n26965;
  assign new_n30275 = new_n30274 ^ new_n30272;
  assign new_n30276 = new_n30275 ^ new_n30249;
  assign new_n30277 = new_n30276 ^ new_n30267;
  assign new_n30278 = new_n30275 ^ new_n30224;
  assign new_n30279 = ~new_n30277 & new_n30278;
  assign new_n30280 = new_n30275 ^ new_n30263;
  assign new_n30281 = new_n30244 & new_n30280;
  assign new_n30282 = new_n30281 ^ new_n30279;
  assign new_n30283 = new_n30249 ^ new_n30236;
  assign new_n30284 = new_n30283 ^ new_n30282;
  assign new_n30285 = new_n30284 ^ new_n30268;
  assign new_n30286 = new_n30280 ^ new_n30237;
  assign new_n30287 = new_n30275 ^ new_n30230;
  assign new_n30288 = new_n30287 ^ new_n30267;
  assign new_n30289 = ~new_n30286 & ~new_n30288;
  assign new_n30290 = new_n30289 ^ new_n30243;
  assign new_n30291 = new_n30290 ^ new_n30286;
  assign new_n30292 = new_n30286 ^ new_n30254;
  assign new_n30293 = new_n30255 ^ new_n30230;
  assign new_n30294 = new_n30293 ^ new_n30267;
  assign new_n30295 = new_n30292 & new_n30294;
  assign new_n30296 = new_n30295 ^ new_n30282;
  assign new_n30297 = new_n30296 ^ new_n30224;
  assign new_n30298 = new_n30297 ^ new_n30291;
  assign new_n30299 = ~new_n30285 & new_n30298;
  assign new_n30300 = new_n30286 ^ new_n30250;
  assign new_n30301 = ~new_n30300 & new_n30267;
  assign new_n30302 = new_n30301 ^ new_n30281;
  assign new_n30303 = new_n30302 ^ new_n30258;
  assign new_n30304 = new_n30263 ^ new_n30255;
  assign new_n30305 = new_n30254 ^ new_n30244;
  assign new_n30306 = ~new_n30304 & ~new_n30305;
  assign new_n30307 = new_n30306 ^ new_n30265;
  assign new_n30308 = new_n30307 ^ new_n30263;
  assign new_n30309 = new_n30308 ^ new_n30303;
  assign new_n30310 = new_n30309 ^ new_n30299;
  assign new_n30311 = new_n30263 ^ new_n30249;
  assign new_n30312 = new_n30275 ^ new_n30255;
  assign new_n30313 = ~new_n30254 & ~new_n30312;
  assign new_n30314 = new_n30313 ^ new_n30295;
  assign new_n30315 = new_n30301 ^ new_n30279;
  assign new_n30316 = new_n30315 ^ new_n30314;
  assign new_n30317 = new_n30316 ^ new_n30311;
  assign new_n30318 = ~new_n30317 & new_n30310;
  assign new_n30319 = new_n30313 ^ new_n30275;
  assign new_n30320 = new_n30319 ^ new_n30290;
  assign new_n30321 = new_n30320 ^ new_n30299;
  assign new_n30322 = new_n30321 ^ new_n30303;
  assign new_n30323 = new_n30306 ^ new_n30256;
  assign new_n30324 = new_n30323 ^ new_n30315;
  assign new_n30325 = ~new_n30322 & ~new_n30324;
  assign new_n30326 = new_n30325 ^ new_n30318;
  assign new_n30327 = new_n30320 ^ new_n30308;
  assign new_n30328 = new_n30327 ^ new_n30326;
  assign new_n30329 = ~new_n30328 & new_n30244;
  assign new_n30330 = ~new_n30328 & new_n30280;
  assign new_n30331 = new_n30330 ^ new_n30329;
  assign new_n30332 = new_n30325 ^ new_n30263;
  assign new_n30333 = new_n30313 ^ new_n30306;
  assign new_n30334 = new_n30249 ^ new_n30230;
  assign new_n30335 = new_n30295 ^ new_n30257;
  assign new_n30336 = new_n30320 ^ new_n30318;
  assign new_n30337 = new_n30336 ^ new_n30303;
  assign new_n30338 = new_n30325 ^ new_n30299;
  assign new_n30339 = ~new_n30338 & new_n30309;
  assign new_n30340 = new_n30339 ^ new_n30299;
  assign new_n30341 = ~new_n30337 & new_n30340;
  assign new_n30342 = new_n30339 ^ new_n30309;
  assign new_n30343 = new_n30342 ^ new_n30341;
  assign new_n30344 = new_n30343 ^ new_n30335;
  assign new_n30345 = new_n30344 ^ new_n30334;
  assign new_n30346 = new_n30345 ^ new_n30333;
  assign new_n30347 = new_n30346 ^ new_n30332;
  assign new_n30348 = new_n30267 & new_n30347;
  assign new_n30349 = ~new_n30304 & ~new_n30337;
  assign new_n30350 = ~new_n30300 & new_n30347;
  assign new_n30351 = new_n30350 ^ new_n30349;
  assign new_n30352 = new_n30341 ^ new_n30318;
  assign new_n30353 = new_n30352 ^ new_n30298;
  assign new_n30354 = ~new_n30264 & new_n30353;
  assign new_n30355 = new_n30325 ^ new_n30309;
  assign new_n30356 = ~new_n30254 & new_n30355;
  assign new_n30357 = new_n30342 ^ new_n30285;
  assign new_n30358 = ~new_n30286 & ~new_n30357;
  assign new_n30359 = new_n30358 ^ new_n30356;
  assign new_n30360 = new_n30359 ^ new_n30354;
  assign new_n30361 = new_n30360 ^ new_n30351;
  assign new_n30362 = new_n30361 ^ new_n30348;
  assign new_n30363 = new_n30362 ^ new_n30331;
  assign new_n30364 = new_n28192 ^ new_n28064;
  assign new_n30365 = new_n26036 ^ new_n22447;
  assign new_n30366 = new_n30365 ^ new_n28175;
  assign new_n30367 = new_n30366 ^ new_n28125;
  assign new_n30368 = new_n30367 ^ new_n30364;
  assign new_n30369 = new_n28229 ^ new_n28085;
  assign new_n30370 = new_n30369 ^ new_n28095;
  assign new_n30371 = new_n25010 ^ new_n22472;
  assign new_n30372 = new_n28168 ^ new_n28110;
  assign new_n30373 = new_n30372 ^ new_n30371;
  assign new_n30374 = new_n30373 ^ new_n30370;
  assign new_n30375 = new_n28168 ^ new_n28141;
  assign new_n30376 = new_n30375 ^ new_n28198;
  assign new_n30377 = new_n30376 ^ new_n28129;
  assign new_n30378 = new_n25968 ^ new_n21187;
  assign new_n30379 = new_n30378 ^ new_n28149;
  assign new_n30380 = new_n30379 ^ new_n28080;
  assign new_n30381 = new_n30380 ^ new_n30377;
  assign new_n30382 = new_n28234 ^ new_n27707;
  assign new_n30383 = new_n30382 ^ new_n28218;
  assign new_n30384 = new_n26006 ^ new_n22393;
  assign new_n30385 = new_n30384 ^ new_n28129;
  assign new_n30386 = new_n30385 ^ new_n28089;
  assign new_n30387 = new_n30386 ^ new_n30383;
  assign new_n30388 = new_n30387 ^ new_n30381;
  assign new_n30389 = new_n30388 ^ new_n30374;
  assign new_n30390 = new_n30389 ^ new_n30368;
  assign new_n30391 = new_n26076 ^ new_n22362;
  assign new_n30392 = new_n30391 ^ new_n28198;
  assign new_n30393 = new_n28205 ^ new_n28147;
  assign new_n30394 = new_n30393 ^ new_n28129;
  assign new_n30395 = new_n30394 ^ new_n30392;
  assign new_n30396 = new_n26110 ^ new_n22417;
  assign new_n30397 = new_n30396 ^ new_n28129;
  assign new_n30398 = new_n30397 ^ new_n28235;
  assign new_n30399 = new_n27863 ^ new_n27407;
  assign new_n30400 = new_n30399 ^ new_n28029;
  assign new_n30401 = new_n30400 ^ new_n30398;
  assign new_n30402 = new_n28048 ^ new_n27556;
  assign new_n30403 = new_n26064 ^ new_n22330;
  assign new_n30404 = new_n30403 ^ new_n28004;
  assign new_n30405 = new_n30404 ^ new_n28188;
  assign new_n30406 = new_n30405 ^ new_n30402;
  assign new_n30407 = new_n30406 ^ new_n30368;
  assign new_n30408 = new_n30407 ^ new_n30395;
  assign new_n30409 = new_n30408 ^ new_n30401;
  assign new_n30410 = ~new_n30395 & ~new_n30409;
  assign new_n30411 = new_n30410 ^ new_n30401;
  assign new_n30412 = new_n26100 ^ new_n22261;
  assign new_n30413 = new_n30412 ^ new_n28193;
  assign new_n30414 = new_n28128 ^ new_n28114;
  assign new_n30415 = new_n30414 ^ new_n27978;
  assign new_n30416 = new_n30415 ^ new_n30413;
  assign new_n30417 = new_n30416 ^ new_n30401;
  assign new_n30418 = new_n30417 ^ new_n30388;
  assign new_n30419 = new_n30416 ^ new_n30381;
  assign new_n30420 = new_n30401 ^ new_n30374;
  assign new_n30421 = new_n30420 ^ new_n30419;
  assign new_n30422 = ~new_n30418 & ~new_n30421;
  assign new_n30423 = new_n30422 ^ new_n30368;
  assign new_n30424 = new_n30423 ^ new_n30411;
  assign new_n30425 = new_n30381 & new_n30408;
  assign new_n30426 = new_n30425 ^ new_n30381;
  assign new_n30427 = new_n30406 ^ new_n30389;
  assign new_n30428 = ~new_n30419 & new_n30427;
  assign new_n30429 = new_n30428 ^ new_n30426;
  assign new_n30430 = new_n30416 ^ new_n30374;
  assign new_n30431 = new_n30430 ^ new_n30429;
  assign new_n30432 = new_n30390 & new_n30417;
  assign new_n30433 = new_n30406 ^ new_n30401;
  assign new_n30434 = new_n30433 ^ new_n30430;
  assign new_n30435 = ~new_n30434 & new_n30420;
  assign new_n30436 = new_n30435 ^ new_n30432;
  assign new_n30437 = new_n30406 ^ new_n30387;
  assign new_n30438 = new_n30437 ^ new_n30436;
  assign new_n30439 = new_n30438 ^ new_n30431;
  assign new_n30440 = new_n30423 ^ new_n30418;
  assign new_n30441 = new_n30408 ^ new_n30381;
  assign new_n30442 = new_n30441 ^ new_n30430;
  assign new_n30443 = new_n30418 ^ new_n30395;
  assign new_n30444 = new_n30442 & new_n30443;
  assign new_n30445 = new_n30444 ^ new_n30436;
  assign new_n30446 = new_n30445 ^ new_n30374;
  assign new_n30447 = new_n30446 ^ new_n30440;
  assign new_n30448 = ~new_n30439 & new_n30447;
  assign new_n30449 = new_n30448 ^ new_n30424;
  assign new_n30450 = new_n30418 ^ new_n30407;
  assign new_n30451 = ~new_n30450 & new_n30430;
  assign new_n30452 = new_n30451 ^ new_n30432;
  assign new_n30453 = new_n30452 ^ new_n30427;
  assign new_n30454 = new_n30453 ^ new_n30449;
  assign new_n30455 = new_n30416 ^ new_n30408;
  assign new_n30456 = new_n30395 ^ new_n30390;
  assign new_n30457 = ~new_n30455 & ~new_n30456;
  assign new_n30458 = new_n30457 ^ new_n30425;
  assign new_n30459 = new_n30451 ^ new_n30435;
  assign new_n30460 = new_n30459 ^ new_n30458;
  assign new_n30461 = ~new_n30454 & ~new_n30460;
  assign new_n30462 = new_n30416 ^ new_n30406;
  assign new_n30463 = new_n30444 ^ new_n30410;
  assign new_n30464 = new_n30463 ^ new_n30459;
  assign new_n30465 = new_n30464 ^ new_n30462;
  assign new_n30466 = new_n30457 ^ new_n30428;
  assign new_n30467 = new_n30466 ^ new_n30416;
  assign new_n30468 = new_n30467 ^ new_n30453;
  assign new_n30469 = new_n30468 ^ new_n30448;
  assign new_n30470 = ~new_n30465 & new_n30469;
  assign new_n30471 = new_n30470 ^ new_n30461;
  assign new_n30472 = new_n30467 ^ new_n30424;
  assign new_n30473 = new_n30472 ^ new_n30471;
  assign new_n30474 = ~new_n30473 & new_n30390;
  assign new_n30475 = ~new_n30473 & new_n30417;
  assign new_n30476 = new_n30475 ^ new_n30474;
  assign new_n30477 = new_n30461 ^ new_n30416;
  assign new_n30478 = new_n30457 ^ new_n30410;
  assign new_n30479 = new_n30406 ^ new_n30381;
  assign new_n30480 = new_n30444 ^ new_n30426;
  assign new_n30481 = new_n30470 ^ new_n30424;
  assign new_n30482 = new_n30481 ^ new_n30453;
  assign new_n30483 = new_n30461 ^ new_n30448;
  assign new_n30484 = new_n30468 & new_n30483;
  assign new_n30485 = new_n30484 ^ new_n30469;
  assign new_n30486 = ~new_n30482 & new_n30485;
  assign new_n30487 = new_n30486 ^ new_n30484;
  assign new_n30488 = new_n30487 ^ new_n30480;
  assign new_n30489 = new_n30488 ^ new_n30479;
  assign new_n30490 = new_n30489 ^ new_n30478;
  assign new_n30491 = new_n30490 ^ new_n30477;
  assign new_n30492 = new_n30430 & new_n30491;
  assign new_n30493 = ~new_n30455 & ~new_n30482;
  assign new_n30494 = ~new_n30450 & new_n30491;
  assign new_n30495 = new_n30494 ^ new_n30493;
  assign new_n30496 = new_n30486 ^ new_n30470;
  assign new_n30497 = new_n30496 ^ new_n30447;
  assign new_n30498 = ~new_n30419 & new_n30497;
  assign new_n30499 = new_n30468 ^ new_n30461;
  assign new_n30500 = ~new_n30395 & new_n30499;
  assign new_n30501 = new_n30484 ^ new_n30439;
  assign new_n30502 = ~new_n30418 & ~new_n30501;
  assign new_n30503 = new_n30502 ^ new_n30500;
  assign new_n30504 = new_n30503 ^ new_n30498;
  assign new_n30505 = new_n30504 ^ new_n30495;
  assign new_n30506 = new_n30505 ^ new_n30492;
  assign new_n30507 = new_n30506 ^ new_n30476;
  assign new_n30508 = new_n30507 ^ new_n30363;
  assign new_n30509 = new_n30489 ^ new_n30401;
  assign new_n30510 = new_n30470 ^ new_n30428;
  assign new_n30511 = new_n30510 ^ new_n30423;
  assign new_n30512 = new_n30511 ^ new_n30509;
  assign new_n30513 = ~new_n30434 & ~new_n30512;
  assign new_n30514 = new_n30513 ^ new_n30474;
  assign new_n30515 = new_n30484 ^ new_n30461;
  assign new_n30516 = new_n30515 ^ new_n30460;
  assign new_n30517 = ~new_n30516 & new_n30443;
  assign new_n30518 = new_n30517 ^ new_n30502;
  assign new_n30519 = ~new_n30421 & ~new_n30501;
  assign new_n30520 = new_n30519 ^ new_n30518;
  assign new_n30521 = ~new_n30516 & new_n30442;
  assign new_n30522 = ~new_n30512 & new_n30420;
  assign new_n30523 = new_n30522 ^ new_n30475;
  assign new_n30524 = new_n30523 ^ new_n30521;
  assign new_n30525 = new_n30524 ^ new_n30520;
  assign new_n30526 = new_n30525 ^ new_n30514;
  assign new_n30527 = new_n30526 ^ new_n30508;
  assign new_n30528 = new_n28439 ^ new_n25469;
  assign new_n30529 = new_n26113 ^ new_n26069;
  assign new_n30530 = new_n30529 ^ new_n30528;
  assign new_n30531 = new_n26094 ^ new_n25929;
  assign new_n30532 = new_n30531 ^ new_n30530;
  assign new_n30533 = new_n26112 ^ new_n25993;
  assign new_n30534 = new_n30533 ^ new_n25985;
  assign new_n30535 = new_n30534 ^ new_n30532;
  assign new_n30536 = new_n28458 ^ new_n25486;
  assign new_n30537 = new_n26112 ^ new_n26070;
  assign new_n30538 = new_n30537 ^ new_n30536;
  assign new_n30539 = new_n26054 ^ new_n26016;
  assign new_n30540 = new_n30539 ^ new_n26058;
  assign new_n30541 = new_n30540 ^ new_n30538;
  assign new_n30542 = new_n30541 ^ new_n30535;
  assign new_n30543 = new_n25980 ^ new_n24738;
  assign new_n30544 = new_n30543 ^ new_n25914;
  assign new_n30545 = new_n28465 ^ new_n25453;
  assign new_n30546 = new_n30545 ^ new_n23663;
  assign new_n30547 = new_n30546 ^ new_n25958;
  assign new_n30548 = new_n30547 ^ new_n30544;
  assign new_n30549 = new_n26096 ^ new_n25940;
  assign new_n30550 = new_n30549 ^ new_n26042;
  assign new_n30551 = new_n28468 ^ new_n25465;
  assign new_n30552 = new_n30551 ^ new_n26094;
  assign new_n30553 = new_n30552 ^ new_n26028;
  assign new_n30554 = new_n30553 ^ new_n30550;
  assign new_n30555 = new_n30554 ^ new_n30548;
  assign new_n30556 = new_n30555 ^ new_n30542;
  assign new_n30557 = new_n25950 ^ new_n22574;
  assign new_n30558 = new_n30557 ^ new_n25972;
  assign new_n30559 = new_n30558 ^ new_n30531;
  assign new_n30560 = new_n28479 ^ new_n25447;
  assign new_n30561 = new_n30560 ^ new_n25958;
  assign new_n30562 = new_n30561 ^ new_n26082;
  assign new_n30563 = new_n30562 ^ new_n30559;
  assign new_n30564 = new_n30563 ^ new_n30541;
  assign new_n30565 = new_n26092 ^ new_n26022;
  assign new_n30566 = new_n30565 ^ new_n26047;
  assign new_n30567 = new_n28484 ^ new_n25459;
  assign new_n30568 = new_n30567 ^ new_n26028;
  assign new_n30569 = new_n30568 ^ new_n26058;
  assign new_n30570 = new_n30569 ^ new_n30566;
  assign new_n30571 = new_n30570 ^ new_n30541;
  assign new_n30572 = new_n28488 ^ new_n25482;
  assign new_n30573 = new_n30572 ^ new_n26082;
  assign new_n30574 = new_n26080 ^ new_n25925;
  assign new_n30575 = new_n30574 ^ new_n30531;
  assign new_n30576 = new_n30575 ^ new_n30573;
  assign new_n30577 = new_n30576 ^ new_n30571;
  assign new_n30578 = ~new_n30563 & ~new_n30577;
  assign new_n30579 = new_n30578 ^ new_n30563;
  assign new_n30580 = new_n30577 ^ new_n30563;
  assign new_n30581 = new_n30580 ^ new_n30555;
  assign new_n30582 = new_n30554 ^ new_n30535;
  assign new_n30583 = new_n28499 ^ new_n25438;
  assign new_n30584 = new_n26120 ^ new_n25999;
  assign new_n30585 = new_n30584 ^ new_n30583;
  assign new_n30586 = new_n30585 ^ new_n30531;
  assign new_n30587 = new_n25993 ^ new_n23663;
  assign new_n30588 = new_n30587 ^ new_n25905;
  assign new_n30589 = new_n30588 ^ new_n30586;
  assign new_n30590 = new_n30589 ^ new_n30563;
  assign new_n30591 = new_n30590 ^ new_n30582;
  assign new_n30592 = new_n30591 ^ new_n30576;
  assign new_n30593 = ~new_n30581 & ~new_n30592;
  assign new_n30594 = new_n30593 ^ new_n30579;
  assign new_n30595 = new_n30563 ^ new_n30535;
  assign new_n30596 = new_n30595 ^ new_n30555;
  assign new_n30597 = ~new_n30596 & new_n30591;
  assign new_n30598 = new_n30597 ^ new_n30570;
  assign new_n30599 = ~new_n30576 & new_n30571;
  assign new_n30600 = new_n30535 & new_n30576;
  assign new_n30601 = new_n30600 ^ new_n30599;
  assign new_n30602 = new_n30601 ^ new_n30598;
  assign new_n30603 = new_n30554 ^ new_n30541;
  assign new_n30604 = new_n30591 ^ new_n30571;
  assign new_n30605 = ~new_n30555 & ~new_n30604;
  assign new_n30606 = new_n30548 ^ new_n30535;
  assign new_n30607 = ~new_n30556 & new_n30606;
  assign new_n30608 = new_n30607 ^ new_n30605;
  assign new_n30609 = new_n30601 ^ new_n30535;
  assign new_n30610 = new_n30609 ^ new_n30593;
  assign new_n30611 = new_n30610 ^ new_n30608;
  assign new_n30612 = new_n30611 ^ new_n30603;
  assign new_n30613 = new_n30589 ^ new_n30548;
  assign new_n30614 = new_n30613 ^ new_n30563;
  assign new_n30615 = new_n30614 ^ new_n30570;
  assign new_n30616 = ~new_n30582 & new_n30615;
  assign new_n30617 = new_n30616 ^ new_n30605;
  assign new_n30618 = new_n30614 ^ new_n30541;
  assign new_n30619 = new_n30618 ^ new_n30617;
  assign new_n30620 = new_n30563 ^ new_n30554;
  assign new_n30621 = ~new_n30618 & ~new_n30620;
  assign new_n30622 = new_n30577 ^ new_n30554;
  assign new_n30623 = new_n30615 ^ new_n30576;
  assign new_n30624 = ~new_n30622 & ~new_n30623;
  assign new_n30625 = new_n30624 ^ new_n30621;
  assign new_n30626 = new_n30625 ^ new_n30554;
  assign new_n30627 = new_n30626 ^ new_n30619;
  assign new_n30628 = new_n30621 ^ new_n30579;
  assign new_n30629 = new_n30628 ^ new_n30555;
  assign new_n30630 = new_n30616 ^ new_n30607;
  assign new_n30631 = new_n30589 ^ new_n30541;
  assign new_n30632 = new_n30631 ^ new_n30630;
  assign new_n30633 = new_n30632 ^ new_n30629;
  assign new_n30634 = new_n30598 ^ new_n30591;
  assign new_n30635 = new_n30630 ^ new_n30593;
  assign new_n30636 = new_n30635 ^ new_n30548;
  assign new_n30637 = new_n30636 ^ new_n30634;
  assign new_n30638 = ~new_n30633 & ~new_n30637;
  assign new_n30639 = new_n30638 ^ new_n30627;
  assign new_n30640 = ~new_n30612 & new_n30639;
  assign new_n30641 = new_n30640 ^ new_n30602;
  assign new_n30642 = new_n30641 ^ new_n30619;
  assign new_n30643 = new_n30638 ^ new_n30602;
  assign new_n30644 = new_n30643 ^ new_n30619;
  assign new_n30645 = new_n30624 ^ new_n30578;
  assign new_n30646 = new_n30645 ^ new_n30608;
  assign new_n30647 = ~new_n30646 & new_n30644;
  assign new_n30648 = new_n30647 ^ new_n30638;
  assign new_n30649 = new_n30627 & new_n30648;
  assign new_n30650 = new_n30649 ^ new_n30639;
  assign new_n30651 = new_n30642 & new_n30650;
  assign new_n30652 = new_n30651 ^ new_n30649;
  assign new_n30653 = new_n30652 ^ new_n30594;
  assign new_n30654 = new_n30653 ^ new_n30564;
  assign new_n30655 = new_n30654 ^ new_n30535;
  assign new_n30656 = new_n30640 ^ new_n30621;
  assign new_n30657 = new_n30656 ^ new_n30598;
  assign new_n30658 = new_n30657 ^ new_n30655;
  assign new_n30659 = ~new_n30556 & new_n30658;
  assign new_n30660 = new_n30647 ^ new_n30640;
  assign new_n30661 = new_n30626 ^ new_n30602;
  assign new_n30662 = new_n30661 ^ new_n30660;
  assign new_n30663 = new_n30615 & new_n30662;
  assign new_n30664 = new_n30663 ^ new_n30659;
  assign new_n30665 = new_n30649 ^ new_n30647;
  assign new_n30666 = new_n30665 ^ new_n30646;
  assign new_n30667 = ~new_n30592 & ~new_n30666;
  assign new_n30668 = new_n30649 ^ new_n30633;
  assign new_n30669 = ~new_n30668 & new_n30591;
  assign new_n30670 = new_n30669 ^ new_n30667;
  assign new_n30671 = ~new_n30596 & ~new_n30668;
  assign new_n30672 = new_n30671 ^ new_n30670;
  assign new_n30673 = ~new_n30581 & ~new_n30666;
  assign new_n30674 = new_n30606 & new_n30658;
  assign new_n30675 = ~new_n30582 & new_n30662;
  assign new_n30676 = new_n30675 ^ new_n30674;
  assign new_n30677 = new_n30676 ^ new_n30673;
  assign new_n30678 = new_n30677 ^ new_n30672;
  assign new_n30679 = new_n30678 ^ new_n30664;
  assign new_n30680 = new_n26110 ^ new_n13835;
  assign new_n30681 = new_n26064 ^ new_n13831;
  assign new_n30682 = new_n30681 ^ new_n30680;
  assign new_n30683 = new_n25010 ^ new_n13845;
  assign new_n30684 = new_n26100 ^ new_n13838;
  assign new_n30685 = new_n30684 ^ new_n30683;
  assign new_n30686 = new_n30685 ^ new_n30682;
  assign new_n30687 = new_n25968 ^ new_n13840;
  assign new_n30688 = new_n30687 ^ new_n30681;
  assign new_n30689 = new_n26036 ^ new_n13832;
  assign new_n30690 = new_n30689 ^ new_n30681;
  assign new_n30691 = new_n26076 ^ new_n13830;
  assign new_n30692 = new_n30691 ^ new_n30690;
  assign new_n30693 = ~new_n30687 & ~new_n30692;
  assign new_n30694 = new_n30693 ^ new_n30687;
  assign new_n30695 = new_n30692 ^ new_n30687;
  assign new_n30696 = new_n30695 ^ new_n30685;
  assign new_n30697 = new_n30684 ^ new_n30680;
  assign new_n30698 = new_n26006 ^ new_n13841;
  assign new_n30699 = new_n30698 ^ new_n30687;
  assign new_n30700 = new_n30699 ^ new_n30697;
  assign new_n30701 = new_n30700 ^ new_n30691;
  assign new_n30702 = new_n30696 & new_n30701;
  assign new_n30703 = new_n30702 ^ new_n30694;
  assign new_n30704 = new_n30687 ^ new_n30680;
  assign new_n30705 = new_n30704 ^ new_n30685;
  assign new_n30706 = new_n30700 & new_n30705;
  assign new_n30707 = new_n30706 ^ new_n30689;
  assign new_n30708 = ~new_n30690 & new_n30691;
  assign new_n30709 = ~new_n30691 & new_n30680;
  assign new_n30710 = new_n30709 ^ new_n30708;
  assign new_n30711 = new_n30710 ^ new_n30707;
  assign new_n30712 = new_n30684 ^ new_n30681;
  assign new_n30713 = new_n30700 ^ new_n30690;
  assign new_n30714 = new_n30685 & new_n30713;
  assign new_n30715 = new_n30683 ^ new_n30680;
  assign new_n30716 = new_n30686 & new_n30715;
  assign new_n30717 = new_n30716 ^ new_n30714;
  assign new_n30718 = new_n30710 ^ new_n30680;
  assign new_n30719 = new_n30718 ^ new_n30702;
  assign new_n30720 = new_n30719 ^ new_n30717;
  assign new_n30721 = new_n30720 ^ new_n30712;
  assign new_n30722 = new_n30699 ^ new_n30683;
  assign new_n30723 = new_n30722 ^ new_n30689;
  assign new_n30724 = new_n30697 & new_n30723;
  assign new_n30725 = new_n30724 ^ new_n30714;
  assign new_n30726 = new_n30722 ^ new_n30681;
  assign new_n30727 = new_n30726 ^ new_n30725;
  assign new_n30728 = new_n30687 ^ new_n30684;
  assign new_n30729 = new_n30726 & new_n30728;
  assign new_n30730 = new_n30692 ^ new_n30684;
  assign new_n30731 = new_n30723 ^ new_n30691;
  assign new_n30732 = new_n30730 & new_n30731;
  assign new_n30733 = new_n30732 ^ new_n30729;
  assign new_n30734 = new_n30733 ^ new_n30684;
  assign new_n30735 = new_n30734 ^ new_n30727;
  assign new_n30736 = new_n30729 ^ new_n30694;
  assign new_n30737 = new_n30736 ^ new_n30685;
  assign new_n30738 = new_n30724 ^ new_n30716;
  assign new_n30739 = new_n30698 ^ new_n30681;
  assign new_n30740 = new_n30739 ^ new_n30738;
  assign new_n30741 = new_n30740 ^ new_n30737;
  assign new_n30742 = new_n30707 ^ new_n30700;
  assign new_n30743 = new_n30724 ^ new_n30702;
  assign new_n30744 = new_n30716 ^ new_n30683;
  assign new_n30745 = new_n30744 ^ new_n30743;
  assign new_n30746 = new_n30745 ^ new_n30742;
  assign new_n30747 = ~new_n30741 & new_n30746;
  assign new_n30748 = new_n30747 ^ new_n30735;
  assign new_n30749 = new_n30721 & new_n30748;
  assign new_n30750 = new_n30749 ^ new_n30711;
  assign new_n30751 = new_n30750 ^ new_n30727;
  assign new_n30752 = new_n30747 ^ new_n30711;
  assign new_n30753 = new_n30752 ^ new_n30727;
  assign new_n30754 = new_n30732 ^ new_n30693;
  assign new_n30755 = new_n30754 ^ new_n30717;
  assign new_n30756 = ~new_n30755 & new_n30753;
  assign new_n30757 = new_n30756 ^ new_n30747;
  assign new_n30758 = new_n30735 & new_n30757;
  assign new_n30759 = new_n30758 ^ new_n30748;
  assign new_n30760 = new_n30751 & new_n30759;
  assign new_n30761 = new_n30760 ^ new_n30758;
  assign new_n30762 = new_n30761 ^ new_n30703;
  assign new_n30763 = new_n30762 ^ new_n30688;
  assign new_n30764 = new_n30763 ^ new_n30680;
  assign new_n30765 = new_n30749 ^ new_n30729;
  assign new_n30766 = new_n30765 ^ new_n30707;
  assign new_n30767 = new_n30766 ^ new_n30764;
  assign new_n30768 = ~new_n30767 & new_n30686;
  assign new_n30769 = new_n30756 ^ new_n30749;
  assign new_n30770 = new_n30734 ^ new_n30711;
  assign new_n30771 = new_n30770 ^ new_n30769;
  assign new_n30772 = new_n30723 & new_n30771;
  assign new_n30773 = new_n30772 ^ new_n30768;
  assign new_n30774 = new_n30758 ^ new_n30756;
  assign new_n30775 = new_n30774 ^ new_n30755;
  assign new_n30776 = ~new_n30775 & new_n30701;
  assign new_n30777 = new_n30758 ^ new_n30741;
  assign new_n30778 = ~new_n30777 & new_n30700;
  assign new_n30779 = new_n30778 ^ new_n30776;
  assign new_n30780 = ~new_n30777 & new_n30705;
  assign new_n30781 = new_n30780 ^ new_n30779;
  assign new_n30782 = ~new_n30775 & new_n30696;
  assign new_n30783 = ~new_n30767 & new_n30715;
  assign new_n30784 = new_n30697 & new_n30771;
  assign new_n30785 = new_n30784 ^ new_n30783;
  assign new_n30786 = new_n30785 ^ new_n30782;
  assign new_n30787 = new_n30786 ^ new_n30781;
  assign new_n30788 = new_n30787 ^ new_n30773;
  assign new_n30789 = new_n30788 ^ new_n26397;
  assign new_n30790 = new_n29375 ^ new_n29176;
  assign new_n30791 = new_n30790 ^ new_n28870;
  assign new_n30792 = new_n26604 ^ new_n23442;
  assign new_n30793 = new_n30792 ^ new_n18149;
  assign new_n30794 = new_n30793 ^ new_n29238;
  assign new_n30795 = new_n29246 ^ new_n29002;
  assign new_n30796 = new_n30795 ^ new_n30794;
  assign new_n30797 = new_n30796 ^ new_n30791;
  assign new_n30798 = new_n26959 ^ new_n22682;
  assign new_n30799 = new_n30798 ^ new_n18174;
  assign new_n30800 = new_n30799 ^ new_n29341;
  assign new_n30801 = new_n29169 ^ new_n28725;
  assign new_n30802 = new_n30801 ^ new_n29231;
  assign new_n30803 = new_n30802 ^ new_n30800;
  assign new_n30804 = new_n30803 ^ new_n30797;
  assign new_n30805 = new_n27036 ^ new_n23537;
  assign new_n30806 = new_n30805 ^ new_n18187;
  assign new_n30807 = new_n30806 ^ new_n29385;
  assign new_n30808 = new_n29309 ^ new_n29277;
  assign new_n30809 = new_n30808 ^ new_n29270;
  assign new_n30810 = new_n30809 ^ new_n30807;
  assign new_n30811 = new_n27051 ^ new_n23457;
  assign new_n30812 = new_n30811 ^ new_n18153;
  assign new_n30813 = new_n30812 ^ new_n29154;
  assign new_n30814 = new_n29346 ^ new_n29254;
  assign new_n30815 = new_n30814 ^ new_n29251;
  assign new_n30816 = new_n30815 ^ new_n30813;
  assign new_n30817 = new_n30816 ^ new_n30810;
  assign new_n30818 = new_n30817 ^ new_n30804;
  assign new_n30819 = new_n29358 ^ new_n29320;
  assign new_n30820 = new_n30819 ^ new_n29318;
  assign new_n30821 = new_n27098 ^ new_n23522;
  assign new_n30822 = new_n30821 ^ new_n18159;
  assign new_n30823 = new_n30822 ^ new_n29291;
  assign new_n30824 = new_n30823 ^ new_n30795;
  assign new_n30825 = new_n30824 ^ new_n30820;
  assign new_n30826 = new_n30825 ^ new_n30803;
  assign new_n30827 = new_n27111 ^ new_n23311;
  assign new_n30828 = new_n30827 ^ new_n18170;
  assign new_n30829 = new_n30828 ^ new_n29258;
  assign new_n30830 = new_n29212 ^ new_n29194;
  assign new_n30831 = new_n30830 ^ new_n29350;
  assign new_n30832 = new_n30831 ^ new_n30829;
  assign new_n30833 = new_n30832 ^ new_n30803;
  assign new_n30834 = new_n27130 ^ new_n23385;
  assign new_n30835 = new_n30834 ^ new_n18180;
  assign new_n30836 = new_n30835 ^ new_n29328;
  assign new_n30837 = new_n30795 ^ new_n29361;
  assign new_n30838 = new_n30837 ^ new_n30836;
  assign new_n30839 = new_n30838 ^ new_n30833;
  assign new_n30840 = new_n30825 & new_n30839;
  assign new_n30841 = new_n30840 ^ new_n30825;
  assign new_n30842 = new_n30839 ^ new_n30825;
  assign new_n30843 = new_n30842 ^ new_n30817;
  assign new_n30844 = new_n30816 ^ new_n30797;
  assign new_n30845 = new_n27163 ^ new_n23478;
  assign new_n30846 = new_n30845 ^ new_n18163;
  assign new_n30847 = new_n30846 ^ new_n29164;
  assign new_n30848 = new_n30847 ^ new_n30795;
  assign new_n30849 = new_n29296 ^ new_n29266;
  assign new_n30850 = new_n30849 ^ new_n29380;
  assign new_n30851 = new_n30850 ^ new_n30848;
  assign new_n30852 = new_n30851 ^ new_n30825;
  assign new_n30853 = new_n30852 ^ new_n30844;
  assign new_n30854 = new_n30853 ^ new_n30838;
  assign new_n30855 = new_n30843 & new_n30854;
  assign new_n30856 = new_n30855 ^ new_n30841;
  assign new_n30857 = new_n30825 ^ new_n30797;
  assign new_n30858 = new_n30857 ^ new_n30817;
  assign new_n30859 = ~new_n30853 & ~new_n30858;
  assign new_n30860 = new_n30859 ^ new_n30832;
  assign new_n30861 = ~new_n30833 & ~new_n30838;
  assign new_n30862 = new_n30797 & new_n30838;
  assign new_n30863 = new_n30862 ^ new_n30861;
  assign new_n30864 = new_n30863 ^ new_n30860;
  assign new_n30865 = new_n30816 ^ new_n30803;
  assign new_n30866 = new_n30853 ^ new_n30833;
  assign new_n30867 = ~new_n30866 & new_n30817;
  assign new_n30868 = new_n30810 ^ new_n30797;
  assign new_n30869 = ~new_n30818 & new_n30868;
  assign new_n30870 = new_n30869 ^ new_n30867;
  assign new_n30871 = new_n30863 ^ new_n30797;
  assign new_n30872 = new_n30871 ^ new_n30855;
  assign new_n30873 = new_n30872 ^ new_n30870;
  assign new_n30874 = new_n30873 ^ new_n30865;
  assign new_n30875 = new_n30852 ^ new_n30810;
  assign new_n30876 = new_n30875 ^ new_n30832;
  assign new_n30877 = new_n30844 & new_n30876;
  assign new_n30878 = new_n30877 ^ new_n30867;
  assign new_n30879 = new_n30875 ^ new_n30803;
  assign new_n30880 = new_n30879 ^ new_n30878;
  assign new_n30881 = new_n30825 ^ new_n30816;
  assign new_n30882 = ~new_n30881 & new_n30879;
  assign new_n30883 = new_n30839 ^ new_n30816;
  assign new_n30884 = new_n30876 ^ new_n30838;
  assign new_n30885 = ~new_n30883 & ~new_n30884;
  assign new_n30886 = new_n30885 ^ new_n30882;
  assign new_n30887 = new_n30886 ^ new_n30816;
  assign new_n30888 = new_n30887 ^ new_n30880;
  assign new_n30889 = new_n30882 ^ new_n30841;
  assign new_n30890 = new_n30889 ^ new_n30817;
  assign new_n30891 = new_n30877 ^ new_n30869;
  assign new_n30892 = new_n30851 ^ new_n30803;
  assign new_n30893 = new_n30892 ^ new_n30891;
  assign new_n30894 = new_n30893 ^ new_n30890;
  assign new_n30895 = new_n30860 ^ new_n30853;
  assign new_n30896 = new_n30891 ^ new_n30855;
  assign new_n30897 = new_n30896 ^ new_n30810;
  assign new_n30898 = new_n30897 ^ new_n30895;
  assign new_n30899 = ~new_n30894 & new_n30898;
  assign new_n30900 = new_n30899 ^ new_n30888;
  assign new_n30901 = ~new_n30874 & new_n30900;
  assign new_n30902 = new_n30901 ^ new_n30864;
  assign new_n30903 = new_n30902 ^ new_n30880;
  assign new_n30904 = new_n30899 ^ new_n30864;
  assign new_n30905 = new_n30904 ^ new_n30880;
  assign new_n30906 = new_n30885 ^ new_n30840;
  assign new_n30907 = new_n30906 ^ new_n30870;
  assign new_n30908 = ~new_n30905 & ~new_n30907;
  assign new_n30909 = new_n30908 ^ new_n30899;
  assign new_n30910 = new_n30888 & new_n30909;
  assign new_n30911 = new_n30910 ^ new_n30900;
  assign new_n30912 = ~new_n30903 & new_n30911;
  assign new_n30913 = new_n30912 ^ new_n30910;
  assign new_n30914 = new_n30913 ^ new_n30856;
  assign new_n30915 = new_n30914 ^ new_n30826;
  assign new_n30916 = new_n30915 ^ new_n30797;
  assign new_n30917 = new_n30901 ^ new_n30882;
  assign new_n30918 = new_n30917 ^ new_n30860;
  assign new_n30919 = new_n30918 ^ new_n30916;
  assign new_n30920 = ~new_n30818 & ~new_n30919;
  assign new_n30921 = new_n30908 ^ new_n30901;
  assign new_n30922 = new_n30887 ^ new_n30864;
  assign new_n30923 = new_n30922 ^ new_n30921;
  assign new_n30924 = ~new_n30923 & new_n30876;
  assign new_n30925 = new_n30924 ^ new_n30920;
  assign new_n30926 = new_n30910 ^ new_n30908;
  assign new_n30927 = new_n30926 ^ new_n30907;
  assign new_n30928 = ~new_n30927 & new_n30854;
  assign new_n30929 = new_n30910 ^ new_n30894;
  assign new_n30930 = ~new_n30853 & ~new_n30929;
  assign new_n30931 = new_n30930 ^ new_n30928;
  assign new_n30932 = ~new_n30858 & ~new_n30929;
  assign new_n30933 = new_n30932 ^ new_n30931;
  assign new_n30934 = ~new_n30927 & new_n30843;
  assign new_n30935 = ~new_n30919 & new_n30868;
  assign new_n30936 = ~new_n30923 & new_n30844;
  assign new_n30937 = new_n30936 ^ new_n30935;
  assign new_n30938 = new_n30937 ^ new_n30934;
  assign new_n30939 = new_n30938 ^ new_n30933;
  assign new_n30940 = new_n30939 ^ new_n30925;
  assign new_n30941 = new_n30940 ^ new_n30789;
  assign new_n30942 = new_n30941 ^ new_n30679;
  assign new_n30943 = new_n30942 ^ new_n30527;
  assign new_n30944 = new_n30647 ^ new_n30627;
  assign new_n30945 = new_n30577 ^ new_n30535;
  assign new_n30946 = new_n30944 & new_n30945;
  assign new_n30947 = new_n30651 ^ new_n30640;
  assign new_n30948 = new_n30947 ^ new_n30637;
  assign new_n30949 = ~new_n30618 & ~new_n30948;
  assign new_n30950 = new_n30651 ^ new_n30612;
  assign new_n30951 = ~new_n30950 & new_n30577;
  assign new_n30952 = new_n30951 ^ new_n30677;
  assign new_n30953 = new_n30952 ^ new_n30949;
  assign new_n30954 = new_n30953 ^ new_n30659;
  assign new_n30955 = new_n30954 ^ new_n30946;
  assign new_n30956 = ~new_n30576 & new_n30944;
  assign new_n30957 = new_n30956 ^ new_n30669;
  assign new_n30958 = ~new_n30620 & ~new_n30948;
  assign new_n30959 = new_n30958 ^ new_n30957;
  assign new_n30960 = ~new_n30622 & new_n30642;
  assign new_n30961 = new_n30647 ^ new_n30554;
  assign new_n30962 = new_n30624 ^ new_n30609;
  assign new_n30963 = new_n30962 ^ new_n30654;
  assign new_n30964 = new_n30963 ^ new_n30961;
  assign new_n30965 = ~new_n30604 & new_n30964;
  assign new_n30966 = new_n30965 ^ new_n30960;
  assign new_n30967 = new_n30966 ^ new_n30959;
  assign new_n30968 = new_n30967 ^ new_n30955;
  assign new_n30969 = new_n30908 ^ new_n30888;
  assign new_n30970 = new_n30839 ^ new_n30797;
  assign new_n30971 = ~new_n30970 & new_n30969;
  assign new_n30972 = new_n30912 ^ new_n30901;
  assign new_n30973 = new_n30972 ^ new_n30898;
  assign new_n30974 = new_n30879 & new_n30973;
  assign new_n30975 = new_n30912 ^ new_n30874;
  assign new_n30976 = ~new_n30839 & ~new_n30975;
  assign new_n30977 = new_n30976 ^ new_n30938;
  assign new_n30978 = new_n30977 ^ new_n30974;
  assign new_n30979 = new_n30978 ^ new_n30920;
  assign new_n30980 = new_n30979 ^ new_n30971;
  assign new_n30981 = ~new_n30838 & new_n30969;
  assign new_n30982 = new_n30981 ^ new_n30930;
  assign new_n30983 = ~new_n30881 & new_n30973;
  assign new_n30984 = new_n30983 ^ new_n30982;
  assign new_n30985 = ~new_n30883 & ~new_n30903;
  assign new_n30986 = new_n30908 ^ new_n30816;
  assign new_n30987 = new_n30885 ^ new_n30871;
  assign new_n30988 = new_n30987 ^ new_n30915;
  assign new_n30989 = new_n30988 ^ new_n30986;
  assign new_n30990 = ~new_n30866 & new_n30989;
  assign new_n30991 = new_n30990 ^ new_n30985;
  assign new_n30992 = new_n30991 ^ new_n30984;
  assign new_n30993 = new_n30992 ^ new_n30980;
  assign new_n30994 = ~new_n30409 & new_n30499;
  assign new_n30995 = new_n30486 ^ new_n30465;
  assign new_n30996 = ~new_n30408 & ~new_n30995;
  assign new_n30997 = new_n30996 ^ new_n30524;
  assign new_n30998 = new_n30427 & new_n30497;
  assign new_n30999 = new_n30998 ^ new_n30997;
  assign new_n31000 = new_n30999 ^ new_n30513;
  assign new_n31001 = new_n31000 ^ new_n30994;
  assign new_n31002 = new_n31001 ^ new_n30505;
  assign new_n31003 = new_n31002 ^ new_n30993;
  assign new_n31004 = new_n31003 ^ new_n30968;
  assign new_n31005 = new_n30756 ^ new_n30735;
  assign new_n31006 = new_n30692 ^ new_n30680;
  assign new_n31007 = new_n31005 & new_n31006;
  assign new_n31008 = new_n30760 ^ new_n30749;
  assign new_n31009 = new_n31008 ^ new_n30746;
  assign new_n31010 = new_n30726 & new_n31009;
  assign new_n31011 = new_n30760 ^ new_n30721;
  assign new_n31012 = new_n30692 & new_n31011;
  assign new_n31013 = new_n31012 ^ new_n30786;
  assign new_n31014 = new_n31013 ^ new_n31010;
  assign new_n31015 = new_n31014 ^ new_n30768;
  assign new_n31016 = new_n31015 ^ new_n31007;
  assign new_n31017 = new_n30691 & new_n31005;
  assign new_n31018 = new_n31017 ^ new_n30778;
  assign new_n31019 = new_n30728 & new_n31009;
  assign new_n31020 = new_n31019 ^ new_n31018;
  assign new_n31021 = new_n30730 & new_n30751;
  assign new_n31022 = new_n30756 ^ new_n30684;
  assign new_n31023 = new_n30732 ^ new_n30718;
  assign new_n31024 = new_n31023 ^ new_n30763;
  assign new_n31025 = new_n31024 ^ new_n31022;
  assign new_n31026 = ~new_n31025 & new_n30713;
  assign new_n31027 = new_n31026 ^ new_n31021;
  assign new_n31028 = new_n31027 ^ new_n31020;
  assign new_n31029 = new_n31028 ^ new_n31016;
  assign new_n31030 = new_n31029 ^ new_n26376;
  assign new_n31031 = new_n30354 ^ new_n30350;
  assign new_n31032 = new_n30345 ^ new_n30275;
  assign new_n31033 = new_n30318 ^ new_n30265;
  assign new_n31034 = new_n31033 ^ new_n30290;
  assign new_n31035 = new_n31034 ^ new_n31032;
  assign new_n31036 = ~new_n30277 & ~new_n31035;
  assign new_n31037 = new_n30341 ^ new_n30317;
  assign new_n31038 = ~new_n30255 & ~new_n31037;
  assign new_n31039 = new_n31038 ^ new_n31036;
  assign new_n31040 = ~new_n30305 & ~new_n30337;
  assign new_n31041 = ~new_n31037 & new_n30293;
  assign new_n31042 = new_n31041 ^ new_n31040;
  assign new_n31043 = ~new_n31035 & new_n30278;
  assign new_n31044 = new_n31043 ^ new_n30330;
  assign new_n31045 = new_n31044 ^ new_n31042;
  assign new_n31046 = new_n31045 ^ new_n31039;
  assign new_n31047 = new_n31046 ^ new_n31031;
  assign new_n31048 = new_n30498 ^ new_n30494;
  assign new_n31049 = new_n30996 ^ new_n30513;
  assign new_n31050 = ~new_n30456 & ~new_n30482;
  assign new_n31051 = ~new_n30995 & new_n30441;
  assign new_n31052 = new_n31051 ^ new_n31050;
  assign new_n31053 = new_n31052 ^ new_n30523;
  assign new_n31054 = new_n31053 ^ new_n31049;
  assign new_n31055 = new_n31054 ^ new_n31048;
  assign new_n31056 = new_n31055 ^ new_n31047;
  assign new_n31057 = new_n31056 ^ new_n31030;
  assign new_n31058 = new_n31057 ^ new_n31004;
  assign new_n31059 = ~new_n30623 & new_n30642;
  assign new_n31060 = new_n31059 ^ new_n30671;
  assign new_n31061 = new_n30956 ^ new_n30667;
  assign new_n31062 = new_n31061 ^ new_n30952;
  assign new_n31063 = new_n31062 ^ new_n31060;
  assign new_n31064 = ~new_n30884 & ~new_n30903;
  assign new_n31065 = new_n31064 ^ new_n30932;
  assign new_n31066 = new_n30981 ^ new_n30928;
  assign new_n31067 = new_n31066 ^ new_n30977;
  assign new_n31068 = new_n31067 ^ new_n31065;
  assign new_n31069 = new_n31050 ^ new_n30519;
  assign new_n31070 = new_n30517 ^ new_n30500;
  assign new_n31071 = new_n31070 ^ new_n30997;
  assign new_n31072 = new_n31071 ^ new_n31069;
  assign new_n31073 = new_n31072 ^ new_n31068;
  assign new_n31074 = new_n31073 ^ new_n31063;
  assign new_n31075 = ~new_n30312 & new_n30355;
  assign new_n31076 = new_n30342 ^ new_n30325;
  assign new_n31077 = new_n31076 ^ new_n30324;
  assign new_n31078 = ~new_n31077 & new_n30294;
  assign new_n31079 = new_n31078 ^ new_n31044;
  assign new_n31080 = new_n31079 ^ new_n31038;
  assign new_n31081 = new_n30258 & new_n30353;
  assign new_n31082 = new_n31081 ^ new_n31080;
  assign new_n31083 = new_n31082 ^ new_n31036;
  assign new_n31084 = new_n31083 ^ new_n31075;
  assign new_n31085 = new_n31084 ^ new_n30361;
  assign new_n31086 = new_n31085 ^ new_n31002;
  assign new_n31087 = new_n30731 & new_n30751;
  assign new_n31088 = new_n31087 ^ new_n30780;
  assign new_n31089 = new_n31017 ^ new_n30776;
  assign new_n31090 = new_n31089 ^ new_n31013;
  assign new_n31091 = new_n31090 ^ new_n31088;
  assign new_n31092 = new_n31091 ^ new_n26369;
  assign new_n31093 = ~new_n30288 & ~new_n30357;
  assign new_n31094 = new_n31093 ^ new_n30329;
  assign new_n31095 = new_n31094 ^ new_n31083;
  assign new_n31096 = new_n30519 ^ new_n30474;
  assign new_n31097 = new_n31096 ^ new_n31000;
  assign new_n31098 = new_n31097 ^ new_n31095;
  assign new_n31099 = new_n31098 ^ new_n31092;
  assign new_n31100 = new_n31099 ^ new_n31086;
  assign new_n31101 = new_n31100 ^ new_n31074;
  assign new_n31102 = new_n31098 ^ new_n31055;
  assign new_n31103 = new_n30998 ^ new_n30504;
  assign new_n31104 = new_n31103 ^ new_n31053;
  assign new_n31105 = new_n31081 ^ new_n30360;
  assign new_n31106 = new_n31105 ^ new_n31045;
  assign new_n31107 = new_n31106 ^ new_n31104;
  assign new_n31108 = new_n31107 ^ new_n31102;
  assign new_n31109 = new_n30965 ^ new_n30958;
  assign new_n31110 = ~new_n30950 & new_n30580;
  assign new_n31111 = new_n31110 ^ new_n31059;
  assign new_n31112 = new_n31111 ^ new_n30676;
  assign new_n31113 = new_n30951 ^ new_n30659;
  assign new_n31114 = new_n31113 ^ new_n31112;
  assign new_n31115 = new_n31114 ^ new_n31109;
  assign new_n31116 = new_n31026 ^ new_n31019;
  assign new_n31117 = new_n30695 & new_n31011;
  assign new_n31118 = new_n31117 ^ new_n31087;
  assign new_n31119 = new_n31118 ^ new_n30785;
  assign new_n31120 = new_n31012 ^ new_n30768;
  assign new_n31121 = new_n31120 ^ new_n31119;
  assign new_n31122 = new_n31121 ^ new_n31116;
  assign new_n31123 = new_n31122 ^ new_n26363;
  assign new_n31124 = new_n30990 ^ new_n30983;
  assign new_n31125 = ~new_n30975 & new_n30842;
  assign new_n31126 = new_n31125 ^ new_n31064;
  assign new_n31127 = new_n31126 ^ new_n30937;
  assign new_n31128 = new_n30976 ^ new_n30920;
  assign new_n31129 = new_n31128 ^ new_n31127;
  assign new_n31130 = new_n31129 ^ new_n31124;
  assign new_n31131 = new_n31130 ^ new_n31123;
  assign new_n31132 = new_n31131 ^ new_n31115;
  assign new_n31133 = new_n31132 ^ new_n31108;
  assign new_n31134 = new_n31133 ^ new_n31101;
  assign new_n31135 = new_n31134 ^ new_n31058;
  assign new_n31136 = new_n31135 ^ new_n30943;
  assign new_n31137 = new_n31104 ^ new_n31098;
  assign new_n31138 = new_n30959 ^ new_n30949;
  assign new_n31139 = new_n31138 ^ new_n31112;
  assign new_n31140 = new_n31020 ^ new_n31010;
  assign new_n31141 = new_n31140 ^ new_n31119;
  assign new_n31142 = new_n31141 ^ new_n26410;
  assign new_n31143 = new_n30984 ^ new_n30974;
  assign new_n31144 = new_n31143 ^ new_n31127;
  assign new_n31145 = new_n31144 ^ new_n31142;
  assign new_n31146 = new_n31145 ^ new_n31139;
  assign new_n31147 = new_n31146 ^ new_n31137;
  assign new_n31148 = new_n31093 ^ new_n31040;
  assign new_n31149 = ~new_n31077 & new_n30292;
  assign new_n31150 = new_n31149 ^ new_n30356;
  assign new_n31151 = new_n31150 ^ new_n31080;
  assign new_n31152 = new_n31151 ^ new_n31148;
  assign new_n31153 = new_n31152 ^ new_n31072;
  assign new_n31154 = new_n31014 ^ new_n30781;
  assign new_n31155 = new_n31154 ^ new_n26388;
  assign new_n31156 = new_n31155 ^ new_n31098;
  assign new_n31157 = new_n31156 ^ new_n31153;
  assign new_n31158 = new_n30978 ^ new_n30933;
  assign new_n31159 = new_n30953 ^ new_n30672;
  assign new_n31160 = new_n30999 ^ new_n30520;
  assign new_n31161 = new_n31160 ^ new_n31159;
  assign new_n31162 = new_n31161 ^ new_n31158;
  assign new_n31163 = new_n31162 ^ new_n31157;
  assign new_n31164 = new_n31149 ^ new_n30358;
  assign new_n31165 = new_n31164 ^ new_n31093;
  assign new_n31166 = new_n31165 ^ new_n31082;
  assign new_n31167 = new_n31166 ^ new_n31160;
  assign new_n31168 = new_n31167 ^ new_n30507;
  assign new_n31169 = new_n30675 ^ new_n30663;
  assign new_n31170 = ~new_n30555 & new_n30964;
  assign new_n31171 = new_n31170 ^ new_n30967;
  assign new_n31172 = new_n31171 ^ new_n31169;
  assign new_n31173 = new_n30784 ^ new_n30772;
  assign new_n31174 = ~new_n31025 & new_n30685;
  assign new_n31175 = new_n31174 ^ new_n31028;
  assign new_n31176 = new_n31175 ^ new_n31173;
  assign new_n31177 = new_n31176 ^ new_n26357;
  assign new_n31178 = new_n30936 ^ new_n30924;
  assign new_n31179 = new_n30817 & new_n30989;
  assign new_n31180 = new_n31179 ^ new_n30992;
  assign new_n31181 = new_n31180 ^ new_n31178;
  assign new_n31182 = new_n31181 ^ new_n31177;
  assign new_n31183 = new_n31182 ^ new_n31172;
  assign new_n31184 = new_n31183 ^ new_n31168;
  assign new_n31185 = new_n31184 ^ new_n30943;
  assign new_n31186 = new_n31185 ^ new_n31147;
  assign new_n31187 = new_n31186 ^ new_n31163;
  assign new_n31188 = new_n31147 & new_n31187;
  assign new_n31189 = new_n31188 ^ new_n31163;
  assign new_n31190 = new_n30780 ^ new_n30772;
  assign new_n31191 = new_n31190 ^ new_n31015;
  assign new_n31192 = new_n31191 ^ new_n26381;
  assign new_n31193 = new_n31036 ^ new_n30329;
  assign new_n31194 = new_n31165 ^ new_n31079;
  assign new_n31195 = new_n31194 ^ new_n31193;
  assign new_n31196 = new_n31195 ^ new_n30526;
  assign new_n31197 = new_n31196 ^ new_n31192;
  assign new_n31198 = new_n30932 ^ new_n30924;
  assign new_n31199 = new_n31198 ^ new_n30979;
  assign new_n31200 = new_n30671 ^ new_n30663;
  assign new_n31201 = new_n31200 ^ new_n30954;
  assign new_n31202 = new_n31201 ^ new_n31097;
  assign new_n31203 = new_n31202 ^ new_n31199;
  assign new_n31204 = new_n31203 ^ new_n31197;
  assign new_n31205 = new_n31204 ^ new_n31163;
  assign new_n31206 = new_n31205 ^ new_n31134;
  assign new_n31207 = new_n31204 ^ new_n31133;
  assign new_n31208 = new_n31163 ^ new_n31058;
  assign new_n31209 = new_n31208 ^ new_n31207;
  assign new_n31210 = new_n31206 & new_n31209;
  assign new_n31211 = new_n31210 ^ new_n30943;
  assign new_n31212 = new_n31211 ^ new_n31189;
  assign new_n31213 = ~new_n31133 & ~new_n31186;
  assign new_n31214 = new_n31213 ^ new_n31133;
  assign new_n31215 = new_n31184 ^ new_n31135;
  assign new_n31216 = new_n31207 & new_n31215;
  assign new_n31217 = new_n31216 ^ new_n31214;
  assign new_n31218 = new_n31204 ^ new_n31058;
  assign new_n31219 = new_n31218 ^ new_n31217;
  assign new_n31220 = new_n31136 & new_n31205;
  assign new_n31221 = new_n31184 ^ new_n31163;
  assign new_n31222 = new_n31221 ^ new_n31218;
  assign new_n31223 = new_n31208 & new_n31222;
  assign new_n31224 = new_n31223 ^ new_n31220;
  assign new_n31225 = new_n31184 ^ new_n31101;
  assign new_n31226 = new_n31225 ^ new_n31224;
  assign new_n31227 = new_n31226 ^ new_n31219;
  assign new_n31228 = new_n31211 ^ new_n31206;
  assign new_n31229 = new_n31186 ^ new_n31133;
  assign new_n31230 = new_n31229 ^ new_n31218;
  assign new_n31231 = new_n31206 ^ new_n31147;
  assign new_n31232 = new_n31230 & new_n31231;
  assign new_n31233 = new_n31232 ^ new_n31220;
  assign new_n31234 = new_n31223 ^ new_n31058;
  assign new_n31235 = new_n31234 ^ new_n31233;
  assign new_n31236 = new_n31235 ^ new_n31228;
  assign new_n31237 = ~new_n31227 & new_n31236;
  assign new_n31238 = new_n31237 ^ new_n31212;
  assign new_n31239 = new_n31206 ^ new_n31185;
  assign new_n31240 = new_n31218 & new_n31239;
  assign new_n31241 = new_n31240 ^ new_n31220;
  assign new_n31242 = new_n31241 ^ new_n31215;
  assign new_n31243 = new_n31242 ^ new_n31238;
  assign new_n31244 = new_n31204 ^ new_n31186;
  assign new_n31245 = new_n31147 ^ new_n31136;
  assign new_n31246 = new_n31244 & new_n31245;
  assign new_n31247 = new_n31246 ^ new_n31213;
  assign new_n31248 = new_n31240 ^ new_n31223;
  assign new_n31249 = new_n31248 ^ new_n31247;
  assign new_n31250 = ~new_n31249 & new_n31243;
  assign new_n31251 = new_n31204 ^ new_n31184;
  assign new_n31252 = new_n31232 ^ new_n31188;
  assign new_n31253 = new_n31252 ^ new_n31248;
  assign new_n31254 = new_n31253 ^ new_n31251;
  assign new_n31255 = new_n31246 ^ new_n31216;
  assign new_n31256 = new_n31255 ^ new_n31204;
  assign new_n31257 = new_n31256 ^ new_n31242;
  assign new_n31258 = new_n31257 ^ new_n31237;
  assign new_n31259 = new_n31254 & new_n31258;
  assign new_n31260 = new_n31259 ^ new_n31250;
  assign new_n31261 = new_n31256 ^ new_n31212;
  assign new_n31262 = new_n31261 ^ new_n31260;
  assign new_n31263 = new_n31136 & new_n31262;
  assign new_n31264 = new_n31250 ^ new_n31237;
  assign new_n31265 = new_n31257 & new_n31264;
  assign new_n31266 = new_n31265 ^ new_n31227;
  assign new_n31267 = ~new_n31266 & new_n31209;
  assign new_n31268 = new_n31267 ^ new_n31263;
  assign new_n31269 = new_n31184 ^ new_n31133;
  assign new_n31270 = new_n31232 ^ new_n31214;
  assign new_n31271 = new_n31259 ^ new_n31212;
  assign new_n31272 = new_n31271 ^ new_n31242;
  assign new_n31273 = new_n31265 ^ new_n31258;
  assign new_n31274 = new_n31272 & new_n31273;
  assign new_n31275 = new_n31274 ^ new_n31265;
  assign new_n31276 = new_n31275 ^ new_n31270;
  assign new_n31277 = new_n31276 ^ new_n31269;
  assign new_n31278 = new_n31277 ^ new_n31163;
  assign new_n31279 = new_n31259 ^ new_n31216;
  assign new_n31280 = new_n31279 ^ new_n31211;
  assign new_n31281 = new_n31280 ^ new_n31278;
  assign new_n31282 = ~new_n31281 & new_n31222;
  assign new_n31283 = new_n31274 ^ new_n31254;
  assign new_n31284 = new_n31186 & new_n31283;
  assign new_n31285 = new_n31265 ^ new_n31250;
  assign new_n31286 = new_n31285 ^ new_n31249;
  assign new_n31287 = ~new_n31286 & new_n31230;
  assign new_n31288 = ~new_n31281 & new_n31208;
  assign new_n31289 = new_n31205 & new_n31262;
  assign new_n31290 = new_n31289 ^ new_n31288;
  assign new_n31291 = new_n31290 ^ new_n31287;
  assign new_n31292 = new_n31291 ^ new_n31284;
  assign new_n31293 = new_n31274 ^ new_n31259;
  assign new_n31294 = new_n31293 ^ new_n31236;
  assign new_n31295 = new_n31215 & new_n31294;
  assign new_n31296 = new_n31295 ^ new_n31292;
  assign new_n31297 = new_n31296 ^ new_n31282;
  assign new_n31298 = new_n31297 ^ new_n31268;
  assign new_n31299 = new_n28590 ^ new_n16210;
  assign new_n31300 = new_n29593 ^ new_n15733;
  assign new_n31301 = new_n29649 ^ new_n16149;
  assign new_n31302 = new_n29688 ^ new_n16131;
  assign new_n31303 = new_n31302 ^ new_n31301;
  assign new_n31304 = new_n31303 ^ new_n31300;
  assign new_n31305 = new_n31304 ^ new_n31299;
  assign new_n31306 = new_n29698 ^ new_n16279;
  assign new_n31307 = new_n29709 ^ new_n16263;
  assign new_n31308 = new_n29739 ^ new_n16254;
  assign new_n31309 = new_n31308 ^ new_n31299;
  assign new_n31310 = new_n31309 ^ new_n31306;
  assign new_n31311 = new_n31310 ^ new_n31307;
  assign new_n31312 = ~new_n31306 & ~new_n31311;
  assign new_n31313 = new_n31312 ^ new_n31307;
  assign new_n31314 = new_n29763 ^ new_n16233;
  assign new_n31315 = new_n31314 ^ new_n31307;
  assign new_n31316 = new_n31315 ^ new_n31303;
  assign new_n31317 = new_n31307 ^ new_n31302;
  assign new_n31318 = new_n31314 ^ new_n31300;
  assign new_n31319 = new_n31318 ^ new_n31317;
  assign new_n31320 = ~new_n31316 & ~new_n31319;
  assign new_n31321 = new_n31320 ^ new_n31299;
  assign new_n31322 = new_n31321 ^ new_n31313;
  assign new_n31323 = new_n31302 & new_n31310;
  assign new_n31324 = new_n31323 ^ new_n31302;
  assign new_n31325 = new_n31308 ^ new_n31304;
  assign new_n31326 = new_n31314 ^ new_n31302;
  assign new_n31327 = ~new_n31326 & new_n31325;
  assign new_n31328 = new_n31327 ^ new_n31324;
  assign new_n31329 = new_n31328 ^ new_n31318;
  assign new_n31330 = new_n31305 & new_n31315;
  assign new_n31331 = new_n31308 ^ new_n31307;
  assign new_n31332 = new_n31331 ^ new_n31318;
  assign new_n31333 = new_n31307 ^ new_n31300;
  assign new_n31334 = ~new_n31332 & new_n31333;
  assign new_n31335 = new_n31334 ^ new_n31330;
  assign new_n31336 = new_n31308 ^ new_n31301;
  assign new_n31337 = new_n31336 ^ new_n31335;
  assign new_n31338 = new_n31337 ^ new_n31329;
  assign new_n31339 = new_n31321 ^ new_n31316;
  assign new_n31340 = new_n31310 ^ new_n31302;
  assign new_n31341 = new_n31340 ^ new_n31318;
  assign new_n31342 = new_n31316 ^ new_n31306;
  assign new_n31343 = new_n31341 & new_n31342;
  assign new_n31344 = new_n31343 ^ new_n31300;
  assign new_n31345 = new_n31344 ^ new_n31335;
  assign new_n31346 = new_n31345 ^ new_n31339;
  assign new_n31347 = ~new_n31338 & new_n31346;
  assign new_n31348 = new_n31347 ^ new_n31322;
  assign new_n31349 = new_n31316 ^ new_n31309;
  assign new_n31350 = ~new_n31349 & new_n31318;
  assign new_n31351 = new_n31350 ^ new_n31330;
  assign new_n31352 = new_n31351 ^ new_n31325;
  assign new_n31353 = new_n31352 ^ new_n31348;
  assign new_n31354 = new_n31314 ^ new_n31310;
  assign new_n31355 = new_n31306 ^ new_n31305;
  assign new_n31356 = ~new_n31354 & ~new_n31355;
  assign new_n31357 = new_n31356 ^ new_n31323;
  assign new_n31358 = new_n31350 ^ new_n31334;
  assign new_n31359 = new_n31358 ^ new_n31357;
  assign new_n31360 = ~new_n31353 & ~new_n31359;
  assign new_n31361 = new_n31314 ^ new_n31308;
  assign new_n31362 = new_n31343 ^ new_n31312;
  assign new_n31363 = new_n31362 ^ new_n31358;
  assign new_n31364 = new_n31363 ^ new_n31361;
  assign new_n31365 = new_n31356 ^ new_n31327;
  assign new_n31366 = new_n31365 ^ new_n31314;
  assign new_n31367 = new_n31366 ^ new_n31352;
  assign new_n31368 = new_n31367 ^ new_n31347;
  assign new_n31369 = ~new_n31364 & new_n31368;
  assign new_n31370 = new_n31369 ^ new_n31360;
  assign new_n31371 = new_n31366 ^ new_n31322;
  assign new_n31372 = new_n31371 ^ new_n31370;
  assign new_n31373 = ~new_n31372 & new_n31305;
  assign new_n31374 = new_n31360 ^ new_n31347;
  assign new_n31375 = new_n31367 & new_n31374;
  assign new_n31376 = new_n31375 ^ new_n31338;
  assign new_n31377 = ~new_n31319 & ~new_n31376;
  assign new_n31378 = new_n31377 ^ new_n31373;
  assign new_n31379 = new_n31308 ^ new_n31302;
  assign new_n31380 = new_n31343 ^ new_n31324;
  assign new_n31381 = new_n31369 ^ new_n31322;
  assign new_n31382 = new_n31381 ^ new_n31352;
  assign new_n31383 = new_n31375 ^ new_n31368;
  assign new_n31384 = ~new_n31382 & new_n31383;
  assign new_n31385 = new_n31384 ^ new_n31375;
  assign new_n31386 = new_n31385 ^ new_n31380;
  assign new_n31387 = new_n31386 ^ new_n31379;
  assign new_n31388 = new_n31387 ^ new_n31307;
  assign new_n31389 = new_n31369 ^ new_n31327;
  assign new_n31390 = new_n31389 ^ new_n31321;
  assign new_n31391 = new_n31390 ^ new_n31388;
  assign new_n31392 = ~new_n31332 & ~new_n31391;
  assign new_n31393 = new_n31384 ^ new_n31364;
  assign new_n31394 = ~new_n31310 & ~new_n31393;
  assign new_n31395 = new_n31375 ^ new_n31360;
  assign new_n31396 = new_n31395 ^ new_n31359;
  assign new_n31397 = ~new_n31396 & new_n31341;
  assign new_n31398 = ~new_n31391 & new_n31333;
  assign new_n31399 = ~new_n31372 & new_n31315;
  assign new_n31400 = new_n31399 ^ new_n31398;
  assign new_n31401 = new_n31400 ^ new_n31397;
  assign new_n31402 = new_n31401 ^ new_n31394;
  assign new_n31403 = new_n31384 ^ new_n31369;
  assign new_n31404 = new_n31403 ^ new_n31346;
  assign new_n31405 = new_n31325 & new_n31404;
  assign new_n31406 = new_n31405 ^ new_n31402;
  assign new_n31407 = new_n31406 ^ new_n31392;
  assign new_n31408 = new_n31407 ^ new_n31378;
  assign new_n31409 = new_n31408 ^ new_n22590;
  assign new_n31410 = new_n31409 ^ new_n31298;
  assign new_n31411 = new_n31392 ^ new_n31373;
  assign new_n31412 = ~new_n31316 & ~new_n31376;
  assign new_n31413 = ~new_n31396 & new_n31342;
  assign new_n31414 = new_n31413 ^ new_n31412;
  assign new_n31415 = new_n31414 ^ new_n31377;
  assign new_n31416 = new_n31415 ^ new_n31401;
  assign new_n31417 = new_n31416 ^ new_n31411;
  assign new_n31418 = new_n31417 ^ new_n22580;
  assign new_n31419 = new_n31282 ^ new_n31263;
  assign new_n31420 = ~new_n31266 & new_n31206;
  assign new_n31421 = ~new_n31286 & new_n31231;
  assign new_n31422 = new_n31421 ^ new_n31420;
  assign new_n31423 = new_n31422 ^ new_n31267;
  assign new_n31424 = new_n31423 ^ new_n31291;
  assign new_n31425 = new_n31424 ^ new_n31419;
  assign new_n31426 = new_n31425 ^ new_n31418;
  assign new_n31427 = new_n31399 ^ new_n31373;
  assign new_n31428 = new_n31360 ^ new_n31314;
  assign new_n31429 = new_n31356 ^ new_n31312;
  assign new_n31430 = new_n31429 ^ new_n31387;
  assign new_n31431 = new_n31430 ^ new_n31428;
  assign new_n31432 = new_n31318 & new_n31431;
  assign new_n31433 = ~new_n31326 & new_n31404;
  assign new_n31434 = new_n31367 ^ new_n31360;
  assign new_n31435 = ~new_n31306 & new_n31434;
  assign new_n31436 = new_n31435 ^ new_n31412;
  assign new_n31437 = new_n31436 ^ new_n31433;
  assign new_n31438 = ~new_n31349 & new_n31431;
  assign new_n31439 = ~new_n31354 & ~new_n31382;
  assign new_n31440 = new_n31439 ^ new_n31438;
  assign new_n31441 = new_n31440 ^ new_n31437;
  assign new_n31442 = new_n31441 ^ new_n31432;
  assign new_n31443 = new_n31442 ^ new_n31427;
  assign new_n31444 = new_n31443 ^ new_n22583;
  assign new_n31445 = new_n31289 ^ new_n31263;
  assign new_n31446 = new_n31250 ^ new_n31204;
  assign new_n31447 = new_n31246 ^ new_n31188;
  assign new_n31448 = new_n31447 ^ new_n31277;
  assign new_n31449 = new_n31448 ^ new_n31446;
  assign new_n31450 = ~new_n31449 & new_n31218;
  assign new_n31451 = new_n31207 & new_n31294;
  assign new_n31452 = new_n31257 ^ new_n31250;
  assign new_n31453 = new_n31147 & new_n31452;
  assign new_n31454 = new_n31453 ^ new_n31420;
  assign new_n31455 = new_n31454 ^ new_n31451;
  assign new_n31456 = ~new_n31449 & new_n31239;
  assign new_n31457 = new_n31244 & new_n31272;
  assign new_n31458 = new_n31457 ^ new_n31456;
  assign new_n31459 = new_n31458 ^ new_n31455;
  assign new_n31460 = new_n31459 ^ new_n31450;
  assign new_n31461 = new_n31460 ^ new_n31445;
  assign new_n31462 = new_n31461 ^ new_n31444;
  assign new_n31463 = new_n31423 ^ new_n31296;
  assign new_n31464 = new_n31415 ^ new_n31406;
  assign new_n31465 = new_n31464 ^ new_n22586;
  assign new_n31466 = new_n31465 ^ new_n31463;
  assign new_n31467 = new_n31245 & new_n31272;
  assign new_n31468 = new_n31467 ^ new_n31267;
  assign new_n31469 = new_n31453 ^ new_n31421;
  assign new_n31470 = new_n31469 ^ new_n31292;
  assign new_n31471 = new_n31470 ^ new_n31468;
  assign new_n31472 = ~new_n31355 & ~new_n31382;
  assign new_n31473 = new_n31472 ^ new_n31377;
  assign new_n31474 = new_n31435 ^ new_n31413;
  assign new_n31475 = new_n31474 ^ new_n31402;
  assign new_n31476 = new_n31475 ^ new_n31473;
  assign new_n31477 = new_n31476 ^ new_n22575;
  assign new_n31478 = new_n31477 ^ new_n31471;
  assign new_n31479 = new_n31187 & new_n31452;
  assign new_n31480 = new_n31479 ^ new_n31297;
  assign new_n31481 = new_n31480 ^ new_n31459;
  assign new_n31482 = ~new_n31311 & new_n31434;
  assign new_n31483 = new_n31482 ^ new_n31407;
  assign new_n31484 = new_n31483 ^ new_n31441;
  assign new_n31485 = new_n31484 ^ new_n22578;
  assign new_n31486 = new_n31485 ^ new_n31481;
  assign new_n31487 = new_n31438 ^ new_n31433;
  assign new_n31488 = ~new_n31393 & new_n31340;
  assign new_n31489 = new_n31488 ^ new_n31472;
  assign new_n31490 = new_n31489 ^ new_n31400;
  assign new_n31491 = new_n31394 ^ new_n31392;
  assign new_n31492 = new_n31491 ^ new_n31490;
  assign new_n31493 = new_n31492 ^ new_n31487;
  assign new_n31494 = new_n31493 ^ new_n22576;
  assign new_n31495 = new_n31456 ^ new_n31451;
  assign new_n31496 = new_n31229 & new_n31283;
  assign new_n31497 = new_n31496 ^ new_n31467;
  assign new_n31498 = new_n31497 ^ new_n31290;
  assign new_n31499 = new_n31284 ^ new_n31282;
  assign new_n31500 = new_n31499 ^ new_n31498;
  assign new_n31501 = new_n31500 ^ new_n31495;
  assign new_n31502 = new_n31501 ^ new_n31494;
  assign new_n31503 = new_n31437 ^ new_n31405;
  assign new_n31504 = new_n31503 ^ new_n31490;
  assign new_n31505 = new_n31504 ^ new_n22582;
  assign new_n31506 = new_n31455 ^ new_n31295;
  assign new_n31507 = new_n31506 ^ new_n31498;
  assign new_n31508 = new_n31507 ^ new_n31505;
  assign new_n31509 = new_n28439 ^ new_n27262;
  assign new_n31510 = new_n31509 ^ new_n28030;
  assign new_n31511 = new_n31510 ^ new_n30414;
  assign new_n31512 = new_n28234 ^ new_n27863;
  assign new_n31513 = new_n31512 ^ new_n28218;
  assign new_n31514 = new_n31513 ^ new_n31511;
  assign new_n31515 = new_n28458 ^ new_n27308;
  assign new_n31516 = new_n31515 ^ new_n30399;
  assign new_n31517 = new_n28189 ^ new_n28004;
  assign new_n31518 = new_n31517 ^ new_n31516;
  assign new_n31519 = new_n31518 ^ new_n31514;
  assign new_n31520 = new_n28465 ^ new_n27293;
  assign new_n31521 = new_n31520 ^ new_n28095;
  assign new_n31522 = new_n30375 ^ new_n28230;
  assign new_n31523 = new_n31522 ^ new_n31521;
  assign new_n31524 = new_n28192 ^ new_n27984;
  assign new_n31525 = new_n28468 ^ new_n27258;
  assign new_n31526 = new_n31525 ^ new_n28114;
  assign new_n31527 = new_n31526 ^ new_n28175;
  assign new_n31528 = new_n31527 ^ new_n31524;
  assign new_n31529 = new_n31528 ^ new_n31523;
  assign new_n31530 = new_n31529 ^ new_n31519;
  assign new_n31531 = new_n30414 ^ new_n28198;
  assign new_n31532 = new_n31531 ^ new_n28142;
  assign new_n31533 = new_n28479 ^ new_n27281;
  assign new_n31534 = new_n31533 ^ new_n28205;
  assign new_n31535 = new_n31534 ^ new_n28080;
  assign new_n31536 = new_n31535 ^ new_n31532;
  assign new_n31537 = new_n31536 ^ new_n31518;
  assign new_n31538 = new_n28484 ^ new_n27299;
  assign new_n31539 = new_n31538 ^ new_n28175;
  assign new_n31540 = new_n31539 ^ new_n28004;
  assign new_n31541 = new_n28126 ^ new_n28048;
  assign new_n31542 = new_n31541 ^ new_n31540;
  assign new_n31543 = new_n31542 ^ new_n31518;
  assign new_n31544 = new_n28488 ^ new_n27287;
  assign new_n31545 = new_n31544 ^ new_n28147;
  assign new_n31546 = new_n30414 ^ new_n28206;
  assign new_n31547 = new_n31546 ^ new_n31545;
  assign new_n31548 = new_n31547 ^ new_n31543;
  assign new_n31549 = ~new_n31536 & ~new_n31548;
  assign new_n31550 = new_n31549 ^ new_n31536;
  assign new_n31551 = new_n31548 ^ new_n31536;
  assign new_n31552 = new_n31551 ^ new_n31529;
  assign new_n31553 = new_n31528 ^ new_n31514;
  assign new_n31554 = new_n28499 ^ new_n27271;
  assign new_n31555 = new_n31554 ^ new_n30414;
  assign new_n31556 = new_n31555 ^ new_n27715;
  assign new_n31557 = new_n28218 ^ new_n28085;
  assign new_n31558 = new_n31557 ^ new_n28095;
  assign new_n31559 = new_n31558 ^ new_n31556;
  assign new_n31560 = new_n31559 ^ new_n31536;
  assign new_n31561 = new_n31560 ^ new_n31553;
  assign new_n31562 = new_n31561 ^ new_n31547;
  assign new_n31563 = ~new_n31562 & new_n31552;
  assign new_n31564 = new_n31563 ^ new_n31550;
  assign new_n31565 = new_n31536 ^ new_n31514;
  assign new_n31566 = new_n31565 ^ new_n31529;
  assign new_n31567 = ~new_n31561 & ~new_n31566;
  assign new_n31568 = new_n31567 ^ new_n31542;
  assign new_n31569 = ~new_n31543 & new_n31547;
  assign new_n31570 = ~new_n31514 & ~new_n31547;
  assign new_n31571 = new_n31570 ^ new_n31569;
  assign new_n31572 = new_n31571 ^ new_n31568;
  assign new_n31573 = new_n31528 ^ new_n31518;
  assign new_n31574 = new_n31561 ^ new_n31543;
  assign new_n31575 = ~new_n31574 & new_n31529;
  assign new_n31576 = new_n31523 ^ new_n31514;
  assign new_n31577 = ~new_n31530 & new_n31576;
  assign new_n31578 = new_n31577 ^ new_n31575;
  assign new_n31579 = new_n31571 ^ new_n31514;
  assign new_n31580 = new_n31579 ^ new_n31563;
  assign new_n31581 = new_n31580 ^ new_n31578;
  assign new_n31582 = new_n31581 ^ new_n31573;
  assign new_n31583 = new_n31560 ^ new_n31523;
  assign new_n31584 = new_n31583 ^ new_n31542;
  assign new_n31585 = new_n31553 & new_n31584;
  assign new_n31586 = new_n31585 ^ new_n31575;
  assign new_n31587 = new_n31583 ^ new_n31518;
  assign new_n31588 = new_n31587 ^ new_n31586;
  assign new_n31589 = new_n31536 ^ new_n31528;
  assign new_n31590 = ~new_n31589 & new_n31587;
  assign new_n31591 = new_n31548 ^ new_n31528;
  assign new_n31592 = new_n31584 ^ new_n31547;
  assign new_n31593 = ~new_n31591 & new_n31592;
  assign new_n31594 = new_n31593 ^ new_n31590;
  assign new_n31595 = new_n31594 ^ new_n31528;
  assign new_n31596 = new_n31595 ^ new_n31588;
  assign new_n31597 = new_n31590 ^ new_n31550;
  assign new_n31598 = new_n31597 ^ new_n31529;
  assign new_n31599 = new_n31585 ^ new_n31577;
  assign new_n31600 = new_n31559 ^ new_n31518;
  assign new_n31601 = new_n31600 ^ new_n31599;
  assign new_n31602 = new_n31601 ^ new_n31598;
  assign new_n31603 = new_n31568 ^ new_n31561;
  assign new_n31604 = new_n31563 ^ new_n31523;
  assign new_n31605 = new_n31604 ^ new_n31599;
  assign new_n31606 = new_n31605 ^ new_n31603;
  assign new_n31607 = new_n31602 & new_n31606;
  assign new_n31608 = new_n31607 ^ new_n31596;
  assign new_n31609 = ~new_n31608 & new_n31582;
  assign new_n31610 = new_n31609 ^ new_n31572;
  assign new_n31611 = new_n31610 ^ new_n31588;
  assign new_n31612 = new_n31607 ^ new_n31572;
  assign new_n31613 = new_n31612 ^ new_n31588;
  assign new_n31614 = new_n31593 ^ new_n31549;
  assign new_n31615 = new_n31614 ^ new_n31578;
  assign new_n31616 = ~new_n31615 & new_n31613;
  assign new_n31617 = new_n31616 ^ new_n31607;
  assign new_n31618 = ~new_n31596 & new_n31617;
  assign new_n31619 = new_n31618 ^ new_n31608;
  assign new_n31620 = ~new_n31619 & new_n31611;
  assign new_n31621 = new_n31620 ^ new_n31618;
  assign new_n31622 = new_n31621 ^ new_n31564;
  assign new_n31623 = new_n31622 ^ new_n31537;
  assign new_n31624 = new_n31623 ^ new_n31514;
  assign new_n31625 = new_n31609 ^ new_n31590;
  assign new_n31626 = new_n31625 ^ new_n31568;
  assign new_n31627 = new_n31626 ^ new_n31624;
  assign new_n31628 = ~new_n31530 & new_n31627;
  assign new_n31629 = new_n31616 ^ new_n31609;
  assign new_n31630 = new_n31595 ^ new_n31572;
  assign new_n31631 = new_n31630 ^ new_n31629;
  assign new_n31632 = ~new_n31631 & new_n31584;
  assign new_n31633 = new_n31632 ^ new_n31628;
  assign new_n31634 = new_n31618 ^ new_n31616;
  assign new_n31635 = new_n31634 ^ new_n31615;
  assign new_n31636 = ~new_n31562 & ~new_n31635;
  assign new_n31637 = new_n31618 ^ new_n31602;
  assign new_n31638 = ~new_n31561 & new_n31637;
  assign new_n31639 = new_n31638 ^ new_n31636;
  assign new_n31640 = ~new_n31566 & new_n31637;
  assign new_n31641 = new_n31640 ^ new_n31639;
  assign new_n31642 = ~new_n31635 & new_n31552;
  assign new_n31643 = new_n31576 & new_n31627;
  assign new_n31644 = ~new_n31631 & new_n31553;
  assign new_n31645 = new_n31644 ^ new_n31643;
  assign new_n31646 = new_n31645 ^ new_n31642;
  assign new_n31647 = new_n31646 ^ new_n31641;
  assign new_n31648 = new_n31647 ^ new_n31633;
  assign new_n31649 = new_n30261 ^ new_n26966;
  assign new_n31650 = new_n30680 ^ new_n26905;
  assign new_n31651 = new_n31650 ^ new_n27159;
  assign new_n31652 = new_n31651 ^ new_n31649;
  assign new_n31653 = new_n27121 ^ new_n26941;
  assign new_n31654 = new_n30681 ^ new_n30273;
  assign new_n31655 = new_n31654 ^ new_n31653;
  assign new_n31656 = new_n31655 ^ new_n31652;
  assign new_n31657 = new_n30683 ^ new_n27089;
  assign new_n31658 = new_n27031 ^ new_n27026;
  assign new_n31659 = new_n31658 ^ new_n27148;
  assign new_n31660 = new_n31659 ^ new_n31657;
  assign new_n31661 = new_n27124 ^ new_n26501;
  assign new_n31662 = new_n30684 ^ new_n27049;
  assign new_n31663 = new_n31662 ^ new_n27108;
  assign new_n31664 = new_n31663 ^ new_n31661;
  assign new_n31665 = new_n31664 ^ new_n31660;
  assign new_n31666 = new_n31665 ^ new_n31656;
  assign new_n31667 = new_n30261 ^ new_n27088;
  assign new_n31668 = new_n31667 ^ new_n27137;
  assign new_n31669 = new_n30687 ^ new_n27045;
  assign new_n31670 = new_n31669 ^ new_n27016;
  assign new_n31671 = new_n31670 ^ new_n31668;
  assign new_n31672 = new_n31671 ^ new_n31655;
  assign new_n31673 = new_n27060 ^ new_n26984;
  assign new_n31674 = new_n30689 ^ new_n27108;
  assign new_n31675 = new_n31674 ^ new_n26941;
  assign new_n31676 = new_n31675 ^ new_n31673;
  assign new_n31677 = new_n31676 ^ new_n31655;
  assign new_n31678 = new_n30261 ^ new_n27136;
  assign new_n31679 = new_n30691 ^ new_n27102;
  assign new_n31680 = new_n31679 ^ new_n27071;
  assign new_n31681 = new_n31680 ^ new_n31678;
  assign new_n31682 = new_n31681 ^ new_n31677;
  assign new_n31683 = new_n31671 & new_n31682;
  assign new_n31684 = new_n31683 ^ new_n31671;
  assign new_n31685 = new_n31682 ^ new_n31671;
  assign new_n31686 = new_n31685 ^ new_n31665;
  assign new_n31687 = new_n31664 ^ new_n31652;
  assign new_n31688 = new_n30698 ^ new_n30261;
  assign new_n31689 = new_n31688 ^ new_n27027;
  assign new_n31690 = new_n27158 ^ new_n26921;
  assign new_n31691 = new_n31690 ^ new_n31689;
  assign new_n31692 = new_n31691 ^ new_n31671;
  assign new_n31693 = new_n31692 ^ new_n31687;
  assign new_n31694 = new_n31693 ^ new_n31681;
  assign new_n31695 = new_n31686 & new_n31694;
  assign new_n31696 = new_n31695 ^ new_n31684;
  assign new_n31697 = new_n31671 ^ new_n31652;
  assign new_n31698 = new_n31697 ^ new_n31665;
  assign new_n31699 = ~new_n31693 & ~new_n31698;
  assign new_n31700 = new_n31699 ^ new_n31676;
  assign new_n31701 = ~new_n31677 & ~new_n31681;
  assign new_n31702 = new_n31652 & new_n31681;
  assign new_n31703 = new_n31702 ^ new_n31701;
  assign new_n31704 = new_n31703 ^ new_n31700;
  assign new_n31705 = new_n31664 ^ new_n31655;
  assign new_n31706 = new_n31693 ^ new_n31677;
  assign new_n31707 = ~new_n31706 & new_n31665;
  assign new_n31708 = new_n31660 ^ new_n31652;
  assign new_n31709 = ~new_n31666 & new_n31708;
  assign new_n31710 = new_n31709 ^ new_n31707;
  assign new_n31711 = new_n31703 ^ new_n31652;
  assign new_n31712 = new_n31711 ^ new_n31695;
  assign new_n31713 = new_n31712 ^ new_n31710;
  assign new_n31714 = new_n31713 ^ new_n31705;
  assign new_n31715 = new_n31692 ^ new_n31660;
  assign new_n31716 = new_n31715 ^ new_n31676;
  assign new_n31717 = new_n31687 & new_n31716;
  assign new_n31718 = new_n31717 ^ new_n31707;
  assign new_n31719 = new_n31715 ^ new_n31655;
  assign new_n31720 = new_n31719 ^ new_n31718;
  assign new_n31721 = new_n31671 ^ new_n31664;
  assign new_n31722 = ~new_n31721 & new_n31719;
  assign new_n31723 = new_n31682 ^ new_n31664;
  assign new_n31724 = new_n31716 ^ new_n31681;
  assign new_n31725 = ~new_n31723 & ~new_n31724;
  assign new_n31726 = new_n31725 ^ new_n31722;
  assign new_n31727 = new_n31726 ^ new_n31664;
  assign new_n31728 = new_n31727 ^ new_n31720;
  assign new_n31729 = new_n31722 ^ new_n31684;
  assign new_n31730 = new_n31729 ^ new_n31665;
  assign new_n31731 = new_n31717 ^ new_n31709;
  assign new_n31732 = new_n31691 ^ new_n31655;
  assign new_n31733 = new_n31732 ^ new_n31731;
  assign new_n31734 = new_n31733 ^ new_n31730;
  assign new_n31735 = new_n31700 ^ new_n31693;
  assign new_n31736 = new_n31731 ^ new_n31695;
  assign new_n31737 = new_n31736 ^ new_n31660;
  assign new_n31738 = new_n31737 ^ new_n31735;
  assign new_n31739 = ~new_n31734 & new_n31738;
  assign new_n31740 = new_n31739 ^ new_n31728;
  assign new_n31741 = ~new_n31714 & new_n31740;
  assign new_n31742 = new_n31741 ^ new_n31704;
  assign new_n31743 = new_n31742 ^ new_n31720;
  assign new_n31744 = new_n31739 ^ new_n31704;
  assign new_n31745 = new_n31744 ^ new_n31720;
  assign new_n31746 = new_n31725 ^ new_n31683;
  assign new_n31747 = new_n31746 ^ new_n31710;
  assign new_n31748 = ~new_n31745 & ~new_n31747;
  assign new_n31749 = new_n31748 ^ new_n31739;
  assign new_n31750 = new_n31728 & new_n31749;
  assign new_n31751 = new_n31750 ^ new_n31740;
  assign new_n31752 = ~new_n31743 & new_n31751;
  assign new_n31753 = new_n31752 ^ new_n31750;
  assign new_n31754 = new_n31753 ^ new_n31696;
  assign new_n31755 = new_n31754 ^ new_n31672;
  assign new_n31756 = new_n31755 ^ new_n31652;
  assign new_n31757 = new_n31741 ^ new_n31722;
  assign new_n31758 = new_n31757 ^ new_n31700;
  assign new_n31759 = new_n31758 ^ new_n31756;
  assign new_n31760 = ~new_n31666 & ~new_n31759;
  assign new_n31761 = new_n31748 ^ new_n31741;
  assign new_n31762 = new_n31727 ^ new_n31704;
  assign new_n31763 = new_n31762 ^ new_n31761;
  assign new_n31764 = ~new_n31763 & new_n31716;
  assign new_n31765 = new_n31764 ^ new_n31760;
  assign new_n31766 = new_n31750 ^ new_n31748;
  assign new_n31767 = new_n31766 ^ new_n31747;
  assign new_n31768 = ~new_n31767 & new_n31694;
  assign new_n31769 = new_n31750 ^ new_n31734;
  assign new_n31770 = ~new_n31693 & ~new_n31769;
  assign new_n31771 = new_n31770 ^ new_n31768;
  assign new_n31772 = ~new_n31698 & ~new_n31769;
  assign new_n31773 = new_n31772 ^ new_n31771;
  assign new_n31774 = ~new_n31767 & new_n31686;
  assign new_n31775 = ~new_n31759 & new_n31708;
  assign new_n31776 = ~new_n31763 & new_n31687;
  assign new_n31777 = new_n31776 ^ new_n31775;
  assign new_n31778 = new_n31777 ^ new_n31774;
  assign new_n31779 = new_n31778 ^ new_n31773;
  assign new_n31780 = new_n31779 ^ new_n31765;
  assign new_n31781 = new_n31780 ^ new_n31648;
  assign new_n31782 = new_n29254 ^ new_n29231;
  assign new_n31783 = new_n28178 ^ new_n24436;
  assign new_n31784 = new_n31783 ^ new_n16812;
  assign new_n31785 = new_n31784 ^ new_n29258;
  assign new_n31786 = new_n31785 ^ new_n29349;
  assign new_n31787 = new_n31786 ^ new_n31782;
  assign new_n31788 = new_n29379 ^ new_n29176;
  assign new_n31789 = new_n31788 ^ new_n29164;
  assign new_n31790 = new_n28222 ^ new_n24561;
  assign new_n31791 = new_n31790 ^ new_n16854;
  assign new_n31792 = new_n31791 ^ new_n29251;
  assign new_n31793 = new_n31792 ^ new_n29270;
  assign new_n31794 = new_n31793 ^ new_n31789;
  assign new_n31795 = new_n29277 ^ new_n29251;
  assign new_n31796 = new_n31795 ^ new_n29361;
  assign new_n31797 = new_n28158 ^ new_n24596;
  assign new_n31798 = new_n31797 ^ new_n16836;
  assign new_n31799 = new_n31798 ^ new_n29291;
  assign new_n31800 = new_n31799 ^ new_n29317;
  assign new_n31801 = new_n31800 ^ new_n31796;
  assign new_n31802 = new_n31801 ^ new_n31794;
  assign new_n31803 = new_n29296 ^ new_n29269;
  assign new_n31804 = new_n31803 ^ new_n29385;
  assign new_n31805 = new_n28100 ^ new_n24616;
  assign new_n31806 = new_n31805 ^ new_n16849;
  assign new_n31807 = new_n31806 ^ new_n29318;
  assign new_n31808 = new_n31807 ^ new_n31804;
  assign new_n31809 = new_n31808 ^ new_n31802;
  assign new_n31810 = new_n31809 ^ new_n31787;
  assign new_n31811 = new_n29320 ^ new_n29251;
  assign new_n31812 = new_n28200 ^ new_n24475;
  assign new_n31813 = new_n31812 ^ new_n16823;
  assign new_n31814 = new_n31813 ^ new_n29328;
  assign new_n31815 = new_n31814 ^ new_n29360;
  assign new_n31816 = new_n31815 ^ new_n31811;
  assign new_n31817 = new_n27966 ^ new_n24517;
  assign new_n31818 = new_n31817 ^ new_n16828;
  assign new_n31819 = new_n31818 ^ new_n29251;
  assign new_n31820 = new_n31819 ^ new_n29380;
  assign new_n31821 = new_n29239 ^ new_n28869;
  assign new_n31822 = new_n31821 ^ new_n31820;
  assign new_n31823 = new_n29194 ^ new_n28870;
  assign new_n31824 = new_n28022 ^ new_n24230;
  assign new_n31825 = new_n31824 ^ new_n16817;
  assign new_n31826 = new_n31825 ^ new_n29341;
  assign new_n31827 = new_n31826 ^ new_n29230;
  assign new_n31828 = new_n31827 ^ new_n31823;
  assign new_n31829 = new_n31828 ^ new_n31787;
  assign new_n31830 = new_n31829 ^ new_n31816;
  assign new_n31831 = new_n31830 ^ new_n31822;
  assign new_n31832 = ~new_n31816 & ~new_n31831;
  assign new_n31833 = new_n31832 ^ new_n31822;
  assign new_n31834 = new_n28116 ^ new_n24541;
  assign new_n31835 = new_n31834 ^ new_n16842;
  assign new_n31836 = new_n31835 ^ new_n29350;
  assign new_n31837 = new_n29250 ^ new_n29154;
  assign new_n31838 = new_n31837 ^ new_n29002;
  assign new_n31839 = new_n31838 ^ new_n31836;
  assign new_n31840 = new_n31839 ^ new_n31822;
  assign new_n31841 = new_n31840 ^ new_n31802;
  assign new_n31842 = new_n31839 ^ new_n31801;
  assign new_n31843 = new_n31822 ^ new_n31808;
  assign new_n31844 = new_n31843 ^ new_n31842;
  assign new_n31845 = ~new_n31841 & ~new_n31844;
  assign new_n31846 = new_n31845 ^ new_n31787;
  assign new_n31847 = new_n31846 ^ new_n31833;
  assign new_n31848 = new_n31801 & new_n31830;
  assign new_n31849 = new_n31848 ^ new_n31801;
  assign new_n31850 = new_n31828 ^ new_n31809;
  assign new_n31851 = ~new_n31842 & new_n31850;
  assign new_n31852 = new_n31851 ^ new_n31849;
  assign new_n31853 = new_n31839 ^ new_n31808;
  assign new_n31854 = new_n31853 ^ new_n31852;
  assign new_n31855 = new_n31810 & new_n31840;
  assign new_n31856 = new_n31828 ^ new_n31822;
  assign new_n31857 = new_n31856 ^ new_n31853;
  assign new_n31858 = ~new_n31857 & new_n31843;
  assign new_n31859 = new_n31858 ^ new_n31855;
  assign new_n31860 = new_n31828 ^ new_n31794;
  assign new_n31861 = new_n31860 ^ new_n31859;
  assign new_n31862 = new_n31861 ^ new_n31854;
  assign new_n31863 = new_n31846 ^ new_n31841;
  assign new_n31864 = new_n31830 ^ new_n31801;
  assign new_n31865 = new_n31864 ^ new_n31853;
  assign new_n31866 = new_n31841 ^ new_n31816;
  assign new_n31867 = new_n31865 & new_n31866;
  assign new_n31868 = new_n31867 ^ new_n31859;
  assign new_n31869 = new_n31868 ^ new_n31808;
  assign new_n31870 = new_n31869 ^ new_n31863;
  assign new_n31871 = ~new_n31862 & new_n31870;
  assign new_n31872 = new_n31871 ^ new_n31847;
  assign new_n31873 = new_n31841 ^ new_n31829;
  assign new_n31874 = ~new_n31873 & new_n31853;
  assign new_n31875 = new_n31874 ^ new_n31855;
  assign new_n31876 = new_n31875 ^ new_n31850;
  assign new_n31877 = new_n31876 ^ new_n31872;
  assign new_n31878 = new_n31839 ^ new_n31830;
  assign new_n31879 = new_n31816 ^ new_n31810;
  assign new_n31880 = ~new_n31878 & ~new_n31879;
  assign new_n31881 = new_n31880 ^ new_n31848;
  assign new_n31882 = new_n31874 ^ new_n31858;
  assign new_n31883 = new_n31882 ^ new_n31881;
  assign new_n31884 = ~new_n31877 & ~new_n31883;
  assign new_n31885 = new_n31839 ^ new_n31828;
  assign new_n31886 = new_n31867 ^ new_n31832;
  assign new_n31887 = new_n31886 ^ new_n31882;
  assign new_n31888 = new_n31887 ^ new_n31885;
  assign new_n31889 = new_n31880 ^ new_n31851;
  assign new_n31890 = new_n31889 ^ new_n31839;
  assign new_n31891 = new_n31890 ^ new_n31876;
  assign new_n31892 = new_n31891 ^ new_n31871;
  assign new_n31893 = ~new_n31888 & new_n31892;
  assign new_n31894 = new_n31893 ^ new_n31884;
  assign new_n31895 = new_n31890 ^ new_n31847;
  assign new_n31896 = new_n31895 ^ new_n31894;
  assign new_n31897 = ~new_n31896 & new_n31810;
  assign new_n31898 = ~new_n31896 & new_n31840;
  assign new_n31899 = new_n31898 ^ new_n31897;
  assign new_n31900 = new_n31884 ^ new_n31839;
  assign new_n31901 = new_n31880 ^ new_n31832;
  assign new_n31902 = new_n31828 ^ new_n31801;
  assign new_n31903 = new_n31867 ^ new_n31849;
  assign new_n31904 = new_n31893 ^ new_n31847;
  assign new_n31905 = new_n31904 ^ new_n31876;
  assign new_n31906 = new_n31884 ^ new_n31871;
  assign new_n31907 = new_n31891 & new_n31906;
  assign new_n31908 = new_n31907 ^ new_n31892;
  assign new_n31909 = ~new_n31905 & new_n31908;
  assign new_n31910 = new_n31909 ^ new_n31907;
  assign new_n31911 = new_n31910 ^ new_n31903;
  assign new_n31912 = new_n31911 ^ new_n31902;
  assign new_n31913 = new_n31912 ^ new_n31901;
  assign new_n31914 = new_n31913 ^ new_n31900;
  assign new_n31915 = new_n31853 & new_n31914;
  assign new_n31916 = ~new_n31878 & ~new_n31905;
  assign new_n31917 = ~new_n31873 & new_n31914;
  assign new_n31918 = new_n31917 ^ new_n31916;
  assign new_n31919 = new_n31891 ^ new_n31884;
  assign new_n31920 = ~new_n31816 & new_n31919;
  assign new_n31921 = new_n31907 ^ new_n31862;
  assign new_n31922 = ~new_n31841 & ~new_n31921;
  assign new_n31923 = new_n31922 ^ new_n31920;
  assign new_n31924 = new_n31909 ^ new_n31893;
  assign new_n31925 = new_n31924 ^ new_n31870;
  assign new_n31926 = ~new_n31842 & new_n31925;
  assign new_n31927 = new_n31926 ^ new_n31923;
  assign new_n31928 = new_n31927 ^ new_n31918;
  assign new_n31929 = new_n31928 ^ new_n31915;
  assign new_n31930 = new_n31929 ^ new_n31899;
  assign new_n31931 = new_n31930 ^ new_n31781;
  assign new_n31932 = new_n30270 ^ new_n30246;
  assign new_n31933 = new_n30259 ^ new_n30220;
  assign new_n31934 = new_n31933 ^ new_n31932;
  assign new_n31935 = new_n30246 ^ new_n30227;
  assign new_n31936 = new_n30246 ^ new_n30240;
  assign new_n31937 = new_n31936 ^ new_n30251;
  assign new_n31938 = ~new_n30227 & ~new_n31937;
  assign new_n31939 = new_n31938 ^ new_n30227;
  assign new_n31940 = new_n31937 ^ new_n30227;
  assign new_n31941 = new_n31940 ^ new_n31933;
  assign new_n31942 = new_n30270 ^ new_n30259;
  assign new_n31943 = new_n30232 ^ new_n30227;
  assign new_n31944 = new_n31943 ^ new_n31942;
  assign new_n31945 = new_n31944 ^ new_n30251;
  assign new_n31946 = new_n31941 & new_n31945;
  assign new_n31947 = new_n31946 ^ new_n31939;
  assign new_n31948 = new_n30270 ^ new_n30227;
  assign new_n31949 = new_n31948 ^ new_n31933;
  assign new_n31950 = new_n31944 & new_n31949;
  assign new_n31951 = new_n31950 ^ new_n30240;
  assign new_n31952 = ~new_n31936 & new_n30251;
  assign new_n31953 = ~new_n30251 & new_n30270;
  assign new_n31954 = new_n31953 ^ new_n31952;
  assign new_n31955 = new_n31954 ^ new_n31951;
  assign new_n31956 = new_n30259 ^ new_n30246;
  assign new_n31957 = new_n31944 ^ new_n31936;
  assign new_n31958 = new_n31933 & new_n31957;
  assign new_n31959 = new_n30270 ^ new_n30220;
  assign new_n31960 = new_n31934 & new_n31959;
  assign new_n31961 = new_n31960 ^ new_n31958;
  assign new_n31962 = new_n31954 ^ new_n30270;
  assign new_n31963 = new_n31962 ^ new_n31946;
  assign new_n31964 = new_n31963 ^ new_n31961;
  assign new_n31965 = new_n31964 ^ new_n31956;
  assign new_n31966 = new_n30232 ^ new_n30220;
  assign new_n31967 = new_n31966 ^ new_n30227;
  assign new_n31968 = new_n31967 ^ new_n30240;
  assign new_n31969 = new_n31942 & new_n31968;
  assign new_n31970 = new_n31969 ^ new_n31958;
  assign new_n31971 = new_n31967 ^ new_n30246;
  assign new_n31972 = new_n31971 ^ new_n31970;
  assign new_n31973 = new_n30259 ^ new_n30227;
  assign new_n31974 = new_n31971 & new_n31973;
  assign new_n31975 = new_n31937 ^ new_n30259;
  assign new_n31976 = new_n31968 ^ new_n30251;
  assign new_n31977 = new_n31975 & new_n31976;
  assign new_n31978 = new_n31977 ^ new_n31974;
  assign new_n31979 = new_n31978 ^ new_n30259;
  assign new_n31980 = new_n31979 ^ new_n31972;
  assign new_n31981 = new_n31974 ^ new_n31939;
  assign new_n31982 = new_n31981 ^ new_n31933;
  assign new_n31983 = new_n31969 ^ new_n31960;
  assign new_n31984 = new_n30246 ^ new_n30232;
  assign new_n31985 = new_n31984 ^ new_n31983;
  assign new_n31986 = new_n31985 ^ new_n31982;
  assign new_n31987 = new_n31951 ^ new_n31944;
  assign new_n31988 = new_n31969 ^ new_n31946;
  assign new_n31989 = new_n31960 ^ new_n30220;
  assign new_n31990 = new_n31989 ^ new_n31988;
  assign new_n31991 = new_n31990 ^ new_n31987;
  assign new_n31992 = ~new_n31986 & new_n31991;
  assign new_n31993 = new_n31992 ^ new_n31980;
  assign new_n31994 = new_n31965 & new_n31993;
  assign new_n31995 = new_n31994 ^ new_n31955;
  assign new_n31996 = new_n31995 ^ new_n31972;
  assign new_n31997 = new_n31992 ^ new_n31955;
  assign new_n31998 = new_n31997 ^ new_n31972;
  assign new_n31999 = new_n31977 ^ new_n31938;
  assign new_n32000 = new_n31999 ^ new_n31961;
  assign new_n32001 = ~new_n32000 & new_n31998;
  assign new_n32002 = new_n32001 ^ new_n31992;
  assign new_n32003 = new_n31980 & new_n32002;
  assign new_n32004 = new_n32003 ^ new_n31993;
  assign new_n32005 = new_n31996 & new_n32004;
  assign new_n32006 = new_n32005 ^ new_n32003;
  assign new_n32007 = new_n32006 ^ new_n31947;
  assign new_n32008 = new_n32007 ^ new_n31935;
  assign new_n32009 = new_n32008 ^ new_n30270;
  assign new_n32010 = new_n31994 ^ new_n31974;
  assign new_n32011 = new_n32010 ^ new_n31951;
  assign new_n32012 = new_n32011 ^ new_n32009;
  assign new_n32013 = ~new_n32012 & new_n31934;
  assign new_n32014 = new_n32001 ^ new_n31994;
  assign new_n32015 = new_n31979 ^ new_n31955;
  assign new_n32016 = new_n32015 ^ new_n32014;
  assign new_n32017 = new_n31968 & new_n32016;
  assign new_n32018 = new_n32017 ^ new_n32013;
  assign new_n32019 = new_n32003 ^ new_n32001;
  assign new_n32020 = new_n32019 ^ new_n32000;
  assign new_n32021 = ~new_n32020 & new_n31945;
  assign new_n32022 = new_n32003 ^ new_n31986;
  assign new_n32023 = ~new_n32022 & new_n31944;
  assign new_n32024 = new_n32023 ^ new_n32021;
  assign new_n32025 = ~new_n32022 & new_n31949;
  assign new_n32026 = new_n32025 ^ new_n32024;
  assign new_n32027 = ~new_n32020 & new_n31941;
  assign new_n32028 = ~new_n32012 & new_n31959;
  assign new_n32029 = new_n31942 & new_n32016;
  assign new_n32030 = new_n32029 ^ new_n32028;
  assign new_n32031 = new_n32030 ^ new_n32027;
  assign new_n32032 = new_n32031 ^ new_n32026;
  assign new_n32033 = new_n32032 ^ new_n32018;
  assign new_n32034 = new_n27111 ^ new_n26230;
  assign new_n32035 = new_n32034 ^ new_n32033;
  assign new_n32036 = new_n27036 ^ new_n19879;
  assign new_n32037 = new_n32036 ^ new_n25905;
  assign new_n32038 = new_n30543 ^ new_n25959;
  assign new_n32039 = new_n32038 ^ new_n32037;
  assign new_n32040 = new_n30557 ^ new_n26083;
  assign new_n32041 = new_n27098 ^ new_n19819;
  assign new_n32042 = new_n32041 ^ new_n25914;
  assign new_n32043 = new_n32042 ^ new_n26097;
  assign new_n32044 = new_n32043 ^ new_n32040;
  assign new_n32045 = new_n27163 ^ new_n19835;
  assign new_n32046 = new_n32045 ^ new_n25985;
  assign new_n32047 = new_n32046 ^ new_n26097;
  assign new_n32048 = new_n30584 ^ new_n24739;
  assign new_n32049 = new_n32048 ^ new_n32047;
  assign new_n32050 = new_n32049 ^ new_n32044;
  assign new_n32051 = new_n32050 ^ new_n32039;
  assign new_n32052 = new_n27111 ^ new_n19030;
  assign new_n32053 = new_n32052 ^ new_n26042;
  assign new_n32054 = new_n30565 ^ new_n26059;
  assign new_n32055 = new_n32054 ^ new_n32053;
  assign new_n32056 = new_n32055 ^ new_n32051;
  assign new_n32057 = new_n26959 ^ new_n19653;
  assign new_n32058 = new_n32057 ^ new_n26047;
  assign new_n32059 = new_n30539 ^ new_n26114;
  assign new_n32060 = new_n32059 ^ new_n32058;
  assign new_n32061 = new_n32060 ^ new_n32055;
  assign new_n32062 = new_n27130 ^ new_n19862;
  assign new_n32063 = new_n32062 ^ new_n25972;
  assign new_n32064 = new_n30574 ^ new_n26097;
  assign new_n32065 = new_n32064 ^ new_n32063;
  assign new_n32066 = new_n32065 ^ new_n32061;
  assign new_n32067 = new_n32044 & new_n32066;
  assign new_n32068 = new_n32067 ^ new_n32044;
  assign new_n32069 = new_n32060 ^ new_n32051;
  assign new_n32070 = new_n27051 ^ new_n19732;
  assign new_n32071 = new_n32070 ^ new_n25929;
  assign new_n32072 = new_n30549 ^ new_n26029;
  assign new_n32073 = new_n32072 ^ new_n32071;
  assign new_n32074 = new_n32073 ^ new_n32044;
  assign new_n32075 = ~new_n32074 & new_n32069;
  assign new_n32076 = new_n32075 ^ new_n32068;
  assign new_n32077 = new_n32073 ^ new_n32039;
  assign new_n32078 = new_n32077 ^ new_n32076;
  assign new_n32079 = new_n30529 ^ new_n26000;
  assign new_n32080 = new_n26604 ^ new_n19776;
  assign new_n32081 = new_n32080 ^ new_n26070;
  assign new_n32082 = new_n32081 ^ new_n26097;
  assign new_n32083 = new_n32082 ^ new_n32079;
  assign new_n32084 = new_n32083 ^ new_n32060;
  assign new_n32085 = new_n32084 ^ new_n32077;
  assign new_n32086 = new_n32083 ^ new_n32039;
  assign new_n32087 = ~new_n32085 & new_n32086;
  assign new_n32088 = new_n32083 ^ new_n32073;
  assign new_n32089 = new_n32056 & new_n32088;
  assign new_n32090 = new_n32089 ^ new_n32087;
  assign new_n32091 = new_n32060 ^ new_n32049;
  assign new_n32092 = new_n32091 ^ new_n32090;
  assign new_n32093 = new_n32092 ^ new_n32078;
  assign new_n32094 = new_n32088 ^ new_n32050;
  assign new_n32095 = new_n32083 ^ new_n32044;
  assign new_n32096 = new_n32095 ^ new_n32077;
  assign new_n32097 = ~new_n32094 & ~new_n32096;
  assign new_n32098 = new_n32097 ^ new_n32055;
  assign new_n32099 = new_n32098 ^ new_n32094;
  assign new_n32100 = new_n32094 ^ new_n32065;
  assign new_n32101 = new_n32066 ^ new_n32044;
  assign new_n32102 = new_n32101 ^ new_n32077;
  assign new_n32103 = new_n32100 & new_n32102;
  assign new_n32104 = new_n32103 ^ new_n32090;
  assign new_n32105 = new_n32104 ^ new_n32039;
  assign new_n32106 = new_n32105 ^ new_n32099;
  assign new_n32107 = ~new_n32093 & new_n32106;
  assign new_n32108 = new_n32094 ^ new_n32061;
  assign new_n32109 = ~new_n32108 & new_n32077;
  assign new_n32110 = new_n32109 ^ new_n32089;
  assign new_n32111 = new_n32110 ^ new_n32069;
  assign new_n32112 = new_n32073 ^ new_n32066;
  assign new_n32113 = new_n32065 ^ new_n32056;
  assign new_n32114 = ~new_n32112 & ~new_n32113;
  assign new_n32115 = new_n32114 ^ new_n32075;
  assign new_n32116 = new_n32115 ^ new_n32073;
  assign new_n32117 = new_n32116 ^ new_n32111;
  assign new_n32118 = new_n32117 ^ new_n32107;
  assign new_n32119 = new_n32073 ^ new_n32060;
  assign new_n32120 = new_n32083 ^ new_n32066;
  assign new_n32121 = ~new_n32065 & ~new_n32120;
  assign new_n32122 = new_n32121 ^ new_n32103;
  assign new_n32123 = new_n32109 ^ new_n32087;
  assign new_n32124 = new_n32123 ^ new_n32122;
  assign new_n32125 = new_n32124 ^ new_n32119;
  assign new_n32126 = ~new_n32125 & new_n32118;
  assign new_n32127 = new_n32121 ^ new_n32083;
  assign new_n32128 = new_n32127 ^ new_n32098;
  assign new_n32129 = new_n32128 ^ new_n32107;
  assign new_n32130 = new_n32129 ^ new_n32111;
  assign new_n32131 = new_n32114 ^ new_n32067;
  assign new_n32132 = new_n32131 ^ new_n32123;
  assign new_n32133 = ~new_n32130 & ~new_n32132;
  assign new_n32134 = new_n32133 ^ new_n32126;
  assign new_n32135 = new_n32128 ^ new_n32116;
  assign new_n32136 = new_n32135 ^ new_n32134;
  assign new_n32137 = ~new_n32136 & new_n32056;
  assign new_n32138 = ~new_n32136 & new_n32088;
  assign new_n32139 = new_n32138 ^ new_n32137;
  assign new_n32140 = new_n32133 ^ new_n32073;
  assign new_n32141 = new_n32121 ^ new_n32114;
  assign new_n32142 = new_n32060 ^ new_n32044;
  assign new_n32143 = new_n32103 ^ new_n32068;
  assign new_n32144 = new_n32128 ^ new_n32126;
  assign new_n32145 = new_n32144 ^ new_n32111;
  assign new_n32146 = new_n32133 ^ new_n32107;
  assign new_n32147 = ~new_n32146 & new_n32117;
  assign new_n32148 = new_n32147 ^ new_n32107;
  assign new_n32149 = ~new_n32145 & new_n32148;
  assign new_n32150 = new_n32147 ^ new_n32117;
  assign new_n32151 = new_n32150 ^ new_n32149;
  assign new_n32152 = new_n32151 ^ new_n32143;
  assign new_n32153 = new_n32152 ^ new_n32142;
  assign new_n32154 = new_n32153 ^ new_n32141;
  assign new_n32155 = new_n32154 ^ new_n32140;
  assign new_n32156 = new_n32077 & new_n32155;
  assign new_n32157 = ~new_n32112 & ~new_n32145;
  assign new_n32158 = ~new_n32108 & new_n32155;
  assign new_n32159 = new_n32158 ^ new_n32157;
  assign new_n32160 = new_n32149 ^ new_n32126;
  assign new_n32161 = new_n32160 ^ new_n32106;
  assign new_n32162 = ~new_n32074 & new_n32161;
  assign new_n32163 = new_n32133 ^ new_n32117;
  assign new_n32164 = ~new_n32065 & new_n32163;
  assign new_n32165 = new_n32150 ^ new_n32093;
  assign new_n32166 = ~new_n32094 & ~new_n32165;
  assign new_n32167 = new_n32166 ^ new_n32164;
  assign new_n32168 = new_n32167 ^ new_n32162;
  assign new_n32169 = new_n32168 ^ new_n32159;
  assign new_n32170 = new_n32169 ^ new_n32156;
  assign new_n32171 = new_n32170 ^ new_n32139;
  assign new_n32172 = new_n32171 ^ new_n32035;
  assign new_n32173 = new_n31912 ^ new_n31822;
  assign new_n32174 = new_n31893 ^ new_n31851;
  assign new_n32175 = new_n32174 ^ new_n31846;
  assign new_n32176 = new_n32175 ^ new_n32173;
  assign new_n32177 = ~new_n31857 & ~new_n32176;
  assign new_n32178 = new_n32177 ^ new_n31897;
  assign new_n32179 = new_n31907 ^ new_n31884;
  assign new_n32180 = new_n32179 ^ new_n31883;
  assign new_n32181 = ~new_n32180 & new_n31866;
  assign new_n32182 = new_n32181 ^ new_n31922;
  assign new_n32183 = ~new_n31844 & ~new_n31921;
  assign new_n32184 = new_n32183 ^ new_n32182;
  assign new_n32185 = ~new_n32180 & new_n31865;
  assign new_n32186 = ~new_n32176 & new_n31843;
  assign new_n32187 = new_n32186 ^ new_n31898;
  assign new_n32188 = new_n32187 ^ new_n32185;
  assign new_n32189 = new_n32188 ^ new_n32184;
  assign new_n32190 = new_n32189 ^ new_n32178;
  assign new_n32191 = new_n32190 ^ new_n32172;
  assign new_n32192 = new_n32191 ^ new_n31931;
  assign new_n32193 = new_n31748 ^ new_n31728;
  assign new_n32194 = new_n31682 ^ new_n31652;
  assign new_n32195 = ~new_n32194 & new_n32193;
  assign new_n32196 = new_n31752 ^ new_n31741;
  assign new_n32197 = new_n32196 ^ new_n31738;
  assign new_n32198 = new_n31719 & new_n32197;
  assign new_n32199 = new_n31752 ^ new_n31714;
  assign new_n32200 = ~new_n31682 & ~new_n32199;
  assign new_n32201 = new_n32200 ^ new_n31778;
  assign new_n32202 = new_n32201 ^ new_n32198;
  assign new_n32203 = new_n32202 ^ new_n31760;
  assign new_n32204 = new_n32203 ^ new_n32195;
  assign new_n32205 = ~new_n31681 & new_n32193;
  assign new_n32206 = new_n32205 ^ new_n31770;
  assign new_n32207 = ~new_n31721 & new_n32197;
  assign new_n32208 = new_n32207 ^ new_n32206;
  assign new_n32209 = ~new_n31723 & ~new_n31743;
  assign new_n32210 = new_n31748 ^ new_n31664;
  assign new_n32211 = new_n31725 ^ new_n31711;
  assign new_n32212 = new_n32211 ^ new_n31755;
  assign new_n32213 = new_n32212 ^ new_n32210;
  assign new_n32214 = ~new_n31706 & new_n32213;
  assign new_n32215 = new_n32214 ^ new_n32209;
  assign new_n32216 = new_n32215 ^ new_n32208;
  assign new_n32217 = new_n32216 ^ new_n32204;
  assign new_n32218 = new_n31616 ^ new_n31596;
  assign new_n32219 = new_n31548 ^ new_n31514;
  assign new_n32220 = ~new_n32218 & ~new_n32219;
  assign new_n32221 = new_n31620 ^ new_n31609;
  assign new_n32222 = new_n32221 ^ new_n31606;
  assign new_n32223 = new_n31587 & new_n32222;
  assign new_n32224 = new_n31620 ^ new_n31582;
  assign new_n32225 = new_n31548 & new_n32224;
  assign new_n32226 = new_n32225 ^ new_n31646;
  assign new_n32227 = new_n32226 ^ new_n32223;
  assign new_n32228 = new_n32227 ^ new_n31628;
  assign new_n32229 = new_n32228 ^ new_n32220;
  assign new_n32230 = ~new_n32218 & new_n31547;
  assign new_n32231 = new_n32230 ^ new_n31638;
  assign new_n32232 = ~new_n31589 & new_n32222;
  assign new_n32233 = new_n32232 ^ new_n32231;
  assign new_n32234 = ~new_n31591 & new_n31611;
  assign new_n32235 = new_n31616 ^ new_n31528;
  assign new_n32236 = new_n31593 ^ new_n31579;
  assign new_n32237 = new_n32236 ^ new_n31623;
  assign new_n32238 = new_n32237 ^ new_n32235;
  assign new_n32239 = ~new_n31574 & ~new_n32238;
  assign new_n32240 = new_n32239 ^ new_n32234;
  assign new_n32241 = new_n32240 ^ new_n32233;
  assign new_n32242 = new_n32241 ^ new_n32229;
  assign new_n32243 = new_n32242 ^ new_n32217;
  assign new_n32244 = new_n31926 ^ new_n31917;
  assign new_n32245 = ~new_n31879 & ~new_n31905;
  assign new_n32246 = new_n31909 ^ new_n31888;
  assign new_n32247 = ~new_n32246 & new_n31864;
  assign new_n32248 = new_n32247 ^ new_n32245;
  assign new_n32249 = new_n32248 ^ new_n32187;
  assign new_n32250 = ~new_n31830 & ~new_n32246;
  assign new_n32251 = new_n32250 ^ new_n32177;
  assign new_n32252 = new_n32251 ^ new_n32249;
  assign new_n32253 = new_n32252 ^ new_n32244;
  assign new_n32254 = new_n32253 ^ new_n32243;
  assign new_n32255 = new_n32162 ^ new_n32158;
  assign new_n32256 = new_n32153 ^ new_n32083;
  assign new_n32257 = new_n32126 ^ new_n32075;
  assign new_n32258 = new_n32257 ^ new_n32098;
  assign new_n32259 = new_n32258 ^ new_n32256;
  assign new_n32260 = ~new_n32085 & ~new_n32259;
  assign new_n32261 = new_n32149 ^ new_n32125;
  assign new_n32262 = ~new_n32066 & ~new_n32261;
  assign new_n32263 = new_n32262 ^ new_n32260;
  assign new_n32264 = ~new_n32113 & ~new_n32145;
  assign new_n32265 = ~new_n32261 & new_n32101;
  assign new_n32266 = new_n32265 ^ new_n32264;
  assign new_n32267 = ~new_n32259 & new_n32086;
  assign new_n32268 = new_n32267 ^ new_n32138;
  assign new_n32269 = new_n32268 ^ new_n32266;
  assign new_n32270 = new_n32269 ^ new_n32263;
  assign new_n32271 = new_n32270 ^ new_n32255;
  assign new_n32272 = new_n32001 ^ new_n31980;
  assign new_n32273 = new_n31937 ^ new_n30270;
  assign new_n32274 = new_n32272 & new_n32273;
  assign new_n32275 = new_n32005 ^ new_n31994;
  assign new_n32276 = new_n32275 ^ new_n31991;
  assign new_n32277 = new_n31971 & new_n32276;
  assign new_n32278 = new_n32005 ^ new_n31965;
  assign new_n32279 = new_n31937 & new_n32278;
  assign new_n32280 = new_n32279 ^ new_n32031;
  assign new_n32281 = new_n32280 ^ new_n32277;
  assign new_n32282 = new_n32281 ^ new_n32013;
  assign new_n32283 = new_n32282 ^ new_n32274;
  assign new_n32284 = new_n30251 & new_n32272;
  assign new_n32285 = new_n32284 ^ new_n32023;
  assign new_n32286 = new_n31973 & new_n32276;
  assign new_n32287 = new_n32286 ^ new_n32285;
  assign new_n32288 = new_n31975 & new_n31996;
  assign new_n32289 = new_n32001 ^ new_n30259;
  assign new_n32290 = new_n31977 ^ new_n31962;
  assign new_n32291 = new_n32290 ^ new_n32008;
  assign new_n32292 = new_n32291 ^ new_n32289;
  assign new_n32293 = ~new_n32292 & new_n31957;
  assign new_n32294 = new_n32293 ^ new_n32288;
  assign new_n32295 = new_n32294 ^ new_n32287;
  assign new_n32296 = new_n32295 ^ new_n32283;
  assign new_n32297 = new_n27036 ^ new_n26211;
  assign new_n32298 = new_n32297 ^ new_n32296;
  assign new_n32299 = ~new_n31831 & new_n31919;
  assign new_n32300 = new_n32250 ^ new_n32188;
  assign new_n32301 = new_n31850 & new_n31925;
  assign new_n32302 = new_n32301 ^ new_n32300;
  assign new_n32303 = new_n32302 ^ new_n32177;
  assign new_n32304 = new_n32303 ^ new_n32299;
  assign new_n32305 = new_n32304 ^ new_n31928;
  assign new_n32306 = new_n32305 ^ new_n32298;
  assign new_n32307 = new_n32306 ^ new_n32271;
  assign new_n32308 = new_n32307 ^ new_n32254;
  assign new_n32309 = ~new_n32120 & new_n32163;
  assign new_n32310 = new_n32150 ^ new_n32133;
  assign new_n32311 = new_n32310 ^ new_n32132;
  assign new_n32312 = ~new_n32311 & new_n32102;
  assign new_n32313 = new_n32312 ^ new_n32268;
  assign new_n32314 = new_n32313 ^ new_n32262;
  assign new_n32315 = new_n32069 & new_n32161;
  assign new_n32316 = new_n32315 ^ new_n32314;
  assign new_n32317 = new_n32316 ^ new_n32260;
  assign new_n32318 = new_n32317 ^ new_n32309;
  assign new_n32319 = new_n32318 ^ new_n32169;
  assign new_n32320 = new_n32245 ^ new_n32183;
  assign new_n32321 = new_n32181 ^ new_n31920;
  assign new_n32322 = new_n32321 ^ new_n32300;
  assign new_n32323 = new_n32322 ^ new_n32320;
  assign new_n32324 = new_n32323 ^ new_n32305;
  assign new_n32325 = new_n32324 ^ new_n32319;
  assign new_n32326 = ~new_n31724 & ~new_n31743;
  assign new_n32327 = new_n32326 ^ new_n31772;
  assign new_n32328 = new_n32205 ^ new_n31768;
  assign new_n32329 = new_n32328 ^ new_n32201;
  assign new_n32330 = new_n32329 ^ new_n32327;
  assign new_n32331 = new_n31592 & new_n31611;
  assign new_n32332 = new_n32331 ^ new_n31640;
  assign new_n32333 = new_n32230 ^ new_n31636;
  assign new_n32334 = new_n32333 ^ new_n32226;
  assign new_n32335 = new_n32334 ^ new_n32332;
  assign new_n32336 = new_n32335 ^ new_n32330;
  assign new_n32337 = new_n31976 & new_n31996;
  assign new_n32338 = new_n32337 ^ new_n32025;
  assign new_n32339 = new_n32284 ^ new_n32021;
  assign new_n32340 = new_n32339 ^ new_n32280;
  assign new_n32341 = new_n32340 ^ new_n32338;
  assign new_n32342 = new_n27163 ^ new_n26223;
  assign new_n32343 = new_n32342 ^ new_n32341;
  assign new_n32344 = ~new_n32096 & ~new_n32165;
  assign new_n32345 = new_n32344 ^ new_n32137;
  assign new_n32346 = new_n32345 ^ new_n32317;
  assign new_n32347 = new_n32183 ^ new_n31897;
  assign new_n32348 = new_n32347 ^ new_n32303;
  assign new_n32349 = new_n32348 ^ new_n32346;
  assign new_n32350 = new_n32349 ^ new_n32343;
  assign new_n32351 = new_n32350 ^ new_n32336;
  assign new_n32352 = new_n32351 ^ new_n32325;
  assign new_n32353 = new_n32239 ^ new_n32232;
  assign new_n32354 = new_n31551 & new_n32224;
  assign new_n32355 = new_n32354 ^ new_n32331;
  assign new_n32356 = new_n32355 ^ new_n31645;
  assign new_n32357 = new_n32225 ^ new_n31628;
  assign new_n32358 = new_n32357 ^ new_n32356;
  assign new_n32359 = new_n32358 ^ new_n32353;
  assign new_n32360 = new_n32214 ^ new_n32207;
  assign new_n32361 = ~new_n32199 & new_n31685;
  assign new_n32362 = new_n32361 ^ new_n32326;
  assign new_n32363 = new_n32362 ^ new_n31777;
  assign new_n32364 = new_n32200 ^ new_n31760;
  assign new_n32365 = new_n32364 ^ new_n32363;
  assign new_n32366 = new_n32365 ^ new_n32360;
  assign new_n32367 = new_n32366 ^ new_n32359;
  assign new_n32368 = new_n32367 ^ new_n32349;
  assign new_n32369 = new_n32301 ^ new_n31927;
  assign new_n32370 = new_n32369 ^ new_n32249;
  assign new_n32371 = new_n32315 ^ new_n32168;
  assign new_n32372 = new_n32371 ^ new_n32269;
  assign new_n32373 = new_n32372 ^ new_n32370;
  assign new_n32374 = new_n32293 ^ new_n32286;
  assign new_n32375 = new_n31940 & new_n32278;
  assign new_n32376 = new_n32375 ^ new_n32337;
  assign new_n32377 = new_n32376 ^ new_n32030;
  assign new_n32378 = new_n32279 ^ new_n32013;
  assign new_n32379 = new_n32378 ^ new_n32377;
  assign new_n32380 = new_n32379 ^ new_n32374;
  assign new_n32381 = new_n27098 ^ new_n26217;
  assign new_n32382 = new_n32381 ^ new_n32380;
  assign new_n32383 = new_n32382 ^ new_n32253;
  assign new_n32384 = new_n32383 ^ new_n32373;
  assign new_n32385 = new_n32384 ^ new_n32368;
  assign new_n32386 = new_n32385 ^ new_n32352;
  assign new_n32387 = new_n32386 ^ new_n32308;
  assign new_n32388 = new_n32387 ^ new_n32192;
  assign new_n32389 = new_n32233 ^ new_n32223;
  assign new_n32390 = new_n32389 ^ new_n32356;
  assign new_n32391 = new_n32287 ^ new_n32277;
  assign new_n32392 = new_n32391 ^ new_n32377;
  assign new_n32393 = new_n27130 ^ new_n26261;
  assign new_n32394 = new_n32393 ^ new_n32392;
  assign new_n32395 = new_n32394 ^ new_n32390;
  assign new_n32396 = new_n32208 ^ new_n32198;
  assign new_n32397 = new_n32396 ^ new_n32363;
  assign new_n32398 = new_n32397 ^ new_n32370;
  assign new_n32399 = new_n32398 ^ new_n32349;
  assign new_n32400 = new_n32399 ^ new_n32395;
  assign new_n32401 = new_n32202 ^ new_n31773;
  assign new_n32402 = new_n32227 ^ new_n31641;
  assign new_n32403 = new_n32402 ^ new_n32401;
  assign new_n32404 = new_n32281 ^ new_n32026;
  assign new_n32405 = new_n26604 ^ new_n26247;
  assign new_n32406 = new_n32405 ^ new_n32404;
  assign new_n32407 = new_n32406 ^ new_n32349;
  assign new_n32408 = new_n32407 ^ new_n32403;
  assign new_n32409 = new_n32344 ^ new_n32264;
  assign new_n32410 = ~new_n32311 & new_n32100;
  assign new_n32411 = new_n32410 ^ new_n32164;
  assign new_n32412 = new_n32411 ^ new_n32314;
  assign new_n32413 = new_n32412 ^ new_n32409;
  assign new_n32414 = new_n32302 ^ new_n32184;
  assign new_n32415 = new_n32414 ^ new_n32323;
  assign new_n32416 = new_n32415 ^ new_n32413;
  assign new_n32417 = new_n32416 ^ new_n32408;
  assign new_n32418 = new_n31644 ^ new_n31632;
  assign new_n32419 = ~new_n32238 & new_n31529;
  assign new_n32420 = new_n32419 ^ new_n32241;
  assign new_n32421 = new_n32420 ^ new_n32418;
  assign new_n32422 = new_n31776 ^ new_n31764;
  assign new_n32423 = new_n31665 & new_n32213;
  assign new_n32424 = new_n32423 ^ new_n32216;
  assign new_n32425 = new_n32424 ^ new_n32422;
  assign new_n32426 = new_n32425 ^ new_n32421;
  assign new_n32427 = new_n32426 ^ new_n31930;
  assign new_n32428 = new_n32029 ^ new_n32017;
  assign new_n32429 = ~new_n32292 & new_n31933;
  assign new_n32430 = new_n32429 ^ new_n32295;
  assign new_n32431 = new_n32430 ^ new_n32428;
  assign new_n32432 = new_n26959 ^ new_n26242;
  assign new_n32433 = new_n32432 ^ new_n32431;
  assign new_n32434 = new_n32410 ^ new_n32166;
  assign new_n32435 = new_n32434 ^ new_n32344;
  assign new_n32436 = new_n32435 ^ new_n32316;
  assign new_n32437 = new_n32436 ^ new_n32414;
  assign new_n32438 = new_n32437 ^ new_n32433;
  assign new_n32439 = new_n32438 ^ new_n32427;
  assign new_n32440 = new_n32439 ^ new_n32192;
  assign new_n32441 = new_n32440 ^ new_n32400;
  assign new_n32442 = new_n32441 ^ new_n32417;
  assign new_n32443 = new_n32400 & new_n32442;
  assign new_n32444 = new_n32443 ^ new_n32417;
  assign new_n32445 = new_n31772 ^ new_n31764;
  assign new_n32446 = new_n32445 ^ new_n32203;
  assign new_n32447 = new_n31640 ^ new_n31632;
  assign new_n32448 = new_n32447 ^ new_n32228;
  assign new_n32449 = new_n32448 ^ new_n32446;
  assign new_n32450 = new_n32449 ^ new_n32190;
  assign new_n32451 = new_n32260 ^ new_n32137;
  assign new_n32452 = new_n32435 ^ new_n32313;
  assign new_n32453 = new_n32452 ^ new_n32451;
  assign new_n32454 = new_n32025 ^ new_n32017;
  assign new_n32455 = new_n32454 ^ new_n32282;
  assign new_n32456 = new_n27051 ^ new_n26236;
  assign new_n32457 = new_n32456 ^ new_n32455;
  assign new_n32458 = new_n32457 ^ new_n32348;
  assign new_n32459 = new_n32458 ^ new_n32453;
  assign new_n32460 = new_n32459 ^ new_n32450;
  assign new_n32461 = new_n32460 ^ new_n32417;
  assign new_n32462 = new_n32461 ^ new_n32386;
  assign new_n32463 = new_n32417 ^ new_n32385;
  assign new_n32464 = new_n32460 ^ new_n32308;
  assign new_n32465 = new_n32464 ^ new_n32463;
  assign new_n32466 = new_n32462 & new_n32465;
  assign new_n32467 = new_n32466 ^ new_n32192;
  assign new_n32468 = new_n32467 ^ new_n32444;
  assign new_n32469 = ~new_n32385 & ~new_n32441;
  assign new_n32470 = new_n32469 ^ new_n32385;
  assign new_n32471 = new_n32439 ^ new_n32387;
  assign new_n32472 = new_n32460 ^ new_n32385;
  assign new_n32473 = new_n32471 & new_n32472;
  assign new_n32474 = new_n32473 ^ new_n32470;
  assign new_n32475 = new_n32474 ^ new_n32464;
  assign new_n32476 = new_n32388 & new_n32461;
  assign new_n32477 = new_n32439 ^ new_n32417;
  assign new_n32478 = new_n32477 ^ new_n32464;
  assign new_n32479 = new_n32417 ^ new_n32308;
  assign new_n32480 = new_n32478 & new_n32479;
  assign new_n32481 = new_n32480 ^ new_n32476;
  assign new_n32482 = new_n32439 ^ new_n32352;
  assign new_n32483 = new_n32482 ^ new_n32481;
  assign new_n32484 = new_n32483 ^ new_n32475;
  assign new_n32485 = new_n32467 ^ new_n32462;
  assign new_n32486 = new_n32441 ^ new_n32385;
  assign new_n32487 = new_n32486 ^ new_n32464;
  assign new_n32488 = new_n32462 ^ new_n32400;
  assign new_n32489 = new_n32487 & new_n32488;
  assign new_n32490 = new_n32489 ^ new_n32476;
  assign new_n32491 = new_n32480 ^ new_n32308;
  assign new_n32492 = new_n32491 ^ new_n32490;
  assign new_n32493 = new_n32492 ^ new_n32485;
  assign new_n32494 = ~new_n32484 & new_n32493;
  assign new_n32495 = new_n32494 ^ new_n32468;
  assign new_n32496 = new_n32462 ^ new_n32440;
  assign new_n32497 = new_n32464 & new_n32496;
  assign new_n32498 = new_n32497 ^ new_n32476;
  assign new_n32499 = new_n32498 ^ new_n32471;
  assign new_n32500 = new_n32499 ^ new_n32495;
  assign new_n32501 = new_n32460 ^ new_n32441;
  assign new_n32502 = new_n32400 ^ new_n32388;
  assign new_n32503 = new_n32501 & new_n32502;
  assign new_n32504 = new_n32503 ^ new_n32469;
  assign new_n32505 = new_n32497 ^ new_n32480;
  assign new_n32506 = new_n32505 ^ new_n32504;
  assign new_n32507 = ~new_n32506 & new_n32500;
  assign new_n32508 = new_n32460 ^ new_n32439;
  assign new_n32509 = new_n32489 ^ new_n32443;
  assign new_n32510 = new_n32509 ^ new_n32505;
  assign new_n32511 = new_n32510 ^ new_n32508;
  assign new_n32512 = new_n32503 ^ new_n32473;
  assign new_n32513 = new_n32512 ^ new_n32460;
  assign new_n32514 = new_n32513 ^ new_n32499;
  assign new_n32515 = new_n32514 ^ new_n32494;
  assign new_n32516 = new_n32511 & new_n32515;
  assign new_n32517 = new_n32516 ^ new_n32507;
  assign new_n32518 = new_n32513 ^ new_n32468;
  assign new_n32519 = new_n32518 ^ new_n32517;
  assign new_n32520 = new_n32388 & new_n32519;
  assign new_n32521 = new_n32507 ^ new_n32494;
  assign new_n32522 = new_n32514 & new_n32521;
  assign new_n32523 = new_n32522 ^ new_n32484;
  assign new_n32524 = ~new_n32523 & new_n32465;
  assign new_n32525 = new_n32524 ^ new_n32520;
  assign new_n32526 = new_n32439 ^ new_n32385;
  assign new_n32527 = new_n32489 ^ new_n32470;
  assign new_n32528 = new_n32516 ^ new_n32468;
  assign new_n32529 = new_n32528 ^ new_n32499;
  assign new_n32530 = new_n32522 ^ new_n32515;
  assign new_n32531 = new_n32529 & new_n32530;
  assign new_n32532 = new_n32531 ^ new_n32522;
  assign new_n32533 = new_n32532 ^ new_n32527;
  assign new_n32534 = new_n32533 ^ new_n32526;
  assign new_n32535 = new_n32534 ^ new_n32417;
  assign new_n32536 = new_n32516 ^ new_n32473;
  assign new_n32537 = new_n32536 ^ new_n32467;
  assign new_n32538 = new_n32537 ^ new_n32535;
  assign new_n32539 = ~new_n32538 & new_n32478;
  assign new_n32540 = new_n32531 ^ new_n32511;
  assign new_n32541 = new_n32441 & new_n32540;
  assign new_n32542 = new_n32522 ^ new_n32507;
  assign new_n32543 = new_n32542 ^ new_n32506;
  assign new_n32544 = ~new_n32543 & new_n32487;
  assign new_n32545 = ~new_n32538 & new_n32479;
  assign new_n32546 = new_n32461 & new_n32519;
  assign new_n32547 = new_n32546 ^ new_n32545;
  assign new_n32548 = new_n32547 ^ new_n32544;
  assign new_n32549 = new_n32548 ^ new_n32541;
  assign new_n32550 = new_n32531 ^ new_n32516;
  assign new_n32551 = new_n32550 ^ new_n32493;
  assign new_n32552 = new_n32471 & new_n32551;
  assign new_n32553 = new_n32552 ^ new_n32549;
  assign new_n32554 = new_n32553 ^ new_n32539;
  assign new_n32555 = new_n32554 ^ new_n32525;
  assign new_n32556 = new_n30788 ^ new_n18928;
  assign new_n32557 = new_n31029 ^ new_n18926;
  assign new_n32558 = new_n31091 ^ new_n18923;
  assign new_n32559 = new_n31122 ^ new_n18924;
  assign new_n32560 = new_n32559 ^ new_n32558;
  assign new_n32561 = new_n32560 ^ new_n32557;
  assign new_n32562 = new_n32561 ^ new_n32556;
  assign new_n32563 = new_n31141 ^ new_n18930;
  assign new_n32564 = new_n31154 ^ new_n18934;
  assign new_n32565 = new_n31176 ^ new_n18931;
  assign new_n32566 = new_n32565 ^ new_n32556;
  assign new_n32567 = new_n32566 ^ new_n32563;
  assign new_n32568 = new_n32567 ^ new_n32564;
  assign new_n32569 = ~new_n32563 & ~new_n32568;
  assign new_n32570 = new_n32569 ^ new_n32564;
  assign new_n32571 = new_n31191 ^ new_n18938;
  assign new_n32572 = new_n32571 ^ new_n32564;
  assign new_n32573 = new_n32572 ^ new_n32560;
  assign new_n32574 = new_n32564 ^ new_n32559;
  assign new_n32575 = new_n32571 ^ new_n32557;
  assign new_n32576 = new_n32575 ^ new_n32574;
  assign new_n32577 = ~new_n32573 & ~new_n32576;
  assign new_n32578 = new_n32577 ^ new_n32556;
  assign new_n32579 = new_n32578 ^ new_n32570;
  assign new_n32580 = new_n32559 & new_n32567;
  assign new_n32581 = new_n32580 ^ new_n32559;
  assign new_n32582 = new_n32565 ^ new_n32561;
  assign new_n32583 = new_n32571 ^ new_n32559;
  assign new_n32584 = ~new_n32583 & new_n32582;
  assign new_n32585 = new_n32584 ^ new_n32581;
  assign new_n32586 = new_n32585 ^ new_n32575;
  assign new_n32587 = new_n32562 & new_n32572;
  assign new_n32588 = new_n32565 ^ new_n32564;
  assign new_n32589 = new_n32588 ^ new_n32575;
  assign new_n32590 = new_n32564 ^ new_n32557;
  assign new_n32591 = ~new_n32589 & new_n32590;
  assign new_n32592 = new_n32591 ^ new_n32587;
  assign new_n32593 = new_n32565 ^ new_n32558;
  assign new_n32594 = new_n32593 ^ new_n32592;
  assign new_n32595 = new_n32594 ^ new_n32586;
  assign new_n32596 = new_n32578 ^ new_n32573;
  assign new_n32597 = new_n32567 ^ new_n32559;
  assign new_n32598 = new_n32597 ^ new_n32575;
  assign new_n32599 = new_n32573 ^ new_n32563;
  assign new_n32600 = new_n32598 & new_n32599;
  assign new_n32601 = new_n32600 ^ new_n32557;
  assign new_n32602 = new_n32601 ^ new_n32592;
  assign new_n32603 = new_n32602 ^ new_n32596;
  assign new_n32604 = ~new_n32595 & new_n32603;
  assign new_n32605 = new_n32604 ^ new_n32579;
  assign new_n32606 = new_n32573 ^ new_n32566;
  assign new_n32607 = ~new_n32606 & new_n32575;
  assign new_n32608 = new_n32607 ^ new_n32587;
  assign new_n32609 = new_n32608 ^ new_n32582;
  assign new_n32610 = new_n32609 ^ new_n32605;
  assign new_n32611 = new_n32571 ^ new_n32567;
  assign new_n32612 = new_n32563 ^ new_n32562;
  assign new_n32613 = ~new_n32611 & ~new_n32612;
  assign new_n32614 = new_n32613 ^ new_n32580;
  assign new_n32615 = new_n32607 ^ new_n32591;
  assign new_n32616 = new_n32615 ^ new_n32614;
  assign new_n32617 = ~new_n32610 & ~new_n32616;
  assign new_n32618 = new_n32571 ^ new_n32565;
  assign new_n32619 = new_n32600 ^ new_n32569;
  assign new_n32620 = new_n32619 ^ new_n32615;
  assign new_n32621 = new_n32620 ^ new_n32618;
  assign new_n32622 = new_n32613 ^ new_n32584;
  assign new_n32623 = new_n32622 ^ new_n32571;
  assign new_n32624 = new_n32623 ^ new_n32609;
  assign new_n32625 = new_n32624 ^ new_n32604;
  assign new_n32626 = ~new_n32621 & new_n32625;
  assign new_n32627 = new_n32626 ^ new_n32617;
  assign new_n32628 = new_n32623 ^ new_n32579;
  assign new_n32629 = new_n32628 ^ new_n32627;
  assign new_n32630 = ~new_n32629 & new_n32562;
  assign new_n32631 = new_n32617 ^ new_n32604;
  assign new_n32632 = new_n32624 & new_n32631;
  assign new_n32633 = new_n32632 ^ new_n32595;
  assign new_n32634 = ~new_n32576 & ~new_n32633;
  assign new_n32635 = new_n32634 ^ new_n32630;
  assign new_n32636 = new_n32565 ^ new_n32559;
  assign new_n32637 = new_n32600 ^ new_n32581;
  assign new_n32638 = new_n32626 ^ new_n32579;
  assign new_n32639 = new_n32638 ^ new_n32609;
  assign new_n32640 = new_n32632 ^ new_n32625;
  assign new_n32641 = ~new_n32639 & new_n32640;
  assign new_n32642 = new_n32641 ^ new_n32632;
  assign new_n32643 = new_n32642 ^ new_n32637;
  assign new_n32644 = new_n32643 ^ new_n32636;
  assign new_n32645 = new_n32644 ^ new_n32564;
  assign new_n32646 = new_n32626 ^ new_n32584;
  assign new_n32647 = new_n32646 ^ new_n32578;
  assign new_n32648 = new_n32647 ^ new_n32645;
  assign new_n32649 = ~new_n32589 & ~new_n32648;
  assign new_n32650 = new_n32641 ^ new_n32621;
  assign new_n32651 = ~new_n32567 & ~new_n32650;
  assign new_n32652 = new_n32632 ^ new_n32617;
  assign new_n32653 = new_n32652 ^ new_n32616;
  assign new_n32654 = ~new_n32653 & new_n32598;
  assign new_n32655 = ~new_n32648 & new_n32590;
  assign new_n32656 = ~new_n32629 & new_n32572;
  assign new_n32657 = new_n32656 ^ new_n32655;
  assign new_n32658 = new_n32657 ^ new_n32654;
  assign new_n32659 = new_n32658 ^ new_n32651;
  assign new_n32660 = new_n32641 ^ new_n32626;
  assign new_n32661 = new_n32660 ^ new_n32603;
  assign new_n32662 = new_n32582 & new_n32661;
  assign new_n32663 = new_n32662 ^ new_n32659;
  assign new_n32664 = new_n32663 ^ new_n32649;
  assign new_n32665 = new_n32664 ^ new_n32635;
  assign new_n32666 = new_n32665 ^ new_n22837;
  assign new_n32667 = new_n32666 ^ new_n32555;
  assign new_n32668 = new_n32649 ^ new_n32630;
  assign new_n32669 = ~new_n32573 & ~new_n32633;
  assign new_n32670 = ~new_n32653 & new_n32599;
  assign new_n32671 = new_n32670 ^ new_n32669;
  assign new_n32672 = new_n32671 ^ new_n32634;
  assign new_n32673 = new_n32672 ^ new_n32658;
  assign new_n32674 = new_n32673 ^ new_n32668;
  assign new_n32675 = new_n32674 ^ new_n22874;
  assign new_n32676 = new_n32539 ^ new_n32520;
  assign new_n32677 = ~new_n32523 & new_n32462;
  assign new_n32678 = ~new_n32543 & new_n32488;
  assign new_n32679 = new_n32678 ^ new_n32677;
  assign new_n32680 = new_n32679 ^ new_n32524;
  assign new_n32681 = new_n32680 ^ new_n32548;
  assign new_n32682 = new_n32681 ^ new_n32676;
  assign new_n32683 = new_n32682 ^ new_n32675;
  assign new_n32684 = new_n32656 ^ new_n32630;
  assign new_n32685 = new_n32617 ^ new_n32571;
  assign new_n32686 = new_n32613 ^ new_n32569;
  assign new_n32687 = new_n32686 ^ new_n32644;
  assign new_n32688 = new_n32687 ^ new_n32685;
  assign new_n32689 = new_n32575 & new_n32688;
  assign new_n32690 = ~new_n32583 & new_n32661;
  assign new_n32691 = new_n32624 ^ new_n32617;
  assign new_n32692 = ~new_n32563 & new_n32691;
  assign new_n32693 = new_n32692 ^ new_n32669;
  assign new_n32694 = new_n32693 ^ new_n32690;
  assign new_n32695 = ~new_n32606 & new_n32688;
  assign new_n32696 = ~new_n32611 & ~new_n32639;
  assign new_n32697 = new_n32696 ^ new_n32695;
  assign new_n32698 = new_n32697 ^ new_n32694;
  assign new_n32699 = new_n32698 ^ new_n32689;
  assign new_n32700 = new_n32699 ^ new_n32684;
  assign new_n32701 = new_n32700 ^ new_n22882;
  assign new_n32702 = new_n32546 ^ new_n32520;
  assign new_n32703 = new_n32507 ^ new_n32460;
  assign new_n32704 = new_n32503 ^ new_n32443;
  assign new_n32705 = new_n32704 ^ new_n32534;
  assign new_n32706 = new_n32705 ^ new_n32703;
  assign new_n32707 = ~new_n32706 & new_n32464;
  assign new_n32708 = new_n32472 & new_n32551;
  assign new_n32709 = new_n32514 ^ new_n32507;
  assign new_n32710 = new_n32400 & new_n32709;
  assign new_n32711 = new_n32710 ^ new_n32677;
  assign new_n32712 = new_n32711 ^ new_n32708;
  assign new_n32713 = ~new_n32706 & new_n32496;
  assign new_n32714 = new_n32501 & new_n32529;
  assign new_n32715 = new_n32714 ^ new_n32713;
  assign new_n32716 = new_n32715 ^ new_n32712;
  assign new_n32717 = new_n32716 ^ new_n32707;
  assign new_n32718 = new_n32717 ^ new_n32702;
  assign new_n32719 = new_n32718 ^ new_n32701;
  assign new_n32720 = new_n32680 ^ new_n32553;
  assign new_n32721 = new_n32672 ^ new_n32663;
  assign new_n32722 = new_n32721 ^ new_n22842;
  assign new_n32723 = new_n32722 ^ new_n32720;
  assign new_n32724 = new_n32502 & new_n32529;
  assign new_n32725 = new_n32724 ^ new_n32524;
  assign new_n32726 = new_n32710 ^ new_n32678;
  assign new_n32727 = new_n32726 ^ new_n32549;
  assign new_n32728 = new_n32727 ^ new_n32725;
  assign new_n32729 = ~new_n32612 & ~new_n32639;
  assign new_n32730 = new_n32729 ^ new_n32634;
  assign new_n32731 = new_n32692 ^ new_n32670;
  assign new_n32732 = new_n32731 ^ new_n32659;
  assign new_n32733 = new_n32732 ^ new_n32730;
  assign new_n32734 = new_n32733 ^ new_n22857;
  assign new_n32735 = new_n32734 ^ new_n32728;
  assign new_n32736 = new_n32442 & new_n32709;
  assign new_n32737 = new_n32736 ^ new_n32554;
  assign new_n32738 = new_n32737 ^ new_n32716;
  assign new_n32739 = ~new_n32568 & new_n32691;
  assign new_n32740 = new_n32739 ^ new_n32664;
  assign new_n32741 = new_n32740 ^ new_n32698;
  assign new_n32742 = new_n32741 ^ new_n22869;
  assign new_n32743 = new_n32742 ^ new_n32738;
  assign new_n32744 = new_n32695 ^ new_n32690;
  assign new_n32745 = ~new_n32650 & new_n32597;
  assign new_n32746 = new_n32745 ^ new_n32729;
  assign new_n32747 = new_n32746 ^ new_n32657;
  assign new_n32748 = new_n32651 ^ new_n32649;
  assign new_n32749 = new_n32748 ^ new_n32747;
  assign new_n32750 = new_n32749 ^ new_n32744;
  assign new_n32751 = new_n32750 ^ new_n22851;
  assign new_n32752 = new_n32713 ^ new_n32708;
  assign new_n32753 = new_n32486 & new_n32540;
  assign new_n32754 = new_n32753 ^ new_n32724;
  assign new_n32755 = new_n32754 ^ new_n32547;
  assign new_n32756 = new_n32541 ^ new_n32539;
  assign new_n32757 = new_n32756 ^ new_n32755;
  assign new_n32758 = new_n32757 ^ new_n32752;
  assign new_n32759 = new_n32758 ^ new_n32751;
  assign new_n32760 = new_n32694 ^ new_n32662;
  assign new_n32761 = new_n32760 ^ new_n32747;
  assign new_n32762 = new_n32761 ^ new_n22863;
  assign new_n32763 = new_n32712 ^ new_n32552;
  assign new_n32764 = new_n32763 ^ new_n32755;
  assign new_n32765 = new_n32764 ^ new_n32762;
  assign new_n32766 = new_n30231 ^ new_n27088;
  assign new_n32767 = new_n28466 ^ new_n27148;
  assign new_n32768 = new_n32767 ^ new_n27016;
  assign new_n32769 = new_n32768 ^ new_n32766;
  assign new_n32770 = new_n27049 ^ new_n26355;
  assign new_n32771 = new_n32770 ^ new_n27136;
  assign new_n32772 = new_n32771 ^ new_n30222;
  assign new_n32773 = new_n28480 ^ new_n27016;
  assign new_n32774 = new_n32773 ^ new_n27071;
  assign new_n32775 = new_n32774 ^ new_n32772;
  assign new_n32776 = new_n30269 ^ new_n28500;
  assign new_n32777 = new_n32776 ^ new_n32770;
  assign new_n32778 = new_n27026 ^ new_n26913;
  assign new_n32779 = new_n32778 ^ new_n27148;
  assign new_n32780 = new_n32779 ^ new_n32777;
  assign new_n32781 = new_n32780 ^ new_n32775;
  assign new_n32782 = new_n32781 ^ new_n32769;
  assign new_n32783 = new_n27125 ^ new_n26941;
  assign new_n32784 = new_n28485 ^ new_n27059;
  assign new_n32785 = new_n32784 ^ new_n27120;
  assign new_n32786 = new_n32785 ^ new_n32783;
  assign new_n32787 = new_n32786 ^ new_n32782;
  assign new_n32788 = new_n27120 ^ new_n27000;
  assign new_n32789 = new_n26965 ^ new_n26905;
  assign new_n32790 = new_n32789 ^ new_n28459;
  assign new_n32791 = new_n32790 ^ new_n32788;
  assign new_n32792 = new_n32791 ^ new_n32786;
  assign new_n32793 = new_n28489 ^ new_n27071;
  assign new_n32794 = new_n32770 ^ new_n30226;
  assign new_n32795 = new_n32794 ^ new_n32793;
  assign new_n32796 = new_n32795 ^ new_n32792;
  assign new_n32797 = new_n32775 & new_n32796;
  assign new_n32798 = new_n32797 ^ new_n32775;
  assign new_n32799 = new_n32791 ^ new_n32782;
  assign new_n32800 = new_n27108 ^ new_n27063;
  assign new_n32801 = new_n28469 ^ new_n26355;
  assign new_n32802 = new_n32801 ^ new_n27059;
  assign new_n32803 = new_n32802 ^ new_n32800;
  assign new_n32804 = new_n32803 ^ new_n32775;
  assign new_n32805 = ~new_n32799 & new_n32804;
  assign new_n32806 = new_n32805 ^ new_n32798;
  assign new_n32807 = new_n32803 ^ new_n32769;
  assign new_n32808 = new_n32807 ^ new_n32806;
  assign new_n32809 = new_n32770 ^ new_n28440;
  assign new_n32810 = new_n32809 ^ new_n26766;
  assign new_n32811 = new_n27158 ^ new_n26965;
  assign new_n32812 = new_n32811 ^ new_n26913;
  assign new_n32813 = new_n32812 ^ new_n32810;
  assign new_n32814 = new_n32813 ^ new_n32791;
  assign new_n32815 = new_n32814 ^ new_n32807;
  assign new_n32816 = new_n32813 ^ new_n32769;
  assign new_n32817 = new_n32815 & new_n32816;
  assign new_n32818 = new_n32813 ^ new_n32803;
  assign new_n32819 = ~new_n32787 & ~new_n32818;
  assign new_n32820 = new_n32819 ^ new_n32817;
  assign new_n32821 = new_n32791 ^ new_n32780;
  assign new_n32822 = new_n32821 ^ new_n32820;
  assign new_n32823 = new_n32822 ^ new_n32808;
  assign new_n32824 = new_n32818 ^ new_n32781;
  assign new_n32825 = new_n32813 ^ new_n32775;
  assign new_n32826 = new_n32825 ^ new_n32807;
  assign new_n32827 = ~new_n32824 & new_n32826;
  assign new_n32828 = new_n32827 ^ new_n32786;
  assign new_n32829 = new_n32828 ^ new_n32824;
  assign new_n32830 = new_n32824 ^ new_n32795;
  assign new_n32831 = new_n32796 ^ new_n32775;
  assign new_n32832 = new_n32831 ^ new_n32807;
  assign new_n32833 = ~new_n32832 & new_n32830;
  assign new_n32834 = new_n32833 ^ new_n32820;
  assign new_n32835 = new_n32834 ^ new_n32769;
  assign new_n32836 = new_n32835 ^ new_n32829;
  assign new_n32837 = ~new_n32823 & new_n32836;
  assign new_n32838 = new_n32824 ^ new_n32792;
  assign new_n32839 = ~new_n32807 & ~new_n32838;
  assign new_n32840 = new_n32839 ^ new_n32819;
  assign new_n32841 = new_n32840 ^ new_n32799;
  assign new_n32842 = new_n32803 ^ new_n32796;
  assign new_n32843 = new_n32795 ^ new_n32787;
  assign new_n32844 = new_n32842 & new_n32843;
  assign new_n32845 = new_n32844 ^ new_n32805;
  assign new_n32846 = new_n32845 ^ new_n32803;
  assign new_n32847 = new_n32846 ^ new_n32841;
  assign new_n32848 = new_n32847 ^ new_n32837;
  assign new_n32849 = new_n32803 ^ new_n32791;
  assign new_n32850 = new_n32813 ^ new_n32796;
  assign new_n32851 = ~new_n32795 & ~new_n32850;
  assign new_n32852 = new_n32851 ^ new_n32833;
  assign new_n32853 = new_n32839 ^ new_n32817;
  assign new_n32854 = new_n32853 ^ new_n32852;
  assign new_n32855 = new_n32854 ^ new_n32849;
  assign new_n32856 = new_n32848 & new_n32855;
  assign new_n32857 = new_n32851 ^ new_n32813;
  assign new_n32858 = new_n32857 ^ new_n32828;
  assign new_n32859 = new_n32858 ^ new_n32837;
  assign new_n32860 = new_n32859 ^ new_n32841;
  assign new_n32861 = new_n32844 ^ new_n32797;
  assign new_n32862 = new_n32861 ^ new_n32853;
  assign new_n32863 = ~new_n32862 & new_n32860;
  assign new_n32864 = new_n32863 ^ new_n32856;
  assign new_n32865 = new_n32858 ^ new_n32846;
  assign new_n32866 = new_n32865 ^ new_n32864;
  assign new_n32867 = ~new_n32787 & new_n32866;
  assign new_n32868 = ~new_n32818 & new_n32866;
  assign new_n32869 = new_n32868 ^ new_n32867;
  assign new_n32870 = new_n32863 ^ new_n32803;
  assign new_n32871 = new_n32851 ^ new_n32844;
  assign new_n32872 = new_n32791 ^ new_n32775;
  assign new_n32873 = new_n32833 ^ new_n32798;
  assign new_n32874 = new_n32858 ^ new_n32856;
  assign new_n32875 = new_n32874 ^ new_n32841;
  assign new_n32876 = new_n32863 ^ new_n32837;
  assign new_n32877 = ~new_n32876 & new_n32847;
  assign new_n32878 = new_n32877 ^ new_n32837;
  assign new_n32879 = new_n32875 & new_n32878;
  assign new_n32880 = new_n32877 ^ new_n32847;
  assign new_n32881 = new_n32880 ^ new_n32879;
  assign new_n32882 = new_n32881 ^ new_n32873;
  assign new_n32883 = new_n32882 ^ new_n32872;
  assign new_n32884 = new_n32883 ^ new_n32871;
  assign new_n32885 = new_n32884 ^ new_n32870;
  assign new_n32886 = ~new_n32807 & ~new_n32885;
  assign new_n32887 = new_n32842 & new_n32875;
  assign new_n32888 = ~new_n32838 & ~new_n32885;
  assign new_n32889 = new_n32888 ^ new_n32887;
  assign new_n32890 = new_n32879 ^ new_n32856;
  assign new_n32891 = new_n32890 ^ new_n32836;
  assign new_n32892 = new_n32804 & new_n32891;
  assign new_n32893 = new_n32863 ^ new_n32847;
  assign new_n32894 = ~new_n32795 & new_n32893;
  assign new_n32895 = new_n32880 ^ new_n32823;
  assign new_n32896 = ~new_n32824 & ~new_n32895;
  assign new_n32897 = new_n32896 ^ new_n32894;
  assign new_n32898 = new_n32897 ^ new_n32892;
  assign new_n32899 = new_n32898 ^ new_n32889;
  assign new_n32900 = new_n32899 ^ new_n32886;
  assign new_n32901 = new_n32900 ^ new_n32869;
  assign new_n32902 = new_n26110 ^ new_n22415;
  assign new_n32903 = new_n32902 ^ new_n15496;
  assign new_n32904 = new_n32903 ^ new_n30801;
  assign new_n32905 = new_n32904 ^ new_n31837;
  assign new_n32906 = new_n29379 ^ new_n29238;
  assign new_n32907 = new_n32906 ^ new_n29164;
  assign new_n32908 = new_n32907 ^ new_n32905;
  assign new_n32909 = new_n30830 ^ new_n29341;
  assign new_n32910 = new_n26064 ^ new_n22328;
  assign new_n32911 = new_n32910 ^ new_n15463;
  assign new_n32912 = new_n29238 ^ new_n28869;
  assign new_n32913 = new_n32912 ^ new_n32911;
  assign new_n32914 = new_n32913 ^ new_n32909;
  assign new_n32915 = new_n32914 ^ new_n32908;
  assign new_n32916 = new_n30849 ^ new_n29317;
  assign new_n32917 = new_n25010 ^ new_n22470;
  assign new_n32918 = new_n32917 ^ new_n15508;
  assign new_n32919 = new_n32918 ^ new_n29385;
  assign new_n32920 = new_n32919 ^ new_n29291;
  assign new_n32921 = new_n32920 ^ new_n32916;
  assign new_n32922 = new_n30795 ^ new_n29349;
  assign new_n32923 = new_n26100 ^ new_n22259;
  assign new_n32924 = new_n32923 ^ new_n15492;
  assign new_n32925 = new_n32924 ^ new_n29154;
  assign new_n32926 = new_n32925 ^ new_n29258;
  assign new_n32927 = new_n32926 ^ new_n32922;
  assign new_n32928 = new_n32927 ^ new_n32921;
  assign new_n32929 = new_n32928 ^ new_n32915;
  assign new_n32930 = new_n31837 ^ new_n29360;
  assign new_n32931 = new_n32930 ^ new_n30808;
  assign new_n32932 = new_n25968 ^ new_n21185;
  assign new_n32933 = new_n32932 ^ new_n15478;
  assign new_n32934 = new_n32933 ^ new_n29291;
  assign new_n32935 = new_n32934 ^ new_n29328;
  assign new_n32936 = new_n32935 ^ new_n32931;
  assign new_n32937 = new_n32936 ^ new_n32914;
  assign new_n32938 = new_n30814 ^ new_n29230;
  assign new_n32939 = new_n26036 ^ new_n22445;
  assign new_n32940 = new_n32939 ^ new_n15469;
  assign new_n32941 = new_n32940 ^ new_n29258;
  assign new_n32942 = new_n32941 ^ new_n29341;
  assign new_n32943 = new_n32942 ^ new_n32938;
  assign new_n32944 = new_n32943 ^ new_n32914;
  assign new_n32945 = new_n26076 ^ new_n22360;
  assign new_n32946 = new_n32945 ^ new_n15518;
  assign new_n32947 = new_n32946 ^ new_n29328;
  assign new_n32948 = new_n31837 ^ new_n30819;
  assign new_n32949 = new_n32948 ^ new_n32947;
  assign new_n32950 = new_n32949 ^ new_n32944;
  assign new_n32951 = new_n32936 & new_n32950;
  assign new_n32952 = new_n32951 ^ new_n32936;
  assign new_n32953 = new_n32950 ^ new_n32936;
  assign new_n32954 = new_n32953 ^ new_n32928;
  assign new_n32955 = new_n32927 ^ new_n32908;
  assign new_n32956 = new_n29269 ^ new_n29164;
  assign new_n32957 = new_n32956 ^ new_n29385;
  assign new_n32958 = new_n26006 ^ new_n22391;
  assign new_n32959 = new_n32958 ^ new_n15484;
  assign new_n32960 = new_n32959 ^ new_n31837;
  assign new_n32961 = new_n32960 ^ new_n30790;
  assign new_n32962 = new_n32961 ^ new_n32957;
  assign new_n32963 = new_n32962 ^ new_n32936;
  assign new_n32964 = new_n32963 ^ new_n32955;
  assign new_n32965 = new_n32964 ^ new_n32949;
  assign new_n32966 = new_n32954 & new_n32965;
  assign new_n32967 = new_n32966 ^ new_n32952;
  assign new_n32968 = new_n32936 ^ new_n32927;
  assign new_n32969 = new_n32921 ^ new_n32908;
  assign new_n32970 = new_n32969 ^ new_n32968;
  assign new_n32971 = ~new_n32964 & ~new_n32970;
  assign new_n32972 = new_n32971 ^ new_n32943;
  assign new_n32973 = ~new_n32944 & ~new_n32949;
  assign new_n32974 = new_n32908 & new_n32949;
  assign new_n32975 = new_n32974 ^ new_n32973;
  assign new_n32976 = new_n32975 ^ new_n32972;
  assign new_n32977 = new_n32927 ^ new_n32914;
  assign new_n32978 = new_n32964 ^ new_n32944;
  assign new_n32979 = ~new_n32978 & new_n32928;
  assign new_n32980 = ~new_n32929 & new_n32969;
  assign new_n32981 = new_n32980 ^ new_n32979;
  assign new_n32982 = new_n32975 ^ new_n32908;
  assign new_n32983 = new_n32982 ^ new_n32966;
  assign new_n32984 = new_n32983 ^ new_n32981;
  assign new_n32985 = new_n32984 ^ new_n32977;
  assign new_n32986 = new_n32963 ^ new_n32921;
  assign new_n32987 = new_n32986 ^ new_n32943;
  assign new_n32988 = new_n32955 & new_n32987;
  assign new_n32989 = new_n32988 ^ new_n32979;
  assign new_n32990 = new_n32986 ^ new_n32914;
  assign new_n32991 = new_n32990 ^ new_n32989;
  assign new_n32992 = ~new_n32968 & new_n32990;
  assign new_n32993 = new_n32950 ^ new_n32927;
  assign new_n32994 = new_n32987 ^ new_n32949;
  assign new_n32995 = ~new_n32993 & ~new_n32994;
  assign new_n32996 = new_n32995 ^ new_n32992;
  assign new_n32997 = new_n32996 ^ new_n32927;
  assign new_n32998 = new_n32997 ^ new_n32991;
  assign new_n32999 = new_n32992 ^ new_n32952;
  assign new_n33000 = new_n32999 ^ new_n32928;
  assign new_n33001 = new_n32988 ^ new_n32980;
  assign new_n33002 = new_n32962 ^ new_n32914;
  assign new_n33003 = new_n33002 ^ new_n33001;
  assign new_n33004 = new_n33003 ^ new_n33000;
  assign new_n33005 = new_n32972 ^ new_n32964;
  assign new_n33006 = new_n33001 ^ new_n32966;
  assign new_n33007 = new_n33006 ^ new_n32921;
  assign new_n33008 = new_n33007 ^ new_n33005;
  assign new_n33009 = ~new_n33004 & new_n33008;
  assign new_n33010 = new_n33009 ^ new_n32998;
  assign new_n33011 = ~new_n32985 & new_n33010;
  assign new_n33012 = new_n33011 ^ new_n32976;
  assign new_n33013 = new_n33012 ^ new_n32991;
  assign new_n33014 = new_n33009 ^ new_n32976;
  assign new_n33015 = new_n33014 ^ new_n32991;
  assign new_n33016 = new_n32995 ^ new_n32951;
  assign new_n33017 = new_n33016 ^ new_n32981;
  assign new_n33018 = ~new_n33015 & ~new_n33017;
  assign new_n33019 = new_n33018 ^ new_n33009;
  assign new_n33020 = new_n32998 & new_n33019;
  assign new_n33021 = new_n33020 ^ new_n33010;
  assign new_n33022 = ~new_n33013 & new_n33021;
  assign new_n33023 = new_n33022 ^ new_n33020;
  assign new_n33024 = new_n33023 ^ new_n32967;
  assign new_n33025 = new_n33024 ^ new_n32937;
  assign new_n33026 = new_n33025 ^ new_n32908;
  assign new_n33027 = new_n33011 ^ new_n32992;
  assign new_n33028 = new_n33027 ^ new_n32972;
  assign new_n33029 = new_n33028 ^ new_n33026;
  assign new_n33030 = ~new_n32929 & ~new_n33029;
  assign new_n33031 = new_n33018 ^ new_n33011;
  assign new_n33032 = new_n32997 ^ new_n32976;
  assign new_n33033 = new_n33032 ^ new_n33031;
  assign new_n33034 = ~new_n33033 & new_n32987;
  assign new_n33035 = new_n33034 ^ new_n33030;
  assign new_n33036 = new_n33020 ^ new_n33018;
  assign new_n33037 = new_n33036 ^ new_n33017;
  assign new_n33038 = ~new_n33037 & new_n32965;
  assign new_n33039 = new_n33020 ^ new_n33004;
  assign new_n33040 = ~new_n32964 & ~new_n33039;
  assign new_n33041 = new_n33040 ^ new_n33038;
  assign new_n33042 = ~new_n32970 & ~new_n33039;
  assign new_n33043 = new_n33042 ^ new_n33041;
  assign new_n33044 = ~new_n33037 & new_n32954;
  assign new_n33045 = ~new_n33029 & new_n32969;
  assign new_n33046 = ~new_n33033 & new_n32955;
  assign new_n33047 = new_n33046 ^ new_n33045;
  assign new_n33048 = new_n33047 ^ new_n33044;
  assign new_n33049 = new_n33048 ^ new_n33043;
  assign new_n33050 = new_n33049 ^ new_n33035;
  assign new_n33051 = new_n27966 ^ new_n23681;
  assign new_n33052 = new_n33051 ^ new_n30549;
  assign new_n33053 = new_n33052 ^ new_n30584;
  assign new_n33054 = new_n26112 ^ new_n26071;
  assign new_n33055 = new_n33054 ^ new_n33053;
  assign new_n33056 = new_n30529 ^ new_n26016;
  assign new_n33057 = new_n28022 ^ new_n23708;
  assign new_n33058 = new_n33057 ^ new_n26058;
  assign new_n33059 = new_n33058 ^ new_n26047;
  assign new_n33060 = new_n33059 ^ new_n33056;
  assign new_n33061 = new_n33060 ^ new_n33055;
  assign new_n33062 = new_n25980 ^ new_n23663;
  assign new_n33063 = new_n33062 ^ new_n25905;
  assign new_n33064 = new_n28100 ^ new_n23701;
  assign new_n33065 = new_n33064 ^ new_n30557;
  assign new_n33066 = new_n33065 ^ new_n33063;
  assign new_n33067 = new_n28116 ^ new_n23677;
  assign new_n33068 = new_n33067 ^ new_n30565;
  assign new_n33069 = new_n26094 ^ new_n25941;
  assign new_n33070 = new_n33069 ^ new_n33068;
  assign new_n33071 = new_n33070 ^ new_n33066;
  assign new_n33072 = new_n33071 ^ new_n33061;
  assign new_n33073 = new_n30549 ^ new_n22574;
  assign new_n33074 = new_n33073 ^ new_n30574;
  assign new_n33075 = new_n28158 ^ new_n23666;
  assign new_n33076 = new_n33075 ^ new_n25958;
  assign new_n33077 = new_n33076 ^ new_n25914;
  assign new_n33078 = new_n33077 ^ new_n33074;
  assign new_n33079 = new_n33078 ^ new_n33060;
  assign new_n33080 = new_n30539 ^ new_n26092;
  assign new_n33081 = new_n28178 ^ new_n23695;
  assign new_n33082 = new_n33081 ^ new_n26028;
  assign new_n33083 = new_n33082 ^ new_n26042;
  assign new_n33084 = new_n33083 ^ new_n33080;
  assign new_n33085 = new_n33084 ^ new_n33060;
  assign new_n33086 = new_n30549 ^ new_n25925;
  assign new_n33087 = new_n28200 ^ new_n23689;
  assign new_n33088 = new_n33087 ^ new_n26082;
  assign new_n33089 = new_n33088 ^ new_n25972;
  assign new_n33090 = new_n33089 ^ new_n33086;
  assign new_n33091 = new_n33090 ^ new_n33085;
  assign new_n33092 = new_n33078 & new_n33091;
  assign new_n33093 = new_n33092 ^ new_n33078;
  assign new_n33094 = new_n33091 ^ new_n33078;
  assign new_n33095 = new_n33094 ^ new_n33071;
  assign new_n33096 = new_n33070 ^ new_n33055;
  assign new_n33097 = new_n26120 ^ new_n25993;
  assign new_n33098 = new_n33097 ^ new_n25985;
  assign new_n33099 = new_n28222 ^ new_n23672;
  assign new_n33100 = new_n33099 ^ new_n30549;
  assign new_n33101 = new_n33100 ^ new_n30543;
  assign new_n33102 = new_n33101 ^ new_n33098;
  assign new_n33103 = new_n33102 ^ new_n33078;
  assign new_n33104 = new_n33103 ^ new_n33096;
  assign new_n33105 = new_n33104 ^ new_n33090;
  assign new_n33106 = new_n33095 & new_n33105;
  assign new_n33107 = new_n33106 ^ new_n33093;
  assign new_n33108 = new_n33078 ^ new_n33070;
  assign new_n33109 = new_n33066 ^ new_n33055;
  assign new_n33110 = new_n33109 ^ new_n33108;
  assign new_n33111 = ~new_n33104 & ~new_n33110;
  assign new_n33112 = new_n33111 ^ new_n33084;
  assign new_n33113 = ~new_n33085 & ~new_n33090;
  assign new_n33114 = new_n33055 & new_n33090;
  assign new_n33115 = new_n33114 ^ new_n33113;
  assign new_n33116 = new_n33115 ^ new_n33112;
  assign new_n33117 = new_n33070 ^ new_n33060;
  assign new_n33118 = new_n33104 ^ new_n33085;
  assign new_n33119 = ~new_n33118 & new_n33071;
  assign new_n33120 = ~new_n33072 & new_n33109;
  assign new_n33121 = new_n33120 ^ new_n33119;
  assign new_n33122 = new_n33115 ^ new_n33055;
  assign new_n33123 = new_n33122 ^ new_n33106;
  assign new_n33124 = new_n33123 ^ new_n33121;
  assign new_n33125 = new_n33124 ^ new_n33117;
  assign new_n33126 = new_n33103 ^ new_n33066;
  assign new_n33127 = new_n33126 ^ new_n33084;
  assign new_n33128 = new_n33096 & new_n33127;
  assign new_n33129 = new_n33128 ^ new_n33119;
  assign new_n33130 = new_n33126 ^ new_n33060;
  assign new_n33131 = new_n33130 ^ new_n33129;
  assign new_n33132 = ~new_n33108 & new_n33130;
  assign new_n33133 = new_n33091 ^ new_n33070;
  assign new_n33134 = new_n33127 ^ new_n33090;
  assign new_n33135 = ~new_n33133 & ~new_n33134;
  assign new_n33136 = new_n33135 ^ new_n33132;
  assign new_n33137 = new_n33136 ^ new_n33070;
  assign new_n33138 = new_n33137 ^ new_n33131;
  assign new_n33139 = new_n33132 ^ new_n33093;
  assign new_n33140 = new_n33139 ^ new_n33071;
  assign new_n33141 = new_n33128 ^ new_n33120;
  assign new_n33142 = new_n33102 ^ new_n33060;
  assign new_n33143 = new_n33142 ^ new_n33141;
  assign new_n33144 = new_n33143 ^ new_n33140;
  assign new_n33145 = new_n33112 ^ new_n33104;
  assign new_n33146 = new_n33141 ^ new_n33106;
  assign new_n33147 = new_n33146 ^ new_n33066;
  assign new_n33148 = new_n33147 ^ new_n33145;
  assign new_n33149 = ~new_n33144 & new_n33148;
  assign new_n33150 = new_n33149 ^ new_n33138;
  assign new_n33151 = ~new_n33125 & new_n33150;
  assign new_n33152 = new_n33151 ^ new_n33116;
  assign new_n33153 = new_n33152 ^ new_n33131;
  assign new_n33154 = new_n33149 ^ new_n33116;
  assign new_n33155 = new_n33154 ^ new_n33131;
  assign new_n33156 = new_n33135 ^ new_n33092;
  assign new_n33157 = new_n33156 ^ new_n33121;
  assign new_n33158 = ~new_n33155 & ~new_n33157;
  assign new_n33159 = new_n33158 ^ new_n33149;
  assign new_n33160 = new_n33138 & new_n33159;
  assign new_n33161 = new_n33160 ^ new_n33150;
  assign new_n33162 = ~new_n33153 & new_n33161;
  assign new_n33163 = new_n33162 ^ new_n33160;
  assign new_n33164 = new_n33163 ^ new_n33107;
  assign new_n33165 = new_n33164 ^ new_n33079;
  assign new_n33166 = new_n33165 ^ new_n33055;
  assign new_n33167 = new_n33151 ^ new_n33132;
  assign new_n33168 = new_n33167 ^ new_n33112;
  assign new_n33169 = new_n33168 ^ new_n33166;
  assign new_n33170 = ~new_n33072 & ~new_n33169;
  assign new_n33171 = new_n33158 ^ new_n33151;
  assign new_n33172 = new_n33137 ^ new_n33116;
  assign new_n33173 = new_n33172 ^ new_n33171;
  assign new_n33174 = ~new_n33173 & new_n33127;
  assign new_n33175 = new_n33174 ^ new_n33170;
  assign new_n33176 = new_n33160 ^ new_n33158;
  assign new_n33177 = new_n33176 ^ new_n33157;
  assign new_n33178 = ~new_n33177 & new_n33105;
  assign new_n33179 = new_n33160 ^ new_n33144;
  assign new_n33180 = ~new_n33104 & ~new_n33179;
  assign new_n33181 = new_n33180 ^ new_n33178;
  assign new_n33182 = ~new_n33110 & ~new_n33179;
  assign new_n33183 = new_n33182 ^ new_n33181;
  assign new_n33184 = ~new_n33177 & new_n33095;
  assign new_n33185 = ~new_n33169 & new_n33109;
  assign new_n33186 = ~new_n33173 & new_n33096;
  assign new_n33187 = new_n33186 ^ new_n33185;
  assign new_n33188 = new_n33187 ^ new_n33184;
  assign new_n33189 = new_n33188 ^ new_n33183;
  assign new_n33190 = new_n33189 ^ new_n33175;
  assign new_n33191 = new_n33190 ^ new_n33050;
  assign new_n33192 = new_n33191 ^ new_n32901;
  assign new_n33193 = new_n28114 ^ new_n27978;
  assign new_n33194 = new_n33193 ^ new_n32405;
  assign new_n33195 = new_n33194 ^ new_n27556;
  assign new_n33196 = new_n28029 ^ new_n27707;
  assign new_n33197 = new_n33196 ^ new_n28218;
  assign new_n33198 = new_n33197 ^ new_n33195;
  assign new_n33199 = new_n28188 ^ new_n28064;
  assign new_n33200 = new_n28029 ^ new_n27863;
  assign new_n33201 = new_n33200 ^ new_n32432;
  assign new_n33202 = new_n33201 ^ new_n33199;
  assign new_n33203 = new_n33202 ^ new_n33198;
  assign new_n33204 = new_n28129 ^ new_n28125;
  assign new_n33205 = new_n32456 ^ new_n27978;
  assign new_n33206 = new_n33205 ^ new_n28175;
  assign new_n33207 = new_n33206 ^ new_n33204;
  assign new_n33208 = new_n32297 ^ new_n28229;
  assign new_n33209 = new_n33208 ^ new_n28141;
  assign new_n33210 = new_n33209 ^ new_n28090;
  assign new_n33211 = new_n33210 ^ new_n33207;
  assign new_n33212 = new_n33211 ^ new_n33203;
  assign new_n33213 = new_n33193 ^ new_n30372;
  assign new_n33214 = new_n32381 ^ new_n28080;
  assign new_n33215 = new_n33214 ^ new_n30393;
  assign new_n33216 = new_n33215 ^ new_n33213;
  assign new_n33217 = new_n33216 ^ new_n33202;
  assign new_n33218 = new_n28193 ^ new_n28188;
  assign new_n33219 = new_n32034 ^ new_n28004;
  assign new_n33220 = new_n33219 ^ new_n28125;
  assign new_n33221 = new_n33220 ^ new_n33218;
  assign new_n33222 = new_n33221 ^ new_n33202;
  assign new_n33223 = new_n32393 ^ new_n28198;
  assign new_n33224 = new_n33193 ^ new_n28150;
  assign new_n33225 = new_n33224 ^ new_n33223;
  assign new_n33226 = new_n33225 ^ new_n33222;
  assign new_n33227 = new_n33216 & new_n33226;
  assign new_n33228 = new_n33227 ^ new_n33216;
  assign new_n33229 = new_n33226 ^ new_n33216;
  assign new_n33230 = new_n33229 ^ new_n33211;
  assign new_n33231 = new_n33207 ^ new_n33198;
  assign new_n33232 = new_n28229 ^ new_n27707;
  assign new_n33233 = new_n33232 ^ new_n28095;
  assign new_n33234 = new_n33193 ^ new_n32342;
  assign new_n33235 = new_n33234 ^ new_n28235;
  assign new_n33236 = new_n33235 ^ new_n33233;
  assign new_n33237 = new_n33236 ^ new_n33216;
  assign new_n33238 = new_n33237 ^ new_n33231;
  assign new_n33239 = new_n33238 ^ new_n33225;
  assign new_n33240 = new_n33230 & new_n33239;
  assign new_n33241 = new_n33240 ^ new_n33228;
  assign new_n33242 = new_n33216 ^ new_n33198;
  assign new_n33243 = new_n33242 ^ new_n33211;
  assign new_n33244 = ~new_n33238 & ~new_n33243;
  assign new_n33245 = new_n33244 ^ new_n33221;
  assign new_n33246 = ~new_n33222 & ~new_n33225;
  assign new_n33247 = new_n33198 & new_n33225;
  assign new_n33248 = new_n33247 ^ new_n33246;
  assign new_n33249 = new_n33248 ^ new_n33245;
  assign new_n33250 = new_n33207 ^ new_n33202;
  assign new_n33251 = new_n33238 ^ new_n33222;
  assign new_n33252 = ~new_n33251 & new_n33211;
  assign new_n33253 = new_n33210 ^ new_n33198;
  assign new_n33254 = ~new_n33212 & new_n33253;
  assign new_n33255 = new_n33254 ^ new_n33252;
  assign new_n33256 = new_n33248 ^ new_n33198;
  assign new_n33257 = new_n33256 ^ new_n33240;
  assign new_n33258 = new_n33257 ^ new_n33255;
  assign new_n33259 = new_n33258 ^ new_n33250;
  assign new_n33260 = new_n33237 ^ new_n33210;
  assign new_n33261 = new_n33260 ^ new_n33221;
  assign new_n33262 = new_n33231 & new_n33261;
  assign new_n33263 = new_n33262 ^ new_n33252;
  assign new_n33264 = new_n33260 ^ new_n33202;
  assign new_n33265 = new_n33264 ^ new_n33263;
  assign new_n33266 = new_n33226 ^ new_n33207;
  assign new_n33267 = new_n33261 ^ new_n33225;
  assign new_n33268 = ~new_n33266 & ~new_n33267;
  assign new_n33269 = new_n33216 ^ new_n33207;
  assign new_n33270 = ~new_n33269 & new_n33264;
  assign new_n33271 = new_n33270 ^ new_n33268;
  assign new_n33272 = new_n33271 ^ new_n33207;
  assign new_n33273 = new_n33272 ^ new_n33265;
  assign new_n33274 = new_n33270 ^ new_n33228;
  assign new_n33275 = new_n33274 ^ new_n33211;
  assign new_n33276 = new_n33262 ^ new_n33254;
  assign new_n33277 = new_n33236 ^ new_n33202;
  assign new_n33278 = new_n33277 ^ new_n33276;
  assign new_n33279 = new_n33278 ^ new_n33275;
  assign new_n33280 = new_n33245 ^ new_n33238;
  assign new_n33281 = new_n33276 ^ new_n33240;
  assign new_n33282 = new_n33281 ^ new_n33210;
  assign new_n33283 = new_n33282 ^ new_n33280;
  assign new_n33284 = ~new_n33279 & new_n33283;
  assign new_n33285 = new_n33284 ^ new_n33273;
  assign new_n33286 = ~new_n33259 & new_n33285;
  assign new_n33287 = new_n33286 ^ new_n33249;
  assign new_n33288 = new_n33287 ^ new_n33265;
  assign new_n33289 = new_n33284 ^ new_n33249;
  assign new_n33290 = new_n33289 ^ new_n33265;
  assign new_n33291 = new_n33268 ^ new_n33227;
  assign new_n33292 = new_n33291 ^ new_n33255;
  assign new_n33293 = ~new_n33290 & ~new_n33292;
  assign new_n33294 = new_n33293 ^ new_n33284;
  assign new_n33295 = new_n33273 & new_n33294;
  assign new_n33296 = new_n33295 ^ new_n33285;
  assign new_n33297 = ~new_n33288 & new_n33296;
  assign new_n33298 = new_n33297 ^ new_n33295;
  assign new_n33299 = new_n33298 ^ new_n33241;
  assign new_n33300 = new_n33299 ^ new_n33217;
  assign new_n33301 = new_n33300 ^ new_n33198;
  assign new_n33302 = new_n33286 ^ new_n33270;
  assign new_n33303 = new_n33302 ^ new_n33245;
  assign new_n33304 = new_n33303 ^ new_n33301;
  assign new_n33305 = ~new_n33212 & ~new_n33304;
  assign new_n33306 = new_n33293 ^ new_n33286;
  assign new_n33307 = new_n33272 ^ new_n33249;
  assign new_n33308 = new_n33307 ^ new_n33306;
  assign new_n33309 = ~new_n33308 & new_n33261;
  assign new_n33310 = new_n33309 ^ new_n33305;
  assign new_n33311 = new_n33295 ^ new_n33293;
  assign new_n33312 = new_n33311 ^ new_n33292;
  assign new_n33313 = ~new_n33312 & new_n33239;
  assign new_n33314 = new_n33295 ^ new_n33279;
  assign new_n33315 = ~new_n33238 & ~new_n33314;
  assign new_n33316 = new_n33315 ^ new_n33313;
  assign new_n33317 = ~new_n33243 & ~new_n33314;
  assign new_n33318 = new_n33317 ^ new_n33316;
  assign new_n33319 = ~new_n33312 & new_n33230;
  assign new_n33320 = ~new_n33308 & new_n33231;
  assign new_n33321 = ~new_n33304 & new_n33253;
  assign new_n33322 = new_n33321 ^ new_n33320;
  assign new_n33323 = new_n33322 ^ new_n33319;
  assign new_n33324 = new_n33323 ^ new_n33318;
  assign new_n33325 = new_n33324 ^ new_n33310;
  assign new_n33326 = new_n33325 ^ new_n29964;
  assign new_n33327 = new_n33320 ^ new_n33309;
  assign new_n33328 = new_n33293 ^ new_n33207;
  assign new_n33329 = new_n33268 ^ new_n33256;
  assign new_n33330 = new_n33329 ^ new_n33300;
  assign new_n33331 = new_n33330 ^ new_n33328;
  assign new_n33332 = new_n33211 & new_n33331;
  assign new_n33333 = ~new_n33266 & ~new_n33288;
  assign new_n33334 = ~new_n33251 & new_n33331;
  assign new_n33335 = new_n33334 ^ new_n33333;
  assign new_n33336 = new_n33293 ^ new_n33273;
  assign new_n33337 = ~new_n33225 & new_n33336;
  assign new_n33338 = new_n33337 ^ new_n33315;
  assign new_n33339 = new_n33297 ^ new_n33286;
  assign new_n33340 = new_n33339 ^ new_n33283;
  assign new_n33341 = ~new_n33269 & new_n33340;
  assign new_n33342 = new_n33341 ^ new_n33338;
  assign new_n33343 = new_n33342 ^ new_n33335;
  assign new_n33344 = new_n33343 ^ new_n33332;
  assign new_n33345 = new_n33344 ^ new_n33327;
  assign new_n33346 = new_n33345 ^ new_n33326;
  assign new_n33347 = new_n33346 ^ new_n33192;
  assign new_n33348 = new_n32892 ^ new_n32888;
  assign new_n33349 = new_n32883 ^ new_n32813;
  assign new_n33350 = new_n32856 ^ new_n32805;
  assign new_n33351 = new_n33350 ^ new_n32828;
  assign new_n33352 = new_n33351 ^ new_n33349;
  assign new_n33353 = ~new_n33352 & new_n32815;
  assign new_n33354 = new_n32879 ^ new_n32855;
  assign new_n33355 = ~new_n32796 & new_n33354;
  assign new_n33356 = new_n33355 ^ new_n33353;
  assign new_n33357 = new_n32843 & new_n32875;
  assign new_n33358 = new_n32831 & new_n33354;
  assign new_n33359 = new_n33358 ^ new_n33357;
  assign new_n33360 = ~new_n33352 & new_n32816;
  assign new_n33361 = new_n33360 ^ new_n32868;
  assign new_n33362 = new_n33361 ^ new_n33359;
  assign new_n33363 = new_n33362 ^ new_n33356;
  assign new_n33364 = new_n33363 ^ new_n33348;
  assign new_n33365 = new_n33158 ^ new_n33138;
  assign new_n33366 = new_n33091 ^ new_n33055;
  assign new_n33367 = ~new_n33366 & new_n33365;
  assign new_n33368 = new_n33162 ^ new_n33151;
  assign new_n33369 = new_n33368 ^ new_n33148;
  assign new_n33370 = new_n33130 & new_n33369;
  assign new_n33371 = new_n33162 ^ new_n33125;
  assign new_n33372 = ~new_n33091 & ~new_n33371;
  assign new_n33373 = new_n33372 ^ new_n33188;
  assign new_n33374 = new_n33373 ^ new_n33370;
  assign new_n33375 = new_n33374 ^ new_n33170;
  assign new_n33376 = new_n33375 ^ new_n33367;
  assign new_n33377 = ~new_n33090 & new_n33365;
  assign new_n33378 = new_n33377 ^ new_n33180;
  assign new_n33379 = ~new_n33108 & new_n33369;
  assign new_n33380 = new_n33379 ^ new_n33378;
  assign new_n33381 = ~new_n33133 & ~new_n33153;
  assign new_n33382 = new_n33158 ^ new_n33070;
  assign new_n33383 = new_n33135 ^ new_n33122;
  assign new_n33384 = new_n33383 ^ new_n33165;
  assign new_n33385 = new_n33384 ^ new_n33382;
  assign new_n33386 = ~new_n33118 & new_n33385;
  assign new_n33387 = new_n33386 ^ new_n33381;
  assign new_n33388 = new_n33387 ^ new_n33380;
  assign new_n33389 = new_n33388 ^ new_n33376;
  assign new_n33390 = new_n33018 ^ new_n32998;
  assign new_n33391 = new_n32950 ^ new_n32908;
  assign new_n33392 = ~new_n33391 & new_n33390;
  assign new_n33393 = new_n33022 ^ new_n33011;
  assign new_n33394 = new_n33393 ^ new_n33008;
  assign new_n33395 = new_n32990 & new_n33394;
  assign new_n33396 = new_n33022 ^ new_n32985;
  assign new_n33397 = ~new_n32950 & ~new_n33396;
  assign new_n33398 = new_n33397 ^ new_n33048;
  assign new_n33399 = new_n33398 ^ new_n33395;
  assign new_n33400 = new_n33399 ^ new_n33030;
  assign new_n33401 = new_n33400 ^ new_n33392;
  assign new_n33402 = ~new_n32949 & new_n33390;
  assign new_n33403 = new_n33402 ^ new_n33040;
  assign new_n33404 = ~new_n32968 & new_n33394;
  assign new_n33405 = new_n33404 ^ new_n33403;
  assign new_n33406 = ~new_n32993 & ~new_n33013;
  assign new_n33407 = new_n33018 ^ new_n32927;
  assign new_n33408 = new_n32995 ^ new_n32982;
  assign new_n33409 = new_n33408 ^ new_n33025;
  assign new_n33410 = new_n33409 ^ new_n33407;
  assign new_n33411 = ~new_n32978 & new_n33410;
  assign new_n33412 = new_n33411 ^ new_n33406;
  assign new_n33413 = new_n33412 ^ new_n33405;
  assign new_n33414 = new_n33413 ^ new_n33401;
  assign new_n33415 = new_n33414 ^ new_n33389;
  assign new_n33416 = new_n33415 ^ new_n33364;
  assign new_n33417 = new_n33226 ^ new_n33198;
  assign new_n33418 = ~new_n33417 & new_n33336;
  assign new_n33419 = new_n33297 ^ new_n33259;
  assign new_n33420 = ~new_n33226 & ~new_n33419;
  assign new_n33421 = new_n33420 ^ new_n33323;
  assign new_n33422 = new_n33264 & new_n33340;
  assign new_n33423 = new_n33422 ^ new_n33421;
  assign new_n33424 = new_n33423 ^ new_n33305;
  assign new_n33425 = new_n33424 ^ new_n33418;
  assign new_n33426 = new_n33425 ^ new_n33343;
  assign new_n33427 = new_n33426 ^ new_n29990;
  assign new_n33428 = new_n33341 ^ new_n33334;
  assign new_n33429 = ~new_n33267 & ~new_n33288;
  assign new_n33430 = ~new_n33419 & new_n33229;
  assign new_n33431 = new_n33430 ^ new_n33429;
  assign new_n33432 = new_n33431 ^ new_n33322;
  assign new_n33433 = new_n33420 ^ new_n33305;
  assign new_n33434 = new_n33433 ^ new_n33432;
  assign new_n33435 = new_n33434 ^ new_n33428;
  assign new_n33436 = new_n33435 ^ new_n33427;
  assign new_n33437 = new_n33436 ^ new_n33416;
  assign new_n33438 = ~new_n33134 & ~new_n33153;
  assign new_n33439 = new_n33438 ^ new_n33182;
  assign new_n33440 = new_n33377 ^ new_n33178;
  assign new_n33441 = new_n33440 ^ new_n33373;
  assign new_n33442 = new_n33441 ^ new_n33439;
  assign new_n33443 = ~new_n32994 & ~new_n33013;
  assign new_n33444 = new_n33443 ^ new_n33042;
  assign new_n33445 = new_n33402 ^ new_n33038;
  assign new_n33446 = new_n33445 ^ new_n33398;
  assign new_n33447 = new_n33446 ^ new_n33444;
  assign new_n33448 = new_n33447 ^ new_n33442;
  assign new_n33449 = new_n33448 ^ new_n29996;
  assign new_n33450 = new_n32880 ^ new_n32863;
  assign new_n33451 = new_n33450 ^ new_n32862;
  assign new_n33452 = ~new_n32832 & ~new_n33451;
  assign new_n33453 = new_n33452 ^ new_n33361;
  assign new_n33454 = new_n33453 ^ new_n33355;
  assign new_n33455 = ~new_n32799 & new_n32891;
  assign new_n33456 = new_n33455 ^ new_n33454;
  assign new_n33457 = new_n33456 ^ new_n33353;
  assign new_n33458 = ~new_n32895 & new_n32826;
  assign new_n33459 = new_n33458 ^ new_n32867;
  assign new_n33460 = new_n33459 ^ new_n33457;
  assign new_n33461 = new_n33317 ^ new_n33309;
  assign new_n33462 = new_n33461 ^ new_n33424;
  assign new_n33463 = new_n33462 ^ new_n33460;
  assign new_n33464 = new_n33463 ^ new_n33449;
  assign new_n33465 = ~new_n32850 & new_n32893;
  assign new_n33466 = new_n33465 ^ new_n33457;
  assign new_n33467 = new_n33466 ^ new_n32899;
  assign new_n33468 = new_n33429 ^ new_n33317;
  assign new_n33469 = new_n33337 ^ new_n33313;
  assign new_n33470 = new_n33469 ^ new_n33421;
  assign new_n33471 = new_n33470 ^ new_n33468;
  assign new_n33472 = new_n33471 ^ new_n33467;
  assign new_n33473 = new_n33472 ^ new_n33426;
  assign new_n33474 = new_n33473 ^ new_n33464;
  assign new_n33475 = new_n33455 ^ new_n32898;
  assign new_n33476 = new_n33475 ^ new_n33362;
  assign new_n33477 = new_n33476 ^ new_n33463;
  assign new_n33478 = new_n33411 ^ new_n33404;
  assign new_n33479 = ~new_n33396 & new_n32953;
  assign new_n33480 = new_n33479 ^ new_n33443;
  assign new_n33481 = new_n33480 ^ new_n33047;
  assign new_n33482 = new_n33397 ^ new_n33030;
  assign new_n33483 = new_n33482 ^ new_n33481;
  assign new_n33484 = new_n33483 ^ new_n33478;
  assign new_n33485 = new_n33386 ^ new_n33379;
  assign new_n33486 = ~new_n33371 & new_n33094;
  assign new_n33487 = new_n33486 ^ new_n33438;
  assign new_n33488 = new_n33487 ^ new_n33187;
  assign new_n33489 = new_n33372 ^ new_n33170;
  assign new_n33490 = new_n33489 ^ new_n33488;
  assign new_n33491 = new_n33490 ^ new_n33485;
  assign new_n33492 = new_n33491 ^ new_n33484;
  assign new_n33493 = new_n33492 ^ new_n33477;
  assign new_n33494 = new_n33422 ^ new_n33342;
  assign new_n33495 = new_n33494 ^ new_n33432;
  assign new_n33496 = new_n33435 ^ new_n30004;
  assign new_n33497 = new_n33496 ^ new_n33495;
  assign new_n33498 = new_n33497 ^ new_n33493;
  assign new_n33499 = new_n33498 ^ new_n33474;
  assign new_n33500 = new_n33499 ^ new_n33437;
  assign new_n33501 = new_n33500 ^ new_n33347;
  assign new_n33502 = new_n33495 ^ new_n30010;
  assign new_n33503 = new_n33405 ^ new_n33395;
  assign new_n33504 = new_n33503 ^ new_n33481;
  assign new_n33505 = new_n33380 ^ new_n33370;
  assign new_n33506 = new_n33505 ^ new_n33488;
  assign new_n33507 = new_n33506 ^ new_n33504;
  assign new_n33508 = new_n33507 ^ new_n33463;
  assign new_n33509 = new_n33508 ^ new_n33502;
  assign new_n33510 = new_n33463 ^ new_n30012;
  assign new_n33511 = new_n33374 ^ new_n33183;
  assign new_n33512 = new_n33399 ^ new_n33043;
  assign new_n33513 = new_n33512 ^ new_n33511;
  assign new_n33514 = new_n33513 ^ new_n33510;
  assign new_n33515 = new_n33458 ^ new_n33357;
  assign new_n33516 = ~new_n33451 & new_n32830;
  assign new_n33517 = new_n33516 ^ new_n32894;
  assign new_n33518 = new_n33517 ^ new_n33454;
  assign new_n33519 = new_n33518 ^ new_n33515;
  assign new_n33520 = new_n33423 ^ new_n33318;
  assign new_n33521 = new_n33520 ^ new_n33519;
  assign new_n33522 = new_n33521 ^ new_n33471;
  assign new_n33523 = new_n33522 ^ new_n33514;
  assign new_n33524 = new_n33046 ^ new_n33034;
  assign new_n33525 = new_n32928 & new_n33410;
  assign new_n33526 = new_n33525 ^ new_n33413;
  assign new_n33527 = new_n33526 ^ new_n33524;
  assign new_n33528 = new_n33186 ^ new_n33174;
  assign new_n33529 = new_n33071 & new_n33385;
  assign new_n33530 = new_n33529 ^ new_n33388;
  assign new_n33531 = new_n33530 ^ new_n33528;
  assign new_n33532 = new_n33531 ^ new_n33527;
  assign new_n33533 = new_n33532 ^ new_n33345;
  assign new_n33534 = new_n33516 ^ new_n32896;
  assign new_n33535 = new_n33534 ^ new_n33458;
  assign new_n33536 = new_n33535 ^ new_n33456;
  assign new_n33537 = new_n33536 ^ new_n33520;
  assign new_n33538 = new_n33537 ^ new_n30017;
  assign new_n33539 = new_n33538 ^ new_n33533;
  assign new_n33540 = new_n33539 ^ new_n33347;
  assign new_n33541 = new_n33540 ^ new_n33509;
  assign new_n33542 = new_n33541 ^ new_n33523;
  assign new_n33543 = new_n33509 & new_n33542;
  assign new_n33544 = new_n33543 ^ new_n33523;
  assign new_n33545 = new_n33353 ^ new_n32867;
  assign new_n33546 = new_n33535 ^ new_n33453;
  assign new_n33547 = new_n33546 ^ new_n33545;
  assign new_n33548 = new_n33182 ^ new_n33174;
  assign new_n33549 = new_n33548 ^ new_n33375;
  assign new_n33550 = new_n33042 ^ new_n33034;
  assign new_n33551 = new_n33550 ^ new_n33400;
  assign new_n33552 = new_n33551 ^ new_n33549;
  assign new_n33553 = new_n33552 ^ new_n33547;
  assign new_n33554 = new_n33462 ^ new_n30025;
  assign new_n33555 = new_n33554 ^ new_n33325;
  assign new_n33556 = new_n33555 ^ new_n33553;
  assign new_n33557 = new_n33556 ^ new_n33523;
  assign new_n33558 = new_n33557 ^ new_n33499;
  assign new_n33559 = new_n33523 ^ new_n33498;
  assign new_n33560 = new_n33556 ^ new_n33437;
  assign new_n33561 = new_n33560 ^ new_n33559;
  assign new_n33562 = ~new_n33561 & new_n33558;
  assign new_n33563 = new_n33562 ^ new_n33347;
  assign new_n33564 = new_n33563 ^ new_n33544;
  assign new_n33565 = ~new_n33541 & new_n33498;
  assign new_n33566 = new_n33565 ^ new_n33498;
  assign new_n33567 = new_n33539 ^ new_n33500;
  assign new_n33568 = new_n33556 ^ new_n33498;
  assign new_n33569 = ~new_n33568 & new_n33567;
  assign new_n33570 = new_n33569 ^ new_n33566;
  assign new_n33571 = new_n33570 ^ new_n33560;
  assign new_n33572 = new_n33501 & new_n33557;
  assign new_n33573 = new_n33539 ^ new_n33523;
  assign new_n33574 = new_n33573 ^ new_n33560;
  assign new_n33575 = new_n33523 ^ new_n33437;
  assign new_n33576 = new_n33574 & new_n33575;
  assign new_n33577 = new_n33576 ^ new_n33572;
  assign new_n33578 = new_n33539 ^ new_n33474;
  assign new_n33579 = new_n33578 ^ new_n33577;
  assign new_n33580 = new_n33579 ^ new_n33571;
  assign new_n33581 = new_n33563 ^ new_n33558;
  assign new_n33582 = new_n33541 ^ new_n33498;
  assign new_n33583 = new_n33582 ^ new_n33560;
  assign new_n33584 = new_n33558 ^ new_n33509;
  assign new_n33585 = ~new_n33583 & new_n33584;
  assign new_n33586 = new_n33585 ^ new_n33572;
  assign new_n33587 = new_n33576 ^ new_n33437;
  assign new_n33588 = new_n33587 ^ new_n33586;
  assign new_n33589 = new_n33588 ^ new_n33581;
  assign new_n33590 = ~new_n33580 & new_n33589;
  assign new_n33591 = new_n33590 ^ new_n33564;
  assign new_n33592 = new_n33558 ^ new_n33540;
  assign new_n33593 = new_n33560 & new_n33592;
  assign new_n33594 = new_n33593 ^ new_n33572;
  assign new_n33595 = new_n33594 ^ new_n33567;
  assign new_n33596 = new_n33595 ^ new_n33591;
  assign new_n33597 = new_n33556 ^ new_n33541;
  assign new_n33598 = new_n33509 ^ new_n33501;
  assign new_n33599 = new_n33597 & new_n33598;
  assign new_n33600 = new_n33599 ^ new_n33565;
  assign new_n33601 = new_n33593 ^ new_n33576;
  assign new_n33602 = new_n33601 ^ new_n33600;
  assign new_n33603 = ~new_n33602 & new_n33596;
  assign new_n33604 = new_n33556 ^ new_n33539;
  assign new_n33605 = new_n33585 ^ new_n33543;
  assign new_n33606 = new_n33605 ^ new_n33601;
  assign new_n33607 = new_n33606 ^ new_n33604;
  assign new_n33608 = new_n33599 ^ new_n33569;
  assign new_n33609 = new_n33608 ^ new_n33556;
  assign new_n33610 = new_n33609 ^ new_n33595;
  assign new_n33611 = new_n33610 ^ new_n33590;
  assign new_n33612 = new_n33607 & new_n33611;
  assign new_n33613 = new_n33612 ^ new_n33603;
  assign new_n33614 = new_n33609 ^ new_n33564;
  assign new_n33615 = new_n33614 ^ new_n33613;
  assign new_n33616 = new_n33501 & new_n33615;
  assign new_n33617 = new_n33603 ^ new_n33590;
  assign new_n33618 = new_n33610 & new_n33617;
  assign new_n33619 = new_n33618 ^ new_n33580;
  assign new_n33620 = ~new_n33561 & ~new_n33619;
  assign new_n33621 = new_n33620 ^ new_n33616;
  assign new_n33622 = new_n33539 ^ new_n33498;
  assign new_n33623 = new_n33585 ^ new_n33566;
  assign new_n33624 = new_n33612 ^ new_n33564;
  assign new_n33625 = new_n33624 ^ new_n33595;
  assign new_n33626 = new_n33618 ^ new_n33611;
  assign new_n33627 = new_n33625 & new_n33626;
  assign new_n33628 = new_n33627 ^ new_n33618;
  assign new_n33629 = new_n33628 ^ new_n33623;
  assign new_n33630 = new_n33629 ^ new_n33622;
  assign new_n33631 = new_n33630 ^ new_n33523;
  assign new_n33632 = new_n33612 ^ new_n33569;
  assign new_n33633 = new_n33632 ^ new_n33563;
  assign new_n33634 = new_n33633 ^ new_n33631;
  assign new_n33635 = ~new_n33634 & new_n33574;
  assign new_n33636 = new_n33627 ^ new_n33607;
  assign new_n33637 = new_n33541 & new_n33636;
  assign new_n33638 = new_n33618 ^ new_n33603;
  assign new_n33639 = new_n33638 ^ new_n33602;
  assign new_n33640 = ~new_n33583 & ~new_n33639;
  assign new_n33641 = ~new_n33634 & new_n33575;
  assign new_n33642 = new_n33557 & new_n33615;
  assign new_n33643 = new_n33642 ^ new_n33641;
  assign new_n33644 = new_n33643 ^ new_n33640;
  assign new_n33645 = new_n33644 ^ new_n33637;
  assign new_n33646 = new_n33627 ^ new_n33612;
  assign new_n33647 = new_n33646 ^ new_n33589;
  assign new_n33648 = new_n33567 & new_n33647;
  assign new_n33649 = new_n33648 ^ new_n33645;
  assign new_n33650 = new_n33649 ^ new_n33635;
  assign new_n33651 = new_n33650 ^ new_n33621;
  assign new_n33652 = new_n32033 ^ new_n17564;
  assign new_n33653 = new_n32296 ^ new_n17556;
  assign new_n33654 = new_n32341 ^ new_n17525;
  assign new_n33655 = new_n32380 ^ new_n17542;
  assign new_n33656 = new_n33655 ^ new_n33654;
  assign new_n33657 = new_n33656 ^ new_n33653;
  assign new_n33658 = new_n33657 ^ new_n33652;
  assign new_n33659 = new_n32392 ^ new_n17581;
  assign new_n33660 = new_n32404 ^ new_n17576;
  assign new_n33661 = new_n32431 ^ new_n17573;
  assign new_n33662 = new_n33661 ^ new_n33652;
  assign new_n33663 = new_n33662 ^ new_n33659;
  assign new_n33664 = new_n33663 ^ new_n33660;
  assign new_n33665 = ~new_n33659 & ~new_n33664;
  assign new_n33666 = new_n33665 ^ new_n33660;
  assign new_n33667 = new_n32455 ^ new_n17568;
  assign new_n33668 = new_n33667 ^ new_n33660;
  assign new_n33669 = new_n33668 ^ new_n33656;
  assign new_n33670 = new_n33660 ^ new_n33655;
  assign new_n33671 = new_n33667 ^ new_n33653;
  assign new_n33672 = new_n33671 ^ new_n33670;
  assign new_n33673 = ~new_n33669 & ~new_n33672;
  assign new_n33674 = new_n33673 ^ new_n33652;
  assign new_n33675 = new_n33674 ^ new_n33666;
  assign new_n33676 = new_n33655 & new_n33663;
  assign new_n33677 = new_n33676 ^ new_n33655;
  assign new_n33678 = new_n33661 ^ new_n33657;
  assign new_n33679 = new_n33667 ^ new_n33655;
  assign new_n33680 = ~new_n33679 & new_n33678;
  assign new_n33681 = new_n33680 ^ new_n33677;
  assign new_n33682 = new_n33681 ^ new_n33671;
  assign new_n33683 = new_n33658 & new_n33668;
  assign new_n33684 = new_n33661 ^ new_n33660;
  assign new_n33685 = new_n33684 ^ new_n33671;
  assign new_n33686 = new_n33660 ^ new_n33653;
  assign new_n33687 = ~new_n33685 & new_n33686;
  assign new_n33688 = new_n33687 ^ new_n33683;
  assign new_n33689 = new_n33661 ^ new_n33654;
  assign new_n33690 = new_n33689 ^ new_n33688;
  assign new_n33691 = new_n33690 ^ new_n33682;
  assign new_n33692 = new_n33674 ^ new_n33669;
  assign new_n33693 = new_n33663 ^ new_n33655;
  assign new_n33694 = new_n33693 ^ new_n33671;
  assign new_n33695 = new_n33669 ^ new_n33659;
  assign new_n33696 = new_n33694 & new_n33695;
  assign new_n33697 = new_n33696 ^ new_n33653;
  assign new_n33698 = new_n33697 ^ new_n33688;
  assign new_n33699 = new_n33698 ^ new_n33692;
  assign new_n33700 = ~new_n33691 & new_n33699;
  assign new_n33701 = new_n33700 ^ new_n33675;
  assign new_n33702 = new_n33669 ^ new_n33662;
  assign new_n33703 = ~new_n33702 & new_n33671;
  assign new_n33704 = new_n33703 ^ new_n33683;
  assign new_n33705 = new_n33704 ^ new_n33678;
  assign new_n33706 = new_n33705 ^ new_n33701;
  assign new_n33707 = new_n33667 ^ new_n33663;
  assign new_n33708 = new_n33659 ^ new_n33658;
  assign new_n33709 = ~new_n33707 & ~new_n33708;
  assign new_n33710 = new_n33709 ^ new_n33676;
  assign new_n33711 = new_n33703 ^ new_n33687;
  assign new_n33712 = new_n33711 ^ new_n33710;
  assign new_n33713 = ~new_n33706 & ~new_n33712;
  assign new_n33714 = new_n33667 ^ new_n33661;
  assign new_n33715 = new_n33696 ^ new_n33665;
  assign new_n33716 = new_n33715 ^ new_n33711;
  assign new_n33717 = new_n33716 ^ new_n33714;
  assign new_n33718 = new_n33709 ^ new_n33680;
  assign new_n33719 = new_n33718 ^ new_n33667;
  assign new_n33720 = new_n33719 ^ new_n33705;
  assign new_n33721 = new_n33720 ^ new_n33700;
  assign new_n33722 = ~new_n33717 & new_n33721;
  assign new_n33723 = new_n33722 ^ new_n33713;
  assign new_n33724 = new_n33719 ^ new_n33675;
  assign new_n33725 = new_n33724 ^ new_n33723;
  assign new_n33726 = ~new_n33725 & new_n33658;
  assign new_n33727 = new_n33713 ^ new_n33700;
  assign new_n33728 = new_n33720 & new_n33727;
  assign new_n33729 = new_n33728 ^ new_n33691;
  assign new_n33730 = ~new_n33672 & ~new_n33729;
  assign new_n33731 = new_n33730 ^ new_n33726;
  assign new_n33732 = new_n33661 ^ new_n33655;
  assign new_n33733 = new_n33696 ^ new_n33677;
  assign new_n33734 = new_n33722 ^ new_n33675;
  assign new_n33735 = new_n33734 ^ new_n33705;
  assign new_n33736 = new_n33728 ^ new_n33721;
  assign new_n33737 = ~new_n33735 & new_n33736;
  assign new_n33738 = new_n33737 ^ new_n33728;
  assign new_n33739 = new_n33738 ^ new_n33733;
  assign new_n33740 = new_n33739 ^ new_n33732;
  assign new_n33741 = new_n33740 ^ new_n33660;
  assign new_n33742 = new_n33722 ^ new_n33680;
  assign new_n33743 = new_n33742 ^ new_n33674;
  assign new_n33744 = new_n33743 ^ new_n33741;
  assign new_n33745 = ~new_n33685 & ~new_n33744;
  assign new_n33746 = new_n33737 ^ new_n33717;
  assign new_n33747 = ~new_n33663 & ~new_n33746;
  assign new_n33748 = new_n33728 ^ new_n33713;
  assign new_n33749 = new_n33748 ^ new_n33712;
  assign new_n33750 = ~new_n33749 & new_n33694;
  assign new_n33751 = ~new_n33744 & new_n33686;
  assign new_n33752 = ~new_n33725 & new_n33668;
  assign new_n33753 = new_n33752 ^ new_n33751;
  assign new_n33754 = new_n33753 ^ new_n33750;
  assign new_n33755 = new_n33754 ^ new_n33747;
  assign new_n33756 = new_n33737 ^ new_n33722;
  assign new_n33757 = new_n33756 ^ new_n33699;
  assign new_n33758 = new_n33678 & new_n33757;
  assign new_n33759 = new_n33758 ^ new_n33755;
  assign new_n33760 = new_n33759 ^ new_n33745;
  assign new_n33761 = new_n33760 ^ new_n33731;
  assign new_n33762 = new_n33761 ^ new_n21077;
  assign new_n33763 = new_n33762 ^ new_n33651;
  assign new_n33764 = new_n33745 ^ new_n33726;
  assign new_n33765 = ~new_n33669 & ~new_n33729;
  assign new_n33766 = ~new_n33749 & new_n33695;
  assign new_n33767 = new_n33766 ^ new_n33765;
  assign new_n33768 = new_n33767 ^ new_n33730;
  assign new_n33769 = new_n33768 ^ new_n33754;
  assign new_n33770 = new_n33769 ^ new_n33764;
  assign new_n33771 = new_n33770 ^ new_n21074;
  assign new_n33772 = new_n33635 ^ new_n33616;
  assign new_n33773 = ~new_n33619 & new_n33558;
  assign new_n33774 = ~new_n33639 & new_n33584;
  assign new_n33775 = new_n33774 ^ new_n33773;
  assign new_n33776 = new_n33775 ^ new_n33620;
  assign new_n33777 = new_n33776 ^ new_n33644;
  assign new_n33778 = new_n33777 ^ new_n33772;
  assign new_n33779 = new_n33778 ^ new_n33771;
  assign new_n33780 = new_n33752 ^ new_n33726;
  assign new_n33781 = new_n33713 ^ new_n33667;
  assign new_n33782 = new_n33709 ^ new_n33665;
  assign new_n33783 = new_n33782 ^ new_n33740;
  assign new_n33784 = new_n33783 ^ new_n33781;
  assign new_n33785 = new_n33671 & new_n33784;
  assign new_n33786 = ~new_n33679 & new_n33757;
  assign new_n33787 = new_n33720 ^ new_n33713;
  assign new_n33788 = ~new_n33659 & new_n33787;
  assign new_n33789 = new_n33788 ^ new_n33765;
  assign new_n33790 = new_n33789 ^ new_n33786;
  assign new_n33791 = ~new_n33702 & new_n33784;
  assign new_n33792 = ~new_n33707 & ~new_n33735;
  assign new_n33793 = new_n33792 ^ new_n33791;
  assign new_n33794 = new_n33793 ^ new_n33790;
  assign new_n33795 = new_n33794 ^ new_n33785;
  assign new_n33796 = new_n33795 ^ new_n33780;
  assign new_n33797 = new_n33796 ^ new_n21075;
  assign new_n33798 = new_n33642 ^ new_n33616;
  assign new_n33799 = new_n33603 ^ new_n33556;
  assign new_n33800 = new_n33599 ^ new_n33543;
  assign new_n33801 = new_n33800 ^ new_n33630;
  assign new_n33802 = new_n33801 ^ new_n33799;
  assign new_n33803 = ~new_n33802 & new_n33560;
  assign new_n33804 = ~new_n33568 & new_n33647;
  assign new_n33805 = new_n33610 ^ new_n33603;
  assign new_n33806 = new_n33509 & new_n33805;
  assign new_n33807 = new_n33806 ^ new_n33773;
  assign new_n33808 = new_n33807 ^ new_n33804;
  assign new_n33809 = ~new_n33802 & new_n33592;
  assign new_n33810 = new_n33597 & new_n33625;
  assign new_n33811 = new_n33810 ^ new_n33809;
  assign new_n33812 = new_n33811 ^ new_n33808;
  assign new_n33813 = new_n33812 ^ new_n33803;
  assign new_n33814 = new_n33813 ^ new_n33798;
  assign new_n33815 = new_n33814 ^ new_n33797;
  assign new_n33816 = new_n33776 ^ new_n33649;
  assign new_n33817 = new_n33768 ^ new_n33759;
  assign new_n33818 = new_n33817 ^ new_n21078;
  assign new_n33819 = new_n33818 ^ new_n33816;
  assign new_n33820 = new_n33598 & new_n33625;
  assign new_n33821 = new_n33820 ^ new_n33620;
  assign new_n33822 = new_n33806 ^ new_n33774;
  assign new_n33823 = new_n33822 ^ new_n33645;
  assign new_n33824 = new_n33823 ^ new_n33821;
  assign new_n33825 = ~new_n33708 & ~new_n33735;
  assign new_n33826 = new_n33825 ^ new_n33730;
  assign new_n33827 = new_n33788 ^ new_n33766;
  assign new_n33828 = new_n33827 ^ new_n33755;
  assign new_n33829 = new_n33828 ^ new_n33826;
  assign new_n33830 = new_n33829 ^ new_n21081;
  assign new_n33831 = new_n33830 ^ new_n33824;
  assign new_n33832 = new_n33542 & new_n33805;
  assign new_n33833 = new_n33832 ^ new_n33650;
  assign new_n33834 = new_n33833 ^ new_n33812;
  assign new_n33835 = ~new_n33664 & new_n33787;
  assign new_n33836 = new_n33835 ^ new_n33760;
  assign new_n33837 = new_n33836 ^ new_n33794;
  assign new_n33838 = new_n33837 ^ new_n21091;
  assign new_n33839 = new_n33838 ^ new_n33834;
  assign new_n33840 = new_n33791 ^ new_n33786;
  assign new_n33841 = ~new_n33746 & new_n33693;
  assign new_n33842 = new_n33841 ^ new_n33825;
  assign new_n33843 = new_n33842 ^ new_n33753;
  assign new_n33844 = new_n33747 ^ new_n33745;
  assign new_n33845 = new_n33844 ^ new_n33843;
  assign new_n33846 = new_n33845 ^ new_n33840;
  assign new_n33847 = new_n33846 ^ new_n21080;
  assign new_n33848 = new_n33809 ^ new_n33804;
  assign new_n33849 = ~new_n33582 & new_n33636;
  assign new_n33850 = new_n33849 ^ new_n33820;
  assign new_n33851 = new_n33850 ^ new_n33643;
  assign new_n33852 = new_n33637 ^ new_n33635;
  assign new_n33853 = new_n33852 ^ new_n33851;
  assign new_n33854 = new_n33853 ^ new_n33848;
  assign new_n33855 = new_n33854 ^ new_n33847;
  assign new_n33856 = new_n33790 ^ new_n33758;
  assign new_n33857 = new_n33856 ^ new_n33843;
  assign new_n33858 = new_n33857 ^ new_n21085;
  assign new_n33859 = new_n33808 ^ new_n33648;
  assign new_n33860 = new_n33859 ^ new_n33851;
  assign new_n33861 = new_n33860 ^ new_n33858;
  assign new_n33862 = new_n31195 ^ new_n30940;
  assign new_n33863 = new_n33862 ^ new_n30507;
  assign new_n33864 = new_n28753 ^ new_n28590;
  assign new_n33865 = new_n33864 ^ new_n30679;
  assign new_n33866 = new_n33865 ^ new_n31172;
  assign new_n33867 = new_n33866 ^ new_n33863;
  assign new_n33868 = new_n31085 ^ new_n30993;
  assign new_n33869 = new_n33868 ^ new_n31055;
  assign new_n33870 = new_n29593 ^ new_n28769;
  assign new_n33871 = new_n33870 ^ new_n30968;
  assign new_n33872 = new_n33871 ^ new_n31115;
  assign new_n33873 = new_n33872 ^ new_n33869;
  assign new_n33874 = new_n31063 ^ new_n31002;
  assign new_n33875 = new_n33874 ^ new_n30968;
  assign new_n33876 = new_n31152 ^ new_n31068;
  assign new_n33877 = new_n29649 ^ new_n28734;
  assign new_n33878 = new_n33877 ^ new_n31202;
  assign new_n33879 = new_n33878 ^ new_n33876;
  assign new_n33880 = new_n33879 ^ new_n33875;
  assign new_n33881 = new_n31202 ^ new_n31104;
  assign new_n33882 = new_n31130 ^ new_n31047;
  assign new_n33883 = new_n33882 ^ new_n33881;
  assign new_n33884 = new_n29688 ^ new_n28728;
  assign new_n33885 = new_n33884 ^ new_n31115;
  assign new_n33886 = new_n33885 ^ new_n31139;
  assign new_n33887 = new_n33886 ^ new_n33883;
  assign new_n33888 = new_n33887 ^ new_n33880;
  assign new_n33889 = new_n33888 ^ new_n33873;
  assign new_n33890 = new_n33889 ^ new_n33867;
  assign new_n33891 = new_n29698 ^ new_n28762;
  assign new_n33892 = new_n33891 ^ new_n31139;
  assign new_n33893 = new_n31144 ^ new_n31106;
  assign new_n33894 = new_n33893 ^ new_n31202;
  assign new_n33895 = new_n33894 ^ new_n33892;
  assign new_n33896 = new_n29709 ^ new_n28744;
  assign new_n33897 = new_n31166 ^ new_n31158;
  assign new_n33898 = new_n33897 ^ new_n33896;
  assign new_n33899 = new_n33898 ^ new_n31202;
  assign new_n33900 = new_n31159 ^ new_n31072;
  assign new_n33901 = new_n33900 ^ new_n31063;
  assign new_n33902 = new_n33901 ^ new_n33899;
  assign new_n33903 = new_n31181 ^ new_n30363;
  assign new_n33904 = new_n33903 ^ new_n31172;
  assign new_n33905 = new_n29739 ^ new_n28758;
  assign new_n33906 = new_n33905 ^ new_n31161;
  assign new_n33907 = new_n33906 ^ new_n33904;
  assign new_n33908 = new_n33907 ^ new_n33867;
  assign new_n33909 = new_n33908 ^ new_n33895;
  assign new_n33910 = new_n33909 ^ new_n33902;
  assign new_n33911 = new_n33895 & new_n33910;
  assign new_n33912 = new_n33911 ^ new_n33902;
  assign new_n33913 = new_n31199 ^ new_n31095;
  assign new_n33914 = new_n33913 ^ new_n30526;
  assign new_n33915 = new_n29763 ^ new_n28740;
  assign new_n33916 = new_n33915 ^ new_n31201;
  assign new_n33917 = new_n33916 ^ new_n30679;
  assign new_n33918 = new_n33917 ^ new_n33914;
  assign new_n33919 = new_n33918 ^ new_n33902;
  assign new_n33920 = new_n33919 ^ new_n33888;
  assign new_n33921 = new_n33918 ^ new_n33887;
  assign new_n33922 = new_n33902 ^ new_n33873;
  assign new_n33923 = new_n33922 ^ new_n33921;
  assign new_n33924 = new_n33920 & new_n33923;
  assign new_n33925 = new_n33924 ^ new_n33867;
  assign new_n33926 = new_n33925 ^ new_n33912;
  assign new_n33927 = ~new_n33887 & ~new_n33909;
  assign new_n33928 = new_n33927 ^ new_n33887;
  assign new_n33929 = new_n33907 ^ new_n33889;
  assign new_n33930 = new_n33921 & new_n33929;
  assign new_n33931 = new_n33930 ^ new_n33928;
  assign new_n33932 = new_n33918 ^ new_n33873;
  assign new_n33933 = new_n33932 ^ new_n33931;
  assign new_n33934 = new_n33890 & new_n33919;
  assign new_n33935 = new_n33907 ^ new_n33902;
  assign new_n33936 = new_n33935 ^ new_n33932;
  assign new_n33937 = new_n33922 & new_n33936;
  assign new_n33938 = new_n33937 ^ new_n33934;
  assign new_n33939 = new_n33907 ^ new_n33880;
  assign new_n33940 = new_n33939 ^ new_n33938;
  assign new_n33941 = new_n33940 ^ new_n33933;
  assign new_n33942 = new_n33925 ^ new_n33920;
  assign new_n33943 = new_n33909 ^ new_n33887;
  assign new_n33944 = new_n33943 ^ new_n33932;
  assign new_n33945 = new_n33920 ^ new_n33895;
  assign new_n33946 = new_n33944 & new_n33945;
  assign new_n33947 = new_n33946 ^ new_n33934;
  assign new_n33948 = new_n33937 ^ new_n33873;
  assign new_n33949 = new_n33948 ^ new_n33947;
  assign new_n33950 = new_n33949 ^ new_n33942;
  assign new_n33951 = ~new_n33941 & new_n33950;
  assign new_n33952 = new_n33951 ^ new_n33926;
  assign new_n33953 = new_n33920 ^ new_n33908;
  assign new_n33954 = new_n33932 & new_n33953;
  assign new_n33955 = new_n33954 ^ new_n33934;
  assign new_n33956 = new_n33955 ^ new_n33929;
  assign new_n33957 = new_n33956 ^ new_n33952;
  assign new_n33958 = new_n33918 ^ new_n33909;
  assign new_n33959 = new_n33895 ^ new_n33890;
  assign new_n33960 = new_n33958 & new_n33959;
  assign new_n33961 = new_n33960 ^ new_n33927;
  assign new_n33962 = new_n33954 ^ new_n33937;
  assign new_n33963 = new_n33962 ^ new_n33961;
  assign new_n33964 = ~new_n33963 & new_n33957;
  assign new_n33965 = new_n33918 ^ new_n33907;
  assign new_n33966 = new_n33946 ^ new_n33911;
  assign new_n33967 = new_n33966 ^ new_n33962;
  assign new_n33968 = new_n33967 ^ new_n33965;
  assign new_n33969 = new_n33960 ^ new_n33930;
  assign new_n33970 = new_n33969 ^ new_n33918;
  assign new_n33971 = new_n33970 ^ new_n33956;
  assign new_n33972 = new_n33971 ^ new_n33951;
  assign new_n33973 = new_n33968 & new_n33972;
  assign new_n33974 = new_n33973 ^ new_n33964;
  assign new_n33975 = new_n33970 ^ new_n33926;
  assign new_n33976 = new_n33975 ^ new_n33974;
  assign new_n33977 = new_n33890 & new_n33976;
  assign new_n33978 = new_n33964 ^ new_n33951;
  assign new_n33979 = new_n33971 & new_n33978;
  assign new_n33980 = new_n33979 ^ new_n33941;
  assign new_n33981 = ~new_n33980 & new_n33923;
  assign new_n33982 = new_n33981 ^ new_n33977;
  assign new_n33983 = new_n33907 ^ new_n33887;
  assign new_n33984 = new_n33946 ^ new_n33928;
  assign new_n33985 = new_n33973 ^ new_n33926;
  assign new_n33986 = new_n33985 ^ new_n33956;
  assign new_n33987 = new_n33979 ^ new_n33972;
  assign new_n33988 = new_n33986 & new_n33987;
  assign new_n33989 = new_n33988 ^ new_n33979;
  assign new_n33990 = new_n33989 ^ new_n33984;
  assign new_n33991 = new_n33990 ^ new_n33983;
  assign new_n33992 = new_n33991 ^ new_n33902;
  assign new_n33993 = new_n33973 ^ new_n33930;
  assign new_n33994 = new_n33993 ^ new_n33925;
  assign new_n33995 = new_n33994 ^ new_n33992;
  assign new_n33996 = ~new_n33995 & new_n33936;
  assign new_n33997 = new_n33988 ^ new_n33968;
  assign new_n33998 = new_n33909 & new_n33997;
  assign new_n33999 = new_n33979 ^ new_n33964;
  assign new_n34000 = new_n33999 ^ new_n33963;
  assign new_n34001 = ~new_n34000 & new_n33944;
  assign new_n34002 = ~new_n33995 & new_n33922;
  assign new_n34003 = new_n33919 & new_n33976;
  assign new_n34004 = new_n34003 ^ new_n34002;
  assign new_n34005 = new_n34004 ^ new_n34001;
  assign new_n34006 = new_n34005 ^ new_n33998;
  assign new_n34007 = new_n33988 ^ new_n33973;
  assign new_n34008 = new_n34007 ^ new_n33950;
  assign new_n34009 = new_n33929 & new_n34008;
  assign new_n34010 = new_n34009 ^ new_n34006;
  assign new_n34011 = new_n34010 ^ new_n33996;
  assign new_n34012 = new_n34011 ^ new_n33982;
  assign new_n34013 = new_n30119 ^ new_n29763;
  assign new_n34014 = new_n34013 ^ new_n23827;
  assign new_n34015 = new_n34014 ^ new_n34012;
  assign new_n34016 = new_n30128 ^ new_n28590;
  assign new_n34017 = new_n34016 ^ new_n23859;
  assign new_n34018 = new_n33996 ^ new_n33977;
  assign new_n34019 = ~new_n33980 & new_n33920;
  assign new_n34020 = ~new_n34000 & new_n33945;
  assign new_n34021 = new_n34020 ^ new_n34019;
  assign new_n34022 = new_n34021 ^ new_n33981;
  assign new_n34023 = new_n34022 ^ new_n34005;
  assign new_n34024 = new_n34023 ^ new_n34018;
  assign new_n34025 = new_n34024 ^ new_n34017;
  assign new_n34026 = new_n30154 ^ new_n29739;
  assign new_n34027 = new_n34026 ^ new_n23868;
  assign new_n34028 = new_n34003 ^ new_n33977;
  assign new_n34029 = new_n33964 ^ new_n33918;
  assign new_n34030 = new_n33960 ^ new_n33911;
  assign new_n34031 = new_n34030 ^ new_n33991;
  assign new_n34032 = new_n34031 ^ new_n34029;
  assign new_n34033 = ~new_n34032 & new_n33932;
  assign new_n34034 = new_n33921 & new_n34008;
  assign new_n34035 = new_n33971 ^ new_n33964;
  assign new_n34036 = new_n33895 & new_n34035;
  assign new_n34037 = new_n34036 ^ new_n34019;
  assign new_n34038 = new_n34037 ^ new_n34034;
  assign new_n34039 = ~new_n34032 & new_n33953;
  assign new_n34040 = new_n33958 & new_n33986;
  assign new_n34041 = new_n34040 ^ new_n34039;
  assign new_n34042 = new_n34041 ^ new_n34038;
  assign new_n34043 = new_n34042 ^ new_n34033;
  assign new_n34044 = new_n34043 ^ new_n34028;
  assign new_n34045 = new_n34044 ^ new_n34027;
  assign new_n34046 = new_n34022 ^ new_n34010;
  assign new_n34047 = new_n30175 ^ new_n29709;
  assign new_n34048 = new_n34047 ^ new_n23832;
  assign new_n34049 = new_n34048 ^ new_n34046;
  assign new_n34050 = new_n33959 & new_n33986;
  assign new_n34051 = new_n34050 ^ new_n33981;
  assign new_n34052 = new_n34036 ^ new_n34020;
  assign new_n34053 = new_n34052 ^ new_n34006;
  assign new_n34054 = new_n34053 ^ new_n34051;
  assign new_n34055 = new_n30187 ^ new_n29649;
  assign new_n34056 = new_n34055 ^ new_n23818;
  assign new_n34057 = new_n34056 ^ new_n34054;
  assign new_n34058 = new_n33910 & new_n34035;
  assign new_n34059 = new_n34058 ^ new_n34011;
  assign new_n34060 = new_n34059 ^ new_n34042;
  assign new_n34061 = new_n30195 ^ new_n29593;
  assign new_n34062 = new_n34061 ^ new_n23851;
  assign new_n34063 = new_n34062 ^ new_n34060;
  assign new_n34064 = new_n30204 ^ new_n29688;
  assign new_n34065 = new_n34064 ^ new_n23811;
  assign new_n34066 = new_n34039 ^ new_n34034;
  assign new_n34067 = new_n33943 & new_n33997;
  assign new_n34068 = new_n34067 ^ new_n34050;
  assign new_n34069 = new_n34068 ^ new_n34004;
  assign new_n34070 = new_n33998 ^ new_n33996;
  assign new_n34071 = new_n34070 ^ new_n34069;
  assign new_n34072 = new_n34071 ^ new_n34066;
  assign new_n34073 = new_n34072 ^ new_n34065;
  assign new_n34074 = new_n30215 ^ new_n29698;
  assign new_n34075 = new_n34074 ^ new_n23842;
  assign new_n34076 = new_n34038 ^ new_n34009;
  assign new_n34077 = new_n34076 ^ new_n34069;
  assign new_n34078 = new_n34077 ^ new_n34075;
  assign new_n34079 = new_n30788 ^ new_n28180;
  assign new_n34080 = new_n34079 ^ new_n32453;
  assign new_n34081 = new_n32425 ^ new_n31930;
  assign new_n34082 = new_n34081 ^ new_n31781;
  assign new_n34083 = new_n34082 ^ new_n34080;
  assign new_n34084 = new_n31029 ^ new_n28102;
  assign new_n34085 = new_n34084 ^ new_n32319;
  assign new_n34086 = new_n34085 ^ new_n32366;
  assign new_n34087 = new_n34086 ^ new_n32254;
  assign new_n34088 = new_n31091 ^ new_n28224;
  assign new_n34089 = new_n34088 ^ new_n32413;
  assign new_n34090 = new_n32446 ^ new_n32348;
  assign new_n34091 = new_n34090 ^ new_n34089;
  assign new_n34092 = new_n32305 ^ new_n32217;
  assign new_n34093 = new_n34092 ^ new_n32336;
  assign new_n34094 = new_n34093 ^ new_n34091;
  assign new_n34095 = new_n32366 ^ new_n32271;
  assign new_n34096 = new_n34095 ^ new_n34090;
  assign new_n34097 = new_n31122 ^ new_n28160;
  assign new_n34098 = new_n34097 ^ new_n32359;
  assign new_n34099 = new_n34098 ^ new_n32398;
  assign new_n34100 = new_n34099 ^ new_n34096;
  assign new_n34101 = new_n34100 ^ new_n34094;
  assign new_n34102 = new_n34101 ^ new_n34087;
  assign new_n34103 = new_n34102 ^ new_n34083;
  assign new_n34104 = new_n31141 ^ new_n28202;
  assign new_n34105 = new_n34104 ^ new_n32390;
  assign new_n34106 = new_n32397 ^ new_n32372;
  assign new_n34107 = new_n34106 ^ new_n34090;
  assign new_n34108 = new_n34107 ^ new_n34105;
  assign new_n34109 = new_n32330 ^ new_n32323;
  assign new_n34110 = new_n34109 ^ new_n32403;
  assign new_n34111 = new_n31154 ^ new_n27968;
  assign new_n34112 = new_n34111 ^ new_n32436;
  assign new_n34113 = new_n34112 ^ new_n34090;
  assign new_n34114 = new_n34113 ^ new_n34110;
  assign new_n34115 = new_n31176 ^ new_n28024;
  assign new_n34116 = new_n34115 ^ new_n32171;
  assign new_n34117 = new_n32414 ^ new_n32401;
  assign new_n34118 = new_n34117 ^ new_n32426;
  assign new_n34119 = new_n34118 ^ new_n34116;
  assign new_n34120 = new_n34119 ^ new_n34083;
  assign new_n34121 = new_n34120 ^ new_n34108;
  assign new_n34122 = new_n34121 ^ new_n34114;
  assign new_n34123 = new_n34108 & new_n34122;
  assign new_n34124 = new_n34123 ^ new_n34114;
  assign new_n34125 = new_n31191 ^ new_n28118;
  assign new_n34126 = new_n34125 ^ new_n32346;
  assign new_n34127 = new_n32190 ^ new_n31780;
  assign new_n34128 = new_n34127 ^ new_n32449;
  assign new_n34129 = new_n34128 ^ new_n34126;
  assign new_n34130 = new_n34129 ^ new_n34114;
  assign new_n34131 = new_n34130 ^ new_n34101;
  assign new_n34132 = new_n34114 ^ new_n34100;
  assign new_n34133 = new_n34129 ^ new_n34087;
  assign new_n34134 = new_n34133 ^ new_n34132;
  assign new_n34135 = new_n34131 & new_n34134;
  assign new_n34136 = new_n34135 ^ new_n34083;
  assign new_n34137 = new_n34136 ^ new_n34124;
  assign new_n34138 = ~new_n34100 & ~new_n34121;
  assign new_n34139 = new_n34138 ^ new_n34100;
  assign new_n34140 = new_n34119 ^ new_n34102;
  assign new_n34141 = new_n34129 ^ new_n34100;
  assign new_n34142 = new_n34140 & new_n34141;
  assign new_n34143 = new_n34142 ^ new_n34139;
  assign new_n34144 = new_n34143 ^ new_n34133;
  assign new_n34145 = new_n34103 & new_n34130;
  assign new_n34146 = new_n34119 ^ new_n34114;
  assign new_n34147 = new_n34146 ^ new_n34133;
  assign new_n34148 = new_n34114 ^ new_n34087;
  assign new_n34149 = new_n34147 & new_n34148;
  assign new_n34150 = new_n34149 ^ new_n34145;
  assign new_n34151 = new_n34119 ^ new_n34094;
  assign new_n34152 = new_n34151 ^ new_n34150;
  assign new_n34153 = new_n34152 ^ new_n34144;
  assign new_n34154 = new_n34136 ^ new_n34131;
  assign new_n34155 = new_n34121 ^ new_n34100;
  assign new_n34156 = new_n34155 ^ new_n34133;
  assign new_n34157 = new_n34131 ^ new_n34108;
  assign new_n34158 = new_n34156 & new_n34157;
  assign new_n34159 = new_n34158 ^ new_n34145;
  assign new_n34160 = new_n34149 ^ new_n34087;
  assign new_n34161 = new_n34160 ^ new_n34159;
  assign new_n34162 = new_n34161 ^ new_n34154;
  assign new_n34163 = ~new_n34153 & new_n34162;
  assign new_n34164 = new_n34163 ^ new_n34137;
  assign new_n34165 = new_n34131 ^ new_n34120;
  assign new_n34166 = new_n34133 & new_n34165;
  assign new_n34167 = new_n34166 ^ new_n34145;
  assign new_n34168 = new_n34167 ^ new_n34140;
  assign new_n34169 = new_n34168 ^ new_n34164;
  assign new_n34170 = new_n34129 ^ new_n34121;
  assign new_n34171 = new_n34108 ^ new_n34103;
  assign new_n34172 = new_n34170 & new_n34171;
  assign new_n34173 = new_n34172 ^ new_n34138;
  assign new_n34174 = new_n34166 ^ new_n34149;
  assign new_n34175 = new_n34174 ^ new_n34173;
  assign new_n34176 = ~new_n34175 & new_n34169;
  assign new_n34177 = new_n34129 ^ new_n34119;
  assign new_n34178 = new_n34158 ^ new_n34123;
  assign new_n34179 = new_n34178 ^ new_n34174;
  assign new_n34180 = new_n34179 ^ new_n34177;
  assign new_n34181 = new_n34172 ^ new_n34142;
  assign new_n34182 = new_n34181 ^ new_n34129;
  assign new_n34183 = new_n34182 ^ new_n34168;
  assign new_n34184 = new_n34183 ^ new_n34163;
  assign new_n34185 = new_n34180 & new_n34184;
  assign new_n34186 = new_n34185 ^ new_n34176;
  assign new_n34187 = new_n34182 ^ new_n34137;
  assign new_n34188 = new_n34187 ^ new_n34186;
  assign new_n34189 = new_n34103 & new_n34188;
  assign new_n34190 = new_n34176 ^ new_n34163;
  assign new_n34191 = new_n34183 & new_n34190;
  assign new_n34192 = new_n34191 ^ new_n34153;
  assign new_n34193 = ~new_n34192 & new_n34134;
  assign new_n34194 = new_n34193 ^ new_n34189;
  assign new_n34195 = new_n34119 ^ new_n34100;
  assign new_n34196 = new_n34158 ^ new_n34139;
  assign new_n34197 = new_n34185 ^ new_n34137;
  assign new_n34198 = new_n34197 ^ new_n34168;
  assign new_n34199 = new_n34191 ^ new_n34184;
  assign new_n34200 = new_n34198 & new_n34199;
  assign new_n34201 = new_n34200 ^ new_n34191;
  assign new_n34202 = new_n34201 ^ new_n34196;
  assign new_n34203 = new_n34202 ^ new_n34195;
  assign new_n34204 = new_n34203 ^ new_n34114;
  assign new_n34205 = new_n34185 ^ new_n34142;
  assign new_n34206 = new_n34205 ^ new_n34136;
  assign new_n34207 = new_n34206 ^ new_n34204;
  assign new_n34208 = ~new_n34207 & new_n34147;
  assign new_n34209 = new_n34200 ^ new_n34180;
  assign new_n34210 = new_n34121 & new_n34209;
  assign new_n34211 = new_n34191 ^ new_n34176;
  assign new_n34212 = new_n34211 ^ new_n34175;
  assign new_n34213 = ~new_n34212 & new_n34156;
  assign new_n34214 = ~new_n34207 & new_n34148;
  assign new_n34215 = new_n34130 & new_n34188;
  assign new_n34216 = new_n34215 ^ new_n34214;
  assign new_n34217 = new_n34216 ^ new_n34213;
  assign new_n34218 = new_n34217 ^ new_n34210;
  assign new_n34219 = new_n34200 ^ new_n34185;
  assign new_n34220 = new_n34219 ^ new_n34162;
  assign new_n34221 = new_n34140 & new_n34220;
  assign new_n34222 = new_n34221 ^ new_n34218;
  assign new_n34223 = new_n34222 ^ new_n34208;
  assign new_n34224 = new_n34223 ^ new_n34194;
  assign new_n34225 = new_n31408 ^ new_n31191;
  assign new_n34226 = new_n34225 ^ new_n21305;
  assign new_n34227 = new_n34226 ^ new_n34224;
  assign new_n34228 = new_n31417 ^ new_n30788;
  assign new_n34229 = new_n34228 ^ new_n22058;
  assign new_n34230 = new_n34208 ^ new_n34189;
  assign new_n34231 = ~new_n34192 & new_n34131;
  assign new_n34232 = ~new_n34212 & new_n34157;
  assign new_n34233 = new_n34232 ^ new_n34231;
  assign new_n34234 = new_n34233 ^ new_n34193;
  assign new_n34235 = new_n34234 ^ new_n34217;
  assign new_n34236 = new_n34235 ^ new_n34230;
  assign new_n34237 = new_n34236 ^ new_n34229;
  assign new_n34238 = new_n31443 ^ new_n31176;
  assign new_n34239 = new_n34238 ^ new_n22081;
  assign new_n34240 = new_n34215 ^ new_n34189;
  assign new_n34241 = new_n34176 ^ new_n34129;
  assign new_n34242 = new_n34172 ^ new_n34123;
  assign new_n34243 = new_n34242 ^ new_n34203;
  assign new_n34244 = new_n34243 ^ new_n34241;
  assign new_n34245 = ~new_n34244 & new_n34133;
  assign new_n34246 = new_n34141 & new_n34220;
  assign new_n34247 = new_n34183 ^ new_n34176;
  assign new_n34248 = new_n34108 & new_n34247;
  assign new_n34249 = new_n34248 ^ new_n34231;
  assign new_n34250 = new_n34249 ^ new_n34246;
  assign new_n34251 = ~new_n34244 & new_n34165;
  assign new_n34252 = new_n34170 & new_n34198;
  assign new_n34253 = new_n34252 ^ new_n34251;
  assign new_n34254 = new_n34253 ^ new_n34250;
  assign new_n34255 = new_n34254 ^ new_n34245;
  assign new_n34256 = new_n34255 ^ new_n34240;
  assign new_n34257 = new_n34256 ^ new_n34239;
  assign new_n34258 = new_n34234 ^ new_n34222;
  assign new_n34259 = new_n31464 ^ new_n31154;
  assign new_n34260 = new_n34259 ^ new_n22092;
  assign new_n34261 = new_n34260 ^ new_n34258;
  assign new_n34262 = new_n34171 & new_n34198;
  assign new_n34263 = new_n34262 ^ new_n34193;
  assign new_n34264 = new_n34248 ^ new_n34232;
  assign new_n34265 = new_n34264 ^ new_n34218;
  assign new_n34266 = new_n34265 ^ new_n34263;
  assign new_n34267 = new_n31476 ^ new_n31091;
  assign new_n34268 = new_n34267 ^ new_n22125;
  assign new_n34269 = new_n34268 ^ new_n34266;
  assign new_n34270 = new_n34122 & new_n34247;
  assign new_n34271 = new_n34270 ^ new_n34223;
  assign new_n34272 = new_n34271 ^ new_n34254;
  assign new_n34273 = new_n31484 ^ new_n31029;
  assign new_n34274 = new_n34273 ^ new_n22018;
  assign new_n34275 = new_n34274 ^ new_n34272;
  assign new_n34276 = new_n31493 ^ new_n31122;
  assign new_n34277 = new_n34276 ^ new_n21957;
  assign new_n34278 = new_n34251 ^ new_n34246;
  assign new_n34279 = new_n34155 & new_n34209;
  assign new_n34280 = new_n34279 ^ new_n34262;
  assign new_n34281 = new_n34280 ^ new_n34216;
  assign new_n34282 = new_n34210 ^ new_n34208;
  assign new_n34283 = new_n34282 ^ new_n34281;
  assign new_n34284 = new_n34283 ^ new_n34278;
  assign new_n34285 = new_n34284 ^ new_n34277;
  assign new_n34286 = new_n31504 ^ new_n31141;
  assign new_n34287 = new_n34286 ^ new_n22149;
  assign new_n34288 = new_n34250 ^ new_n34221;
  assign new_n34289 = new_n34288 ^ new_n34281;
  assign new_n34290 = new_n34289 ^ new_n34287;
  assign new_n34291 = new_n33652 ^ new_n33547;
  assign new_n34292 = new_n33531 ^ new_n33345;
  assign new_n34293 = new_n34292 ^ new_n33191;
  assign new_n34294 = new_n34293 ^ new_n34291;
  assign new_n34295 = new_n33467 ^ new_n33414;
  assign new_n34296 = new_n34295 ^ new_n33435;
  assign new_n34297 = new_n33653 ^ new_n33389;
  assign new_n34298 = new_n34297 ^ new_n33491;
  assign new_n34299 = new_n34298 ^ new_n34296;
  assign new_n34300 = new_n33442 ^ new_n33389;
  assign new_n34301 = new_n34300 ^ new_n33426;
  assign new_n34302 = new_n33519 ^ new_n33447;
  assign new_n34303 = new_n33549 ^ new_n33462;
  assign new_n34304 = new_n34303 ^ new_n33654;
  assign new_n34305 = new_n34304 ^ new_n34302;
  assign new_n34306 = new_n34305 ^ new_n34301;
  assign new_n34307 = new_n34303 ^ new_n33495;
  assign new_n34308 = new_n33484 ^ new_n33364;
  assign new_n34309 = new_n34308 ^ new_n34307;
  assign new_n34310 = new_n33655 ^ new_n33491;
  assign new_n34311 = new_n34310 ^ new_n33506;
  assign new_n34312 = new_n34311 ^ new_n34309;
  assign new_n34313 = new_n34312 ^ new_n34306;
  assign new_n34314 = new_n34313 ^ new_n34299;
  assign new_n34315 = new_n34314 ^ new_n34294;
  assign new_n34316 = new_n33659 ^ new_n33506;
  assign new_n34317 = new_n33504 ^ new_n33476;
  assign new_n34318 = new_n34317 ^ new_n34303;
  assign new_n34319 = new_n34318 ^ new_n34316;
  assign new_n34320 = new_n34303 ^ new_n33660;
  assign new_n34321 = new_n34320 ^ new_n33513;
  assign new_n34322 = new_n33471 ^ new_n33442;
  assign new_n34323 = new_n34322 ^ new_n33536;
  assign new_n34324 = new_n34323 ^ new_n34321;
  assign new_n34325 = new_n33661 ^ new_n32901;
  assign new_n34326 = new_n33520 ^ new_n33511;
  assign new_n34327 = new_n34326 ^ new_n33532;
  assign new_n34328 = new_n34327 ^ new_n34325;
  assign new_n34329 = new_n34328 ^ new_n34294;
  assign new_n34330 = new_n34329 ^ new_n34319;
  assign new_n34331 = new_n34330 ^ new_n34324;
  assign new_n34332 = new_n34319 & new_n34331;
  assign new_n34333 = new_n34332 ^ new_n34324;
  assign new_n34334 = new_n33667 ^ new_n33460;
  assign new_n34335 = new_n33325 ^ new_n33190;
  assign new_n34336 = new_n34335 ^ new_n33552;
  assign new_n34337 = new_n34336 ^ new_n34334;
  assign new_n34338 = new_n34337 ^ new_n34324;
  assign new_n34339 = new_n34338 ^ new_n34313;
  assign new_n34340 = new_n34337 ^ new_n34312;
  assign new_n34341 = new_n34324 ^ new_n34299;
  assign new_n34342 = new_n34341 ^ new_n34340;
  assign new_n34343 = new_n34339 & new_n34342;
  assign new_n34344 = new_n34343 ^ new_n34294;
  assign new_n34345 = new_n34344 ^ new_n34333;
  assign new_n34346 = ~new_n34312 & ~new_n34330;
  assign new_n34347 = new_n34346 ^ new_n34312;
  assign new_n34348 = new_n34328 ^ new_n34314;
  assign new_n34349 = new_n34340 & new_n34348;
  assign new_n34350 = new_n34349 ^ new_n34347;
  assign new_n34351 = new_n34337 ^ new_n34299;
  assign new_n34352 = new_n34351 ^ new_n34350;
  assign new_n34353 = new_n34315 & new_n34338;
  assign new_n34354 = new_n34328 ^ new_n34324;
  assign new_n34355 = new_n34354 ^ new_n34351;
  assign new_n34356 = new_n34341 & new_n34355;
  assign new_n34357 = new_n34356 ^ new_n34353;
  assign new_n34358 = new_n34328 ^ new_n34306;
  assign new_n34359 = new_n34358 ^ new_n34357;
  assign new_n34360 = new_n34359 ^ new_n34352;
  assign new_n34361 = new_n34344 ^ new_n34339;
  assign new_n34362 = new_n34330 ^ new_n34312;
  assign new_n34363 = new_n34362 ^ new_n34351;
  assign new_n34364 = new_n34339 ^ new_n34319;
  assign new_n34365 = new_n34363 & new_n34364;
  assign new_n34366 = new_n34365 ^ new_n34353;
  assign new_n34367 = new_n34356 ^ new_n34299;
  assign new_n34368 = new_n34367 ^ new_n34366;
  assign new_n34369 = new_n34368 ^ new_n34361;
  assign new_n34370 = ~new_n34360 & new_n34369;
  assign new_n34371 = new_n34370 ^ new_n34345;
  assign new_n34372 = new_n34339 ^ new_n34329;
  assign new_n34373 = new_n34351 & new_n34372;
  assign new_n34374 = new_n34373 ^ new_n34353;
  assign new_n34375 = new_n34374 ^ new_n34348;
  assign new_n34376 = new_n34375 ^ new_n34371;
  assign new_n34377 = new_n34337 ^ new_n34330;
  assign new_n34378 = new_n34319 ^ new_n34315;
  assign new_n34379 = new_n34377 & new_n34378;
  assign new_n34380 = new_n34379 ^ new_n34346;
  assign new_n34381 = new_n34373 ^ new_n34356;
  assign new_n34382 = new_n34381 ^ new_n34380;
  assign new_n34383 = ~new_n34382 & new_n34376;
  assign new_n34384 = new_n34337 ^ new_n34328;
  assign new_n34385 = new_n34365 ^ new_n34332;
  assign new_n34386 = new_n34385 ^ new_n34381;
  assign new_n34387 = new_n34386 ^ new_n34384;
  assign new_n34388 = new_n34379 ^ new_n34349;
  assign new_n34389 = new_n34388 ^ new_n34337;
  assign new_n34390 = new_n34389 ^ new_n34375;
  assign new_n34391 = new_n34390 ^ new_n34370;
  assign new_n34392 = new_n34387 & new_n34391;
  assign new_n34393 = new_n34392 ^ new_n34383;
  assign new_n34394 = new_n34389 ^ new_n34345;
  assign new_n34395 = new_n34394 ^ new_n34393;
  assign new_n34396 = new_n34315 & new_n34395;
  assign new_n34397 = new_n34383 ^ new_n34370;
  assign new_n34398 = new_n34390 & new_n34397;
  assign new_n34399 = new_n34398 ^ new_n34360;
  assign new_n34400 = ~new_n34399 & new_n34342;
  assign new_n34401 = new_n34400 ^ new_n34396;
  assign new_n34402 = new_n34328 ^ new_n34312;
  assign new_n34403 = new_n34365 ^ new_n34347;
  assign new_n34404 = new_n34392 ^ new_n34345;
  assign new_n34405 = new_n34404 ^ new_n34375;
  assign new_n34406 = new_n34398 ^ new_n34391;
  assign new_n34407 = new_n34405 & new_n34406;
  assign new_n34408 = new_n34407 ^ new_n34398;
  assign new_n34409 = new_n34408 ^ new_n34403;
  assign new_n34410 = new_n34409 ^ new_n34402;
  assign new_n34411 = new_n34410 ^ new_n34324;
  assign new_n34412 = new_n34392 ^ new_n34349;
  assign new_n34413 = new_n34412 ^ new_n34344;
  assign new_n34414 = new_n34413 ^ new_n34411;
  assign new_n34415 = ~new_n34414 & new_n34355;
  assign new_n34416 = new_n34407 ^ new_n34387;
  assign new_n34417 = new_n34330 & new_n34416;
  assign new_n34418 = new_n34398 ^ new_n34383;
  assign new_n34419 = new_n34418 ^ new_n34382;
  assign new_n34420 = ~new_n34419 & new_n34363;
  assign new_n34421 = ~new_n34414 & new_n34341;
  assign new_n34422 = new_n34338 & new_n34395;
  assign new_n34423 = new_n34422 ^ new_n34421;
  assign new_n34424 = new_n34423 ^ new_n34420;
  assign new_n34425 = new_n34424 ^ new_n34417;
  assign new_n34426 = new_n34407 ^ new_n34392;
  assign new_n34427 = new_n34426 ^ new_n34369;
  assign new_n34428 = new_n34348 & new_n34427;
  assign new_n34429 = new_n34428 ^ new_n34425;
  assign new_n34430 = new_n34429 ^ new_n34415;
  assign new_n34431 = new_n34430 ^ new_n34401;
  assign new_n34432 = new_n32665 ^ new_n32455;
  assign new_n34433 = new_n34432 ^ new_n25060;
  assign new_n34434 = new_n34433 ^ new_n34431;
  assign new_n34435 = new_n32674 ^ new_n32033;
  assign new_n34436 = new_n34435 ^ new_n25014;
  assign new_n34437 = new_n34415 ^ new_n34396;
  assign new_n34438 = ~new_n34399 & new_n34339;
  assign new_n34439 = ~new_n34419 & new_n34364;
  assign new_n34440 = new_n34439 ^ new_n34438;
  assign new_n34441 = new_n34440 ^ new_n34400;
  assign new_n34442 = new_n34441 ^ new_n34424;
  assign new_n34443 = new_n34442 ^ new_n34437;
  assign new_n34444 = new_n34443 ^ new_n34436;
  assign new_n34445 = new_n32700 ^ new_n32431;
  assign new_n34446 = new_n34445 ^ new_n25050;
  assign new_n34447 = new_n34422 ^ new_n34396;
  assign new_n34448 = new_n34383 ^ new_n34337;
  assign new_n34449 = new_n34379 ^ new_n34332;
  assign new_n34450 = new_n34449 ^ new_n34410;
  assign new_n34451 = new_n34450 ^ new_n34448;
  assign new_n34452 = ~new_n34451 & new_n34351;
  assign new_n34453 = new_n34340 & new_n34427;
  assign new_n34454 = new_n34390 ^ new_n34383;
  assign new_n34455 = new_n34319 & new_n34454;
  assign new_n34456 = new_n34455 ^ new_n34438;
  assign new_n34457 = new_n34456 ^ new_n34453;
  assign new_n34458 = ~new_n34451 & new_n34372;
  assign new_n34459 = new_n34377 & new_n34405;
  assign new_n34460 = new_n34459 ^ new_n34458;
  assign new_n34461 = new_n34460 ^ new_n34457;
  assign new_n34462 = new_n34461 ^ new_n34452;
  assign new_n34463 = new_n34462 ^ new_n34447;
  assign new_n34464 = new_n34463 ^ new_n34446;
  assign new_n34465 = new_n34441 ^ new_n34429;
  assign new_n34466 = new_n32721 ^ new_n32404;
  assign new_n34467 = new_n34466 ^ new_n25045;
  assign new_n34468 = new_n34467 ^ new_n34465;
  assign new_n34469 = new_n34378 & new_n34405;
  assign new_n34470 = new_n34469 ^ new_n34400;
  assign new_n34471 = new_n34455 ^ new_n34439;
  assign new_n34472 = new_n34471 ^ new_n34425;
  assign new_n34473 = new_n34472 ^ new_n34470;
  assign new_n34474 = new_n32733 ^ new_n32341;
  assign new_n34475 = new_n34474 ^ new_n25019;
  assign new_n34476 = new_n34475 ^ new_n34473;
  assign new_n34477 = new_n34331 & new_n34454;
  assign new_n34478 = new_n34477 ^ new_n34430;
  assign new_n34479 = new_n34478 ^ new_n34461;
  assign new_n34480 = new_n32741 ^ new_n32296;
  assign new_n34481 = new_n34480 ^ new_n25032;
  assign new_n34482 = new_n34481 ^ new_n34479;
  assign new_n34483 = new_n32750 ^ new_n32380;
  assign new_n34484 = new_n34483 ^ new_n25026;
  assign new_n34485 = new_n34458 ^ new_n34453;
  assign new_n34486 = new_n34362 & new_n34416;
  assign new_n34487 = new_n34486 ^ new_n34469;
  assign new_n34488 = new_n34487 ^ new_n34423;
  assign new_n34489 = new_n34417 ^ new_n34415;
  assign new_n34490 = new_n34489 ^ new_n34488;
  assign new_n34491 = new_n34490 ^ new_n34485;
  assign new_n34492 = new_n34491 ^ new_n34484;
  assign new_n34493 = new_n32761 ^ new_n32392;
  assign new_n34494 = new_n34493 ^ new_n25039;
  assign new_n34495 = new_n34457 ^ new_n34428;
  assign new_n34496 = new_n34495 ^ new_n34488;
  assign new_n34497 = new_n34496 ^ new_n34494;
  assign new_n34498 = new_n29755 ^ new_n28326;
  assign new_n34499 = new_n34498 ^ new_n29729;
  assign new_n34500 = new_n29963 ^ new_n28484;
  assign new_n34501 = new_n34500 ^ new_n21607;
  assign new_n34502 = new_n34501 ^ new_n29497;
  assign new_n34503 = new_n34502 ^ new_n27255;
  assign new_n34504 = new_n34503 ^ new_n34499;
  assign new_n34505 = new_n29627 ^ new_n29566;
  assign new_n34506 = new_n34505 ^ new_n29670;
  assign new_n34507 = new_n29989 ^ new_n28465;
  assign new_n34508 = new_n34507 ^ new_n21585;
  assign new_n34509 = new_n34508 ^ new_n29541;
  assign new_n34510 = new_n34509 ^ new_n29614;
  assign new_n34511 = new_n34510 ^ new_n34506;
  assign new_n34512 = new_n29638 ^ new_n29541;
  assign new_n34513 = new_n34512 ^ new_n29605;
  assign new_n34514 = new_n29995 ^ new_n28499;
  assign new_n34515 = new_n34514 ^ new_n21590;
  assign new_n34516 = new_n29721 ^ new_n29643;
  assign new_n34517 = new_n34516 ^ new_n34515;
  assign new_n34518 = new_n29757 ^ new_n29653;
  assign new_n34519 = new_n34518 ^ new_n34517;
  assign new_n34520 = new_n34519 ^ new_n34513;
  assign new_n34521 = new_n29677 ^ new_n29516;
  assign new_n34522 = new_n34521 ^ new_n29703;
  assign new_n34523 = new_n34522 ^ new_n34518;
  assign new_n34524 = new_n30003 ^ new_n28479;
  assign new_n34525 = new_n34524 ^ new_n21599;
  assign new_n34526 = new_n34525 ^ new_n29681;
  assign new_n34527 = new_n34526 ^ new_n29670;
  assign new_n34528 = new_n34527 ^ new_n34523;
  assign new_n34529 = new_n34528 ^ new_n34520;
  assign new_n34530 = new_n34529 ^ new_n34511;
  assign new_n34531 = new_n34530 ^ new_n34504;
  assign new_n34532 = new_n30009 ^ new_n28488;
  assign new_n34533 = new_n34532 ^ new_n21626;
  assign new_n34534 = new_n34533 ^ new_n29703;
  assign new_n34535 = new_n29705 ^ new_n29662;
  assign new_n34536 = new_n34535 ^ new_n34518;
  assign new_n34537 = new_n34536 ^ new_n34534;
  assign new_n34538 = new_n30011 ^ new_n28439;
  assign new_n34539 = new_n34538 ^ new_n21641;
  assign new_n34540 = new_n29744 ^ new_n29713;
  assign new_n34541 = new_n34540 ^ new_n34539;
  assign new_n34542 = new_n34541 ^ new_n34518;
  assign new_n34543 = new_n29712 ^ new_n29638;
  assign new_n34544 = new_n34543 ^ new_n29631;
  assign new_n34545 = new_n34544 ^ new_n34542;
  assign new_n34546 = new_n29733 ^ new_n26210;
  assign new_n34547 = new_n34546 ^ new_n29729;
  assign new_n34548 = new_n30016 ^ new_n28458;
  assign new_n34549 = new_n34548 ^ new_n21620;
  assign new_n34550 = new_n29722 ^ new_n29712;
  assign new_n34551 = new_n34550 ^ new_n34549;
  assign new_n34552 = new_n34551 ^ new_n34547;
  assign new_n34553 = new_n34552 ^ new_n34504;
  assign new_n34554 = new_n34553 ^ new_n34537;
  assign new_n34555 = new_n34554 ^ new_n34545;
  assign new_n34556 = new_n34537 & new_n34555;
  assign new_n34557 = new_n34556 ^ new_n34545;
  assign new_n34558 = new_n29759 ^ new_n29656;
  assign new_n34559 = new_n34558 ^ new_n27255;
  assign new_n34560 = new_n30024 ^ new_n28468;
  assign new_n34561 = new_n34560 ^ new_n21614;
  assign new_n34562 = new_n34561 ^ new_n29757;
  assign new_n34563 = new_n34562 ^ new_n29477;
  assign new_n34564 = new_n34563 ^ new_n34559;
  assign new_n34565 = new_n34564 ^ new_n34545;
  assign new_n34566 = new_n34565 ^ new_n34529;
  assign new_n34567 = new_n34545 ^ new_n34528;
  assign new_n34568 = new_n34564 ^ new_n34511;
  assign new_n34569 = new_n34568 ^ new_n34567;
  assign new_n34570 = new_n34566 & new_n34569;
  assign new_n34571 = new_n34570 ^ new_n34504;
  assign new_n34572 = new_n34571 ^ new_n34557;
  assign new_n34573 = ~new_n34554 & new_n34528;
  assign new_n34574 = new_n34573 ^ new_n34528;
  assign new_n34575 = new_n34552 ^ new_n34530;
  assign new_n34576 = new_n34564 ^ new_n34528;
  assign new_n34577 = ~new_n34575 & new_n34576;
  assign new_n34578 = new_n34577 ^ new_n34574;
  assign new_n34579 = new_n34578 ^ new_n34568;
  assign new_n34580 = ~new_n34531 & ~new_n34565;
  assign new_n34581 = new_n34552 ^ new_n34545;
  assign new_n34582 = new_n34581 ^ new_n34568;
  assign new_n34583 = new_n34545 ^ new_n34511;
  assign new_n34584 = ~new_n34582 & new_n34583;
  assign new_n34585 = new_n34584 ^ new_n34580;
  assign new_n34586 = new_n34552 ^ new_n34520;
  assign new_n34587 = new_n34586 ^ new_n34585;
  assign new_n34588 = new_n34587 ^ new_n34579;
  assign new_n34589 = new_n34571 ^ new_n34566;
  assign new_n34590 = new_n34554 ^ new_n34528;
  assign new_n34591 = new_n34590 ^ new_n34568;
  assign new_n34592 = new_n34566 ^ new_n34537;
  assign new_n34593 = new_n34591 & new_n34592;
  assign new_n34594 = new_n34593 ^ new_n34580;
  assign new_n34595 = new_n34584 ^ new_n34511;
  assign new_n34596 = new_n34595 ^ new_n34594;
  assign new_n34597 = new_n34596 ^ new_n34589;
  assign new_n34598 = ~new_n34588 & new_n34597;
  assign new_n34599 = new_n34598 ^ new_n34572;
  assign new_n34600 = new_n34566 ^ new_n34553;
  assign new_n34601 = ~new_n34568 & new_n34600;
  assign new_n34602 = new_n34601 ^ new_n34580;
  assign new_n34603 = new_n34602 ^ new_n34575;
  assign new_n34604 = new_n34603 ^ new_n34599;
  assign new_n34605 = new_n34564 ^ new_n34554;
  assign new_n34606 = new_n34537 ^ new_n34531;
  assign new_n34607 = ~new_n34605 & ~new_n34606;
  assign new_n34608 = new_n34607 ^ new_n34573;
  assign new_n34609 = new_n34601 ^ new_n34584;
  assign new_n34610 = new_n34609 ^ new_n34608;
  assign new_n34611 = ~new_n34604 & ~new_n34610;
  assign new_n34612 = new_n34564 ^ new_n34552;
  assign new_n34613 = new_n34593 ^ new_n34556;
  assign new_n34614 = new_n34613 ^ new_n34609;
  assign new_n34615 = new_n34614 ^ new_n34612;
  assign new_n34616 = new_n34607 ^ new_n34577;
  assign new_n34617 = new_n34616 ^ new_n34564;
  assign new_n34618 = new_n34617 ^ new_n34603;
  assign new_n34619 = new_n34618 ^ new_n34598;
  assign new_n34620 = ~new_n34615 & new_n34619;
  assign new_n34621 = new_n34620 ^ new_n34611;
  assign new_n34622 = new_n34617 ^ new_n34572;
  assign new_n34623 = new_n34622 ^ new_n34621;
  assign new_n34624 = ~new_n34531 & ~new_n34623;
  assign new_n34625 = new_n34611 ^ new_n34598;
  assign new_n34626 = new_n34618 & new_n34625;
  assign new_n34627 = new_n34626 ^ new_n34588;
  assign new_n34628 = ~new_n34627 & new_n34569;
  assign new_n34629 = new_n34628 ^ new_n34624;
  assign new_n34630 = new_n34552 ^ new_n34528;
  assign new_n34631 = new_n34593 ^ new_n34574;
  assign new_n34632 = new_n34620 ^ new_n34572;
  assign new_n34633 = new_n34632 ^ new_n34603;
  assign new_n34634 = new_n34626 ^ new_n34619;
  assign new_n34635 = ~new_n34633 & new_n34634;
  assign new_n34636 = new_n34635 ^ new_n34626;
  assign new_n34637 = new_n34636 ^ new_n34631;
  assign new_n34638 = new_n34637 ^ new_n34630;
  assign new_n34639 = new_n34638 ^ new_n34545;
  assign new_n34640 = new_n34620 ^ new_n34577;
  assign new_n34641 = new_n34640 ^ new_n34571;
  assign new_n34642 = new_n34641 ^ new_n34639;
  assign new_n34643 = ~new_n34582 & ~new_n34642;
  assign new_n34644 = new_n34635 ^ new_n34615;
  assign new_n34645 = ~new_n34644 & new_n34554;
  assign new_n34646 = new_n34626 ^ new_n34611;
  assign new_n34647 = new_n34646 ^ new_n34610;
  assign new_n34648 = ~new_n34647 & new_n34591;
  assign new_n34649 = ~new_n34642 & new_n34583;
  assign new_n34650 = ~new_n34565 & ~new_n34623;
  assign new_n34651 = new_n34650 ^ new_n34649;
  assign new_n34652 = new_n34651 ^ new_n34648;
  assign new_n34653 = new_n34652 ^ new_n34645;
  assign new_n34654 = new_n34635 ^ new_n34620;
  assign new_n34655 = new_n34654 ^ new_n34597;
  assign new_n34656 = ~new_n34575 & new_n34655;
  assign new_n34657 = new_n34656 ^ new_n34653;
  assign new_n34658 = new_n34657 ^ new_n34643;
  assign new_n34659 = new_n34658 ^ new_n34629;
  assign new_n34660 = new_n33761 ^ new_n30024;
  assign new_n34661 = new_n34660 ^ new_n22740;
  assign new_n34662 = new_n34661 ^ new_n34659;
  assign new_n34663 = new_n33770 ^ new_n29963;
  assign new_n34664 = new_n34663 ^ new_n22710;
  assign new_n34665 = new_n34643 ^ new_n34624;
  assign new_n34666 = ~new_n34627 & new_n34566;
  assign new_n34667 = ~new_n34647 & new_n34592;
  assign new_n34668 = new_n34667 ^ new_n34666;
  assign new_n34669 = new_n34668 ^ new_n34628;
  assign new_n34670 = new_n34669 ^ new_n34652;
  assign new_n34671 = new_n34670 ^ new_n34665;
  assign new_n34672 = new_n34671 ^ new_n34664;
  assign new_n34673 = new_n33796 ^ new_n30016;
  assign new_n34674 = new_n34673 ^ new_n22728;
  assign new_n34675 = new_n34650 ^ new_n34624;
  assign new_n34676 = new_n34611 ^ new_n34564;
  assign new_n34677 = new_n34607 ^ new_n34556;
  assign new_n34678 = new_n34677 ^ new_n34638;
  assign new_n34679 = new_n34678 ^ new_n34676;
  assign new_n34680 = ~new_n34568 & new_n34679;
  assign new_n34681 = new_n34576 & new_n34655;
  assign new_n34682 = new_n34618 ^ new_n34611;
  assign new_n34683 = new_n34537 & new_n34682;
  assign new_n34684 = new_n34683 ^ new_n34666;
  assign new_n34685 = new_n34684 ^ new_n34681;
  assign new_n34686 = new_n34600 & new_n34679;
  assign new_n34687 = ~new_n34605 & ~new_n34633;
  assign new_n34688 = new_n34687 ^ new_n34686;
  assign new_n34689 = new_n34688 ^ new_n34685;
  assign new_n34690 = new_n34689 ^ new_n34680;
  assign new_n34691 = new_n34690 ^ new_n34675;
  assign new_n34692 = new_n34691 ^ new_n34674;
  assign new_n34693 = new_n34669 ^ new_n34657;
  assign new_n34694 = new_n33817 ^ new_n30011;
  assign new_n34695 = new_n34694 ^ new_n22721;
  assign new_n34696 = new_n34695 ^ new_n34693;
  assign new_n34697 = ~new_n34606 & ~new_n34633;
  assign new_n34698 = new_n34697 ^ new_n34628;
  assign new_n34699 = new_n34683 ^ new_n34667;
  assign new_n34700 = new_n34699 ^ new_n34653;
  assign new_n34701 = new_n34700 ^ new_n34698;
  assign new_n34702 = new_n33829 ^ new_n29995;
  assign new_n34703 = new_n34702 ^ new_n22694;
  assign new_n34704 = new_n34703 ^ new_n34701;
  assign new_n34705 = new_n34555 & new_n34682;
  assign new_n34706 = new_n34705 ^ new_n34658;
  assign new_n34707 = new_n34706 ^ new_n34689;
  assign new_n34708 = new_n33837 ^ new_n29989;
  assign new_n34709 = new_n34708 ^ new_n22687;
  assign new_n34710 = new_n34709 ^ new_n34707;
  assign new_n34711 = new_n33846 ^ new_n30003;
  assign new_n34712 = new_n34711 ^ new_n22702;
  assign new_n34713 = new_n34686 ^ new_n34681;
  assign new_n34714 = ~new_n34590 & ~new_n34644;
  assign new_n34715 = new_n34714 ^ new_n34697;
  assign new_n34716 = new_n34715 ^ new_n34651;
  assign new_n34717 = new_n34645 ^ new_n34643;
  assign new_n34718 = new_n34717 ^ new_n34716;
  assign new_n34719 = new_n34718 ^ new_n34713;
  assign new_n34720 = new_n34719 ^ new_n34712;
  assign new_n34721 = new_n33857 ^ new_n30009;
  assign new_n34722 = new_n34721 ^ new_n22716;
  assign new_n34723 = new_n34685 ^ new_n34656;
  assign new_n34724 = new_n34723 ^ new_n34716;
  assign new_n34725 = new_n34724 ^ new_n34722;
  assign new_n34726 = new_n32426 ^ new_n31648;
  assign new_n34727 = new_n30365 ^ new_n28590;
  assign new_n34728 = new_n34727 ^ new_n32453;
  assign new_n34729 = new_n34728 ^ new_n32190;
  assign new_n34730 = new_n34729 ^ new_n34726;
  assign new_n34731 = new_n32305 ^ new_n32242;
  assign new_n34732 = new_n34731 ^ new_n32319;
  assign new_n34733 = new_n30371 ^ new_n29593;
  assign new_n34734 = new_n34733 ^ new_n32367;
  assign new_n34735 = new_n34734 ^ new_n34732;
  assign new_n34736 = new_n32335 ^ new_n32323;
  assign new_n34737 = new_n34736 ^ new_n32413;
  assign new_n34738 = new_n30384 ^ new_n29649;
  assign new_n34739 = new_n34738 ^ new_n32449;
  assign new_n34740 = new_n34739 ^ new_n32243;
  assign new_n34741 = new_n34740 ^ new_n34737;
  assign new_n34742 = new_n32359 ^ new_n32271;
  assign new_n34743 = new_n34742 ^ new_n32390;
  assign new_n34744 = new_n34743 ^ new_n32449;
  assign new_n34745 = new_n30378 ^ new_n29688;
  assign new_n34746 = new_n34745 ^ new_n32397;
  assign new_n34747 = new_n34746 ^ new_n32253;
  assign new_n34748 = new_n34747 ^ new_n34744;
  assign new_n34749 = new_n34748 ^ new_n34741;
  assign new_n34750 = new_n34749 ^ new_n34735;
  assign new_n34751 = new_n34750 ^ new_n34730;
  assign new_n34752 = new_n30391 ^ new_n29698;
  assign new_n34753 = new_n34752 ^ new_n32390;
  assign new_n34754 = new_n32449 ^ new_n32373;
  assign new_n34755 = new_n34754 ^ new_n34753;
  assign new_n34756 = new_n30396 ^ new_n29709;
  assign new_n34757 = new_n34756 ^ new_n32449;
  assign new_n34758 = new_n34757 ^ new_n32336;
  assign new_n34759 = new_n32436 ^ new_n32402;
  assign new_n34760 = new_n34759 ^ new_n32414;
  assign new_n34761 = new_n34760 ^ new_n34758;
  assign new_n34762 = new_n32421 ^ new_n32403;
  assign new_n34763 = new_n30403 ^ new_n29739;
  assign new_n34764 = new_n34763 ^ new_n32171;
  assign new_n34765 = new_n34764 ^ new_n31930;
  assign new_n34766 = new_n34765 ^ new_n34762;
  assign new_n34767 = new_n34766 ^ new_n34730;
  assign new_n34768 = new_n34767 ^ new_n34755;
  assign new_n34769 = new_n34768 ^ new_n34761;
  assign new_n34770 = new_n34755 & new_n34769;
  assign new_n34771 = new_n34770 ^ new_n34761;
  assign new_n34772 = new_n30412 ^ new_n29763;
  assign new_n34773 = new_n34772 ^ new_n31781;
  assign new_n34774 = new_n32448 ^ new_n32349;
  assign new_n34775 = new_n34774 ^ new_n34773;
  assign new_n34776 = new_n34775 ^ new_n34761;
  assign new_n34777 = new_n34776 ^ new_n34749;
  assign new_n34778 = new_n34775 ^ new_n34748;
  assign new_n34779 = new_n34761 ^ new_n34735;
  assign new_n34780 = new_n34779 ^ new_n34778;
  assign new_n34781 = new_n34777 & new_n34780;
  assign new_n34782 = new_n34781 ^ new_n34730;
  assign new_n34783 = new_n34782 ^ new_n34771;
  assign new_n34784 = ~new_n34748 & ~new_n34768;
  assign new_n34785 = new_n34784 ^ new_n34748;
  assign new_n34786 = new_n34766 ^ new_n34750;
  assign new_n34787 = new_n34778 & new_n34786;
  assign new_n34788 = new_n34787 ^ new_n34785;
  assign new_n34789 = new_n34775 ^ new_n34735;
  assign new_n34790 = new_n34789 ^ new_n34788;
  assign new_n34791 = new_n34751 & new_n34776;
  assign new_n34792 = new_n34766 ^ new_n34761;
  assign new_n34793 = new_n34792 ^ new_n34789;
  assign new_n34794 = new_n34779 & new_n34793;
  assign new_n34795 = new_n34794 ^ new_n34791;
  assign new_n34796 = new_n34766 ^ new_n34741;
  assign new_n34797 = new_n34796 ^ new_n34795;
  assign new_n34798 = new_n34797 ^ new_n34790;
  assign new_n34799 = new_n34782 ^ new_n34777;
  assign new_n34800 = new_n34768 ^ new_n34748;
  assign new_n34801 = new_n34800 ^ new_n34789;
  assign new_n34802 = new_n34777 ^ new_n34755;
  assign new_n34803 = new_n34801 & new_n34802;
  assign new_n34804 = new_n34803 ^ new_n34791;
  assign new_n34805 = new_n34794 ^ new_n34735;
  assign new_n34806 = new_n34805 ^ new_n34804;
  assign new_n34807 = new_n34806 ^ new_n34799;
  assign new_n34808 = ~new_n34798 & new_n34807;
  assign new_n34809 = new_n34808 ^ new_n34783;
  assign new_n34810 = new_n34777 ^ new_n34767;
  assign new_n34811 = new_n34789 & new_n34810;
  assign new_n34812 = new_n34811 ^ new_n34791;
  assign new_n34813 = new_n34812 ^ new_n34786;
  assign new_n34814 = new_n34813 ^ new_n34809;
  assign new_n34815 = new_n34775 ^ new_n34768;
  assign new_n34816 = new_n34755 ^ new_n34751;
  assign new_n34817 = new_n34815 & new_n34816;
  assign new_n34818 = new_n34817 ^ new_n34784;
  assign new_n34819 = new_n34811 ^ new_n34794;
  assign new_n34820 = new_n34819 ^ new_n34818;
  assign new_n34821 = ~new_n34820 & new_n34814;
  assign new_n34822 = new_n34775 ^ new_n34766;
  assign new_n34823 = new_n34803 ^ new_n34770;
  assign new_n34824 = new_n34823 ^ new_n34819;
  assign new_n34825 = new_n34824 ^ new_n34822;
  assign new_n34826 = new_n34817 ^ new_n34787;
  assign new_n34827 = new_n34826 ^ new_n34775;
  assign new_n34828 = new_n34827 ^ new_n34813;
  assign new_n34829 = new_n34828 ^ new_n34808;
  assign new_n34830 = new_n34825 & new_n34829;
  assign new_n34831 = new_n34830 ^ new_n34821;
  assign new_n34832 = new_n34827 ^ new_n34783;
  assign new_n34833 = new_n34832 ^ new_n34831;
  assign new_n34834 = new_n34751 & new_n34833;
  assign new_n34835 = new_n34821 ^ new_n34808;
  assign new_n34836 = new_n34828 & new_n34835;
  assign new_n34837 = new_n34836 ^ new_n34798;
  assign new_n34838 = ~new_n34837 & new_n34780;
  assign new_n34839 = new_n34838 ^ new_n34834;
  assign new_n34840 = new_n34766 ^ new_n34748;
  assign new_n34841 = new_n34803 ^ new_n34785;
  assign new_n34842 = new_n34830 ^ new_n34783;
  assign new_n34843 = new_n34842 ^ new_n34813;
  assign new_n34844 = new_n34836 ^ new_n34829;
  assign new_n34845 = new_n34843 & new_n34844;
  assign new_n34846 = new_n34845 ^ new_n34836;
  assign new_n34847 = new_n34846 ^ new_n34841;
  assign new_n34848 = new_n34847 ^ new_n34840;
  assign new_n34849 = new_n34848 ^ new_n34761;
  assign new_n34850 = new_n34830 ^ new_n34787;
  assign new_n34851 = new_n34850 ^ new_n34782;
  assign new_n34852 = new_n34851 ^ new_n34849;
  assign new_n34853 = ~new_n34852 & new_n34793;
  assign new_n34854 = new_n34845 ^ new_n34825;
  assign new_n34855 = new_n34768 & new_n34854;
  assign new_n34856 = new_n34836 ^ new_n34821;
  assign new_n34857 = new_n34856 ^ new_n34820;
  assign new_n34858 = ~new_n34857 & new_n34801;
  assign new_n34859 = ~new_n34852 & new_n34779;
  assign new_n34860 = new_n34776 & new_n34833;
  assign new_n34861 = new_n34860 ^ new_n34859;
  assign new_n34862 = new_n34861 ^ new_n34858;
  assign new_n34863 = new_n34862 ^ new_n34855;
  assign new_n34864 = new_n34845 ^ new_n34830;
  assign new_n34865 = new_n34864 ^ new_n34807;
  assign new_n34866 = new_n34786 & new_n34865;
  assign new_n34867 = new_n34866 ^ new_n34863;
  assign new_n34868 = new_n34867 ^ new_n34853;
  assign new_n34869 = new_n34868 ^ new_n34839;
  assign new_n34870 = new_n30119 ^ new_n26101;
  assign new_n34871 = new_n34870 ^ new_n34869;
  assign new_n34872 = new_n30128 ^ new_n26037;
  assign new_n34873 = new_n34853 ^ new_n34834;
  assign new_n34874 = ~new_n34837 & new_n34777;
  assign new_n34875 = ~new_n34857 & new_n34802;
  assign new_n34876 = new_n34875 ^ new_n34874;
  assign new_n34877 = new_n34876 ^ new_n34838;
  assign new_n34878 = new_n34877 ^ new_n34862;
  assign new_n34879 = new_n34878 ^ new_n34873;
  assign new_n34880 = new_n34879 ^ new_n34872;
  assign new_n34881 = new_n30154 ^ new_n26065;
  assign new_n34882 = new_n34860 ^ new_n34834;
  assign new_n34883 = new_n34821 ^ new_n34775;
  assign new_n34884 = new_n34817 ^ new_n34770;
  assign new_n34885 = new_n34884 ^ new_n34848;
  assign new_n34886 = new_n34885 ^ new_n34883;
  assign new_n34887 = ~new_n34886 & new_n34789;
  assign new_n34888 = new_n34778 & new_n34865;
  assign new_n34889 = new_n34828 ^ new_n34821;
  assign new_n34890 = new_n34755 & new_n34889;
  assign new_n34891 = new_n34890 ^ new_n34874;
  assign new_n34892 = new_n34891 ^ new_n34888;
  assign new_n34893 = ~new_n34886 & new_n34810;
  assign new_n34894 = new_n34815 & new_n34843;
  assign new_n34895 = new_n34894 ^ new_n34893;
  assign new_n34896 = new_n34895 ^ new_n34892;
  assign new_n34897 = new_n34896 ^ new_n34887;
  assign new_n34898 = new_n34897 ^ new_n34882;
  assign new_n34899 = new_n34898 ^ new_n34881;
  assign new_n34900 = new_n34877 ^ new_n34867;
  assign new_n34901 = new_n30175 ^ new_n26111;
  assign new_n34902 = new_n34901 ^ new_n34900;
  assign new_n34903 = new_n34816 & new_n34843;
  assign new_n34904 = new_n34903 ^ new_n34838;
  assign new_n34905 = new_n34890 ^ new_n34875;
  assign new_n34906 = new_n34905 ^ new_n34863;
  assign new_n34907 = new_n34906 ^ new_n34904;
  assign new_n34908 = new_n30187 ^ new_n26007;
  assign new_n34909 = new_n34908 ^ new_n34907;
  assign new_n34910 = new_n34769 & new_n34889;
  assign new_n34911 = new_n34910 ^ new_n34868;
  assign new_n34912 = new_n34911 ^ new_n34896;
  assign new_n34913 = new_n30195 ^ new_n25011;
  assign new_n34914 = new_n34913 ^ new_n34912;
  assign new_n34915 = new_n30204 ^ new_n25969;
  assign new_n34916 = new_n34893 ^ new_n34888;
  assign new_n34917 = new_n34800 & new_n34854;
  assign new_n34918 = new_n34917 ^ new_n34903;
  assign new_n34919 = new_n34918 ^ new_n34861;
  assign new_n34920 = new_n34855 ^ new_n34853;
  assign new_n34921 = new_n34920 ^ new_n34919;
  assign new_n34922 = new_n34921 ^ new_n34916;
  assign new_n34923 = new_n34922 ^ new_n34915;
  assign new_n34924 = new_n30215 ^ new_n26077;
  assign new_n34925 = new_n34892 ^ new_n34866;
  assign new_n34926 = new_n34925 ^ new_n34919;
  assign new_n34927 = new_n34926 ^ new_n34924;
  assign new_n34928 = new_n33532 ^ new_n33050;
  assign new_n34929 = new_n33325 ^ new_n32556;
  assign new_n34930 = new_n34929 ^ new_n33547;
  assign new_n34931 = new_n34930 ^ new_n34928;
  assign new_n34932 = new_n33426 ^ new_n32557;
  assign new_n34933 = new_n34295 ^ new_n33492;
  assign new_n34934 = new_n34933 ^ new_n34932;
  assign new_n34935 = new_n33471 ^ new_n32558;
  assign new_n34936 = new_n34935 ^ new_n33415;
  assign new_n34937 = new_n34302 ^ new_n33552;
  assign new_n34938 = new_n34937 ^ new_n34936;
  assign new_n34939 = new_n34308 ^ new_n33552;
  assign new_n34940 = new_n33435 ^ new_n32559;
  assign new_n34941 = new_n34940 ^ new_n33507;
  assign new_n34942 = new_n34941 ^ new_n34939;
  assign new_n34943 = new_n34942 ^ new_n34938;
  assign new_n34944 = new_n34943 ^ new_n34934;
  assign new_n34945 = new_n34944 ^ new_n34931;
  assign new_n34946 = new_n33495 ^ new_n32563;
  assign new_n34947 = new_n34317 ^ new_n33552;
  assign new_n34948 = new_n34947 ^ new_n34946;
  assign new_n34949 = new_n33448 ^ new_n32564;
  assign new_n34950 = new_n34949 ^ new_n33552;
  assign new_n34951 = new_n33536 ^ new_n33512;
  assign new_n34952 = new_n34951 ^ new_n33520;
  assign new_n34953 = new_n34952 ^ new_n34950;
  assign new_n34954 = new_n33527 ^ new_n33513;
  assign new_n34955 = new_n33345 ^ new_n32565;
  assign new_n34956 = new_n34955 ^ new_n32901;
  assign new_n34957 = new_n34956 ^ new_n34954;
  assign new_n34958 = new_n34957 ^ new_n34931;
  assign new_n34959 = new_n34958 ^ new_n34948;
  assign new_n34960 = new_n34959 ^ new_n34953;
  assign new_n34961 = new_n34948 & new_n34960;
  assign new_n34962 = new_n34961 ^ new_n34953;
  assign new_n34963 = new_n33191 ^ new_n32571;
  assign new_n34964 = new_n33551 ^ new_n33463;
  assign new_n34965 = new_n34964 ^ new_n34963;
  assign new_n34966 = new_n34965 ^ new_n34953;
  assign new_n34967 = new_n34966 ^ new_n34943;
  assign new_n34968 = new_n34953 ^ new_n34942;
  assign new_n34969 = new_n34965 ^ new_n34934;
  assign new_n34970 = new_n34969 ^ new_n34968;
  assign new_n34971 = new_n34967 & new_n34970;
  assign new_n34972 = new_n34971 ^ new_n34931;
  assign new_n34973 = new_n34972 ^ new_n34962;
  assign new_n34974 = ~new_n34942 & ~new_n34959;
  assign new_n34975 = new_n34974 ^ new_n34942;
  assign new_n34976 = new_n34957 ^ new_n34944;
  assign new_n34977 = new_n34965 ^ new_n34942;
  assign new_n34978 = new_n34976 & new_n34977;
  assign new_n34979 = new_n34978 ^ new_n34975;
  assign new_n34980 = new_n34979 ^ new_n34969;
  assign new_n34981 = new_n34945 & new_n34966;
  assign new_n34982 = new_n34957 ^ new_n34953;
  assign new_n34983 = new_n34982 ^ new_n34969;
  assign new_n34984 = new_n34953 ^ new_n34934;
  assign new_n34985 = new_n34983 & new_n34984;
  assign new_n34986 = new_n34985 ^ new_n34981;
  assign new_n34987 = new_n34957 ^ new_n34938;
  assign new_n34988 = new_n34987 ^ new_n34986;
  assign new_n34989 = new_n34988 ^ new_n34980;
  assign new_n34990 = new_n34972 ^ new_n34967;
  assign new_n34991 = new_n34959 ^ new_n34942;
  assign new_n34992 = new_n34991 ^ new_n34969;
  assign new_n34993 = new_n34967 ^ new_n34948;
  assign new_n34994 = new_n34992 & new_n34993;
  assign new_n34995 = new_n34994 ^ new_n34981;
  assign new_n34996 = new_n34985 ^ new_n34934;
  assign new_n34997 = new_n34996 ^ new_n34995;
  assign new_n34998 = new_n34997 ^ new_n34990;
  assign new_n34999 = ~new_n34989 & new_n34998;
  assign new_n35000 = new_n34999 ^ new_n34973;
  assign new_n35001 = new_n34967 ^ new_n34958;
  assign new_n35002 = new_n34969 & new_n35001;
  assign new_n35003 = new_n35002 ^ new_n34981;
  assign new_n35004 = new_n35003 ^ new_n34976;
  assign new_n35005 = new_n35004 ^ new_n35000;
  assign new_n35006 = new_n34965 ^ new_n34959;
  assign new_n35007 = new_n34948 ^ new_n34945;
  assign new_n35008 = new_n35006 & new_n35007;
  assign new_n35009 = new_n35008 ^ new_n34974;
  assign new_n35010 = new_n35002 ^ new_n34985;
  assign new_n35011 = new_n35010 ^ new_n35009;
  assign new_n35012 = ~new_n35011 & new_n35005;
  assign new_n35013 = new_n34965 ^ new_n34957;
  assign new_n35014 = new_n34994 ^ new_n34961;
  assign new_n35015 = new_n35014 ^ new_n35010;
  assign new_n35016 = new_n35015 ^ new_n35013;
  assign new_n35017 = new_n35008 ^ new_n34978;
  assign new_n35018 = new_n35017 ^ new_n34965;
  assign new_n35019 = new_n35018 ^ new_n35004;
  assign new_n35020 = new_n35019 ^ new_n34999;
  assign new_n35021 = new_n35016 & new_n35020;
  assign new_n35022 = new_n35021 ^ new_n35012;
  assign new_n35023 = new_n35018 ^ new_n34973;
  assign new_n35024 = new_n35023 ^ new_n35022;
  assign new_n35025 = new_n34945 & new_n35024;
  assign new_n35026 = new_n35012 ^ new_n34999;
  assign new_n35027 = new_n35019 & new_n35026;
  assign new_n35028 = new_n35027 ^ new_n34989;
  assign new_n35029 = ~new_n35028 & new_n34970;
  assign new_n35030 = new_n35029 ^ new_n35025;
  assign new_n35031 = new_n34957 ^ new_n34942;
  assign new_n35032 = new_n34994 ^ new_n34975;
  assign new_n35033 = new_n35021 ^ new_n34973;
  assign new_n35034 = new_n35033 ^ new_n35004;
  assign new_n35035 = new_n35027 ^ new_n35020;
  assign new_n35036 = new_n35034 & new_n35035;
  assign new_n35037 = new_n35036 ^ new_n35027;
  assign new_n35038 = new_n35037 ^ new_n35032;
  assign new_n35039 = new_n35038 ^ new_n35031;
  assign new_n35040 = new_n35039 ^ new_n34953;
  assign new_n35041 = new_n35021 ^ new_n34978;
  assign new_n35042 = new_n35041 ^ new_n34972;
  assign new_n35043 = new_n35042 ^ new_n35040;
  assign new_n35044 = ~new_n35043 & new_n34983;
  assign new_n35045 = new_n35036 ^ new_n35016;
  assign new_n35046 = new_n34959 & new_n35045;
  assign new_n35047 = new_n35027 ^ new_n35012;
  assign new_n35048 = new_n35047 ^ new_n35011;
  assign new_n35049 = ~new_n35048 & new_n34992;
  assign new_n35050 = ~new_n35043 & new_n34984;
  assign new_n35051 = new_n34966 & new_n35024;
  assign new_n35052 = new_n35051 ^ new_n35050;
  assign new_n35053 = new_n35052 ^ new_n35049;
  assign new_n35054 = new_n35053 ^ new_n35046;
  assign new_n35055 = new_n35036 ^ new_n35021;
  assign new_n35056 = new_n35055 ^ new_n34998;
  assign new_n35057 = new_n34976 & new_n35056;
  assign new_n35058 = new_n35057 ^ new_n35054;
  assign new_n35059 = new_n35058 ^ new_n35044;
  assign new_n35060 = new_n35059 ^ new_n35030;
  assign new_n35061 = new_n33067 ^ new_n31408;
  assign new_n35062 = new_n35061 ^ new_n35060;
  assign new_n35063 = new_n33081 ^ new_n31417;
  assign new_n35064 = new_n35044 ^ new_n35025;
  assign new_n35065 = ~new_n35028 & new_n34967;
  assign new_n35066 = ~new_n35048 & new_n34993;
  assign new_n35067 = new_n35066 ^ new_n35065;
  assign new_n35068 = new_n35067 ^ new_n35029;
  assign new_n35069 = new_n35068 ^ new_n35053;
  assign new_n35070 = new_n35069 ^ new_n35064;
  assign new_n35071 = new_n35070 ^ new_n35063;
  assign new_n35072 = new_n33057 ^ new_n31443;
  assign new_n35073 = new_n35051 ^ new_n35025;
  assign new_n35074 = new_n35012 ^ new_n34965;
  assign new_n35075 = new_n35008 ^ new_n34961;
  assign new_n35076 = new_n35075 ^ new_n35039;
  assign new_n35077 = new_n35076 ^ new_n35074;
  assign new_n35078 = ~new_n35077 & new_n34969;
  assign new_n35079 = new_n34977 & new_n35056;
  assign new_n35080 = new_n35019 ^ new_n35012;
  assign new_n35081 = new_n34948 & new_n35080;
  assign new_n35082 = new_n35081 ^ new_n35065;
  assign new_n35083 = new_n35082 ^ new_n35079;
  assign new_n35084 = ~new_n35077 & new_n35001;
  assign new_n35085 = new_n35006 & new_n35034;
  assign new_n35086 = new_n35085 ^ new_n35084;
  assign new_n35087 = new_n35086 ^ new_n35083;
  assign new_n35088 = new_n35087 ^ new_n35078;
  assign new_n35089 = new_n35088 ^ new_n35073;
  assign new_n35090 = new_n35089 ^ new_n35072;
  assign new_n35091 = new_n35068 ^ new_n35058;
  assign new_n35092 = new_n33051 ^ new_n31464;
  assign new_n35093 = new_n35092 ^ new_n35091;
  assign new_n35094 = new_n35007 & new_n35034;
  assign new_n35095 = new_n35094 ^ new_n35029;
  assign new_n35096 = new_n35081 ^ new_n35066;
  assign new_n35097 = new_n35096 ^ new_n35054;
  assign new_n35098 = new_n35097 ^ new_n35095;
  assign new_n35099 = new_n33099 ^ new_n31476;
  assign new_n35100 = new_n35099 ^ new_n35098;
  assign new_n35101 = new_n34960 & new_n35080;
  assign new_n35102 = new_n35101 ^ new_n35059;
  assign new_n35103 = new_n35102 ^ new_n35087;
  assign new_n35104 = new_n33064 ^ new_n31484;
  assign new_n35105 = new_n35104 ^ new_n35103;
  assign new_n35106 = new_n33075 ^ new_n31493;
  assign new_n35107 = new_n35084 ^ new_n35079;
  assign new_n35108 = new_n34991 & new_n35045;
  assign new_n35109 = new_n35108 ^ new_n35094;
  assign new_n35110 = new_n35109 ^ new_n35052;
  assign new_n35111 = new_n35046 ^ new_n35044;
  assign new_n35112 = new_n35111 ^ new_n35110;
  assign new_n35113 = new_n35112 ^ new_n35107;
  assign new_n35114 = new_n35113 ^ new_n35106;
  assign new_n35115 = new_n33087 ^ new_n31504;
  assign new_n35116 = new_n35083 ^ new_n35057;
  assign new_n35117 = new_n35116 ^ new_n35110;
  assign new_n35118 = new_n35117 ^ new_n35115;
  assign new_n35119 = new_n32033 ^ new_n27111;
  assign new_n35120 = new_n35119 ^ new_n19197;
  assign new_n35121 = new_n35120 ^ new_n29477;
  assign new_n35122 = new_n34498 ^ new_n29734;
  assign new_n35123 = new_n35122 ^ new_n35121;
  assign new_n35124 = new_n32296 ^ new_n27036;
  assign new_n35125 = new_n35124 ^ new_n19190;
  assign new_n35126 = new_n35125 ^ new_n29605;
  assign new_n35127 = new_n34505 ^ new_n29678;
  assign new_n35128 = new_n35127 ^ new_n35126;
  assign new_n35129 = new_n32341 ^ new_n27163;
  assign new_n35130 = new_n35129 ^ new_n19174;
  assign new_n35131 = new_n35130 ^ new_n29631;
  assign new_n35132 = new_n35131 ^ new_n29760;
  assign new_n35133 = new_n34516 ^ new_n29567;
  assign new_n35134 = new_n35133 ^ new_n35132;
  assign new_n35135 = new_n34521 ^ new_n29706;
  assign new_n35136 = new_n32380 ^ new_n27098;
  assign new_n35137 = new_n35136 ^ new_n19184;
  assign new_n35138 = new_n35137 ^ new_n29614;
  assign new_n35139 = new_n35138 ^ new_n29760;
  assign new_n35140 = new_n35139 ^ new_n35135;
  assign new_n35141 = new_n35140 ^ new_n35134;
  assign new_n35142 = new_n35141 ^ new_n35128;
  assign new_n35143 = new_n35142 ^ new_n35123;
  assign new_n35144 = new_n32392 ^ new_n27130;
  assign new_n35145 = new_n35144 ^ new_n19224;
  assign new_n35146 = new_n35145 ^ new_n29681;
  assign new_n35147 = new_n34535 ^ new_n29760;
  assign new_n35148 = new_n35147 ^ new_n35146;
  assign new_n35149 = new_n34540 ^ new_n29644;
  assign new_n35150 = new_n32404 ^ new_n26604;
  assign new_n35151 = new_n35150 ^ new_n19212;
  assign new_n35152 = new_n35151 ^ new_n29722;
  assign new_n35153 = new_n35152 ^ new_n29760;
  assign new_n35154 = new_n35153 ^ new_n35149;
  assign new_n35155 = new_n32431 ^ new_n26959;
  assign new_n35156 = new_n35155 ^ new_n19229;
  assign new_n35157 = new_n35156 ^ new_n29497;
  assign new_n35158 = new_n34546 ^ new_n29714;
  assign new_n35159 = new_n35158 ^ new_n35157;
  assign new_n35160 = new_n35159 ^ new_n35123;
  assign new_n35161 = new_n35160 ^ new_n35148;
  assign new_n35162 = new_n35161 ^ new_n35154;
  assign new_n35163 = new_n35148 & new_n35162;
  assign new_n35164 = new_n35163 ^ new_n35154;
  assign new_n35165 = new_n32455 ^ new_n27051;
  assign new_n35166 = new_n35165 ^ new_n19204;
  assign new_n35167 = new_n35166 ^ new_n29653;
  assign new_n35168 = new_n34558 ^ new_n28327;
  assign new_n35169 = new_n35168 ^ new_n35167;
  assign new_n35170 = new_n35169 ^ new_n35154;
  assign new_n35171 = new_n35170 ^ new_n35141;
  assign new_n35172 = new_n35154 ^ new_n35140;
  assign new_n35173 = new_n35169 ^ new_n35128;
  assign new_n35174 = new_n35173 ^ new_n35172;
  assign new_n35175 = new_n35171 & new_n35174;
  assign new_n35176 = new_n35175 ^ new_n35123;
  assign new_n35177 = new_n35176 ^ new_n35164;
  assign new_n35178 = ~new_n35140 & ~new_n35161;
  assign new_n35179 = new_n35178 ^ new_n35140;
  assign new_n35180 = new_n35159 ^ new_n35142;
  assign new_n35181 = new_n35169 ^ new_n35140;
  assign new_n35182 = new_n35180 & new_n35181;
  assign new_n35183 = new_n35182 ^ new_n35179;
  assign new_n35184 = new_n35183 ^ new_n35173;
  assign new_n35185 = new_n35143 & new_n35170;
  assign new_n35186 = new_n35159 ^ new_n35154;
  assign new_n35187 = new_n35186 ^ new_n35173;
  assign new_n35188 = new_n35154 ^ new_n35128;
  assign new_n35189 = new_n35187 & new_n35188;
  assign new_n35190 = new_n35189 ^ new_n35185;
  assign new_n35191 = new_n35159 ^ new_n35134;
  assign new_n35192 = new_n35191 ^ new_n35190;
  assign new_n35193 = new_n35192 ^ new_n35184;
  assign new_n35194 = new_n35176 ^ new_n35171;
  assign new_n35195 = new_n35161 ^ new_n35140;
  assign new_n35196 = new_n35195 ^ new_n35173;
  assign new_n35197 = new_n35171 ^ new_n35148;
  assign new_n35198 = new_n35196 & new_n35197;
  assign new_n35199 = new_n35198 ^ new_n35185;
  assign new_n35200 = new_n35189 ^ new_n35128;
  assign new_n35201 = new_n35200 ^ new_n35199;
  assign new_n35202 = new_n35201 ^ new_n35194;
  assign new_n35203 = ~new_n35193 & new_n35202;
  assign new_n35204 = new_n35203 ^ new_n35177;
  assign new_n35205 = new_n35171 ^ new_n35160;
  assign new_n35206 = new_n35173 & new_n35205;
  assign new_n35207 = new_n35206 ^ new_n35185;
  assign new_n35208 = new_n35207 ^ new_n35180;
  assign new_n35209 = new_n35208 ^ new_n35204;
  assign new_n35210 = new_n35169 ^ new_n35161;
  assign new_n35211 = new_n35148 ^ new_n35143;
  assign new_n35212 = new_n35210 & new_n35211;
  assign new_n35213 = new_n35212 ^ new_n35178;
  assign new_n35214 = new_n35206 ^ new_n35189;
  assign new_n35215 = new_n35214 ^ new_n35213;
  assign new_n35216 = ~new_n35215 & new_n35209;
  assign new_n35217 = new_n35169 ^ new_n35159;
  assign new_n35218 = new_n35198 ^ new_n35163;
  assign new_n35219 = new_n35218 ^ new_n35214;
  assign new_n35220 = new_n35219 ^ new_n35217;
  assign new_n35221 = new_n35212 ^ new_n35182;
  assign new_n35222 = new_n35221 ^ new_n35169;
  assign new_n35223 = new_n35222 ^ new_n35208;
  assign new_n35224 = new_n35223 ^ new_n35203;
  assign new_n35225 = new_n35220 & new_n35224;
  assign new_n35226 = new_n35225 ^ new_n35216;
  assign new_n35227 = new_n35222 ^ new_n35177;
  assign new_n35228 = new_n35227 ^ new_n35226;
  assign new_n35229 = new_n35143 & new_n35228;
  assign new_n35230 = new_n35216 ^ new_n35203;
  assign new_n35231 = new_n35223 & new_n35230;
  assign new_n35232 = new_n35231 ^ new_n35193;
  assign new_n35233 = ~new_n35232 & new_n35174;
  assign new_n35234 = new_n35233 ^ new_n35229;
  assign new_n35235 = new_n35159 ^ new_n35140;
  assign new_n35236 = new_n35198 ^ new_n35179;
  assign new_n35237 = new_n35225 ^ new_n35177;
  assign new_n35238 = new_n35237 ^ new_n35208;
  assign new_n35239 = new_n35231 ^ new_n35224;
  assign new_n35240 = new_n35238 & new_n35239;
  assign new_n35241 = new_n35240 ^ new_n35231;
  assign new_n35242 = new_n35241 ^ new_n35236;
  assign new_n35243 = new_n35242 ^ new_n35235;
  assign new_n35244 = new_n35243 ^ new_n35154;
  assign new_n35245 = new_n35225 ^ new_n35182;
  assign new_n35246 = new_n35245 ^ new_n35176;
  assign new_n35247 = new_n35246 ^ new_n35244;
  assign new_n35248 = ~new_n35247 & new_n35187;
  assign new_n35249 = new_n35240 ^ new_n35220;
  assign new_n35250 = new_n35161 & new_n35249;
  assign new_n35251 = new_n35231 ^ new_n35216;
  assign new_n35252 = new_n35251 ^ new_n35215;
  assign new_n35253 = ~new_n35252 & new_n35196;
  assign new_n35254 = ~new_n35247 & new_n35188;
  assign new_n35255 = new_n35170 & new_n35228;
  assign new_n35256 = new_n35255 ^ new_n35254;
  assign new_n35257 = new_n35256 ^ new_n35253;
  assign new_n35258 = new_n35257 ^ new_n35250;
  assign new_n35259 = new_n35240 ^ new_n35225;
  assign new_n35260 = new_n35259 ^ new_n35202;
  assign new_n35261 = new_n35180 & new_n35260;
  assign new_n35262 = new_n35261 ^ new_n35258;
  assign new_n35263 = new_n35262 ^ new_n35248;
  assign new_n35264 = new_n35263 ^ new_n35234;
  assign new_n35265 = new_n32665 ^ new_n32070;
  assign new_n35266 = new_n35265 ^ new_n35264;
  assign new_n35267 = new_n32674 ^ new_n32052;
  assign new_n35268 = new_n35248 ^ new_n35229;
  assign new_n35269 = ~new_n35232 & new_n35171;
  assign new_n35270 = ~new_n35252 & new_n35197;
  assign new_n35271 = new_n35270 ^ new_n35269;
  assign new_n35272 = new_n35271 ^ new_n35233;
  assign new_n35273 = new_n35272 ^ new_n35257;
  assign new_n35274 = new_n35273 ^ new_n35268;
  assign new_n35275 = new_n35274 ^ new_n35267;
  assign new_n35276 = new_n32700 ^ new_n32057;
  assign new_n35277 = new_n35255 ^ new_n35229;
  assign new_n35278 = new_n35216 ^ new_n35169;
  assign new_n35279 = new_n35212 ^ new_n35163;
  assign new_n35280 = new_n35279 ^ new_n35243;
  assign new_n35281 = new_n35280 ^ new_n35278;
  assign new_n35282 = ~new_n35281 & new_n35173;
  assign new_n35283 = new_n35181 & new_n35260;
  assign new_n35284 = new_n35223 ^ new_n35216;
  assign new_n35285 = new_n35148 & new_n35284;
  assign new_n35286 = new_n35285 ^ new_n35269;
  assign new_n35287 = new_n35286 ^ new_n35283;
  assign new_n35288 = ~new_n35281 & new_n35205;
  assign new_n35289 = new_n35210 & new_n35238;
  assign new_n35290 = new_n35289 ^ new_n35288;
  assign new_n35291 = new_n35290 ^ new_n35287;
  assign new_n35292 = new_n35291 ^ new_n35282;
  assign new_n35293 = new_n35292 ^ new_n35277;
  assign new_n35294 = new_n35293 ^ new_n35276;
  assign new_n35295 = new_n35272 ^ new_n35262;
  assign new_n35296 = new_n32721 ^ new_n32080;
  assign new_n35297 = new_n35296 ^ new_n35295;
  assign new_n35298 = new_n35211 & new_n35238;
  assign new_n35299 = new_n35298 ^ new_n35233;
  assign new_n35300 = new_n35285 ^ new_n35270;
  assign new_n35301 = new_n35300 ^ new_n35258;
  assign new_n35302 = new_n35301 ^ new_n35299;
  assign new_n35303 = new_n32733 ^ new_n32045;
  assign new_n35304 = new_n35303 ^ new_n35302;
  assign new_n35305 = new_n35162 & new_n35284;
  assign new_n35306 = new_n35305 ^ new_n35263;
  assign new_n35307 = new_n35306 ^ new_n35291;
  assign new_n35308 = new_n32741 ^ new_n32036;
  assign new_n35309 = new_n35308 ^ new_n35307;
  assign new_n35310 = new_n32750 ^ new_n32041;
  assign new_n35311 = new_n35288 ^ new_n35283;
  assign new_n35312 = new_n35195 & new_n35249;
  assign new_n35313 = new_n35312 ^ new_n35298;
  assign new_n35314 = new_n35313 ^ new_n35256;
  assign new_n35315 = new_n35250 ^ new_n35248;
  assign new_n35316 = new_n35315 ^ new_n35314;
  assign new_n35317 = new_n35316 ^ new_n35311;
  assign new_n35318 = new_n35317 ^ new_n35310;
  assign new_n35319 = new_n32761 ^ new_n32062;
  assign new_n35320 = new_n35287 ^ new_n35261;
  assign new_n35321 = new_n35320 ^ new_n35314;
  assign new_n35322 = new_n35321 ^ new_n35319;
  assign new_n35323 = new_n29963 ^ new_n25012;
  assign new_n35324 = new_n35323 ^ new_n30940;
  assign new_n35325 = new_n35324 ^ new_n31181;
  assign new_n35326 = new_n31196 ^ new_n31172;
  assign new_n35327 = new_n35326 ^ new_n35325;
  assign new_n35328 = new_n31115 ^ new_n31086;
  assign new_n35329 = new_n29989 ^ new_n25796;
  assign new_n35330 = new_n35329 ^ new_n30993;
  assign new_n35331 = new_n35330 ^ new_n31130;
  assign new_n35332 = new_n35331 ^ new_n35328;
  assign new_n35333 = new_n29995 ^ new_n25755;
  assign new_n35334 = new_n35333 ^ new_n31153;
  assign new_n35335 = new_n31201 ^ new_n31199;
  assign new_n35336 = new_n35335 ^ new_n35334;
  assign new_n35337 = new_n31068 ^ new_n30993;
  assign new_n35338 = new_n35337 ^ new_n30968;
  assign new_n35339 = new_n35338 ^ new_n35336;
  assign new_n35340 = new_n31139 ^ new_n31056;
  assign new_n35341 = new_n35340 ^ new_n35335;
  assign new_n35342 = new_n30003 ^ new_n25740;
  assign new_n35343 = new_n35342 ^ new_n31130;
  assign new_n35344 = new_n35343 ^ new_n31144;
  assign new_n35345 = new_n35344 ^ new_n35341;
  assign new_n35346 = new_n35345 ^ new_n35339;
  assign new_n35347 = new_n35346 ^ new_n35332;
  assign new_n35348 = new_n35347 ^ new_n35327;
  assign new_n35349 = new_n30009 ^ new_n25771;
  assign new_n35350 = new_n35349 ^ new_n31144;
  assign new_n35351 = new_n35335 ^ new_n31107;
  assign new_n35352 = new_n35351 ^ new_n35350;
  assign new_n35353 = new_n30011 ^ new_n25685;
  assign new_n35354 = new_n35353 ^ new_n31167;
  assign new_n35355 = new_n35354 ^ new_n35335;
  assign new_n35356 = new_n31158 ^ new_n31068;
  assign new_n35357 = new_n35356 ^ new_n31063;
  assign new_n35358 = new_n35357 ^ new_n35355;
  assign new_n35359 = new_n31181 ^ new_n30508;
  assign new_n35360 = new_n30016 ^ new_n25625;
  assign new_n35361 = new_n31159 ^ new_n31158;
  assign new_n35362 = new_n35361 ^ new_n35360;
  assign new_n35363 = new_n35362 ^ new_n35359;
  assign new_n35364 = new_n35363 ^ new_n35327;
  assign new_n35365 = new_n35364 ^ new_n35352;
  assign new_n35366 = new_n35365 ^ new_n35358;
  assign new_n35367 = ~new_n35366 & new_n35352;
  assign new_n35368 = new_n35367 ^ new_n35358;
  assign new_n35369 = new_n31098 ^ new_n30679;
  assign new_n35370 = new_n30024 ^ new_n25678;
  assign new_n35371 = new_n35370 ^ new_n31199;
  assign new_n35372 = new_n35371 ^ new_n30940;
  assign new_n35373 = new_n35372 ^ new_n35369;
  assign new_n35374 = new_n35373 ^ new_n35358;
  assign new_n35375 = new_n35374 ^ new_n35346;
  assign new_n35376 = new_n35358 ^ new_n35345;
  assign new_n35377 = new_n35373 ^ new_n35332;
  assign new_n35378 = new_n35377 ^ new_n35376;
  assign new_n35379 = new_n35375 & new_n35378;
  assign new_n35380 = new_n35379 ^ new_n35327;
  assign new_n35381 = new_n35380 ^ new_n35368;
  assign new_n35382 = new_n35345 & new_n35365;
  assign new_n35383 = new_n35382 ^ new_n35345;
  assign new_n35384 = new_n35363 ^ new_n35347;
  assign new_n35385 = new_n35373 ^ new_n35345;
  assign new_n35386 = ~new_n35384 & ~new_n35385;
  assign new_n35387 = new_n35386 ^ new_n35383;
  assign new_n35388 = new_n35387 ^ new_n35377;
  assign new_n35389 = new_n35348 & new_n35374;
  assign new_n35390 = new_n35363 ^ new_n35358;
  assign new_n35391 = new_n35390 ^ new_n35377;
  assign new_n35392 = new_n35358 ^ new_n35332;
  assign new_n35393 = ~new_n35391 & ~new_n35392;
  assign new_n35394 = new_n35393 ^ new_n35389;
  assign new_n35395 = new_n35363 ^ new_n35339;
  assign new_n35396 = new_n35395 ^ new_n35394;
  assign new_n35397 = new_n35396 ^ new_n35388;
  assign new_n35398 = new_n35380 ^ new_n35375;
  assign new_n35399 = new_n35365 ^ new_n35345;
  assign new_n35400 = new_n35399 ^ new_n35377;
  assign new_n35401 = new_n35375 ^ new_n35352;
  assign new_n35402 = ~new_n35400 & new_n35401;
  assign new_n35403 = new_n35402 ^ new_n35332;
  assign new_n35404 = new_n35403 ^ new_n35394;
  assign new_n35405 = new_n35404 ^ new_n35398;
  assign new_n35406 = new_n35397 & new_n35405;
  assign new_n35407 = new_n35406 ^ new_n35381;
  assign new_n35408 = new_n35375 ^ new_n35364;
  assign new_n35409 = ~new_n35377 & ~new_n35408;
  assign new_n35410 = new_n35409 ^ new_n35389;
  assign new_n35411 = new_n35410 ^ new_n35384;
  assign new_n35412 = new_n35411 ^ new_n35407;
  assign new_n35413 = new_n35373 ^ new_n35365;
  assign new_n35414 = new_n35352 ^ new_n35348;
  assign new_n35415 = ~new_n35413 & new_n35414;
  assign new_n35416 = new_n35415 ^ new_n35382;
  assign new_n35417 = new_n35409 ^ new_n35393;
  assign new_n35418 = new_n35417 ^ new_n35416;
  assign new_n35419 = ~new_n35418 & new_n35412;
  assign new_n35420 = new_n35373 ^ new_n35363;
  assign new_n35421 = new_n35402 ^ new_n35367;
  assign new_n35422 = new_n35421 ^ new_n35417;
  assign new_n35423 = new_n35422 ^ new_n35420;
  assign new_n35424 = new_n35415 ^ new_n35386;
  assign new_n35425 = new_n35424 ^ new_n35373;
  assign new_n35426 = new_n35425 ^ new_n35411;
  assign new_n35427 = new_n35426 ^ new_n35406;
  assign new_n35428 = ~new_n35427 & new_n35423;
  assign new_n35429 = new_n35428 ^ new_n35419;
  assign new_n35430 = new_n35425 ^ new_n35381;
  assign new_n35431 = new_n35430 ^ new_n35429;
  assign new_n35432 = ~new_n35431 & new_n35348;
  assign new_n35433 = new_n35419 ^ new_n35406;
  assign new_n35434 = ~new_n35426 & new_n35433;
  assign new_n35435 = new_n35434 ^ new_n35397;
  assign new_n35436 = new_n35378 & new_n35435;
  assign new_n35437 = new_n35436 ^ new_n35432;
  assign new_n35438 = new_n35363 ^ new_n35345;
  assign new_n35439 = new_n35402 ^ new_n35383;
  assign new_n35440 = new_n35428 ^ new_n35381;
  assign new_n35441 = new_n35440 ^ new_n35411;
  assign new_n35442 = new_n35434 ^ new_n35427;
  assign new_n35443 = ~new_n35442 & new_n35441;
  assign new_n35444 = new_n35443 ^ new_n35434;
  assign new_n35445 = new_n35444 ^ new_n35439;
  assign new_n35446 = new_n35445 ^ new_n35438;
  assign new_n35447 = new_n35446 ^ new_n35358;
  assign new_n35448 = new_n35428 ^ new_n35386;
  assign new_n35449 = new_n35448 ^ new_n35380;
  assign new_n35450 = new_n35449 ^ new_n35447;
  assign new_n35451 = ~new_n35391 & new_n35450;
  assign new_n35452 = new_n35443 ^ new_n35423;
  assign new_n35453 = ~new_n35365 & new_n35452;
  assign new_n35454 = new_n35434 ^ new_n35419;
  assign new_n35455 = new_n35454 ^ new_n35418;
  assign new_n35456 = ~new_n35400 & ~new_n35455;
  assign new_n35457 = ~new_n35392 & new_n35450;
  assign new_n35458 = ~new_n35431 & new_n35374;
  assign new_n35459 = new_n35458 ^ new_n35457;
  assign new_n35460 = new_n35459 ^ new_n35456;
  assign new_n35461 = new_n35460 ^ new_n35453;
  assign new_n35462 = new_n35443 ^ new_n35428;
  assign new_n35463 = new_n35462 ^ new_n35405;
  assign new_n35464 = ~new_n35384 & new_n35463;
  assign new_n35465 = new_n35464 ^ new_n35461;
  assign new_n35466 = new_n35465 ^ new_n35451;
  assign new_n35467 = new_n35466 ^ new_n35437;
  assign new_n35468 = new_n33761 ^ new_n30551;
  assign new_n35469 = new_n35468 ^ new_n35467;
  assign new_n35470 = new_n33770 ^ new_n30567;
  assign new_n35471 = new_n35451 ^ new_n35432;
  assign new_n35472 = new_n35375 & new_n35435;
  assign new_n35473 = ~new_n35455 & new_n35401;
  assign new_n35474 = new_n35473 ^ new_n35472;
  assign new_n35475 = new_n35474 ^ new_n35436;
  assign new_n35476 = new_n35475 ^ new_n35460;
  assign new_n35477 = new_n35476 ^ new_n35471;
  assign new_n35478 = new_n35477 ^ new_n35470;
  assign new_n35479 = new_n33796 ^ new_n30536;
  assign new_n35480 = new_n35458 ^ new_n35432;
  assign new_n35481 = new_n35419 ^ new_n35373;
  assign new_n35482 = new_n35415 ^ new_n35367;
  assign new_n35483 = new_n35482 ^ new_n35446;
  assign new_n35484 = new_n35483 ^ new_n35481;
  assign new_n35485 = ~new_n35377 & ~new_n35484;
  assign new_n35486 = ~new_n35385 & new_n35463;
  assign new_n35487 = new_n35426 ^ new_n35419;
  assign new_n35488 = ~new_n35487 & new_n35352;
  assign new_n35489 = new_n35488 ^ new_n35472;
  assign new_n35490 = new_n35489 ^ new_n35486;
  assign new_n35491 = ~new_n35408 & ~new_n35484;
  assign new_n35492 = ~new_n35413 & new_n35441;
  assign new_n35493 = new_n35492 ^ new_n35491;
  assign new_n35494 = new_n35493 ^ new_n35490;
  assign new_n35495 = new_n35494 ^ new_n35485;
  assign new_n35496 = new_n35495 ^ new_n35480;
  assign new_n35497 = new_n35496 ^ new_n35479;
  assign new_n35498 = new_n35475 ^ new_n35465;
  assign new_n35499 = new_n33817 ^ new_n30528;
  assign new_n35500 = new_n35499 ^ new_n35498;
  assign new_n35501 = new_n35414 & new_n35441;
  assign new_n35502 = new_n35501 ^ new_n35436;
  assign new_n35503 = new_n35488 ^ new_n35473;
  assign new_n35504 = new_n35503 ^ new_n35461;
  assign new_n35505 = new_n35504 ^ new_n35502;
  assign new_n35506 = new_n33829 ^ new_n30583;
  assign new_n35507 = new_n35506 ^ new_n35505;
  assign new_n35508 = ~new_n35366 & ~new_n35487;
  assign new_n35509 = new_n35508 ^ new_n35466;
  assign new_n35510 = new_n35509 ^ new_n35494;
  assign new_n35511 = new_n33837 ^ new_n30545;
  assign new_n35512 = new_n35511 ^ new_n35510;
  assign new_n35513 = new_n33846 ^ new_n30560;
  assign new_n35514 = new_n35491 ^ new_n35486;
  assign new_n35515 = new_n35399 & new_n35452;
  assign new_n35516 = new_n35515 ^ new_n35501;
  assign new_n35517 = new_n35516 ^ new_n35459;
  assign new_n35518 = new_n35453 ^ new_n35451;
  assign new_n35519 = new_n35518 ^ new_n35517;
  assign new_n35520 = new_n35519 ^ new_n35514;
  assign new_n35521 = new_n35520 ^ new_n35513;
  assign new_n35522 = new_n33857 ^ new_n30572;
  assign new_n35523 = new_n35490 ^ new_n35464;
  assign new_n35524 = new_n35523 ^ new_n35517;
  assign new_n35525 = new_n35524 ^ new_n35522;
  assign new_n35526 = new_n34335 ^ new_n33527;
  assign new_n35527 = new_n33547 ^ new_n31299;
  assign new_n35528 = new_n35527 ^ new_n32901;
  assign new_n35529 = new_n35528 ^ new_n35526;
  assign new_n35530 = new_n34308 ^ new_n31300;
  assign new_n35531 = new_n33467 ^ new_n33389;
  assign new_n35532 = new_n35531 ^ new_n33426;
  assign new_n35533 = new_n35532 ^ new_n35530;
  assign new_n35534 = new_n33551 ^ new_n33460;
  assign new_n35535 = new_n35534 ^ new_n31301;
  assign new_n35536 = new_n35535 ^ new_n34295;
  assign new_n35537 = new_n34322 ^ new_n33519;
  assign new_n35538 = new_n35537 ^ new_n35536;
  assign new_n35539 = new_n35534 ^ new_n33364;
  assign new_n35540 = new_n35539 ^ new_n34317;
  assign new_n35541 = new_n33491 ^ new_n31302;
  assign new_n35542 = new_n35541 ^ new_n33435;
  assign new_n35543 = new_n35542 ^ new_n35540;
  assign new_n35544 = new_n35543 ^ new_n35538;
  assign new_n35545 = new_n35544 ^ new_n35533;
  assign new_n35546 = new_n35545 ^ new_n35529;
  assign new_n35547 = new_n35534 ^ new_n33476;
  assign new_n35548 = new_n33506 ^ new_n31306;
  assign new_n35549 = new_n35548 ^ new_n33495;
  assign new_n35550 = new_n35549 ^ new_n35547;
  assign new_n35551 = new_n35534 ^ new_n34326;
  assign new_n35552 = new_n33536 ^ new_n31307;
  assign new_n35553 = new_n35552 ^ new_n34302;
  assign new_n35554 = new_n35553 ^ new_n35551;
  assign new_n35555 = new_n34292 ^ new_n32901;
  assign new_n35556 = new_n34951 ^ new_n31308;
  assign new_n35557 = new_n35556 ^ new_n35555;
  assign new_n35558 = new_n35557 ^ new_n35529;
  assign new_n35559 = new_n35558 ^ new_n35550;
  assign new_n35560 = new_n35559 ^ new_n35554;
  assign new_n35561 = new_n35550 & new_n35560;
  assign new_n35562 = new_n35561 ^ new_n35554;
  assign new_n35563 = new_n34303 ^ new_n33050;
  assign new_n35564 = new_n33460 ^ new_n31314;
  assign new_n35565 = new_n35564 ^ new_n33547;
  assign new_n35566 = new_n35565 ^ new_n35563;
  assign new_n35567 = new_n35566 ^ new_n35554;
  assign new_n35568 = new_n35567 ^ new_n35544;
  assign new_n35569 = new_n35554 ^ new_n35543;
  assign new_n35570 = new_n35566 ^ new_n35533;
  assign new_n35571 = new_n35570 ^ new_n35569;
  assign new_n35572 = new_n35568 & new_n35571;
  assign new_n35573 = new_n35572 ^ new_n35529;
  assign new_n35574 = new_n35573 ^ new_n35562;
  assign new_n35575 = ~new_n35543 & ~new_n35559;
  assign new_n35576 = new_n35575 ^ new_n35543;
  assign new_n35577 = new_n35557 ^ new_n35545;
  assign new_n35578 = new_n35566 ^ new_n35543;
  assign new_n35579 = new_n35577 & new_n35578;
  assign new_n35580 = new_n35579 ^ new_n35576;
  assign new_n35581 = new_n35580 ^ new_n35570;
  assign new_n35582 = new_n35546 & new_n35567;
  assign new_n35583 = new_n35557 ^ new_n35554;
  assign new_n35584 = new_n35583 ^ new_n35570;
  assign new_n35585 = new_n35554 ^ new_n35533;
  assign new_n35586 = new_n35584 & new_n35585;
  assign new_n35587 = new_n35586 ^ new_n35582;
  assign new_n35588 = new_n35557 ^ new_n35538;
  assign new_n35589 = new_n35588 ^ new_n35587;
  assign new_n35590 = new_n35589 ^ new_n35581;
  assign new_n35591 = new_n35573 ^ new_n35568;
  assign new_n35592 = new_n35559 ^ new_n35543;
  assign new_n35593 = new_n35592 ^ new_n35570;
  assign new_n35594 = new_n35568 ^ new_n35550;
  assign new_n35595 = new_n35593 & new_n35594;
  assign new_n35596 = new_n35595 ^ new_n35582;
  assign new_n35597 = new_n35586 ^ new_n35533;
  assign new_n35598 = new_n35597 ^ new_n35596;
  assign new_n35599 = new_n35598 ^ new_n35591;
  assign new_n35600 = ~new_n35590 & new_n35599;
  assign new_n35601 = new_n35600 ^ new_n35574;
  assign new_n35602 = new_n35568 ^ new_n35558;
  assign new_n35603 = new_n35570 & new_n35602;
  assign new_n35604 = new_n35603 ^ new_n35582;
  assign new_n35605 = new_n35604 ^ new_n35577;
  assign new_n35606 = new_n35605 ^ new_n35601;
  assign new_n35607 = new_n35566 ^ new_n35559;
  assign new_n35608 = new_n35550 ^ new_n35546;
  assign new_n35609 = new_n35607 & new_n35608;
  assign new_n35610 = new_n35609 ^ new_n35575;
  assign new_n35611 = new_n35603 ^ new_n35586;
  assign new_n35612 = new_n35611 ^ new_n35610;
  assign new_n35613 = ~new_n35612 & new_n35606;
  assign new_n35614 = new_n35566 ^ new_n35557;
  assign new_n35615 = new_n35595 ^ new_n35561;
  assign new_n35616 = new_n35615 ^ new_n35611;
  assign new_n35617 = new_n35616 ^ new_n35614;
  assign new_n35618 = new_n35609 ^ new_n35579;
  assign new_n35619 = new_n35618 ^ new_n35566;
  assign new_n35620 = new_n35619 ^ new_n35605;
  assign new_n35621 = new_n35620 ^ new_n35600;
  assign new_n35622 = new_n35617 & new_n35621;
  assign new_n35623 = new_n35622 ^ new_n35613;
  assign new_n35624 = new_n35619 ^ new_n35574;
  assign new_n35625 = new_n35624 ^ new_n35623;
  assign new_n35626 = new_n35546 & new_n35625;
  assign new_n35627 = new_n35613 ^ new_n35600;
  assign new_n35628 = new_n35620 & new_n35627;
  assign new_n35629 = new_n35628 ^ new_n35590;
  assign new_n35630 = ~new_n35629 & new_n35571;
  assign new_n35631 = new_n35630 ^ new_n35626;
  assign new_n35632 = new_n35557 ^ new_n35543;
  assign new_n35633 = new_n35595 ^ new_n35576;
  assign new_n35634 = new_n35622 ^ new_n35574;
  assign new_n35635 = new_n35634 ^ new_n35605;
  assign new_n35636 = new_n35628 ^ new_n35621;
  assign new_n35637 = new_n35635 & new_n35636;
  assign new_n35638 = new_n35637 ^ new_n35628;
  assign new_n35639 = new_n35638 ^ new_n35633;
  assign new_n35640 = new_n35639 ^ new_n35632;
  assign new_n35641 = new_n35640 ^ new_n35554;
  assign new_n35642 = new_n35622 ^ new_n35579;
  assign new_n35643 = new_n35642 ^ new_n35573;
  assign new_n35644 = new_n35643 ^ new_n35641;
  assign new_n35645 = ~new_n35644 & new_n35584;
  assign new_n35646 = new_n35637 ^ new_n35617;
  assign new_n35647 = new_n35559 & new_n35646;
  assign new_n35648 = new_n35628 ^ new_n35613;
  assign new_n35649 = new_n35648 ^ new_n35612;
  assign new_n35650 = ~new_n35649 & new_n35593;
  assign new_n35651 = ~new_n35644 & new_n35585;
  assign new_n35652 = new_n35567 & new_n35625;
  assign new_n35653 = new_n35652 ^ new_n35651;
  assign new_n35654 = new_n35653 ^ new_n35650;
  assign new_n35655 = new_n35654 ^ new_n35647;
  assign new_n35656 = new_n35637 ^ new_n35622;
  assign new_n35657 = new_n35656 ^ new_n35599;
  assign new_n35658 = new_n35577 & new_n35657;
  assign new_n35659 = new_n35658 ^ new_n35655;
  assign new_n35660 = new_n35659 ^ new_n35645;
  assign new_n35661 = new_n35660 ^ new_n35631;
  assign new_n35662 = new_n34772 ^ new_n30119;
  assign new_n35663 = new_n35662 ^ new_n35661;
  assign new_n35664 = new_n34727 ^ new_n30128;
  assign new_n35665 = new_n35645 ^ new_n35626;
  assign new_n35666 = ~new_n35629 & new_n35568;
  assign new_n35667 = ~new_n35649 & new_n35594;
  assign new_n35668 = new_n35667 ^ new_n35666;
  assign new_n35669 = new_n35668 ^ new_n35630;
  assign new_n35670 = new_n35669 ^ new_n35654;
  assign new_n35671 = new_n35670 ^ new_n35665;
  assign new_n35672 = new_n35671 ^ new_n35664;
  assign new_n35673 = new_n34763 ^ new_n30154;
  assign new_n35674 = new_n35652 ^ new_n35626;
  assign new_n35675 = new_n35613 ^ new_n35566;
  assign new_n35676 = new_n35609 ^ new_n35561;
  assign new_n35677 = new_n35676 ^ new_n35640;
  assign new_n35678 = new_n35677 ^ new_n35675;
  assign new_n35679 = ~new_n35678 & new_n35570;
  assign new_n35680 = new_n35578 & new_n35657;
  assign new_n35681 = new_n35620 ^ new_n35613;
  assign new_n35682 = new_n35550 & new_n35681;
  assign new_n35683 = new_n35682 ^ new_n35666;
  assign new_n35684 = new_n35683 ^ new_n35680;
  assign new_n35685 = ~new_n35678 & new_n35602;
  assign new_n35686 = new_n35607 & new_n35635;
  assign new_n35687 = new_n35686 ^ new_n35685;
  assign new_n35688 = new_n35687 ^ new_n35684;
  assign new_n35689 = new_n35688 ^ new_n35679;
  assign new_n35690 = new_n35689 ^ new_n35674;
  assign new_n35691 = new_n35690 ^ new_n35673;
  assign new_n35692 = new_n35669 ^ new_n35659;
  assign new_n35693 = new_n34756 ^ new_n30175;
  assign new_n35694 = new_n35693 ^ new_n35692;
  assign new_n35695 = new_n35608 & new_n35635;
  assign new_n35696 = new_n35695 ^ new_n35630;
  assign new_n35697 = new_n35682 ^ new_n35667;
  assign new_n35698 = new_n35697 ^ new_n35655;
  assign new_n35699 = new_n35698 ^ new_n35696;
  assign new_n35700 = new_n34738 ^ new_n30187;
  assign new_n35701 = new_n35700 ^ new_n35699;
  assign new_n35702 = new_n35560 & new_n35681;
  assign new_n35703 = new_n35702 ^ new_n35660;
  assign new_n35704 = new_n35703 ^ new_n35688;
  assign new_n35705 = new_n34733 ^ new_n30195;
  assign new_n35706 = new_n35705 ^ new_n35704;
  assign new_n35707 = new_n34745 ^ new_n30204;
  assign new_n35708 = new_n35685 ^ new_n35680;
  assign new_n35709 = new_n35592 & new_n35646;
  assign new_n35710 = new_n35709 ^ new_n35695;
  assign new_n35711 = new_n35710 ^ new_n35653;
  assign new_n35712 = new_n35647 ^ new_n35645;
  assign new_n35713 = new_n35712 ^ new_n35711;
  assign new_n35714 = new_n35713 ^ new_n35708;
  assign new_n35715 = new_n35714 ^ new_n35707;
  assign new_n35716 = new_n34752 ^ new_n30215;
  assign new_n35717 = new_n35684 ^ new_n35658;
  assign new_n35718 = new_n35717 ^ new_n35711;
  assign new_n35719 = new_n35718 ^ new_n35716;
  assign new_n35720 = new_n34546 ^ new_n27255;
  assign new_n35721 = new_n30788 ^ new_n28178;
  assign new_n35722 = new_n35721 ^ new_n15128;
  assign new_n35723 = new_n35722 ^ new_n29477;
  assign new_n35724 = new_n35723 ^ new_n29755;
  assign new_n35725 = new_n35724 ^ new_n35720;
  assign new_n35726 = new_n29627 ^ new_n29541;
  assign new_n35727 = new_n35726 ^ new_n29605;
  assign new_n35728 = new_n31029 ^ new_n28100;
  assign new_n35729 = new_n35728 ^ new_n14081;
  assign new_n35730 = new_n35729 ^ new_n34521;
  assign new_n35731 = new_n35730 ^ new_n35727;
  assign new_n35732 = new_n29721 ^ new_n29638;
  assign new_n35733 = new_n35732 ^ new_n29631;
  assign new_n35734 = new_n31091 ^ new_n28222;
  assign new_n35735 = new_n35734 ^ new_n15037;
  assign new_n35736 = new_n35735 ^ new_n34558;
  assign new_n35737 = new_n35736 ^ new_n34505;
  assign new_n35738 = new_n35737 ^ new_n35733;
  assign new_n35739 = new_n34558 ^ new_n29670;
  assign new_n35740 = new_n35739 ^ new_n34535;
  assign new_n35741 = new_n31122 ^ new_n28158;
  assign new_n35742 = new_n35741 ^ new_n15092;
  assign new_n35743 = new_n35742 ^ new_n29614;
  assign new_n35744 = new_n35743 ^ new_n29516;
  assign new_n35745 = new_n35744 ^ new_n35740;
  assign new_n35746 = new_n35745 ^ new_n35738;
  assign new_n35747 = new_n35746 ^ new_n35731;
  assign new_n35748 = new_n35747 ^ new_n35725;
  assign new_n35749 = new_n34558 ^ new_n29703;
  assign new_n35750 = new_n31141 ^ new_n28200;
  assign new_n35751 = new_n35750 ^ new_n15208;
  assign new_n35752 = new_n35751 ^ new_n29681;
  assign new_n35753 = new_n35752 ^ new_n29662;
  assign new_n35754 = new_n35753 ^ new_n35749;
  assign new_n35755 = new_n31154 ^ new_n27966;
  assign new_n35756 = new_n35755 ^ new_n15187;
  assign new_n35757 = new_n35756 ^ new_n34558;
  assign new_n35758 = new_n35757 ^ new_n34516;
  assign new_n35759 = new_n29745 ^ new_n29712;
  assign new_n35760 = new_n35759 ^ new_n35758;
  assign new_n35761 = new_n34540 ^ new_n29729;
  assign new_n35762 = new_n31176 ^ new_n28022;
  assign new_n35763 = new_n35762 ^ new_n15176;
  assign new_n35764 = new_n35763 ^ new_n29497;
  assign new_n35765 = new_n35764 ^ new_n26210;
  assign new_n35766 = new_n35765 ^ new_n35761;
  assign new_n35767 = new_n35766 ^ new_n35725;
  assign new_n35768 = new_n35767 ^ new_n35754;
  assign new_n35769 = new_n35768 ^ new_n35760;
  assign new_n35770 = new_n35754 & new_n35769;
  assign new_n35771 = new_n35770 ^ new_n35760;
  assign new_n35772 = new_n31191 ^ new_n28116;
  assign new_n35773 = new_n35772 ^ new_n15147;
  assign new_n35774 = new_n35773 ^ new_n34498;
  assign new_n35775 = new_n29757 ^ new_n29657;
  assign new_n35776 = new_n35775 ^ new_n35774;
  assign new_n35777 = new_n35776 ^ new_n35760;
  assign new_n35778 = new_n35777 ^ new_n35746;
  assign new_n35779 = new_n35776 ^ new_n35745;
  assign new_n35780 = new_n35760 ^ new_n35731;
  assign new_n35781 = new_n35780 ^ new_n35779;
  assign new_n35782 = new_n35778 & new_n35781;
  assign new_n35783 = new_n35782 ^ new_n35725;
  assign new_n35784 = new_n35783 ^ new_n35771;
  assign new_n35785 = ~new_n35745 & ~new_n35768;
  assign new_n35786 = new_n35785 ^ new_n35745;
  assign new_n35787 = new_n35766 ^ new_n35747;
  assign new_n35788 = new_n35779 & new_n35787;
  assign new_n35789 = new_n35788 ^ new_n35786;
  assign new_n35790 = new_n35776 ^ new_n35731;
  assign new_n35791 = new_n35790 ^ new_n35789;
  assign new_n35792 = new_n35748 & new_n35777;
  assign new_n35793 = new_n35766 ^ new_n35760;
  assign new_n35794 = new_n35793 ^ new_n35790;
  assign new_n35795 = new_n35780 & new_n35794;
  assign new_n35796 = new_n35795 ^ new_n35792;
  assign new_n35797 = new_n35766 ^ new_n35738;
  assign new_n35798 = new_n35797 ^ new_n35796;
  assign new_n35799 = new_n35798 ^ new_n35791;
  assign new_n35800 = new_n35783 ^ new_n35778;
  assign new_n35801 = new_n35768 ^ new_n35745;
  assign new_n35802 = new_n35801 ^ new_n35790;
  assign new_n35803 = new_n35778 ^ new_n35754;
  assign new_n35804 = new_n35802 & new_n35803;
  assign new_n35805 = new_n35804 ^ new_n35792;
  assign new_n35806 = new_n35795 ^ new_n35731;
  assign new_n35807 = new_n35806 ^ new_n35805;
  assign new_n35808 = new_n35807 ^ new_n35800;
  assign new_n35809 = ~new_n35799 & new_n35808;
  assign new_n35810 = new_n35809 ^ new_n35784;
  assign new_n35811 = new_n35778 ^ new_n35767;
  assign new_n35812 = new_n35790 & new_n35811;
  assign new_n35813 = new_n35812 ^ new_n35792;
  assign new_n35814 = new_n35813 ^ new_n35787;
  assign new_n35815 = new_n35814 ^ new_n35810;
  assign new_n35816 = new_n35776 ^ new_n35768;
  assign new_n35817 = new_n35754 ^ new_n35748;
  assign new_n35818 = new_n35816 & new_n35817;
  assign new_n35819 = new_n35818 ^ new_n35785;
  assign new_n35820 = new_n35812 ^ new_n35795;
  assign new_n35821 = new_n35820 ^ new_n35819;
  assign new_n35822 = ~new_n35821 & new_n35815;
  assign new_n35823 = new_n35776 ^ new_n35766;
  assign new_n35824 = new_n35804 ^ new_n35770;
  assign new_n35825 = new_n35824 ^ new_n35820;
  assign new_n35826 = new_n35825 ^ new_n35823;
  assign new_n35827 = new_n35818 ^ new_n35788;
  assign new_n35828 = new_n35827 ^ new_n35776;
  assign new_n35829 = new_n35828 ^ new_n35814;
  assign new_n35830 = new_n35829 ^ new_n35809;
  assign new_n35831 = new_n35826 & new_n35830;
  assign new_n35832 = new_n35831 ^ new_n35822;
  assign new_n35833 = new_n35828 ^ new_n35784;
  assign new_n35834 = new_n35833 ^ new_n35832;
  assign new_n35835 = new_n35748 & new_n35834;
  assign new_n35836 = new_n35822 ^ new_n35809;
  assign new_n35837 = new_n35829 & new_n35836;
  assign new_n35838 = new_n35837 ^ new_n35799;
  assign new_n35839 = ~new_n35838 & new_n35781;
  assign new_n35840 = new_n35839 ^ new_n35835;
  assign new_n35841 = new_n35766 ^ new_n35745;
  assign new_n35842 = new_n35804 ^ new_n35786;
  assign new_n35843 = new_n35831 ^ new_n35784;
  assign new_n35844 = new_n35843 ^ new_n35814;
  assign new_n35845 = new_n35837 ^ new_n35830;
  assign new_n35846 = new_n35844 & new_n35845;
  assign new_n35847 = new_n35846 ^ new_n35837;
  assign new_n35848 = new_n35847 ^ new_n35842;
  assign new_n35849 = new_n35848 ^ new_n35841;
  assign new_n35850 = new_n35849 ^ new_n35760;
  assign new_n35851 = new_n35831 ^ new_n35788;
  assign new_n35852 = new_n35851 ^ new_n35783;
  assign new_n35853 = new_n35852 ^ new_n35850;
  assign new_n35854 = ~new_n35853 & new_n35794;
  assign new_n35855 = new_n35846 ^ new_n35826;
  assign new_n35856 = new_n35768 & new_n35855;
  assign new_n35857 = new_n35837 ^ new_n35822;
  assign new_n35858 = new_n35857 ^ new_n35821;
  assign new_n35859 = ~new_n35858 & new_n35802;
  assign new_n35860 = ~new_n35853 & new_n35780;
  assign new_n35861 = new_n35777 & new_n35834;
  assign new_n35862 = new_n35861 ^ new_n35860;
  assign new_n35863 = new_n35862 ^ new_n35859;
  assign new_n35864 = new_n35863 ^ new_n35856;
  assign new_n35865 = new_n35846 ^ new_n35831;
  assign new_n35866 = new_n35865 ^ new_n35808;
  assign new_n35867 = new_n35787 & new_n35866;
  assign new_n35868 = new_n35867 ^ new_n35864;
  assign new_n35869 = new_n35868 ^ new_n35854;
  assign new_n35870 = new_n35869 ^ new_n35840;
  assign new_n35871 = new_n34125 ^ new_n31408;
  assign new_n35872 = new_n35871 ^ new_n35870;
  assign new_n35873 = new_n34079 ^ new_n31417;
  assign new_n35874 = new_n35854 ^ new_n35835;
  assign new_n35875 = ~new_n35838 & new_n35778;
  assign new_n35876 = ~new_n35858 & new_n35803;
  assign new_n35877 = new_n35876 ^ new_n35875;
  assign new_n35878 = new_n35877 ^ new_n35839;
  assign new_n35879 = new_n35878 ^ new_n35863;
  assign new_n35880 = new_n35879 ^ new_n35874;
  assign new_n35881 = new_n35880 ^ new_n35873;
  assign new_n35882 = new_n34115 ^ new_n31443;
  assign new_n35883 = new_n35861 ^ new_n35835;
  assign new_n35884 = new_n35822 ^ new_n35776;
  assign new_n35885 = new_n35818 ^ new_n35770;
  assign new_n35886 = new_n35885 ^ new_n35849;
  assign new_n35887 = new_n35886 ^ new_n35884;
  assign new_n35888 = ~new_n35887 & new_n35790;
  assign new_n35889 = new_n35779 & new_n35866;
  assign new_n35890 = new_n35829 ^ new_n35822;
  assign new_n35891 = new_n35754 & new_n35890;
  assign new_n35892 = new_n35891 ^ new_n35875;
  assign new_n35893 = new_n35892 ^ new_n35889;
  assign new_n35894 = ~new_n35887 & new_n35811;
  assign new_n35895 = new_n35816 & new_n35844;
  assign new_n35896 = new_n35895 ^ new_n35894;
  assign new_n35897 = new_n35896 ^ new_n35893;
  assign new_n35898 = new_n35897 ^ new_n35888;
  assign new_n35899 = new_n35898 ^ new_n35883;
  assign new_n35900 = new_n35899 ^ new_n35882;
  assign new_n35901 = new_n35878 ^ new_n35868;
  assign new_n35902 = new_n34111 ^ new_n31464;
  assign new_n35903 = new_n35902 ^ new_n35901;
  assign new_n35904 = new_n35817 & new_n35844;
  assign new_n35905 = new_n35904 ^ new_n35839;
  assign new_n35906 = new_n35891 ^ new_n35876;
  assign new_n35907 = new_n35906 ^ new_n35864;
  assign new_n35908 = new_n35907 ^ new_n35905;
  assign new_n35909 = new_n34088 ^ new_n31476;
  assign new_n35910 = new_n35909 ^ new_n35908;
  assign new_n35911 = new_n35769 & new_n35890;
  assign new_n35912 = new_n35911 ^ new_n35869;
  assign new_n35913 = new_n35912 ^ new_n35897;
  assign new_n35914 = new_n34084 ^ new_n31484;
  assign new_n35915 = new_n35914 ^ new_n35913;
  assign new_n35916 = new_n34097 ^ new_n31493;
  assign new_n35917 = new_n35894 ^ new_n35889;
  assign new_n35918 = new_n35801 & new_n35855;
  assign new_n35919 = new_n35918 ^ new_n35904;
  assign new_n35920 = new_n35919 ^ new_n35862;
  assign new_n35921 = new_n35856 ^ new_n35854;
  assign new_n35922 = new_n35921 ^ new_n35920;
  assign new_n35923 = new_n35922 ^ new_n35917;
  assign new_n35924 = new_n35923 ^ new_n35916;
  assign new_n35925 = new_n34104 ^ new_n31504;
  assign new_n35926 = new_n35893 ^ new_n35867;
  assign new_n35927 = new_n35926 ^ new_n35920;
  assign new_n35928 = new_n35927 ^ new_n35925;
  assign new_n35929 = new_n32033 ^ new_n27755;
  assign new_n35930 = new_n35929 ^ new_n30679;
  assign new_n35931 = new_n33903 ^ new_n31196;
  assign new_n35932 = new_n35931 ^ new_n35930;
  assign new_n35933 = new_n32296 ^ new_n27749;
  assign new_n35934 = new_n35933 ^ new_n30968;
  assign new_n35935 = new_n33882 ^ new_n31086;
  assign new_n35936 = new_n35935 ^ new_n35934;
  assign new_n35937 = new_n32341 ^ new_n27730;
  assign new_n35938 = new_n35937 ^ new_n31063;
  assign new_n35939 = new_n35938 ^ new_n33913;
  assign new_n35940 = new_n33868 ^ new_n31153;
  assign new_n35941 = new_n35940 ^ new_n35939;
  assign new_n35942 = new_n33893 ^ new_n31056;
  assign new_n35943 = new_n32380 ^ new_n27738;
  assign new_n35944 = new_n35943 ^ new_n31115;
  assign new_n35945 = new_n35944 ^ new_n33913;
  assign new_n35946 = new_n35945 ^ new_n35942;
  assign new_n35947 = new_n35946 ^ new_n35941;
  assign new_n35948 = new_n35947 ^ new_n35936;
  assign new_n35949 = new_n35948 ^ new_n35932;
  assign new_n35950 = new_n32392 ^ new_n27744;
  assign new_n35951 = new_n35950 ^ new_n31139;
  assign new_n35952 = new_n33913 ^ new_n31107;
  assign new_n35953 = new_n35952 ^ new_n35951;
  assign new_n35954 = new_n33876 ^ new_n31167;
  assign new_n35955 = new_n32404 ^ new_n27724;
  assign new_n35956 = new_n35955 ^ new_n31159;
  assign new_n35957 = new_n35956 ^ new_n33913;
  assign new_n35958 = new_n35957 ^ new_n35954;
  assign new_n35959 = new_n32431 ^ new_n27763;
  assign new_n35960 = new_n35959 ^ new_n31172;
  assign new_n35961 = new_n33897 ^ new_n30508;
  assign new_n35962 = new_n35961 ^ new_n35960;
  assign new_n35963 = new_n35962 ^ new_n35932;
  assign new_n35964 = new_n35963 ^ new_n35953;
  assign new_n35965 = new_n35964 ^ new_n35958;
  assign new_n35966 = new_n35953 & new_n35965;
  assign new_n35967 = new_n35966 ^ new_n35958;
  assign new_n35968 = new_n32455 ^ new_n27717;
  assign new_n35969 = new_n35968 ^ new_n31201;
  assign new_n35970 = new_n33862 ^ new_n31098;
  assign new_n35971 = new_n35970 ^ new_n35969;
  assign new_n35972 = new_n35971 ^ new_n35958;
  assign new_n35973 = new_n35972 ^ new_n35947;
  assign new_n35974 = new_n35958 ^ new_n35946;
  assign new_n35975 = new_n35971 ^ new_n35936;
  assign new_n35976 = new_n35975 ^ new_n35974;
  assign new_n35977 = new_n35973 & new_n35976;
  assign new_n35978 = new_n35977 ^ new_n35932;
  assign new_n35979 = new_n35978 ^ new_n35967;
  assign new_n35980 = ~new_n35946 & ~new_n35964;
  assign new_n35981 = new_n35980 ^ new_n35946;
  assign new_n35982 = new_n35962 ^ new_n35948;
  assign new_n35983 = new_n35971 ^ new_n35946;
  assign new_n35984 = new_n35982 & new_n35983;
  assign new_n35985 = new_n35984 ^ new_n35981;
  assign new_n35986 = new_n35985 ^ new_n35975;
  assign new_n35987 = new_n35949 & new_n35972;
  assign new_n35988 = new_n35962 ^ new_n35958;
  assign new_n35989 = new_n35988 ^ new_n35975;
  assign new_n35990 = new_n35958 ^ new_n35936;
  assign new_n35991 = new_n35989 & new_n35990;
  assign new_n35992 = new_n35991 ^ new_n35987;
  assign new_n35993 = new_n35962 ^ new_n35941;
  assign new_n35994 = new_n35993 ^ new_n35992;
  assign new_n35995 = new_n35994 ^ new_n35986;
  assign new_n35996 = new_n35978 ^ new_n35973;
  assign new_n35997 = new_n35964 ^ new_n35946;
  assign new_n35998 = new_n35997 ^ new_n35975;
  assign new_n35999 = new_n35973 ^ new_n35953;
  assign new_n36000 = new_n35998 & new_n35999;
  assign new_n36001 = new_n36000 ^ new_n35987;
  assign new_n36002 = new_n35991 ^ new_n35936;
  assign new_n36003 = new_n36002 ^ new_n36001;
  assign new_n36004 = new_n36003 ^ new_n35996;
  assign new_n36005 = ~new_n35995 & new_n36004;
  assign new_n36006 = new_n36005 ^ new_n35979;
  assign new_n36007 = new_n35973 ^ new_n35963;
  assign new_n36008 = new_n35975 & new_n36007;
  assign new_n36009 = new_n36008 ^ new_n35987;
  assign new_n36010 = new_n36009 ^ new_n35982;
  assign new_n36011 = new_n36010 ^ new_n36006;
  assign new_n36012 = new_n35971 ^ new_n35964;
  assign new_n36013 = new_n35953 ^ new_n35949;
  assign new_n36014 = new_n36012 & new_n36013;
  assign new_n36015 = new_n36014 ^ new_n35980;
  assign new_n36016 = new_n36008 ^ new_n35991;
  assign new_n36017 = new_n36016 ^ new_n36015;
  assign new_n36018 = ~new_n36017 & new_n36011;
  assign new_n36019 = new_n35971 ^ new_n35962;
  assign new_n36020 = new_n36000 ^ new_n35966;
  assign new_n36021 = new_n36020 ^ new_n36016;
  assign new_n36022 = new_n36021 ^ new_n36019;
  assign new_n36023 = new_n36014 ^ new_n35984;
  assign new_n36024 = new_n36023 ^ new_n35971;
  assign new_n36025 = new_n36024 ^ new_n36010;
  assign new_n36026 = new_n36025 ^ new_n36005;
  assign new_n36027 = new_n36022 & new_n36026;
  assign new_n36028 = new_n36027 ^ new_n36018;
  assign new_n36029 = new_n36024 ^ new_n35979;
  assign new_n36030 = new_n36029 ^ new_n36028;
  assign new_n36031 = new_n35949 & new_n36030;
  assign new_n36032 = new_n36018 ^ new_n36005;
  assign new_n36033 = new_n36025 & new_n36032;
  assign new_n36034 = new_n36033 ^ new_n35995;
  assign new_n36035 = ~new_n36034 & new_n35976;
  assign new_n36036 = new_n36035 ^ new_n36031;
  assign new_n36037 = new_n35962 ^ new_n35946;
  assign new_n36038 = new_n36000 ^ new_n35981;
  assign new_n36039 = new_n36027 ^ new_n35979;
  assign new_n36040 = new_n36039 ^ new_n36010;
  assign new_n36041 = new_n36033 ^ new_n36026;
  assign new_n36042 = new_n36040 & new_n36041;
  assign new_n36043 = new_n36042 ^ new_n36033;
  assign new_n36044 = new_n36043 ^ new_n36038;
  assign new_n36045 = new_n36044 ^ new_n36037;
  assign new_n36046 = new_n36045 ^ new_n35958;
  assign new_n36047 = new_n36027 ^ new_n35984;
  assign new_n36048 = new_n36047 ^ new_n35978;
  assign new_n36049 = new_n36048 ^ new_n36046;
  assign new_n36050 = ~new_n36049 & new_n35989;
  assign new_n36051 = new_n36042 ^ new_n36022;
  assign new_n36052 = new_n35964 & new_n36051;
  assign new_n36053 = new_n36033 ^ new_n36018;
  assign new_n36054 = new_n36053 ^ new_n36017;
  assign new_n36055 = ~new_n36054 & new_n35998;
  assign new_n36056 = ~new_n36049 & new_n35990;
  assign new_n36057 = new_n35972 & new_n36030;
  assign new_n36058 = new_n36057 ^ new_n36056;
  assign new_n36059 = new_n36058 ^ new_n36055;
  assign new_n36060 = new_n36059 ^ new_n36052;
  assign new_n36061 = new_n36042 ^ new_n36027;
  assign new_n36062 = new_n36061 ^ new_n36004;
  assign new_n36063 = new_n35982 & new_n36062;
  assign new_n36064 = new_n36063 ^ new_n36060;
  assign new_n36065 = new_n36064 ^ new_n36050;
  assign new_n36066 = new_n36065 ^ new_n36036;
  assign new_n36067 = new_n32665 ^ new_n32457;
  assign new_n36068 = new_n36067 ^ new_n36066;
  assign new_n36069 = new_n32674 ^ new_n32035;
  assign new_n36070 = new_n36050 ^ new_n36031;
  assign new_n36071 = ~new_n36034 & new_n35973;
  assign new_n36072 = ~new_n36054 & new_n35999;
  assign new_n36073 = new_n36072 ^ new_n36071;
  assign new_n36074 = new_n36073 ^ new_n36035;
  assign new_n36075 = new_n36074 ^ new_n36059;
  assign new_n36076 = new_n36075 ^ new_n36070;
  assign new_n36077 = new_n36076 ^ new_n36069;
  assign new_n36078 = new_n32700 ^ new_n32433;
  assign new_n36079 = new_n36057 ^ new_n36031;
  assign new_n36080 = new_n36018 ^ new_n35971;
  assign new_n36081 = new_n36014 ^ new_n35966;
  assign new_n36082 = new_n36081 ^ new_n36045;
  assign new_n36083 = new_n36082 ^ new_n36080;
  assign new_n36084 = ~new_n36083 & new_n35975;
  assign new_n36085 = new_n35983 & new_n36062;
  assign new_n36086 = new_n36025 ^ new_n36018;
  assign new_n36087 = new_n35953 & new_n36086;
  assign new_n36088 = new_n36087 ^ new_n36071;
  assign new_n36089 = new_n36088 ^ new_n36085;
  assign new_n36090 = ~new_n36083 & new_n36007;
  assign new_n36091 = new_n36012 & new_n36040;
  assign new_n36092 = new_n36091 ^ new_n36090;
  assign new_n36093 = new_n36092 ^ new_n36089;
  assign new_n36094 = new_n36093 ^ new_n36084;
  assign new_n36095 = new_n36094 ^ new_n36079;
  assign new_n36096 = new_n36095 ^ new_n36078;
  assign new_n36097 = new_n36074 ^ new_n36064;
  assign new_n36098 = new_n32721 ^ new_n32406;
  assign new_n36099 = new_n36098 ^ new_n36097;
  assign new_n36100 = new_n36013 & new_n36040;
  assign new_n36101 = new_n36100 ^ new_n36035;
  assign new_n36102 = new_n36087 ^ new_n36072;
  assign new_n36103 = new_n36102 ^ new_n36060;
  assign new_n36104 = new_n36103 ^ new_n36101;
  assign new_n36105 = new_n32733 ^ new_n32343;
  assign new_n36106 = new_n36105 ^ new_n36104;
  assign new_n36107 = new_n35965 & new_n36086;
  assign new_n36108 = new_n36107 ^ new_n36065;
  assign new_n36109 = new_n36108 ^ new_n36093;
  assign new_n36110 = new_n32741 ^ new_n32298;
  assign new_n36111 = new_n36110 ^ new_n36109;
  assign new_n36112 = new_n32750 ^ new_n32382;
  assign new_n36113 = new_n36090 ^ new_n36085;
  assign new_n36114 = new_n35997 & new_n36051;
  assign new_n36115 = new_n36114 ^ new_n36100;
  assign new_n36116 = new_n36115 ^ new_n36058;
  assign new_n36117 = new_n36052 ^ new_n36050;
  assign new_n36118 = new_n36117 ^ new_n36116;
  assign new_n36119 = new_n36118 ^ new_n36113;
  assign new_n36120 = new_n36119 ^ new_n36112;
  assign new_n36121 = new_n32761 ^ new_n32394;
  assign new_n36122 = new_n36089 ^ new_n36063;
  assign new_n36123 = new_n36122 ^ new_n36116;
  assign new_n36124 = new_n36123 ^ new_n36121;
  assign new_n36125 = new_n31538 ^ new_n29963;
  assign new_n36126 = new_n36125 ^ new_n32453;
  assign new_n36127 = new_n36126 ^ new_n32171;
  assign new_n36128 = new_n34127 ^ new_n32421;
  assign new_n36129 = new_n36128 ^ new_n36127;
  assign new_n36130 = new_n31520 ^ new_n29989;
  assign new_n36131 = new_n36130 ^ new_n32319;
  assign new_n36132 = new_n34742 ^ new_n34092;
  assign new_n36133 = new_n36132 ^ new_n36131;
  assign new_n36134 = new_n32413 ^ new_n32242;
  assign new_n36135 = new_n36134 ^ new_n32319;
  assign new_n36136 = new_n31554 ^ new_n29995;
  assign new_n36137 = new_n32448 ^ new_n32346;
  assign new_n36138 = new_n36137 ^ new_n36136;
  assign new_n36139 = new_n36138 ^ new_n34109;
  assign new_n36140 = new_n36139 ^ new_n36135;
  assign new_n36141 = new_n36137 ^ new_n32390;
  assign new_n36142 = new_n36141 ^ new_n34095;
  assign new_n36143 = new_n31533 ^ new_n30003;
  assign new_n36144 = new_n36143 ^ new_n32372;
  assign new_n36145 = new_n36144 ^ new_n32253;
  assign new_n36146 = new_n36145 ^ new_n36142;
  assign new_n36147 = new_n36146 ^ new_n36140;
  assign new_n36148 = new_n36147 ^ new_n36133;
  assign new_n36149 = new_n36148 ^ new_n36129;
  assign new_n36150 = new_n31544 ^ new_n30009;
  assign new_n36151 = new_n36150 ^ new_n32370;
  assign new_n36152 = new_n36137 ^ new_n34106;
  assign new_n36153 = new_n36152 ^ new_n36151;
  assign new_n36154 = new_n31509 ^ new_n30011;
  assign new_n36155 = new_n36154 ^ new_n34117;
  assign new_n36156 = new_n36155 ^ new_n36137;
  assign new_n36157 = new_n32436 ^ new_n32335;
  assign new_n36158 = new_n36157 ^ new_n32413;
  assign new_n36159 = new_n36158 ^ new_n36156;
  assign new_n36160 = new_n31515 ^ new_n30016;
  assign new_n36161 = new_n36160 ^ new_n34759;
  assign new_n36162 = new_n34081 ^ new_n32171;
  assign new_n36163 = new_n36162 ^ new_n36161;
  assign new_n36164 = new_n36163 ^ new_n36129;
  assign new_n36165 = new_n36164 ^ new_n36153;
  assign new_n36166 = new_n36165 ^ new_n36159;
  assign new_n36167 = new_n36153 & new_n36166;
  assign new_n36168 = new_n36167 ^ new_n36159;
  assign new_n36169 = new_n34090 ^ new_n31648;
  assign new_n36170 = new_n31525 ^ new_n30024;
  assign new_n36171 = new_n36170 ^ new_n32346;
  assign new_n36172 = new_n36171 ^ new_n32453;
  assign new_n36173 = new_n36172 ^ new_n36169;
  assign new_n36174 = new_n36173 ^ new_n36159;
  assign new_n36175 = new_n36174 ^ new_n36147;
  assign new_n36176 = new_n36159 ^ new_n36146;
  assign new_n36177 = new_n36173 ^ new_n36133;
  assign new_n36178 = new_n36177 ^ new_n36176;
  assign new_n36179 = ~new_n36175 & new_n36178;
  assign new_n36180 = new_n36179 ^ new_n36129;
  assign new_n36181 = new_n36180 ^ new_n36168;
  assign new_n36182 = ~new_n36146 & ~new_n36165;
  assign new_n36183 = new_n36182 ^ new_n36146;
  assign new_n36184 = new_n36163 ^ new_n36148;
  assign new_n36185 = new_n36173 ^ new_n36146;
  assign new_n36186 = ~new_n36185 & new_n36184;
  assign new_n36187 = new_n36186 ^ new_n36183;
  assign new_n36188 = new_n36187 ^ new_n36177;
  assign new_n36189 = ~new_n36174 & new_n36149;
  assign new_n36190 = new_n36163 ^ new_n36159;
  assign new_n36191 = new_n36190 ^ new_n36177;
  assign new_n36192 = new_n36159 ^ new_n36133;
  assign new_n36193 = ~new_n36191 & ~new_n36192;
  assign new_n36194 = new_n36193 ^ new_n36189;
  assign new_n36195 = new_n36163 ^ new_n36140;
  assign new_n36196 = new_n36195 ^ new_n36194;
  assign new_n36197 = new_n36196 ^ new_n36188;
  assign new_n36198 = new_n36180 ^ new_n36175;
  assign new_n36199 = new_n36165 ^ new_n36146;
  assign new_n36200 = new_n36199 ^ new_n36177;
  assign new_n36201 = new_n36175 ^ new_n36153;
  assign new_n36202 = ~new_n36201 & new_n36200;
  assign new_n36203 = new_n36202 ^ new_n36133;
  assign new_n36204 = new_n36203 ^ new_n36194;
  assign new_n36205 = new_n36204 ^ new_n36198;
  assign new_n36206 = ~new_n36205 & new_n36197;
  assign new_n36207 = new_n36206 ^ new_n36181;
  assign new_n36208 = new_n36175 ^ new_n36164;
  assign new_n36209 = ~new_n36208 & new_n36177;
  assign new_n36210 = new_n36209 ^ new_n36189;
  assign new_n36211 = new_n36210 ^ new_n36184;
  assign new_n36212 = new_n36211 ^ new_n36207;
  assign new_n36213 = new_n36173 ^ new_n36165;
  assign new_n36214 = new_n36153 ^ new_n36149;
  assign new_n36215 = ~new_n36213 & new_n36214;
  assign new_n36216 = new_n36215 ^ new_n36182;
  assign new_n36217 = new_n36209 ^ new_n36193;
  assign new_n36218 = new_n36217 ^ new_n36216;
  assign new_n36219 = ~new_n36212 & ~new_n36218;
  assign new_n36220 = new_n36173 ^ new_n36163;
  assign new_n36221 = new_n36202 ^ new_n36167;
  assign new_n36222 = new_n36221 ^ new_n36217;
  assign new_n36223 = new_n36222 ^ new_n36220;
  assign new_n36224 = new_n36215 ^ new_n36186;
  assign new_n36225 = new_n36224 ^ new_n36173;
  assign new_n36226 = new_n36225 ^ new_n36211;
  assign new_n36227 = new_n36226 ^ new_n36206;
  assign new_n36228 = ~new_n36227 & new_n36223;
  assign new_n36229 = new_n36228 ^ new_n36219;
  assign new_n36230 = new_n36225 ^ new_n36181;
  assign new_n36231 = new_n36230 ^ new_n36229;
  assign new_n36232 = new_n36149 & new_n36231;
  assign new_n36233 = new_n36219 ^ new_n36206;
  assign new_n36234 = ~new_n36226 & new_n36233;
  assign new_n36235 = new_n36234 ^ new_n36197;
  assign new_n36236 = new_n36178 & new_n36235;
  assign new_n36237 = new_n36236 ^ new_n36232;
  assign new_n36238 = new_n36163 ^ new_n36146;
  assign new_n36239 = new_n36202 ^ new_n36183;
  assign new_n36240 = new_n36228 ^ new_n36181;
  assign new_n36241 = new_n36240 ^ new_n36211;
  assign new_n36242 = new_n36234 ^ new_n36227;
  assign new_n36243 = ~new_n36241 & ~new_n36242;
  assign new_n36244 = new_n36243 ^ new_n36234;
  assign new_n36245 = new_n36244 ^ new_n36239;
  assign new_n36246 = new_n36245 ^ new_n36238;
  assign new_n36247 = new_n36246 ^ new_n36159;
  assign new_n36248 = new_n36228 ^ new_n36186;
  assign new_n36249 = new_n36248 ^ new_n36180;
  assign new_n36250 = new_n36249 ^ new_n36247;
  assign new_n36251 = ~new_n36191 & ~new_n36250;
  assign new_n36252 = new_n36243 ^ new_n36223;
  assign new_n36253 = new_n36165 & new_n36252;
  assign new_n36254 = new_n36234 ^ new_n36219;
  assign new_n36255 = new_n36254 ^ new_n36218;
  assign new_n36256 = ~new_n36255 & new_n36200;
  assign new_n36257 = ~new_n36192 & ~new_n36250;
  assign new_n36258 = ~new_n36174 & new_n36231;
  assign new_n36259 = new_n36258 ^ new_n36257;
  assign new_n36260 = new_n36259 ^ new_n36256;
  assign new_n36261 = new_n36260 ^ new_n36253;
  assign new_n36262 = new_n36243 ^ new_n36228;
  assign new_n36263 = new_n36262 ^ new_n36205;
  assign new_n36264 = ~new_n36263 & new_n36184;
  assign new_n36265 = new_n36264 ^ new_n36261;
  assign new_n36266 = new_n36265 ^ new_n36251;
  assign new_n36267 = new_n36266 ^ new_n36237;
  assign new_n36268 = new_n36170 ^ new_n33761;
  assign new_n36269 = new_n36268 ^ new_n36267;
  assign new_n36270 = new_n36125 ^ new_n33770;
  assign new_n36271 = new_n36251 ^ new_n36232;
  assign new_n36272 = ~new_n36175 & new_n36235;
  assign new_n36273 = ~new_n36201 & ~new_n36255;
  assign new_n36274 = new_n36273 ^ new_n36272;
  assign new_n36275 = new_n36274 ^ new_n36236;
  assign new_n36276 = new_n36275 ^ new_n36260;
  assign new_n36277 = new_n36276 ^ new_n36271;
  assign new_n36278 = new_n36277 ^ new_n36270;
  assign new_n36279 = new_n36160 ^ new_n33796;
  assign new_n36280 = new_n36258 ^ new_n36232;
  assign new_n36281 = new_n36219 ^ new_n36173;
  assign new_n36282 = new_n36215 ^ new_n36167;
  assign new_n36283 = new_n36282 ^ new_n36246;
  assign new_n36284 = new_n36283 ^ new_n36281;
  assign new_n36285 = ~new_n36284 & new_n36177;
  assign new_n36286 = ~new_n36185 & ~new_n36263;
  assign new_n36287 = new_n36226 ^ new_n36219;
  assign new_n36288 = ~new_n36287 & new_n36153;
  assign new_n36289 = new_n36288 ^ new_n36272;
  assign new_n36290 = new_n36289 ^ new_n36286;
  assign new_n36291 = ~new_n36208 & ~new_n36284;
  assign new_n36292 = ~new_n36213 & ~new_n36241;
  assign new_n36293 = new_n36292 ^ new_n36291;
  assign new_n36294 = new_n36293 ^ new_n36290;
  assign new_n36295 = new_n36294 ^ new_n36285;
  assign new_n36296 = new_n36295 ^ new_n36280;
  assign new_n36297 = new_n36296 ^ new_n36279;
  assign new_n36298 = new_n36275 ^ new_n36265;
  assign new_n36299 = new_n36154 ^ new_n33817;
  assign new_n36300 = new_n36299 ^ new_n36298;
  assign new_n36301 = ~new_n36241 & new_n36214;
  assign new_n36302 = new_n36301 ^ new_n36236;
  assign new_n36303 = new_n36288 ^ new_n36273;
  assign new_n36304 = new_n36303 ^ new_n36261;
  assign new_n36305 = new_n36304 ^ new_n36302;
  assign new_n36306 = new_n36136 ^ new_n33829;
  assign new_n36307 = new_n36306 ^ new_n36305;
  assign new_n36308 = ~new_n36287 & new_n36166;
  assign new_n36309 = new_n36308 ^ new_n36266;
  assign new_n36310 = new_n36309 ^ new_n36294;
  assign new_n36311 = new_n36130 ^ new_n33837;
  assign new_n36312 = new_n36311 ^ new_n36310;
  assign new_n36313 = new_n36143 ^ new_n33846;
  assign new_n36314 = new_n36291 ^ new_n36286;
  assign new_n36315 = new_n36199 & new_n36252;
  assign new_n36316 = new_n36315 ^ new_n36301;
  assign new_n36317 = new_n36316 ^ new_n36259;
  assign new_n36318 = new_n36253 ^ new_n36251;
  assign new_n36319 = new_n36318 ^ new_n36317;
  assign new_n36320 = new_n36319 ^ new_n36314;
  assign new_n36321 = new_n36320 ^ new_n36313;
  assign new_n36322 = new_n36150 ^ new_n33857;
  assign new_n36323 = new_n36290 ^ new_n36264;
  assign new_n36324 = new_n36323 ^ new_n36317;
  assign new_n36325 = new_n36324 ^ new_n36322;
  assign po0 = new_n30121;
  assign po1 = new_n30137;
  assign po2 = new_n30173;
  assign po3 = new_n30177;
  assign po4 = new_n30189;
  assign po5 = new_n30197;
  assign po6 = new_n30213;
  assign po7 = new_n30219;
  assign po8 = new_n31410;
  assign po9 = new_n31426;
  assign po10 = new_n31462;
  assign po11 = new_n31466;
  assign po12 = new_n31478;
  assign po13 = new_n31486;
  assign po14 = new_n31502;
  assign po15 = new_n31508;
  assign po16 = new_n32667;
  assign po17 = new_n32683;
  assign po18 = new_n32719;
  assign po19 = new_n32723;
  assign po20 = new_n32735;
  assign po21 = new_n32743;
  assign po22 = new_n32759;
  assign po23 = new_n32765;
  assign po24 = new_n33763;
  assign po25 = new_n33779;
  assign po26 = new_n33815;
  assign po27 = ~new_n33819;
  assign po28 = new_n33831;
  assign po29 = ~new_n33839;
  assign po30 = new_n33855;
  assign po31 = new_n33861;
  assign po32 = new_n34015;
  assign po33 = ~new_n34025;
  assign po34 = ~new_n34045;
  assign po35 = new_n34049;
  assign po36 = new_n34057;
  assign po37 = new_n34063;
  assign po38 = ~new_n34073;
  assign po39 = ~new_n34078;
  assign po40 = new_n34227;
  assign po41 = ~new_n34237;
  assign po42 = ~new_n34257;
  assign po43 = new_n34261;
  assign po44 = new_n34269;
  assign po45 = new_n34275;
  assign po46 = ~new_n34285;
  assign po47 = ~new_n34290;
  assign po48 = new_n34434;
  assign po49 = ~new_n34444;
  assign po50 = ~new_n34464;
  assign po51 = new_n34468;
  assign po52 = new_n34476;
  assign po53 = new_n34482;
  assign po54 = ~new_n34492;
  assign po55 = ~new_n34497;
  assign po56 = new_n34662;
  assign po57 = ~new_n34672;
  assign po58 = ~new_n34692;
  assign po59 = ~new_n34696;
  assign po60 = ~new_n34704;
  assign po61 = ~new_n34710;
  assign po62 = new_n34720;
  assign po63 = ~new_n34725;
  assign po64 = new_n34871;
  assign po65 = new_n34880;
  assign po66 = new_n34899;
  assign po67 = new_n34902;
  assign po68 = new_n34909;
  assign po69 = new_n34914;
  assign po70 = new_n34923;
  assign po71 = new_n34927;
  assign po72 = new_n35062;
  assign po73 = new_n35071;
  assign po74 = new_n35090;
  assign po75 = new_n35093;
  assign po76 = new_n35100;
  assign po77 = new_n35105;
  assign po78 = new_n35114;
  assign po79 = new_n35118;
  assign po80 = new_n35266;
  assign po81 = new_n35275;
  assign po82 = new_n35294;
  assign po83 = new_n35297;
  assign po84 = new_n35304;
  assign po85 = new_n35309;
  assign po86 = new_n35318;
  assign po87 = new_n35322;
  assign po88 = ~new_n35469;
  assign po89 = new_n35478;
  assign po90 = new_n35497;
  assign po91 = ~new_n35500;
  assign po92 = ~new_n35507;
  assign po93 = ~new_n35512;
  assign po94 = new_n35521;
  assign po95 = new_n35525;
  assign po96 = new_n35663;
  assign po97 = ~new_n35672;
  assign po98 = ~new_n35691;
  assign po99 = new_n35694;
  assign po100 = new_n35701;
  assign po101 = new_n35706;
  assign po102 = ~new_n35715;
  assign po103 = ~new_n35719;
  assign po104 = new_n35872;
  assign po105 = ~new_n35881;
  assign po106 = ~new_n35900;
  assign po107 = new_n35903;
  assign po108 = new_n35910;
  assign po109 = new_n35915;
  assign po110 = ~new_n35924;
  assign po111 = ~new_n35928;
  assign po112 = new_n36068;
  assign po113 = ~new_n36077;
  assign po114 = ~new_n36096;
  assign po115 = new_n36099;
  assign po116 = new_n36106;
  assign po117 = new_n36111;
  assign po118 = ~new_n36120;
  assign po119 = ~new_n36124;
  assign po120 = ~new_n36269;
  assign po121 = new_n36278;
  assign po122 = ~new_n36297;
  assign po123 = ~new_n36300;
  assign po124 = new_n36307;
  assign po125 = new_n36312;
  assign po126 = new_n36321;
  assign po127 = ~new_n36325;
endmodule


