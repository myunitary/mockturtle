module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 ;
  assign n49 = ~x42 & ~x43 ;
  assign n50 = ~x44 & n49 ;
  assign n51 = ~x39 & ~x40 ;
  assign n52 = ~x41 & n51 ;
  assign n53 = ~n50 & ~n52 ;
  assign n54 = ~x45 & ~x46 ;
  assign n55 = ~x47 & n54 ;
  assign n56 = n50 & n52 ;
  assign n57 = ~n53 & ~n56 ;
  assign n58 = ~n55 & n57 ;
  assign n59 = ~n53 & ~n58 ;
  assign n60 = n55 & ~n57 ;
  assign n61 = ~n58 & ~n60 ;
  assign n62 = ~x27 & ~x28 ;
  assign n63 = ~x29 & n62 ;
  assign n64 = ~n61 & n63 ;
  assign n65 = n61 & ~n63 ;
  assign n66 = ~x36 & ~x37 ;
  assign n67 = ~x38 & n66 ;
  assign n68 = ~x33 & ~x34 ;
  assign n69 = ~x35 & n68 ;
  assign n70 = ~x30 & ~x31 ;
  assign n71 = ~x32 & n70 ;
  assign n72 = ~n69 & ~n71 ;
  assign n73 = n69 & n71 ;
  assign n74 = ~n72 & ~n73 ;
  assign n75 = ~n67 & n74 ;
  assign n76 = n67 & ~n74 ;
  assign n77 = ~n75 & ~n76 ;
  assign n78 = ~n65 & ~n77 ;
  assign n79 = ~n64 & ~n78 ;
  assign n80 = n59 & ~n79 ;
  assign n81 = ~n72 & ~n75 ;
  assign n82 = ~n59 & n79 ;
  assign n83 = ~n80 & ~n82 ;
  assign n84 = n81 & n83 ;
  assign n85 = ~n80 & ~n84 ;
  assign n86 = ~n81 & ~n83 ;
  assign n87 = ~n84 & ~n86 ;
  assign n88 = ~x3 & ~x4 ;
  assign n89 = ~x5 & n88 ;
  assign n90 = ~n64 & ~n65 ;
  assign n91 = ~n77 & n90 ;
  assign n92 = n77 & ~n90 ;
  assign n93 = ~n91 & ~n92 ;
  assign n94 = n89 & n93 ;
  assign n95 = ~n89 & ~n93 ;
  assign n96 = ~x15 & ~x16 ;
  assign n97 = ~x17 & n96 ;
  assign n98 = ~x12 & ~x13 ;
  assign n99 = ~x14 & n98 ;
  assign n100 = ~x9 & ~x10 ;
  assign n101 = ~x11 & n100 ;
  assign n102 = n99 & n101 ;
  assign n103 = ~n99 & ~n101 ;
  assign n104 = ~n102 & ~n103 ;
  assign n105 = ~n97 & n104 ;
  assign n106 = n97 & ~n104 ;
  assign n107 = ~n105 & ~n106 ;
  assign n108 = ~x24 & ~x25 ;
  assign n109 = ~x26 & n108 ;
  assign n110 = ~x21 & ~x22 ;
  assign n111 = ~x23 & n110 ;
  assign n112 = ~x18 & ~x19 ;
  assign n113 = ~x20 & n112 ;
  assign n114 = n111 & n113 ;
  assign n115 = ~n111 & ~n113 ;
  assign n116 = ~n114 & ~n115 ;
  assign n117 = ~n109 & n116 ;
  assign n118 = n109 & ~n116 ;
  assign n119 = ~n117 & ~n118 ;
  assign n120 = ~x6 & ~x7 ;
  assign n121 = ~x8 & n120 ;
  assign n122 = n119 & ~n121 ;
  assign n123 = ~n119 & n121 ;
  assign n124 = ~n122 & ~n123 ;
  assign n125 = n107 & ~n124 ;
  assign n126 = ~n107 & n124 ;
  assign n127 = ~n125 & ~n126 ;
  assign n128 = ~n95 & n127 ;
  assign n129 = ~n94 & ~n128 ;
  assign n130 = n87 & ~n129 ;
  assign n131 = ~n87 & n129 ;
  assign n132 = ~n115 & ~n117 ;
  assign n133 = ~n123 & ~n126 ;
  assign n134 = n132 & ~n133 ;
  assign n135 = ~n132 & n133 ;
  assign n136 = ~n134 & ~n135 ;
  assign n137 = ~n103 & ~n105 ;
  assign n138 = ~n136 & n137 ;
  assign n139 = n136 & ~n137 ;
  assign n140 = ~n138 & ~n139 ;
  assign n141 = ~n131 & ~n140 ;
  assign n142 = ~n130 & ~n141 ;
  assign n143 = n85 & n142 ;
  assign n144 = ~n134 & ~n137 ;
  assign n145 = ~n135 & ~n144 ;
  assign n146 = ~n85 & ~n142 ;
  assign n147 = ~n143 & ~n146 ;
  assign n148 = ~n145 & n147 ;
  assign n149 = ~n143 & ~n148 ;
  assign n150 = n145 & ~n147 ;
  assign n151 = ~n148 & ~n150 ;
  assign n152 = ~x0 & ~x1 ;
  assign n153 = ~x2 & n152 ;
  assign n154 = ~n94 & ~n95 ;
  assign n155 = n127 & n154 ;
  assign n156 = ~n127 & ~n154 ;
  assign n157 = ~n155 & ~n156 ;
  assign n158 = n153 & n157 ;
  assign n159 = ~n130 & ~n131 ;
  assign n160 = ~n140 & n159 ;
  assign n161 = n140 & ~n159 ;
  assign n162 = ~n160 & ~n161 ;
  assign n163 = n158 & n162 ;
  assign n164 = ~n151 & n163 ;
  assign n165 = n149 & n164 ;
  assign n166 = x3 & ~x4 ;
  assign n167 = ~x5 & n166 ;
  assign n168 = x27 & ~x28 ;
  assign n169 = ~x29 & n168 ;
  assign n170 = x45 & ~x46 ;
  assign n171 = ~x47 & n170 ;
  assign n172 = x42 & ~x43 ;
  assign n173 = ~x44 & n172 ;
  assign n174 = x39 & ~x40 ;
  assign n175 = ~x41 & n174 ;
  assign n176 = ~n173 & ~n175 ;
  assign n177 = n173 & n175 ;
  assign n178 = ~n176 & ~n177 ;
  assign n179 = n171 & ~n178 ;
  assign n180 = ~n171 & n178 ;
  assign n181 = ~n179 & ~n180 ;
  assign n182 = n169 & ~n181 ;
  assign n183 = ~n169 & n181 ;
  assign n184 = ~n182 & ~n183 ;
  assign n185 = x36 & ~x37 ;
  assign n186 = ~x38 & n185 ;
  assign n187 = x33 & ~x34 ;
  assign n188 = ~x35 & n187 ;
  assign n189 = x30 & ~x31 ;
  assign n190 = ~x32 & n189 ;
  assign n191 = n188 & n190 ;
  assign n192 = ~n188 & ~n190 ;
  assign n193 = ~n191 & ~n192 ;
  assign n194 = n186 & ~n193 ;
  assign n195 = ~n186 & n193 ;
  assign n196 = ~n194 & ~n195 ;
  assign n197 = n184 & ~n196 ;
  assign n198 = ~n184 & n196 ;
  assign n199 = ~n197 & ~n198 ;
  assign n200 = n167 & n199 ;
  assign n201 = x6 & ~x7 ;
  assign n202 = ~x8 & n201 ;
  assign n203 = x24 & ~x25 ;
  assign n204 = ~x26 & n203 ;
  assign n205 = x21 & ~x22 ;
  assign n206 = ~x23 & n205 ;
  assign n207 = x18 & ~x19 ;
  assign n208 = ~x20 & n207 ;
  assign n209 = n206 & n208 ;
  assign n210 = ~n206 & ~n208 ;
  assign n211 = ~n209 & ~n210 ;
  assign n212 = n204 & ~n211 ;
  assign n213 = ~n204 & n211 ;
  assign n214 = ~n212 & ~n213 ;
  assign n215 = ~n202 & n214 ;
  assign n216 = n202 & ~n214 ;
  assign n217 = ~n215 & ~n216 ;
  assign n218 = x15 & ~x16 ;
  assign n219 = ~x17 & n218 ;
  assign n220 = x12 & ~x13 ;
  assign n221 = ~x14 & n220 ;
  assign n222 = x9 & ~x10 ;
  assign n223 = ~x11 & n222 ;
  assign n224 = n221 & n223 ;
  assign n225 = ~n221 & ~n223 ;
  assign n226 = ~n224 & ~n225 ;
  assign n227 = n219 & ~n226 ;
  assign n228 = ~n219 & n226 ;
  assign n229 = ~n227 & ~n228 ;
  assign n230 = n217 & ~n229 ;
  assign n231 = ~n217 & n229 ;
  assign n232 = ~n230 & ~n231 ;
  assign n233 = ~n167 & ~n199 ;
  assign n234 = ~n200 & ~n233 ;
  assign n235 = n232 & n234 ;
  assign n236 = ~n200 & ~n235 ;
  assign n237 = ~n186 & ~n191 ;
  assign n238 = ~n192 & ~n237 ;
  assign n239 = ~n171 & ~n177 ;
  assign n240 = ~n176 & ~n239 ;
  assign n241 = ~n182 & ~n197 ;
  assign n242 = ~n240 & n241 ;
  assign n243 = n240 & ~n241 ;
  assign n244 = ~n242 & ~n243 ;
  assign n245 = n238 & n244 ;
  assign n246 = ~n238 & ~n244 ;
  assign n247 = ~n245 & ~n246 ;
  assign n248 = n236 & ~n247 ;
  assign n249 = ~n236 & n247 ;
  assign n250 = ~n219 & ~n224 ;
  assign n251 = ~n225 & ~n250 ;
  assign n252 = ~n204 & ~n209 ;
  assign n253 = ~n210 & ~n252 ;
  assign n254 = ~n216 & ~n230 ;
  assign n255 = n253 & ~n254 ;
  assign n256 = ~n253 & n254 ;
  assign n257 = ~n255 & ~n256 ;
  assign n258 = n251 & n257 ;
  assign n259 = ~n251 & ~n257 ;
  assign n260 = ~n258 & ~n259 ;
  assign n261 = ~n249 & ~n260 ;
  assign n262 = ~n248 & ~n261 ;
  assign n263 = ~n243 & ~n245 ;
  assign n264 = ~n262 & n263 ;
  assign n265 = n262 & ~n263 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = ~n255 & ~n258 ;
  assign n268 = n266 & n267 ;
  assign n269 = ~n264 & ~n268 ;
  assign n270 = ~n266 & ~n267 ;
  assign n271 = ~n268 & ~n270 ;
  assign n272 = x0 & ~x1 ;
  assign n273 = ~x2 & n272 ;
  assign n274 = ~n232 & ~n234 ;
  assign n275 = ~n235 & ~n274 ;
  assign n276 = n273 & n275 ;
  assign n277 = ~n248 & ~n249 ;
  assign n278 = ~n260 & n277 ;
  assign n279 = n260 & ~n277 ;
  assign n280 = ~n278 & ~n279 ;
  assign n281 = n276 & ~n280 ;
  assign n282 = ~n271 & n281 ;
  assign n283 = n269 & n282 ;
  assign n284 = ~n165 & n283 ;
  assign n285 = ~n149 & ~n164 ;
  assign n286 = ~n165 & ~n285 ;
  assign n287 = ~n269 & ~n282 ;
  assign n288 = ~n283 & ~n287 ;
  assign n289 = ~n286 & n288 ;
  assign n290 = n151 & ~n163 ;
  assign n291 = ~n164 & ~n290 ;
  assign n292 = ~n273 & ~n275 ;
  assign n293 = ~n276 & ~n292 ;
  assign n294 = ~n153 & ~n157 ;
  assign n295 = ~n158 & ~n294 ;
  assign n296 = ~n293 & n295 ;
  assign n297 = n162 & n296 ;
  assign n298 = ~n158 & ~n162 ;
  assign n299 = ~n163 & ~n298 ;
  assign n300 = ~n296 & ~n299 ;
  assign n301 = ~n276 & n280 ;
  assign n302 = ~n281 & ~n301 ;
  assign n303 = ~n300 & ~n302 ;
  assign n304 = ~n297 & ~n303 ;
  assign n305 = ~n291 & n304 ;
  assign n306 = n271 & ~n281 ;
  assign n307 = ~n282 & ~n306 ;
  assign n308 = n291 & ~n304 ;
  assign n309 = n307 & ~n308 ;
  assign n310 = ~n305 & ~n309 ;
  assign n311 = ~n289 & n310 ;
  assign n312 = n165 & ~n283 ;
  assign n313 = n286 & ~n288 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = ~n311 & n314 ;
  assign n316 = ~n284 & ~n315 ;
  assign n317 = ~x42 & x43 ;
  assign n318 = x44 & n317 ;
  assign n319 = ~x39 & x40 ;
  assign n320 = x41 & n319 ;
  assign n321 = ~n318 & ~n320 ;
  assign n322 = ~x45 & x46 ;
  assign n323 = x47 & n322 ;
  assign n324 = n318 & n320 ;
  assign n325 = ~n323 & ~n324 ;
  assign n326 = ~n321 & ~n325 ;
  assign n327 = ~x27 & x28 ;
  assign n328 = x29 & n327 ;
  assign n329 = ~n321 & ~n324 ;
  assign n330 = n323 & ~n329 ;
  assign n331 = ~n323 & n329 ;
  assign n332 = ~n330 & ~n331 ;
  assign n333 = n328 & ~n332 ;
  assign n334 = ~n328 & n332 ;
  assign n335 = ~n333 & ~n334 ;
  assign n336 = ~x36 & x37 ;
  assign n337 = x38 & n336 ;
  assign n338 = ~x33 & x34 ;
  assign n339 = x35 & n338 ;
  assign n340 = ~x30 & x31 ;
  assign n341 = x32 & n340 ;
  assign n342 = ~n339 & ~n341 ;
  assign n343 = n339 & n341 ;
  assign n344 = ~n342 & ~n343 ;
  assign n345 = n337 & ~n344 ;
  assign n346 = ~n337 & n344 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = n335 & ~n347 ;
  assign n349 = ~n333 & ~n348 ;
  assign n350 = n326 & ~n349 ;
  assign n351 = ~n337 & ~n343 ;
  assign n352 = ~n342 & ~n351 ;
  assign n353 = ~n326 & n349 ;
  assign n354 = ~n350 & ~n353 ;
  assign n355 = n352 & n354 ;
  assign n356 = ~n350 & ~n355 ;
  assign n357 = ~n352 & ~n354 ;
  assign n358 = ~n355 & ~n357 ;
  assign n359 = ~x3 & x4 ;
  assign n360 = x5 & n359 ;
  assign n361 = ~n335 & n347 ;
  assign n362 = ~n348 & ~n361 ;
  assign n363 = n360 & n362 ;
  assign n364 = ~x6 & x7 ;
  assign n365 = x8 & n364 ;
  assign n366 = ~x24 & x25 ;
  assign n367 = x26 & n366 ;
  assign n368 = ~x21 & x22 ;
  assign n369 = x23 & n368 ;
  assign n370 = ~x18 & x19 ;
  assign n371 = x20 & n370 ;
  assign n372 = n369 & n371 ;
  assign n373 = ~n369 & ~n371 ;
  assign n374 = ~n372 & ~n373 ;
  assign n375 = n367 & ~n374 ;
  assign n376 = ~n367 & n374 ;
  assign n377 = ~n375 & ~n376 ;
  assign n378 = ~n365 & n377 ;
  assign n379 = n365 & ~n377 ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = ~x15 & x16 ;
  assign n382 = x17 & n381 ;
  assign n383 = ~x12 & x13 ;
  assign n384 = x14 & n383 ;
  assign n385 = ~x9 & x10 ;
  assign n386 = x11 & n385 ;
  assign n387 = n384 & n386 ;
  assign n388 = ~n384 & ~n386 ;
  assign n389 = ~n387 & ~n388 ;
  assign n390 = n382 & ~n389 ;
  assign n391 = ~n382 & n389 ;
  assign n392 = ~n390 & ~n391 ;
  assign n393 = n380 & ~n392 ;
  assign n394 = ~n380 & n392 ;
  assign n395 = ~n393 & ~n394 ;
  assign n396 = ~n360 & ~n362 ;
  assign n397 = ~n363 & ~n396 ;
  assign n398 = n395 & n397 ;
  assign n399 = ~n363 & ~n398 ;
  assign n400 = n358 & ~n399 ;
  assign n401 = ~n382 & ~n387 ;
  assign n402 = ~n388 & ~n401 ;
  assign n403 = ~n367 & ~n372 ;
  assign n404 = ~n373 & ~n403 ;
  assign n405 = ~n379 & ~n393 ;
  assign n406 = n404 & ~n405 ;
  assign n407 = ~n404 & n405 ;
  assign n408 = ~n406 & ~n407 ;
  assign n409 = n402 & n408 ;
  assign n410 = ~n402 & ~n408 ;
  assign n411 = ~n409 & ~n410 ;
  assign n412 = ~n358 & n399 ;
  assign n413 = ~n400 & ~n412 ;
  assign n414 = n411 & n413 ;
  assign n415 = ~n400 & ~n414 ;
  assign n416 = n356 & n415 ;
  assign n417 = ~n356 & ~n415 ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = ~n406 & ~n409 ;
  assign n420 = n418 & n419 ;
  assign n421 = ~n416 & ~n420 ;
  assign n422 = ~n418 & ~n419 ;
  assign n423 = ~n420 & ~n422 ;
  assign n424 = ~x0 & x1 ;
  assign n425 = x2 & n424 ;
  assign n426 = ~n395 & ~n397 ;
  assign n427 = ~n398 & ~n426 ;
  assign n428 = n425 & n427 ;
  assign n429 = ~n411 & ~n413 ;
  assign n430 = ~n414 & ~n429 ;
  assign n431 = n428 & n430 ;
  assign n432 = ~n423 & n431 ;
  assign n433 = n421 & n432 ;
  assign n434 = x0 & x1 ;
  assign n435 = x2 & n434 ;
  assign n436 = x6 & x7 ;
  assign n437 = x8 & n436 ;
  assign n438 = x24 & x25 ;
  assign n439 = x26 & n438 ;
  assign n440 = x21 & x22 ;
  assign n441 = x23 & n440 ;
  assign n442 = x18 & x19 ;
  assign n443 = x20 & n442 ;
  assign n444 = n441 & n443 ;
  assign n445 = ~n441 & ~n443 ;
  assign n446 = ~n444 & ~n445 ;
  assign n447 = n439 & ~n446 ;
  assign n448 = ~n439 & n446 ;
  assign n449 = ~n447 & ~n448 ;
  assign n450 = ~n437 & n449 ;
  assign n451 = n437 & ~n449 ;
  assign n452 = ~n450 & ~n451 ;
  assign n453 = x15 & x16 ;
  assign n454 = x17 & n453 ;
  assign n455 = x12 & x13 ;
  assign n456 = x14 & n455 ;
  assign n457 = x9 & x10 ;
  assign n458 = x11 & n457 ;
  assign n459 = n456 & n458 ;
  assign n460 = ~n456 & ~n458 ;
  assign n461 = ~n459 & ~n460 ;
  assign n462 = n454 & ~n461 ;
  assign n463 = ~n454 & n461 ;
  assign n464 = ~n462 & ~n463 ;
  assign n465 = n452 & ~n464 ;
  assign n466 = ~n452 & n464 ;
  assign n467 = ~n465 & ~n466 ;
  assign n468 = x3 & x4 ;
  assign n469 = x5 & n468 ;
  assign n470 = x27 & x28 ;
  assign n471 = x29 & n470 ;
  assign n472 = x45 & x46 ;
  assign n473 = x47 & n472 ;
  assign n474 = x42 & x43 ;
  assign n475 = x44 & n474 ;
  assign n476 = x39 & x40 ;
  assign n477 = x41 & n476 ;
  assign n478 = ~n475 & ~n477 ;
  assign n479 = n475 & n477 ;
  assign n480 = ~n478 & ~n479 ;
  assign n481 = n473 & ~n480 ;
  assign n482 = ~n473 & n480 ;
  assign n483 = ~n481 & ~n482 ;
  assign n484 = n471 & ~n483 ;
  assign n485 = ~n471 & n483 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = x36 & x37 ;
  assign n488 = x38 & n487 ;
  assign n489 = x33 & x34 ;
  assign n490 = x35 & n489 ;
  assign n491 = x30 & x31 ;
  assign n492 = x32 & n491 ;
  assign n493 = ~n490 & ~n492 ;
  assign n494 = n490 & n492 ;
  assign n495 = ~n493 & ~n494 ;
  assign n496 = n488 & ~n495 ;
  assign n497 = ~n488 & n495 ;
  assign n498 = ~n496 & ~n497 ;
  assign n499 = n486 & ~n498 ;
  assign n500 = ~n486 & n498 ;
  assign n501 = ~n499 & ~n500 ;
  assign n502 = n469 & n501 ;
  assign n503 = ~n469 & ~n501 ;
  assign n504 = ~n502 & ~n503 ;
  assign n505 = n467 & n504 ;
  assign n506 = ~n467 & ~n504 ;
  assign n507 = ~n505 & ~n506 ;
  assign n508 = n435 & n507 ;
  assign n509 = ~n454 & ~n459 ;
  assign n510 = ~n460 & ~n509 ;
  assign n511 = ~n439 & ~n444 ;
  assign n512 = ~n445 & ~n511 ;
  assign n513 = ~n451 & ~n465 ;
  assign n514 = n512 & ~n513 ;
  assign n515 = ~n512 & n513 ;
  assign n516 = ~n514 & ~n515 ;
  assign n517 = n510 & n516 ;
  assign n518 = ~n510 & ~n516 ;
  assign n519 = ~n517 & ~n518 ;
  assign n520 = ~n488 & ~n494 ;
  assign n521 = ~n493 & ~n520 ;
  assign n522 = ~n473 & ~n479 ;
  assign n523 = ~n478 & ~n522 ;
  assign n524 = ~n484 & ~n499 ;
  assign n525 = n523 & ~n524 ;
  assign n526 = ~n523 & n524 ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = n521 & n527 ;
  assign n529 = ~n521 & ~n527 ;
  assign n530 = ~n528 & ~n529 ;
  assign n531 = ~n502 & ~n505 ;
  assign n532 = n530 & ~n531 ;
  assign n533 = ~n530 & n531 ;
  assign n534 = ~n532 & ~n533 ;
  assign n535 = n519 & n534 ;
  assign n536 = ~n519 & ~n534 ;
  assign n537 = ~n535 & ~n536 ;
  assign n538 = n508 & n537 ;
  assign n539 = ~n525 & ~n528 ;
  assign n540 = ~n532 & ~n535 ;
  assign n541 = n539 & n540 ;
  assign n542 = ~n539 & ~n540 ;
  assign n543 = ~n541 & ~n542 ;
  assign n544 = ~n514 & ~n517 ;
  assign n545 = n543 & n544 ;
  assign n546 = ~n543 & ~n544 ;
  assign n547 = ~n545 & ~n546 ;
  assign n548 = n538 & ~n547 ;
  assign n549 = ~n541 & ~n545 ;
  assign n550 = n548 & n549 ;
  assign n551 = ~n433 & ~n550 ;
  assign n552 = x2 & n152 ;
  assign n553 = x8 & n120 ;
  assign n554 = x26 & n108 ;
  assign n555 = x23 & n110 ;
  assign n556 = x20 & n112 ;
  assign n557 = ~n555 & ~n556 ;
  assign n558 = n555 & n556 ;
  assign n559 = ~n557 & ~n558 ;
  assign n560 = n554 & ~n559 ;
  assign n561 = ~n554 & n559 ;
  assign n562 = ~n560 & ~n561 ;
  assign n563 = n553 & ~n562 ;
  assign n564 = ~n553 & n562 ;
  assign n565 = ~n563 & ~n564 ;
  assign n566 = x17 & n96 ;
  assign n567 = x14 & n98 ;
  assign n568 = x11 & n100 ;
  assign n569 = n567 & n568 ;
  assign n570 = ~n567 & ~n568 ;
  assign n571 = ~n569 & ~n570 ;
  assign n572 = n566 & ~n571 ;
  assign n573 = ~n566 & n571 ;
  assign n574 = ~n572 & ~n573 ;
  assign n575 = n565 & ~n574 ;
  assign n576 = ~n565 & n574 ;
  assign n577 = ~n575 & ~n576 ;
  assign n578 = x5 & n88 ;
  assign n579 = x29 & n62 ;
  assign n580 = x47 & n54 ;
  assign n581 = x44 & n49 ;
  assign n582 = x41 & n51 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = n581 & n582 ;
  assign n585 = ~n583 & ~n584 ;
  assign n586 = n580 & ~n585 ;
  assign n587 = ~n580 & n585 ;
  assign n588 = ~n586 & ~n587 ;
  assign n589 = n579 & ~n588 ;
  assign n590 = ~n579 & n588 ;
  assign n591 = ~n589 & ~n590 ;
  assign n592 = x38 & n66 ;
  assign n593 = x35 & n68 ;
  assign n594 = x32 & n70 ;
  assign n595 = ~n593 & ~n594 ;
  assign n596 = n593 & n594 ;
  assign n597 = ~n595 & ~n596 ;
  assign n598 = n592 & ~n597 ;
  assign n599 = ~n592 & n597 ;
  assign n600 = ~n598 & ~n599 ;
  assign n601 = n591 & ~n600 ;
  assign n602 = ~n591 & n600 ;
  assign n603 = ~n601 & ~n602 ;
  assign n604 = n578 & n603 ;
  assign n605 = ~n578 & ~n603 ;
  assign n606 = ~n604 & ~n605 ;
  assign n607 = n577 & n606 ;
  assign n608 = ~n577 & ~n606 ;
  assign n609 = ~n607 & ~n608 ;
  assign n610 = n552 & n609 ;
  assign n611 = ~n566 & ~n569 ;
  assign n612 = ~n570 & ~n611 ;
  assign n613 = ~n554 & ~n558 ;
  assign n614 = ~n557 & ~n613 ;
  assign n615 = ~n563 & ~n575 ;
  assign n616 = ~n614 & n615 ;
  assign n617 = n614 & ~n615 ;
  assign n618 = ~n616 & ~n617 ;
  assign n619 = n612 & n618 ;
  assign n620 = ~n612 & ~n618 ;
  assign n621 = ~n619 & ~n620 ;
  assign n622 = ~n592 & ~n596 ;
  assign n623 = ~n595 & ~n622 ;
  assign n624 = ~n580 & ~n584 ;
  assign n625 = ~n583 & ~n624 ;
  assign n626 = ~n589 & ~n601 ;
  assign n627 = n625 & ~n626 ;
  assign n628 = ~n625 & n626 ;
  assign n629 = ~n627 & ~n628 ;
  assign n630 = n623 & n629 ;
  assign n631 = ~n623 & ~n629 ;
  assign n632 = ~n630 & ~n631 ;
  assign n633 = ~n604 & ~n607 ;
  assign n634 = n632 & ~n633 ;
  assign n635 = ~n632 & n633 ;
  assign n636 = ~n634 & ~n635 ;
  assign n637 = n621 & n636 ;
  assign n638 = ~n621 & ~n636 ;
  assign n639 = ~n637 & ~n638 ;
  assign n640 = n610 & n639 ;
  assign n641 = ~n627 & ~n630 ;
  assign n642 = ~n634 & ~n637 ;
  assign n643 = n641 & n642 ;
  assign n644 = ~n641 & ~n642 ;
  assign n645 = ~n643 & ~n644 ;
  assign n646 = ~n617 & ~n619 ;
  assign n647 = n645 & n646 ;
  assign n648 = ~n645 & ~n646 ;
  assign n649 = ~n647 & ~n648 ;
  assign n650 = n640 & ~n649 ;
  assign n651 = ~n643 & ~n647 ;
  assign n652 = n650 & n651 ;
  assign n653 = x44 & n172 ;
  assign n654 = x41 & n174 ;
  assign n655 = ~n653 & ~n654 ;
  assign n656 = x47 & n170 ;
  assign n657 = n653 & n654 ;
  assign n658 = ~n656 & ~n657 ;
  assign n659 = ~n655 & ~n658 ;
  assign n660 = x29 & n168 ;
  assign n661 = ~n655 & ~n657 ;
  assign n662 = n656 & ~n661 ;
  assign n663 = ~n656 & n661 ;
  assign n664 = ~n662 & ~n663 ;
  assign n665 = n660 & ~n664 ;
  assign n666 = ~n660 & n664 ;
  assign n667 = ~n665 & ~n666 ;
  assign n668 = x38 & n185 ;
  assign n669 = x35 & n187 ;
  assign n670 = x32 & n189 ;
  assign n671 = n669 & n670 ;
  assign n672 = ~n669 & ~n670 ;
  assign n673 = ~n671 & ~n672 ;
  assign n674 = n668 & ~n673 ;
  assign n675 = ~n668 & n673 ;
  assign n676 = ~n674 & ~n675 ;
  assign n677 = n667 & ~n676 ;
  assign n678 = ~n665 & ~n677 ;
  assign n679 = n659 & ~n678 ;
  assign n680 = ~n668 & ~n671 ;
  assign n681 = ~n672 & ~n680 ;
  assign n682 = ~n659 & n678 ;
  assign n683 = ~n679 & ~n682 ;
  assign n684 = n681 & n683 ;
  assign n685 = ~n679 & ~n684 ;
  assign n686 = x5 & n166 ;
  assign n687 = ~n667 & n676 ;
  assign n688 = ~n677 & ~n687 ;
  assign n689 = n686 & n688 ;
  assign n690 = x8 & n201 ;
  assign n691 = x26 & n203 ;
  assign n692 = x23 & n205 ;
  assign n693 = x20 & n207 ;
  assign n694 = n692 & n693 ;
  assign n695 = ~n692 & ~n693 ;
  assign n696 = ~n694 & ~n695 ;
  assign n697 = n691 & ~n696 ;
  assign n698 = ~n691 & n696 ;
  assign n699 = ~n697 & ~n698 ;
  assign n700 = ~n690 & n699 ;
  assign n701 = n690 & ~n699 ;
  assign n702 = ~n700 & ~n701 ;
  assign n703 = x17 & n218 ;
  assign n704 = x14 & n220 ;
  assign n705 = x11 & n222 ;
  assign n706 = n704 & n705 ;
  assign n707 = ~n704 & ~n705 ;
  assign n708 = ~n706 & ~n707 ;
  assign n709 = n703 & ~n708 ;
  assign n710 = ~n703 & n708 ;
  assign n711 = ~n709 & ~n710 ;
  assign n712 = n702 & ~n711 ;
  assign n713 = ~n702 & n711 ;
  assign n714 = ~n712 & ~n713 ;
  assign n715 = ~n686 & ~n688 ;
  assign n716 = ~n689 & ~n715 ;
  assign n717 = n714 & n716 ;
  assign n718 = ~n689 & ~n717 ;
  assign n719 = ~n681 & ~n683 ;
  assign n720 = ~n684 & ~n719 ;
  assign n721 = n718 & ~n720 ;
  assign n722 = ~n703 & ~n706 ;
  assign n723 = ~n707 & ~n722 ;
  assign n724 = ~n691 & ~n694 ;
  assign n725 = ~n695 & ~n724 ;
  assign n726 = ~n701 & ~n712 ;
  assign n727 = n725 & ~n726 ;
  assign n728 = ~n725 & n726 ;
  assign n729 = ~n727 & ~n728 ;
  assign n730 = n723 & n729 ;
  assign n731 = ~n723 & ~n729 ;
  assign n732 = ~n730 & ~n731 ;
  assign n733 = ~n718 & n720 ;
  assign n734 = ~n721 & ~n733 ;
  assign n735 = ~n732 & n734 ;
  assign n736 = ~n721 & ~n735 ;
  assign n737 = n685 & ~n736 ;
  assign n738 = ~n685 & n736 ;
  assign n739 = ~n737 & ~n738 ;
  assign n740 = ~n727 & ~n730 ;
  assign n741 = n739 & n740 ;
  assign n742 = ~n737 & ~n741 ;
  assign n743 = ~n739 & ~n740 ;
  assign n744 = ~n741 & ~n743 ;
  assign n745 = x2 & n272 ;
  assign n746 = ~n714 & ~n716 ;
  assign n747 = ~n717 & ~n746 ;
  assign n748 = n745 & n747 ;
  assign n749 = n732 & ~n734 ;
  assign n750 = ~n735 & ~n749 ;
  assign n751 = n748 & ~n750 ;
  assign n752 = ~n744 & n751 ;
  assign n753 = n742 & n752 ;
  assign n754 = ~n652 & ~n753 ;
  assign n755 = n551 & ~n754 ;
  assign n756 = ~n435 & ~n507 ;
  assign n757 = ~n508 & ~n756 ;
  assign n758 = ~n433 & n550 ;
  assign n759 = ~n538 & n547 ;
  assign n760 = ~n548 & ~n759 ;
  assign n761 = n423 & ~n431 ;
  assign n762 = ~n432 & ~n761 ;
  assign n763 = ~n760 & n762 ;
  assign n764 = ~n508 & ~n537 ;
  assign n765 = ~n538 & ~n764 ;
  assign n766 = ~n428 & ~n430 ;
  assign n767 = ~n431 & ~n766 ;
  assign n768 = ~n765 & n767 ;
  assign n769 = n765 & ~n767 ;
  assign n770 = ~n425 & ~n427 ;
  assign n771 = ~n428 & ~n770 ;
  assign n772 = ~n757 & n771 ;
  assign n773 = ~n769 & n772 ;
  assign n774 = ~n768 & ~n773 ;
  assign n775 = ~n763 & n774 ;
  assign n776 = ~n421 & ~n432 ;
  assign n777 = ~n433 & ~n776 ;
  assign n778 = ~n548 & ~n549 ;
  assign n779 = ~n550 & ~n778 ;
  assign n780 = ~n777 & n779 ;
  assign n781 = n760 & ~n762 ;
  assign n782 = ~n780 & ~n781 ;
  assign n783 = ~n775 & n782 ;
  assign n784 = n433 & ~n550 ;
  assign n785 = n777 & ~n779 ;
  assign n786 = ~n784 & ~n785 ;
  assign n787 = ~n783 & n786 ;
  assign n788 = ~n758 & ~n787 ;
  assign n789 = ~n757 & ~n788 ;
  assign n790 = ~n771 & n788 ;
  assign n791 = ~n789 & ~n790 ;
  assign n792 = ~n745 & ~n747 ;
  assign n793 = ~n748 & ~n792 ;
  assign n794 = ~n652 & n753 ;
  assign n795 = ~n650 & ~n651 ;
  assign n796 = ~n652 & ~n795 ;
  assign n797 = ~n742 & ~n752 ;
  assign n798 = ~n753 & ~n797 ;
  assign n799 = ~n796 & n798 ;
  assign n800 = n744 & ~n751 ;
  assign n801 = ~n752 & ~n800 ;
  assign n802 = ~n640 & n649 ;
  assign n803 = ~n650 & ~n802 ;
  assign n804 = ~n610 & ~n639 ;
  assign n805 = ~n640 & ~n804 ;
  assign n806 = ~n748 & n750 ;
  assign n807 = ~n751 & ~n806 ;
  assign n808 = n805 & ~n807 ;
  assign n809 = ~n639 & n807 ;
  assign n810 = ~n552 & ~n609 ;
  assign n811 = ~n610 & ~n810 ;
  assign n812 = ~n793 & n811 ;
  assign n813 = ~n809 & n812 ;
  assign n814 = ~n808 & ~n813 ;
  assign n815 = n803 & ~n814 ;
  assign n816 = n801 & ~n815 ;
  assign n817 = ~n803 & n814 ;
  assign n818 = ~n816 & ~n817 ;
  assign n819 = ~n799 & n818 ;
  assign n820 = n652 & ~n753 ;
  assign n821 = n796 & ~n798 ;
  assign n822 = ~n820 & ~n821 ;
  assign n823 = ~n819 & n822 ;
  assign n824 = ~n794 & ~n823 ;
  assign n825 = ~n793 & ~n824 ;
  assign n826 = ~n811 & n824 ;
  assign n827 = ~n825 & ~n826 ;
  assign n828 = ~n791 & n827 ;
  assign n829 = n807 & ~n824 ;
  assign n830 = n805 & n824 ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = n767 & n788 ;
  assign n833 = n765 & ~n788 ;
  assign n834 = ~n832 & ~n833 ;
  assign n835 = ~n831 & n834 ;
  assign n836 = ~n828 & ~n835 ;
  assign n837 = n831 & ~n834 ;
  assign n838 = ~n801 & ~n824 ;
  assign n839 = ~n803 & n824 ;
  assign n840 = ~n838 & ~n839 ;
  assign n841 = n762 & n788 ;
  assign n842 = n760 & ~n788 ;
  assign n843 = ~n841 & ~n842 ;
  assign n844 = ~n840 & ~n843 ;
  assign n845 = ~n837 & ~n844 ;
  assign n846 = ~n836 & n845 ;
  assign n847 = n840 & n843 ;
  assign n848 = n776 & n778 ;
  assign n849 = n551 & ~n848 ;
  assign n850 = n795 & n797 ;
  assign n851 = n754 & ~n850 ;
  assign n852 = ~n849 & n851 ;
  assign n853 = ~n847 & ~n852 ;
  assign n854 = ~n846 & n853 ;
  assign n855 = ~n551 & n754 ;
  assign n856 = n849 & ~n851 ;
  assign n857 = ~n855 & ~n856 ;
  assign n858 = ~n854 & n857 ;
  assign n859 = ~n755 & ~n858 ;
  assign n860 = ~n302 & ~n316 ;
  assign n861 = ~n299 & n316 ;
  assign n862 = ~n860 & ~n861 ;
  assign n863 = ~x2 & n424 ;
  assign n864 = ~x8 & n364 ;
  assign n865 = ~x26 & n366 ;
  assign n866 = ~x23 & n368 ;
  assign n867 = ~x20 & n370 ;
  assign n868 = n866 & n867 ;
  assign n869 = ~n866 & ~n867 ;
  assign n870 = ~n868 & ~n869 ;
  assign n871 = n865 & ~n870 ;
  assign n872 = ~n865 & n870 ;
  assign n873 = ~n871 & ~n872 ;
  assign n874 = ~n864 & n873 ;
  assign n875 = n864 & ~n873 ;
  assign n876 = ~n874 & ~n875 ;
  assign n877 = ~x17 & n381 ;
  assign n878 = ~x14 & n383 ;
  assign n879 = ~x11 & n385 ;
  assign n880 = n878 & n879 ;
  assign n881 = ~n878 & ~n879 ;
  assign n882 = ~n880 & ~n881 ;
  assign n883 = n877 & ~n882 ;
  assign n884 = ~n877 & n882 ;
  assign n885 = ~n883 & ~n884 ;
  assign n886 = n876 & ~n885 ;
  assign n887 = ~n876 & n885 ;
  assign n888 = ~n886 & ~n887 ;
  assign n889 = ~x5 & n359 ;
  assign n890 = ~x29 & n327 ;
  assign n891 = ~x47 & n322 ;
  assign n892 = ~x44 & n317 ;
  assign n893 = ~x41 & n319 ;
  assign n894 = ~n892 & ~n893 ;
  assign n895 = n892 & n893 ;
  assign n896 = ~n894 & ~n895 ;
  assign n897 = n891 & ~n896 ;
  assign n898 = ~n891 & n896 ;
  assign n899 = ~n897 & ~n898 ;
  assign n900 = ~n890 & n899 ;
  assign n901 = n890 & ~n899 ;
  assign n902 = ~n900 & ~n901 ;
  assign n903 = ~x38 & n336 ;
  assign n904 = ~x35 & n338 ;
  assign n905 = ~x32 & n340 ;
  assign n906 = ~n904 & ~n905 ;
  assign n907 = n904 & n905 ;
  assign n908 = ~n906 & ~n907 ;
  assign n909 = n903 & ~n908 ;
  assign n910 = ~n903 & n908 ;
  assign n911 = ~n909 & ~n910 ;
  assign n912 = n902 & n911 ;
  assign n913 = ~n902 & ~n911 ;
  assign n914 = ~n912 & ~n913 ;
  assign n915 = ~n889 & n914 ;
  assign n916 = n889 & ~n914 ;
  assign n917 = ~n915 & ~n916 ;
  assign n918 = n888 & ~n917 ;
  assign n919 = ~n888 & n917 ;
  assign n920 = ~n918 & ~n919 ;
  assign n921 = n863 & ~n920 ;
  assign n922 = ~n877 & ~n880 ;
  assign n923 = ~n881 & ~n922 ;
  assign n924 = ~n865 & ~n868 ;
  assign n925 = ~n869 & ~n924 ;
  assign n926 = ~n875 & ~n886 ;
  assign n927 = n925 & ~n926 ;
  assign n928 = ~n925 & n926 ;
  assign n929 = ~n927 & ~n928 ;
  assign n930 = n923 & n929 ;
  assign n931 = ~n923 & ~n929 ;
  assign n932 = ~n930 & ~n931 ;
  assign n933 = ~n903 & ~n907 ;
  assign n934 = ~n906 & ~n933 ;
  assign n935 = ~n891 & ~n895 ;
  assign n936 = ~n894 & ~n935 ;
  assign n937 = ~n900 & ~n911 ;
  assign n938 = ~n901 & ~n937 ;
  assign n939 = n936 & ~n938 ;
  assign n940 = ~n936 & n938 ;
  assign n941 = ~n939 & ~n940 ;
  assign n942 = n934 & n941 ;
  assign n943 = ~n934 & ~n941 ;
  assign n944 = ~n942 & ~n943 ;
  assign n945 = n888 & ~n915 ;
  assign n946 = ~n916 & ~n945 ;
  assign n947 = ~n944 & n946 ;
  assign n948 = n944 & ~n946 ;
  assign n949 = ~n947 & ~n948 ;
  assign n950 = n932 & n949 ;
  assign n951 = ~n932 & ~n949 ;
  assign n952 = ~n950 & ~n951 ;
  assign n953 = n921 & n952 ;
  assign n954 = ~n939 & ~n942 ;
  assign n955 = n932 & ~n947 ;
  assign n956 = ~n948 & ~n955 ;
  assign n957 = n954 & n956 ;
  assign n958 = ~n954 & ~n956 ;
  assign n959 = ~n957 & ~n958 ;
  assign n960 = ~n927 & ~n930 ;
  assign n961 = n959 & n960 ;
  assign n962 = ~n959 & ~n960 ;
  assign n963 = ~n961 & ~n962 ;
  assign n964 = n953 & ~n963 ;
  assign n965 = ~n957 & ~n961 ;
  assign n966 = n964 & n965 ;
  assign n967 = ~x5 & n468 ;
  assign n968 = ~x29 & n470 ;
  assign n969 = ~x47 & n472 ;
  assign n970 = ~x44 & n474 ;
  assign n971 = ~x41 & n476 ;
  assign n972 = ~n970 & ~n971 ;
  assign n973 = n970 & n971 ;
  assign n974 = ~n972 & ~n973 ;
  assign n975 = n969 & ~n974 ;
  assign n976 = ~n969 & n974 ;
  assign n977 = ~n975 & ~n976 ;
  assign n978 = n968 & ~n977 ;
  assign n979 = ~n968 & n977 ;
  assign n980 = ~n978 & ~n979 ;
  assign n981 = ~x38 & n487 ;
  assign n982 = ~x35 & n489 ;
  assign n983 = ~x32 & n491 ;
  assign n984 = n982 & n983 ;
  assign n985 = ~n982 & ~n983 ;
  assign n986 = ~n984 & ~n985 ;
  assign n987 = n981 & ~n986 ;
  assign n988 = ~n981 & n986 ;
  assign n989 = ~n987 & ~n988 ;
  assign n990 = n980 & ~n989 ;
  assign n991 = ~n980 & n989 ;
  assign n992 = ~n990 & ~n991 ;
  assign n993 = n967 & n992 ;
  assign n994 = ~x8 & n436 ;
  assign n995 = ~x26 & n438 ;
  assign n996 = ~x23 & n440 ;
  assign n997 = ~x20 & n442 ;
  assign n998 = n996 & n997 ;
  assign n999 = ~n996 & ~n997 ;
  assign n1000 = ~n998 & ~n999 ;
  assign n1001 = n995 & ~n1000 ;
  assign n1002 = ~n995 & n1000 ;
  assign n1003 = ~n1001 & ~n1002 ;
  assign n1004 = ~n994 & n1003 ;
  assign n1005 = n994 & ~n1003 ;
  assign n1006 = ~n1004 & ~n1005 ;
  assign n1007 = ~x17 & n453 ;
  assign n1008 = ~x14 & n455 ;
  assign n1009 = ~x11 & n457 ;
  assign n1010 = n1008 & n1009 ;
  assign n1011 = ~n1008 & ~n1009 ;
  assign n1012 = ~n1010 & ~n1011 ;
  assign n1013 = n1007 & ~n1012 ;
  assign n1014 = ~n1007 & n1012 ;
  assign n1015 = ~n1013 & ~n1014 ;
  assign n1016 = n1006 & ~n1015 ;
  assign n1017 = ~n1006 & n1015 ;
  assign n1018 = ~n1016 & ~n1017 ;
  assign n1019 = ~n967 & ~n992 ;
  assign n1020 = ~n993 & ~n1019 ;
  assign n1021 = n1018 & n1020 ;
  assign n1022 = ~n993 & ~n1021 ;
  assign n1023 = ~n981 & ~n984 ;
  assign n1024 = ~n985 & ~n1023 ;
  assign n1025 = ~n969 & ~n973 ;
  assign n1026 = ~n972 & ~n1025 ;
  assign n1027 = ~n978 & ~n990 ;
  assign n1028 = ~n1026 & n1027 ;
  assign n1029 = n1026 & ~n1027 ;
  assign n1030 = ~n1028 & ~n1029 ;
  assign n1031 = n1024 & n1030 ;
  assign n1032 = ~n1024 & ~n1030 ;
  assign n1033 = ~n1031 & ~n1032 ;
  assign n1034 = n1022 & ~n1033 ;
  assign n1035 = ~n1022 & n1033 ;
  assign n1036 = ~n1007 & ~n1010 ;
  assign n1037 = ~n1011 & ~n1036 ;
  assign n1038 = ~n995 & ~n998 ;
  assign n1039 = ~n999 & ~n1038 ;
  assign n1040 = ~n1005 & ~n1016 ;
  assign n1041 = n1039 & ~n1040 ;
  assign n1042 = ~n1039 & n1040 ;
  assign n1043 = ~n1041 & ~n1042 ;
  assign n1044 = n1037 & n1043 ;
  assign n1045 = ~n1037 & ~n1043 ;
  assign n1046 = ~n1044 & ~n1045 ;
  assign n1047 = ~n1035 & ~n1046 ;
  assign n1048 = ~n1034 & ~n1047 ;
  assign n1049 = ~n1029 & ~n1031 ;
  assign n1050 = ~n1048 & n1049 ;
  assign n1051 = n1048 & ~n1049 ;
  assign n1052 = ~n1050 & ~n1051 ;
  assign n1053 = ~n1041 & ~n1044 ;
  assign n1054 = n1052 & n1053 ;
  assign n1055 = ~n1050 & ~n1054 ;
  assign n1056 = ~n1052 & ~n1053 ;
  assign n1057 = ~n1054 & ~n1056 ;
  assign n1058 = ~x2 & n434 ;
  assign n1059 = ~n1018 & ~n1020 ;
  assign n1060 = ~n1021 & ~n1059 ;
  assign n1061 = n1058 & n1060 ;
  assign n1062 = ~n1034 & ~n1035 ;
  assign n1063 = ~n1046 & n1062 ;
  assign n1064 = n1046 & ~n1062 ;
  assign n1065 = ~n1063 & ~n1064 ;
  assign n1066 = n1061 & ~n1065 ;
  assign n1067 = ~n1057 & n1066 ;
  assign n1068 = n1055 & n1067 ;
  assign n1069 = ~n966 & ~n1068 ;
  assign n1070 = ~n165 & ~n283 ;
  assign n1071 = n1069 & ~n1070 ;
  assign n1072 = ~n1055 & ~n1067 ;
  assign n1073 = ~n964 & ~n965 ;
  assign n1074 = n1072 & n1073 ;
  assign n1075 = n1069 & ~n1074 ;
  assign n1076 = n285 & n287 ;
  assign n1077 = n1070 & ~n1076 ;
  assign n1078 = ~n1075 & n1077 ;
  assign n1079 = n1057 & ~n1066 ;
  assign n1080 = ~n1067 & ~n1079 ;
  assign n1081 = ~n966 & n1068 ;
  assign n1082 = ~n1068 & ~n1072 ;
  assign n1083 = ~n966 & ~n1073 ;
  assign n1084 = n1082 & ~n1083 ;
  assign n1085 = ~n953 & n963 ;
  assign n1086 = ~n964 & ~n1085 ;
  assign n1087 = ~n1058 & ~n1060 ;
  assign n1088 = ~n1061 & ~n1087 ;
  assign n1089 = ~n863 & n920 ;
  assign n1090 = ~n921 & ~n1089 ;
  assign n1091 = ~n1088 & n1090 ;
  assign n1092 = n952 & n1091 ;
  assign n1093 = ~n921 & ~n952 ;
  assign n1094 = ~n953 & ~n1093 ;
  assign n1095 = ~n1091 & ~n1094 ;
  assign n1096 = ~n1061 & n1065 ;
  assign n1097 = ~n1066 & ~n1096 ;
  assign n1098 = ~n1095 & ~n1097 ;
  assign n1099 = ~n1092 & ~n1098 ;
  assign n1100 = n1086 & ~n1099 ;
  assign n1101 = ~n1086 & n1099 ;
  assign n1102 = ~n1080 & ~n1101 ;
  assign n1103 = ~n1100 & ~n1102 ;
  assign n1104 = ~n1084 & ~n1103 ;
  assign n1105 = n966 & ~n1068 ;
  assign n1106 = ~n1082 & n1083 ;
  assign n1107 = ~n1105 & ~n1106 ;
  assign n1108 = ~n1104 & n1107 ;
  assign n1109 = ~n1081 & ~n1108 ;
  assign n1110 = ~n1080 & ~n1109 ;
  assign n1111 = ~n1086 & n1109 ;
  assign n1112 = ~n1110 & ~n1111 ;
  assign n1113 = ~n307 & ~n316 ;
  assign n1114 = ~n291 & n316 ;
  assign n1115 = ~n1113 & ~n1114 ;
  assign n1116 = n1112 & ~n1115 ;
  assign n1117 = ~n1088 & ~n1109 ;
  assign n1118 = ~n1090 & n1109 ;
  assign n1119 = ~n1117 & ~n1118 ;
  assign n1120 = ~n293 & ~n316 ;
  assign n1121 = ~n295 & n316 ;
  assign n1122 = ~n1120 & ~n1121 ;
  assign n1123 = ~n1119 & n1122 ;
  assign n1124 = ~n1097 & ~n1109 ;
  assign n1125 = ~n1094 & n1109 ;
  assign n1126 = ~n1124 & ~n1125 ;
  assign n1127 = ~n1123 & n1126 ;
  assign n1128 = n862 & ~n1127 ;
  assign n1129 = ~n1112 & n1115 ;
  assign n1130 = n1123 & ~n1126 ;
  assign n1131 = ~n1129 & ~n1130 ;
  assign n1132 = ~n1128 & n1131 ;
  assign n1133 = ~n1116 & ~n1132 ;
  assign n1134 = ~n1078 & ~n1133 ;
  assign n1135 = ~n1069 & n1070 ;
  assign n1136 = n1075 & ~n1077 ;
  assign n1137 = ~n1135 & ~n1136 ;
  assign n1138 = ~n1134 & n1137 ;
  assign n1139 = ~n1071 & ~n1138 ;
  assign n1140 = ~n862 & ~n1139 ;
  assign n1141 = ~n1126 & n1139 ;
  assign n1142 = ~n1140 & ~n1141 ;
  assign n1143 = ~n834 & n859 ;
  assign n1144 = ~n831 & ~n859 ;
  assign n1145 = ~n1143 & ~n1144 ;
  assign n1146 = ~n1142 & ~n1145 ;
  assign n1147 = ~n827 & ~n859 ;
  assign n1148 = ~n791 & n859 ;
  assign n1149 = ~n1147 & ~n1148 ;
  assign n1150 = n1119 & n1139 ;
  assign n1151 = n1122 & ~n1139 ;
  assign n1152 = ~n1150 & ~n1151 ;
  assign n1153 = ~n1149 & ~n1152 ;
  assign n1154 = ~n1146 & n1153 ;
  assign n1155 = ~n1115 & ~n1139 ;
  assign n1156 = ~n1112 & n1139 ;
  assign n1157 = ~n1155 & ~n1156 ;
  assign n1158 = ~n843 & n859 ;
  assign n1159 = n840 & ~n859 ;
  assign n1160 = ~n1158 & ~n1159 ;
  assign n1161 = n1157 & n1160 ;
  assign n1162 = n1142 & n1145 ;
  assign n1163 = ~n1161 & ~n1162 ;
  assign n1164 = ~n1154 & n1163 ;
  assign n1165 = n849 & n859 ;
  assign n1166 = n851 & n858 ;
  assign n1167 = ~n1165 & ~n1166 ;
  assign n1168 = n1075 & n1139 ;
  assign n1169 = n1077 & n1138 ;
  assign n1170 = ~n1168 & ~n1169 ;
  assign n1171 = ~n1167 & n1170 ;
  assign n1172 = ~n1157 & ~n1160 ;
  assign n1173 = ~n1171 & ~n1172 ;
  assign n1174 = ~n1164 & n1173 ;
  assign n1175 = n1167 & ~n1170 ;
  assign n1176 = n1069 & n1070 ;
  assign n1177 = n551 & n754 ;
  assign n1178 = ~n1176 & n1177 ;
  assign n1179 = ~n1175 & ~n1178 ;
  assign n1180 = ~n1174 & n1179 ;
  assign n1181 = n1176 & ~n1177 ;
  assign n1182 = ~n1180 & ~n1181 ;
  assign n1183 = n859 & ~n1182 ;
  assign n1184 = n1139 & n1182 ;
  assign n1185 = ~n1183 & ~n1184 ;
  assign n1186 = n316 & n1185 ;
  assign n1187 = n1109 & n1139 ;
  assign n1188 = n1182 & ~n1187 ;
  assign n1189 = ~n1186 & n1188 ;
  assign n1190 = n824 & n1185 ;
  assign n1191 = n788 & n859 ;
  assign n1192 = ~n1182 & ~n1191 ;
  assign n1193 = ~n1190 & n1192 ;
  assign n1194 = ~n1189 & ~n1193 ;
  assign y0 = ~n1194 ;
  assign y1 = ~n1185 ;
  assign y2 = ~n1182 ;
endmodule
