module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 ;
  assign n513 = ~x287 & ~x319 ;
  assign n514 = ~x351 & ~x383 ;
  assign n515 = n513 & n514 ;
  assign n516 = ~x415 & ~x447 ;
  assign n517 = ~x479 & ~x511 ;
  assign n518 = n516 & n517 ;
  assign n519 = n515 & n518 ;
  assign n520 = ~x31 & ~x63 ;
  assign n521 = ~x95 & ~x127 ;
  assign n522 = n520 & n521 ;
  assign n523 = ~x159 & ~x191 ;
  assign n524 = ~x223 & ~x255 ;
  assign n525 = n523 & n524 ;
  assign n526 = n522 & n525 ;
  assign n527 = n519 & ~n526 ;
  assign n528 = ~x31 & x63 ;
  assign n529 = x31 & ~x63 ;
  assign n530 = ~x30 & x62 ;
  assign n531 = x30 & ~x62 ;
  assign n532 = ~x29 & x61 ;
  assign n533 = x29 & ~x61 ;
  assign n534 = ~x28 & x60 ;
  assign n535 = x28 & ~x60 ;
  assign n536 = ~x27 & x59 ;
  assign n537 = x27 & ~x59 ;
  assign n538 = ~x26 & x58 ;
  assign n539 = x26 & ~x58 ;
  assign n540 = ~x25 & x57 ;
  assign n541 = x25 & ~x57 ;
  assign n542 = ~x24 & x56 ;
  assign n543 = x24 & ~x56 ;
  assign n544 = ~x23 & x55 ;
  assign n545 = x23 & ~x55 ;
  assign n546 = ~x22 & x54 ;
  assign n547 = x22 & ~x54 ;
  assign n548 = ~x21 & x53 ;
  assign n549 = x21 & ~x53 ;
  assign n550 = ~x20 & x52 ;
  assign n551 = x20 & ~x52 ;
  assign n552 = ~x19 & x51 ;
  assign n553 = x19 & ~x51 ;
  assign n554 = ~x18 & x50 ;
  assign n555 = x18 & ~x50 ;
  assign n556 = ~x17 & x49 ;
  assign n557 = x17 & ~x49 ;
  assign n558 = ~x16 & x48 ;
  assign n559 = x16 & ~x48 ;
  assign n560 = ~x15 & x47 ;
  assign n561 = x15 & ~x47 ;
  assign n562 = ~x14 & x46 ;
  assign n563 = x14 & ~x46 ;
  assign n564 = ~x13 & x45 ;
  assign n565 = x13 & ~x45 ;
  assign n566 = ~x12 & x44 ;
  assign n567 = x12 & ~x44 ;
  assign n568 = ~x11 & x43 ;
  assign n569 = x11 & ~x43 ;
  assign n570 = ~x10 & x42 ;
  assign n571 = x10 & ~x42 ;
  assign n572 = ~x9 & x41 ;
  assign n573 = x9 & ~x41 ;
  assign n574 = ~x8 & x40 ;
  assign n575 = x8 & ~x40 ;
  assign n576 = ~x7 & x39 ;
  assign n577 = x7 & ~x39 ;
  assign n578 = ~x6 & x38 ;
  assign n579 = x6 & ~x38 ;
  assign n580 = ~x5 & x37 ;
  assign n581 = x5 & ~x37 ;
  assign n582 = ~x4 & x36 ;
  assign n583 = x4 & ~x36 ;
  assign n584 = ~x3 & x35 ;
  assign n585 = x3 & ~x35 ;
  assign n586 = ~x2 & x34 ;
  assign n587 = x2 & ~x34 ;
  assign n588 = ~x1 & x33 ;
  assign n589 = x1 & ~x33 ;
  assign n590 = x0 & ~x32 ;
  assign n591 = ~n589 & ~n590 ;
  assign n592 = ~n588 & ~n591 ;
  assign n593 = ~n587 & ~n592 ;
  assign n594 = ~n586 & ~n593 ;
  assign n595 = ~n585 & ~n594 ;
  assign n596 = ~n584 & ~n595 ;
  assign n597 = ~n583 & ~n596 ;
  assign n598 = ~n582 & ~n597 ;
  assign n599 = ~n581 & ~n598 ;
  assign n600 = ~n580 & ~n599 ;
  assign n601 = ~n579 & ~n600 ;
  assign n602 = ~n578 & ~n601 ;
  assign n603 = ~n577 & ~n602 ;
  assign n604 = ~n576 & ~n603 ;
  assign n605 = ~n575 & ~n604 ;
  assign n606 = ~n574 & ~n605 ;
  assign n607 = ~n573 & ~n606 ;
  assign n608 = ~n572 & ~n607 ;
  assign n609 = ~n571 & ~n608 ;
  assign n610 = ~n570 & ~n609 ;
  assign n611 = ~n569 & ~n610 ;
  assign n612 = ~n568 & ~n611 ;
  assign n613 = ~n567 & ~n612 ;
  assign n614 = ~n566 & ~n613 ;
  assign n615 = ~n565 & ~n614 ;
  assign n616 = ~n564 & ~n615 ;
  assign n617 = ~n563 & ~n616 ;
  assign n618 = ~n562 & ~n617 ;
  assign n619 = ~n561 & ~n618 ;
  assign n620 = ~n560 & ~n619 ;
  assign n621 = ~n559 & ~n620 ;
  assign n622 = ~n558 & ~n621 ;
  assign n623 = ~n557 & ~n622 ;
  assign n624 = ~n556 & ~n623 ;
  assign n625 = ~n555 & ~n624 ;
  assign n626 = ~n554 & ~n625 ;
  assign n627 = ~n553 & ~n626 ;
  assign n628 = ~n552 & ~n627 ;
  assign n629 = ~n551 & ~n628 ;
  assign n630 = ~n550 & ~n629 ;
  assign n631 = ~n549 & ~n630 ;
  assign n632 = ~n548 & ~n631 ;
  assign n633 = ~n547 & ~n632 ;
  assign n634 = ~n546 & ~n633 ;
  assign n635 = ~n545 & ~n634 ;
  assign n636 = ~n544 & ~n635 ;
  assign n637 = ~n543 & ~n636 ;
  assign n638 = ~n542 & ~n637 ;
  assign n639 = ~n541 & ~n638 ;
  assign n640 = ~n540 & ~n639 ;
  assign n641 = ~n539 & ~n640 ;
  assign n642 = ~n538 & ~n641 ;
  assign n643 = ~n537 & ~n642 ;
  assign n644 = ~n536 & ~n643 ;
  assign n645 = ~n535 & ~n644 ;
  assign n646 = ~n534 & ~n645 ;
  assign n647 = ~n533 & ~n646 ;
  assign n648 = ~n532 & ~n647 ;
  assign n649 = ~n531 & ~n648 ;
  assign n650 = ~n530 & ~n649 ;
  assign n651 = ~n529 & ~n650 ;
  assign n652 = ~n528 & ~n651 ;
  assign n653 = x59 & ~n652 ;
  assign n654 = x27 & n652 ;
  assign n655 = ~n653 & ~n654 ;
  assign n656 = n520 & ~n521 ;
  assign n657 = ~n520 & n521 ;
  assign n658 = x33 & ~n652 ;
  assign n659 = x1 & n652 ;
  assign n660 = ~n658 & ~n659 ;
  assign n661 = ~x95 & x127 ;
  assign n662 = x95 & ~x127 ;
  assign n663 = ~x94 & x126 ;
  assign n664 = x94 & ~x126 ;
  assign n665 = ~x93 & x125 ;
  assign n666 = x93 & ~x125 ;
  assign n667 = ~x92 & x124 ;
  assign n668 = x92 & ~x124 ;
  assign n669 = ~x91 & x123 ;
  assign n670 = x91 & ~x123 ;
  assign n671 = ~x90 & x122 ;
  assign n672 = x90 & ~x122 ;
  assign n673 = ~x89 & x121 ;
  assign n674 = x89 & ~x121 ;
  assign n675 = ~x88 & x120 ;
  assign n676 = x88 & ~x120 ;
  assign n677 = ~x87 & x119 ;
  assign n678 = x87 & ~x119 ;
  assign n679 = ~x86 & x118 ;
  assign n680 = x86 & ~x118 ;
  assign n681 = ~x85 & x117 ;
  assign n682 = x85 & ~x117 ;
  assign n683 = ~x84 & x116 ;
  assign n684 = x84 & ~x116 ;
  assign n685 = ~x83 & x115 ;
  assign n686 = x83 & ~x115 ;
  assign n687 = ~x82 & x114 ;
  assign n688 = x82 & ~x114 ;
  assign n689 = ~x81 & x113 ;
  assign n690 = x81 & ~x113 ;
  assign n691 = ~x80 & x112 ;
  assign n692 = x80 & ~x112 ;
  assign n693 = ~x79 & x111 ;
  assign n694 = x79 & ~x111 ;
  assign n695 = ~x78 & x110 ;
  assign n696 = x78 & ~x110 ;
  assign n697 = ~x77 & x109 ;
  assign n698 = x77 & ~x109 ;
  assign n699 = ~x76 & x108 ;
  assign n700 = x76 & ~x108 ;
  assign n701 = ~x75 & x107 ;
  assign n702 = x75 & ~x107 ;
  assign n703 = ~x74 & x106 ;
  assign n704 = x74 & ~x106 ;
  assign n705 = ~x73 & x105 ;
  assign n706 = x73 & ~x105 ;
  assign n707 = ~x72 & x104 ;
  assign n708 = x72 & ~x104 ;
  assign n709 = ~x71 & x103 ;
  assign n710 = x71 & ~x103 ;
  assign n711 = ~x70 & x102 ;
  assign n712 = x70 & ~x102 ;
  assign n713 = ~x69 & x101 ;
  assign n714 = x69 & ~x101 ;
  assign n715 = ~x68 & x100 ;
  assign n716 = x68 & ~x100 ;
  assign n717 = ~x67 & x99 ;
  assign n718 = x67 & ~x99 ;
  assign n719 = ~x66 & x98 ;
  assign n720 = x66 & ~x98 ;
  assign n721 = ~x65 & x97 ;
  assign n722 = x65 & ~x97 ;
  assign n723 = x64 & ~x96 ;
  assign n724 = ~n722 & ~n723 ;
  assign n725 = ~n721 & ~n724 ;
  assign n726 = ~n720 & ~n725 ;
  assign n727 = ~n719 & ~n726 ;
  assign n728 = ~n718 & ~n727 ;
  assign n729 = ~n717 & ~n728 ;
  assign n730 = ~n716 & ~n729 ;
  assign n731 = ~n715 & ~n730 ;
  assign n732 = ~n714 & ~n731 ;
  assign n733 = ~n713 & ~n732 ;
  assign n734 = ~n712 & ~n733 ;
  assign n735 = ~n711 & ~n734 ;
  assign n736 = ~n710 & ~n735 ;
  assign n737 = ~n709 & ~n736 ;
  assign n738 = ~n708 & ~n737 ;
  assign n739 = ~n707 & ~n738 ;
  assign n740 = ~n706 & ~n739 ;
  assign n741 = ~n705 & ~n740 ;
  assign n742 = ~n704 & ~n741 ;
  assign n743 = ~n703 & ~n742 ;
  assign n744 = ~n702 & ~n743 ;
  assign n745 = ~n701 & ~n744 ;
  assign n746 = ~n700 & ~n745 ;
  assign n747 = ~n699 & ~n746 ;
  assign n748 = ~n698 & ~n747 ;
  assign n749 = ~n697 & ~n748 ;
  assign n750 = ~n696 & ~n749 ;
  assign n751 = ~n695 & ~n750 ;
  assign n752 = ~n694 & ~n751 ;
  assign n753 = ~n693 & ~n752 ;
  assign n754 = ~n692 & ~n753 ;
  assign n755 = ~n691 & ~n754 ;
  assign n756 = ~n690 & ~n755 ;
  assign n757 = ~n689 & ~n756 ;
  assign n758 = ~n688 & ~n757 ;
  assign n759 = ~n687 & ~n758 ;
  assign n760 = ~n686 & ~n759 ;
  assign n761 = ~n685 & ~n760 ;
  assign n762 = ~n684 & ~n761 ;
  assign n763 = ~n683 & ~n762 ;
  assign n764 = ~n682 & ~n763 ;
  assign n765 = ~n681 & ~n764 ;
  assign n766 = ~n680 & ~n765 ;
  assign n767 = ~n679 & ~n766 ;
  assign n768 = ~n678 & ~n767 ;
  assign n769 = ~n677 & ~n768 ;
  assign n770 = ~n676 & ~n769 ;
  assign n771 = ~n675 & ~n770 ;
  assign n772 = ~n674 & ~n771 ;
  assign n773 = ~n673 & ~n772 ;
  assign n774 = ~n672 & ~n773 ;
  assign n775 = ~n671 & ~n774 ;
  assign n776 = ~n670 & ~n775 ;
  assign n777 = ~n669 & ~n776 ;
  assign n778 = ~n668 & ~n777 ;
  assign n779 = ~n667 & ~n778 ;
  assign n780 = ~n666 & ~n779 ;
  assign n781 = ~n665 & ~n780 ;
  assign n782 = ~n664 & ~n781 ;
  assign n783 = ~n663 & ~n782 ;
  assign n784 = ~n662 & ~n783 ;
  assign n785 = ~n661 & ~n784 ;
  assign n786 = x97 & ~n785 ;
  assign n787 = x65 & n785 ;
  assign n788 = ~n786 & ~n787 ;
  assign n789 = n660 & ~n788 ;
  assign n790 = x32 & ~n652 ;
  assign n791 = x0 & n652 ;
  assign n792 = ~n790 & ~n791 ;
  assign n793 = x96 & ~n785 ;
  assign n794 = x64 & n785 ;
  assign n795 = ~n793 & ~n794 ;
  assign n796 = ~n792 & n795 ;
  assign n797 = ~n789 & n796 ;
  assign n798 = x98 & ~n785 ;
  assign n799 = x66 & n785 ;
  assign n800 = ~n798 & ~n799 ;
  assign n801 = x34 & ~n652 ;
  assign n802 = x2 & n652 ;
  assign n803 = ~n801 & ~n802 ;
  assign n804 = n800 & ~n803 ;
  assign n805 = ~n660 & n788 ;
  assign n806 = ~n804 & ~n805 ;
  assign n807 = ~n797 & n806 ;
  assign n808 = x35 & ~n652 ;
  assign n809 = x3 & n652 ;
  assign n810 = ~n808 & ~n809 ;
  assign n811 = x99 & ~n785 ;
  assign n812 = x67 & n785 ;
  assign n813 = ~n811 & ~n812 ;
  assign n814 = n810 & ~n813 ;
  assign n815 = ~n800 & n803 ;
  assign n816 = ~n814 & ~n815 ;
  assign n817 = ~n807 & n816 ;
  assign n818 = ~n810 & n813 ;
  assign n819 = x36 & ~n652 ;
  assign n820 = x4 & n652 ;
  assign n821 = ~n819 & ~n820 ;
  assign n822 = x100 & ~n785 ;
  assign n823 = x68 & n785 ;
  assign n824 = ~n822 & ~n823 ;
  assign n825 = ~n821 & n824 ;
  assign n826 = ~n818 & ~n825 ;
  assign n827 = ~n817 & n826 ;
  assign n828 = n821 & ~n824 ;
  assign n829 = x101 & ~n785 ;
  assign n830 = x69 & n785 ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = x37 & ~n652 ;
  assign n833 = x5 & n652 ;
  assign n834 = ~n832 & ~n833 ;
  assign n835 = ~n831 & n834 ;
  assign n836 = ~n828 & ~n835 ;
  assign n837 = ~n827 & n836 ;
  assign n838 = n831 & ~n834 ;
  assign n839 = x102 & ~n785 ;
  assign n840 = x70 & n785 ;
  assign n841 = ~n839 & ~n840 ;
  assign n842 = x38 & ~n652 ;
  assign n843 = x6 & n652 ;
  assign n844 = ~n842 & ~n843 ;
  assign n845 = n841 & ~n844 ;
  assign n846 = ~n838 & ~n845 ;
  assign n847 = ~n837 & n846 ;
  assign n848 = ~n841 & n844 ;
  assign n849 = x39 & ~n652 ;
  assign n850 = x7 & n652 ;
  assign n851 = ~n849 & ~n850 ;
  assign n852 = x103 & ~n785 ;
  assign n853 = x71 & n785 ;
  assign n854 = ~n852 & ~n853 ;
  assign n855 = n851 & ~n854 ;
  assign n856 = ~n848 & ~n855 ;
  assign n857 = ~n847 & n856 ;
  assign n858 = ~n851 & n854 ;
  assign n859 = x104 & ~n785 ;
  assign n860 = x72 & n785 ;
  assign n861 = ~n859 & ~n860 ;
  assign n862 = x40 & ~n652 ;
  assign n863 = x8 & n652 ;
  assign n864 = ~n862 & ~n863 ;
  assign n865 = n861 & ~n864 ;
  assign n866 = ~n858 & ~n865 ;
  assign n867 = ~n857 & n866 ;
  assign n868 = ~n861 & n864 ;
  assign n869 = x105 & ~n785 ;
  assign n870 = x73 & n785 ;
  assign n871 = ~n869 & ~n870 ;
  assign n872 = x41 & ~n652 ;
  assign n873 = x9 & n652 ;
  assign n874 = ~n872 & ~n873 ;
  assign n875 = ~n871 & n874 ;
  assign n876 = ~n868 & ~n875 ;
  assign n877 = ~n867 & n876 ;
  assign n878 = n871 & ~n874 ;
  assign n879 = x42 & ~n652 ;
  assign n880 = x10 & n652 ;
  assign n881 = ~n879 & ~n880 ;
  assign n882 = x106 & ~n785 ;
  assign n883 = x74 & n785 ;
  assign n884 = ~n882 & ~n883 ;
  assign n885 = ~n881 & n884 ;
  assign n886 = ~n878 & ~n885 ;
  assign n887 = ~n877 & n886 ;
  assign n888 = x43 & ~n652 ;
  assign n889 = x11 & n652 ;
  assign n890 = ~n888 & ~n889 ;
  assign n891 = x107 & ~n785 ;
  assign n892 = x75 & n785 ;
  assign n893 = ~n891 & ~n892 ;
  assign n894 = n890 & ~n893 ;
  assign n895 = n881 & ~n884 ;
  assign n896 = ~n894 & ~n895 ;
  assign n897 = ~n887 & n896 ;
  assign n898 = x108 & ~n785 ;
  assign n899 = x76 & n785 ;
  assign n900 = ~n898 & ~n899 ;
  assign n901 = x44 & ~n652 ;
  assign n902 = x12 & n652 ;
  assign n903 = ~n901 & ~n902 ;
  assign n904 = n900 & ~n903 ;
  assign n905 = ~n890 & n893 ;
  assign n906 = ~n904 & ~n905 ;
  assign n907 = ~n897 & n906 ;
  assign n908 = ~n900 & n903 ;
  assign n909 = x109 & ~n785 ;
  assign n910 = x77 & n785 ;
  assign n911 = ~n909 & ~n910 ;
  assign n912 = x45 & ~n652 ;
  assign n913 = x13 & n652 ;
  assign n914 = ~n912 & ~n913 ;
  assign n915 = ~n911 & n914 ;
  assign n916 = ~n908 & ~n915 ;
  assign n917 = ~n907 & n916 ;
  assign n918 = n911 & ~n914 ;
  assign n919 = x46 & ~n652 ;
  assign n920 = x14 & n652 ;
  assign n921 = ~n919 & ~n920 ;
  assign n922 = x110 & ~n785 ;
  assign n923 = x78 & n785 ;
  assign n924 = ~n922 & ~n923 ;
  assign n925 = ~n921 & n924 ;
  assign n926 = ~n918 & ~n925 ;
  assign n927 = ~n917 & n926 ;
  assign n928 = x47 & ~n652 ;
  assign n929 = x15 & n652 ;
  assign n930 = ~n928 & ~n929 ;
  assign n931 = x111 & ~n785 ;
  assign n932 = x79 & n785 ;
  assign n933 = ~n931 & ~n932 ;
  assign n934 = n930 & ~n933 ;
  assign n935 = n921 & ~n924 ;
  assign n936 = ~n934 & ~n935 ;
  assign n937 = ~n927 & n936 ;
  assign n938 = x112 & ~n785 ;
  assign n939 = x80 & n785 ;
  assign n940 = ~n938 & ~n939 ;
  assign n941 = x48 & ~n652 ;
  assign n942 = x16 & n652 ;
  assign n943 = ~n941 & ~n942 ;
  assign n944 = n940 & ~n943 ;
  assign n945 = ~n930 & n933 ;
  assign n946 = ~n944 & ~n945 ;
  assign n947 = ~n937 & n946 ;
  assign n948 = ~n940 & n943 ;
  assign n949 = x113 & ~n785 ;
  assign n950 = x81 & n785 ;
  assign n951 = ~n949 & ~n950 ;
  assign n952 = x49 & ~n652 ;
  assign n953 = x17 & n652 ;
  assign n954 = ~n952 & ~n953 ;
  assign n955 = ~n951 & n954 ;
  assign n956 = ~n948 & ~n955 ;
  assign n957 = ~n947 & n956 ;
  assign n958 = n951 & ~n954 ;
  assign n959 = x50 & ~n652 ;
  assign n960 = x18 & n652 ;
  assign n961 = ~n959 & ~n960 ;
  assign n962 = x114 & ~n785 ;
  assign n963 = x82 & n785 ;
  assign n964 = ~n962 & ~n963 ;
  assign n965 = ~n961 & n964 ;
  assign n966 = ~n958 & ~n965 ;
  assign n967 = ~n957 & n966 ;
  assign n968 = x51 & ~n652 ;
  assign n969 = x19 & n652 ;
  assign n970 = ~n968 & ~n969 ;
  assign n971 = x115 & ~n785 ;
  assign n972 = x83 & n785 ;
  assign n973 = ~n971 & ~n972 ;
  assign n974 = n970 & ~n973 ;
  assign n975 = n961 & ~n964 ;
  assign n976 = ~n974 & ~n975 ;
  assign n977 = ~n967 & n976 ;
  assign n978 = x116 & ~n785 ;
  assign n979 = x84 & n785 ;
  assign n980 = ~n978 & ~n979 ;
  assign n981 = x52 & ~n652 ;
  assign n982 = x20 & n652 ;
  assign n983 = ~n981 & ~n982 ;
  assign n984 = n980 & ~n983 ;
  assign n985 = ~n970 & n973 ;
  assign n986 = ~n984 & ~n985 ;
  assign n987 = ~n977 & n986 ;
  assign n988 = ~n980 & n983 ;
  assign n989 = x117 & ~n785 ;
  assign n990 = x85 & n785 ;
  assign n991 = ~n989 & ~n990 ;
  assign n992 = x53 & ~n652 ;
  assign n993 = x21 & n652 ;
  assign n994 = ~n992 & ~n993 ;
  assign n995 = ~n991 & n994 ;
  assign n996 = ~n988 & ~n995 ;
  assign n997 = ~n987 & n996 ;
  assign n998 = n991 & ~n994 ;
  assign n999 = x54 & ~n652 ;
  assign n1000 = x22 & n652 ;
  assign n1001 = ~n999 & ~n1000 ;
  assign n1002 = x118 & ~n785 ;
  assign n1003 = x86 & n785 ;
  assign n1004 = ~n1002 & ~n1003 ;
  assign n1005 = ~n1001 & n1004 ;
  assign n1006 = ~n998 & ~n1005 ;
  assign n1007 = ~n997 & n1006 ;
  assign n1008 = x55 & ~n652 ;
  assign n1009 = x23 & n652 ;
  assign n1010 = ~n1008 & ~n1009 ;
  assign n1011 = x119 & ~n785 ;
  assign n1012 = x87 & n785 ;
  assign n1013 = ~n1011 & ~n1012 ;
  assign n1014 = n1010 & ~n1013 ;
  assign n1015 = n1001 & ~n1004 ;
  assign n1016 = ~n1014 & ~n1015 ;
  assign n1017 = ~n1007 & n1016 ;
  assign n1018 = x120 & ~n785 ;
  assign n1019 = x88 & n785 ;
  assign n1020 = ~n1018 & ~n1019 ;
  assign n1021 = x56 & ~n652 ;
  assign n1022 = x24 & n652 ;
  assign n1023 = ~n1021 & ~n1022 ;
  assign n1024 = n1020 & ~n1023 ;
  assign n1025 = ~n1010 & n1013 ;
  assign n1026 = ~n1024 & ~n1025 ;
  assign n1027 = ~n1017 & n1026 ;
  assign n1028 = ~n1020 & n1023 ;
  assign n1029 = x121 & ~n785 ;
  assign n1030 = x89 & n785 ;
  assign n1031 = ~n1029 & ~n1030 ;
  assign n1032 = x57 & ~n652 ;
  assign n1033 = x25 & n652 ;
  assign n1034 = ~n1032 & ~n1033 ;
  assign n1035 = ~n1031 & n1034 ;
  assign n1036 = ~n1028 & ~n1035 ;
  assign n1037 = ~n1027 & n1036 ;
  assign n1038 = n1031 & ~n1034 ;
  assign n1039 = x58 & ~n652 ;
  assign n1040 = x26 & n652 ;
  assign n1041 = ~n1039 & ~n1040 ;
  assign n1042 = x122 & ~n785 ;
  assign n1043 = x90 & n785 ;
  assign n1044 = ~n1042 & ~n1043 ;
  assign n1045 = ~n1041 & n1044 ;
  assign n1046 = ~n1038 & ~n1045 ;
  assign n1047 = ~n1037 & n1046 ;
  assign n1048 = x123 & ~n785 ;
  assign n1049 = x91 & n785 ;
  assign n1050 = ~n1048 & ~n1049 ;
  assign n1051 = n655 & ~n1050 ;
  assign n1052 = n1041 & ~n1044 ;
  assign n1053 = ~n1051 & ~n1052 ;
  assign n1054 = ~n1047 & n1053 ;
  assign n1055 = x124 & ~n785 ;
  assign n1056 = x92 & n785 ;
  assign n1057 = ~n1055 & ~n1056 ;
  assign n1058 = x60 & ~n652 ;
  assign n1059 = x28 & n652 ;
  assign n1060 = ~n1058 & ~n1059 ;
  assign n1061 = n1057 & ~n1060 ;
  assign n1062 = ~n655 & n1050 ;
  assign n1063 = ~n1061 & ~n1062 ;
  assign n1064 = ~n1054 & n1063 ;
  assign n1065 = ~n1057 & n1060 ;
  assign n1066 = x125 & ~n785 ;
  assign n1067 = x93 & n785 ;
  assign n1068 = ~n1066 & ~n1067 ;
  assign n1069 = x61 & ~n652 ;
  assign n1070 = x29 & n652 ;
  assign n1071 = ~n1069 & ~n1070 ;
  assign n1072 = ~n1068 & n1071 ;
  assign n1073 = ~n1065 & ~n1072 ;
  assign n1074 = ~n1064 & n1073 ;
  assign n1075 = n1068 & ~n1071 ;
  assign n1076 = x62 & ~n652 ;
  assign n1077 = x30 & n652 ;
  assign n1078 = ~n1076 & ~n1077 ;
  assign n1079 = x126 & ~n785 ;
  assign n1080 = x94 & n785 ;
  assign n1081 = ~n1079 & ~n1080 ;
  assign n1082 = ~n1078 & n1081 ;
  assign n1083 = ~n1075 & ~n1082 ;
  assign n1084 = ~n1074 & n1083 ;
  assign n1085 = n1078 & ~n1081 ;
  assign n1086 = ~n1084 & ~n1085 ;
  assign n1087 = ~n657 & ~n1086 ;
  assign n1088 = ~n656 & ~n1087 ;
  assign n1089 = ~n655 & n1088 ;
  assign n1090 = ~n1050 & ~n1088 ;
  assign n1091 = ~n1089 & ~n1090 ;
  assign n1092 = ~n522 & n525 ;
  assign n1093 = ~n660 & n1088 ;
  assign n1094 = ~n788 & ~n1088 ;
  assign n1095 = ~n1093 & ~n1094 ;
  assign n1096 = ~x159 & x191 ;
  assign n1097 = x159 & ~x191 ;
  assign n1098 = ~x158 & x190 ;
  assign n1099 = x158 & ~x190 ;
  assign n1100 = ~x157 & x189 ;
  assign n1101 = x157 & ~x189 ;
  assign n1102 = ~x156 & x188 ;
  assign n1103 = x156 & ~x188 ;
  assign n1104 = ~x155 & x187 ;
  assign n1105 = x155 & ~x187 ;
  assign n1106 = ~x154 & x186 ;
  assign n1107 = x154 & ~x186 ;
  assign n1108 = ~x153 & x185 ;
  assign n1109 = x153 & ~x185 ;
  assign n1110 = ~x152 & x184 ;
  assign n1111 = x152 & ~x184 ;
  assign n1112 = ~x151 & x183 ;
  assign n1113 = x151 & ~x183 ;
  assign n1114 = ~x150 & x182 ;
  assign n1115 = x150 & ~x182 ;
  assign n1116 = ~x149 & x181 ;
  assign n1117 = x149 & ~x181 ;
  assign n1118 = ~x148 & x180 ;
  assign n1119 = x148 & ~x180 ;
  assign n1120 = ~x147 & x179 ;
  assign n1121 = x147 & ~x179 ;
  assign n1122 = ~x146 & x178 ;
  assign n1123 = x146 & ~x178 ;
  assign n1124 = ~x145 & x177 ;
  assign n1125 = x145 & ~x177 ;
  assign n1126 = ~x144 & x176 ;
  assign n1127 = x144 & ~x176 ;
  assign n1128 = ~x143 & x175 ;
  assign n1129 = x143 & ~x175 ;
  assign n1130 = ~x142 & x174 ;
  assign n1131 = x142 & ~x174 ;
  assign n1132 = ~x141 & x173 ;
  assign n1133 = x141 & ~x173 ;
  assign n1134 = ~x140 & x172 ;
  assign n1135 = x140 & ~x172 ;
  assign n1136 = ~x139 & x171 ;
  assign n1137 = x139 & ~x171 ;
  assign n1138 = ~x138 & x170 ;
  assign n1139 = x138 & ~x170 ;
  assign n1140 = ~x137 & x169 ;
  assign n1141 = x137 & ~x169 ;
  assign n1142 = ~x136 & x168 ;
  assign n1143 = x136 & ~x168 ;
  assign n1144 = ~x135 & x167 ;
  assign n1145 = x135 & ~x167 ;
  assign n1146 = ~x134 & x166 ;
  assign n1147 = x134 & ~x166 ;
  assign n1148 = ~x133 & x165 ;
  assign n1149 = x133 & ~x165 ;
  assign n1150 = ~x132 & x164 ;
  assign n1151 = x132 & ~x164 ;
  assign n1152 = ~x131 & x163 ;
  assign n1153 = x131 & ~x163 ;
  assign n1154 = ~x130 & x162 ;
  assign n1155 = x130 & ~x162 ;
  assign n1156 = ~x129 & x161 ;
  assign n1157 = x129 & ~x161 ;
  assign n1158 = x128 & ~x160 ;
  assign n1159 = ~n1157 & ~n1158 ;
  assign n1160 = ~n1156 & ~n1159 ;
  assign n1161 = ~n1155 & ~n1160 ;
  assign n1162 = ~n1154 & ~n1161 ;
  assign n1163 = ~n1153 & ~n1162 ;
  assign n1164 = ~n1152 & ~n1163 ;
  assign n1165 = ~n1151 & ~n1164 ;
  assign n1166 = ~n1150 & ~n1165 ;
  assign n1167 = ~n1149 & ~n1166 ;
  assign n1168 = ~n1148 & ~n1167 ;
  assign n1169 = ~n1147 & ~n1168 ;
  assign n1170 = ~n1146 & ~n1169 ;
  assign n1171 = ~n1145 & ~n1170 ;
  assign n1172 = ~n1144 & ~n1171 ;
  assign n1173 = ~n1143 & ~n1172 ;
  assign n1174 = ~n1142 & ~n1173 ;
  assign n1175 = ~n1141 & ~n1174 ;
  assign n1176 = ~n1140 & ~n1175 ;
  assign n1177 = ~n1139 & ~n1176 ;
  assign n1178 = ~n1138 & ~n1177 ;
  assign n1179 = ~n1137 & ~n1178 ;
  assign n1180 = ~n1136 & ~n1179 ;
  assign n1181 = ~n1135 & ~n1180 ;
  assign n1182 = ~n1134 & ~n1181 ;
  assign n1183 = ~n1133 & ~n1182 ;
  assign n1184 = ~n1132 & ~n1183 ;
  assign n1185 = ~n1131 & ~n1184 ;
  assign n1186 = ~n1130 & ~n1185 ;
  assign n1187 = ~n1129 & ~n1186 ;
  assign n1188 = ~n1128 & ~n1187 ;
  assign n1189 = ~n1127 & ~n1188 ;
  assign n1190 = ~n1126 & ~n1189 ;
  assign n1191 = ~n1125 & ~n1190 ;
  assign n1192 = ~n1124 & ~n1191 ;
  assign n1193 = ~n1123 & ~n1192 ;
  assign n1194 = ~n1122 & ~n1193 ;
  assign n1195 = ~n1121 & ~n1194 ;
  assign n1196 = ~n1120 & ~n1195 ;
  assign n1197 = ~n1119 & ~n1196 ;
  assign n1198 = ~n1118 & ~n1197 ;
  assign n1199 = ~n1117 & ~n1198 ;
  assign n1200 = ~n1116 & ~n1199 ;
  assign n1201 = ~n1115 & ~n1200 ;
  assign n1202 = ~n1114 & ~n1201 ;
  assign n1203 = ~n1113 & ~n1202 ;
  assign n1204 = ~n1112 & ~n1203 ;
  assign n1205 = ~n1111 & ~n1204 ;
  assign n1206 = ~n1110 & ~n1205 ;
  assign n1207 = ~n1109 & ~n1206 ;
  assign n1208 = ~n1108 & ~n1207 ;
  assign n1209 = ~n1107 & ~n1208 ;
  assign n1210 = ~n1106 & ~n1209 ;
  assign n1211 = ~n1105 & ~n1210 ;
  assign n1212 = ~n1104 & ~n1211 ;
  assign n1213 = ~n1103 & ~n1212 ;
  assign n1214 = ~n1102 & ~n1213 ;
  assign n1215 = ~n1101 & ~n1214 ;
  assign n1216 = ~n1100 & ~n1215 ;
  assign n1217 = ~n1099 & ~n1216 ;
  assign n1218 = ~n1098 & ~n1217 ;
  assign n1219 = ~n1097 & ~n1218 ;
  assign n1220 = ~n1096 & ~n1219 ;
  assign n1221 = x161 & ~n1220 ;
  assign n1222 = x129 & n1220 ;
  assign n1223 = ~n1221 & ~n1222 ;
  assign n1224 = n523 & ~n524 ;
  assign n1225 = ~n523 & n524 ;
  assign n1226 = ~x223 & x255 ;
  assign n1227 = x223 & ~x255 ;
  assign n1228 = ~x222 & x254 ;
  assign n1229 = x222 & ~x254 ;
  assign n1230 = ~x221 & x253 ;
  assign n1231 = x221 & ~x253 ;
  assign n1232 = ~x220 & x252 ;
  assign n1233 = x220 & ~x252 ;
  assign n1234 = ~x219 & x251 ;
  assign n1235 = x219 & ~x251 ;
  assign n1236 = ~x218 & x250 ;
  assign n1237 = x218 & ~x250 ;
  assign n1238 = ~x217 & x249 ;
  assign n1239 = x217 & ~x249 ;
  assign n1240 = ~x216 & x248 ;
  assign n1241 = x216 & ~x248 ;
  assign n1242 = ~x215 & x247 ;
  assign n1243 = x215 & ~x247 ;
  assign n1244 = ~x214 & x246 ;
  assign n1245 = x214 & ~x246 ;
  assign n1246 = ~x213 & x245 ;
  assign n1247 = x213 & ~x245 ;
  assign n1248 = ~x212 & x244 ;
  assign n1249 = x212 & ~x244 ;
  assign n1250 = ~x211 & x243 ;
  assign n1251 = x211 & ~x243 ;
  assign n1252 = ~x210 & x242 ;
  assign n1253 = x210 & ~x242 ;
  assign n1254 = ~x209 & x241 ;
  assign n1255 = x209 & ~x241 ;
  assign n1256 = ~x208 & x240 ;
  assign n1257 = x208 & ~x240 ;
  assign n1258 = ~x207 & x239 ;
  assign n1259 = x207 & ~x239 ;
  assign n1260 = ~x206 & x238 ;
  assign n1261 = x206 & ~x238 ;
  assign n1262 = ~x205 & x237 ;
  assign n1263 = x205 & ~x237 ;
  assign n1264 = ~x204 & x236 ;
  assign n1265 = x204 & ~x236 ;
  assign n1266 = ~x203 & x235 ;
  assign n1267 = x203 & ~x235 ;
  assign n1268 = ~x202 & x234 ;
  assign n1269 = x202 & ~x234 ;
  assign n1270 = ~x201 & x233 ;
  assign n1271 = x201 & ~x233 ;
  assign n1272 = ~x200 & x232 ;
  assign n1273 = x200 & ~x232 ;
  assign n1274 = ~x199 & x231 ;
  assign n1275 = x199 & ~x231 ;
  assign n1276 = ~x198 & x230 ;
  assign n1277 = x198 & ~x230 ;
  assign n1278 = ~x197 & x229 ;
  assign n1279 = x197 & ~x229 ;
  assign n1280 = ~x196 & x228 ;
  assign n1281 = x196 & ~x228 ;
  assign n1282 = ~x195 & x227 ;
  assign n1283 = x195 & ~x227 ;
  assign n1284 = ~x194 & x226 ;
  assign n1285 = x194 & ~x226 ;
  assign n1286 = ~x193 & x225 ;
  assign n1287 = x193 & ~x225 ;
  assign n1288 = x192 & ~x224 ;
  assign n1289 = ~n1287 & ~n1288 ;
  assign n1290 = ~n1286 & ~n1289 ;
  assign n1291 = ~n1285 & ~n1290 ;
  assign n1292 = ~n1284 & ~n1291 ;
  assign n1293 = ~n1283 & ~n1292 ;
  assign n1294 = ~n1282 & ~n1293 ;
  assign n1295 = ~n1281 & ~n1294 ;
  assign n1296 = ~n1280 & ~n1295 ;
  assign n1297 = ~n1279 & ~n1296 ;
  assign n1298 = ~n1278 & ~n1297 ;
  assign n1299 = ~n1277 & ~n1298 ;
  assign n1300 = ~n1276 & ~n1299 ;
  assign n1301 = ~n1275 & ~n1300 ;
  assign n1302 = ~n1274 & ~n1301 ;
  assign n1303 = ~n1273 & ~n1302 ;
  assign n1304 = ~n1272 & ~n1303 ;
  assign n1305 = ~n1271 & ~n1304 ;
  assign n1306 = ~n1270 & ~n1305 ;
  assign n1307 = ~n1269 & ~n1306 ;
  assign n1308 = ~n1268 & ~n1307 ;
  assign n1309 = ~n1267 & ~n1308 ;
  assign n1310 = ~n1266 & ~n1309 ;
  assign n1311 = ~n1265 & ~n1310 ;
  assign n1312 = ~n1264 & ~n1311 ;
  assign n1313 = ~n1263 & ~n1312 ;
  assign n1314 = ~n1262 & ~n1313 ;
  assign n1315 = ~n1261 & ~n1314 ;
  assign n1316 = ~n1260 & ~n1315 ;
  assign n1317 = ~n1259 & ~n1316 ;
  assign n1318 = ~n1258 & ~n1317 ;
  assign n1319 = ~n1257 & ~n1318 ;
  assign n1320 = ~n1256 & ~n1319 ;
  assign n1321 = ~n1255 & ~n1320 ;
  assign n1322 = ~n1254 & ~n1321 ;
  assign n1323 = ~n1253 & ~n1322 ;
  assign n1324 = ~n1252 & ~n1323 ;
  assign n1325 = ~n1251 & ~n1324 ;
  assign n1326 = ~n1250 & ~n1325 ;
  assign n1327 = ~n1249 & ~n1326 ;
  assign n1328 = ~n1248 & ~n1327 ;
  assign n1329 = ~n1247 & ~n1328 ;
  assign n1330 = ~n1246 & ~n1329 ;
  assign n1331 = ~n1245 & ~n1330 ;
  assign n1332 = ~n1244 & ~n1331 ;
  assign n1333 = ~n1243 & ~n1332 ;
  assign n1334 = ~n1242 & ~n1333 ;
  assign n1335 = ~n1241 & ~n1334 ;
  assign n1336 = ~n1240 & ~n1335 ;
  assign n1337 = ~n1239 & ~n1336 ;
  assign n1338 = ~n1238 & ~n1337 ;
  assign n1339 = ~n1237 & ~n1338 ;
  assign n1340 = ~n1236 & ~n1339 ;
  assign n1341 = ~n1235 & ~n1340 ;
  assign n1342 = ~n1234 & ~n1341 ;
  assign n1343 = ~n1233 & ~n1342 ;
  assign n1344 = ~n1232 & ~n1343 ;
  assign n1345 = ~n1231 & ~n1344 ;
  assign n1346 = ~n1230 & ~n1345 ;
  assign n1347 = ~n1229 & ~n1346 ;
  assign n1348 = ~n1228 & ~n1347 ;
  assign n1349 = ~n1227 & ~n1348 ;
  assign n1350 = ~n1226 & ~n1349 ;
  assign n1351 = x254 & ~n1350 ;
  assign n1352 = x222 & n1350 ;
  assign n1353 = ~n1351 & ~n1352 ;
  assign n1354 = x190 & ~n1220 ;
  assign n1355 = x158 & n1220 ;
  assign n1356 = ~n1354 & ~n1355 ;
  assign n1357 = ~n1353 & n1356 ;
  assign n1358 = x225 & ~n1350 ;
  assign n1359 = x193 & n1350 ;
  assign n1360 = ~n1358 & ~n1359 ;
  assign n1361 = n1223 & ~n1360 ;
  assign n1362 = x224 & ~n1350 ;
  assign n1363 = x192 & n1350 ;
  assign n1364 = ~n1362 & ~n1363 ;
  assign n1365 = x160 & ~n1220 ;
  assign n1366 = x128 & n1220 ;
  assign n1367 = ~n1365 & ~n1366 ;
  assign n1368 = n1364 & ~n1367 ;
  assign n1369 = ~n1361 & n1368 ;
  assign n1370 = x226 & ~n1350 ;
  assign n1371 = x194 & n1350 ;
  assign n1372 = ~n1370 & ~n1371 ;
  assign n1373 = x162 & ~n1220 ;
  assign n1374 = x130 & n1220 ;
  assign n1375 = ~n1373 & ~n1374 ;
  assign n1376 = n1372 & ~n1375 ;
  assign n1377 = ~n1223 & n1360 ;
  assign n1378 = ~n1376 & ~n1377 ;
  assign n1379 = ~n1369 & n1378 ;
  assign n1380 = x227 & ~n1350 ;
  assign n1381 = x195 & n1350 ;
  assign n1382 = ~n1380 & ~n1381 ;
  assign n1383 = x163 & ~n1220 ;
  assign n1384 = x131 & n1220 ;
  assign n1385 = ~n1383 & ~n1384 ;
  assign n1386 = ~n1382 & n1385 ;
  assign n1387 = ~n1372 & n1375 ;
  assign n1388 = ~n1386 & ~n1387 ;
  assign n1389 = ~n1379 & n1388 ;
  assign n1390 = x228 & ~n1350 ;
  assign n1391 = x196 & n1350 ;
  assign n1392 = ~n1390 & ~n1391 ;
  assign n1393 = x164 & ~n1220 ;
  assign n1394 = x132 & n1220 ;
  assign n1395 = ~n1393 & ~n1394 ;
  assign n1396 = n1392 & ~n1395 ;
  assign n1397 = n1382 & ~n1385 ;
  assign n1398 = ~n1396 & ~n1397 ;
  assign n1399 = ~n1389 & n1398 ;
  assign n1400 = x229 & ~n1350 ;
  assign n1401 = x197 & n1350 ;
  assign n1402 = ~n1400 & ~n1401 ;
  assign n1403 = x165 & ~n1220 ;
  assign n1404 = x133 & n1220 ;
  assign n1405 = ~n1403 & ~n1404 ;
  assign n1406 = ~n1402 & n1405 ;
  assign n1407 = ~n1392 & n1395 ;
  assign n1408 = ~n1406 & ~n1407 ;
  assign n1409 = ~n1399 & n1408 ;
  assign n1410 = n1402 & ~n1405 ;
  assign n1411 = x166 & ~n1220 ;
  assign n1412 = x134 & n1220 ;
  assign n1413 = ~n1411 & ~n1412 ;
  assign n1414 = x230 & ~n1350 ;
  assign n1415 = x198 & n1350 ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = ~n1413 & n1416 ;
  assign n1418 = ~n1410 & ~n1417 ;
  assign n1419 = ~n1409 & n1418 ;
  assign n1420 = x167 & ~n1220 ;
  assign n1421 = x135 & n1220 ;
  assign n1422 = ~n1420 & ~n1421 ;
  assign n1423 = x231 & ~n1350 ;
  assign n1424 = x199 & n1350 ;
  assign n1425 = ~n1423 & ~n1424 ;
  assign n1426 = n1422 & ~n1425 ;
  assign n1427 = n1413 & ~n1416 ;
  assign n1428 = ~n1426 & ~n1427 ;
  assign n1429 = ~n1419 & n1428 ;
  assign n1430 = ~n1422 & n1425 ;
  assign n1431 = x232 & ~n1350 ;
  assign n1432 = x200 & n1350 ;
  assign n1433 = ~n1431 & ~n1432 ;
  assign n1434 = x168 & ~n1220 ;
  assign n1435 = x136 & n1220 ;
  assign n1436 = ~n1434 & ~n1435 ;
  assign n1437 = n1433 & ~n1436 ;
  assign n1438 = ~n1430 & ~n1437 ;
  assign n1439 = ~n1429 & n1438 ;
  assign n1440 = ~n1433 & n1436 ;
  assign n1441 = x233 & ~n1350 ;
  assign n1442 = x201 & n1350 ;
  assign n1443 = ~n1441 & ~n1442 ;
  assign n1444 = x169 & ~n1220 ;
  assign n1445 = x137 & n1220 ;
  assign n1446 = ~n1444 & ~n1445 ;
  assign n1447 = ~n1443 & n1446 ;
  assign n1448 = ~n1440 & ~n1447 ;
  assign n1449 = ~n1439 & n1448 ;
  assign n1450 = n1443 & ~n1446 ;
  assign n1451 = x170 & ~n1220 ;
  assign n1452 = x138 & n1220 ;
  assign n1453 = ~n1451 & ~n1452 ;
  assign n1454 = x234 & ~n1350 ;
  assign n1455 = x202 & n1350 ;
  assign n1456 = ~n1454 & ~n1455 ;
  assign n1457 = ~n1453 & n1456 ;
  assign n1458 = ~n1450 & ~n1457 ;
  assign n1459 = ~n1449 & n1458 ;
  assign n1460 = x171 & ~n1220 ;
  assign n1461 = x139 & n1220 ;
  assign n1462 = ~n1460 & ~n1461 ;
  assign n1463 = x235 & ~n1350 ;
  assign n1464 = x203 & n1350 ;
  assign n1465 = ~n1463 & ~n1464 ;
  assign n1466 = n1462 & ~n1465 ;
  assign n1467 = n1453 & ~n1456 ;
  assign n1468 = ~n1466 & ~n1467 ;
  assign n1469 = ~n1459 & n1468 ;
  assign n1470 = x236 & ~n1350 ;
  assign n1471 = x204 & n1350 ;
  assign n1472 = ~n1470 & ~n1471 ;
  assign n1473 = x172 & ~n1220 ;
  assign n1474 = x140 & n1220 ;
  assign n1475 = ~n1473 & ~n1474 ;
  assign n1476 = n1472 & ~n1475 ;
  assign n1477 = ~n1462 & n1465 ;
  assign n1478 = ~n1476 & ~n1477 ;
  assign n1479 = ~n1469 & n1478 ;
  assign n1480 = ~n1472 & n1475 ;
  assign n1481 = x237 & ~n1350 ;
  assign n1482 = x205 & n1350 ;
  assign n1483 = ~n1481 & ~n1482 ;
  assign n1484 = x173 & ~n1220 ;
  assign n1485 = x141 & n1220 ;
  assign n1486 = ~n1484 & ~n1485 ;
  assign n1487 = ~n1483 & n1486 ;
  assign n1488 = ~n1480 & ~n1487 ;
  assign n1489 = ~n1479 & n1488 ;
  assign n1490 = n1483 & ~n1486 ;
  assign n1491 = x174 & ~n1220 ;
  assign n1492 = x142 & n1220 ;
  assign n1493 = ~n1491 & ~n1492 ;
  assign n1494 = x238 & ~n1350 ;
  assign n1495 = x206 & n1350 ;
  assign n1496 = ~n1494 & ~n1495 ;
  assign n1497 = ~n1493 & n1496 ;
  assign n1498 = ~n1490 & ~n1497 ;
  assign n1499 = ~n1489 & n1498 ;
  assign n1500 = x175 & ~n1220 ;
  assign n1501 = x143 & n1220 ;
  assign n1502 = ~n1500 & ~n1501 ;
  assign n1503 = x239 & ~n1350 ;
  assign n1504 = x207 & n1350 ;
  assign n1505 = ~n1503 & ~n1504 ;
  assign n1506 = n1502 & ~n1505 ;
  assign n1507 = n1493 & ~n1496 ;
  assign n1508 = ~n1506 & ~n1507 ;
  assign n1509 = ~n1499 & n1508 ;
  assign n1510 = x240 & ~n1350 ;
  assign n1511 = x208 & n1350 ;
  assign n1512 = ~n1510 & ~n1511 ;
  assign n1513 = x176 & ~n1220 ;
  assign n1514 = x144 & n1220 ;
  assign n1515 = ~n1513 & ~n1514 ;
  assign n1516 = n1512 & ~n1515 ;
  assign n1517 = ~n1502 & n1505 ;
  assign n1518 = ~n1516 & ~n1517 ;
  assign n1519 = ~n1509 & n1518 ;
  assign n1520 = ~n1512 & n1515 ;
  assign n1521 = x241 & ~n1350 ;
  assign n1522 = x209 & n1350 ;
  assign n1523 = ~n1521 & ~n1522 ;
  assign n1524 = x177 & ~n1220 ;
  assign n1525 = x145 & n1220 ;
  assign n1526 = ~n1524 & ~n1525 ;
  assign n1527 = ~n1523 & n1526 ;
  assign n1528 = ~n1520 & ~n1527 ;
  assign n1529 = ~n1519 & n1528 ;
  assign n1530 = n1523 & ~n1526 ;
  assign n1531 = x178 & ~n1220 ;
  assign n1532 = x146 & n1220 ;
  assign n1533 = ~n1531 & ~n1532 ;
  assign n1534 = x242 & ~n1350 ;
  assign n1535 = x210 & n1350 ;
  assign n1536 = ~n1534 & ~n1535 ;
  assign n1537 = ~n1533 & n1536 ;
  assign n1538 = ~n1530 & ~n1537 ;
  assign n1539 = ~n1529 & n1538 ;
  assign n1540 = x179 & ~n1220 ;
  assign n1541 = x147 & n1220 ;
  assign n1542 = ~n1540 & ~n1541 ;
  assign n1543 = x243 & ~n1350 ;
  assign n1544 = x211 & n1350 ;
  assign n1545 = ~n1543 & ~n1544 ;
  assign n1546 = n1542 & ~n1545 ;
  assign n1547 = n1533 & ~n1536 ;
  assign n1548 = ~n1546 & ~n1547 ;
  assign n1549 = ~n1539 & n1548 ;
  assign n1550 = x244 & ~n1350 ;
  assign n1551 = x212 & n1350 ;
  assign n1552 = ~n1550 & ~n1551 ;
  assign n1553 = x180 & ~n1220 ;
  assign n1554 = x148 & n1220 ;
  assign n1555 = ~n1553 & ~n1554 ;
  assign n1556 = n1552 & ~n1555 ;
  assign n1557 = ~n1542 & n1545 ;
  assign n1558 = ~n1556 & ~n1557 ;
  assign n1559 = ~n1549 & n1558 ;
  assign n1560 = ~n1552 & n1555 ;
  assign n1561 = x245 & ~n1350 ;
  assign n1562 = x213 & n1350 ;
  assign n1563 = ~n1561 & ~n1562 ;
  assign n1564 = x181 & ~n1220 ;
  assign n1565 = x149 & n1220 ;
  assign n1566 = ~n1564 & ~n1565 ;
  assign n1567 = ~n1563 & n1566 ;
  assign n1568 = ~n1560 & ~n1567 ;
  assign n1569 = ~n1559 & n1568 ;
  assign n1570 = n1563 & ~n1566 ;
  assign n1571 = x182 & ~n1220 ;
  assign n1572 = x150 & n1220 ;
  assign n1573 = ~n1571 & ~n1572 ;
  assign n1574 = x246 & ~n1350 ;
  assign n1575 = x214 & n1350 ;
  assign n1576 = ~n1574 & ~n1575 ;
  assign n1577 = ~n1573 & n1576 ;
  assign n1578 = ~n1570 & ~n1577 ;
  assign n1579 = ~n1569 & n1578 ;
  assign n1580 = x183 & ~n1220 ;
  assign n1581 = x151 & n1220 ;
  assign n1582 = ~n1580 & ~n1581 ;
  assign n1583 = x247 & ~n1350 ;
  assign n1584 = x215 & n1350 ;
  assign n1585 = ~n1583 & ~n1584 ;
  assign n1586 = n1582 & ~n1585 ;
  assign n1587 = n1573 & ~n1576 ;
  assign n1588 = ~n1586 & ~n1587 ;
  assign n1589 = ~n1579 & n1588 ;
  assign n1590 = x248 & ~n1350 ;
  assign n1591 = x216 & n1350 ;
  assign n1592 = ~n1590 & ~n1591 ;
  assign n1593 = x184 & ~n1220 ;
  assign n1594 = x152 & n1220 ;
  assign n1595 = ~n1593 & ~n1594 ;
  assign n1596 = n1592 & ~n1595 ;
  assign n1597 = ~n1582 & n1585 ;
  assign n1598 = ~n1596 & ~n1597 ;
  assign n1599 = ~n1589 & n1598 ;
  assign n1600 = ~n1592 & n1595 ;
  assign n1601 = x249 & ~n1350 ;
  assign n1602 = x217 & n1350 ;
  assign n1603 = ~n1601 & ~n1602 ;
  assign n1604 = x185 & ~n1220 ;
  assign n1605 = x153 & n1220 ;
  assign n1606 = ~n1604 & ~n1605 ;
  assign n1607 = ~n1603 & n1606 ;
  assign n1608 = ~n1600 & ~n1607 ;
  assign n1609 = ~n1599 & n1608 ;
  assign n1610 = n1603 & ~n1606 ;
  assign n1611 = x186 & ~n1220 ;
  assign n1612 = x154 & n1220 ;
  assign n1613 = ~n1611 & ~n1612 ;
  assign n1614 = x250 & ~n1350 ;
  assign n1615 = x218 & n1350 ;
  assign n1616 = ~n1614 & ~n1615 ;
  assign n1617 = ~n1613 & n1616 ;
  assign n1618 = ~n1610 & ~n1617 ;
  assign n1619 = ~n1609 & n1618 ;
  assign n1620 = x187 & ~n1220 ;
  assign n1621 = x155 & n1220 ;
  assign n1622 = ~n1620 & ~n1621 ;
  assign n1623 = x251 & ~n1350 ;
  assign n1624 = x219 & n1350 ;
  assign n1625 = ~n1623 & ~n1624 ;
  assign n1626 = n1622 & ~n1625 ;
  assign n1627 = n1613 & ~n1616 ;
  assign n1628 = ~n1626 & ~n1627 ;
  assign n1629 = ~n1619 & n1628 ;
  assign n1630 = x252 & ~n1350 ;
  assign n1631 = x220 & n1350 ;
  assign n1632 = ~n1630 & ~n1631 ;
  assign n1633 = x188 & ~n1220 ;
  assign n1634 = x156 & n1220 ;
  assign n1635 = ~n1633 & ~n1634 ;
  assign n1636 = n1632 & ~n1635 ;
  assign n1637 = ~n1622 & n1625 ;
  assign n1638 = ~n1636 & ~n1637 ;
  assign n1639 = ~n1629 & n1638 ;
  assign n1640 = ~n1632 & n1635 ;
  assign n1641 = x253 & ~n1350 ;
  assign n1642 = x221 & n1350 ;
  assign n1643 = ~n1641 & ~n1642 ;
  assign n1644 = x189 & ~n1220 ;
  assign n1645 = x157 & n1220 ;
  assign n1646 = ~n1644 & ~n1645 ;
  assign n1647 = ~n1643 & n1646 ;
  assign n1648 = ~n1640 & ~n1647 ;
  assign n1649 = ~n1639 & n1648 ;
  assign n1650 = n1353 & ~n1356 ;
  assign n1651 = n1643 & ~n1646 ;
  assign n1652 = ~n1650 & ~n1651 ;
  assign n1653 = ~n1649 & n1652 ;
  assign n1654 = ~n1357 & ~n1653 ;
  assign n1655 = ~n1225 & ~n1654 ;
  assign n1656 = ~n1224 & ~n1655 ;
  assign n1657 = ~n1223 & n1656 ;
  assign n1658 = ~n1360 & ~n1656 ;
  assign n1659 = ~n1657 & ~n1658 ;
  assign n1660 = n1095 & ~n1659 ;
  assign n1661 = ~n1367 & n1656 ;
  assign n1662 = ~n1364 & ~n1656 ;
  assign n1663 = ~n1661 & ~n1662 ;
  assign n1664 = ~n792 & n1088 ;
  assign n1665 = ~n795 & ~n1088 ;
  assign n1666 = ~n1664 & ~n1665 ;
  assign n1667 = n1663 & ~n1666 ;
  assign n1668 = ~n1660 & n1667 ;
  assign n1669 = ~n1375 & n1656 ;
  assign n1670 = ~n1372 & ~n1656 ;
  assign n1671 = ~n1669 & ~n1670 ;
  assign n1672 = ~n803 & n1088 ;
  assign n1673 = ~n800 & ~n1088 ;
  assign n1674 = ~n1672 & ~n1673 ;
  assign n1675 = n1671 & ~n1674 ;
  assign n1676 = ~n1095 & n1659 ;
  assign n1677 = ~n1675 & ~n1676 ;
  assign n1678 = ~n1668 & n1677 ;
  assign n1679 = ~n1671 & n1674 ;
  assign n1680 = ~n810 & n1088 ;
  assign n1681 = ~n813 & ~n1088 ;
  assign n1682 = ~n1680 & ~n1681 ;
  assign n1683 = n1382 & ~n1656 ;
  assign n1684 = n1385 & n1656 ;
  assign n1685 = ~n1683 & ~n1684 ;
  assign n1686 = n1682 & n1685 ;
  assign n1687 = ~n1679 & ~n1686 ;
  assign n1688 = ~n1678 & n1687 ;
  assign n1689 = ~n821 & n1088 ;
  assign n1690 = ~n824 & ~n1088 ;
  assign n1691 = ~n1689 & ~n1690 ;
  assign n1692 = ~n1395 & n1656 ;
  assign n1693 = ~n1392 & ~n1656 ;
  assign n1694 = ~n1692 & ~n1693 ;
  assign n1695 = ~n1691 & n1694 ;
  assign n1696 = ~n1682 & ~n1685 ;
  assign n1697 = ~n1695 & ~n1696 ;
  assign n1698 = ~n1688 & n1697 ;
  assign n1699 = ~n834 & n1088 ;
  assign n1700 = ~n831 & ~n1088 ;
  assign n1701 = ~n1699 & ~n1700 ;
  assign n1702 = ~n1405 & n1656 ;
  assign n1703 = ~n1402 & ~n1656 ;
  assign n1704 = ~n1702 & ~n1703 ;
  assign n1705 = n1701 & ~n1704 ;
  assign n1706 = n1691 & ~n1694 ;
  assign n1707 = ~n1705 & ~n1706 ;
  assign n1708 = ~n1698 & n1707 ;
  assign n1709 = ~n1413 & n1656 ;
  assign n1710 = ~n1416 & ~n1656 ;
  assign n1711 = ~n1709 & ~n1710 ;
  assign n1712 = ~n844 & n1088 ;
  assign n1713 = ~n841 & ~n1088 ;
  assign n1714 = ~n1712 & ~n1713 ;
  assign n1715 = n1711 & ~n1714 ;
  assign n1716 = ~n1701 & n1704 ;
  assign n1717 = ~n1715 & ~n1716 ;
  assign n1718 = ~n1708 & n1717 ;
  assign n1719 = ~n851 & n1088 ;
  assign n1720 = ~n854 & ~n1088 ;
  assign n1721 = ~n1719 & ~n1720 ;
  assign n1722 = ~n1422 & n1656 ;
  assign n1723 = ~n1425 & ~n1656 ;
  assign n1724 = ~n1722 & ~n1723 ;
  assign n1725 = n1721 & ~n1724 ;
  assign n1726 = ~n1711 & n1714 ;
  assign n1727 = ~n1725 & ~n1726 ;
  assign n1728 = ~n1718 & n1727 ;
  assign n1729 = ~n1436 & n1656 ;
  assign n1730 = ~n1433 & ~n1656 ;
  assign n1731 = ~n1729 & ~n1730 ;
  assign n1732 = ~n864 & n1088 ;
  assign n1733 = ~n861 & ~n1088 ;
  assign n1734 = ~n1732 & ~n1733 ;
  assign n1735 = n1731 & ~n1734 ;
  assign n1736 = ~n1721 & n1724 ;
  assign n1737 = ~n1735 & ~n1736 ;
  assign n1738 = ~n1728 & n1737 ;
  assign n1739 = ~n874 & n1088 ;
  assign n1740 = ~n871 & ~n1088 ;
  assign n1741 = ~n1739 & ~n1740 ;
  assign n1742 = ~n1446 & n1656 ;
  assign n1743 = ~n1443 & ~n1656 ;
  assign n1744 = ~n1742 & ~n1743 ;
  assign n1745 = n1741 & ~n1744 ;
  assign n1746 = ~n1731 & n1734 ;
  assign n1747 = ~n1745 & ~n1746 ;
  assign n1748 = ~n1738 & n1747 ;
  assign n1749 = ~n1453 & n1656 ;
  assign n1750 = ~n1456 & ~n1656 ;
  assign n1751 = ~n1749 & ~n1750 ;
  assign n1752 = ~n881 & n1088 ;
  assign n1753 = ~n884 & ~n1088 ;
  assign n1754 = ~n1752 & ~n1753 ;
  assign n1755 = n1751 & ~n1754 ;
  assign n1756 = ~n1741 & n1744 ;
  assign n1757 = ~n1755 & ~n1756 ;
  assign n1758 = ~n1748 & n1757 ;
  assign n1759 = ~n890 & n1088 ;
  assign n1760 = ~n893 & ~n1088 ;
  assign n1761 = ~n1759 & ~n1760 ;
  assign n1762 = ~n1462 & n1656 ;
  assign n1763 = ~n1465 & ~n1656 ;
  assign n1764 = ~n1762 & ~n1763 ;
  assign n1765 = n1761 & ~n1764 ;
  assign n1766 = ~n1751 & n1754 ;
  assign n1767 = ~n1765 & ~n1766 ;
  assign n1768 = ~n1758 & n1767 ;
  assign n1769 = ~n1475 & n1656 ;
  assign n1770 = ~n1472 & ~n1656 ;
  assign n1771 = ~n1769 & ~n1770 ;
  assign n1772 = ~n903 & n1088 ;
  assign n1773 = ~n900 & ~n1088 ;
  assign n1774 = ~n1772 & ~n1773 ;
  assign n1775 = n1771 & ~n1774 ;
  assign n1776 = ~n1761 & n1764 ;
  assign n1777 = ~n1775 & ~n1776 ;
  assign n1778 = ~n1768 & n1777 ;
  assign n1779 = ~n914 & n1088 ;
  assign n1780 = ~n911 & ~n1088 ;
  assign n1781 = ~n1779 & ~n1780 ;
  assign n1782 = ~n1486 & n1656 ;
  assign n1783 = ~n1483 & ~n1656 ;
  assign n1784 = ~n1782 & ~n1783 ;
  assign n1785 = n1781 & ~n1784 ;
  assign n1786 = ~n1771 & n1774 ;
  assign n1787 = ~n1785 & ~n1786 ;
  assign n1788 = ~n1778 & n1787 ;
  assign n1789 = ~n1493 & n1656 ;
  assign n1790 = ~n1496 & ~n1656 ;
  assign n1791 = ~n1789 & ~n1790 ;
  assign n1792 = ~n921 & n1088 ;
  assign n1793 = ~n924 & ~n1088 ;
  assign n1794 = ~n1792 & ~n1793 ;
  assign n1795 = n1791 & ~n1794 ;
  assign n1796 = ~n1781 & n1784 ;
  assign n1797 = ~n1795 & ~n1796 ;
  assign n1798 = ~n1788 & n1797 ;
  assign n1799 = ~n930 & n1088 ;
  assign n1800 = ~n933 & ~n1088 ;
  assign n1801 = ~n1799 & ~n1800 ;
  assign n1802 = ~n1502 & n1656 ;
  assign n1803 = ~n1505 & ~n1656 ;
  assign n1804 = ~n1802 & ~n1803 ;
  assign n1805 = n1801 & ~n1804 ;
  assign n1806 = ~n1791 & n1794 ;
  assign n1807 = ~n1805 & ~n1806 ;
  assign n1808 = ~n1798 & n1807 ;
  assign n1809 = ~n1515 & n1656 ;
  assign n1810 = ~n1512 & ~n1656 ;
  assign n1811 = ~n1809 & ~n1810 ;
  assign n1812 = ~n943 & n1088 ;
  assign n1813 = ~n940 & ~n1088 ;
  assign n1814 = ~n1812 & ~n1813 ;
  assign n1815 = n1811 & ~n1814 ;
  assign n1816 = ~n1801 & n1804 ;
  assign n1817 = ~n1815 & ~n1816 ;
  assign n1818 = ~n1808 & n1817 ;
  assign n1819 = ~n954 & n1088 ;
  assign n1820 = ~n951 & ~n1088 ;
  assign n1821 = ~n1819 & ~n1820 ;
  assign n1822 = ~n1526 & n1656 ;
  assign n1823 = ~n1523 & ~n1656 ;
  assign n1824 = ~n1822 & ~n1823 ;
  assign n1825 = n1821 & ~n1824 ;
  assign n1826 = ~n1811 & n1814 ;
  assign n1827 = ~n1825 & ~n1826 ;
  assign n1828 = ~n1818 & n1827 ;
  assign n1829 = ~n1533 & n1656 ;
  assign n1830 = ~n1536 & ~n1656 ;
  assign n1831 = ~n1829 & ~n1830 ;
  assign n1832 = ~n961 & n1088 ;
  assign n1833 = ~n964 & ~n1088 ;
  assign n1834 = ~n1832 & ~n1833 ;
  assign n1835 = n1831 & ~n1834 ;
  assign n1836 = ~n1821 & n1824 ;
  assign n1837 = ~n1835 & ~n1836 ;
  assign n1838 = ~n1828 & n1837 ;
  assign n1839 = ~n970 & n1088 ;
  assign n1840 = ~n973 & ~n1088 ;
  assign n1841 = ~n1839 & ~n1840 ;
  assign n1842 = ~n1542 & n1656 ;
  assign n1843 = ~n1545 & ~n1656 ;
  assign n1844 = ~n1842 & ~n1843 ;
  assign n1845 = n1841 & ~n1844 ;
  assign n1846 = ~n1831 & n1834 ;
  assign n1847 = ~n1845 & ~n1846 ;
  assign n1848 = ~n1838 & n1847 ;
  assign n1849 = ~n1555 & n1656 ;
  assign n1850 = ~n1552 & ~n1656 ;
  assign n1851 = ~n1849 & ~n1850 ;
  assign n1852 = ~n983 & n1088 ;
  assign n1853 = ~n980 & ~n1088 ;
  assign n1854 = ~n1852 & ~n1853 ;
  assign n1855 = n1851 & ~n1854 ;
  assign n1856 = ~n1841 & n1844 ;
  assign n1857 = ~n1855 & ~n1856 ;
  assign n1858 = ~n1848 & n1857 ;
  assign n1859 = ~n994 & n1088 ;
  assign n1860 = ~n991 & ~n1088 ;
  assign n1861 = ~n1859 & ~n1860 ;
  assign n1862 = ~n1566 & n1656 ;
  assign n1863 = ~n1563 & ~n1656 ;
  assign n1864 = ~n1862 & ~n1863 ;
  assign n1865 = n1861 & ~n1864 ;
  assign n1866 = ~n1851 & n1854 ;
  assign n1867 = ~n1865 & ~n1866 ;
  assign n1868 = ~n1858 & n1867 ;
  assign n1869 = ~n1573 & n1656 ;
  assign n1870 = ~n1576 & ~n1656 ;
  assign n1871 = ~n1869 & ~n1870 ;
  assign n1872 = ~n1001 & n1088 ;
  assign n1873 = ~n1004 & ~n1088 ;
  assign n1874 = ~n1872 & ~n1873 ;
  assign n1875 = n1871 & ~n1874 ;
  assign n1876 = ~n1861 & n1864 ;
  assign n1877 = ~n1875 & ~n1876 ;
  assign n1878 = ~n1868 & n1877 ;
  assign n1879 = ~n1010 & n1088 ;
  assign n1880 = ~n1013 & ~n1088 ;
  assign n1881 = ~n1879 & ~n1880 ;
  assign n1882 = ~n1582 & n1656 ;
  assign n1883 = ~n1585 & ~n1656 ;
  assign n1884 = ~n1882 & ~n1883 ;
  assign n1885 = n1881 & ~n1884 ;
  assign n1886 = ~n1871 & n1874 ;
  assign n1887 = ~n1885 & ~n1886 ;
  assign n1888 = ~n1878 & n1887 ;
  assign n1889 = ~n1595 & n1656 ;
  assign n1890 = ~n1592 & ~n1656 ;
  assign n1891 = ~n1889 & ~n1890 ;
  assign n1892 = ~n1023 & n1088 ;
  assign n1893 = ~n1020 & ~n1088 ;
  assign n1894 = ~n1892 & ~n1893 ;
  assign n1895 = n1891 & ~n1894 ;
  assign n1896 = ~n1881 & n1884 ;
  assign n1897 = ~n1895 & ~n1896 ;
  assign n1898 = ~n1888 & n1897 ;
  assign n1899 = ~n1606 & n1656 ;
  assign n1900 = ~n1603 & ~n1656 ;
  assign n1901 = ~n1899 & ~n1900 ;
  assign n1902 = ~n1034 & n1088 ;
  assign n1903 = ~n1031 & ~n1088 ;
  assign n1904 = ~n1902 & ~n1903 ;
  assign n1905 = ~n1901 & n1904 ;
  assign n1906 = ~n1891 & n1894 ;
  assign n1907 = ~n1905 & ~n1906 ;
  assign n1908 = ~n1898 & n1907 ;
  assign n1909 = ~n1613 & n1656 ;
  assign n1910 = ~n1616 & ~n1656 ;
  assign n1911 = ~n1909 & ~n1910 ;
  assign n1912 = ~n1041 & n1088 ;
  assign n1913 = ~n1044 & ~n1088 ;
  assign n1914 = ~n1912 & ~n1913 ;
  assign n1915 = n1911 & ~n1914 ;
  assign n1916 = n1901 & ~n1904 ;
  assign n1917 = ~n1915 & ~n1916 ;
  assign n1918 = ~n1908 & n1917 ;
  assign n1919 = ~n1911 & n1914 ;
  assign n1920 = ~n1622 & n1656 ;
  assign n1921 = ~n1625 & ~n1656 ;
  assign n1922 = ~n1920 & ~n1921 ;
  assign n1923 = n1091 & ~n1922 ;
  assign n1924 = ~n1919 & ~n1923 ;
  assign n1925 = ~n1918 & n1924 ;
  assign n1926 = ~n1091 & n1922 ;
  assign n1927 = ~n1060 & n1088 ;
  assign n1928 = ~n1057 & ~n1088 ;
  assign n1929 = ~n1927 & ~n1928 ;
  assign n1930 = ~n1635 & n1656 ;
  assign n1931 = ~n1632 & ~n1656 ;
  assign n1932 = ~n1930 & ~n1931 ;
  assign n1933 = ~n1929 & n1932 ;
  assign n1934 = ~n1926 & ~n1933 ;
  assign n1935 = ~n1925 & n1934 ;
  assign n1936 = n1929 & ~n1932 ;
  assign n1937 = ~n1071 & n1088 ;
  assign n1938 = ~n1068 & ~n1088 ;
  assign n1939 = ~n1937 & ~n1938 ;
  assign n1940 = ~n1646 & n1656 ;
  assign n1941 = ~n1643 & ~n1656 ;
  assign n1942 = ~n1940 & ~n1941 ;
  assign n1943 = n1939 & ~n1942 ;
  assign n1944 = ~n1936 & ~n1943 ;
  assign n1945 = ~n1935 & n1944 ;
  assign n1946 = ~n1939 & n1942 ;
  assign n1947 = ~n1078 & n1088 ;
  assign n1948 = ~n1081 & ~n1088 ;
  assign n1949 = ~n1947 & ~n1948 ;
  assign n1950 = ~n1356 & n1656 ;
  assign n1951 = ~n1353 & ~n1656 ;
  assign n1952 = ~n1950 & ~n1951 ;
  assign n1953 = ~n1949 & n1952 ;
  assign n1954 = ~n1946 & ~n1953 ;
  assign n1955 = ~n1945 & n1954 ;
  assign n1956 = n522 & ~n525 ;
  assign n1957 = n1949 & ~n1952 ;
  assign n1958 = ~n1956 & ~n1957 ;
  assign n1959 = ~n1955 & n1958 ;
  assign n1960 = ~n1092 & ~n1959 ;
  assign n1961 = n1091 & ~n1960 ;
  assign n1962 = n1922 & n1960 ;
  assign n1963 = ~n1961 & ~n1962 ;
  assign n1964 = ~x287 & x319 ;
  assign n1965 = x287 & ~x319 ;
  assign n1966 = ~x286 & x318 ;
  assign n1967 = x286 & ~x318 ;
  assign n1968 = ~x285 & x317 ;
  assign n1969 = x285 & ~x317 ;
  assign n1970 = ~x284 & x316 ;
  assign n1971 = x284 & ~x316 ;
  assign n1972 = ~x283 & x315 ;
  assign n1973 = x283 & ~x315 ;
  assign n1974 = ~x282 & x314 ;
  assign n1975 = x282 & ~x314 ;
  assign n1976 = ~x281 & x313 ;
  assign n1977 = x281 & ~x313 ;
  assign n1978 = ~x280 & x312 ;
  assign n1979 = x280 & ~x312 ;
  assign n1980 = ~x279 & x311 ;
  assign n1981 = x279 & ~x311 ;
  assign n1982 = ~x278 & x310 ;
  assign n1983 = x278 & ~x310 ;
  assign n1984 = ~x277 & x309 ;
  assign n1985 = x277 & ~x309 ;
  assign n1986 = ~x276 & x308 ;
  assign n1987 = x276 & ~x308 ;
  assign n1988 = ~x275 & x307 ;
  assign n1989 = x275 & ~x307 ;
  assign n1990 = ~x274 & x306 ;
  assign n1991 = x274 & ~x306 ;
  assign n1992 = ~x273 & x305 ;
  assign n1993 = x273 & ~x305 ;
  assign n1994 = ~x272 & x304 ;
  assign n1995 = x272 & ~x304 ;
  assign n1996 = ~x271 & x303 ;
  assign n1997 = x271 & ~x303 ;
  assign n1998 = ~x270 & x302 ;
  assign n1999 = x270 & ~x302 ;
  assign n2000 = ~x269 & x301 ;
  assign n2001 = x269 & ~x301 ;
  assign n2002 = ~x268 & x300 ;
  assign n2003 = x268 & ~x300 ;
  assign n2004 = ~x267 & x299 ;
  assign n2005 = x267 & ~x299 ;
  assign n2006 = ~x266 & x298 ;
  assign n2007 = x266 & ~x298 ;
  assign n2008 = ~x265 & x297 ;
  assign n2009 = x265 & ~x297 ;
  assign n2010 = ~x264 & x296 ;
  assign n2011 = x264 & ~x296 ;
  assign n2012 = ~x263 & x295 ;
  assign n2013 = x263 & ~x295 ;
  assign n2014 = ~x262 & x294 ;
  assign n2015 = x262 & ~x294 ;
  assign n2016 = ~x261 & x293 ;
  assign n2017 = x261 & ~x293 ;
  assign n2018 = ~x260 & x292 ;
  assign n2019 = x260 & ~x292 ;
  assign n2020 = ~x259 & x291 ;
  assign n2021 = x259 & ~x291 ;
  assign n2022 = ~x258 & x290 ;
  assign n2023 = x258 & ~x290 ;
  assign n2024 = ~x257 & x289 ;
  assign n2025 = x257 & ~x289 ;
  assign n2026 = x256 & ~x288 ;
  assign n2027 = ~n2025 & ~n2026 ;
  assign n2028 = ~n2024 & ~n2027 ;
  assign n2029 = ~n2023 & ~n2028 ;
  assign n2030 = ~n2022 & ~n2029 ;
  assign n2031 = ~n2021 & ~n2030 ;
  assign n2032 = ~n2020 & ~n2031 ;
  assign n2033 = ~n2019 & ~n2032 ;
  assign n2034 = ~n2018 & ~n2033 ;
  assign n2035 = ~n2017 & ~n2034 ;
  assign n2036 = ~n2016 & ~n2035 ;
  assign n2037 = ~n2015 & ~n2036 ;
  assign n2038 = ~n2014 & ~n2037 ;
  assign n2039 = ~n2013 & ~n2038 ;
  assign n2040 = ~n2012 & ~n2039 ;
  assign n2041 = ~n2011 & ~n2040 ;
  assign n2042 = ~n2010 & ~n2041 ;
  assign n2043 = ~n2009 & ~n2042 ;
  assign n2044 = ~n2008 & ~n2043 ;
  assign n2045 = ~n2007 & ~n2044 ;
  assign n2046 = ~n2006 & ~n2045 ;
  assign n2047 = ~n2005 & ~n2046 ;
  assign n2048 = ~n2004 & ~n2047 ;
  assign n2049 = ~n2003 & ~n2048 ;
  assign n2050 = ~n2002 & ~n2049 ;
  assign n2051 = ~n2001 & ~n2050 ;
  assign n2052 = ~n2000 & ~n2051 ;
  assign n2053 = ~n1999 & ~n2052 ;
  assign n2054 = ~n1998 & ~n2053 ;
  assign n2055 = ~n1997 & ~n2054 ;
  assign n2056 = ~n1996 & ~n2055 ;
  assign n2057 = ~n1995 & ~n2056 ;
  assign n2058 = ~n1994 & ~n2057 ;
  assign n2059 = ~n1993 & ~n2058 ;
  assign n2060 = ~n1992 & ~n2059 ;
  assign n2061 = ~n1991 & ~n2060 ;
  assign n2062 = ~n1990 & ~n2061 ;
  assign n2063 = ~n1989 & ~n2062 ;
  assign n2064 = ~n1988 & ~n2063 ;
  assign n2065 = ~n1987 & ~n2064 ;
  assign n2066 = ~n1986 & ~n2065 ;
  assign n2067 = ~n1985 & ~n2066 ;
  assign n2068 = ~n1984 & ~n2067 ;
  assign n2069 = ~n1983 & ~n2068 ;
  assign n2070 = ~n1982 & ~n2069 ;
  assign n2071 = ~n1981 & ~n2070 ;
  assign n2072 = ~n1980 & ~n2071 ;
  assign n2073 = ~n1979 & ~n2072 ;
  assign n2074 = ~n1978 & ~n2073 ;
  assign n2075 = ~n1977 & ~n2074 ;
  assign n2076 = ~n1976 & ~n2075 ;
  assign n2077 = ~n1975 & ~n2076 ;
  assign n2078 = ~n1974 & ~n2077 ;
  assign n2079 = ~n1973 & ~n2078 ;
  assign n2080 = ~n1972 & ~n2079 ;
  assign n2081 = ~n1971 & ~n2080 ;
  assign n2082 = ~n1970 & ~n2081 ;
  assign n2083 = ~n1969 & ~n2082 ;
  assign n2084 = ~n1968 & ~n2083 ;
  assign n2085 = ~n1967 & ~n2084 ;
  assign n2086 = ~n1966 & ~n2085 ;
  assign n2087 = ~n1965 & ~n2086 ;
  assign n2088 = ~n1964 & ~n2087 ;
  assign n2089 = x315 & ~n2088 ;
  assign n2090 = x283 & n2088 ;
  assign n2091 = ~n2089 & ~n2090 ;
  assign n2092 = n513 & ~n514 ;
  assign n2093 = ~n513 & n514 ;
  assign n2094 = x289 & ~n2088 ;
  assign n2095 = x257 & n2088 ;
  assign n2096 = ~n2094 & ~n2095 ;
  assign n2097 = ~x351 & x383 ;
  assign n2098 = x351 & ~x383 ;
  assign n2099 = ~x350 & x382 ;
  assign n2100 = x350 & ~x382 ;
  assign n2101 = ~x349 & x381 ;
  assign n2102 = x349 & ~x381 ;
  assign n2103 = ~x348 & x380 ;
  assign n2104 = x348 & ~x380 ;
  assign n2105 = ~x347 & x379 ;
  assign n2106 = x347 & ~x379 ;
  assign n2107 = ~x346 & x378 ;
  assign n2108 = x346 & ~x378 ;
  assign n2109 = ~x345 & x377 ;
  assign n2110 = x345 & ~x377 ;
  assign n2111 = ~x344 & x376 ;
  assign n2112 = x344 & ~x376 ;
  assign n2113 = ~x343 & x375 ;
  assign n2114 = x343 & ~x375 ;
  assign n2115 = ~x342 & x374 ;
  assign n2116 = x342 & ~x374 ;
  assign n2117 = ~x341 & x373 ;
  assign n2118 = x341 & ~x373 ;
  assign n2119 = ~x340 & x372 ;
  assign n2120 = x340 & ~x372 ;
  assign n2121 = ~x339 & x371 ;
  assign n2122 = x339 & ~x371 ;
  assign n2123 = ~x338 & x370 ;
  assign n2124 = x338 & ~x370 ;
  assign n2125 = ~x337 & x369 ;
  assign n2126 = x337 & ~x369 ;
  assign n2127 = ~x336 & x368 ;
  assign n2128 = x336 & ~x368 ;
  assign n2129 = ~x335 & x367 ;
  assign n2130 = x335 & ~x367 ;
  assign n2131 = ~x334 & x366 ;
  assign n2132 = x334 & ~x366 ;
  assign n2133 = ~x333 & x365 ;
  assign n2134 = x333 & ~x365 ;
  assign n2135 = ~x332 & x364 ;
  assign n2136 = x332 & ~x364 ;
  assign n2137 = ~x331 & x363 ;
  assign n2138 = x331 & ~x363 ;
  assign n2139 = ~x330 & x362 ;
  assign n2140 = x330 & ~x362 ;
  assign n2141 = ~x329 & x361 ;
  assign n2142 = x329 & ~x361 ;
  assign n2143 = ~x328 & x360 ;
  assign n2144 = x328 & ~x360 ;
  assign n2145 = ~x327 & x359 ;
  assign n2146 = x327 & ~x359 ;
  assign n2147 = ~x326 & x358 ;
  assign n2148 = x326 & ~x358 ;
  assign n2149 = ~x325 & x357 ;
  assign n2150 = x325 & ~x357 ;
  assign n2151 = ~x324 & x356 ;
  assign n2152 = x324 & ~x356 ;
  assign n2153 = ~x323 & x355 ;
  assign n2154 = x323 & ~x355 ;
  assign n2155 = ~x322 & x354 ;
  assign n2156 = x322 & ~x354 ;
  assign n2157 = ~x321 & x353 ;
  assign n2158 = x321 & ~x353 ;
  assign n2159 = x320 & ~x352 ;
  assign n2160 = ~n2158 & ~n2159 ;
  assign n2161 = ~n2157 & ~n2160 ;
  assign n2162 = ~n2156 & ~n2161 ;
  assign n2163 = ~n2155 & ~n2162 ;
  assign n2164 = ~n2154 & ~n2163 ;
  assign n2165 = ~n2153 & ~n2164 ;
  assign n2166 = ~n2152 & ~n2165 ;
  assign n2167 = ~n2151 & ~n2166 ;
  assign n2168 = ~n2150 & ~n2167 ;
  assign n2169 = ~n2149 & ~n2168 ;
  assign n2170 = ~n2148 & ~n2169 ;
  assign n2171 = ~n2147 & ~n2170 ;
  assign n2172 = ~n2146 & ~n2171 ;
  assign n2173 = ~n2145 & ~n2172 ;
  assign n2174 = ~n2144 & ~n2173 ;
  assign n2175 = ~n2143 & ~n2174 ;
  assign n2176 = ~n2142 & ~n2175 ;
  assign n2177 = ~n2141 & ~n2176 ;
  assign n2178 = ~n2140 & ~n2177 ;
  assign n2179 = ~n2139 & ~n2178 ;
  assign n2180 = ~n2138 & ~n2179 ;
  assign n2181 = ~n2137 & ~n2180 ;
  assign n2182 = ~n2136 & ~n2181 ;
  assign n2183 = ~n2135 & ~n2182 ;
  assign n2184 = ~n2134 & ~n2183 ;
  assign n2185 = ~n2133 & ~n2184 ;
  assign n2186 = ~n2132 & ~n2185 ;
  assign n2187 = ~n2131 & ~n2186 ;
  assign n2188 = ~n2130 & ~n2187 ;
  assign n2189 = ~n2129 & ~n2188 ;
  assign n2190 = ~n2128 & ~n2189 ;
  assign n2191 = ~n2127 & ~n2190 ;
  assign n2192 = ~n2126 & ~n2191 ;
  assign n2193 = ~n2125 & ~n2192 ;
  assign n2194 = ~n2124 & ~n2193 ;
  assign n2195 = ~n2123 & ~n2194 ;
  assign n2196 = ~n2122 & ~n2195 ;
  assign n2197 = ~n2121 & ~n2196 ;
  assign n2198 = ~n2120 & ~n2197 ;
  assign n2199 = ~n2119 & ~n2198 ;
  assign n2200 = ~n2118 & ~n2199 ;
  assign n2201 = ~n2117 & ~n2200 ;
  assign n2202 = ~n2116 & ~n2201 ;
  assign n2203 = ~n2115 & ~n2202 ;
  assign n2204 = ~n2114 & ~n2203 ;
  assign n2205 = ~n2113 & ~n2204 ;
  assign n2206 = ~n2112 & ~n2205 ;
  assign n2207 = ~n2111 & ~n2206 ;
  assign n2208 = ~n2110 & ~n2207 ;
  assign n2209 = ~n2109 & ~n2208 ;
  assign n2210 = ~n2108 & ~n2209 ;
  assign n2211 = ~n2107 & ~n2210 ;
  assign n2212 = ~n2106 & ~n2211 ;
  assign n2213 = ~n2105 & ~n2212 ;
  assign n2214 = ~n2104 & ~n2213 ;
  assign n2215 = ~n2103 & ~n2214 ;
  assign n2216 = ~n2102 & ~n2215 ;
  assign n2217 = ~n2101 & ~n2216 ;
  assign n2218 = ~n2100 & ~n2217 ;
  assign n2219 = ~n2099 & ~n2218 ;
  assign n2220 = ~n2098 & ~n2219 ;
  assign n2221 = ~n2097 & ~n2220 ;
  assign n2222 = x353 & ~n2221 ;
  assign n2223 = x321 & n2221 ;
  assign n2224 = ~n2222 & ~n2223 ;
  assign n2225 = n2096 & ~n2224 ;
  assign n2226 = x352 & ~n2221 ;
  assign n2227 = x320 & n2221 ;
  assign n2228 = ~n2226 & ~n2227 ;
  assign n2229 = x288 & ~n2088 ;
  assign n2230 = x256 & n2088 ;
  assign n2231 = ~n2229 & ~n2230 ;
  assign n2232 = n2228 & ~n2231 ;
  assign n2233 = ~n2225 & n2232 ;
  assign n2234 = x354 & ~n2221 ;
  assign n2235 = x322 & n2221 ;
  assign n2236 = ~n2234 & ~n2235 ;
  assign n2237 = x290 & ~n2088 ;
  assign n2238 = x258 & n2088 ;
  assign n2239 = ~n2237 & ~n2238 ;
  assign n2240 = n2236 & ~n2239 ;
  assign n2241 = ~n2096 & n2224 ;
  assign n2242 = ~n2240 & ~n2241 ;
  assign n2243 = ~n2233 & n2242 ;
  assign n2244 = x291 & ~n2088 ;
  assign n2245 = x259 & n2088 ;
  assign n2246 = ~n2244 & ~n2245 ;
  assign n2247 = x355 & ~n2221 ;
  assign n2248 = x323 & n2221 ;
  assign n2249 = ~n2247 & ~n2248 ;
  assign n2250 = n2246 & ~n2249 ;
  assign n2251 = ~n2236 & n2239 ;
  assign n2252 = ~n2250 & ~n2251 ;
  assign n2253 = ~n2243 & n2252 ;
  assign n2254 = ~n2246 & n2249 ;
  assign n2255 = x356 & ~n2221 ;
  assign n2256 = x324 & n2221 ;
  assign n2257 = ~n2255 & ~n2256 ;
  assign n2258 = x292 & ~n2088 ;
  assign n2259 = x260 & n2088 ;
  assign n2260 = ~n2258 & ~n2259 ;
  assign n2261 = n2257 & ~n2260 ;
  assign n2262 = ~n2254 & ~n2261 ;
  assign n2263 = ~n2253 & n2262 ;
  assign n2264 = x357 & ~n2221 ;
  assign n2265 = x325 & n2221 ;
  assign n2266 = ~n2264 & ~n2265 ;
  assign n2267 = x293 & ~n2088 ;
  assign n2268 = x261 & n2088 ;
  assign n2269 = ~n2267 & ~n2268 ;
  assign n2270 = ~n2266 & n2269 ;
  assign n2271 = ~n2257 & n2260 ;
  assign n2272 = ~n2270 & ~n2271 ;
  assign n2273 = ~n2263 & n2272 ;
  assign n2274 = x358 & ~n2221 ;
  assign n2275 = x326 & n2221 ;
  assign n2276 = ~n2274 & ~n2275 ;
  assign n2277 = x294 & ~n2088 ;
  assign n2278 = x262 & n2088 ;
  assign n2279 = ~n2277 & ~n2278 ;
  assign n2280 = n2276 & ~n2279 ;
  assign n2281 = n2266 & ~n2269 ;
  assign n2282 = ~n2280 & ~n2281 ;
  assign n2283 = ~n2273 & n2282 ;
  assign n2284 = x295 & ~n2088 ;
  assign n2285 = x263 & n2088 ;
  assign n2286 = ~n2284 & ~n2285 ;
  assign n2287 = x359 & ~n2221 ;
  assign n2288 = x327 & n2221 ;
  assign n2289 = ~n2287 & ~n2288 ;
  assign n2290 = n2286 & ~n2289 ;
  assign n2291 = ~n2276 & n2279 ;
  assign n2292 = ~n2290 & ~n2291 ;
  assign n2293 = ~n2283 & n2292 ;
  assign n2294 = ~n2286 & n2289 ;
  assign n2295 = x360 & ~n2221 ;
  assign n2296 = x328 & n2221 ;
  assign n2297 = ~n2295 & ~n2296 ;
  assign n2298 = x296 & ~n2088 ;
  assign n2299 = x264 & n2088 ;
  assign n2300 = ~n2298 & ~n2299 ;
  assign n2301 = n2297 & ~n2300 ;
  assign n2302 = ~n2294 & ~n2301 ;
  assign n2303 = ~n2293 & n2302 ;
  assign n2304 = ~n2297 & n2300 ;
  assign n2305 = x361 & ~n2221 ;
  assign n2306 = x329 & n2221 ;
  assign n2307 = ~n2305 & ~n2306 ;
  assign n2308 = x297 & ~n2088 ;
  assign n2309 = x265 & n2088 ;
  assign n2310 = ~n2308 & ~n2309 ;
  assign n2311 = ~n2307 & n2310 ;
  assign n2312 = ~n2304 & ~n2311 ;
  assign n2313 = ~n2303 & n2312 ;
  assign n2314 = n2307 & ~n2310 ;
  assign n2315 = x298 & ~n2088 ;
  assign n2316 = x266 & n2088 ;
  assign n2317 = ~n2315 & ~n2316 ;
  assign n2318 = x362 & ~n2221 ;
  assign n2319 = x330 & n2221 ;
  assign n2320 = ~n2318 & ~n2319 ;
  assign n2321 = ~n2317 & n2320 ;
  assign n2322 = ~n2314 & ~n2321 ;
  assign n2323 = ~n2313 & n2322 ;
  assign n2324 = x299 & ~n2088 ;
  assign n2325 = x267 & n2088 ;
  assign n2326 = ~n2324 & ~n2325 ;
  assign n2327 = x363 & ~n2221 ;
  assign n2328 = x331 & n2221 ;
  assign n2329 = ~n2327 & ~n2328 ;
  assign n2330 = n2326 & ~n2329 ;
  assign n2331 = n2317 & ~n2320 ;
  assign n2332 = ~n2330 & ~n2331 ;
  assign n2333 = ~n2323 & n2332 ;
  assign n2334 = x364 & ~n2221 ;
  assign n2335 = x332 & n2221 ;
  assign n2336 = ~n2334 & ~n2335 ;
  assign n2337 = x300 & ~n2088 ;
  assign n2338 = x268 & n2088 ;
  assign n2339 = ~n2337 & ~n2338 ;
  assign n2340 = n2336 & ~n2339 ;
  assign n2341 = ~n2326 & n2329 ;
  assign n2342 = ~n2340 & ~n2341 ;
  assign n2343 = ~n2333 & n2342 ;
  assign n2344 = ~n2336 & n2339 ;
  assign n2345 = x365 & ~n2221 ;
  assign n2346 = x333 & n2221 ;
  assign n2347 = ~n2345 & ~n2346 ;
  assign n2348 = x301 & ~n2088 ;
  assign n2349 = x269 & n2088 ;
  assign n2350 = ~n2348 & ~n2349 ;
  assign n2351 = ~n2347 & n2350 ;
  assign n2352 = ~n2344 & ~n2351 ;
  assign n2353 = ~n2343 & n2352 ;
  assign n2354 = n2347 & ~n2350 ;
  assign n2355 = x302 & ~n2088 ;
  assign n2356 = x270 & n2088 ;
  assign n2357 = ~n2355 & ~n2356 ;
  assign n2358 = x366 & ~n2221 ;
  assign n2359 = x334 & n2221 ;
  assign n2360 = ~n2358 & ~n2359 ;
  assign n2361 = ~n2357 & n2360 ;
  assign n2362 = ~n2354 & ~n2361 ;
  assign n2363 = ~n2353 & n2362 ;
  assign n2364 = x303 & ~n2088 ;
  assign n2365 = x271 & n2088 ;
  assign n2366 = ~n2364 & ~n2365 ;
  assign n2367 = x367 & ~n2221 ;
  assign n2368 = x335 & n2221 ;
  assign n2369 = ~n2367 & ~n2368 ;
  assign n2370 = n2366 & ~n2369 ;
  assign n2371 = n2357 & ~n2360 ;
  assign n2372 = ~n2370 & ~n2371 ;
  assign n2373 = ~n2363 & n2372 ;
  assign n2374 = x368 & ~n2221 ;
  assign n2375 = x336 & n2221 ;
  assign n2376 = ~n2374 & ~n2375 ;
  assign n2377 = x304 & ~n2088 ;
  assign n2378 = x272 & n2088 ;
  assign n2379 = ~n2377 & ~n2378 ;
  assign n2380 = n2376 & ~n2379 ;
  assign n2381 = ~n2366 & n2369 ;
  assign n2382 = ~n2380 & ~n2381 ;
  assign n2383 = ~n2373 & n2382 ;
  assign n2384 = ~n2376 & n2379 ;
  assign n2385 = x369 & ~n2221 ;
  assign n2386 = x337 & n2221 ;
  assign n2387 = ~n2385 & ~n2386 ;
  assign n2388 = x305 & ~n2088 ;
  assign n2389 = x273 & n2088 ;
  assign n2390 = ~n2388 & ~n2389 ;
  assign n2391 = ~n2387 & n2390 ;
  assign n2392 = ~n2384 & ~n2391 ;
  assign n2393 = ~n2383 & n2392 ;
  assign n2394 = n2387 & ~n2390 ;
  assign n2395 = x306 & ~n2088 ;
  assign n2396 = x274 & n2088 ;
  assign n2397 = ~n2395 & ~n2396 ;
  assign n2398 = x370 & ~n2221 ;
  assign n2399 = x338 & n2221 ;
  assign n2400 = ~n2398 & ~n2399 ;
  assign n2401 = ~n2397 & n2400 ;
  assign n2402 = ~n2394 & ~n2401 ;
  assign n2403 = ~n2393 & n2402 ;
  assign n2404 = x307 & ~n2088 ;
  assign n2405 = x275 & n2088 ;
  assign n2406 = ~n2404 & ~n2405 ;
  assign n2407 = x371 & ~n2221 ;
  assign n2408 = x339 & n2221 ;
  assign n2409 = ~n2407 & ~n2408 ;
  assign n2410 = n2406 & ~n2409 ;
  assign n2411 = n2397 & ~n2400 ;
  assign n2412 = ~n2410 & ~n2411 ;
  assign n2413 = ~n2403 & n2412 ;
  assign n2414 = x372 & ~n2221 ;
  assign n2415 = x340 & n2221 ;
  assign n2416 = ~n2414 & ~n2415 ;
  assign n2417 = x308 & ~n2088 ;
  assign n2418 = x276 & n2088 ;
  assign n2419 = ~n2417 & ~n2418 ;
  assign n2420 = n2416 & ~n2419 ;
  assign n2421 = ~n2406 & n2409 ;
  assign n2422 = ~n2420 & ~n2421 ;
  assign n2423 = ~n2413 & n2422 ;
  assign n2424 = ~n2416 & n2419 ;
  assign n2425 = x373 & ~n2221 ;
  assign n2426 = x341 & n2221 ;
  assign n2427 = ~n2425 & ~n2426 ;
  assign n2428 = x309 & ~n2088 ;
  assign n2429 = x277 & n2088 ;
  assign n2430 = ~n2428 & ~n2429 ;
  assign n2431 = ~n2427 & n2430 ;
  assign n2432 = ~n2424 & ~n2431 ;
  assign n2433 = ~n2423 & n2432 ;
  assign n2434 = n2427 & ~n2430 ;
  assign n2435 = x310 & ~n2088 ;
  assign n2436 = x278 & n2088 ;
  assign n2437 = ~n2435 & ~n2436 ;
  assign n2438 = x374 & ~n2221 ;
  assign n2439 = x342 & n2221 ;
  assign n2440 = ~n2438 & ~n2439 ;
  assign n2441 = ~n2437 & n2440 ;
  assign n2442 = ~n2434 & ~n2441 ;
  assign n2443 = ~n2433 & n2442 ;
  assign n2444 = x311 & ~n2088 ;
  assign n2445 = x279 & n2088 ;
  assign n2446 = ~n2444 & ~n2445 ;
  assign n2447 = x375 & ~n2221 ;
  assign n2448 = x343 & n2221 ;
  assign n2449 = ~n2447 & ~n2448 ;
  assign n2450 = n2446 & ~n2449 ;
  assign n2451 = n2437 & ~n2440 ;
  assign n2452 = ~n2450 & ~n2451 ;
  assign n2453 = ~n2443 & n2452 ;
  assign n2454 = x376 & ~n2221 ;
  assign n2455 = x344 & n2221 ;
  assign n2456 = ~n2454 & ~n2455 ;
  assign n2457 = x312 & ~n2088 ;
  assign n2458 = x280 & n2088 ;
  assign n2459 = ~n2457 & ~n2458 ;
  assign n2460 = n2456 & ~n2459 ;
  assign n2461 = ~n2446 & n2449 ;
  assign n2462 = ~n2460 & ~n2461 ;
  assign n2463 = ~n2453 & n2462 ;
  assign n2464 = ~n2456 & n2459 ;
  assign n2465 = x377 & ~n2221 ;
  assign n2466 = x345 & n2221 ;
  assign n2467 = ~n2465 & ~n2466 ;
  assign n2468 = x313 & ~n2088 ;
  assign n2469 = x281 & n2088 ;
  assign n2470 = ~n2468 & ~n2469 ;
  assign n2471 = ~n2467 & n2470 ;
  assign n2472 = ~n2464 & ~n2471 ;
  assign n2473 = ~n2463 & n2472 ;
  assign n2474 = n2467 & ~n2470 ;
  assign n2475 = x314 & ~n2088 ;
  assign n2476 = x282 & n2088 ;
  assign n2477 = ~n2475 & ~n2476 ;
  assign n2478 = x378 & ~n2221 ;
  assign n2479 = x346 & n2221 ;
  assign n2480 = ~n2478 & ~n2479 ;
  assign n2481 = ~n2477 & n2480 ;
  assign n2482 = ~n2474 & ~n2481 ;
  assign n2483 = ~n2473 & n2482 ;
  assign n2484 = x379 & ~n2221 ;
  assign n2485 = x347 & n2221 ;
  assign n2486 = ~n2484 & ~n2485 ;
  assign n2487 = n2091 & ~n2486 ;
  assign n2488 = n2477 & ~n2480 ;
  assign n2489 = ~n2487 & ~n2488 ;
  assign n2490 = ~n2483 & n2489 ;
  assign n2491 = x380 & ~n2221 ;
  assign n2492 = x348 & n2221 ;
  assign n2493 = ~n2491 & ~n2492 ;
  assign n2494 = x316 & ~n2088 ;
  assign n2495 = x284 & n2088 ;
  assign n2496 = ~n2494 & ~n2495 ;
  assign n2497 = n2493 & ~n2496 ;
  assign n2498 = ~n2091 & n2486 ;
  assign n2499 = ~n2497 & ~n2498 ;
  assign n2500 = ~n2490 & n2499 ;
  assign n2501 = ~n2493 & n2496 ;
  assign n2502 = x381 & ~n2221 ;
  assign n2503 = x349 & n2221 ;
  assign n2504 = ~n2502 & ~n2503 ;
  assign n2505 = x317 & ~n2088 ;
  assign n2506 = x285 & n2088 ;
  assign n2507 = ~n2505 & ~n2506 ;
  assign n2508 = ~n2504 & n2507 ;
  assign n2509 = ~n2501 & ~n2508 ;
  assign n2510 = ~n2500 & n2509 ;
  assign n2511 = n2504 & ~n2507 ;
  assign n2512 = x318 & ~n2088 ;
  assign n2513 = x286 & n2088 ;
  assign n2514 = ~n2512 & ~n2513 ;
  assign n2515 = x382 & ~n2221 ;
  assign n2516 = x350 & n2221 ;
  assign n2517 = ~n2515 & ~n2516 ;
  assign n2518 = ~n2514 & n2517 ;
  assign n2519 = ~n2511 & ~n2518 ;
  assign n2520 = ~n2510 & n2519 ;
  assign n2521 = n2514 & ~n2517 ;
  assign n2522 = ~n2520 & ~n2521 ;
  assign n2523 = ~n2093 & ~n2522 ;
  assign n2524 = ~n2092 & ~n2523 ;
  assign n2525 = ~n2091 & n2524 ;
  assign n2526 = ~n2486 & ~n2524 ;
  assign n2527 = ~n2525 & ~n2526 ;
  assign n2528 = ~n515 & n518 ;
  assign n2529 = ~n2096 & n2524 ;
  assign n2530 = ~n2224 & ~n2524 ;
  assign n2531 = ~n2529 & ~n2530 ;
  assign n2532 = ~x415 & x447 ;
  assign n2533 = x415 & ~x447 ;
  assign n2534 = ~x414 & x446 ;
  assign n2535 = x414 & ~x446 ;
  assign n2536 = ~x413 & x445 ;
  assign n2537 = x413 & ~x445 ;
  assign n2538 = ~x412 & x444 ;
  assign n2539 = x412 & ~x444 ;
  assign n2540 = ~x411 & x443 ;
  assign n2541 = x411 & ~x443 ;
  assign n2542 = ~x410 & x442 ;
  assign n2543 = x410 & ~x442 ;
  assign n2544 = ~x409 & x441 ;
  assign n2545 = x409 & ~x441 ;
  assign n2546 = ~x408 & x440 ;
  assign n2547 = x408 & ~x440 ;
  assign n2548 = ~x407 & x439 ;
  assign n2549 = x407 & ~x439 ;
  assign n2550 = ~x406 & x438 ;
  assign n2551 = x406 & ~x438 ;
  assign n2552 = ~x405 & x437 ;
  assign n2553 = x405 & ~x437 ;
  assign n2554 = ~x404 & x436 ;
  assign n2555 = x404 & ~x436 ;
  assign n2556 = ~x403 & x435 ;
  assign n2557 = x403 & ~x435 ;
  assign n2558 = ~x402 & x434 ;
  assign n2559 = x402 & ~x434 ;
  assign n2560 = ~x401 & x433 ;
  assign n2561 = x401 & ~x433 ;
  assign n2562 = ~x400 & x432 ;
  assign n2563 = x400 & ~x432 ;
  assign n2564 = ~x399 & x431 ;
  assign n2565 = x399 & ~x431 ;
  assign n2566 = ~x398 & x430 ;
  assign n2567 = x398 & ~x430 ;
  assign n2568 = ~x397 & x429 ;
  assign n2569 = x397 & ~x429 ;
  assign n2570 = ~x396 & x428 ;
  assign n2571 = x396 & ~x428 ;
  assign n2572 = ~x395 & x427 ;
  assign n2573 = x395 & ~x427 ;
  assign n2574 = ~x394 & x426 ;
  assign n2575 = x394 & ~x426 ;
  assign n2576 = ~x393 & x425 ;
  assign n2577 = x393 & ~x425 ;
  assign n2578 = ~x392 & x424 ;
  assign n2579 = x392 & ~x424 ;
  assign n2580 = ~x391 & x423 ;
  assign n2581 = x391 & ~x423 ;
  assign n2582 = ~x390 & x422 ;
  assign n2583 = x390 & ~x422 ;
  assign n2584 = ~x389 & x421 ;
  assign n2585 = x389 & ~x421 ;
  assign n2586 = ~x388 & x420 ;
  assign n2587 = x388 & ~x420 ;
  assign n2588 = ~x387 & x419 ;
  assign n2589 = x387 & ~x419 ;
  assign n2590 = ~x386 & x418 ;
  assign n2591 = x386 & ~x418 ;
  assign n2592 = ~x385 & x417 ;
  assign n2593 = x385 & ~x417 ;
  assign n2594 = x384 & ~x416 ;
  assign n2595 = ~n2593 & ~n2594 ;
  assign n2596 = ~n2592 & ~n2595 ;
  assign n2597 = ~n2591 & ~n2596 ;
  assign n2598 = ~n2590 & ~n2597 ;
  assign n2599 = ~n2589 & ~n2598 ;
  assign n2600 = ~n2588 & ~n2599 ;
  assign n2601 = ~n2587 & ~n2600 ;
  assign n2602 = ~n2586 & ~n2601 ;
  assign n2603 = ~n2585 & ~n2602 ;
  assign n2604 = ~n2584 & ~n2603 ;
  assign n2605 = ~n2583 & ~n2604 ;
  assign n2606 = ~n2582 & ~n2605 ;
  assign n2607 = ~n2581 & ~n2606 ;
  assign n2608 = ~n2580 & ~n2607 ;
  assign n2609 = ~n2579 & ~n2608 ;
  assign n2610 = ~n2578 & ~n2609 ;
  assign n2611 = ~n2577 & ~n2610 ;
  assign n2612 = ~n2576 & ~n2611 ;
  assign n2613 = ~n2575 & ~n2612 ;
  assign n2614 = ~n2574 & ~n2613 ;
  assign n2615 = ~n2573 & ~n2614 ;
  assign n2616 = ~n2572 & ~n2615 ;
  assign n2617 = ~n2571 & ~n2616 ;
  assign n2618 = ~n2570 & ~n2617 ;
  assign n2619 = ~n2569 & ~n2618 ;
  assign n2620 = ~n2568 & ~n2619 ;
  assign n2621 = ~n2567 & ~n2620 ;
  assign n2622 = ~n2566 & ~n2621 ;
  assign n2623 = ~n2565 & ~n2622 ;
  assign n2624 = ~n2564 & ~n2623 ;
  assign n2625 = ~n2563 & ~n2624 ;
  assign n2626 = ~n2562 & ~n2625 ;
  assign n2627 = ~n2561 & ~n2626 ;
  assign n2628 = ~n2560 & ~n2627 ;
  assign n2629 = ~n2559 & ~n2628 ;
  assign n2630 = ~n2558 & ~n2629 ;
  assign n2631 = ~n2557 & ~n2630 ;
  assign n2632 = ~n2556 & ~n2631 ;
  assign n2633 = ~n2555 & ~n2632 ;
  assign n2634 = ~n2554 & ~n2633 ;
  assign n2635 = ~n2553 & ~n2634 ;
  assign n2636 = ~n2552 & ~n2635 ;
  assign n2637 = ~n2551 & ~n2636 ;
  assign n2638 = ~n2550 & ~n2637 ;
  assign n2639 = ~n2549 & ~n2638 ;
  assign n2640 = ~n2548 & ~n2639 ;
  assign n2641 = ~n2547 & ~n2640 ;
  assign n2642 = ~n2546 & ~n2641 ;
  assign n2643 = ~n2545 & ~n2642 ;
  assign n2644 = ~n2544 & ~n2643 ;
  assign n2645 = ~n2543 & ~n2644 ;
  assign n2646 = ~n2542 & ~n2645 ;
  assign n2647 = ~n2541 & ~n2646 ;
  assign n2648 = ~n2540 & ~n2647 ;
  assign n2649 = ~n2539 & ~n2648 ;
  assign n2650 = ~n2538 & ~n2649 ;
  assign n2651 = ~n2537 & ~n2650 ;
  assign n2652 = ~n2536 & ~n2651 ;
  assign n2653 = ~n2535 & ~n2652 ;
  assign n2654 = ~n2534 & ~n2653 ;
  assign n2655 = ~n2533 & ~n2654 ;
  assign n2656 = ~n2532 & ~n2655 ;
  assign n2657 = x417 & ~n2656 ;
  assign n2658 = x385 & n2656 ;
  assign n2659 = ~n2657 & ~n2658 ;
  assign n2660 = n516 & ~n517 ;
  assign n2661 = ~n516 & n517 ;
  assign n2662 = ~x479 & x511 ;
  assign n2663 = x479 & ~x511 ;
  assign n2664 = ~x478 & x510 ;
  assign n2665 = x478 & ~x510 ;
  assign n2666 = ~x477 & x509 ;
  assign n2667 = x477 & ~x509 ;
  assign n2668 = ~x476 & x508 ;
  assign n2669 = x476 & ~x508 ;
  assign n2670 = ~x475 & x507 ;
  assign n2671 = x475 & ~x507 ;
  assign n2672 = ~x474 & x506 ;
  assign n2673 = x474 & ~x506 ;
  assign n2674 = ~x473 & x505 ;
  assign n2675 = x473 & ~x505 ;
  assign n2676 = ~x472 & x504 ;
  assign n2677 = x472 & ~x504 ;
  assign n2678 = ~x471 & x503 ;
  assign n2679 = x471 & ~x503 ;
  assign n2680 = ~x470 & x502 ;
  assign n2681 = x470 & ~x502 ;
  assign n2682 = ~x469 & x501 ;
  assign n2683 = x469 & ~x501 ;
  assign n2684 = ~x468 & x500 ;
  assign n2685 = x468 & ~x500 ;
  assign n2686 = ~x467 & x499 ;
  assign n2687 = x467 & ~x499 ;
  assign n2688 = ~x466 & x498 ;
  assign n2689 = x466 & ~x498 ;
  assign n2690 = ~x465 & x497 ;
  assign n2691 = x465 & ~x497 ;
  assign n2692 = ~x464 & x496 ;
  assign n2693 = x464 & ~x496 ;
  assign n2694 = ~x463 & x495 ;
  assign n2695 = x463 & ~x495 ;
  assign n2696 = ~x462 & x494 ;
  assign n2697 = x462 & ~x494 ;
  assign n2698 = ~x461 & x493 ;
  assign n2699 = x461 & ~x493 ;
  assign n2700 = ~x460 & x492 ;
  assign n2701 = x460 & ~x492 ;
  assign n2702 = ~x459 & x491 ;
  assign n2703 = x459 & ~x491 ;
  assign n2704 = ~x458 & x490 ;
  assign n2705 = x458 & ~x490 ;
  assign n2706 = ~x457 & x489 ;
  assign n2707 = x457 & ~x489 ;
  assign n2708 = ~x456 & x488 ;
  assign n2709 = x456 & ~x488 ;
  assign n2710 = ~x455 & x487 ;
  assign n2711 = x455 & ~x487 ;
  assign n2712 = ~x454 & x486 ;
  assign n2713 = x454 & ~x486 ;
  assign n2714 = ~x453 & x485 ;
  assign n2715 = x453 & ~x485 ;
  assign n2716 = ~x452 & x484 ;
  assign n2717 = x452 & ~x484 ;
  assign n2718 = ~x451 & x483 ;
  assign n2719 = x451 & ~x483 ;
  assign n2720 = ~x450 & x482 ;
  assign n2721 = x450 & ~x482 ;
  assign n2722 = ~x449 & x481 ;
  assign n2723 = x449 & ~x481 ;
  assign n2724 = x448 & ~x480 ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = ~n2722 & ~n2725 ;
  assign n2727 = ~n2721 & ~n2726 ;
  assign n2728 = ~n2720 & ~n2727 ;
  assign n2729 = ~n2719 & ~n2728 ;
  assign n2730 = ~n2718 & ~n2729 ;
  assign n2731 = ~n2717 & ~n2730 ;
  assign n2732 = ~n2716 & ~n2731 ;
  assign n2733 = ~n2715 & ~n2732 ;
  assign n2734 = ~n2714 & ~n2733 ;
  assign n2735 = ~n2713 & ~n2734 ;
  assign n2736 = ~n2712 & ~n2735 ;
  assign n2737 = ~n2711 & ~n2736 ;
  assign n2738 = ~n2710 & ~n2737 ;
  assign n2739 = ~n2709 & ~n2738 ;
  assign n2740 = ~n2708 & ~n2739 ;
  assign n2741 = ~n2707 & ~n2740 ;
  assign n2742 = ~n2706 & ~n2741 ;
  assign n2743 = ~n2705 & ~n2742 ;
  assign n2744 = ~n2704 & ~n2743 ;
  assign n2745 = ~n2703 & ~n2744 ;
  assign n2746 = ~n2702 & ~n2745 ;
  assign n2747 = ~n2701 & ~n2746 ;
  assign n2748 = ~n2700 & ~n2747 ;
  assign n2749 = ~n2699 & ~n2748 ;
  assign n2750 = ~n2698 & ~n2749 ;
  assign n2751 = ~n2697 & ~n2750 ;
  assign n2752 = ~n2696 & ~n2751 ;
  assign n2753 = ~n2695 & ~n2752 ;
  assign n2754 = ~n2694 & ~n2753 ;
  assign n2755 = ~n2693 & ~n2754 ;
  assign n2756 = ~n2692 & ~n2755 ;
  assign n2757 = ~n2691 & ~n2756 ;
  assign n2758 = ~n2690 & ~n2757 ;
  assign n2759 = ~n2689 & ~n2758 ;
  assign n2760 = ~n2688 & ~n2759 ;
  assign n2761 = ~n2687 & ~n2760 ;
  assign n2762 = ~n2686 & ~n2761 ;
  assign n2763 = ~n2685 & ~n2762 ;
  assign n2764 = ~n2684 & ~n2763 ;
  assign n2765 = ~n2683 & ~n2764 ;
  assign n2766 = ~n2682 & ~n2765 ;
  assign n2767 = ~n2681 & ~n2766 ;
  assign n2768 = ~n2680 & ~n2767 ;
  assign n2769 = ~n2679 & ~n2768 ;
  assign n2770 = ~n2678 & ~n2769 ;
  assign n2771 = ~n2677 & ~n2770 ;
  assign n2772 = ~n2676 & ~n2771 ;
  assign n2773 = ~n2675 & ~n2772 ;
  assign n2774 = ~n2674 & ~n2773 ;
  assign n2775 = ~n2673 & ~n2774 ;
  assign n2776 = ~n2672 & ~n2775 ;
  assign n2777 = ~n2671 & ~n2776 ;
  assign n2778 = ~n2670 & ~n2777 ;
  assign n2779 = ~n2669 & ~n2778 ;
  assign n2780 = ~n2668 & ~n2779 ;
  assign n2781 = ~n2667 & ~n2780 ;
  assign n2782 = ~n2666 & ~n2781 ;
  assign n2783 = ~n2665 & ~n2782 ;
  assign n2784 = ~n2664 & ~n2783 ;
  assign n2785 = ~n2663 & ~n2784 ;
  assign n2786 = ~n2662 & ~n2785 ;
  assign n2787 = x510 & ~n2786 ;
  assign n2788 = x478 & n2786 ;
  assign n2789 = ~n2787 & ~n2788 ;
  assign n2790 = x446 & ~n2656 ;
  assign n2791 = x414 & n2656 ;
  assign n2792 = ~n2790 & ~n2791 ;
  assign n2793 = ~n2789 & n2792 ;
  assign n2794 = x481 & ~n2786 ;
  assign n2795 = x449 & n2786 ;
  assign n2796 = ~n2794 & ~n2795 ;
  assign n2797 = n2659 & ~n2796 ;
  assign n2798 = x480 & ~n2786 ;
  assign n2799 = x448 & n2786 ;
  assign n2800 = ~n2798 & ~n2799 ;
  assign n2801 = x416 & ~n2656 ;
  assign n2802 = x384 & n2656 ;
  assign n2803 = ~n2801 & ~n2802 ;
  assign n2804 = n2800 & ~n2803 ;
  assign n2805 = ~n2797 & n2804 ;
  assign n2806 = x482 & ~n2786 ;
  assign n2807 = x450 & n2786 ;
  assign n2808 = ~n2806 & ~n2807 ;
  assign n2809 = x418 & ~n2656 ;
  assign n2810 = x386 & n2656 ;
  assign n2811 = ~n2809 & ~n2810 ;
  assign n2812 = n2808 & ~n2811 ;
  assign n2813 = ~n2659 & n2796 ;
  assign n2814 = ~n2812 & ~n2813 ;
  assign n2815 = ~n2805 & n2814 ;
  assign n2816 = x419 & ~n2656 ;
  assign n2817 = x387 & n2656 ;
  assign n2818 = ~n2816 & ~n2817 ;
  assign n2819 = x483 & ~n2786 ;
  assign n2820 = x451 & n2786 ;
  assign n2821 = ~n2819 & ~n2820 ;
  assign n2822 = n2818 & ~n2821 ;
  assign n2823 = ~n2808 & n2811 ;
  assign n2824 = ~n2822 & ~n2823 ;
  assign n2825 = ~n2815 & n2824 ;
  assign n2826 = x484 & ~n2786 ;
  assign n2827 = x452 & n2786 ;
  assign n2828 = ~n2826 & ~n2827 ;
  assign n2829 = x420 & ~n2656 ;
  assign n2830 = x388 & n2656 ;
  assign n2831 = ~n2829 & ~n2830 ;
  assign n2832 = n2828 & ~n2831 ;
  assign n2833 = ~n2818 & n2821 ;
  assign n2834 = ~n2832 & ~n2833 ;
  assign n2835 = ~n2825 & n2834 ;
  assign n2836 = ~n2828 & n2831 ;
  assign n2837 = x485 & ~n2786 ;
  assign n2838 = x453 & n2786 ;
  assign n2839 = ~n2837 & ~n2838 ;
  assign n2840 = x421 & ~n2656 ;
  assign n2841 = x389 & n2656 ;
  assign n2842 = ~n2840 & ~n2841 ;
  assign n2843 = ~n2839 & n2842 ;
  assign n2844 = ~n2836 & ~n2843 ;
  assign n2845 = ~n2835 & n2844 ;
  assign n2846 = n2839 & ~n2842 ;
  assign n2847 = x422 & ~n2656 ;
  assign n2848 = x390 & n2656 ;
  assign n2849 = ~n2847 & ~n2848 ;
  assign n2850 = x486 & ~n2786 ;
  assign n2851 = x454 & n2786 ;
  assign n2852 = ~n2850 & ~n2851 ;
  assign n2853 = ~n2849 & n2852 ;
  assign n2854 = ~n2846 & ~n2853 ;
  assign n2855 = ~n2845 & n2854 ;
  assign n2856 = n2849 & ~n2852 ;
  assign n2857 = x423 & ~n2656 ;
  assign n2858 = x391 & n2656 ;
  assign n2859 = ~n2857 & ~n2858 ;
  assign n2860 = x487 & ~n2786 ;
  assign n2861 = x455 & n2786 ;
  assign n2862 = ~n2860 & ~n2861 ;
  assign n2863 = n2859 & ~n2862 ;
  assign n2864 = ~n2856 & ~n2863 ;
  assign n2865 = ~n2855 & n2864 ;
  assign n2866 = x488 & ~n2786 ;
  assign n2867 = x456 & n2786 ;
  assign n2868 = ~n2866 & ~n2867 ;
  assign n2869 = x424 & ~n2656 ;
  assign n2870 = x392 & n2656 ;
  assign n2871 = ~n2869 & ~n2870 ;
  assign n2872 = n2868 & ~n2871 ;
  assign n2873 = ~n2859 & n2862 ;
  assign n2874 = ~n2872 & ~n2873 ;
  assign n2875 = ~n2865 & n2874 ;
  assign n2876 = ~n2868 & n2871 ;
  assign n2877 = x489 & ~n2786 ;
  assign n2878 = x457 & n2786 ;
  assign n2879 = ~n2877 & ~n2878 ;
  assign n2880 = x425 & ~n2656 ;
  assign n2881 = x393 & n2656 ;
  assign n2882 = ~n2880 & ~n2881 ;
  assign n2883 = ~n2879 & n2882 ;
  assign n2884 = ~n2876 & ~n2883 ;
  assign n2885 = ~n2875 & n2884 ;
  assign n2886 = n2879 & ~n2882 ;
  assign n2887 = x426 & ~n2656 ;
  assign n2888 = x394 & n2656 ;
  assign n2889 = ~n2887 & ~n2888 ;
  assign n2890 = x490 & ~n2786 ;
  assign n2891 = x458 & n2786 ;
  assign n2892 = ~n2890 & ~n2891 ;
  assign n2893 = ~n2889 & n2892 ;
  assign n2894 = ~n2886 & ~n2893 ;
  assign n2895 = ~n2885 & n2894 ;
  assign n2896 = x427 & ~n2656 ;
  assign n2897 = x395 & n2656 ;
  assign n2898 = ~n2896 & ~n2897 ;
  assign n2899 = x491 & ~n2786 ;
  assign n2900 = x459 & n2786 ;
  assign n2901 = ~n2899 & ~n2900 ;
  assign n2902 = n2898 & ~n2901 ;
  assign n2903 = n2889 & ~n2892 ;
  assign n2904 = ~n2902 & ~n2903 ;
  assign n2905 = ~n2895 & n2904 ;
  assign n2906 = x492 & ~n2786 ;
  assign n2907 = x460 & n2786 ;
  assign n2908 = ~n2906 & ~n2907 ;
  assign n2909 = x428 & ~n2656 ;
  assign n2910 = x396 & n2656 ;
  assign n2911 = ~n2909 & ~n2910 ;
  assign n2912 = n2908 & ~n2911 ;
  assign n2913 = ~n2898 & n2901 ;
  assign n2914 = ~n2912 & ~n2913 ;
  assign n2915 = ~n2905 & n2914 ;
  assign n2916 = ~n2908 & n2911 ;
  assign n2917 = x493 & ~n2786 ;
  assign n2918 = x461 & n2786 ;
  assign n2919 = ~n2917 & ~n2918 ;
  assign n2920 = x429 & ~n2656 ;
  assign n2921 = x397 & n2656 ;
  assign n2922 = ~n2920 & ~n2921 ;
  assign n2923 = ~n2919 & n2922 ;
  assign n2924 = ~n2916 & ~n2923 ;
  assign n2925 = ~n2915 & n2924 ;
  assign n2926 = n2919 & ~n2922 ;
  assign n2927 = x430 & ~n2656 ;
  assign n2928 = x398 & n2656 ;
  assign n2929 = ~n2927 & ~n2928 ;
  assign n2930 = x494 & ~n2786 ;
  assign n2931 = x462 & n2786 ;
  assign n2932 = ~n2930 & ~n2931 ;
  assign n2933 = ~n2929 & n2932 ;
  assign n2934 = ~n2926 & ~n2933 ;
  assign n2935 = ~n2925 & n2934 ;
  assign n2936 = x431 & ~n2656 ;
  assign n2937 = x399 & n2656 ;
  assign n2938 = ~n2936 & ~n2937 ;
  assign n2939 = x495 & ~n2786 ;
  assign n2940 = x463 & n2786 ;
  assign n2941 = ~n2939 & ~n2940 ;
  assign n2942 = n2938 & ~n2941 ;
  assign n2943 = n2929 & ~n2932 ;
  assign n2944 = ~n2942 & ~n2943 ;
  assign n2945 = ~n2935 & n2944 ;
  assign n2946 = x496 & ~n2786 ;
  assign n2947 = x464 & n2786 ;
  assign n2948 = ~n2946 & ~n2947 ;
  assign n2949 = x432 & ~n2656 ;
  assign n2950 = x400 & n2656 ;
  assign n2951 = ~n2949 & ~n2950 ;
  assign n2952 = n2948 & ~n2951 ;
  assign n2953 = ~n2938 & n2941 ;
  assign n2954 = ~n2952 & ~n2953 ;
  assign n2955 = ~n2945 & n2954 ;
  assign n2956 = ~n2948 & n2951 ;
  assign n2957 = x497 & ~n2786 ;
  assign n2958 = x465 & n2786 ;
  assign n2959 = ~n2957 & ~n2958 ;
  assign n2960 = x433 & ~n2656 ;
  assign n2961 = x401 & n2656 ;
  assign n2962 = ~n2960 & ~n2961 ;
  assign n2963 = ~n2959 & n2962 ;
  assign n2964 = ~n2956 & ~n2963 ;
  assign n2965 = ~n2955 & n2964 ;
  assign n2966 = n2959 & ~n2962 ;
  assign n2967 = x434 & ~n2656 ;
  assign n2968 = x402 & n2656 ;
  assign n2969 = ~n2967 & ~n2968 ;
  assign n2970 = x498 & ~n2786 ;
  assign n2971 = x466 & n2786 ;
  assign n2972 = ~n2970 & ~n2971 ;
  assign n2973 = ~n2969 & n2972 ;
  assign n2974 = ~n2966 & ~n2973 ;
  assign n2975 = ~n2965 & n2974 ;
  assign n2976 = x435 & ~n2656 ;
  assign n2977 = x403 & n2656 ;
  assign n2978 = ~n2976 & ~n2977 ;
  assign n2979 = x499 & ~n2786 ;
  assign n2980 = x467 & n2786 ;
  assign n2981 = ~n2979 & ~n2980 ;
  assign n2982 = n2978 & ~n2981 ;
  assign n2983 = n2969 & ~n2972 ;
  assign n2984 = ~n2982 & ~n2983 ;
  assign n2985 = ~n2975 & n2984 ;
  assign n2986 = x500 & ~n2786 ;
  assign n2987 = x468 & n2786 ;
  assign n2988 = ~n2986 & ~n2987 ;
  assign n2989 = x436 & ~n2656 ;
  assign n2990 = x404 & n2656 ;
  assign n2991 = ~n2989 & ~n2990 ;
  assign n2992 = n2988 & ~n2991 ;
  assign n2993 = ~n2978 & n2981 ;
  assign n2994 = ~n2992 & ~n2993 ;
  assign n2995 = ~n2985 & n2994 ;
  assign n2996 = ~n2988 & n2991 ;
  assign n2997 = x501 & ~n2786 ;
  assign n2998 = x469 & n2786 ;
  assign n2999 = ~n2997 & ~n2998 ;
  assign n3000 = x437 & ~n2656 ;
  assign n3001 = x405 & n2656 ;
  assign n3002 = ~n3000 & ~n3001 ;
  assign n3003 = ~n2999 & n3002 ;
  assign n3004 = ~n2996 & ~n3003 ;
  assign n3005 = ~n2995 & n3004 ;
  assign n3006 = n2999 & ~n3002 ;
  assign n3007 = x438 & ~n2656 ;
  assign n3008 = x406 & n2656 ;
  assign n3009 = ~n3007 & ~n3008 ;
  assign n3010 = x502 & ~n2786 ;
  assign n3011 = x470 & n2786 ;
  assign n3012 = ~n3010 & ~n3011 ;
  assign n3013 = ~n3009 & n3012 ;
  assign n3014 = ~n3006 & ~n3013 ;
  assign n3015 = ~n3005 & n3014 ;
  assign n3016 = x439 & ~n2656 ;
  assign n3017 = x407 & n2656 ;
  assign n3018 = ~n3016 & ~n3017 ;
  assign n3019 = x503 & ~n2786 ;
  assign n3020 = x471 & n2786 ;
  assign n3021 = ~n3019 & ~n3020 ;
  assign n3022 = n3018 & ~n3021 ;
  assign n3023 = n3009 & ~n3012 ;
  assign n3024 = ~n3022 & ~n3023 ;
  assign n3025 = ~n3015 & n3024 ;
  assign n3026 = x504 & ~n2786 ;
  assign n3027 = x472 & n2786 ;
  assign n3028 = ~n3026 & ~n3027 ;
  assign n3029 = x440 & ~n2656 ;
  assign n3030 = x408 & n2656 ;
  assign n3031 = ~n3029 & ~n3030 ;
  assign n3032 = n3028 & ~n3031 ;
  assign n3033 = ~n3018 & n3021 ;
  assign n3034 = ~n3032 & ~n3033 ;
  assign n3035 = ~n3025 & n3034 ;
  assign n3036 = ~n3028 & n3031 ;
  assign n3037 = x441 & ~n2656 ;
  assign n3038 = x409 & n2656 ;
  assign n3039 = ~n3037 & ~n3038 ;
  assign n3040 = x505 & ~n2786 ;
  assign n3041 = x473 & n2786 ;
  assign n3042 = ~n3040 & ~n3041 ;
  assign n3043 = n3039 & ~n3042 ;
  assign n3044 = ~n3036 & ~n3043 ;
  assign n3045 = ~n3035 & n3044 ;
  assign n3046 = ~n3039 & n3042 ;
  assign n3047 = x442 & ~n2656 ;
  assign n3048 = x410 & n2656 ;
  assign n3049 = ~n3047 & ~n3048 ;
  assign n3050 = x506 & ~n2786 ;
  assign n3051 = x474 & n2786 ;
  assign n3052 = ~n3050 & ~n3051 ;
  assign n3053 = ~n3049 & n3052 ;
  assign n3054 = ~n3046 & ~n3053 ;
  assign n3055 = ~n3045 & n3054 ;
  assign n3056 = x443 & ~n2656 ;
  assign n3057 = x411 & n2656 ;
  assign n3058 = ~n3056 & ~n3057 ;
  assign n3059 = x507 & ~n2786 ;
  assign n3060 = x475 & n2786 ;
  assign n3061 = ~n3059 & ~n3060 ;
  assign n3062 = n3058 & ~n3061 ;
  assign n3063 = n3049 & ~n3052 ;
  assign n3064 = ~n3062 & ~n3063 ;
  assign n3065 = ~n3055 & n3064 ;
  assign n3066 = x508 & ~n2786 ;
  assign n3067 = x476 & n2786 ;
  assign n3068 = ~n3066 & ~n3067 ;
  assign n3069 = x444 & ~n2656 ;
  assign n3070 = x412 & n2656 ;
  assign n3071 = ~n3069 & ~n3070 ;
  assign n3072 = n3068 & ~n3071 ;
  assign n3073 = ~n3058 & n3061 ;
  assign n3074 = ~n3072 & ~n3073 ;
  assign n3075 = ~n3065 & n3074 ;
  assign n3076 = ~n3068 & n3071 ;
  assign n3077 = x509 & ~n2786 ;
  assign n3078 = x477 & n2786 ;
  assign n3079 = ~n3077 & ~n3078 ;
  assign n3080 = x445 & ~n2656 ;
  assign n3081 = x413 & n2656 ;
  assign n3082 = ~n3080 & ~n3081 ;
  assign n3083 = ~n3079 & n3082 ;
  assign n3084 = ~n3076 & ~n3083 ;
  assign n3085 = ~n3075 & n3084 ;
  assign n3086 = n2789 & ~n2792 ;
  assign n3087 = n3079 & ~n3082 ;
  assign n3088 = ~n3086 & ~n3087 ;
  assign n3089 = ~n3085 & n3088 ;
  assign n3090 = ~n2793 & ~n3089 ;
  assign n3091 = ~n2661 & ~n3090 ;
  assign n3092 = ~n2660 & ~n3091 ;
  assign n3093 = ~n2659 & n3092 ;
  assign n3094 = ~n2796 & ~n3092 ;
  assign n3095 = ~n3093 & ~n3094 ;
  assign n3096 = n2531 & ~n3095 ;
  assign n3097 = ~n2803 & n3092 ;
  assign n3098 = ~n2800 & ~n3092 ;
  assign n3099 = ~n3097 & ~n3098 ;
  assign n3100 = ~n2231 & n2524 ;
  assign n3101 = ~n2228 & ~n2524 ;
  assign n3102 = ~n3100 & ~n3101 ;
  assign n3103 = n3099 & ~n3102 ;
  assign n3104 = ~n3096 & n3103 ;
  assign n3105 = ~n2811 & n3092 ;
  assign n3106 = ~n2808 & ~n3092 ;
  assign n3107 = ~n3105 & ~n3106 ;
  assign n3108 = ~n2239 & n2524 ;
  assign n3109 = ~n2236 & ~n2524 ;
  assign n3110 = ~n3108 & ~n3109 ;
  assign n3111 = n3107 & ~n3110 ;
  assign n3112 = ~n2531 & n3095 ;
  assign n3113 = ~n3111 & ~n3112 ;
  assign n3114 = ~n3104 & n3113 ;
  assign n3115 = ~n3107 & n3110 ;
  assign n3116 = ~n2818 & n3092 ;
  assign n3117 = ~n2821 & ~n3092 ;
  assign n3118 = ~n3116 & ~n3117 ;
  assign n3119 = ~n2246 & n2524 ;
  assign n3120 = ~n2249 & ~n2524 ;
  assign n3121 = ~n3119 & ~n3120 ;
  assign n3122 = ~n3118 & n3121 ;
  assign n3123 = ~n3115 & ~n3122 ;
  assign n3124 = ~n3114 & n3123 ;
  assign n3125 = ~n2831 & n3092 ;
  assign n3126 = ~n2828 & ~n3092 ;
  assign n3127 = ~n3125 & ~n3126 ;
  assign n3128 = ~n2260 & n2524 ;
  assign n3129 = ~n2257 & ~n2524 ;
  assign n3130 = ~n3128 & ~n3129 ;
  assign n3131 = n3127 & ~n3130 ;
  assign n3132 = n3118 & ~n3121 ;
  assign n3133 = ~n3131 & ~n3132 ;
  assign n3134 = ~n3124 & n3133 ;
  assign n3135 = ~n2269 & n2524 ;
  assign n3136 = ~n2266 & ~n2524 ;
  assign n3137 = ~n3135 & ~n3136 ;
  assign n3138 = ~n2842 & n3092 ;
  assign n3139 = ~n2839 & ~n3092 ;
  assign n3140 = ~n3138 & ~n3139 ;
  assign n3141 = n3137 & ~n3140 ;
  assign n3142 = ~n3127 & n3130 ;
  assign n3143 = ~n3141 & ~n3142 ;
  assign n3144 = ~n3134 & n3143 ;
  assign n3145 = ~n2849 & n3092 ;
  assign n3146 = ~n2852 & ~n3092 ;
  assign n3147 = ~n3145 & ~n3146 ;
  assign n3148 = ~n2279 & n2524 ;
  assign n3149 = ~n2276 & ~n2524 ;
  assign n3150 = ~n3148 & ~n3149 ;
  assign n3151 = n3147 & ~n3150 ;
  assign n3152 = ~n3137 & n3140 ;
  assign n3153 = ~n3151 & ~n3152 ;
  assign n3154 = ~n3144 & n3153 ;
  assign n3155 = ~n2286 & n2524 ;
  assign n3156 = ~n2289 & ~n2524 ;
  assign n3157 = ~n3155 & ~n3156 ;
  assign n3158 = ~n2859 & n3092 ;
  assign n3159 = ~n2862 & ~n3092 ;
  assign n3160 = ~n3158 & ~n3159 ;
  assign n3161 = n3157 & ~n3160 ;
  assign n3162 = ~n3147 & n3150 ;
  assign n3163 = ~n3161 & ~n3162 ;
  assign n3164 = ~n3154 & n3163 ;
  assign n3165 = ~n2871 & n3092 ;
  assign n3166 = ~n2868 & ~n3092 ;
  assign n3167 = ~n3165 & ~n3166 ;
  assign n3168 = ~n2300 & n2524 ;
  assign n3169 = ~n2297 & ~n2524 ;
  assign n3170 = ~n3168 & ~n3169 ;
  assign n3171 = n3167 & ~n3170 ;
  assign n3172 = ~n3157 & n3160 ;
  assign n3173 = ~n3171 & ~n3172 ;
  assign n3174 = ~n3164 & n3173 ;
  assign n3175 = ~n2310 & n2524 ;
  assign n3176 = ~n2307 & ~n2524 ;
  assign n3177 = ~n3175 & ~n3176 ;
  assign n3178 = ~n2882 & n3092 ;
  assign n3179 = ~n2879 & ~n3092 ;
  assign n3180 = ~n3178 & ~n3179 ;
  assign n3181 = n3177 & ~n3180 ;
  assign n3182 = ~n3167 & n3170 ;
  assign n3183 = ~n3181 & ~n3182 ;
  assign n3184 = ~n3174 & n3183 ;
  assign n3185 = ~n2889 & n3092 ;
  assign n3186 = ~n2892 & ~n3092 ;
  assign n3187 = ~n3185 & ~n3186 ;
  assign n3188 = ~n2317 & n2524 ;
  assign n3189 = ~n2320 & ~n2524 ;
  assign n3190 = ~n3188 & ~n3189 ;
  assign n3191 = n3187 & ~n3190 ;
  assign n3192 = ~n3177 & n3180 ;
  assign n3193 = ~n3191 & ~n3192 ;
  assign n3194 = ~n3184 & n3193 ;
  assign n3195 = ~n2326 & n2524 ;
  assign n3196 = ~n2329 & ~n2524 ;
  assign n3197 = ~n3195 & ~n3196 ;
  assign n3198 = ~n2898 & n3092 ;
  assign n3199 = ~n2901 & ~n3092 ;
  assign n3200 = ~n3198 & ~n3199 ;
  assign n3201 = n3197 & ~n3200 ;
  assign n3202 = ~n3187 & n3190 ;
  assign n3203 = ~n3201 & ~n3202 ;
  assign n3204 = ~n3194 & n3203 ;
  assign n3205 = ~n2911 & n3092 ;
  assign n3206 = ~n2908 & ~n3092 ;
  assign n3207 = ~n3205 & ~n3206 ;
  assign n3208 = ~n2339 & n2524 ;
  assign n3209 = ~n2336 & ~n2524 ;
  assign n3210 = ~n3208 & ~n3209 ;
  assign n3211 = n3207 & ~n3210 ;
  assign n3212 = ~n3197 & n3200 ;
  assign n3213 = ~n3211 & ~n3212 ;
  assign n3214 = ~n3204 & n3213 ;
  assign n3215 = ~n2350 & n2524 ;
  assign n3216 = ~n2347 & ~n2524 ;
  assign n3217 = ~n3215 & ~n3216 ;
  assign n3218 = ~n2922 & n3092 ;
  assign n3219 = ~n2919 & ~n3092 ;
  assign n3220 = ~n3218 & ~n3219 ;
  assign n3221 = n3217 & ~n3220 ;
  assign n3222 = ~n3207 & n3210 ;
  assign n3223 = ~n3221 & ~n3222 ;
  assign n3224 = ~n3214 & n3223 ;
  assign n3225 = ~n2929 & n3092 ;
  assign n3226 = ~n2932 & ~n3092 ;
  assign n3227 = ~n3225 & ~n3226 ;
  assign n3228 = ~n2357 & n2524 ;
  assign n3229 = ~n2360 & ~n2524 ;
  assign n3230 = ~n3228 & ~n3229 ;
  assign n3231 = n3227 & ~n3230 ;
  assign n3232 = ~n3217 & n3220 ;
  assign n3233 = ~n3231 & ~n3232 ;
  assign n3234 = ~n3224 & n3233 ;
  assign n3235 = ~n2366 & n2524 ;
  assign n3236 = ~n2369 & ~n2524 ;
  assign n3237 = ~n3235 & ~n3236 ;
  assign n3238 = ~n2938 & n3092 ;
  assign n3239 = ~n2941 & ~n3092 ;
  assign n3240 = ~n3238 & ~n3239 ;
  assign n3241 = n3237 & ~n3240 ;
  assign n3242 = ~n3227 & n3230 ;
  assign n3243 = ~n3241 & ~n3242 ;
  assign n3244 = ~n3234 & n3243 ;
  assign n3245 = ~n2951 & n3092 ;
  assign n3246 = ~n2948 & ~n3092 ;
  assign n3247 = ~n3245 & ~n3246 ;
  assign n3248 = ~n2379 & n2524 ;
  assign n3249 = ~n2376 & ~n2524 ;
  assign n3250 = ~n3248 & ~n3249 ;
  assign n3251 = n3247 & ~n3250 ;
  assign n3252 = ~n3237 & n3240 ;
  assign n3253 = ~n3251 & ~n3252 ;
  assign n3254 = ~n3244 & n3253 ;
  assign n3255 = ~n2390 & n2524 ;
  assign n3256 = ~n2387 & ~n2524 ;
  assign n3257 = ~n3255 & ~n3256 ;
  assign n3258 = ~n2962 & n3092 ;
  assign n3259 = ~n2959 & ~n3092 ;
  assign n3260 = ~n3258 & ~n3259 ;
  assign n3261 = n3257 & ~n3260 ;
  assign n3262 = ~n3247 & n3250 ;
  assign n3263 = ~n3261 & ~n3262 ;
  assign n3264 = ~n3254 & n3263 ;
  assign n3265 = ~n2969 & n3092 ;
  assign n3266 = ~n2972 & ~n3092 ;
  assign n3267 = ~n3265 & ~n3266 ;
  assign n3268 = ~n2397 & n2524 ;
  assign n3269 = ~n2400 & ~n2524 ;
  assign n3270 = ~n3268 & ~n3269 ;
  assign n3271 = n3267 & ~n3270 ;
  assign n3272 = ~n3257 & n3260 ;
  assign n3273 = ~n3271 & ~n3272 ;
  assign n3274 = ~n3264 & n3273 ;
  assign n3275 = ~n2406 & n2524 ;
  assign n3276 = ~n2409 & ~n2524 ;
  assign n3277 = ~n3275 & ~n3276 ;
  assign n3278 = ~n2978 & n3092 ;
  assign n3279 = ~n2981 & ~n3092 ;
  assign n3280 = ~n3278 & ~n3279 ;
  assign n3281 = n3277 & ~n3280 ;
  assign n3282 = ~n3267 & n3270 ;
  assign n3283 = ~n3281 & ~n3282 ;
  assign n3284 = ~n3274 & n3283 ;
  assign n3285 = ~n2991 & n3092 ;
  assign n3286 = ~n2988 & ~n3092 ;
  assign n3287 = ~n3285 & ~n3286 ;
  assign n3288 = ~n2419 & n2524 ;
  assign n3289 = ~n2416 & ~n2524 ;
  assign n3290 = ~n3288 & ~n3289 ;
  assign n3291 = n3287 & ~n3290 ;
  assign n3292 = ~n3277 & n3280 ;
  assign n3293 = ~n3291 & ~n3292 ;
  assign n3294 = ~n3284 & n3293 ;
  assign n3295 = ~n2430 & n2524 ;
  assign n3296 = ~n2427 & ~n2524 ;
  assign n3297 = ~n3295 & ~n3296 ;
  assign n3298 = ~n3002 & n3092 ;
  assign n3299 = ~n2999 & ~n3092 ;
  assign n3300 = ~n3298 & ~n3299 ;
  assign n3301 = n3297 & ~n3300 ;
  assign n3302 = ~n3287 & n3290 ;
  assign n3303 = ~n3301 & ~n3302 ;
  assign n3304 = ~n3294 & n3303 ;
  assign n3305 = ~n3009 & n3092 ;
  assign n3306 = ~n3012 & ~n3092 ;
  assign n3307 = ~n3305 & ~n3306 ;
  assign n3308 = ~n2437 & n2524 ;
  assign n3309 = ~n2440 & ~n2524 ;
  assign n3310 = ~n3308 & ~n3309 ;
  assign n3311 = n3307 & ~n3310 ;
  assign n3312 = ~n3297 & n3300 ;
  assign n3313 = ~n3311 & ~n3312 ;
  assign n3314 = ~n3304 & n3313 ;
  assign n3315 = ~n2446 & n2524 ;
  assign n3316 = ~n2449 & ~n2524 ;
  assign n3317 = ~n3315 & ~n3316 ;
  assign n3318 = ~n3018 & n3092 ;
  assign n3319 = ~n3021 & ~n3092 ;
  assign n3320 = ~n3318 & ~n3319 ;
  assign n3321 = n3317 & ~n3320 ;
  assign n3322 = ~n3307 & n3310 ;
  assign n3323 = ~n3321 & ~n3322 ;
  assign n3324 = ~n3314 & n3323 ;
  assign n3325 = ~n3031 & n3092 ;
  assign n3326 = ~n3028 & ~n3092 ;
  assign n3327 = ~n3325 & ~n3326 ;
  assign n3328 = ~n2459 & n2524 ;
  assign n3329 = ~n2456 & ~n2524 ;
  assign n3330 = ~n3328 & ~n3329 ;
  assign n3331 = n3327 & ~n3330 ;
  assign n3332 = ~n3317 & n3320 ;
  assign n3333 = ~n3331 & ~n3332 ;
  assign n3334 = ~n3324 & n3333 ;
  assign n3335 = ~n3039 & n3092 ;
  assign n3336 = ~n3042 & ~n3092 ;
  assign n3337 = ~n3335 & ~n3336 ;
  assign n3338 = ~n2470 & n2524 ;
  assign n3339 = ~n2467 & ~n2524 ;
  assign n3340 = ~n3338 & ~n3339 ;
  assign n3341 = ~n3337 & n3340 ;
  assign n3342 = ~n3327 & n3330 ;
  assign n3343 = ~n3341 & ~n3342 ;
  assign n3344 = ~n3334 & n3343 ;
  assign n3345 = ~n3049 & n3092 ;
  assign n3346 = ~n3052 & ~n3092 ;
  assign n3347 = ~n3345 & ~n3346 ;
  assign n3348 = ~n2477 & n2524 ;
  assign n3349 = ~n2480 & ~n2524 ;
  assign n3350 = ~n3348 & ~n3349 ;
  assign n3351 = n3347 & ~n3350 ;
  assign n3352 = n3337 & ~n3340 ;
  assign n3353 = ~n3351 & ~n3352 ;
  assign n3354 = ~n3344 & n3353 ;
  assign n3355 = ~n3347 & n3350 ;
  assign n3356 = ~n3058 & n3092 ;
  assign n3357 = ~n3061 & ~n3092 ;
  assign n3358 = ~n3356 & ~n3357 ;
  assign n3359 = n2527 & ~n3358 ;
  assign n3360 = ~n3355 & ~n3359 ;
  assign n3361 = ~n3354 & n3360 ;
  assign n3362 = ~n2527 & n3358 ;
  assign n3363 = ~n2496 & n2524 ;
  assign n3364 = ~n2493 & ~n2524 ;
  assign n3365 = ~n3363 & ~n3364 ;
  assign n3366 = ~n3071 & n3092 ;
  assign n3367 = ~n3068 & ~n3092 ;
  assign n3368 = ~n3366 & ~n3367 ;
  assign n3369 = ~n3365 & n3368 ;
  assign n3370 = ~n3362 & ~n3369 ;
  assign n3371 = ~n3361 & n3370 ;
  assign n3372 = n3365 & ~n3368 ;
  assign n3373 = ~n2507 & n2524 ;
  assign n3374 = ~n2504 & ~n2524 ;
  assign n3375 = ~n3373 & ~n3374 ;
  assign n3376 = ~n3082 & n3092 ;
  assign n3377 = ~n3079 & ~n3092 ;
  assign n3378 = ~n3376 & ~n3377 ;
  assign n3379 = n3375 & ~n3378 ;
  assign n3380 = ~n3372 & ~n3379 ;
  assign n3381 = ~n3371 & n3380 ;
  assign n3382 = ~n3375 & n3378 ;
  assign n3383 = ~n2514 & n2524 ;
  assign n3384 = ~n2517 & ~n2524 ;
  assign n3385 = ~n3383 & ~n3384 ;
  assign n3386 = ~n2792 & n3092 ;
  assign n3387 = ~n2789 & ~n3092 ;
  assign n3388 = ~n3386 & ~n3387 ;
  assign n3389 = ~n3385 & n3388 ;
  assign n3390 = ~n3382 & ~n3389 ;
  assign n3391 = ~n3381 & n3390 ;
  assign n3392 = n515 & ~n518 ;
  assign n3393 = n3385 & ~n3388 ;
  assign n3394 = ~n3392 & ~n3393 ;
  assign n3395 = ~n3391 & n3394 ;
  assign n3396 = ~n2528 & ~n3395 ;
  assign n3397 = n2527 & ~n3396 ;
  assign n3398 = n3358 & n3396 ;
  assign n3399 = ~n3397 & ~n3398 ;
  assign n3400 = ~n1963 & n3399 ;
  assign n3401 = n3350 & ~n3396 ;
  assign n3402 = n3347 & n3396 ;
  assign n3403 = ~n3401 & ~n3402 ;
  assign n3404 = n1914 & ~n1960 ;
  assign n3405 = n1911 & n1960 ;
  assign n3406 = ~n3404 & ~n3405 ;
  assign n3407 = ~n3403 & n3406 ;
  assign n3408 = ~n1904 & ~n1960 ;
  assign n3409 = ~n1901 & n1960 ;
  assign n3410 = ~n3408 & ~n3409 ;
  assign n3411 = ~n3340 & ~n3396 ;
  assign n3412 = ~n3337 & n3396 ;
  assign n3413 = ~n3411 & ~n3412 ;
  assign n3414 = ~n3410 & n3413 ;
  assign n3415 = ~n1894 & ~n1960 ;
  assign n3416 = ~n1891 & n1960 ;
  assign n3417 = ~n3415 & ~n3416 ;
  assign n3418 = ~n3330 & ~n3396 ;
  assign n3419 = ~n3327 & n3396 ;
  assign n3420 = ~n3418 & ~n3419 ;
  assign n3421 = n3417 & ~n3420 ;
  assign n3422 = ~n3317 & ~n3396 ;
  assign n3423 = ~n3320 & n3396 ;
  assign n3424 = ~n3422 & ~n3423 ;
  assign n3425 = ~n3277 & ~n3396 ;
  assign n3426 = ~n3280 & n3396 ;
  assign n3427 = ~n3425 & ~n3426 ;
  assign n3428 = ~n3237 & ~n3396 ;
  assign n3429 = ~n3240 & n3396 ;
  assign n3430 = ~n3428 & ~n3429 ;
  assign n3431 = ~n3197 & ~n3396 ;
  assign n3432 = ~n3200 & n3396 ;
  assign n3433 = ~n3431 & ~n3432 ;
  assign n3434 = ~n3150 & ~n3396 ;
  assign n3435 = ~n3147 & n3396 ;
  assign n3436 = ~n3434 & ~n3435 ;
  assign n3437 = ~n1714 & ~n1960 ;
  assign n3438 = ~n1711 & n1960 ;
  assign n3439 = ~n3437 & ~n3438 ;
  assign n3440 = n3436 & ~n3439 ;
  assign n3441 = ~n1701 & ~n1960 ;
  assign n3442 = ~n1704 & n1960 ;
  assign n3443 = ~n3441 & ~n3442 ;
  assign n3444 = ~n3137 & ~n3396 ;
  assign n3445 = ~n3140 & n3396 ;
  assign n3446 = ~n3444 & ~n3445 ;
  assign n3447 = n3443 & ~n3446 ;
  assign n3448 = ~n3443 & n3446 ;
  assign n3449 = ~n3130 & ~n3396 ;
  assign n3450 = ~n3127 & n3396 ;
  assign n3451 = ~n3449 & ~n3450 ;
  assign n3452 = ~n1694 & n1960 ;
  assign n3453 = ~n1691 & ~n1960 ;
  assign n3454 = ~n3452 & ~n3453 ;
  assign n3455 = ~n3451 & n3454 ;
  assign n3456 = ~n1095 & ~n1960 ;
  assign n3457 = ~n1659 & n1960 ;
  assign n3458 = ~n3456 & ~n3457 ;
  assign n3459 = ~n3095 & n3396 ;
  assign n3460 = ~n2531 & ~n3396 ;
  assign n3461 = ~n3459 & ~n3460 ;
  assign n3462 = n3458 & ~n3461 ;
  assign n3463 = ~n3102 & ~n3396 ;
  assign n3464 = ~n3099 & n3396 ;
  assign n3465 = ~n3463 & ~n3464 ;
  assign n3466 = ~n1666 & ~n1960 ;
  assign n3467 = ~n1663 & n1960 ;
  assign n3468 = ~n3466 & ~n3467 ;
  assign n3469 = n3465 & ~n3468 ;
  assign n3470 = ~n3462 & n3469 ;
  assign n3471 = ~n3110 & ~n3396 ;
  assign n3472 = ~n3107 & n3396 ;
  assign n3473 = ~n3471 & ~n3472 ;
  assign n3474 = ~n1674 & ~n1960 ;
  assign n3475 = ~n1671 & n1960 ;
  assign n3476 = ~n3474 & ~n3475 ;
  assign n3477 = n3473 & ~n3476 ;
  assign n3478 = ~n3458 & n3461 ;
  assign n3479 = ~n3477 & ~n3478 ;
  assign n3480 = ~n3470 & n3479 ;
  assign n3481 = n3121 & ~n3396 ;
  assign n3482 = n3118 & n3396 ;
  assign n3483 = ~n3481 & ~n3482 ;
  assign n3484 = ~n1682 & ~n1960 ;
  assign n3485 = n1685 & n1960 ;
  assign n3486 = ~n3484 & ~n3485 ;
  assign n3487 = n3483 & n3486 ;
  assign n3488 = ~n3473 & n3476 ;
  assign n3489 = ~n3487 & ~n3488 ;
  assign n3490 = ~n3480 & n3489 ;
  assign n3491 = n3451 & ~n3454 ;
  assign n3492 = ~n3483 & ~n3486 ;
  assign n3493 = ~n3491 & ~n3492 ;
  assign n3494 = ~n3490 & n3493 ;
  assign n3495 = ~n3455 & ~n3494 ;
  assign n3496 = ~n3448 & ~n3495 ;
  assign n3497 = ~n3447 & ~n3496 ;
  assign n3498 = ~n3440 & ~n3497 ;
  assign n3499 = ~n3436 & n3439 ;
  assign n3500 = ~n1721 & ~n1960 ;
  assign n3501 = ~n1724 & n1960 ;
  assign n3502 = ~n3500 & ~n3501 ;
  assign n3503 = ~n3157 & ~n3396 ;
  assign n3504 = ~n3160 & n3396 ;
  assign n3505 = ~n3503 & ~n3504 ;
  assign n3506 = n3502 & ~n3505 ;
  assign n3507 = ~n3499 & ~n3506 ;
  assign n3508 = ~n3498 & n3507 ;
  assign n3509 = ~n3502 & n3505 ;
  assign n3510 = ~n3170 & ~n3396 ;
  assign n3511 = ~n3167 & n3396 ;
  assign n3512 = ~n3510 & ~n3511 ;
  assign n3513 = ~n1734 & ~n1960 ;
  assign n3514 = ~n1731 & n1960 ;
  assign n3515 = ~n3513 & ~n3514 ;
  assign n3516 = n3512 & ~n3515 ;
  assign n3517 = ~n3509 & ~n3516 ;
  assign n3518 = ~n3508 & n3517 ;
  assign n3519 = ~n3512 & n3515 ;
  assign n3520 = ~n1741 & ~n1960 ;
  assign n3521 = ~n1744 & n1960 ;
  assign n3522 = ~n3520 & ~n3521 ;
  assign n3523 = ~n3177 & ~n3396 ;
  assign n3524 = ~n3180 & n3396 ;
  assign n3525 = ~n3523 & ~n3524 ;
  assign n3526 = n3522 & ~n3525 ;
  assign n3527 = ~n3519 & ~n3526 ;
  assign n3528 = ~n3518 & n3527 ;
  assign n3529 = ~n3522 & n3525 ;
  assign n3530 = n3190 & ~n3396 ;
  assign n3531 = n3187 & n3396 ;
  assign n3532 = ~n3530 & ~n3531 ;
  assign n3533 = n1754 & ~n1960 ;
  assign n3534 = n1751 & n1960 ;
  assign n3535 = ~n3533 & ~n3534 ;
  assign n3536 = ~n3532 & n3535 ;
  assign n3537 = ~n3529 & ~n3536 ;
  assign n3538 = ~n3528 & n3537 ;
  assign n3539 = n3532 & ~n3535 ;
  assign n3540 = ~n3538 & ~n3539 ;
  assign n3541 = ~n1761 & ~n1960 ;
  assign n3542 = ~n1764 & n1960 ;
  assign n3543 = ~n3541 & ~n3542 ;
  assign n3544 = ~n3540 & n3543 ;
  assign n3545 = n3433 & ~n3544 ;
  assign n3546 = ~n1774 & ~n1960 ;
  assign n3547 = ~n1771 & n1960 ;
  assign n3548 = ~n3546 & ~n3547 ;
  assign n3549 = ~n3210 & ~n3396 ;
  assign n3550 = ~n3207 & n3396 ;
  assign n3551 = ~n3549 & ~n3550 ;
  assign n3552 = ~n3548 & n3551 ;
  assign n3553 = n3540 & ~n3543 ;
  assign n3554 = ~n3552 & ~n3553 ;
  assign n3555 = ~n3545 & n3554 ;
  assign n3556 = n3548 & ~n3551 ;
  assign n3557 = ~n1781 & ~n1960 ;
  assign n3558 = ~n1784 & n1960 ;
  assign n3559 = ~n3557 & ~n3558 ;
  assign n3560 = ~n3217 & ~n3396 ;
  assign n3561 = ~n3220 & n3396 ;
  assign n3562 = ~n3560 & ~n3561 ;
  assign n3563 = n3559 & ~n3562 ;
  assign n3564 = ~n3556 & ~n3563 ;
  assign n3565 = ~n3555 & n3564 ;
  assign n3566 = ~n3559 & n3562 ;
  assign n3567 = n3230 & ~n3396 ;
  assign n3568 = n3227 & n3396 ;
  assign n3569 = ~n3567 & ~n3568 ;
  assign n3570 = n1794 & ~n1960 ;
  assign n3571 = n1791 & n1960 ;
  assign n3572 = ~n3570 & ~n3571 ;
  assign n3573 = ~n3569 & n3572 ;
  assign n3574 = ~n3566 & ~n3573 ;
  assign n3575 = ~n3565 & n3574 ;
  assign n3576 = n3569 & ~n3572 ;
  assign n3577 = ~n3575 & ~n3576 ;
  assign n3578 = ~n1801 & ~n1960 ;
  assign n3579 = ~n1804 & n1960 ;
  assign n3580 = ~n3578 & ~n3579 ;
  assign n3581 = ~n3577 & n3580 ;
  assign n3582 = n3430 & ~n3581 ;
  assign n3583 = ~n1814 & ~n1960 ;
  assign n3584 = ~n1811 & n1960 ;
  assign n3585 = ~n3583 & ~n3584 ;
  assign n3586 = ~n3250 & ~n3396 ;
  assign n3587 = ~n3247 & n3396 ;
  assign n3588 = ~n3586 & ~n3587 ;
  assign n3589 = ~n3585 & n3588 ;
  assign n3590 = n3577 & ~n3580 ;
  assign n3591 = ~n3589 & ~n3590 ;
  assign n3592 = ~n3582 & n3591 ;
  assign n3593 = n3585 & ~n3588 ;
  assign n3594 = ~n1821 & ~n1960 ;
  assign n3595 = ~n1824 & n1960 ;
  assign n3596 = ~n3594 & ~n3595 ;
  assign n3597 = ~n3257 & ~n3396 ;
  assign n3598 = ~n3260 & n3396 ;
  assign n3599 = ~n3597 & ~n3598 ;
  assign n3600 = n3596 & ~n3599 ;
  assign n3601 = ~n3593 & ~n3600 ;
  assign n3602 = ~n3592 & n3601 ;
  assign n3603 = ~n3596 & n3599 ;
  assign n3604 = n3270 & ~n3396 ;
  assign n3605 = n3267 & n3396 ;
  assign n3606 = ~n3604 & ~n3605 ;
  assign n3607 = n1834 & ~n1960 ;
  assign n3608 = n1831 & n1960 ;
  assign n3609 = ~n3607 & ~n3608 ;
  assign n3610 = ~n3606 & n3609 ;
  assign n3611 = ~n3603 & ~n3610 ;
  assign n3612 = ~n3602 & n3611 ;
  assign n3613 = n3606 & ~n3609 ;
  assign n3614 = ~n3612 & ~n3613 ;
  assign n3615 = ~n1841 & ~n1960 ;
  assign n3616 = ~n1844 & n1960 ;
  assign n3617 = ~n3615 & ~n3616 ;
  assign n3618 = ~n3614 & n3617 ;
  assign n3619 = n3427 & ~n3618 ;
  assign n3620 = ~n1854 & ~n1960 ;
  assign n3621 = ~n1851 & n1960 ;
  assign n3622 = ~n3620 & ~n3621 ;
  assign n3623 = ~n3290 & ~n3396 ;
  assign n3624 = ~n3287 & n3396 ;
  assign n3625 = ~n3623 & ~n3624 ;
  assign n3626 = ~n3622 & n3625 ;
  assign n3627 = n3614 & ~n3617 ;
  assign n3628 = ~n3626 & ~n3627 ;
  assign n3629 = ~n3619 & n3628 ;
  assign n3630 = n3622 & ~n3625 ;
  assign n3631 = ~n1861 & ~n1960 ;
  assign n3632 = ~n1864 & n1960 ;
  assign n3633 = ~n3631 & ~n3632 ;
  assign n3634 = ~n3297 & ~n3396 ;
  assign n3635 = ~n3300 & n3396 ;
  assign n3636 = ~n3634 & ~n3635 ;
  assign n3637 = n3633 & ~n3636 ;
  assign n3638 = ~n3630 & ~n3637 ;
  assign n3639 = ~n3629 & n3638 ;
  assign n3640 = ~n3633 & n3636 ;
  assign n3641 = n3310 & ~n3396 ;
  assign n3642 = n3307 & n3396 ;
  assign n3643 = ~n3641 & ~n3642 ;
  assign n3644 = n1874 & ~n1960 ;
  assign n3645 = n1871 & n1960 ;
  assign n3646 = ~n3644 & ~n3645 ;
  assign n3647 = ~n3643 & n3646 ;
  assign n3648 = ~n3640 & ~n3647 ;
  assign n3649 = ~n3639 & n3648 ;
  assign n3650 = n3643 & ~n3646 ;
  assign n3651 = ~n3649 & ~n3650 ;
  assign n3652 = ~n1881 & ~n1960 ;
  assign n3653 = ~n1884 & n1960 ;
  assign n3654 = ~n3652 & ~n3653 ;
  assign n3655 = ~n3651 & n3654 ;
  assign n3656 = n3424 & ~n3655 ;
  assign n3657 = ~n3417 & n3420 ;
  assign n3658 = n3651 & ~n3654 ;
  assign n3659 = ~n3657 & ~n3658 ;
  assign n3660 = ~n3656 & n3659 ;
  assign n3661 = ~n3421 & ~n3660 ;
  assign n3662 = ~n3414 & ~n3661 ;
  assign n3663 = n3410 & ~n3413 ;
  assign n3664 = n3403 & ~n3406 ;
  assign n3665 = ~n3663 & ~n3664 ;
  assign n3666 = ~n3662 & n3665 ;
  assign n3667 = ~n3407 & ~n3666 ;
  assign n3668 = ~n3400 & ~n3667 ;
  assign n3669 = n1963 & ~n3399 ;
  assign n3670 = ~n3365 & ~n3396 ;
  assign n3671 = ~n3368 & n3396 ;
  assign n3672 = ~n3670 & ~n3671 ;
  assign n3673 = ~n1929 & ~n1960 ;
  assign n3674 = ~n1932 & n1960 ;
  assign n3675 = ~n3673 & ~n3674 ;
  assign n3676 = n3672 & ~n3675 ;
  assign n3677 = ~n3669 & ~n3676 ;
  assign n3678 = ~n3668 & n3677 ;
  assign n3679 = ~n3672 & n3675 ;
  assign n3680 = ~n1939 & ~n1960 ;
  assign n3681 = ~n1942 & n1960 ;
  assign n3682 = ~n3680 & ~n3681 ;
  assign n3683 = ~n3375 & ~n3396 ;
  assign n3684 = ~n3378 & n3396 ;
  assign n3685 = ~n3683 & ~n3684 ;
  assign n3686 = n3682 & ~n3685 ;
  assign n3687 = ~n3679 & ~n3686 ;
  assign n3688 = ~n3678 & n3687 ;
  assign n3689 = ~n3682 & n3685 ;
  assign n3690 = ~n3388 & n3396 ;
  assign n3691 = ~n3385 & ~n3396 ;
  assign n3692 = ~n3690 & ~n3691 ;
  assign n3693 = ~n1952 & n1960 ;
  assign n3694 = ~n1949 & ~n1960 ;
  assign n3695 = ~n3693 & ~n3694 ;
  assign n3696 = n3692 & ~n3695 ;
  assign n3697 = ~n3689 & ~n3696 ;
  assign n3698 = ~n3688 & n3697 ;
  assign n3699 = ~n519 & n526 ;
  assign n3700 = ~n3692 & n3695 ;
  assign n3701 = ~n3699 & ~n3700 ;
  assign n3702 = ~n3698 & n3701 ;
  assign n3703 = ~n527 & ~n3702 ;
  assign n3704 = n1960 & ~n3703 ;
  assign n3705 = n3396 & n3703 ;
  assign n3706 = ~n3704 & ~n3705 ;
  assign n3707 = ~n2524 & n3706 ;
  assign n3708 = ~n3092 & n3396 ;
  assign n3709 = ~n3707 & ~n3708 ;
  assign n3710 = n3703 & ~n3709 ;
  assign n3711 = ~n1088 & n3706 ;
  assign n3712 = ~n1656 & n1960 ;
  assign n3713 = ~n3711 & ~n3712 ;
  assign n3714 = ~n3703 & ~n3713 ;
  assign n3715 = ~n3710 & ~n3714 ;
  assign n3716 = n2088 & n3715 ;
  assign n3717 = n2221 & ~n3715 ;
  assign n3718 = n3706 & ~n3717 ;
  assign n3719 = ~n3716 & n3718 ;
  assign n3720 = n2656 & n3715 ;
  assign n3721 = n2786 & ~n3715 ;
  assign n3722 = ~n3706 & ~n3721 ;
  assign n3723 = ~n3720 & n3722 ;
  assign n3724 = ~n3719 & ~n3723 ;
  assign n3725 = n3703 & ~n3724 ;
  assign n3726 = n652 & n3715 ;
  assign n3727 = n785 & ~n3715 ;
  assign n3728 = n3706 & ~n3727 ;
  assign n3729 = ~n3726 & n3728 ;
  assign n3730 = n1220 & n3715 ;
  assign n3731 = n1350 & ~n3715 ;
  assign n3732 = ~n3706 & ~n3731 ;
  assign n3733 = ~n3730 & n3732 ;
  assign n3734 = ~n3729 & ~n3733 ;
  assign n3735 = ~n3703 & ~n3734 ;
  assign n3736 = ~n3725 & ~n3735 ;
  assign n3737 = ~n3465 & n3703 ;
  assign n3738 = ~n3468 & ~n3703 ;
  assign n3739 = ~n3737 & ~n3738 ;
  assign n3740 = n3458 & ~n3703 ;
  assign n3741 = n3461 & n3703 ;
  assign n3742 = ~n3740 & ~n3741 ;
  assign n3743 = ~n3473 & n3703 ;
  assign n3744 = ~n3476 & ~n3703 ;
  assign n3745 = ~n3743 & ~n3744 ;
  assign n3746 = ~n3486 & ~n3703 ;
  assign n3747 = n3483 & n3703 ;
  assign n3748 = ~n3746 & ~n3747 ;
  assign n3749 = ~n3451 & n3703 ;
  assign n3750 = ~n3454 & ~n3703 ;
  assign n3751 = ~n3749 & ~n3750 ;
  assign n3752 = ~n3446 & n3703 ;
  assign n3753 = ~n3443 & ~n3703 ;
  assign n3754 = ~n3752 & ~n3753 ;
  assign n3755 = ~n3436 & n3703 ;
  assign n3756 = ~n3439 & ~n3703 ;
  assign n3757 = ~n3755 & ~n3756 ;
  assign n3758 = ~n3505 & n3703 ;
  assign n3759 = ~n3502 & ~n3703 ;
  assign n3760 = ~n3758 & ~n3759 ;
  assign n3761 = ~n3512 & n3703 ;
  assign n3762 = ~n3515 & ~n3703 ;
  assign n3763 = ~n3761 & ~n3762 ;
  assign n3764 = ~n3525 & n3703 ;
  assign n3765 = ~n3522 & ~n3703 ;
  assign n3766 = ~n3764 & ~n3765 ;
  assign n3767 = ~n3532 & n3703 ;
  assign n3768 = ~n3535 & ~n3703 ;
  assign n3769 = ~n3767 & ~n3768 ;
  assign n3770 = ~n3433 & n3703 ;
  assign n3771 = ~n3543 & ~n3703 ;
  assign n3772 = ~n3770 & ~n3771 ;
  assign n3773 = ~n3551 & n3703 ;
  assign n3774 = ~n3548 & ~n3703 ;
  assign n3775 = ~n3773 & ~n3774 ;
  assign n3776 = ~n3562 & n3703 ;
  assign n3777 = ~n3559 & ~n3703 ;
  assign n3778 = ~n3776 & ~n3777 ;
  assign n3779 = ~n3569 & n3703 ;
  assign n3780 = ~n3572 & ~n3703 ;
  assign n3781 = ~n3779 & ~n3780 ;
  assign n3782 = ~n3430 & n3703 ;
  assign n3783 = ~n3580 & ~n3703 ;
  assign n3784 = ~n3782 & ~n3783 ;
  assign n3785 = ~n3588 & n3703 ;
  assign n3786 = ~n3585 & ~n3703 ;
  assign n3787 = ~n3785 & ~n3786 ;
  assign n3788 = ~n3599 & n3703 ;
  assign n3789 = ~n3596 & ~n3703 ;
  assign n3790 = ~n3788 & ~n3789 ;
  assign n3791 = ~n3606 & n3703 ;
  assign n3792 = ~n3609 & ~n3703 ;
  assign n3793 = ~n3791 & ~n3792 ;
  assign n3794 = ~n3427 & n3703 ;
  assign n3795 = ~n3617 & ~n3703 ;
  assign n3796 = ~n3794 & ~n3795 ;
  assign n3797 = ~n3625 & n3703 ;
  assign n3798 = ~n3622 & ~n3703 ;
  assign n3799 = ~n3797 & ~n3798 ;
  assign n3800 = ~n3636 & n3703 ;
  assign n3801 = ~n3633 & ~n3703 ;
  assign n3802 = ~n3800 & ~n3801 ;
  assign n3803 = ~n3643 & n3703 ;
  assign n3804 = ~n3646 & ~n3703 ;
  assign n3805 = ~n3803 & ~n3804 ;
  assign n3806 = ~n3424 & n3703 ;
  assign n3807 = ~n3654 & ~n3703 ;
  assign n3808 = ~n3806 & ~n3807 ;
  assign n3809 = ~n3420 & n3703 ;
  assign n3810 = ~n3417 & ~n3703 ;
  assign n3811 = ~n3809 & ~n3810 ;
  assign n3812 = ~n3413 & n3703 ;
  assign n3813 = ~n3410 & ~n3703 ;
  assign n3814 = ~n3812 & ~n3813 ;
  assign n3815 = ~n3403 & n3703 ;
  assign n3816 = ~n3406 & ~n3703 ;
  assign n3817 = ~n3815 & ~n3816 ;
  assign n3818 = n1963 & ~n3703 ;
  assign n3819 = n3399 & n3703 ;
  assign n3820 = ~n3818 & ~n3819 ;
  assign n3821 = ~n3672 & n3703 ;
  assign n3822 = ~n3675 & ~n3703 ;
  assign n3823 = ~n3821 & ~n3822 ;
  assign n3824 = ~n3685 & n3703 ;
  assign n3825 = ~n3682 & ~n3703 ;
  assign n3826 = ~n3824 & ~n3825 ;
  assign n3827 = ~n3692 & n3703 ;
  assign n3828 = ~n3695 & ~n3703 ;
  assign n3829 = ~n3827 & ~n3828 ;
  assign n3830 = n519 & n526 ;
  assign y0 = ~n3736 ;
  assign y1 = ~n3715 ;
  assign y2 = ~n3706 ;
  assign y3 = n3703 ;
  assign y4 = ~n3739 ;
  assign y5 = n3742 ;
  assign y6 = ~n3745 ;
  assign y7 = ~n3748 ;
  assign y8 = ~n3751 ;
  assign y9 = ~n3754 ;
  assign y10 = ~n3757 ;
  assign y11 = ~n3760 ;
  assign y12 = ~n3763 ;
  assign y13 = ~n3766 ;
  assign y14 = n3769 ;
  assign y15 = ~n3772 ;
  assign y16 = ~n3775 ;
  assign y17 = ~n3778 ;
  assign y18 = n3781 ;
  assign y19 = ~n3784 ;
  assign y20 = ~n3787 ;
  assign y21 = ~n3790 ;
  assign y22 = n3793 ;
  assign y23 = ~n3796 ;
  assign y24 = ~n3799 ;
  assign y25 = ~n3802 ;
  assign y26 = n3805 ;
  assign y27 = ~n3808 ;
  assign y28 = ~n3811 ;
  assign y29 = ~n3814 ;
  assign y30 = n3817 ;
  assign y31 = ~n3820 ;
  assign y32 = ~n3823 ;
  assign y33 = ~n3826 ;
  assign y34 = ~n3829 ;
  assign y35 = ~n3830 ;
endmodule
