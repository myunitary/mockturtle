module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 ;
  assign n61 = x27 & x28 ;
  assign n62 = x29 & n61 ;
  assign n64 = x9 & x10 ;
  assign n65 = n64 ^ x9 ;
  assign n66 = n65 ^ x10 ;
  assign n67 = x11 & ~n66 ;
  assign n68 = n67 ^ x11 ;
  assign n63 = ~x12 & ~x13 ;
  assign n69 = n68 ^ n63 ;
  assign n70 = n63 ^ x14 ;
  assign n71 = ~x14 & ~n70 ;
  assign n72 = n71 ^ x14 ;
  assign n73 = n72 ^ n68 ;
  assign n74 = ~n69 & n73 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = n75 ^ n68 ;
  assign n77 = x15 & ~x16 ;
  assign n78 = n76 & n77 ;
  assign n79 = n78 ^ x16 ;
  assign n80 = x17 & ~x18 ;
  assign n81 = n79 & n80 ;
  assign n82 = n81 ^ x18 ;
  assign n83 = x19 & x20 ;
  assign n84 = ~n82 & n83 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = ~x21 & ~x22 ;
  assign n87 = n85 & n86 ;
  assign n88 = n87 ^ n86 ;
  assign n89 = x23 & x24 ;
  assign n90 = x25 & ~x26 ;
  assign n91 = n89 & n90 ;
  assign n92 = ~n88 & n91 ;
  assign n93 = n92 ^ x26 ;
  assign n94 = n62 & ~n93 ;
  assign n95 = n94 ^ n62 ;
  assign n96 = x17 & ~n79 ;
  assign n97 = n96 ^ x17 ;
  assign n98 = n76 ^ x15 ;
  assign n99 = x15 & n76 ;
  assign n100 = x16 & n99 ;
  assign n101 = ~x12 & n68 ;
  assign n102 = ~x11 & x12 ;
  assign n103 = ~n66 & n102 ;
  assign n104 = ~n101 & ~n103 ;
  assign n105 = x20 & ~x21 ;
  assign n106 = ~x22 & x23 ;
  assign n107 = ~x1 & ~x2 ;
  assign n108 = n106 & n107 ;
  assign n109 = n105 & n108 ;
  assign n110 = ~x7 & ~x8 ;
  assign n111 = x9 & ~x10 ;
  assign n112 = n110 & n111 ;
  assign n113 = ~x3 & ~x4 ;
  assign n114 = ~x5 & ~x6 ;
  assign n115 = n113 & n114 ;
  assign n116 = n112 & n115 ;
  assign n117 = x24 & x25 ;
  assign n118 = ~x26 & n117 ;
  assign n119 = ~x13 & x14 ;
  assign n120 = ~x18 & x19 ;
  assign n121 = n119 & n120 ;
  assign n122 = n118 & n121 ;
  assign n123 = n116 & n122 ;
  assign n124 = n109 & n123 ;
  assign n125 = ~n104 & n124 ;
  assign n126 = ~n100 & n125 ;
  assign n127 = ~n98 & n126 ;
  assign n128 = n97 & n127 ;
  assign n129 = n95 & n128 ;
  assign n130 = n129 ^ n95 ;
  assign n131 = ~x17 & ~n79 ;
  assign n132 = x19 & x25 ;
  assign n133 = ~x26 & n132 ;
  assign n134 = n63 & n77 ;
  assign n135 = n133 & n134 ;
  assign n136 = n62 & n135 ;
  assign n137 = x0 & x1 ;
  assign n138 = ~n66 & n137 ;
  assign n139 = n105 & n106 ;
  assign n140 = n138 & n139 ;
  assign n141 = x6 & x7 ;
  assign n142 = x8 & x11 ;
  assign n143 = n141 & n142 ;
  assign n144 = x2 & x3 ;
  assign n145 = x4 & x5 ;
  assign n146 = n144 & n145 ;
  assign n147 = n143 & n146 ;
  assign n148 = n140 & n147 ;
  assign n149 = n136 & n148 ;
  assign n150 = n63 & n68 ;
  assign n151 = n150 ^ n63 ;
  assign n152 = n151 ^ x14 ;
  assign n153 = n149 & ~n152 ;
  assign n154 = ~n131 & n153 ;
  assign n155 = ~n82 & n154 ;
  assign n159 = n86 ^ n83 ;
  assign n168 = n159 ^ x23 ;
  assign n160 = n86 ^ x18 ;
  assign n161 = n159 & ~n160 ;
  assign n162 = n161 ^ x18 ;
  assign n163 = n162 ^ n97 ;
  assign n169 = n168 ^ n163 ;
  assign n170 = n97 ^ n83 ;
  assign n171 = n170 ^ n162 ;
  assign n172 = n169 & n171 ;
  assign n164 = n162 ^ n83 ;
  assign n157 = n86 ^ x23 ;
  assign n165 = n164 ^ n157 ;
  assign n166 = n163 & ~n165 ;
  assign n173 = n172 ^ n166 ;
  assign n174 = n173 ^ n162 ;
  assign n175 = n174 ^ n168 ;
  assign n176 = n166 ^ n97 ;
  assign n177 = n176 ^ x23 ;
  assign n178 = ~n175 & ~n177 ;
  assign n179 = n178 ^ n172 ;
  assign n167 = n166 ^ n161 ;
  assign n180 = n179 ^ n167 ;
  assign n156 = n83 ^ x18 ;
  assign n158 = n157 ^ n156 ;
  assign n181 = n180 ^ n158 ;
  assign n182 = n181 ^ x23 ;
  assign n183 = n182 ^ x24 ;
  assign n184 = ~n95 & ~n183 ;
  assign n185 = n155 & n184 ;
  assign n186 = n185 ^ n95 ;
  assign n187 = n130 & ~n186 ;
  assign n188 = n187 ^ n130 ;
  assign n189 = n188 ^ n186 ;
  assign n227 = x54 & x55 ;
  assign n245 = x53 & n227 ;
  assign n244 = ~x51 & ~x52 ;
  assign n249 = n245 ^ n244 ;
  assign n250 = n245 & n249 ;
  assign n190 = x39 & x40 ;
  assign n191 = n190 ^ x39 ;
  assign n192 = n191 ^ x40 ;
  assign n193 = x41 & x42 ;
  assign n194 = n193 ^ x41 ;
  assign n195 = n192 & n194 ;
  assign n196 = n195 ^ x42 ;
  assign n197 = ~x43 & x44 ;
  assign n198 = n196 & n197 ;
  assign n199 = n198 ^ n197 ;
  assign n200 = n199 ^ x44 ;
  assign n201 = x45 & ~x46 ;
  assign n202 = n200 & n201 ;
  assign n203 = n202 ^ x46 ;
  assign n240 = x47 & ~x48 ;
  assign n241 = n203 & n240 ;
  assign n242 = n241 ^ x48 ;
  assign n243 = n242 ^ x49 ;
  assign n220 = x49 & x50 ;
  assign n246 = n244 & n245 ;
  assign n247 = n220 & n246 ;
  assign n248 = ~n243 & n247 ;
  assign n251 = n250 ^ n248 ;
  assign n252 = n251 ^ n245 ;
  assign n253 = n252 ^ n245 ;
  assign n254 = x57 & x58 ;
  assign n255 = x59 & n254 ;
  assign n256 = ~x56 & n255 ;
  assign n257 = n253 & n256 ;
  assign n258 = n257 ^ n256 ;
  assign n259 = n258 ^ n255 ;
  assign n260 = ~x0 & ~x51 ;
  assign n261 = n259 & n260 ;
  assign n262 = n261 ^ n259 ;
  assign n263 = n262 ^ n260 ;
  assign n264 = n220 & ~n242 ;
  assign n265 = n264 ^ n220 ;
  assign n266 = x52 & ~x53 ;
  assign n267 = n265 & ~n266 ;
  assign n268 = n263 & n267 ;
  assign n269 = n268 ^ n263 ;
  assign n221 = ~x52 & x53 ;
  assign n270 = ~n221 & ~n265 ;
  assign n204 = x47 & ~n203 ;
  assign n205 = n204 ^ x47 ;
  assign n272 = ~x49 & n205 ;
  assign n273 = n242 & ~n272 ;
  assign n274 = n200 ^ x45 ;
  assign n232 = x41 & ~n192 ;
  assign n233 = n232 ^ x41 ;
  assign n275 = x42 & n233 ;
  assign n276 = x43 & n275 ;
  assign n277 = ~x44 & ~n276 ;
  assign n278 = x36 & x37 ;
  assign n279 = x38 & x41 ;
  assign n280 = n278 & n279 ;
  assign n281 = x32 & x33 ;
  assign n282 = x34 & x35 ;
  assign n283 = n281 & n282 ;
  assign n284 = n280 & n283 ;
  assign n285 = x46 & x47 ;
  assign n286 = n285 ^ x47 ;
  assign n287 = x50 & x56 ;
  assign n288 = n287 ^ x50 ;
  assign n289 = n286 & n288 ;
  assign n290 = n255 & n289 ;
  assign n291 = n284 & n290 ;
  assign n292 = x30 & x31 ;
  assign n293 = n227 & n292 ;
  assign n294 = ~x48 & ~x49 ;
  assign n295 = ~n192 & ~n294 ;
  assign n296 = n293 & n295 ;
  assign n297 = ~n200 & n296 ;
  assign n298 = n291 & n297 ;
  assign n299 = n277 & n298 ;
  assign n300 = n299 ^ n298 ;
  assign n301 = n274 & n300 ;
  assign n308 = n273 & n301 ;
  assign n309 = n308 ^ n301 ;
  assign n310 = n270 & n309 ;
  assign n311 = n310 ^ n309 ;
  assign n312 = n269 & n311 ;
  assign n206 = x48 & ~n203 ;
  assign n207 = ~n205 & ~n206 ;
  assign n208 = ~x46 & ~x51 ;
  assign n209 = ~x56 & x57 ;
  assign n210 = n208 & n209 ;
  assign n211 = x44 & x45 ;
  assign n212 = x41 & ~x43 ;
  assign n213 = n211 & n212 ;
  assign n214 = ~x37 & ~x38 ;
  assign n215 = x39 & ~x40 ;
  assign n216 = n214 & n215 ;
  assign n217 = n213 & n216 ;
  assign n218 = n210 & n217 ;
  assign n219 = x47 & x48 ;
  assign n222 = n220 & n221 ;
  assign n223 = ~n219 & n222 ;
  assign n224 = ~x33 & ~x34 ;
  assign n225 = ~x35 & ~x36 ;
  assign n226 = n224 & n225 ;
  assign n228 = ~x31 & ~x32 ;
  assign n229 = n227 & n228 ;
  assign n230 = n226 & n229 ;
  assign n231 = n223 & n230 ;
  assign n234 = n233 ^ x42 ;
  assign n235 = n231 & n234 ;
  assign n236 = n218 & n235 ;
  assign n237 = ~n207 & n236 ;
  assign n238 = ~x0 & ~x30 ;
  assign n239 = n237 & n238 ;
  assign n271 = n259 & ~n270 ;
  assign n302 = ~n273 & n301 ;
  assign n303 = n271 & n302 ;
  assign n304 = n269 & n303 ;
  assign n305 = n304 ^ n259 ;
  assign n306 = n239 & n305 ;
  assign n307 = n306 ^ n305 ;
  assign n313 = n312 ^ n307 ;
  assign n314 = n313 ^ n95 ;
  assign n315 = ~x24 & n182 ;
  assign n316 = x24 & ~n182 ;
  assign n317 = n155 & ~n316 ;
  assign n318 = ~n315 & n317 ;
  assign n321 = n318 ^ n313 ;
  assign n319 = n318 ^ n128 ;
  assign n320 = n319 ^ n318 ;
  assign n322 = n321 ^ n320 ;
  assign n323 = n321 ^ n318 ;
  assign n324 = n322 & n323 ;
  assign n325 = n324 ^ n322 ;
  assign n326 = n325 ^ n323 ;
  assign n327 = n326 ^ n321 ;
  assign n328 = n314 & ~n327 ;
  assign n329 = n328 ^ n314 ;
  assign n330 = n329 ^ n314 ;
  assign n331 = n330 ^ n313 ;
  assign n332 = n186 ^ n130 ;
  assign n333 = x0 & x30 ;
  assign n334 = n237 & ~n333 ;
  assign n335 = n259 & ~n334 ;
  assign n336 = n335 ^ n130 ;
  assign n337 = ~n335 & ~n336 ;
  assign n338 = n337 ^ n130 ;
  assign n339 = ~n332 & n338 ;
  assign n340 = n339 ^ n337 ;
  assign n341 = n340 ^ n186 ;
  assign y0 = ~n189 ;
  assign y1 = ~n331 ;
  assign y2 = n341 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
