module voting_N_1_M_4_opt( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 ;
  assign n39 = x14 ^ x13 ;
  assign n40 = n39 ^ x15 ;
  assign n49 = n40 ^ x9 ;
  assign n33 = x11 ^ x10 ;
  assign n37 = n33 ^ x12 ;
  assign n50 = n49 ^ n37 ;
  assign n51 = n50 ^ x1 ;
  assign n17 = x7 ^ x6 ;
  assign n24 = n17 ^ x8 ;
  assign n52 = n24 ^ x2 ;
  assign n21 = x4 ^ x3 ;
  assign n22 = n21 ^ x5 ;
  assign n53 = n52 ^ n22 ;
  assign n54 = n53 ^ n50 ;
  assign n55 = n51 & ~n54 ;
  assign n56 = n55 ^ x1 ;
  assign n44 = x15 ^ x14 ;
  assign n45 = n39 & ~n44 ;
  assign n46 = n45 ^ x13 ;
  assign n38 = n37 ^ x9 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n38 & ~n41 ;
  assign n43 = n42 ^ x9 ;
  assign n47 = n46 ^ n43 ;
  assign n34 = x12 ^ x11 ;
  assign n35 = n33 & ~n34 ;
  assign n36 = n35 ^ x10 ;
  assign n48 = n47 ^ n36 ;
  assign n57 = n56 ^ n48 ;
  assign n29 = x5 ^ x3 ;
  assign n30 = n21 & n29 ;
  assign n31 = n30 ^ x3 ;
  assign n23 = n22 ^ x2 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n23 & ~n25 ;
  assign n27 = n26 ^ x2 ;
  assign n18 = x8 ^ x7 ;
  assign n19 = n17 & ~n18 ;
  assign n20 = n19 ^ x6 ;
  assign n28 = n27 ^ n20 ;
  assign n32 = n31 ^ n28 ;
  assign n70 = n56 ^ n32 ;
  assign n71 = n57 & ~n70 ;
  assign n72 = n71 ^ n48 ;
  assign n66 = n46 ^ n36 ;
  assign n67 = n47 & ~n66 ;
  assign n68 = n67 ^ n43 ;
  assign n73 = n72 ^ n68 ;
  assign n62 = n31 ^ n27 ;
  assign n63 = n28 & ~n62 ;
  assign n64 = n63 ^ n20 ;
  assign n58 = n57 ^ n32 ;
  assign n59 = n53 ^ n51 ;
  assign n60 = x0 & n59 ;
  assign n61 = n58 & n60 ;
  assign n65 = n64 ^ n61 ;
  assign n69 = n68 ^ n65 ;
  assign n74 = n73 ^ n69 ;
  assign n75 = n72 ^ n64 ;
  assign n76 = n75 ^ n68 ;
  assign n77 = ~n65 & n75 ;
  assign n78 = n77 ^ n65 ;
  assign n79 = n76 & ~n78 ;
  assign n80 = n79 ^ n68 ;
  assign n81 = n74 & n80 ;
  assign n82 = n81 ^ n77 ;
  assign n83 = n82 ^ n68 ;
  assign n84 = n83 ^ n73 ;
  assign y0 = n84 ;
endmodule
