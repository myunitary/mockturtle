// Benchmark "/tmp/tmp" written by ABC on Wed Nov 12 17:58:22 2025

module FP-lt_opt ( 
    n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
    n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63  );
  input  n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
    n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
    n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63;
  wire new_n129, new_n130, new_n131, new_n132, new_n133, new_n134, new_n135,
    new_n136, new_n137, new_n138, new_n139, new_n140, new_n141, new_n142,
    new_n143, new_n144, new_n145, new_n146, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n182, new_n183, new_n184,
    new_n185, new_n186, new_n187, new_n188, new_n189, new_n190, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771;
  assign new_n129 = n128 ^ n64;
  assign new_n130 = n127 ^ n124;
  assign new_n131 = ~n125 & new_n130;
  assign new_n132 = new_n131 ^ n125;
  assign new_n133 = new_n131 ^ n126;
  assign new_n134 = ~n127 & ~new_n133;
  assign new_n135 = new_n134 ^ n127;
  assign new_n136 = new_n135 ^ n124;
  assign new_n137 = ~new_n132 & new_n136;
  assign new_n138 = ~n62 & ~n63;
  assign new_n139 = ~n60 & ~n61;
  assign new_n140 = new_n138 & new_n139;
  assign new_n141 = new_n137 & new_n140;
  assign new_n142 = n123 ^ n120;
  assign new_n143 = ~n121 & new_n142;
  assign new_n144 = new_n143 ^ n121;
  assign new_n145 = new_n143 ^ n122;
  assign new_n146 = ~n123 & ~new_n145;
  assign new_n147 = new_n146 ^ n123;
  assign new_n148 = new_n147 ^ n120;
  assign new_n149 = ~new_n144 & new_n148;
  assign new_n150 = ~n58 & ~n59;
  assign new_n151 = ~n56 & ~n57;
  assign new_n152 = new_n150 & new_n151;
  assign new_n153 = new_n149 & new_n152;
  assign new_n154 = new_n141 & new_n153;
  assign new_n155 = n119 ^ n116;
  assign new_n156 = ~n117 & new_n155;
  assign new_n157 = new_n156 ^ n117;
  assign new_n158 = new_n156 ^ n118;
  assign new_n159 = ~n119 & ~new_n158;
  assign new_n160 = new_n159 ^ n119;
  assign new_n161 = new_n160 ^ n116;
  assign new_n162 = ~new_n157 & new_n161;
  assign new_n163 = ~n54 & ~n55;
  assign new_n164 = ~n52 & ~n53;
  assign new_n165 = new_n163 & new_n164;
  assign new_n166 = new_n162 & new_n165;
  assign new_n167 = n115 ^ n112;
  assign new_n168 = ~n113 & new_n167;
  assign new_n169 = new_n168 ^ n113;
  assign new_n170 = new_n168 ^ n114;
  assign new_n171 = ~n115 & ~new_n170;
  assign new_n172 = new_n171 ^ n115;
  assign new_n173 = new_n172 ^ n112;
  assign new_n174 = ~new_n169 & new_n173;
  assign new_n175 = ~n50 & ~n51;
  assign new_n176 = ~n48 & ~n49;
  assign new_n177 = new_n175 & new_n176;
  assign new_n178 = new_n174 & new_n177;
  assign new_n179 = new_n166 & new_n178;
  assign new_n180 = new_n154 & new_n179;
  assign new_n181 = n111 ^ n108;
  assign new_n182 = ~n109 & new_n181;
  assign new_n183 = new_n182 ^ n109;
  assign new_n184 = new_n182 ^ n110;
  assign new_n185 = ~n111 & ~new_n184;
  assign new_n186 = new_n185 ^ n111;
  assign new_n187 = new_n186 ^ n108;
  assign new_n188 = ~new_n183 & new_n187;
  assign new_n189 = ~n46 & ~n47;
  assign new_n190 = ~n44 & ~n45;
  assign new_n191 = new_n189 & new_n190;
  assign new_n192 = new_n188 & new_n191;
  assign new_n193 = n107 ^ n104;
  assign new_n194 = ~n105 & new_n193;
  assign new_n195 = new_n194 ^ n105;
  assign new_n196 = new_n194 ^ n106;
  assign new_n197 = ~n107 & ~new_n196;
  assign new_n198 = new_n197 ^ n107;
  assign new_n199 = new_n198 ^ n104;
  assign new_n200 = ~new_n195 & new_n199;
  assign new_n201 = ~n42 & ~n43;
  assign new_n202 = ~n40 & ~n41;
  assign new_n203 = new_n201 & new_n202;
  assign new_n204 = new_n200 & new_n203;
  assign new_n205 = new_n192 & new_n204;
  assign new_n206 = n103 ^ n100;
  assign new_n207 = ~n101 & new_n206;
  assign new_n208 = new_n207 ^ n101;
  assign new_n209 = new_n207 ^ n102;
  assign new_n210 = ~n103 & ~new_n209;
  assign new_n211 = new_n210 ^ n103;
  assign new_n212 = new_n211 ^ n100;
  assign new_n213 = ~new_n208 & new_n212;
  assign new_n214 = ~n38 & ~n39;
  assign new_n215 = ~n36 & ~n37;
  assign new_n216 = new_n214 & new_n215;
  assign new_n217 = new_n213 & new_n216;
  assign new_n218 = n99 ^ n96;
  assign new_n219 = ~n97 & new_n218;
  assign new_n220 = new_n219 ^ n97;
  assign new_n221 = new_n219 ^ n98;
  assign new_n222 = ~n99 & ~new_n221;
  assign new_n223 = new_n222 ^ n99;
  assign new_n224 = new_n223 ^ n96;
  assign new_n225 = ~new_n220 & new_n224;
  assign new_n226 = ~n34 & ~n35;
  assign new_n227 = ~n32 & ~n33;
  assign new_n228 = new_n226 & new_n227;
  assign new_n229 = new_n225 & new_n228;
  assign new_n230 = new_n217 & new_n229;
  assign new_n231 = new_n205 & new_n230;
  assign new_n232 = new_n180 & new_n231;
  assign new_n233 = n95 ^ n92;
  assign new_n234 = ~n93 & new_n233;
  assign new_n235 = new_n234 ^ n93;
  assign new_n236 = new_n234 ^ n94;
  assign new_n237 = ~n95 & ~new_n236;
  assign new_n238 = new_n237 ^ n95;
  assign new_n239 = new_n238 ^ n92;
  assign new_n240 = ~new_n235 & new_n239;
  assign new_n241 = ~n30 & ~n31;
  assign new_n242 = ~n28 & ~n29;
  assign new_n243 = new_n241 & new_n242;
  assign new_n244 = new_n240 & new_n243;
  assign new_n245 = n91 ^ n88;
  assign new_n246 = ~n89 & new_n245;
  assign new_n247 = new_n246 ^ n89;
  assign new_n248 = new_n246 ^ n90;
  assign new_n249 = ~n91 & ~new_n248;
  assign new_n250 = new_n249 ^ n91;
  assign new_n251 = new_n250 ^ n88;
  assign new_n252 = ~new_n247 & new_n251;
  assign new_n253 = ~n26 & ~n27;
  assign new_n254 = ~n24 & ~n25;
  assign new_n255 = new_n253 & new_n254;
  assign new_n256 = new_n252 & new_n255;
  assign new_n257 = new_n244 & new_n256;
  assign new_n258 = n87 ^ n84;
  assign new_n259 = ~n85 & new_n258;
  assign new_n260 = new_n259 ^ n85;
  assign new_n261 = new_n259 ^ n86;
  assign new_n262 = ~n87 & ~new_n261;
  assign new_n263 = new_n262 ^ n87;
  assign new_n264 = new_n263 ^ n84;
  assign new_n265 = ~new_n260 & new_n264;
  assign new_n266 = ~n22 & ~n23;
  assign new_n267 = ~n20 & ~n21;
  assign new_n268 = new_n266 & new_n267;
  assign new_n269 = new_n265 & new_n268;
  assign new_n270 = n83 ^ n80;
  assign new_n271 = ~n81 & new_n270;
  assign new_n272 = new_n271 ^ n81;
  assign new_n273 = new_n271 ^ n82;
  assign new_n274 = ~n83 & ~new_n273;
  assign new_n275 = new_n274 ^ n83;
  assign new_n276 = new_n275 ^ n80;
  assign new_n277 = ~new_n272 & new_n276;
  assign new_n278 = ~n18 & ~n19;
  assign new_n279 = ~n16 & ~n17;
  assign new_n280 = new_n278 & new_n279;
  assign new_n281 = new_n277 & new_n280;
  assign new_n282 = new_n269 & new_n281;
  assign new_n283 = new_n257 & new_n282;
  assign new_n284 = n79 ^ n76;
  assign new_n285 = ~n77 & new_n284;
  assign new_n286 = new_n285 ^ n77;
  assign new_n287 = new_n285 ^ n78;
  assign new_n288 = ~n79 & ~new_n287;
  assign new_n289 = new_n288 ^ n79;
  assign new_n290 = new_n289 ^ n76;
  assign new_n291 = ~new_n286 & new_n290;
  assign new_n292 = ~n14 & ~n15;
  assign new_n293 = ~n12 & ~n13;
  assign new_n294 = new_n292 & new_n293;
  assign new_n295 = new_n291 & new_n294;
  assign new_n296 = n75 ^ n72;
  assign new_n297 = ~n73 & new_n296;
  assign new_n298 = new_n297 ^ n73;
  assign new_n299 = new_n297 ^ n74;
  assign new_n300 = ~n75 & ~new_n299;
  assign new_n301 = new_n300 ^ n75;
  assign new_n302 = new_n301 ^ n72;
  assign new_n303 = ~new_n298 & new_n302;
  assign new_n304 = ~n10 & ~n11;
  assign new_n305 = ~n8 & ~n9;
  assign new_n306 = new_n304 & new_n305;
  assign new_n307 = new_n303 & new_n306;
  assign new_n308 = new_n295 & new_n307;
  assign new_n309 = n71 ^ n68;
  assign new_n310 = ~n69 & new_n309;
  assign new_n311 = new_n310 ^ n69;
  assign new_n312 = new_n310 ^ n70;
  assign new_n313 = ~n71 & ~new_n312;
  assign new_n314 = new_n313 ^ n71;
  assign new_n315 = new_n314 ^ n68;
  assign new_n316 = ~new_n311 & new_n315;
  assign new_n317 = n67 ^ n3;
  assign new_n318 = n66 ^ n2;
  assign new_n319 = ~n1 & n65;
  assign new_n320 = new_n319 ^ n66;
  assign new_n321 = ~new_n318 & ~new_n320;
  assign new_n322 = new_n321 ^ n2;
  assign new_n323 = new_n322 ^ n67;
  assign new_n324 = ~new_n323 & new_n317;
  assign new_n325 = new_n324 ^ new_n322;
  assign new_n326 = ~n1 & ~n2;
  assign new_n327 = ~n3 & new_n326;
  assign new_n328 = ~n6 & ~n7;
  assign new_n329 = ~n4 & ~n5;
  assign new_n330 = new_n328 & new_n329;
  assign new_n331 = new_n327 & new_n330;
  assign new_n332 = new_n325 & new_n331;
  assign new_n333 = new_n316 & new_n332;
  assign new_n334 = new_n308 & new_n333;
  assign new_n335 = new_n283 & new_n334;
  assign new_n336 = new_n232 & new_n335;
  assign new_n337 = ~new_n336 & n64;
  assign new_n338 = n127 ^ n63;
  assign new_n339 = ~new_n129 & ~new_n338;
  assign new_n340 = n126 ^ n62;
  assign new_n341 = n125 ^ n61;
  assign new_n342 = ~new_n340 & ~new_n341;
  assign new_n343 = new_n339 & new_n342;
  assign new_n344 = n124 ^ n60;
  assign new_n345 = n123 ^ n59;
  assign new_n346 = ~new_n344 & ~new_n345;
  assign new_n347 = n122 ^ n58;
  assign new_n348 = n121 ^ n57;
  assign new_n349 = ~new_n347 & ~new_n348;
  assign new_n350 = new_n346 & new_n349;
  assign new_n351 = new_n343 & new_n350;
  assign new_n352 = n120 ^ n56;
  assign new_n353 = n119 ^ n55;
  assign new_n354 = ~new_n352 & ~new_n353;
  assign new_n355 = n118 ^ n54;
  assign new_n356 = n117 ^ n53;
  assign new_n357 = ~new_n355 & ~new_n356;
  assign new_n358 = new_n354 & new_n357;
  assign new_n359 = n116 ^ n52;
  assign new_n360 = n115 ^ n51;
  assign new_n361 = ~new_n359 & ~new_n360;
  assign new_n362 = n114 ^ n50;
  assign new_n363 = n113 ^ n49;
  assign new_n364 = ~new_n362 & ~new_n363;
  assign new_n365 = new_n361 & new_n364;
  assign new_n366 = new_n358 & new_n365;
  assign new_n367 = new_n351 & new_n366;
  assign new_n368 = n112 ^ n48;
  assign new_n369 = n111 ^ n47;
  assign new_n370 = ~new_n368 & ~new_n369;
  assign new_n371 = n110 ^ n46;
  assign new_n372 = n109 ^ n45;
  assign new_n373 = ~new_n371 & ~new_n372;
  assign new_n374 = new_n370 & new_n373;
  assign new_n375 = n108 ^ n44;
  assign new_n376 = n107 ^ n43;
  assign new_n377 = ~new_n375 & ~new_n376;
  assign new_n378 = n106 ^ n42;
  assign new_n379 = n105 ^ n41;
  assign new_n380 = ~new_n378 & ~new_n379;
  assign new_n381 = new_n377 & new_n380;
  assign new_n382 = new_n374 & new_n381;
  assign new_n383 = n104 ^ n40;
  assign new_n384 = n103 ^ n39;
  assign new_n385 = ~new_n383 & ~new_n384;
  assign new_n386 = n102 ^ n38;
  assign new_n387 = n101 ^ n37;
  assign new_n388 = ~new_n386 & ~new_n387;
  assign new_n389 = new_n385 & new_n388;
  assign new_n390 = n100 ^ n36;
  assign new_n391 = n99 ^ n35;
  assign new_n392 = ~new_n390 & ~new_n391;
  assign new_n393 = n98 ^ n34;
  assign new_n394 = n97 ^ n33;
  assign new_n395 = ~new_n393 & ~new_n394;
  assign new_n396 = new_n392 & new_n395;
  assign new_n397 = new_n389 & new_n396;
  assign new_n398 = new_n382 & new_n397;
  assign new_n399 = new_n367 & new_n398;
  assign new_n400 = n96 ^ n32;
  assign new_n401 = n95 ^ n31;
  assign new_n402 = ~new_n400 & ~new_n401;
  assign new_n403 = n94 ^ n30;
  assign new_n404 = n93 ^ n29;
  assign new_n405 = ~new_n403 & ~new_n404;
  assign new_n406 = new_n402 & new_n405;
  assign new_n407 = n92 ^ n28;
  assign new_n408 = n91 ^ n27;
  assign new_n409 = ~new_n407 & ~new_n408;
  assign new_n410 = n90 ^ n26;
  assign new_n411 = n89 ^ n25;
  assign new_n412 = ~new_n410 & ~new_n411;
  assign new_n413 = new_n409 & new_n412;
  assign new_n414 = new_n406 & new_n413;
  assign new_n415 = n88 ^ n24;
  assign new_n416 = n87 ^ n23;
  assign new_n417 = ~new_n415 & ~new_n416;
  assign new_n418 = n86 ^ n22;
  assign new_n419 = n85 ^ n21;
  assign new_n420 = ~new_n418 & ~new_n419;
  assign new_n421 = new_n417 & new_n420;
  assign new_n422 = n84 ^ n20;
  assign new_n423 = n83 ^ n19;
  assign new_n424 = ~new_n422 & ~new_n423;
  assign new_n425 = n82 ^ n18;
  assign new_n426 = n81 ^ n17;
  assign new_n427 = ~new_n425 & ~new_n426;
  assign new_n428 = new_n424 & new_n427;
  assign new_n429 = new_n421 & new_n428;
  assign new_n430 = new_n414 & new_n429;
  assign new_n431 = n80 ^ n16;
  assign new_n432 = n79 ^ n15;
  assign new_n433 = ~new_n431 & ~new_n432;
  assign new_n434 = n78 ^ n14;
  assign new_n435 = n77 ^ n13;
  assign new_n436 = ~new_n434 & ~new_n435;
  assign new_n437 = new_n433 & new_n436;
  assign new_n438 = n76 ^ n12;
  assign new_n439 = n75 ^ n11;
  assign new_n440 = ~new_n438 & ~new_n439;
  assign new_n441 = n74 ^ n10;
  assign new_n442 = n73 ^ n9;
  assign new_n443 = ~new_n441 & ~new_n442;
  assign new_n444 = new_n440 & new_n443;
  assign new_n445 = new_n437 & new_n444;
  assign new_n446 = n72 ^ n8;
  assign new_n447 = n71 ^ n7;
  assign new_n448 = ~new_n446 & ~new_n447;
  assign new_n449 = n70 ^ n6;
  assign new_n450 = n69 ^ n5;
  assign new_n451 = ~new_n449 & ~new_n450;
  assign new_n452 = new_n448 & new_n451;
  assign new_n453 = n68 ^ n4;
  assign new_n454 = ~new_n317 & ~new_n453;
  assign new_n455 = n65 ^ n1;
  assign new_n456 = ~new_n318 & ~new_n455;
  assign new_n457 = new_n454 & new_n456;
  assign new_n458 = new_n452 & new_n457;
  assign new_n459 = new_n445 & new_n458;
  assign new_n460 = new_n430 & new_n459;
  assign new_n461 = new_n399 & new_n460;
  assign new_n462 = new_n325 ^ n68;
  assign new_n463 = ~new_n453 & new_n462;
  assign new_n464 = new_n463 ^ n4;
  assign new_n465 = new_n464 ^ n69;
  assign new_n466 = ~new_n465 & new_n450;
  assign new_n467 = new_n466 ^ new_n464;
  assign new_n468 = new_n467 ^ n70;
  assign new_n469 = ~new_n449 & new_n468;
  assign new_n470 = new_n469 ^ n6;
  assign new_n471 = new_n470 ^ n71;
  assign new_n472 = ~new_n471 & new_n447;
  assign new_n473 = new_n472 ^ new_n470;
  assign new_n474 = new_n473 ^ n72;
  assign new_n475 = ~new_n446 & new_n474;
  assign new_n476 = new_n475 ^ n8;
  assign new_n477 = new_n476 ^ n73;
  assign new_n478 = ~new_n477 & new_n442;
  assign new_n479 = new_n478 ^ new_n476;
  assign new_n480 = new_n479 ^ n74;
  assign new_n481 = ~new_n441 & new_n480;
  assign new_n482 = new_n481 ^ n10;
  assign new_n483 = new_n482 ^ n75;
  assign new_n484 = ~new_n483 & new_n439;
  assign new_n485 = new_n484 ^ new_n482;
  assign new_n486 = new_n485 ^ n76;
  assign new_n487 = ~new_n438 & new_n486;
  assign new_n488 = new_n487 ^ n12;
  assign new_n489 = new_n488 ^ n77;
  assign new_n490 = ~new_n489 & new_n435;
  assign new_n491 = new_n490 ^ new_n488;
  assign new_n492 = new_n491 ^ n78;
  assign new_n493 = ~new_n434 & new_n492;
  assign new_n494 = new_n493 ^ n14;
  assign new_n495 = new_n494 ^ n79;
  assign new_n496 = ~new_n495 & new_n432;
  assign new_n497 = new_n496 ^ new_n494;
  assign new_n498 = new_n497 ^ n80;
  assign new_n499 = ~new_n431 & new_n498;
  assign new_n500 = new_n499 ^ n16;
  assign new_n501 = new_n500 ^ n81;
  assign new_n502 = ~new_n501 & new_n426;
  assign new_n503 = new_n502 ^ new_n500;
  assign new_n504 = new_n503 ^ n82;
  assign new_n505 = ~new_n425 & new_n504;
  assign new_n506 = new_n505 ^ n18;
  assign new_n507 = new_n506 ^ n83;
  assign new_n508 = ~new_n507 & new_n423;
  assign new_n509 = new_n508 ^ new_n506;
  assign new_n510 = new_n509 ^ n84;
  assign new_n511 = ~new_n422 & new_n510;
  assign new_n512 = new_n511 ^ n20;
  assign new_n513 = new_n512 ^ n85;
  assign new_n514 = ~new_n513 & new_n419;
  assign new_n515 = new_n514 ^ new_n512;
  assign new_n516 = new_n515 ^ n86;
  assign new_n517 = ~new_n418 & new_n516;
  assign new_n518 = new_n517 ^ n22;
  assign new_n519 = new_n518 ^ n87;
  assign new_n520 = ~new_n519 & new_n416;
  assign new_n521 = new_n520 ^ new_n518;
  assign new_n522 = new_n521 ^ n88;
  assign new_n523 = ~new_n415 & new_n522;
  assign new_n524 = new_n523 ^ n24;
  assign new_n525 = new_n524 ^ n89;
  assign new_n526 = ~new_n525 & new_n411;
  assign new_n527 = new_n526 ^ new_n524;
  assign new_n528 = new_n527 ^ n90;
  assign new_n529 = ~new_n410 & new_n528;
  assign new_n530 = new_n529 ^ n26;
  assign new_n531 = new_n530 ^ n91;
  assign new_n532 = ~new_n531 & new_n408;
  assign new_n533 = new_n532 ^ new_n530;
  assign new_n534 = new_n533 ^ n92;
  assign new_n535 = ~new_n407 & new_n534;
  assign new_n536 = new_n535 ^ n28;
  assign new_n537 = new_n536 ^ n93;
  assign new_n538 = ~new_n537 & new_n404;
  assign new_n539 = new_n538 ^ new_n536;
  assign new_n540 = new_n539 ^ n94;
  assign new_n541 = ~new_n403 & new_n540;
  assign new_n542 = new_n541 ^ n30;
  assign new_n543 = new_n542 ^ n95;
  assign new_n544 = ~new_n543 & new_n401;
  assign new_n545 = new_n544 ^ new_n542;
  assign new_n546 = new_n545 ^ n96;
  assign new_n547 = ~new_n400 & new_n546;
  assign new_n548 = new_n547 ^ n32;
  assign new_n549 = new_n548 ^ n97;
  assign new_n550 = ~new_n549 & new_n394;
  assign new_n551 = new_n550 ^ new_n548;
  assign new_n552 = new_n551 ^ n98;
  assign new_n553 = ~new_n393 & new_n552;
  assign new_n554 = new_n553 ^ n34;
  assign new_n555 = new_n554 ^ n99;
  assign new_n556 = ~new_n555 & new_n391;
  assign new_n557 = new_n556 ^ new_n554;
  assign new_n558 = new_n557 ^ n100;
  assign new_n559 = ~new_n390 & new_n558;
  assign new_n560 = new_n559 ^ n36;
  assign new_n561 = new_n560 ^ n101;
  assign new_n562 = ~new_n561 & new_n387;
  assign new_n563 = new_n562 ^ new_n560;
  assign new_n564 = new_n563 ^ n102;
  assign new_n565 = ~new_n386 & new_n564;
  assign new_n566 = new_n565 ^ n38;
  assign new_n567 = new_n566 ^ n103;
  assign new_n568 = ~new_n567 & new_n384;
  assign new_n569 = new_n568 ^ new_n566;
  assign new_n570 = new_n569 ^ n104;
  assign new_n571 = ~new_n383 & new_n570;
  assign new_n572 = new_n571 ^ n40;
  assign new_n573 = new_n572 ^ n105;
  assign new_n574 = ~new_n573 & new_n379;
  assign new_n575 = new_n574 ^ new_n572;
  assign new_n576 = new_n575 ^ n106;
  assign new_n577 = ~new_n378 & new_n576;
  assign new_n578 = new_n577 ^ n42;
  assign new_n579 = new_n578 ^ n107;
  assign new_n580 = ~new_n579 & new_n376;
  assign new_n581 = new_n580 ^ new_n578;
  assign new_n582 = new_n581 ^ n108;
  assign new_n583 = ~new_n375 & new_n582;
  assign new_n584 = new_n583 ^ n44;
  assign new_n585 = new_n584 ^ n109;
  assign new_n586 = ~new_n585 & new_n372;
  assign new_n587 = new_n586 ^ new_n584;
  assign new_n588 = new_n587 ^ n110;
  assign new_n589 = ~new_n371 & new_n588;
  assign new_n590 = new_n589 ^ n46;
  assign new_n591 = new_n590 ^ n111;
  assign new_n592 = ~new_n591 & new_n369;
  assign new_n593 = new_n592 ^ new_n590;
  assign new_n594 = new_n593 ^ n112;
  assign new_n595 = ~new_n368 & new_n594;
  assign new_n596 = new_n595 ^ n48;
  assign new_n597 = new_n596 ^ n113;
  assign new_n598 = ~new_n597 & new_n363;
  assign new_n599 = new_n598 ^ new_n596;
  assign new_n600 = new_n599 ^ n114;
  assign new_n601 = ~new_n362 & new_n600;
  assign new_n602 = new_n601 ^ n50;
  assign new_n603 = new_n602 ^ n115;
  assign new_n604 = ~new_n603 & new_n360;
  assign new_n605 = new_n604 ^ new_n602;
  assign new_n606 = new_n605 ^ n116;
  assign new_n607 = ~new_n359 & new_n606;
  assign new_n608 = new_n607 ^ n52;
  assign new_n609 = new_n608 ^ n117;
  assign new_n610 = ~new_n609 & new_n356;
  assign new_n611 = new_n610 ^ new_n608;
  assign new_n612 = new_n611 ^ n118;
  assign new_n613 = ~new_n355 & new_n612;
  assign new_n614 = new_n613 ^ n54;
  assign new_n615 = new_n614 ^ n119;
  assign new_n616 = ~new_n615 & new_n353;
  assign new_n617 = new_n616 ^ new_n614;
  assign new_n618 = new_n617 ^ n120;
  assign new_n619 = ~new_n352 & new_n618;
  assign new_n620 = new_n619 ^ n56;
  assign new_n621 = new_n620 ^ n121;
  assign new_n622 = ~new_n621 & new_n348;
  assign new_n623 = new_n622 ^ new_n620;
  assign new_n624 = new_n623 ^ n122;
  assign new_n625 = ~new_n347 & new_n624;
  assign new_n626 = new_n625 ^ n58;
  assign new_n627 = new_n626 ^ n123;
  assign new_n628 = ~new_n627 & new_n345;
  assign new_n629 = new_n628 ^ new_n626;
  assign new_n630 = new_n629 ^ n124;
  assign new_n631 = ~new_n344 & new_n630;
  assign new_n632 = new_n631 ^ n60;
  assign new_n633 = new_n632 ^ n125;
  assign new_n634 = ~new_n633 & new_n341;
  assign new_n635 = new_n634 ^ new_n632;
  assign new_n636 = new_n635 ^ n126;
  assign new_n637 = ~new_n340 & new_n636;
  assign new_n638 = new_n637 ^ n62;
  assign new_n639 = new_n638 ^ n127;
  assign new_n640 = ~new_n639 & new_n338;
  assign new_n641 = new_n640 ^ new_n638;
  assign new_n642 = new_n641 ^ n128;
  assign new_n643 = ~new_n129 & new_n642;
  assign new_n644 = ~new_n461 & ~new_n643;
  assign new_n645 = new_n644 ^ new_n337;
  assign new_n646 = new_n129 & new_n645;
  assign new_n647 = new_n646 ^ new_n644;
  assign new_n648 = ~n51 & ~n52;
  assign new_n649 = ~n49 & ~n50;
  assign new_n650 = new_n648 & new_n649;
  assign new_n651 = ~n47 & ~n48;
  assign new_n652 = ~n45 & ~n46;
  assign new_n653 = new_n651 & new_n652;
  assign new_n654 = ~n43 & ~n44;
  assign new_n655 = ~n41 & ~n42;
  assign new_n656 = new_n654 & new_n655;
  assign new_n657 = new_n653 & new_n656;
  assign new_n658 = ~n39 & ~n40;
  assign new_n659 = ~n37 & ~n38;
  assign new_n660 = new_n658 & new_n659;
  assign new_n661 = ~n35 & ~n36;
  assign new_n662 = ~n33 & ~n34;
  assign new_n663 = new_n661 & new_n662;
  assign new_n664 = new_n660 & new_n663;
  assign new_n665 = new_n657 & new_n664;
  assign new_n666 = new_n650 & new_n665;
  assign new_n667 = ~n31 & ~n32;
  assign new_n668 = ~n29 & ~n30;
  assign new_n669 = new_n667 & new_n668;
  assign new_n670 = ~n27 & ~n28;
  assign new_n671 = ~n25 & ~n26;
  assign new_n672 = new_n670 & new_n671;
  assign new_n673 = new_n669 & new_n672;
  assign new_n674 = ~n23 & ~n24;
  assign new_n675 = ~n21 & ~n22;
  assign new_n676 = new_n674 & new_n675;
  assign new_n677 = ~n19 & ~n20;
  assign new_n678 = ~n17 & ~n18;
  assign new_n679 = new_n677 & new_n678;
  assign new_n680 = new_n676 & new_n679;
  assign new_n681 = new_n673 & new_n680;
  assign new_n682 = ~n15 & ~n16;
  assign new_n683 = ~n13 & ~n14;
  assign new_n684 = new_n682 & new_n683;
  assign new_n685 = ~n11 & ~n12;
  assign new_n686 = ~n9 & ~n10;
  assign new_n687 = new_n685 & new_n686;
  assign new_n688 = new_n684 & new_n687;
  assign new_n689 = ~n7 & ~n8;
  assign new_n690 = ~n5 & ~n6;
  assign new_n691 = new_n689 & new_n690;
  assign new_n692 = ~n4 & new_n327;
  assign new_n693 = new_n691 & new_n692;
  assign new_n694 = new_n688 & new_n693;
  assign new_n695 = new_n681 & new_n694;
  assign new_n696 = new_n666 & new_n695;
  assign new_n697 = n61 & n62;
  assign new_n698 = n63 & new_n697;
  assign new_n699 = n59 & n60;
  assign new_n700 = n57 & n58;
  assign new_n701 = new_n699 & new_n700;
  assign new_n702 = n53 & n54;
  assign new_n703 = n55 & n56;
  assign new_n704 = new_n702 & new_n703;
  assign new_n705 = new_n701 & new_n704;
  assign new_n706 = new_n698 & new_n705;
  assign new_n707 = ~new_n696 & new_n706;
  assign new_n708 = ~n115 & ~n116;
  assign new_n709 = ~n113 & ~n114;
  assign new_n710 = new_n708 & new_n709;
  assign new_n711 = ~n111 & ~n112;
  assign new_n712 = ~n109 & ~n110;
  assign new_n713 = new_n711 & new_n712;
  assign new_n714 = ~n107 & ~n108;
  assign new_n715 = ~n105 & ~n106;
  assign new_n716 = new_n714 & new_n715;
  assign new_n717 = new_n713 & new_n716;
  assign new_n718 = ~n103 & ~n104;
  assign new_n719 = ~n101 & ~n102;
  assign new_n720 = new_n718 & new_n719;
  assign new_n721 = ~n99 & ~n100;
  assign new_n722 = ~n97 & ~n98;
  assign new_n723 = new_n721 & new_n722;
  assign new_n724 = new_n720 & new_n723;
  assign new_n725 = new_n717 & new_n724;
  assign new_n726 = new_n710 & new_n725;
  assign new_n727 = ~n95 & ~n96;
  assign new_n728 = ~n93 & ~n94;
  assign new_n729 = new_n727 & new_n728;
  assign new_n730 = ~n91 & ~n92;
  assign new_n731 = ~n89 & ~n90;
  assign new_n732 = new_n730 & new_n731;
  assign new_n733 = new_n729 & new_n732;
  assign new_n734 = ~n87 & ~n88;
  assign new_n735 = ~n85 & ~n86;
  assign new_n736 = new_n734 & new_n735;
  assign new_n737 = ~n83 & ~n84;
  assign new_n738 = ~n81 & ~n82;
  assign new_n739 = new_n737 & new_n738;
  assign new_n740 = new_n736 & new_n739;
  assign new_n741 = new_n733 & new_n740;
  assign new_n742 = ~n79 & ~n80;
  assign new_n743 = ~n77 & ~n78;
  assign new_n744 = new_n742 & new_n743;
  assign new_n745 = ~n75 & ~n76;
  assign new_n746 = ~n73 & ~n74;
  assign new_n747 = new_n745 & new_n746;
  assign new_n748 = new_n744 & new_n747;
  assign new_n749 = ~n71 & ~n72;
  assign new_n750 = ~n69 & ~n70;
  assign new_n751 = new_n749 & new_n750;
  assign new_n752 = ~n67 & ~n68;
  assign new_n753 = ~n65 & ~n66;
  assign new_n754 = new_n752 & new_n753;
  assign new_n755 = new_n751 & new_n754;
  assign new_n756 = new_n748 & new_n755;
  assign new_n757 = new_n741 & new_n756;
  assign new_n758 = new_n726 & new_n757;
  assign new_n759 = n125 & n126;
  assign new_n760 = n127 & new_n759;
  assign new_n761 = n123 & n124;
  assign new_n762 = n121 & n122;
  assign new_n763 = new_n761 & new_n762;
  assign new_n764 = n119 & n120;
  assign new_n765 = n117 & n118;
  assign new_n766 = new_n764 & new_n765;
  assign new_n767 = new_n763 & new_n766;
  assign new_n768 = new_n760 & new_n767;
  assign new_n769 = ~new_n758 & new_n768;
  assign new_n770 = ~new_n707 & ~new_n769;
  assign new_n771 = new_n647 & new_n770;
  assign po0 = new_n771;
  assign po1 = 1'b0;
  assign po2 = 1'b0;
  assign po3 = 1'b0;
  assign po4 = 1'b0;
  assign po5 = 1'b0;
  assign po6 = 1'b0;
  assign po7 = 1'b0;
  assign po8 = 1'b0;
  assign po9 = 1'b0;
  assign po10 = 1'b0;
  assign po11 = 1'b0;
  assign po12 = 1'b0;
  assign po13 = 1'b0;
  assign po14 = 1'b0;
  assign po15 = 1'b0;
  assign po16 = 1'b0;
  assign po17 = 1'b0;
  assign po18 = 1'b0;
  assign po19 = 1'b0;
  assign po20 = 1'b0;
  assign po21 = 1'b0;
  assign po22 = 1'b0;
  assign po23 = 1'b0;
  assign po24 = 1'b0;
  assign po25 = 1'b0;
  assign po26 = 1'b0;
  assign po27 = 1'b0;
  assign po28 = 1'b0;
  assign po29 = 1'b0;
  assign po30 = 1'b0;
  assign po31 = 1'b0;
  assign po32 = 1'b0;
  assign po33 = 1'b0;
  assign po34 = 1'b0;
  assign po35 = 1'b0;
  assign po36 = 1'b0;
  assign po37 = 1'b0;
  assign po38 = 1'b0;
  assign po39 = 1'b0;
  assign po40 = 1'b0;
  assign po41 = 1'b0;
  assign po42 = 1'b0;
  assign po43 = 1'b0;
  assign po44 = 1'b0;
  assign po45 = 1'b0;
  assign po46 = 1'b0;
  assign po47 = 1'b0;
  assign po48 = 1'b0;
  assign po49 = 1'b0;
  assign po50 = 1'b0;
  assign po51 = 1'b0;
  assign po52 = 1'b0;
  assign po53 = 1'b0;
  assign po54 = 1'b0;
  assign po55 = 1'b0;
  assign po56 = 1'b0;
  assign po57 = 1'b0;
  assign po58 = 1'b0;
  assign po59 = 1'b0;
  assign po60 = 1'b0;
  assign po61 = 1'b0;
  assign po62 = 1'b0;
  assign po63 = 1'b0;
endmodule


