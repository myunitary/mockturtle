module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 ;
  assign n44 = x25 & x26 ;
  assign n53 = x24 & x25 ;
  assign n253 = n44 & n53 ;
  assign n54 = x22 & x23 ;
  assign n105 = x23 & x24 ;
  assign n254 = n54 & n105 ;
  assign n255 = n253 & n254 ;
  assign n256 = n255 ^ n253 ;
  assign n257 = n256 ^ n254 ;
  assign n45 = x27 & x28 ;
  assign n76 = x26 & x27 ;
  assign n164 = n45 & n76 ;
  assign n73 = x30 & x31 ;
  assign n122 = x29 & x30 ;
  assign n258 = n73 & n122 ;
  assign n259 = n164 & n258 ;
  assign n260 = n259 ^ n258 ;
  assign n261 = n260 ^ n164 ;
  assign n262 = n257 & n261 ;
  assign n263 = n262 ^ n257 ;
  assign n264 = n263 ^ n261 ;
  assign n81 = x9 & x10 ;
  assign n83 = x8 & x9 ;
  assign n185 = n81 & n83 ;
  assign n33 = x13 & x14 ;
  assign n112 = x14 & x15 ;
  assign n265 = n33 & n112 ;
  assign n266 = n185 & n265 ;
  assign n267 = n266 ^ n265 ;
  assign n268 = n267 ^ n185 ;
  assign n74 = x28 & x29 ;
  assign n144 = n74 & n122 ;
  assign n62 = x15 & x16 ;
  assign n269 = n62 & n112 ;
  assign n270 = n144 & n269 ;
  assign n271 = n270 ^ n269 ;
  assign n272 = n271 ^ n144 ;
  assign n273 = ~n268 & ~n272 ;
  assign n274 = ~n264 & n273 ;
  assign n113 = x16 & x17 ;
  assign n235 = n62 & n113 ;
  assign n63 = x17 & x18 ;
  assign n64 = n62 & n63 ;
  assign n236 = n235 ^ n64 ;
  assign n234 = n63 & n113 ;
  assign n237 = n236 ^ n234 ;
  assign n89 = x1 & x2 ;
  assign n220 = ~x0 & ~x3 ;
  assign n238 = n89 & ~n220 ;
  assign n239 = ~n237 & n238 ;
  assign n240 = n239 ^ n237 ;
  assign n241 = n53 & n105 ;
  assign n242 = n44 & n76 ;
  assign n243 = ~n241 & ~n242 ;
  assign n244 = ~n240 & n243 ;
  assign n102 = x20 & x21 ;
  assign n245 = x19 & n102 ;
  assign n246 = n45 & n74 ;
  assign n251 = ~n245 & ~n246 ;
  assign n252 = n244 & n251 ;
  assign n275 = n274 ^ n252 ;
  assign n276 = ~n185 & ~n265 ;
  assign n277 = n276 ^ n272 ;
  assign n278 = ~n276 & ~n277 ;
  assign n279 = n278 ^ n272 ;
  assign n280 = n279 ^ n264 ;
  assign n281 = n264 & n280 ;
  assign n282 = n281 ^ n278 ;
  assign n283 = n282 ^ n272 ;
  assign n284 = ~x17 & x18 ;
  assign n285 = x19 & ~x20 ;
  assign n286 = n284 & n285 ;
  assign n103 = x18 & x19 ;
  assign n287 = n286 ^ n103 ;
  assign n37 = x5 & x6 ;
  assign n84 = x6 & x7 ;
  assign n173 = n37 & n84 ;
  assign n36 = x3 & x4 ;
  assign n91 = x4 & x5 ;
  assign n195 = n36 & n91 ;
  assign n288 = n173 & n195 ;
  assign n289 = n288 ^ n195 ;
  assign n290 = n289 ^ n173 ;
  assign n291 = n287 & n290 ;
  assign n292 = n291 ^ n287 ;
  assign n293 = n292 ^ n290 ;
  assign n106 = x21 & x22 ;
  assign n127 = n54 & n102 ;
  assign n177 = n127 ^ n102 ;
  assign n178 = n177 ^ n54 ;
  assign n294 = n106 & n178 ;
  assign n295 = n293 & n294 ;
  assign n296 = n295 ^ n294 ;
  assign n297 = n296 ^ n293 ;
  assign n34 = x11 & x12 ;
  assign n299 = n34 & n81 ;
  assign n65 = x10 & x11 ;
  assign n298 = n65 & n81 ;
  assign n300 = n299 ^ n298 ;
  assign n148 = n34 & n65 ;
  assign n301 = n300 ^ n148 ;
  assign n66 = x12 & x13 ;
  assign n151 = n33 & n66 ;
  assign n35 = n33 & n34 ;
  assign n303 = n151 ^ n35 ;
  assign n302 = n34 & n66 ;
  assign n304 = n303 ^ n302 ;
  assign n305 = ~n301 & ~n304 ;
  assign n42 = x7 & x8 ;
  assign n306 = n42 & n84 ;
  assign n307 = n37 & n91 ;
  assign n308 = n306 & n307 ;
  assign n309 = n308 ^ n306 ;
  assign n310 = n309 ^ n307 ;
  assign n56 = x2 & x3 ;
  assign n311 = n36 & n56 ;
  assign n312 = x7 & n83 ;
  assign n313 = n311 & n312 ;
  assign n314 = n313 ^ n312 ;
  assign n315 = n314 ^ n311 ;
  assign n316 = n310 & n315 ;
  assign n317 = n316 ^ n310 ;
  assign n318 = n317 ^ n315 ;
  assign n319 = n305 & n318 ;
  assign n320 = n319 ^ n305 ;
  assign n321 = n297 & n320 ;
  assign n322 = n321 ^ n320 ;
  assign n323 = ~n283 & n322 ;
  assign n324 = n323 ^ n283 ;
  assign n325 = n324 ^ n274 ;
  assign n326 = n275 & ~n325 ;
  assign n327 = n326 ^ n275 ;
  assign n328 = n327 ^ n324 ;
  assign n247 = n245 & n246 ;
  assign n248 = n247 ^ n245 ;
  assign n249 = n248 ^ n246 ;
  assign n250 = n244 & ~n249 ;
  assign n329 = n328 ^ n250 ;
  assign n202 = ~x18 & ~x19 ;
  assign n203 = ~x21 & ~x22 ;
  assign n204 = n202 & n203 ;
  assign n205 = ~x14 & ~x15 ;
  assign n206 = ~x16 & ~x17 ;
  assign n207 = n205 & n206 ;
  assign n208 = n204 & n207 ;
  assign n209 = ~x28 & ~x29 ;
  assign n210 = ~x30 & ~x31 ;
  assign n211 = n209 & n210 ;
  assign n212 = ~x23 & ~x24 ;
  assign n213 = ~x25 & ~x27 ;
  assign n214 = n212 & n213 ;
  assign n215 = n211 & n214 ;
  assign n216 = n208 & n215 ;
  assign n217 = ~x1 & ~x2 ;
  assign n218 = ~x4 & ~x5 ;
  assign n219 = n217 & n218 ;
  assign n221 = ~x20 & ~x26 ;
  assign n222 = n220 & n221 ;
  assign n223 = n219 & n222 ;
  assign n224 = ~x10 & ~x11 ;
  assign n225 = ~x12 & ~x13 ;
  assign n226 = n224 & n225 ;
  assign n227 = ~x6 & ~x7 ;
  assign n228 = ~x8 & ~x9 ;
  assign n229 = n227 & n228 ;
  assign n230 = n226 & n229 ;
  assign n231 = n223 & n230 ;
  assign n232 = n216 & n231 ;
  assign n533 = n329 ^ n232 ;
  assign n141 = n56 & n62 ;
  assign n142 = n141 ^ n62 ;
  assign n143 = n142 ^ n56 ;
  assign n145 = n144 ^ n74 ;
  assign n146 = n145 ^ n122 ;
  assign n147 = ~n143 & ~n146 ;
  assign n149 = n148 ^ n34 ;
  assign n150 = n149 ^ n65 ;
  assign n152 = n151 ^ n33 ;
  assign n153 = n152 ^ n66 ;
  assign n154 = ~n150 & ~n153 ;
  assign n155 = n147 & n154 ;
  assign n156 = n73 & n106 ;
  assign n157 = n156 ^ n73 ;
  assign n158 = n157 ^ n106 ;
  assign n159 = n53 & ~n158 ;
  assign n160 = n159 ^ n158 ;
  assign n161 = n44 & n103 ;
  assign n162 = n161 ^ n44 ;
  assign n163 = n162 ^ n103 ;
  assign n165 = n164 ^ n76 ;
  assign n166 = n165 ^ n45 ;
  assign n167 = ~n163 & ~n166 ;
  assign n168 = ~n160 & n167 ;
  assign n169 = n155 & n168 ;
  assign n170 = n105 & n113 ;
  assign n171 = n170 ^ n113 ;
  assign n172 = n171 ^ n105 ;
  assign n174 = n173 ^ n37 ;
  assign n175 = n174 ^ n84 ;
  assign n176 = ~n172 & ~n175 ;
  assign n128 = x19 & x20 ;
  assign n179 = n63 & n128 ;
  assign n180 = n179 ^ n63 ;
  assign n181 = n180 ^ n128 ;
  assign n182 = ~n178 & n181 ;
  assign n183 = n182 ^ n178 ;
  assign n184 = n176 & ~n183 ;
  assign n186 = n185 ^ n81 ;
  assign n187 = n186 ^ n83 ;
  assign n57 = x0 & x1 ;
  assign n188 = n57 & n89 ;
  assign n189 = n188 ^ n89 ;
  assign n190 = n189 ^ n57 ;
  assign n191 = ~n187 & ~n190 ;
  assign n192 = n42 & n112 ;
  assign n193 = n192 ^ n112 ;
  assign n194 = n193 ^ n42 ;
  assign n196 = n195 ^ n36 ;
  assign n197 = n196 ^ n91 ;
  assign n198 = ~n194 & ~n197 ;
  assign n199 = n191 & n198 ;
  assign n200 = n184 & n199 ;
  assign n201 = n169 & n200 ;
  assign n534 = n533 ^ n201 ;
  assign n75 = n73 & n74 ;
  assign n77 = n53 & n76 ;
  assign n78 = n75 & n77 ;
  assign n79 = n78 ^ n75 ;
  assign n80 = n79 ^ n77 ;
  assign n82 = n42 & n81 ;
  assign n85 = n83 & n84 ;
  assign n86 = n82 & n85 ;
  assign n87 = n86 ^ n82 ;
  assign n88 = n87 ^ n85 ;
  assign n90 = n36 & n89 ;
  assign n92 = n56 & n91 ;
  assign n93 = n90 & n92 ;
  assign n94 = n93 ^ n90 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = n88 & n95 ;
  assign n97 = n96 ^ n88 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = n80 & n98 ;
  assign n100 = n99 ^ n80 ;
  assign n101 = n100 ^ n98 ;
  assign n104 = n102 & n103 ;
  assign n107 = n105 & n106 ;
  assign n108 = n104 & n107 ;
  assign n109 = n108 ^ n104 ;
  assign n110 = n109 ^ n107 ;
  assign n111 = n74 & n76 ;
  assign n114 = n112 & n113 ;
  assign n115 = n111 & n114 ;
  assign n116 = n115 ^ n111 ;
  assign n117 = n116 ^ n114 ;
  assign n118 = n110 & n117 ;
  assign n119 = n118 ^ n110 ;
  assign n120 = n119 ^ n117 ;
  assign n121 = n65 & n83 ;
  assign n123 = n45 & n122 ;
  assign n124 = n121 & n123 ;
  assign n125 = n124 ^ n123 ;
  assign n126 = n125 ^ n121 ;
  assign n129 = n106 & n128 ;
  assign n130 = n127 & n129 ;
  assign n131 = n130 ^ n129 ;
  assign n132 = n131 ^ n127 ;
  assign n133 = n126 & n132 ;
  assign n134 = n133 ^ n126 ;
  assign n135 = n134 ^ n132 ;
  assign n136 = n120 & n135 ;
  assign n137 = n136 ^ n120 ;
  assign n138 = n137 ^ n135 ;
  assign n139 = ~n101 & ~n138 ;
  assign n38 = n36 & n37 ;
  assign n39 = n35 & n38 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n40 ^ n38 ;
  assign n43 = n37 & n42 ;
  assign n46 = n44 & n45 ;
  assign n47 = n43 & n46 ;
  assign n48 = n47 ^ n43 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = n41 & n49 ;
  assign n51 = n50 ^ n41 ;
  assign n52 = n51 ^ n49 ;
  assign n55 = n53 & n54 ;
  assign n58 = n56 & n57 ;
  assign n59 = n55 & n58 ;
  assign n60 = n59 ^ n58 ;
  assign n61 = n60 ^ n55 ;
  assign n67 = n65 & n66 ;
  assign n68 = n64 & n67 ;
  assign n69 = n68 ^ n64 ;
  assign n70 = n69 ^ n67 ;
  assign n71 = ~n61 & ~n70 ;
  assign n72 = ~n52 & n71 ;
  assign n338 = n84 & n91 ;
  assign n339 = n103 & n113 ;
  assign n340 = n338 & n339 ;
  assign n341 = n340 ^ n339 ;
  assign n342 = n341 ^ n338 ;
  assign n343 = n103 & n128 ;
  assign n344 = n63 & n343 ;
  assign n345 = ~n342 & n344 ;
  assign n346 = n345 ^ n342 ;
  assign n347 = n33 & n62 ;
  assign n348 = ~n299 & ~n347 ;
  assign n350 = n44 & n105 ;
  assign n351 = n66 & n112 ;
  assign n356 = n350 & n351 ;
  assign n357 = n356 ^ n351 ;
  assign n358 = n357 ^ n350 ;
  assign n535 = n348 & ~n358 ;
  assign n536 = ~n346 & n535 ;
  assign n537 = n72 & n536 ;
  assign n538 = n139 & n537 ;
  assign n539 = n538 ^ n232 ;
  assign n540 = n539 ^ n201 ;
  assign n541 = ~n534 & n540 ;
  assign n542 = n541 ^ n540 ;
  assign n543 = n542 ^ n540 ;
  assign n544 = n543 ^ n538 ;
  assign n532 = ~n201 & ~n232 ;
  assign n545 = n544 ^ n532 ;
  assign n546 = n545 ^ n534 ;
  assign n371 = n37 & n85 ;
  assign n372 = n307 & n311 ;
  assign n373 = n288 & n372 ;
  assign n374 = n373 ^ n288 ;
  assign n375 = n374 ^ n372 ;
  assign n376 = n371 & n375 ;
  assign n377 = n376 ^ n371 ;
  assign n378 = n377 ^ n375 ;
  assign n379 = n57 & n90 ;
  assign n380 = n82 & n306 ;
  assign n381 = ~n379 & ~n380 ;
  assign n382 = n378 & n381 ;
  assign n383 = n382 ^ n381 ;
  assign n384 = n148 & n185 ;
  assign n385 = n265 & n302 ;
  assign n386 = n384 & n385 ;
  assign n387 = n386 ^ n384 ;
  assign n388 = n387 ^ n385 ;
  assign n389 = n242 & n246 ;
  assign n390 = n164 & n253 ;
  assign n391 = n389 & n390 ;
  assign n392 = n391 ^ n389 ;
  assign n393 = n392 ^ n390 ;
  assign n394 = n388 & n393 ;
  assign n395 = n394 ^ n388 ;
  assign n396 = n395 ^ n393 ;
  assign n397 = n56 & n89 ;
  assign n398 = n195 & n397 ;
  assign n399 = n298 & n312 ;
  assign n400 = n398 & n399 ;
  assign n401 = n400 ^ n398 ;
  assign n402 = n401 ^ n399 ;
  assign n403 = n298 & n302 ;
  assign n404 = n308 & n403 ;
  assign n405 = n404 ^ n308 ;
  assign n406 = n405 ^ n403 ;
  assign n407 = n402 & n406 ;
  assign n408 = n407 ^ n402 ;
  assign n409 = n408 ^ n406 ;
  assign n410 = ~n396 & ~n409 ;
  assign n411 = n383 & n410 ;
  assign n412 = n54 & n106 ;
  assign n413 = n241 & n412 ;
  assign n414 = n148 & n151 ;
  assign n415 = n413 & n414 ;
  assign n416 = n415 ^ n413 ;
  assign n417 = n416 ^ n414 ;
  assign n418 = n234 & n269 ;
  assign n419 = n245 & n412 ;
  assign n420 = n418 & n419 ;
  assign n421 = n420 ^ n418 ;
  assign n422 = n421 ^ n419 ;
  assign n423 = ~n417 & ~n422 ;
  assign n424 = n63 & n103 ;
  assign n425 = n235 & n424 ;
  assign n426 = n151 & n269 ;
  assign n427 = n425 & n426 ;
  assign n428 = n427 ^ n425 ;
  assign n429 = n428 ^ n426 ;
  assign n430 = n235 & n265 ;
  assign n431 = n234 & n343 ;
  assign n432 = n430 & n431 ;
  assign n433 = n432 ^ n430 ;
  assign n434 = n433 ^ n431 ;
  assign n435 = ~n429 & ~n434 ;
  assign n436 = n423 & n435 ;
  assign n437 = n241 & n242 ;
  assign n438 = n45 & n75 ;
  assign n439 = n437 & n438 ;
  assign n440 = n439 ^ n437 ;
  assign n441 = n440 ^ n438 ;
  assign n442 = n76 & n123 ;
  assign n443 = n255 & n442 ;
  assign n444 = n443 ^ n255 ;
  assign n445 = n444 ^ n442 ;
  assign n446 = ~n441 & n445 ;
  assign n447 = n446 ^ n441 ;
  assign n448 = n102 & n107 ;
  assign n449 = n63 & n104 ;
  assign n450 = n129 & n343 ;
  assign n451 = n449 & n450 ;
  assign n452 = n451 ^ n449 ;
  assign n453 = n452 ^ n450 ;
  assign n454 = n448 & ~n453 ;
  assign n455 = n454 ^ n453 ;
  assign n456 = ~n447 & ~n455 ;
  assign n457 = n436 & n456 ;
  assign n458 = n411 & n457 ;
  assign n349 = ~n346 & n348 ;
  assign n352 = ~n350 & ~n351 ;
  assign n353 = n349 & n352 ;
  assign n331 = ~n61 & ~n64 ;
  assign n332 = ~n52 & n67 ;
  assign n333 = n332 ^ n52 ;
  assign n334 = n331 & ~n333 ;
  assign n335 = n139 & n334 ;
  assign n336 = n335 ^ n334 ;
  assign n337 = n336 ^ n139 ;
  assign n354 = n353 ^ n337 ;
  assign n355 = n354 ^ n72 ;
  assign n360 = n358 ^ n349 ;
  assign n361 = n358 & n360 ;
  assign n362 = n361 ^ n360 ;
  assign n363 = n362 ^ n358 ;
  assign n359 = n358 ^ n139 ;
  assign n364 = n363 ^ n359 ;
  assign n365 = n355 & ~n364 ;
  assign n366 = n365 ^ n355 ;
  assign n367 = n366 ^ n364 ;
  assign n368 = n367 ^ n337 ;
  assign n233 = n232 ^ n201 ;
  assign n330 = n329 ^ n233 ;
  assign n369 = n368 ^ n330 ;
  assign n140 = n139 ^ n72 ;
  assign n370 = n369 ^ n140 ;
  assign n459 = n458 ^ n370 ;
  assign n460 = n38 & n397 ;
  assign n461 = n46 & n241 ;
  assign n462 = n460 & n461 ;
  assign n463 = n462 ^ n460 ;
  assign n464 = n463 ^ n461 ;
  assign n465 = n77 & n254 ;
  assign n466 = n148 & n351 ;
  assign n467 = n465 & n466 ;
  assign n468 = n467 ^ n465 ;
  assign n469 = n468 ^ n466 ;
  assign n470 = ~n464 & ~n469 ;
  assign n471 = n35 & n298 ;
  assign n472 = n302 & n347 ;
  assign n473 = n471 & n472 ;
  assign n474 = n473 ^ n471 ;
  assign n475 = n474 ^ n472 ;
  assign n476 = n104 & n234 ;
  assign n477 = n179 & n235 ;
  assign n478 = n476 & n477 ;
  assign n479 = n478 ^ n476 ;
  assign n480 = n479 ^ n477 ;
  assign n481 = ~n475 & ~n480 ;
  assign n482 = n470 & n481 ;
  assign n483 = n82 & n371 ;
  assign n484 = n92 & n379 ;
  assign n485 = n483 & n484 ;
  assign n486 = n485 ^ n483 ;
  assign n487 = n486 ^ n484 ;
  assign n488 = n221 & n413 ;
  assign n489 = n488 ^ n413 ;
  assign n490 = ~x13 & ~x19 ;
  assign n491 = n418 & n490 ;
  assign n492 = n491 ^ n418 ;
  assign n493 = n489 & n492 ;
  assign n494 = n493 ^ n489 ;
  assign n495 = n494 ^ n492 ;
  assign n496 = n107 & n245 ;
  assign n497 = n123 & n242 ;
  assign n498 = n496 & n497 ;
  assign n499 = n498 ^ n496 ;
  assign n500 = n499 ^ n497 ;
  assign n501 = n495 & n500 ;
  assign n502 = n501 ^ n495 ;
  assign n503 = n502 ^ n500 ;
  assign n504 = ~n487 & ~n503 ;
  assign n505 = n482 & n504 ;
  assign n506 = n129 & n449 ;
  assign n507 = n80 & n111 ;
  assign n508 = n66 & ~n114 ;
  assign n509 = ~n384 & n508 ;
  assign n510 = n509 ^ n66 ;
  assign n511 = n507 & n510 ;
  assign n512 = n511 ^ n507 ;
  assign n513 = n512 ^ n510 ;
  assign n514 = n506 & ~n513 ;
  assign n515 = n514 ^ n513 ;
  assign n516 = n43 & n195 ;
  assign n517 = n85 & n307 ;
  assign n518 = ~n516 & ~n517 ;
  assign n519 = n311 & n338 ;
  assign n520 = n299 & n312 ;
  assign n521 = ~n519 & ~n520 ;
  assign n522 = n518 & n521 ;
  assign n523 = n121 & n380 ;
  assign n524 = n127 & n450 ;
  assign n525 = ~n523 & ~n524 ;
  assign n526 = n522 & n525 ;
  assign n527 = ~n515 & n526 ;
  assign n528 = n505 & n527 ;
  assign n529 = n528 ^ n370 ;
  assign n530 = n459 & n529 ;
  assign n531 = n530 ^ n370 ;
  assign n547 = n546 ^ n531 ;
  assign n548 = n379 & n460 ;
  assign n549 = n425 & n476 ;
  assign n550 = n163 & n448 ;
  assign n551 = ~n549 & ~n550 ;
  assign n552 = ~n548 & n551 ;
  assign n553 = ~n76 & ~n128 ;
  assign n554 = n413 & ~n553 ;
  assign n555 = ~n34 & ~n103 ;
  assign n556 = n430 & n555 ;
  assign n557 = n556 ^ n430 ;
  assign n558 = ~n106 & ~n112 ;
  assign n559 = n431 & n558 ;
  assign n560 = n559 ^ n431 ;
  assign n561 = n557 & n560 ;
  assign n562 = n561 ^ n557 ;
  assign n563 = n562 ^ n560 ;
  assign n564 = n554 & n563 ;
  assign n565 = n564 ^ n554 ;
  assign n566 = n565 ^ n563 ;
  assign n567 = n372 & n516 ;
  assign n568 = ~n63 & ~n65 ;
  assign n569 = n426 & n568 ;
  assign n570 = n569 ^ n426 ;
  assign n571 = ~n194 & n403 ;
  assign n572 = n571 ^ n403 ;
  assign n573 = n570 & n572 ;
  assign n574 = n573 ^ n570 ;
  assign n575 = n574 ^ n572 ;
  assign n576 = n567 & n575 ;
  assign n577 = n576 ^ n567 ;
  assign n578 = n577 ^ n575 ;
  assign n579 = n566 & n578 ;
  assign n580 = n579 ^ n566 ;
  assign n581 = n580 ^ n578 ;
  assign n582 = n552 & ~n581 ;
  assign n583 = n308 & n483 ;
  assign n584 = n288 & n517 ;
  assign n585 = n398 & n519 ;
  assign n586 = n584 & n585 ;
  assign n587 = n586 ^ n584 ;
  assign n588 = n587 ^ n585 ;
  assign n589 = n583 & n588 ;
  assign n590 = n589 ^ n583 ;
  assign n591 = n590 ^ n588 ;
  assign n592 = n37 & n83 ;
  assign n593 = n65 & n84 ;
  assign n594 = n592 & n593 ;
  assign n595 = n380 & n594 ;
  assign n596 = n380 & n520 ;
  assign n597 = n384 & n471 ;
  assign n598 = n596 & n597 ;
  assign n599 = n598 ^ n596 ;
  assign n600 = n599 ^ n597 ;
  assign n601 = n595 & n600 ;
  assign n602 = n601 ^ n595 ;
  assign n603 = n602 ^ n600 ;
  assign n604 = n591 & n603 ;
  assign n605 = n604 ^ n591 ;
  assign n606 = n605 ^ n603 ;
  assign n607 = n389 & n441 ;
  assign n608 = n390 & n445 ;
  assign n609 = n608 ^ n390 ;
  assign n610 = n609 ^ n390 ;
  assign n611 = n63 & n102 ;
  assign n612 = n54 & n103 ;
  assign n613 = n611 & n612 ;
  assign n614 = n450 & n613 ;
  assign n615 = n610 & n614 ;
  assign n616 = n615 ^ n610 ;
  assign n617 = n616 ^ n614 ;
  assign n618 = n607 & n617 ;
  assign n619 = n618 ^ n607 ;
  assign n620 = n619 ^ n617 ;
  assign n621 = ~n606 & n620 ;
  assign n622 = n621 ^ n606 ;
  assign n623 = n582 & ~n622 ;
  assign n624 = n528 ^ n459 ;
  assign n625 = n623 & n624 ;
  assign n626 = n625 ^ n623 ;
  assign n627 = n626 ^ n624 ;
  assign n628 = ~n547 & n627 ;
  assign n629 = n628 ^ n547 ;
  assign n660 = n370 & n458 ;
  assign n661 = n660 ^ n458 ;
  assign n662 = n661 ^ n370 ;
  assign n678 = n201 & n232 ;
  assign n679 = n678 ^ n232 ;
  assign n686 = ~n329 & n679 ;
  assign n687 = n686 ^ n679 ;
  assign n688 = n662 & n687 ;
  assign n689 = n537 & n688 ;
  assign n690 = n689 ^ n688 ;
  assign n680 = n139 & n679 ;
  assign n681 = n680 ^ n679 ;
  assign n682 = ~n329 & n681 ;
  assign n683 = n682 ^ n681 ;
  assign n684 = n662 & n683 ;
  assign n685 = n537 & n684 ;
  assign n691 = n690 ^ n685 ;
  assign n673 = n201 & ~n329 ;
  assign n674 = n662 & n673 ;
  assign n675 = n537 & n674 ;
  assign n676 = n675 ^ n674 ;
  assign n669 = ~n139 & n201 ;
  assign n670 = ~n329 & n669 ;
  assign n671 = n662 & n670 ;
  assign n672 = n537 & n671 ;
  assign n677 = n676 ^ n672 ;
  assign n692 = n691 ^ n677 ;
  assign n664 = n139 & n232 ;
  assign n665 = n536 & n664 ;
  assign n666 = n72 & n665 ;
  assign n667 = n662 & n666 ;
  assign n663 = n232 & n662 ;
  assign n668 = n667 ^ n663 ;
  assign n693 = n692 ^ n668 ;
  assign n656 = n233 & n329 ;
  assign n657 = ~n532 & n656 ;
  assign n643 = n546 ^ n370 ;
  assign n644 = ~n546 & ~n643 ;
  assign n645 = n644 ^ n643 ;
  assign n630 = n436 & ~n447 ;
  assign n631 = n630 ^ n411 ;
  assign n639 = n630 ^ n546 ;
  assign n632 = n630 ^ n370 ;
  assign n633 = n630 ^ n455 ;
  assign n634 = n633 ^ n370 ;
  assign n635 = n632 & ~n634 ;
  assign n636 = n635 ^ n632 ;
  assign n637 = n636 ^ n634 ;
  assign n638 = n637 ^ n455 ;
  assign n640 = n639 ^ n638 ;
  assign n641 = n631 & n640 ;
  assign n642 = n641 ^ n631 ;
  assign n646 = n645 ^ n642 ;
  assign n647 = n646 ^ n637 ;
  assign n648 = n647 ^ n634 ;
  assign n649 = n645 ^ n546 ;
  assign n650 = n648 & n649 ;
  assign n651 = n650 ^ n648 ;
  assign n652 = n651 ^ n649 ;
  assign n653 = n652 ^ n645 ;
  assign n654 = n653 ^ n546 ;
  assign n655 = n654 ^ n546 ;
  assign n658 = n657 ^ n655 ;
  assign n659 = n658 ^ n532 ;
  assign n694 = n693 ^ n659 ;
  assign n695 = ~n629 & n694 ;
  assign n696 = n695 ^ n629 ;
  assign n697 = n696 ^ n694 ;
  assign n698 = n624 ^ n623 ;
  assign n699 = n607 & n610 ;
  assign n700 = n477 & n570 ;
  assign n701 = n700 ^ n477 ;
  assign n702 = n701 ^ n570 ;
  assign n703 = n557 & ~n702 ;
  assign n704 = n703 ^ n557 ;
  assign n705 = n549 & n560 ;
  assign n706 = n704 & n705 ;
  assign n707 = n706 ^ n704 ;
  assign n708 = n707 ^ n705 ;
  assign n709 = n699 & ~n708 ;
  assign n710 = n709 ^ n708 ;
  assign n711 = n172 & n614 ;
  assign n712 = ~n461 & ~n550 ;
  assign n713 = n554 & ~n712 ;
  assign n714 = ~n711 & ~n713 ;
  assign n715 = ~n710 & n714 ;
  assign n716 = ~n472 & ~n600 ;
  assign n717 = n572 & ~n716 ;
  assign n718 = ~n487 & n567 ;
  assign n719 = n718 ^ n487 ;
  assign n720 = n588 & ~n719 ;
  assign n721 = n720 ^ n588 ;
  assign n722 = n596 ^ n595 ;
  assign n723 = ~n595 & n722 ;
  assign n724 = n723 ^ n595 ;
  assign n725 = n724 ^ n583 ;
  assign n726 = n596 ^ n583 ;
  assign n727 = n725 & n726 ;
  assign n728 = n727 ^ n723 ;
  assign n729 = n728 ^ n583 ;
  assign n730 = n721 & n729 ;
  assign n731 = n730 ^ n721 ;
  assign n732 = n731 ^ n729 ;
  assign n733 = n717 & ~n732 ;
  assign n734 = n733 ^ n732 ;
  assign n735 = n715 & ~n734 ;
  assign n736 = n698 & n735 ;
  assign n737 = n736 ^ n698 ;
  assign n738 = ~n547 & n737 ;
  assign n739 = ~n697 & n738 ;
  assign n740 = n459 & ~n546 ;
  assign n741 = n740 ^ n459 ;
  assign n742 = n528 & n741 ;
  assign n743 = n742 ^ n741 ;
  assign n744 = n694 & n743 ;
  assign n745 = n744 ^ n743 ;
  assign n752 = ~n547 & n735 ;
  assign n753 = n752 ^ n547 ;
  assign n754 = n753 ^ n735 ;
  assign n755 = n698 & n754 ;
  assign n746 = n459 & n528 ;
  assign n747 = n746 ^ n459 ;
  assign n748 = ~n546 & n747 ;
  assign n749 = n748 ^ n747 ;
  assign n750 = n749 ^ n745 ;
  assign n751 = n750 ^ n737 ;
  assign n756 = n755 ^ n751 ;
  assign n757 = n745 & n756 ;
  assign n758 = n757 ^ n756 ;
  assign n759 = n758 ^ n750 ;
  assign n760 = n759 ^ n749 ;
  assign n761 = n760 ^ n750 ;
  assign n762 = n761 ^ n697 ;
  assign n763 = n735 ^ n624 ;
  assign n764 = n698 & n763 ;
  assign n765 = n764 ^ n624 ;
  assign n766 = n765 ^ n547 ;
  assign n767 = ~n698 & ~n735 ;
  assign n768 = ~n736 & ~n767 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = 1'b0 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = n739 ;
  assign y29 = ~n762 ;
  assign y30 = n766 ;
  assign y31 = ~n768 ;
endmodule
