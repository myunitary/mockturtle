module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 ;
  assign n129 = ~x95 & x127 ;
  assign n130 = x95 & ~x127 ;
  assign n131 = ~x94 & x126 ;
  assign n132 = x94 & ~x126 ;
  assign n133 = ~x93 & x125 ;
  assign n134 = x93 & ~x125 ;
  assign n135 = ~x92 & x124 ;
  assign n136 = x92 & ~x124 ;
  assign n137 = ~x91 & x123 ;
  assign n138 = x91 & ~x123 ;
  assign n139 = ~x90 & x122 ;
  assign n140 = x90 & ~x122 ;
  assign n141 = ~x89 & x121 ;
  assign n142 = x89 & ~x121 ;
  assign n143 = ~x88 & x120 ;
  assign n144 = x88 & ~x120 ;
  assign n145 = ~x87 & x119 ;
  assign n146 = x87 & ~x119 ;
  assign n147 = ~x86 & x118 ;
  assign n148 = x86 & ~x118 ;
  assign n149 = ~x85 & x117 ;
  assign n150 = x85 & ~x117 ;
  assign n151 = ~x84 & x116 ;
  assign n152 = x84 & ~x116 ;
  assign n153 = ~x83 & x115 ;
  assign n154 = x83 & ~x115 ;
  assign n155 = ~x82 & x114 ;
  assign n156 = x82 & ~x114 ;
  assign n157 = ~x81 & x113 ;
  assign n158 = x81 & ~x113 ;
  assign n159 = ~x80 & x112 ;
  assign n160 = x80 & ~x112 ;
  assign n161 = ~x79 & x111 ;
  assign n162 = x79 & ~x111 ;
  assign n163 = ~x78 & x110 ;
  assign n164 = x78 & ~x110 ;
  assign n165 = ~x77 & x109 ;
  assign n166 = x77 & ~x109 ;
  assign n167 = ~x76 & x108 ;
  assign n168 = x76 & ~x108 ;
  assign n169 = ~x75 & x107 ;
  assign n170 = x75 & ~x107 ;
  assign n171 = ~x74 & x106 ;
  assign n172 = x74 & ~x106 ;
  assign n173 = ~x73 & x105 ;
  assign n174 = x73 & ~x105 ;
  assign n175 = ~x72 & x104 ;
  assign n176 = x72 & ~x104 ;
  assign n177 = ~x71 & x103 ;
  assign n178 = x71 & ~x103 ;
  assign n179 = ~x70 & x102 ;
  assign n180 = x70 & ~x102 ;
  assign n181 = ~x69 & x101 ;
  assign n182 = x69 & ~x101 ;
  assign n183 = ~x68 & x100 ;
  assign n184 = x68 & ~x100 ;
  assign n185 = ~x67 & x99 ;
  assign n186 = x67 & ~x99 ;
  assign n187 = ~x66 & x98 ;
  assign n188 = x66 & ~x98 ;
  assign n189 = ~x65 & x97 ;
  assign n190 = x65 & ~x97 ;
  assign n191 = x64 & ~x96 ;
  assign n192 = ~n190 & ~n191 ;
  assign n193 = ~n189 & ~n192 ;
  assign n194 = ~n188 & ~n193 ;
  assign n195 = ~n187 & ~n194 ;
  assign n196 = ~n186 & ~n195 ;
  assign n197 = ~n185 & ~n196 ;
  assign n198 = ~n184 & ~n197 ;
  assign n199 = ~n183 & ~n198 ;
  assign n200 = ~n182 & ~n199 ;
  assign n201 = ~n181 & ~n200 ;
  assign n202 = ~n180 & ~n201 ;
  assign n203 = ~n179 & ~n202 ;
  assign n204 = ~n178 & ~n203 ;
  assign n205 = ~n177 & ~n204 ;
  assign n206 = ~n176 & ~n205 ;
  assign n207 = ~n175 & ~n206 ;
  assign n208 = ~n174 & ~n207 ;
  assign n209 = ~n173 & ~n208 ;
  assign n210 = ~n172 & ~n209 ;
  assign n211 = ~n171 & ~n210 ;
  assign n212 = ~n170 & ~n211 ;
  assign n213 = ~n169 & ~n212 ;
  assign n214 = ~n168 & ~n213 ;
  assign n215 = ~n167 & ~n214 ;
  assign n216 = ~n166 & ~n215 ;
  assign n217 = ~n165 & ~n216 ;
  assign n218 = ~n164 & ~n217 ;
  assign n219 = ~n163 & ~n218 ;
  assign n220 = ~n162 & ~n219 ;
  assign n221 = ~n161 & ~n220 ;
  assign n222 = ~n160 & ~n221 ;
  assign n223 = ~n159 & ~n222 ;
  assign n224 = ~n158 & ~n223 ;
  assign n225 = ~n157 & ~n224 ;
  assign n226 = ~n156 & ~n225 ;
  assign n227 = ~n155 & ~n226 ;
  assign n228 = ~n154 & ~n227 ;
  assign n229 = ~n153 & ~n228 ;
  assign n230 = ~n152 & ~n229 ;
  assign n231 = ~n151 & ~n230 ;
  assign n232 = ~n150 & ~n231 ;
  assign n233 = ~n149 & ~n232 ;
  assign n234 = ~n148 & ~n233 ;
  assign n235 = ~n147 & ~n234 ;
  assign n236 = ~n146 & ~n235 ;
  assign n237 = ~n145 & ~n236 ;
  assign n238 = ~n144 & ~n237 ;
  assign n239 = ~n143 & ~n238 ;
  assign n240 = ~n142 & ~n239 ;
  assign n241 = ~n141 & ~n240 ;
  assign n242 = ~n140 & ~n241 ;
  assign n243 = ~n139 & ~n242 ;
  assign n244 = ~n138 & ~n243 ;
  assign n245 = ~n137 & ~n244 ;
  assign n246 = ~n136 & ~n245 ;
  assign n247 = ~n135 & ~n246 ;
  assign n248 = ~n134 & ~n247 ;
  assign n249 = ~n133 & ~n248 ;
  assign n250 = ~n132 & ~n249 ;
  assign n251 = ~n131 & ~n250 ;
  assign n252 = ~n130 & ~n251 ;
  assign n253 = ~n129 & ~n252 ;
  assign n254 = ~x95 & ~x127 ;
  assign n255 = ~x31 & ~x63 ;
  assign n256 = ~n254 & n255 ;
  assign n257 = n254 & ~n255 ;
  assign n258 = x126 & ~n253 ;
  assign n259 = x94 & n253 ;
  assign n260 = ~n258 & ~n259 ;
  assign n261 = ~x31 & x63 ;
  assign n262 = x31 & ~x63 ;
  assign n263 = ~x30 & x62 ;
  assign n264 = x30 & ~x62 ;
  assign n265 = ~x29 & x61 ;
  assign n266 = x29 & ~x61 ;
  assign n267 = ~x28 & x60 ;
  assign n268 = x28 & ~x60 ;
  assign n269 = ~x27 & x59 ;
  assign n270 = x27 & ~x59 ;
  assign n271 = ~x26 & x58 ;
  assign n272 = x26 & ~x58 ;
  assign n273 = ~x25 & x57 ;
  assign n274 = x25 & ~x57 ;
  assign n275 = ~x24 & x56 ;
  assign n276 = x24 & ~x56 ;
  assign n277 = ~x23 & x55 ;
  assign n278 = x23 & ~x55 ;
  assign n279 = ~x22 & x54 ;
  assign n280 = x22 & ~x54 ;
  assign n281 = ~x21 & x53 ;
  assign n282 = x21 & ~x53 ;
  assign n283 = ~x20 & x52 ;
  assign n284 = x20 & ~x52 ;
  assign n285 = ~x19 & x51 ;
  assign n286 = x19 & ~x51 ;
  assign n287 = ~x18 & x50 ;
  assign n288 = x18 & ~x50 ;
  assign n289 = ~x17 & x49 ;
  assign n290 = x17 & ~x49 ;
  assign n291 = ~x16 & x48 ;
  assign n292 = x16 & ~x48 ;
  assign n293 = ~x15 & x47 ;
  assign n294 = x15 & ~x47 ;
  assign n295 = ~x14 & x46 ;
  assign n296 = x14 & ~x46 ;
  assign n297 = ~x13 & x45 ;
  assign n298 = x13 & ~x45 ;
  assign n299 = ~x12 & x44 ;
  assign n300 = x12 & ~x44 ;
  assign n301 = ~x11 & x43 ;
  assign n302 = x11 & ~x43 ;
  assign n303 = ~x10 & x42 ;
  assign n304 = x10 & ~x42 ;
  assign n305 = ~x9 & x41 ;
  assign n306 = x9 & ~x41 ;
  assign n307 = ~x8 & x40 ;
  assign n308 = x8 & ~x40 ;
  assign n309 = ~x7 & x39 ;
  assign n310 = x7 & ~x39 ;
  assign n311 = ~x6 & x38 ;
  assign n312 = x6 & ~x38 ;
  assign n313 = ~x5 & x37 ;
  assign n314 = x5 & ~x37 ;
  assign n315 = ~x4 & x36 ;
  assign n316 = x4 & ~x36 ;
  assign n317 = ~x3 & x35 ;
  assign n318 = x3 & ~x35 ;
  assign n319 = ~x2 & x34 ;
  assign n320 = x2 & ~x34 ;
  assign n321 = ~x1 & x33 ;
  assign n322 = x1 & ~x33 ;
  assign n323 = x0 & ~x32 ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = ~n321 & ~n324 ;
  assign n326 = ~n320 & ~n325 ;
  assign n327 = ~n319 & ~n326 ;
  assign n328 = ~n318 & ~n327 ;
  assign n329 = ~n317 & ~n328 ;
  assign n330 = ~n316 & ~n329 ;
  assign n331 = ~n315 & ~n330 ;
  assign n332 = ~n314 & ~n331 ;
  assign n333 = ~n313 & ~n332 ;
  assign n334 = ~n312 & ~n333 ;
  assign n335 = ~n311 & ~n334 ;
  assign n336 = ~n310 & ~n335 ;
  assign n337 = ~n309 & ~n336 ;
  assign n338 = ~n308 & ~n337 ;
  assign n339 = ~n307 & ~n338 ;
  assign n340 = ~n306 & ~n339 ;
  assign n341 = ~n305 & ~n340 ;
  assign n342 = ~n304 & ~n341 ;
  assign n343 = ~n303 & ~n342 ;
  assign n344 = ~n302 & ~n343 ;
  assign n345 = ~n301 & ~n344 ;
  assign n346 = ~n300 & ~n345 ;
  assign n347 = ~n299 & ~n346 ;
  assign n348 = ~n298 & ~n347 ;
  assign n349 = ~n297 & ~n348 ;
  assign n350 = ~n296 & ~n349 ;
  assign n351 = ~n295 & ~n350 ;
  assign n352 = ~n294 & ~n351 ;
  assign n353 = ~n293 & ~n352 ;
  assign n354 = ~n292 & ~n353 ;
  assign n355 = ~n291 & ~n354 ;
  assign n356 = ~n290 & ~n355 ;
  assign n357 = ~n289 & ~n356 ;
  assign n358 = ~n288 & ~n357 ;
  assign n359 = ~n287 & ~n358 ;
  assign n360 = ~n286 & ~n359 ;
  assign n361 = ~n285 & ~n360 ;
  assign n362 = ~n284 & ~n361 ;
  assign n363 = ~n283 & ~n362 ;
  assign n364 = ~n282 & ~n363 ;
  assign n365 = ~n281 & ~n364 ;
  assign n366 = ~n280 & ~n365 ;
  assign n367 = ~n279 & ~n366 ;
  assign n368 = ~n278 & ~n367 ;
  assign n369 = ~n277 & ~n368 ;
  assign n370 = ~n276 & ~n369 ;
  assign n371 = ~n275 & ~n370 ;
  assign n372 = ~n274 & ~n371 ;
  assign n373 = ~n273 & ~n372 ;
  assign n374 = ~n272 & ~n373 ;
  assign n375 = ~n271 & ~n374 ;
  assign n376 = ~n270 & ~n375 ;
  assign n377 = ~n269 & ~n376 ;
  assign n378 = ~n268 & ~n377 ;
  assign n379 = ~n267 & ~n378 ;
  assign n380 = ~n266 & ~n379 ;
  assign n381 = ~n265 & ~n380 ;
  assign n382 = ~n264 & ~n381 ;
  assign n383 = ~n263 & ~n382 ;
  assign n384 = ~n262 & ~n383 ;
  assign n385 = ~n261 & ~n384 ;
  assign n386 = x62 & ~n385 ;
  assign n387 = x30 & n385 ;
  assign n388 = ~n386 & ~n387 ;
  assign n389 = ~n260 & n388 ;
  assign n390 = x97 & ~n253 ;
  assign n391 = x65 & n253 ;
  assign n392 = ~n390 & ~n391 ;
  assign n393 = x33 & ~n385 ;
  assign n394 = x1 & n385 ;
  assign n395 = ~n393 & ~n394 ;
  assign n396 = ~n392 & n395 ;
  assign n397 = x96 & ~n253 ;
  assign n398 = x64 & n253 ;
  assign n399 = ~n397 & ~n398 ;
  assign n400 = x32 & ~n385 ;
  assign n401 = x0 & n385 ;
  assign n402 = ~n400 & ~n401 ;
  assign n403 = n399 & ~n402 ;
  assign n404 = ~n396 & n403 ;
  assign n405 = x98 & ~n253 ;
  assign n406 = x66 & n253 ;
  assign n407 = ~n405 & ~n406 ;
  assign n408 = x34 & ~n385 ;
  assign n409 = x2 & n385 ;
  assign n410 = ~n408 & ~n409 ;
  assign n411 = n407 & ~n410 ;
  assign n412 = n392 & ~n395 ;
  assign n413 = ~n411 & ~n412 ;
  assign n414 = ~n404 & n413 ;
  assign n415 = x99 & ~n253 ;
  assign n416 = x67 & n253 ;
  assign n417 = ~n415 & ~n416 ;
  assign n418 = x35 & ~n385 ;
  assign n419 = x3 & n385 ;
  assign n420 = ~n418 & ~n419 ;
  assign n421 = ~n417 & n420 ;
  assign n422 = ~n407 & n410 ;
  assign n423 = ~n421 & ~n422 ;
  assign n424 = ~n414 & n423 ;
  assign n425 = x100 & ~n253 ;
  assign n426 = x68 & n253 ;
  assign n427 = ~n425 & ~n426 ;
  assign n428 = x36 & ~n385 ;
  assign n429 = x4 & n385 ;
  assign n430 = ~n428 & ~n429 ;
  assign n431 = n427 & ~n430 ;
  assign n432 = n417 & ~n420 ;
  assign n433 = ~n431 & ~n432 ;
  assign n434 = ~n424 & n433 ;
  assign n435 = ~n427 & n430 ;
  assign n436 = x101 & ~n253 ;
  assign n437 = x69 & n253 ;
  assign n438 = ~n436 & ~n437 ;
  assign n439 = x37 & ~n385 ;
  assign n440 = x5 & n385 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = ~n438 & n441 ;
  assign n443 = ~n435 & ~n442 ;
  assign n444 = ~n434 & n443 ;
  assign n445 = x102 & ~n253 ;
  assign n446 = x70 & n253 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = x38 & ~n385 ;
  assign n449 = x6 & n385 ;
  assign n450 = ~n448 & ~n449 ;
  assign n451 = n447 & ~n450 ;
  assign n452 = n438 & ~n441 ;
  assign n453 = ~n451 & ~n452 ;
  assign n454 = ~n444 & n453 ;
  assign n455 = x39 & ~n385 ;
  assign n456 = x7 & n385 ;
  assign n457 = ~n455 & ~n456 ;
  assign n458 = x103 & ~n253 ;
  assign n459 = x71 & n253 ;
  assign n460 = ~n458 & ~n459 ;
  assign n461 = n457 & ~n460 ;
  assign n462 = ~n447 & n450 ;
  assign n463 = ~n461 & ~n462 ;
  assign n464 = ~n454 & n463 ;
  assign n465 = ~n457 & n460 ;
  assign n466 = x104 & ~n253 ;
  assign n467 = x72 & n253 ;
  assign n468 = ~n466 & ~n467 ;
  assign n469 = x40 & ~n385 ;
  assign n470 = x8 & n385 ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = n468 & ~n471 ;
  assign n473 = ~n465 & ~n472 ;
  assign n474 = ~n464 & n473 ;
  assign n475 = ~n468 & n471 ;
  assign n476 = x105 & ~n253 ;
  assign n477 = x73 & n253 ;
  assign n478 = ~n476 & ~n477 ;
  assign n479 = x41 & ~n385 ;
  assign n480 = x9 & n385 ;
  assign n481 = ~n479 & ~n480 ;
  assign n482 = ~n478 & n481 ;
  assign n483 = ~n475 & ~n482 ;
  assign n484 = ~n474 & n483 ;
  assign n485 = n478 & ~n481 ;
  assign n486 = x42 & ~n385 ;
  assign n487 = x10 & n385 ;
  assign n488 = ~n486 & ~n487 ;
  assign n489 = x106 & ~n253 ;
  assign n490 = x74 & n253 ;
  assign n491 = ~n489 & ~n490 ;
  assign n492 = ~n488 & n491 ;
  assign n493 = ~n485 & ~n492 ;
  assign n494 = ~n484 & n493 ;
  assign n495 = x43 & ~n385 ;
  assign n496 = x11 & n385 ;
  assign n497 = ~n495 & ~n496 ;
  assign n498 = x107 & ~n253 ;
  assign n499 = x75 & n253 ;
  assign n500 = ~n498 & ~n499 ;
  assign n501 = n497 & ~n500 ;
  assign n502 = n488 & ~n491 ;
  assign n503 = ~n501 & ~n502 ;
  assign n504 = ~n494 & n503 ;
  assign n505 = x108 & ~n253 ;
  assign n506 = x76 & n253 ;
  assign n507 = ~n505 & ~n506 ;
  assign n508 = x44 & ~n385 ;
  assign n509 = x12 & n385 ;
  assign n510 = ~n508 & ~n509 ;
  assign n511 = n507 & ~n510 ;
  assign n512 = ~n497 & n500 ;
  assign n513 = ~n511 & ~n512 ;
  assign n514 = ~n504 & n513 ;
  assign n515 = ~n507 & n510 ;
  assign n516 = x109 & ~n253 ;
  assign n517 = x77 & n253 ;
  assign n518 = ~n516 & ~n517 ;
  assign n519 = x45 & ~n385 ;
  assign n520 = x13 & n385 ;
  assign n521 = ~n519 & ~n520 ;
  assign n522 = ~n518 & n521 ;
  assign n523 = ~n515 & ~n522 ;
  assign n524 = ~n514 & n523 ;
  assign n525 = n518 & ~n521 ;
  assign n526 = x46 & ~n385 ;
  assign n527 = x14 & n385 ;
  assign n528 = ~n526 & ~n527 ;
  assign n529 = x110 & ~n253 ;
  assign n530 = x78 & n253 ;
  assign n531 = ~n529 & ~n530 ;
  assign n532 = ~n528 & n531 ;
  assign n533 = ~n525 & ~n532 ;
  assign n534 = ~n524 & n533 ;
  assign n535 = x47 & ~n385 ;
  assign n536 = x15 & n385 ;
  assign n537 = ~n535 & ~n536 ;
  assign n538 = x111 & ~n253 ;
  assign n539 = x79 & n253 ;
  assign n540 = ~n538 & ~n539 ;
  assign n541 = n537 & ~n540 ;
  assign n542 = n528 & ~n531 ;
  assign n543 = ~n541 & ~n542 ;
  assign n544 = ~n534 & n543 ;
  assign n545 = x112 & ~n253 ;
  assign n546 = x80 & n253 ;
  assign n547 = ~n545 & ~n546 ;
  assign n548 = x48 & ~n385 ;
  assign n549 = x16 & n385 ;
  assign n550 = ~n548 & ~n549 ;
  assign n551 = n547 & ~n550 ;
  assign n552 = ~n537 & n540 ;
  assign n553 = ~n551 & ~n552 ;
  assign n554 = ~n544 & n553 ;
  assign n555 = ~n547 & n550 ;
  assign n556 = x113 & ~n253 ;
  assign n557 = x81 & n253 ;
  assign n558 = ~n556 & ~n557 ;
  assign n559 = x49 & ~n385 ;
  assign n560 = x17 & n385 ;
  assign n561 = ~n559 & ~n560 ;
  assign n562 = ~n558 & n561 ;
  assign n563 = ~n555 & ~n562 ;
  assign n564 = ~n554 & n563 ;
  assign n565 = n558 & ~n561 ;
  assign n566 = x50 & ~n385 ;
  assign n567 = x18 & n385 ;
  assign n568 = ~n566 & ~n567 ;
  assign n569 = x114 & ~n253 ;
  assign n570 = x82 & n253 ;
  assign n571 = ~n569 & ~n570 ;
  assign n572 = ~n568 & n571 ;
  assign n573 = ~n565 & ~n572 ;
  assign n574 = ~n564 & n573 ;
  assign n575 = x51 & ~n385 ;
  assign n576 = x19 & n385 ;
  assign n577 = ~n575 & ~n576 ;
  assign n578 = x115 & ~n253 ;
  assign n579 = x83 & n253 ;
  assign n580 = ~n578 & ~n579 ;
  assign n581 = n577 & ~n580 ;
  assign n582 = n568 & ~n571 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = ~n574 & n583 ;
  assign n585 = x116 & ~n253 ;
  assign n586 = x84 & n253 ;
  assign n587 = ~n585 & ~n586 ;
  assign n588 = x52 & ~n385 ;
  assign n589 = x20 & n385 ;
  assign n590 = ~n588 & ~n589 ;
  assign n591 = n587 & ~n590 ;
  assign n592 = ~n577 & n580 ;
  assign n593 = ~n591 & ~n592 ;
  assign n594 = ~n584 & n593 ;
  assign n595 = ~n587 & n590 ;
  assign n596 = x117 & ~n253 ;
  assign n597 = x85 & n253 ;
  assign n598 = ~n596 & ~n597 ;
  assign n599 = x53 & ~n385 ;
  assign n600 = x21 & n385 ;
  assign n601 = ~n599 & ~n600 ;
  assign n602 = ~n598 & n601 ;
  assign n603 = ~n595 & ~n602 ;
  assign n604 = ~n594 & n603 ;
  assign n605 = n598 & ~n601 ;
  assign n606 = x54 & ~n385 ;
  assign n607 = x22 & n385 ;
  assign n608 = ~n606 & ~n607 ;
  assign n609 = x118 & ~n253 ;
  assign n610 = x86 & n253 ;
  assign n611 = ~n609 & ~n610 ;
  assign n612 = ~n608 & n611 ;
  assign n613 = ~n605 & ~n612 ;
  assign n614 = ~n604 & n613 ;
  assign n615 = x55 & ~n385 ;
  assign n616 = x23 & n385 ;
  assign n617 = ~n615 & ~n616 ;
  assign n618 = x119 & ~n253 ;
  assign n619 = x87 & n253 ;
  assign n620 = ~n618 & ~n619 ;
  assign n621 = n617 & ~n620 ;
  assign n622 = n608 & ~n611 ;
  assign n623 = ~n621 & ~n622 ;
  assign n624 = ~n614 & n623 ;
  assign n625 = x120 & ~n253 ;
  assign n626 = x88 & n253 ;
  assign n627 = ~n625 & ~n626 ;
  assign n628 = x56 & ~n385 ;
  assign n629 = x24 & n385 ;
  assign n630 = ~n628 & ~n629 ;
  assign n631 = n627 & ~n630 ;
  assign n632 = ~n617 & n620 ;
  assign n633 = ~n631 & ~n632 ;
  assign n634 = ~n624 & n633 ;
  assign n635 = ~n627 & n630 ;
  assign n636 = x121 & ~n253 ;
  assign n637 = x89 & n253 ;
  assign n638 = ~n636 & ~n637 ;
  assign n639 = x57 & ~n385 ;
  assign n640 = x25 & n385 ;
  assign n641 = ~n639 & ~n640 ;
  assign n642 = ~n638 & n641 ;
  assign n643 = ~n635 & ~n642 ;
  assign n644 = ~n634 & n643 ;
  assign n645 = n638 & ~n641 ;
  assign n646 = x58 & ~n385 ;
  assign n647 = x26 & n385 ;
  assign n648 = ~n646 & ~n647 ;
  assign n649 = x122 & ~n253 ;
  assign n650 = x90 & n253 ;
  assign n651 = ~n649 & ~n650 ;
  assign n652 = ~n648 & n651 ;
  assign n653 = ~n645 & ~n652 ;
  assign n654 = ~n644 & n653 ;
  assign n655 = x59 & ~n385 ;
  assign n656 = x27 & n385 ;
  assign n657 = ~n655 & ~n656 ;
  assign n658 = x123 & ~n253 ;
  assign n659 = x91 & n253 ;
  assign n660 = ~n658 & ~n659 ;
  assign n661 = n657 & ~n660 ;
  assign n662 = n648 & ~n651 ;
  assign n663 = ~n661 & ~n662 ;
  assign n664 = ~n654 & n663 ;
  assign n665 = x124 & ~n253 ;
  assign n666 = x92 & n253 ;
  assign n667 = ~n665 & ~n666 ;
  assign n668 = x60 & ~n385 ;
  assign n669 = x28 & n385 ;
  assign n670 = ~n668 & ~n669 ;
  assign n671 = n667 & ~n670 ;
  assign n672 = ~n657 & n660 ;
  assign n673 = ~n671 & ~n672 ;
  assign n674 = ~n664 & n673 ;
  assign n675 = ~n667 & n670 ;
  assign n676 = x125 & ~n253 ;
  assign n677 = x93 & n253 ;
  assign n678 = ~n676 & ~n677 ;
  assign n679 = x61 & ~n385 ;
  assign n680 = x29 & n385 ;
  assign n681 = ~n679 & ~n680 ;
  assign n682 = ~n678 & n681 ;
  assign n683 = ~n675 & ~n682 ;
  assign n684 = ~n674 & n683 ;
  assign n685 = n260 & ~n388 ;
  assign n686 = n678 & ~n681 ;
  assign n687 = ~n685 & ~n686 ;
  assign n688 = ~n684 & n687 ;
  assign n689 = ~n389 & ~n688 ;
  assign n690 = ~n257 & ~n689 ;
  assign n691 = ~n256 & ~n690 ;
  assign n692 = ~n253 & ~n691 ;
  assign n693 = ~n385 & n691 ;
  assign n694 = ~n692 & ~n693 ;
  assign n695 = ~n402 & n691 ;
  assign n696 = ~n399 & ~n691 ;
  assign n697 = ~n695 & ~n696 ;
  assign n698 = ~n395 & n691 ;
  assign n699 = ~n392 & ~n691 ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = ~n410 & n691 ;
  assign n702 = ~n407 & ~n691 ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = ~n420 & n691 ;
  assign n705 = ~n417 & ~n691 ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = ~n430 & n691 ;
  assign n708 = ~n427 & ~n691 ;
  assign n709 = ~n707 & ~n708 ;
  assign n710 = ~n441 & n691 ;
  assign n711 = ~n438 & ~n691 ;
  assign n712 = ~n710 & ~n711 ;
  assign n713 = ~n450 & n691 ;
  assign n714 = ~n447 & ~n691 ;
  assign n715 = ~n713 & ~n714 ;
  assign n716 = ~n457 & n691 ;
  assign n717 = ~n460 & ~n691 ;
  assign n718 = ~n716 & ~n717 ;
  assign n719 = ~n471 & n691 ;
  assign n720 = ~n468 & ~n691 ;
  assign n721 = ~n719 & ~n720 ;
  assign n722 = ~n481 & n691 ;
  assign n723 = ~n478 & ~n691 ;
  assign n724 = ~n722 & ~n723 ;
  assign n725 = ~n488 & n691 ;
  assign n726 = ~n491 & ~n691 ;
  assign n727 = ~n725 & ~n726 ;
  assign n728 = ~n497 & n691 ;
  assign n729 = ~n500 & ~n691 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = ~n510 & n691 ;
  assign n732 = ~n507 & ~n691 ;
  assign n733 = ~n731 & ~n732 ;
  assign n734 = ~n521 & n691 ;
  assign n735 = ~n518 & ~n691 ;
  assign n736 = ~n734 & ~n735 ;
  assign n737 = ~n528 & n691 ;
  assign n738 = ~n531 & ~n691 ;
  assign n739 = ~n737 & ~n738 ;
  assign n740 = ~n537 & n691 ;
  assign n741 = ~n540 & ~n691 ;
  assign n742 = ~n740 & ~n741 ;
  assign n743 = ~n550 & n691 ;
  assign n744 = ~n547 & ~n691 ;
  assign n745 = ~n743 & ~n744 ;
  assign n746 = ~n561 & n691 ;
  assign n747 = ~n558 & ~n691 ;
  assign n748 = ~n746 & ~n747 ;
  assign n749 = ~n568 & n691 ;
  assign n750 = ~n571 & ~n691 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = ~n577 & n691 ;
  assign n753 = ~n580 & ~n691 ;
  assign n754 = ~n752 & ~n753 ;
  assign n755 = ~n590 & n691 ;
  assign n756 = ~n587 & ~n691 ;
  assign n757 = ~n755 & ~n756 ;
  assign n758 = ~n601 & n691 ;
  assign n759 = ~n598 & ~n691 ;
  assign n760 = ~n758 & ~n759 ;
  assign n761 = ~n608 & n691 ;
  assign n762 = ~n611 & ~n691 ;
  assign n763 = ~n761 & ~n762 ;
  assign n764 = ~n617 & n691 ;
  assign n765 = ~n620 & ~n691 ;
  assign n766 = ~n764 & ~n765 ;
  assign n767 = ~n630 & n691 ;
  assign n768 = ~n627 & ~n691 ;
  assign n769 = ~n767 & ~n768 ;
  assign n770 = ~n641 & n691 ;
  assign n771 = ~n638 & ~n691 ;
  assign n772 = ~n770 & ~n771 ;
  assign n773 = ~n648 & n691 ;
  assign n774 = ~n651 & ~n691 ;
  assign n775 = ~n773 & ~n774 ;
  assign n776 = ~n657 & n691 ;
  assign n777 = ~n660 & ~n691 ;
  assign n778 = ~n776 & ~n777 ;
  assign n779 = ~n670 & n691 ;
  assign n780 = ~n667 & ~n691 ;
  assign n781 = ~n779 & ~n780 ;
  assign n782 = ~n681 & n691 ;
  assign n783 = ~n678 & ~n691 ;
  assign n784 = ~n782 & ~n783 ;
  assign n785 = ~n388 & n691 ;
  assign n786 = ~n260 & ~n691 ;
  assign n787 = ~n785 & ~n786 ;
  assign n788 = n254 & n255 ;
  assign y0 = ~n694 ;
  assign y1 = ~n691 ;
  assign y2 = ~n697 ;
  assign y3 = ~n700 ;
  assign y4 = ~n703 ;
  assign y5 = ~n706 ;
  assign y6 = ~n709 ;
  assign y7 = ~n712 ;
  assign y8 = ~n715 ;
  assign y9 = ~n718 ;
  assign y10 = ~n721 ;
  assign y11 = ~n724 ;
  assign y12 = ~n727 ;
  assign y13 = ~n730 ;
  assign y14 = ~n733 ;
  assign y15 = ~n736 ;
  assign y16 = ~n739 ;
  assign y17 = ~n742 ;
  assign y18 = ~n745 ;
  assign y19 = ~n748 ;
  assign y20 = ~n751 ;
  assign y21 = ~n754 ;
  assign y22 = ~n757 ;
  assign y23 = ~n760 ;
  assign y24 = ~n763 ;
  assign y25 = ~n766 ;
  assign y26 = ~n769 ;
  assign y27 = ~n772 ;
  assign y28 = ~n775 ;
  assign y29 = ~n778 ;
  assign y30 = ~n781 ;
  assign y31 = ~n784 ;
  assign y32 = ~n787 ;
  assign y33 = ~n788 ;
endmodule
