module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 ;
  assign n11 = x1 & ~x8 ;
  assign n12 = ~x1 & x9 ;
  assign n13 = x2 & ~x3 ;
  assign n14 = n12 & n13 ;
  assign n15 = ~n11 & ~n14 ;
  assign n16 = ~x0 & ~n15 ;
  assign n17 = x2 & x6 ;
  assign n18 = n17 ^ x6 ;
  assign n19 = x3 & n18 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = x2 & x9 ;
  assign n22 = ~x1 & ~x9 ;
  assign n23 = ~n21 & n22 ;
  assign n24 = ~n20 & n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = x8 & ~n25 ;
  assign n27 = n26 ^ x8 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n16 & n28 ;
  assign n30 = n29 ^ n16 ;
  assign n31 = n30 ^ n28 ;
  assign n44 = ~x2 & x5 ;
  assign n45 = x0 & ~x9 ;
  assign n49 = x6 & ~n45 ;
  assign n50 = n44 & n49 ;
  assign n48 = x5 & x6 ;
  assign n51 = n50 ^ n48 ;
  assign n41 = ~x0 & x9 ;
  assign n42 = x1 & ~x3 ;
  assign n43 = ~n41 & n42 ;
  assign n46 = n44 & ~n45 ;
  assign n47 = n43 & n46 ;
  assign n52 = n51 ^ n47 ;
  assign n53 = ~x0 & ~x3 ;
  assign n54 = x6 & n53 ;
  assign n57 = x1 & ~x9 ;
  assign n58 = ~x2 & n57 ;
  assign n59 = n54 & n58 ;
  assign n60 = ~n52 & n59 ;
  assign n61 = n60 ^ n52 ;
  assign n55 = n21 & n54 ;
  assign n56 = ~n52 & n55 ;
  assign n62 = n61 ^ n56 ;
  assign n32 = ~x8 & n22 ;
  assign n33 = x2 & x3 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n34 ^ x3 ;
  assign n36 = ~x0 & ~n35 ;
  assign n37 = n32 & n36 ;
  assign n65 = ~x5 & x8 ;
  assign n66 = ~n37 & n65 ;
  assign n67 = n62 & n66 ;
  assign n68 = n31 & n67 ;
  assign n63 = x8 & ~n37 ;
  assign n64 = n62 & n63 ;
  assign n69 = n68 ^ n64 ;
  assign n38 = ~x5 & ~n37 ;
  assign n39 = n31 & n38 ;
  assign n40 = n39 ^ n37 ;
  assign n70 = n69 ^ n40 ;
  assign n71 = ~x0 & ~x2 ;
  assign n72 = n12 & n71 ;
  assign n73 = ~x5 & x6 ;
  assign n74 = ~n72 & n73 ;
  assign n75 = n74 ^ x6 ;
  assign n82 = x8 & n75 ;
  assign n76 = x1 & x5 ;
  assign n77 = x2 & n76 ;
  assign n78 = x9 ^ x0 ;
  assign n79 = x8 & ~n78 ;
  assign n80 = n77 & n79 ;
  assign n81 = ~n75 & n80 ;
  assign n83 = n82 ^ n81 ;
  assign n92 = x3 & x5 ;
  assign n93 = ~n83 & n92 ;
  assign n94 = n93 ^ x3 ;
  assign n84 = ~x1 & ~n41 ;
  assign n85 = ~x8 & ~n84 ;
  assign n86 = ~x1 & x2 ;
  assign n87 = n45 & n86 ;
  assign n88 = x3 & ~x5 ;
  assign n89 = ~n87 & n88 ;
  assign n90 = ~n85 & n89 ;
  assign n91 = ~n83 & n90 ;
  assign n95 = n94 ^ n91 ;
  assign n98 = x7 & ~n95 ;
  assign n99 = ~n70 & n98 ;
  assign n100 = n99 ^ x7 ;
  assign n96 = ~n70 & n95 ;
  assign n97 = n96 ^ n70 ;
  assign n101 = n100 ^ n97 ;
  assign n143 = x3 & x9 ;
  assign n142 = x1 & x9 ;
  assign n144 = n143 ^ n142 ;
  assign n140 = ~x3 & x9 ;
  assign n141 = n86 & n140 ;
  assign n145 = n144 ^ n141 ;
  assign n128 = x2 ^ x0 ;
  assign n129 = n128 ^ x2 ;
  assign n127 = x9 ^ x2 ;
  assign n130 = n129 ^ n127 ;
  assign n131 = n127 ^ x2 ;
  assign n132 = n130 & ~n131 ;
  assign n133 = n132 ^ n127 ;
  assign n134 = x9 ^ x3 ;
  assign n135 = ~x1 & n134 ;
  assign n136 = ~n133 & n135 ;
  assign n137 = n136 ^ x1 ;
  assign n138 = n137 ^ n134 ;
  assign n139 = n138 ^ x9 ;
  assign n146 = n145 ^ n139 ;
  assign n123 = x0 & ~x1 ;
  assign n124 = x2 & n123 ;
  assign n125 = n124 ^ x2 ;
  assign n122 = x5 & n71 ;
  assign n126 = n125 ^ n122 ;
  assign n147 = n146 ^ n126 ;
  assign n148 = n126 ^ x9 ;
  assign n149 = n147 & ~n148 ;
  assign n150 = n149 ^ n145 ;
  assign n151 = n150 ^ n126 ;
  assign n152 = x7 & ~n151 ;
  assign n153 = n152 ^ x7 ;
  assign n154 = n153 ^ n151 ;
  assign n157 = ~x3 & ~x5 ;
  assign n158 = ~n12 & n157 ;
  assign n164 = ~x7 & ~x9 ;
  assign n165 = n123 & n164 ;
  assign n166 = ~n158 & n165 ;
  assign n160 = ~x0 & x1 ;
  assign n161 = x7 & x9 ;
  assign n162 = n160 & n161 ;
  assign n163 = n158 & n162 ;
  assign n167 = n166 ^ n163 ;
  assign n159 = ~x1 & n158 ;
  assign n168 = n167 ^ n159 ;
  assign n106 = x1 & ~x7 ;
  assign n107 = x9 & n106 ;
  assign n169 = n168 ^ n107 ;
  assign n170 = ~x2 & x6 ;
  assign n171 = ~x8 & n170 ;
  assign n172 = n169 & n171 ;
  assign n173 = ~n154 & n172 ;
  assign n155 = x6 & ~x8 ;
  assign n156 = n154 & n155 ;
  assign n174 = n173 ^ n156 ;
  assign n175 = n174 ^ x6 ;
  assign n102 = x0 & ~x2 ;
  assign n103 = x7 & x8 ;
  assign n104 = x1 & ~x5 ;
  assign n105 = n103 & n104 ;
  assign n108 = n107 ^ n105 ;
  assign n109 = ~x5 & ~x9 ;
  assign n110 = ~n106 & n109 ;
  assign n111 = ~n108 & ~n110 ;
  assign n112 = n102 & ~n111 ;
  assign n113 = ~x5 & x7 ;
  assign n114 = x8 & n113 ;
  assign n115 = ~x0 & ~x1 ;
  assign n116 = x2 & ~x9 ;
  assign n117 = n115 & n116 ;
  assign n118 = n114 & n117 ;
  assign n119 = ~x3 & ~n118 ;
  assign n120 = ~n112 & n119 ;
  assign n121 = n120 ^ x3 ;
  assign n176 = n175 ^ n121 ;
  assign n184 = x8 & ~n154 ;
  assign n181 = ~x2 & x8 ;
  assign n182 = n169 & n181 ;
  assign n183 = ~n154 & n182 ;
  assign n185 = n184 ^ n183 ;
  assign n186 = n185 ^ x8 ;
  assign n177 = ~x2 & n169 ;
  assign n178 = n154 & n177 ;
  assign n179 = n178 ^ n177 ;
  assign n180 = n179 ^ n154 ;
  assign n187 = n186 ^ n180 ;
  assign n188 = n187 ^ n121 ;
  assign n189 = n176 & ~n188 ;
  assign n190 = n189 ^ n174 ;
  assign n191 = n190 ^ n121 ;
  assign n195 = ~x6 & x8 ;
  assign n196 = x5 & ~n195 ;
  assign n197 = ~x6 & ~x9 ;
  assign n198 = x4 & x8 ;
  assign n199 = ~n197 & ~n198 ;
  assign n200 = n196 & ~n199 ;
  assign n201 = x6 & ~x9 ;
  assign n202 = x4 & x9 ;
  assign n203 = ~n201 & ~n202 ;
  assign n204 = ~x8 & ~n48 ;
  assign n205 = ~n203 & n204 ;
  assign n206 = ~n200 & ~n205 ;
  assign n207 = ~x1 & ~x3 ;
  assign n208 = ~x7 & n71 ;
  assign n209 = n207 & n208 ;
  assign n210 = ~n206 & n209 ;
  assign n211 = ~x4 & n210 ;
  assign n212 = n191 & n211 ;
  assign n213 = ~n101 & n212 ;
  assign n214 = n213 ^ n211 ;
  assign n192 = ~x4 & n191 ;
  assign n193 = ~n101 & n192 ;
  assign n194 = n193 ^ x4 ;
  assign n215 = n214 ^ n194 ;
  assign n216 = n215 ^ n210 ;
  assign n224 = x0 & x1 ;
  assign n221 = x5 ^ x0 ;
  assign n225 = ~n181 & ~n221 ;
  assign n226 = n224 & n225 ;
  assign n217 = x3 & x8 ;
  assign n218 = ~x2 & ~n217 ;
  assign n222 = n160 & ~n221 ;
  assign n223 = n218 & n222 ;
  assign n227 = n226 ^ n223 ;
  assign n219 = n115 & ~n218 ;
  assign n220 = n219 ^ x1 ;
  assign n228 = n227 ^ n220 ;
  assign n229 = ~x2 & ~x8 ;
  assign n230 = x5 & n229 ;
  assign n237 = ~x1 & n230 ;
  assign n238 = ~n228 & n237 ;
  assign n239 = n238 ^ n228 ;
  assign n232 = x3 & ~x8 ;
  assign n231 = x5 & x8 ;
  assign n233 = n232 ^ n231 ;
  assign n234 = n123 & n233 ;
  assign n235 = ~n230 & n234 ;
  assign n236 = ~n228 & n235 ;
  assign n240 = n239 ^ n236 ;
  assign n241 = ~x6 & n240 ;
  assign n242 = ~x0 & x8 ;
  assign n243 = ~x2 & ~n242 ;
  assign n244 = ~x1 & ~x6 ;
  assign n245 = ~n224 & ~n244 ;
  assign n246 = n243 & n245 ;
  assign n256 = n109 & n246 ;
  assign n257 = n256 ^ x9 ;
  assign n249 = x6 & x8 ;
  assign n250 = n86 & n249 ;
  assign n247 = ~x1 & ~x2 ;
  assign n248 = ~x8 & n247 ;
  assign n251 = n250 ^ n248 ;
  assign n252 = n251 ^ x2 ;
  assign n253 = ~x9 & n88 ;
  assign n254 = ~n252 & n253 ;
  assign n255 = ~n246 & n254 ;
  assign n258 = n257 ^ n255 ;
  assign n259 = ~n241 & ~n258 ;
  assign n260 = ~x1 & x3 ;
  assign n261 = n229 & n260 ;
  assign n262 = n261 ^ n76 ;
  assign n263 = x0 & n262 ;
  assign n266 = ~x2 & ~x3 ;
  assign n267 = x5 & n266 ;
  assign n264 = x1 & x2 ;
  assign n265 = n88 & n264 ;
  assign n268 = n267 ^ n265 ;
  assign n269 = n268 ^ x5 ;
  assign n270 = x6 & ~n269 ;
  assign n271 = ~n263 & n270 ;
  assign n272 = n271 ^ x6 ;
  assign n273 = x5 & ~x8 ;
  assign n274 = x3 & n264 ;
  assign n275 = n273 & n274 ;
  assign n276 = ~x4 & x9 ;
  assign n277 = ~n275 & n276 ;
  assign n278 = ~n272 & n277 ;
  assign n279 = n278 ^ x4 ;
  assign n280 = ~n259 & ~n279 ;
  assign n300 = ~x0 & ~x5 ;
  assign n301 = ~x6 & n300 ;
  assign n302 = x8 & x9 ;
  assign n322 = n301 & n302 ;
  assign n310 = ~x6 & x9 ;
  assign n284 = ~x8 & x9 ;
  assign n287 = x0 & x6 ;
  assign n288 = n284 & n287 ;
  assign n311 = n310 ^ n288 ;
  assign n323 = n322 ^ n311 ;
  assign n282 = x0 & ~x5 ;
  assign n306 = x8 & ~x9 ;
  assign n307 = n282 & n306 ;
  assign n305 = x5 & ~x9 ;
  assign n308 = n307 ^ n305 ;
  assign n324 = n323 ^ n308 ;
  assign n317 = x0 & x8 ;
  assign n318 = n21 & n317 ;
  assign n315 = ~x0 & ~x9 ;
  assign n316 = n229 & n315 ;
  assign n319 = n318 ^ n316 ;
  assign n325 = x5 & n86 ;
  assign n326 = n319 & n325 ;
  assign n327 = ~n324 & n326 ;
  assign n320 = ~x1 & x5 ;
  assign n321 = n319 & n320 ;
  assign n328 = n327 ^ n321 ;
  assign n312 = n86 & ~n311 ;
  assign n309 = n86 & n308 ;
  assign n313 = n312 ^ n309 ;
  assign n303 = n86 & n302 ;
  assign n304 = n301 & n303 ;
  assign n314 = n313 ^ n304 ;
  assign n329 = n328 ^ n314 ;
  assign n330 = n116 & n195 ;
  assign n335 = ~n329 & ~n330 ;
  assign n336 = ~x4 & ~n335 ;
  assign n285 = ~x0 & x5 ;
  assign n286 = n284 & n285 ;
  assign n289 = n288 ^ n286 ;
  assign n283 = n195 & n282 ;
  assign n290 = n289 ^ n283 ;
  assign n291 = ~x2 & n290 ;
  assign n294 = ~x0 & x6 ;
  assign n295 = ~x2 & ~n294 ;
  assign n296 = ~x9 & n65 ;
  assign n297 = ~n295 & n296 ;
  assign n292 = ~x6 & ~x8 ;
  assign n293 = ~x9 & n292 ;
  assign n298 = n297 ^ n293 ;
  assign n299 = ~n291 & ~n298 ;
  assign n331 = x1 & ~x4 ;
  assign n332 = ~n330 & n331 ;
  assign n333 = ~n329 & n332 ;
  assign n334 = ~n299 & n333 ;
  assign n337 = n336 ^ n334 ;
  assign n338 = ~x2 & n115 ;
  assign n339 = ~n198 & ~n273 ;
  assign n340 = n197 & ~n339 ;
  assign n341 = x6 & x9 ;
  assign n342 = x4 & n341 ;
  assign n343 = ~n340 & ~n342 ;
  assign n344 = n338 & ~n343 ;
  assign n365 = ~x6 & n157 ;
  assign n366 = ~x4 & n365 ;
  assign n369 = ~x7 & n117 ;
  assign n370 = n366 & n369 ;
  assign n372 = ~x3 & n370 ;
  assign n373 = ~n344 & n372 ;
  assign n374 = ~n337 & n373 ;
  assign n371 = x3 & n370 ;
  assign n375 = n374 ^ n371 ;
  assign n376 = ~n280 & n375 ;
  assign n351 = ~x2 & x9 ;
  assign n352 = n123 & n351 ;
  assign n353 = n352 ^ n71 ;
  assign n356 = x2 & ~x8 ;
  assign n357 = ~n115 & n356 ;
  assign n358 = ~n353 & n357 ;
  assign n355 = n57 & n181 ;
  assign n359 = n358 ^ n355 ;
  assign n354 = ~x8 & ~n353 ;
  assign n360 = n359 ^ n354 ;
  assign n363 = ~n117 & ~n360 ;
  assign n361 = ~x7 & ~n117 ;
  assign n362 = n360 & n361 ;
  assign n364 = n363 ^ n362 ;
  assign n367 = x7 & n366 ;
  assign n368 = ~n364 & n367 ;
  assign n377 = n376 ^ n368 ;
  assign n345 = ~x3 & ~x7 ;
  assign n346 = ~n344 & n345 ;
  assign n347 = ~n337 & n346 ;
  assign n281 = x3 & ~x7 ;
  assign n348 = n347 ^ n281 ;
  assign n349 = ~n280 & n348 ;
  assign n350 = n349 ^ x7 ;
  assign n378 = n377 ^ n350 ;
  assign n400 = ~x1 & ~x8 ;
  assign n482 = n45 & n400 ;
  assign n477 = x1 & ~n41 ;
  assign n478 = x0 & x7 ;
  assign n479 = n302 & n478 ;
  assign n480 = n479 ^ x0 ;
  assign n481 = n477 & ~n480 ;
  assign n483 = n482 ^ n481 ;
  assign n484 = ~x5 & ~x6 ;
  assign n485 = ~x4 & ~n35 ;
  assign n486 = n484 & n485 ;
  assign n487 = n483 & n486 ;
  assign n441 = ~x9 & n231 ;
  assign n439 = x5 & x9 ;
  assign n440 = ~n317 & n439 ;
  assign n442 = n441 ^ n440 ;
  assign n443 = ~n21 & n104 ;
  assign n444 = n443 ^ x1 ;
  assign n445 = ~n442 & n444 ;
  assign n450 = ~x3 & n445 ;
  assign n446 = x9 ^ x8 ;
  assign n447 = ~n22 & ~n446 ;
  assign n448 = n13 & ~n447 ;
  assign n449 = ~n445 & n448 ;
  assign n451 = n450 ^ n449 ;
  assign n452 = x5 & ~n260 ;
  assign n453 = ~x8 & ~x9 ;
  assign n463 = n102 & n453 ;
  assign n464 = ~n452 & n463 ;
  assign n465 = ~n451 & n464 ;
  assign n466 = n465 ^ n451 ;
  assign n454 = ~x2 & n453 ;
  assign n455 = ~n452 & n454 ;
  assign n456 = x9 & ~n35 ;
  assign n457 = n456 ^ x9 ;
  assign n458 = ~x1 & x8 ;
  assign n459 = x0 & n458 ;
  assign n460 = n457 & n459 ;
  assign n461 = ~n455 & n460 ;
  assign n462 = ~n451 & n461 ;
  assign n467 = n466 ^ n462 ;
  assign n419 = n264 & n341 ;
  assign n417 = ~x1 & x6 ;
  assign n418 = x8 & n417 ;
  assign n420 = n419 ^ n418 ;
  assign n423 = n232 & ~n420 ;
  assign n424 = n423 ^ x3 ;
  assign n421 = ~x9 & n33 ;
  assign n422 = ~n420 & n421 ;
  assign n425 = n424 ^ n422 ;
  assign n430 = x9 ^ x1 ;
  assign n431 = ~x8 & ~n430 ;
  assign n432 = n266 & n431 ;
  assign n426 = x1 & ~x6 ;
  assign n427 = n426 ^ n12 ;
  assign n428 = n427 ^ n197 ;
  assign n429 = n181 & ~n428 ;
  assign n433 = n432 ^ n429 ;
  assign n468 = ~x4 & ~x6 ;
  assign n470 = n282 & n468 ;
  assign n471 = ~n433 & n470 ;
  assign n472 = ~n425 & n471 ;
  assign n469 = ~n282 & n468 ;
  assign n473 = n472 ^ n469 ;
  assign n498 = n467 & n473 ;
  assign n434 = n282 & ~n433 ;
  assign n435 = ~n425 & n434 ;
  assign n436 = n435 ^ n282 ;
  assign n437 = ~x4 & n436 ;
  assign n499 = n498 ^ n437 ;
  assign n500 = ~x7 & n499 ;
  assign n501 = ~n487 & n500 ;
  assign n502 = n501 ^ n487 ;
  assign n379 = x2 & ~n195 ;
  assign n380 = x1 & ~n379 ;
  assign n381 = x5 & ~n218 ;
  assign n382 = ~n380 & n381 ;
  assign n383 = ~n57 & ~n232 ;
  assign n384 = x3 & ~x9 ;
  assign n385 = ~x6 & ~n384 ;
  assign n386 = ~n383 & n385 ;
  assign n387 = x1 & n140 ;
  assign n388 = ~x4 & n155 ;
  assign n389 = n387 & n388 ;
  assign n390 = n389 ^ x4 ;
  assign n391 = ~n386 & ~n390 ;
  assign n392 = ~n382 & n391 ;
  assign n399 = ~x3 & n73 ;
  assign n401 = ~x9 & n400 ;
  assign n402 = n399 & n401 ;
  assign n395 = ~x5 & ~x8 ;
  assign n393 = ~x2 & x3 ;
  assign n394 = x8 & n393 ;
  assign n396 = n395 ^ n394 ;
  assign n397 = n396 ^ n92 ;
  assign n398 = n57 & ~n397 ;
  assign n403 = n402 ^ n398 ;
  assign n405 = x1 & x8 ;
  assign n407 = ~x9 & n405 ;
  assign n406 = n197 & ~n405 ;
  assign n408 = n407 ^ n406 ;
  assign n410 = n12 & n229 ;
  assign n411 = ~n408 & n410 ;
  assign n409 = ~x2 & ~n408 ;
  assign n412 = n411 ^ n409 ;
  assign n404 = ~x8 & n12 ;
  assign n413 = n412 ^ n404 ;
  assign n414 = x3 & n413 ;
  assign n415 = ~n403 & ~n414 ;
  assign n416 = n392 & n415 ;
  assign n474 = ~x7 & n473 ;
  assign n475 = n467 & n474 ;
  assign n438 = ~x7 & ~n437 ;
  assign n476 = n475 ^ n438 ;
  assign n488 = n306 ^ n292 ;
  assign n489 = ~x5 & ~n488 ;
  assign n490 = ~x2 & x4 ;
  assign n491 = n207 & n490 ;
  assign n492 = ~n489 & n491 ;
  assign n493 = n492 ^ x4 ;
  assign n494 = ~x0 & ~n493 ;
  assign n495 = ~n487 & n494 ;
  assign n496 = n476 & n495 ;
  assign n497 = ~n416 & n496 ;
  assign n503 = n502 ^ n497 ;
  assign n569 = x0 & ~x4 ;
  assign n581 = n44 & n306 ;
  assign n576 = ~x6 & ~n232 ;
  assign n574 = ~x3 & x5 ;
  assign n575 = n284 & n574 ;
  assign n584 = n575 ^ x3 ;
  assign n604 = n576 & ~n584 ;
  assign n605 = n581 & n604 ;
  assign n585 = x2 & n88 ;
  assign n601 = n306 & n393 ;
  assign n600 = n88 & n306 ;
  assign n602 = n601 ^ n600 ;
  assign n603 = n585 & n602 ;
  assign n606 = n605 ^ n603 ;
  assign n597 = x2 & ~n88 ;
  assign n580 = n116 & ~n233 ;
  assign n582 = n581 ^ n580 ;
  assign n598 = n576 & n582 ;
  assign n599 = n597 & n598 ;
  assign n607 = n606 ^ n599 ;
  assign n593 = x2 & ~x6 ;
  assign n594 = ~n232 & n593 ;
  assign n595 = n584 & n594 ;
  assign n591 = ~x2 & n88 ;
  assign n592 = ~n584 & n591 ;
  assign n596 = n595 ^ n592 ;
  assign n608 = n607 ^ n596 ;
  assign n588 = ~n576 & n585 ;
  assign n583 = n576 & ~n582 ;
  assign n586 = ~n584 & n585 ;
  assign n587 = n583 & n586 ;
  assign n589 = n588 ^ n587 ;
  assign n578 = ~x3 & n576 ;
  assign n577 = n575 & n576 ;
  assign n579 = n578 ^ n577 ;
  assign n590 = n589 ^ n579 ;
  assign n609 = n608 ^ n590 ;
  assign n620 = n142 & ~n609 ;
  assign n621 = n620 ^ x9 ;
  assign n610 = n230 & n244 ;
  assign n614 = ~x3 & ~x9 ;
  assign n615 = n73 & n614 ;
  assign n616 = n615 ^ x9 ;
  assign n617 = ~n610 & ~n616 ;
  assign n618 = n609 & n617 ;
  assign n611 = n22 & ~n399 ;
  assign n612 = ~n610 & n611 ;
  assign n613 = ~n609 & n612 ;
  assign n619 = n618 ^ n613 ;
  assign n622 = n621 ^ n619 ;
  assign n623 = n569 & ~n622 ;
  assign n537 = ~n109 & ~n292 ;
  assign n538 = ~x2 & ~n537 ;
  assign n541 = n104 & n310 ;
  assign n539 = x5 & ~x6 ;
  assign n540 = n306 & n539 ;
  assign n542 = n541 ^ n540 ;
  assign n543 = x3 & ~n542 ;
  assign n544 = ~n538 & n543 ;
  assign n545 = n544 ^ x3 ;
  assign n553 = x3 & ~x6 ;
  assign n558 = ~n73 & ~n553 ;
  assign n559 = n453 & n558 ;
  assign n560 = n559 ^ n306 ;
  assign n550 = ~x6 & n33 ;
  assign n549 = n73 & n266 ;
  assign n551 = n550 ^ n549 ;
  assign n552 = n551 ^ n73 ;
  assign n556 = x9 & ~n552 ;
  assign n554 = n284 & n553 ;
  assign n555 = ~n552 & n554 ;
  assign n557 = n556 ^ n555 ;
  assign n561 = n560 ^ n557 ;
  assign n562 = ~x1 & ~n561 ;
  assign n563 = ~n545 & n562 ;
  assign n564 = n563 ^ n545 ;
  assign n546 = ~x9 & n73 ;
  assign n547 = n405 & n546 ;
  assign n548 = ~n545 & n547 ;
  assign n565 = n564 ^ n548 ;
  assign n624 = ~x7 & ~n565 ;
  assign n625 = n623 & n624 ;
  assign n518 = x6 & n35 ;
  assign n519 = ~n384 & ~n518 ;
  assign n520 = x2 & n73 ;
  assign n521 = ~x1 & ~x4 ;
  assign n522 = ~n520 & n521 ;
  assign n523 = n519 & n522 ;
  assign n511 = n195 & n439 ;
  assign n510 = ~x8 & n109 ;
  assign n512 = n511 ^ n510 ;
  assign n513 = n331 & ~n512 ;
  assign n505 = n92 & n195 ;
  assign n506 = n505 ^ n88 ;
  assign n504 = n155 & n157 ;
  assign n507 = n506 ^ n504 ;
  assign n514 = x2 & ~n73 ;
  assign n515 = ~n507 & n514 ;
  assign n516 = n513 & n515 ;
  assign n508 = ~x2 & n331 ;
  assign n509 = ~n507 & n508 ;
  assign n517 = n516 ^ n509 ;
  assign n524 = n523 ^ n517 ;
  assign n526 = ~x3 & x4 ;
  assign n527 = n247 & n526 ;
  assign n528 = x6 ^ x5 ;
  assign n532 = n527 & ~n528 ;
  assign n529 = ~x5 & ~n528 ;
  assign n530 = ~n302 & n529 ;
  assign n531 = n527 & n530 ;
  assign n533 = n532 ^ n531 ;
  assign n566 = ~x0 & ~x4 ;
  assign n567 = ~n533 & n566 ;
  assign n568 = n524 & n567 ;
  assign n570 = n569 ^ n568 ;
  assign n571 = n565 & n570 ;
  assign n525 = n524 ^ x4 ;
  assign n534 = ~x0 & ~n533 ;
  assign n535 = n525 & n534 ;
  assign n536 = n535 ^ x0 ;
  assign n572 = n571 ^ n536 ;
  assign n573 = ~x7 & ~n572 ;
  assign n626 = n625 ^ n573 ;
  assign n627 = x2 & ~n115 ;
  assign n628 = ~x4 & n627 ;
  assign n629 = x4 ^ x3 ;
  assign n630 = n338 & n629 ;
  assign n631 = ~n628 & ~n630 ;
  assign n632 = ~x7 & n48 ;
  assign n633 = ~n631 & n632 ;
  assign n634 = x3 & ~x4 ;
  assign n635 = ~n338 & n634 ;
  assign n636 = n338 & n526 ;
  assign n637 = ~n635 & ~n636 ;
  assign n638 = n632 & ~n637 ;
  assign n639 = x4 & n115 ;
  assign n640 = ~n35 & n639 ;
  assign n641 = ~n48 & ~n640 ;
  assign n642 = ~x7 & ~n641 ;
  assign n651 = ~x0 & ~x8 ;
  assign n657 = n44 & n651 ;
  assign n656 = n44 & n284 ;
  assign n658 = n657 ^ n656 ;
  assign n652 = x9 & n651 ;
  assign n653 = x2 & ~x5 ;
  assign n654 = ~x6 & ~n653 ;
  assign n655 = n652 & ~n654 ;
  assign n659 = n658 ^ n655 ;
  assign n660 = x9 & n317 ;
  assign n664 = x6 & n660 ;
  assign n665 = ~n659 & n664 ;
  assign n666 = n665 ^ n659 ;
  assign n661 = n17 & ~n453 ;
  assign n662 = ~n660 & n661 ;
  assign n663 = ~n659 & n662 ;
  assign n667 = n666 ^ n663 ;
  assign n668 = x1 & ~n667 ;
  assign n643 = x2 & x8 ;
  assign n644 = n41 & n643 ;
  assign n645 = ~x0 & ~n155 ;
  assign n646 = ~x2 & ~x9 ;
  assign n647 = ~n231 & n646 ;
  assign n648 = ~n645 & n647 ;
  assign n649 = ~n644 & ~n648 ;
  assign n650 = ~x1 & n649 ;
  assign n669 = n668 ^ n650 ;
  assign n694 = n345 & n669 ;
  assign n695 = n694 ^ x7 ;
  assign n673 = ~x0 & ~x6 ;
  assign n675 = n400 & n673 ;
  assign n676 = n675 ^ n673 ;
  assign n674 = n264 & ~n673 ;
  assign n677 = n676 ^ n674 ;
  assign n679 = x1 & n677 ;
  assign n678 = x9 & n677 ;
  assign n680 = n679 ^ n678 ;
  assign n671 = x9 & n224 ;
  assign n670 = n123 & n453 ;
  assign n672 = n671 ^ n670 ;
  assign n681 = n680 ^ n672 ;
  assign n682 = ~x5 & n681 ;
  assign n688 = ~n282 & ~n651 ;
  assign n689 = n57 & n688 ;
  assign n684 = n160 & n356 ;
  assign n683 = n102 & n249 ;
  assign n685 = n684 ^ n683 ;
  assign n686 = n685 ^ n11 ;
  assign n687 = x9 & n686 ;
  assign n690 = n689 ^ n687 ;
  assign n691 = n281 & ~n690 ;
  assign n692 = ~n682 & n691 ;
  assign n693 = n669 & n692 ;
  assign n696 = n695 ^ n693 ;
  assign n703 = x9 ^ x5 ;
  assign n711 = n703 ^ x2 ;
  assign n704 = x5 ^ x1 ;
  assign n705 = n704 ^ x9 ;
  assign n706 = n705 ^ x5 ;
  assign n707 = n706 ^ n703 ;
  assign n708 = ~n703 & n707 ;
  assign n697 = x9 ^ x6 ;
  assign n698 = n697 ^ x2 ;
  assign n699 = ~x6 & ~n698 ;
  assign n700 = n699 ^ x2 ;
  assign n701 = n700 ^ x6 ;
  assign n702 = x2 & ~n701 ;
  assign n709 = n708 ^ n702 ;
  assign n710 = n709 ^ n699 ;
  assign n712 = n711 ^ n710 ;
  assign n714 = n697 ^ x6 ;
  assign n713 = n702 ^ x2 ;
  assign n715 = n714 ^ n713 ;
  assign n716 = ~n712 & n715 ;
  assign n717 = n716 ^ n702 ;
  assign n718 = n717 ^ n700 ;
  assign n719 = n718 ^ x1 ;
  assign n720 = n719 ^ x5 ;
  assign n721 = n720 ^ x9 ;
  assign n722 = n721 ^ n705 ;
  assign n723 = ~x0 & x2 ;
  assign n724 = ~n109 & n723 ;
  assign n727 = x8 & ~n724 ;
  assign n728 = ~n722 & n727 ;
  assign n725 = n242 & ~n724 ;
  assign n726 = n722 & n725 ;
  assign n729 = n728 ^ n726 ;
  assign n730 = n729 ^ x8 ;
  assign n731 = x8 ^ x2 ;
  assign n732 = x6 & ~n446 ;
  assign n733 = ~n731 & n732 ;
  assign n735 = n320 & n453 ;
  assign n734 = n439 & n723 ;
  assign n736 = n735 ^ n734 ;
  assign n737 = ~n733 & ~n736 ;
  assign n740 = x7 & n737 ;
  assign n741 = ~n730 & n740 ;
  assign n742 = n741 ^ x7 ;
  assign n738 = n730 & n737 ;
  assign n739 = n738 ^ n737 ;
  assign n743 = n742 ^ n739 ;
  assign n744 = ~x3 & ~x4 ;
  assign n746 = x2 & n115 ;
  assign n747 = x7 & ~x9 ;
  assign n748 = x8 & ~n747 ;
  assign n749 = n746 & ~n748 ;
  assign n745 = n57 & n71 ;
  assign n750 = n749 ^ n745 ;
  assign n757 = n484 & n750 ;
  assign n751 = n142 & n317 ;
  assign n752 = n751 ^ n453 ;
  assign n753 = ~x2 & x7 ;
  assign n754 = n484 & n753 ;
  assign n755 = n752 & n754 ;
  assign n756 = ~n750 & n755 ;
  assign n758 = n757 ^ n756 ;
  assign n759 = n744 & ~n758 ;
  assign n760 = n743 & n759 ;
  assign n761 = n760 ^ n634 ;
  assign n762 = n696 & n761 ;
  assign n763 = n762 ^ x4 ;
  assign n764 = n642 & ~n763 ;
  assign n765 = n764 ^ n642 ;
  assign n766 = n765 ^ n763 ;
  assign n856 = x8 & n747 ;
  assign n857 = n102 & n856 ;
  assign n855 = n446 & n723 ;
  assign n858 = n857 ^ n855 ;
  assign n859 = n207 & n484 ;
  assign n866 = n858 & n859 ;
  assign n867 = ~x4 & x7 ;
  assign n868 = ~n866 & n867 ;
  assign n869 = n868 ^ x4 ;
  assign n789 = x3 & n229 ;
  assign n790 = n201 & n789 ;
  assign n797 = x8 & n294 ;
  assign n795 = ~x2 & ~x6 ;
  assign n796 = n284 & n795 ;
  assign n798 = n797 ^ n796 ;
  assign n793 = n197 & n723 ;
  assign n794 = n793 ^ n315 ;
  assign n799 = n798 ^ n794 ;
  assign n800 = x3 & n799 ;
  assign n801 = ~n790 & ~n800 ;
  assign n802 = x2 & ~n453 ;
  assign n777 = ~x3 & ~x8 ;
  assign n803 = ~x6 & ~n777 ;
  assign n804 = n802 & ~n803 ;
  assign n805 = n45 & n249 ;
  assign n806 = n805 ^ n316 ;
  assign n807 = n76 ^ x1 ;
  assign n808 = n807 ^ x5 ;
  assign n809 = ~n806 & ~n808 ;
  assign n810 = ~n804 & n809 ;
  assign n811 = n801 & n810 ;
  assign n781 = x3 & ~n302 ;
  assign n782 = ~n317 & ~n781 ;
  assign n783 = ~x6 & ~n782 ;
  assign n784 = ~x3 & n302 ;
  assign n778 = n197 & n777 ;
  assign n785 = x2 & ~n778 ;
  assign n786 = ~n784 & n785 ;
  assign n787 = ~n783 & n786 ;
  assign n772 = ~x6 & n53 ;
  assign n773 = n306 & n772 ;
  assign n771 = x9 & n242 ;
  assign n774 = n773 ^ n771 ;
  assign n770 = ~x9 & n155 ;
  assign n775 = n774 ^ n770 ;
  assign n767 = ~x3 & ~x6 ;
  assign n768 = x8 & n767 ;
  assign n769 = n768 ^ x6 ;
  assign n776 = n775 ^ n769 ;
  assign n779 = ~x2 & ~n778 ;
  assign n780 = ~n776 & n779 ;
  assign n788 = n787 ^ n780 ;
  assign n791 = n104 & ~n790 ;
  assign n792 = n788 & n791 ;
  assign n812 = n811 ^ n792 ;
  assign n813 = n812 ^ x5 ;
  assign n843 = x0 & x3 ;
  assign n844 = x2 & n453 ;
  assign n845 = n843 & n844 ;
  assign n846 = ~n33 & n446 ;
  assign n847 = n44 & ~n843 ;
  assign n848 = n847 ^ x5 ;
  assign n849 = ~n846 & n848 ;
  assign n850 = ~n845 & ~n849 ;
  assign n839 = x8 & n439 ;
  assign n840 = n33 & n839 ;
  assign n851 = n244 & ~n840 ;
  assign n852 = n850 & n851 ;
  assign n824 = ~n92 & ~n116 ;
  assign n827 = ~x0 & x3 ;
  assign n828 = n44 & n827 ;
  assign n829 = ~n824 & n828 ;
  assign n826 = x3 & n44 ;
  assign n830 = n829 ^ n826 ;
  assign n825 = ~x0 & ~n824 ;
  assign n831 = n830 ^ n825 ;
  assign n818 = x8 & n102 ;
  assign n816 = x2 & x5 ;
  assign n817 = n284 & n816 ;
  assign n819 = n818 ^ n817 ;
  assign n814 = n300 & n306 ;
  assign n815 = n814 ^ n306 ;
  assign n820 = n819 ^ n815 ;
  assign n834 = n777 & n820 ;
  assign n835 = n834 ^ x8 ;
  assign n832 = ~x8 & n646 ;
  assign n833 = n92 & n832 ;
  assign n836 = n835 ^ n833 ;
  assign n837 = n831 & ~n836 ;
  assign n821 = ~x3 & n820 ;
  assign n822 = n92 & n646 ;
  assign n823 = ~n821 & ~n822 ;
  assign n838 = n837 ^ n823 ;
  assign n841 = n426 & ~n840 ;
  assign n842 = n838 & n841 ;
  assign n853 = n852 ^ n842 ;
  assign n854 = n853 ^ x6 ;
  assign n860 = ~x4 & ~x7 ;
  assign n861 = n859 & n860 ;
  assign n862 = n858 & n861 ;
  assign n863 = n862 ^ n860 ;
  assign n864 = n854 & n863 ;
  assign n865 = n813 & n864 ;
  assign n870 = n869 ^ n865 ;
  assign n871 = ~x5 & ~x7 ;
  assign n872 = n636 & n871 ;
  assign n873 = ~x6 & n872 ;
  assign n874 = n870 & ~n873 ;
  assign n917 = n320 ^ n157 ;
  assign n918 = ~x2 & ~n22 ;
  assign n919 = ~n140 & n918 ;
  assign n920 = n917 & n919 ;
  assign n921 = n22 & n44 ;
  assign n922 = n921 ^ n387 ;
  assign n923 = ~x0 & n922 ;
  assign n924 = n430 & n808 ;
  assign n925 = n13 & ~n924 ;
  assign n926 = ~n923 & ~n925 ;
  assign n927 = ~n920 & n926 ;
  assign n905 = ~n92 & ~n653 ;
  assign n906 = x1 & x3 ;
  assign n907 = ~n181 & n906 ;
  assign n908 = n907 ^ x1 ;
  assign n909 = ~n905 & n908 ;
  assign n910 = n181 & ~n285 ;
  assign n911 = x9 & n260 ;
  assign n912 = n910 & n911 ;
  assign n913 = n912 ^ x9 ;
  assign n914 = ~n909 & n913 ;
  assign n893 = n13 & n123 ;
  assign n892 = n123 & n574 ;
  assign n894 = n893 ^ n892 ;
  assign n891 = n92 & n247 ;
  assign n895 = n894 ^ n891 ;
  assign n890 = n102 & n157 ;
  assign n896 = n895 ^ n890 ;
  assign n897 = ~x9 & ~n896 ;
  assign n886 = ~n92 & n264 ;
  assign n901 = x8 & ~n886 ;
  assign n902 = n897 & ~n901 ;
  assign n898 = x8 & n282 ;
  assign n899 = n886 & n898 ;
  assign n900 = n897 & ~n899 ;
  assign n903 = n902 ^ n900 ;
  assign n887 = n273 & n886 ;
  assign n888 = n887 ^ x8 ;
  assign n889 = ~x9 & ~n888 ;
  assign n904 = n903 ^ n889 ;
  assign n915 = n914 ^ n904 ;
  assign n928 = n292 & n915 ;
  assign n929 = ~n927 & n928 ;
  assign n916 = ~x6 & ~n915 ;
  assign n930 = n929 ^ n916 ;
  assign n933 = x1 & x6 ;
  assign n934 = ~n242 & n933 ;
  assign n932 = ~x9 & n417 ;
  assign n935 = n934 ^ n932 ;
  assign n931 = n201 & n242 ;
  assign n936 = n935 ^ n931 ;
  assign n937 = n591 & ~n936 ;
  assign n938 = n937 ^ n88 ;
  assign n940 = n123 & ~n453 ;
  assign n941 = n940 ^ x0 ;
  assign n942 = ~x6 & ~x7 ;
  assign n943 = ~n11 & n942 ;
  assign n944 = ~n941 & n943 ;
  assign n945 = n938 & n944 ;
  assign n939 = ~x7 & ~n938 ;
  assign n946 = n945 ^ n939 ;
  assign n950 = ~x4 & ~n872 ;
  assign n952 = n946 & n950 ;
  assign n953 = ~n930 & n952 ;
  assign n951 = ~x7 & n950 ;
  assign n954 = n953 ^ n951 ;
  assign n955 = n954 ^ n872 ;
  assign n880 = ~x0 & n229 ;
  assign n881 = n142 & n880 ;
  assign n876 = ~x9 & n181 ;
  assign n877 = n876 ^ n315 ;
  assign n875 = ~x8 & n723 ;
  assign n878 = n877 ^ n875 ;
  assign n879 = ~x1 & n878 ;
  assign n882 = n881 ^ n879 ;
  assign n883 = n366 & n882 ;
  assign n884 = ~n872 & n883 ;
  assign n947 = n884 & n946 ;
  assign n948 = ~n930 & n947 ;
  assign n885 = x7 & n884 ;
  assign n949 = n948 ^ n885 ;
  assign n956 = n955 ^ n949 ;
  assign n957 = ~x1 & ~n453 ;
  assign n958 = x2 & n553 ;
  assign n959 = n282 & n958 ;
  assign n960 = ~x7 & ~n959 ;
  assign n961 = ~n957 & ~n960 ;
  assign n962 = ~x2 & n207 ;
  assign n963 = ~x7 & ~n962 ;
  assign n964 = x0 & ~n963 ;
  assign n965 = ~x5 & ~n13 ;
  assign n966 = x6 & ~n965 ;
  assign n967 = n491 ^ x4 ;
  assign n968 = x7 & ~n13 ;
  assign n969 = ~n967 & ~n968 ;
  assign n970 = ~n966 & n969 ;
  assign n971 = ~n964 & n970 ;
  assign n972 = ~n961 & n971 ;
  assign n987 = x3 & ~n341 ;
  assign n988 = ~x6 & ~n439 ;
  assign n989 = n242 & ~n988 ;
  assign n990 = n987 & ~n989 ;
  assign n991 = ~n484 & n526 ;
  assign n992 = ~x2 & ~n991 ;
  assign n993 = ~n990 & n992 ;
  assign n981 = ~x5 & ~n302 ;
  assign n994 = n13 & ~n453 ;
  assign n995 = ~n981 & n994 ;
  assign n996 = ~x1 & ~n995 ;
  assign n997 = ~n993 & n996 ;
  assign n998 = n972 & n997 ;
  assign n975 = n242 & n341 ;
  assign n976 = n393 & n975 ;
  assign n973 = n109 & ~n242 ;
  assign n974 = n266 & n973 ;
  assign n977 = n976 ^ n974 ;
  assign n978 = n977 ^ n266 ;
  assign n982 = n550 & n981 ;
  assign n979 = n511 ^ x6 ;
  assign n980 = ~x3 & n979 ;
  assign n983 = n982 ^ n980 ;
  assign n984 = ~n978 & ~n983 ;
  assign n985 = x1 & n984 ;
  assign n986 = n972 & n985 ;
  assign n999 = n998 ^ n986 ;
  assign n1000 = ~x7 & n484 ;
  assign n1001 = x8 & ~n477 ;
  assign n1002 = ~x1 & ~n45 ;
  assign n1003 = x2 & n634 ;
  assign n1004 = ~n1002 & n1003 ;
  assign n1005 = ~n1001 & n1004 ;
  assign n1006 = ~n636 & ~n1005 ;
  assign n1007 = n1000 & ~n1006 ;
  assign y0 = ~n216 ;
  assign y1 = ~n378 ;
  assign y2 = n503 ;
  assign y3 = n626 ;
  assign y4 = n633 ;
  assign y5 = n638 ;
  assign y6 = n766 ;
  assign y7 = n874 ;
  assign y8 = ~n956 ;
  assign y9 = n999 ;
  assign y10 = n1007 ;
endmodule
