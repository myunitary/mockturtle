module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 ;
  assign n33 = x2 & ~x3 ;
  assign n34 = x18 & ~x19 ;
  assign n35 = x30 & ~x31 ;
  assign n36 = x28 & ~x29 ;
  assign n37 = x26 & ~x27 ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = n36 & n37 ;
  assign n40 = ~n38 & ~n39 ;
  assign n41 = n35 & ~n40 ;
  assign n42 = ~n35 & n40 ;
  assign n43 = ~n41 & ~n42 ;
  assign n44 = n34 & ~n43 ;
  assign n45 = ~n34 & n43 ;
  assign n46 = ~n44 & ~n45 ;
  assign n47 = x24 & ~x25 ;
  assign n48 = x22 & ~x23 ;
  assign n49 = x20 & ~x21 ;
  assign n50 = n48 & n49 ;
  assign n51 = ~n48 & ~n49 ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = n47 & ~n52 ;
  assign n54 = ~n47 & n52 ;
  assign n55 = ~n53 & ~n54 ;
  assign n56 = n46 & ~n55 ;
  assign n57 = ~n46 & n55 ;
  assign n58 = ~n56 & ~n57 ;
  assign n59 = n33 & n58 ;
  assign n60 = x4 & ~x5 ;
  assign n61 = x16 & ~x17 ;
  assign n62 = x14 & ~x15 ;
  assign n63 = x12 & ~x13 ;
  assign n64 = n62 & n63 ;
  assign n65 = ~n62 & ~n63 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = n61 & ~n66 ;
  assign n68 = ~n61 & n66 ;
  assign n69 = ~n67 & ~n68 ;
  assign n70 = ~n60 & n69 ;
  assign n71 = n60 & ~n69 ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = x10 & ~x11 ;
  assign n74 = x8 & ~x9 ;
  assign n75 = x6 & ~x7 ;
  assign n76 = n74 & n75 ;
  assign n77 = ~n74 & ~n75 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = n73 & ~n78 ;
  assign n80 = ~n73 & n78 ;
  assign n81 = ~n79 & ~n80 ;
  assign n82 = n72 & ~n81 ;
  assign n83 = ~n72 & n81 ;
  assign n84 = ~n82 & ~n83 ;
  assign n85 = ~n33 & ~n58 ;
  assign n86 = ~n59 & ~n85 ;
  assign n87 = n84 & n86 ;
  assign n88 = ~n59 & ~n87 ;
  assign n89 = ~n44 & ~n56 ;
  assign n90 = ~n35 & ~n39 ;
  assign n91 = ~n38 & ~n90 ;
  assign n92 = n89 & ~n91 ;
  assign n93 = ~n89 & n91 ;
  assign n94 = ~n92 & ~n93 ;
  assign n95 = ~n47 & ~n50 ;
  assign n96 = ~n51 & ~n95 ;
  assign n97 = n94 & n96 ;
  assign n98 = ~n94 & ~n96 ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = n88 & ~n99 ;
  assign n101 = ~n88 & n99 ;
  assign n102 = ~n71 & ~n82 ;
  assign n103 = ~n61 & ~n64 ;
  assign n104 = ~n65 & ~n103 ;
  assign n105 = ~n102 & n104 ;
  assign n106 = n102 & ~n104 ;
  assign n107 = ~n105 & ~n106 ;
  assign n108 = ~n73 & ~n76 ;
  assign n109 = ~n77 & ~n108 ;
  assign n110 = n107 & n109 ;
  assign n111 = ~n107 & ~n109 ;
  assign n112 = ~n110 & ~n111 ;
  assign n113 = ~n101 & ~n112 ;
  assign n114 = ~n100 & ~n113 ;
  assign n115 = ~n93 & ~n97 ;
  assign n116 = ~n114 & n115 ;
  assign n117 = n114 & ~n115 ;
  assign n118 = ~n116 & ~n117 ;
  assign n119 = ~n105 & ~n110 ;
  assign n120 = n118 & n119 ;
  assign n121 = ~n116 & ~n120 ;
  assign n122 = ~n118 & ~n119 ;
  assign n123 = ~n120 & ~n122 ;
  assign n124 = x0 & ~x1 ;
  assign n125 = ~n84 & ~n86 ;
  assign n126 = ~n87 & ~n125 ;
  assign n127 = n124 & n126 ;
  assign n128 = ~n100 & ~n101 ;
  assign n129 = ~n112 & n128 ;
  assign n130 = n112 & ~n128 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = n127 & ~n131 ;
  assign n133 = ~n123 & n132 ;
  assign n134 = n121 & n133 ;
  assign n135 = ~x28 & ~x29 ;
  assign n136 = ~x26 & ~x27 ;
  assign n137 = ~n135 & ~n136 ;
  assign n138 = ~x30 & ~x31 ;
  assign n139 = n135 & n136 ;
  assign n140 = ~n137 & ~n139 ;
  assign n141 = ~n138 & n140 ;
  assign n142 = ~n137 & ~n141 ;
  assign n143 = n138 & ~n140 ;
  assign n144 = ~n141 & ~n143 ;
  assign n145 = ~x18 & ~x19 ;
  assign n146 = ~n144 & n145 ;
  assign n147 = n144 & ~n145 ;
  assign n148 = ~x24 & ~x25 ;
  assign n149 = ~x22 & ~x23 ;
  assign n150 = ~x20 & ~x21 ;
  assign n151 = ~n149 & ~n150 ;
  assign n152 = n149 & n150 ;
  assign n153 = ~n151 & ~n152 ;
  assign n154 = ~n148 & n153 ;
  assign n155 = n148 & ~n153 ;
  assign n156 = ~n154 & ~n155 ;
  assign n157 = ~n147 & ~n156 ;
  assign n158 = ~n146 & ~n157 ;
  assign n159 = ~n142 & n158 ;
  assign n160 = ~n151 & ~n154 ;
  assign n161 = n142 & ~n158 ;
  assign n162 = ~n159 & ~n161 ;
  assign n163 = ~n160 & n162 ;
  assign n164 = ~n159 & ~n163 ;
  assign n165 = n160 & ~n162 ;
  assign n166 = ~n163 & ~n165 ;
  assign n167 = ~x2 & ~x3 ;
  assign n168 = ~n146 & ~n147 ;
  assign n169 = n156 & n168 ;
  assign n170 = ~n156 & ~n168 ;
  assign n171 = ~n169 & ~n170 ;
  assign n172 = n167 & ~n171 ;
  assign n173 = ~n167 & n171 ;
  assign n174 = ~x10 & ~x11 ;
  assign n175 = ~x8 & ~x9 ;
  assign n176 = ~x6 & ~x7 ;
  assign n177 = ~n175 & ~n176 ;
  assign n178 = n175 & n176 ;
  assign n179 = ~n177 & ~n178 ;
  assign n180 = ~n174 & n179 ;
  assign n181 = n174 & ~n179 ;
  assign n182 = ~n180 & ~n181 ;
  assign n183 = ~x16 & ~x17 ;
  assign n184 = ~x14 & ~x15 ;
  assign n185 = ~x12 & ~x13 ;
  assign n186 = ~n184 & ~n185 ;
  assign n187 = n184 & n185 ;
  assign n188 = ~n186 & ~n187 ;
  assign n189 = ~n183 & n188 ;
  assign n190 = n183 & ~n188 ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = ~x4 & ~x5 ;
  assign n193 = n191 & ~n192 ;
  assign n194 = ~n191 & n192 ;
  assign n195 = ~n193 & ~n194 ;
  assign n196 = n182 & n195 ;
  assign n197 = ~n182 & ~n195 ;
  assign n198 = ~n196 & ~n197 ;
  assign n199 = ~n173 & ~n198 ;
  assign n200 = ~n172 & ~n199 ;
  assign n201 = ~n166 & ~n200 ;
  assign n202 = n166 & n200 ;
  assign n203 = ~n186 & ~n189 ;
  assign n204 = ~n193 & ~n196 ;
  assign n205 = n203 & n204 ;
  assign n206 = ~n203 & ~n204 ;
  assign n207 = ~n205 & ~n206 ;
  assign n208 = ~n177 & ~n180 ;
  assign n209 = ~n207 & n208 ;
  assign n210 = n207 & ~n208 ;
  assign n211 = ~n209 & ~n210 ;
  assign n212 = ~n202 & ~n211 ;
  assign n213 = ~n201 & ~n212 ;
  assign n214 = n164 & ~n213 ;
  assign n215 = ~x0 & ~x1 ;
  assign n216 = ~n172 & ~n173 ;
  assign n217 = n198 & n216 ;
  assign n218 = ~n198 & ~n216 ;
  assign n219 = ~n217 & ~n218 ;
  assign n220 = n215 & ~n219 ;
  assign n221 = ~n201 & ~n202 ;
  assign n222 = ~n211 & n221 ;
  assign n223 = n211 & ~n221 ;
  assign n224 = ~n222 & ~n223 ;
  assign n225 = n220 & n224 ;
  assign n226 = ~n206 & ~n210 ;
  assign n227 = ~n164 & n213 ;
  assign n228 = ~n214 & ~n227 ;
  assign n229 = n226 & n228 ;
  assign n230 = ~n226 & ~n228 ;
  assign n231 = ~n229 & ~n230 ;
  assign n232 = n225 & n231 ;
  assign n233 = n214 & n232 ;
  assign n234 = n134 & ~n233 ;
  assign n235 = ~n121 & ~n133 ;
  assign n236 = ~n134 & ~n235 ;
  assign n237 = ~n214 & ~n229 ;
  assign n238 = ~n232 & n237 ;
  assign n239 = ~n233 & ~n238 ;
  assign n240 = n236 & ~n239 ;
  assign n241 = ~n225 & ~n231 ;
  assign n242 = ~n232 & ~n241 ;
  assign n243 = ~n215 & n219 ;
  assign n244 = ~n220 & ~n243 ;
  assign n245 = ~n124 & ~n126 ;
  assign n246 = ~n127 & ~n245 ;
  assign n247 = n244 & ~n246 ;
  assign n248 = n224 & n247 ;
  assign n249 = ~n127 & n131 ;
  assign n250 = ~n132 & ~n249 ;
  assign n251 = ~n220 & ~n224 ;
  assign n252 = ~n225 & ~n251 ;
  assign n253 = ~n247 & ~n252 ;
  assign n254 = ~n250 & ~n253 ;
  assign n255 = ~n248 & ~n254 ;
  assign n256 = n242 & ~n255 ;
  assign n257 = n123 & ~n132 ;
  assign n258 = ~n133 & ~n257 ;
  assign n259 = ~n242 & n255 ;
  assign n260 = ~n258 & ~n259 ;
  assign n261 = ~n256 & ~n260 ;
  assign n262 = ~n240 & ~n261 ;
  assign n263 = ~n134 & n233 ;
  assign n264 = ~n236 & n239 ;
  assign n265 = ~n263 & ~n264 ;
  assign n266 = ~n262 & n265 ;
  assign n267 = ~n234 & ~n266 ;
  assign n268 = ~n134 & ~n233 ;
  assign n269 = ~x18 & x19 ;
  assign n270 = ~x30 & x31 ;
  assign n271 = ~x28 & x29 ;
  assign n272 = ~x26 & x27 ;
  assign n273 = ~n271 & ~n272 ;
  assign n274 = n271 & n272 ;
  assign n275 = ~n273 & ~n274 ;
  assign n276 = n270 & ~n275 ;
  assign n277 = ~n270 & n275 ;
  assign n278 = ~n276 & ~n277 ;
  assign n279 = n269 & ~n278 ;
  assign n280 = ~n269 & n278 ;
  assign n281 = ~x24 & x25 ;
  assign n282 = ~x22 & x23 ;
  assign n283 = ~x20 & x21 ;
  assign n284 = ~n282 & ~n283 ;
  assign n285 = n282 & n283 ;
  assign n286 = ~n284 & ~n285 ;
  assign n287 = n281 & ~n286 ;
  assign n288 = ~n281 & n286 ;
  assign n289 = ~n287 & ~n288 ;
  assign n290 = ~n280 & ~n289 ;
  assign n291 = ~n279 & ~n290 ;
  assign n292 = ~n270 & ~n274 ;
  assign n293 = ~n273 & ~n292 ;
  assign n294 = ~n291 & n293 ;
  assign n295 = n291 & ~n293 ;
  assign n296 = ~n294 & ~n295 ;
  assign n297 = ~n281 & ~n285 ;
  assign n298 = ~n284 & ~n297 ;
  assign n299 = n296 & n298 ;
  assign n300 = ~n294 & ~n299 ;
  assign n301 = ~n296 & ~n298 ;
  assign n302 = ~n299 & ~n301 ;
  assign n303 = ~x2 & x3 ;
  assign n304 = ~n279 & ~n280 ;
  assign n305 = n289 & n304 ;
  assign n306 = ~n289 & ~n304 ;
  assign n307 = ~n305 & ~n306 ;
  assign n308 = n303 & ~n307 ;
  assign n309 = ~n303 & n307 ;
  assign n310 = ~x4 & x5 ;
  assign n311 = ~x16 & x17 ;
  assign n312 = ~x14 & x15 ;
  assign n313 = ~x12 & x13 ;
  assign n314 = n312 & n313 ;
  assign n315 = ~n312 & ~n313 ;
  assign n316 = ~n314 & ~n315 ;
  assign n317 = n311 & ~n316 ;
  assign n318 = ~n311 & n316 ;
  assign n319 = ~n317 & ~n318 ;
  assign n320 = n310 & ~n319 ;
  assign n321 = ~n310 & n319 ;
  assign n322 = ~n320 & ~n321 ;
  assign n323 = ~x10 & x11 ;
  assign n324 = ~x8 & x9 ;
  assign n325 = ~x6 & x7 ;
  assign n326 = n324 & n325 ;
  assign n327 = ~n324 & ~n325 ;
  assign n328 = ~n326 & ~n327 ;
  assign n329 = n323 & ~n328 ;
  assign n330 = ~n323 & n328 ;
  assign n331 = ~n329 & ~n330 ;
  assign n332 = n322 & ~n331 ;
  assign n333 = ~n322 & n331 ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = ~n309 & n334 ;
  assign n336 = ~n308 & ~n335 ;
  assign n337 = n302 & ~n336 ;
  assign n338 = ~n302 & n336 ;
  assign n339 = ~n320 & ~n332 ;
  assign n340 = ~n311 & ~n314 ;
  assign n341 = ~n315 & ~n340 ;
  assign n342 = n339 & ~n341 ;
  assign n343 = ~n339 & n341 ;
  assign n344 = ~n342 & ~n343 ;
  assign n345 = ~n323 & ~n326 ;
  assign n346 = ~n327 & ~n345 ;
  assign n347 = n344 & n346 ;
  assign n348 = ~n344 & ~n346 ;
  assign n349 = ~n347 & ~n348 ;
  assign n350 = ~n338 & n349 ;
  assign n351 = ~n337 & ~n350 ;
  assign n352 = n300 & n351 ;
  assign n353 = ~n300 & ~n351 ;
  assign n354 = ~n352 & ~n353 ;
  assign n355 = ~n343 & ~n347 ;
  assign n356 = n354 & n355 ;
  assign n357 = ~n354 & ~n355 ;
  assign n358 = ~n356 & ~n357 ;
  assign n359 = ~x0 & x1 ;
  assign n360 = ~n308 & ~n309 ;
  assign n361 = n334 & n360 ;
  assign n362 = ~n334 & ~n360 ;
  assign n363 = ~n361 & ~n362 ;
  assign n364 = n359 & n363 ;
  assign n365 = ~n337 & ~n338 ;
  assign n366 = n349 & n365 ;
  assign n367 = ~n349 & ~n365 ;
  assign n368 = ~n366 & ~n367 ;
  assign n369 = n364 & n368 ;
  assign n370 = ~n358 & n369 ;
  assign n371 = ~n352 & ~n356 ;
  assign n372 = n370 & n371 ;
  assign n373 = x2 & x3 ;
  assign n374 = x18 & x19 ;
  assign n375 = x30 & x31 ;
  assign n376 = x28 & x29 ;
  assign n377 = x26 & x27 ;
  assign n378 = ~n376 & ~n377 ;
  assign n379 = n376 & n377 ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = n375 & ~n380 ;
  assign n382 = ~n375 & n380 ;
  assign n383 = ~n381 & ~n382 ;
  assign n384 = n374 & ~n383 ;
  assign n385 = ~n374 & n383 ;
  assign n386 = ~n384 & ~n385 ;
  assign n387 = x24 & x25 ;
  assign n388 = x22 & x23 ;
  assign n389 = x20 & x21 ;
  assign n390 = n388 & n389 ;
  assign n391 = ~n388 & ~n389 ;
  assign n392 = ~n390 & ~n391 ;
  assign n393 = n387 & ~n392 ;
  assign n394 = ~n387 & n392 ;
  assign n395 = ~n393 & ~n394 ;
  assign n396 = n386 & ~n395 ;
  assign n397 = ~n386 & n395 ;
  assign n398 = ~n396 & ~n397 ;
  assign n399 = n373 & n398 ;
  assign n400 = x4 & x5 ;
  assign n401 = x16 & x17 ;
  assign n402 = x14 & x15 ;
  assign n403 = x12 & x13 ;
  assign n404 = n402 & n403 ;
  assign n405 = ~n402 & ~n403 ;
  assign n406 = ~n404 & ~n405 ;
  assign n407 = n401 & ~n406 ;
  assign n408 = ~n401 & n406 ;
  assign n409 = ~n407 & ~n408 ;
  assign n410 = ~n400 & n409 ;
  assign n411 = n400 & ~n409 ;
  assign n412 = ~n410 & ~n411 ;
  assign n413 = x10 & x11 ;
  assign n414 = x8 & x9 ;
  assign n415 = x6 & x7 ;
  assign n416 = n414 & n415 ;
  assign n417 = ~n414 & ~n415 ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = n413 & ~n418 ;
  assign n420 = ~n413 & n418 ;
  assign n421 = ~n419 & ~n420 ;
  assign n422 = n412 & ~n421 ;
  assign n423 = ~n412 & n421 ;
  assign n424 = ~n422 & ~n423 ;
  assign n425 = ~n373 & ~n398 ;
  assign n426 = ~n399 & ~n425 ;
  assign n427 = n424 & n426 ;
  assign n428 = ~n399 & ~n427 ;
  assign n429 = ~n384 & ~n396 ;
  assign n430 = ~n375 & ~n379 ;
  assign n431 = ~n378 & ~n430 ;
  assign n432 = n429 & ~n431 ;
  assign n433 = ~n429 & n431 ;
  assign n434 = ~n432 & ~n433 ;
  assign n435 = ~n387 & ~n390 ;
  assign n436 = ~n391 & ~n435 ;
  assign n437 = n434 & n436 ;
  assign n438 = ~n434 & ~n436 ;
  assign n439 = ~n437 & ~n438 ;
  assign n440 = n428 & ~n439 ;
  assign n441 = ~n428 & n439 ;
  assign n442 = ~n411 & ~n422 ;
  assign n443 = ~n401 & ~n404 ;
  assign n444 = ~n405 & ~n443 ;
  assign n445 = ~n442 & n444 ;
  assign n446 = n442 & ~n444 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = ~n413 & ~n416 ;
  assign n449 = ~n417 & ~n448 ;
  assign n450 = n447 & n449 ;
  assign n451 = ~n447 & ~n449 ;
  assign n452 = ~n450 & ~n451 ;
  assign n453 = ~n441 & ~n452 ;
  assign n454 = ~n440 & ~n453 ;
  assign n455 = ~n433 & ~n437 ;
  assign n456 = ~n454 & n455 ;
  assign n457 = n454 & ~n455 ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = ~n445 & ~n450 ;
  assign n460 = n458 & n459 ;
  assign n461 = ~n456 & ~n460 ;
  assign n462 = ~n458 & ~n459 ;
  assign n463 = ~n460 & ~n462 ;
  assign n464 = x0 & x1 ;
  assign n465 = ~n424 & ~n426 ;
  assign n466 = ~n427 & ~n465 ;
  assign n467 = n464 & n466 ;
  assign n468 = ~n440 & ~n441 ;
  assign n469 = ~n452 & n468 ;
  assign n470 = n452 & ~n468 ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = n467 & ~n471 ;
  assign n473 = ~n463 & n472 ;
  assign n474 = n461 & n473 ;
  assign n475 = ~n372 & ~n474 ;
  assign n476 = n268 & ~n475 ;
  assign n477 = ~n467 & n471 ;
  assign n478 = ~n472 & ~n477 ;
  assign n479 = ~n372 & n474 ;
  assign n480 = ~n461 & ~n473 ;
  assign n481 = ~n474 & ~n480 ;
  assign n482 = ~n370 & ~n371 ;
  assign n483 = ~n372 & ~n482 ;
  assign n484 = n481 & ~n483 ;
  assign n485 = n358 & ~n369 ;
  assign n486 = ~n370 & ~n485 ;
  assign n487 = ~n359 & ~n363 ;
  assign n488 = ~n364 & ~n487 ;
  assign n489 = ~n464 & ~n466 ;
  assign n490 = ~n467 & ~n489 ;
  assign n491 = n488 & ~n490 ;
  assign n492 = n368 & n491 ;
  assign n493 = ~n364 & ~n368 ;
  assign n494 = ~n369 & ~n493 ;
  assign n495 = ~n491 & ~n494 ;
  assign n496 = ~n478 & ~n495 ;
  assign n497 = ~n492 & ~n496 ;
  assign n498 = ~n486 & n497 ;
  assign n499 = n463 & ~n472 ;
  assign n500 = ~n473 & ~n499 ;
  assign n501 = n486 & ~n497 ;
  assign n502 = n500 & ~n501 ;
  assign n503 = ~n498 & ~n502 ;
  assign n504 = ~n484 & n503 ;
  assign n505 = n372 & ~n474 ;
  assign n506 = ~n481 & n483 ;
  assign n507 = ~n505 & ~n506 ;
  assign n508 = ~n504 & n507 ;
  assign n509 = ~n479 & ~n508 ;
  assign n510 = ~n478 & ~n509 ;
  assign n511 = ~n494 & n509 ;
  assign n512 = ~n510 & ~n511 ;
  assign n513 = ~n252 & n267 ;
  assign n514 = ~n250 & ~n267 ;
  assign n515 = ~n513 & ~n514 ;
  assign n516 = n512 & ~n515 ;
  assign n517 = ~n490 & ~n509 ;
  assign n518 = ~n488 & n509 ;
  assign n519 = ~n517 & ~n518 ;
  assign n520 = ~n244 & n267 ;
  assign n521 = ~n246 & ~n267 ;
  assign n522 = ~n520 & ~n521 ;
  assign n523 = ~n519 & n522 ;
  assign n524 = ~n516 & n523 ;
  assign n525 = n486 & n509 ;
  assign n526 = n500 & ~n509 ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = n242 & n267 ;
  assign n529 = n258 & ~n267 ;
  assign n530 = ~n528 & ~n529 ;
  assign n531 = n527 & ~n530 ;
  assign n532 = ~n512 & n515 ;
  assign n533 = ~n531 & ~n532 ;
  assign n534 = ~n524 & n533 ;
  assign n535 = n235 & n238 ;
  assign n536 = n268 & ~n535 ;
  assign n537 = n480 & n482 ;
  assign n538 = n475 & ~n537 ;
  assign n539 = ~n536 & n538 ;
  assign n540 = ~n527 & n530 ;
  assign n541 = ~n539 & ~n540 ;
  assign n542 = ~n534 & n541 ;
  assign n543 = ~n268 & n475 ;
  assign n544 = n536 & ~n538 ;
  assign n545 = ~n543 & ~n544 ;
  assign n546 = ~n542 & n545 ;
  assign n547 = ~n476 & ~n546 ;
  assign n548 = ~n267 & n547 ;
  assign n549 = ~n509 & ~n547 ;
  assign n550 = ~n548 & ~n549 ;
  assign y0 = ~n550 ;
  assign y1 = ~n547 ;
endmodule
