module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
  assign n17 = x13 & x14 ;
  assign n18 = ~x13 & ~x14 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = x15 & n19 ;
  assign n21 = ~n17 & ~n20 ;
  assign n22 = ~x15 & ~n19 ;
  assign n23 = ~n20 & ~n22 ;
  assign n24 = x9 & n23 ;
  assign n25 = ~x9 & ~n23 ;
  assign n26 = ~x10 & ~x11 ;
  assign n27 = x10 & x11 ;
  assign n28 = ~n26 & ~n27 ;
  assign n29 = x12 & n28 ;
  assign n30 = ~x12 & ~n28 ;
  assign n31 = ~n29 & ~n30 ;
  assign n32 = ~n25 & n31 ;
  assign n33 = ~n24 & ~n32 ;
  assign n34 = ~n21 & ~n33 ;
  assign n35 = ~n27 & ~n29 ;
  assign n36 = n21 & n33 ;
  assign n37 = ~n34 & ~n36 ;
  assign n38 = ~n35 & n37 ;
  assign n39 = ~n34 & ~n38 ;
  assign n40 = n35 & ~n37 ;
  assign n41 = ~n38 & ~n40 ;
  assign n42 = ~n24 & ~n25 ;
  assign n43 = n31 & ~n42 ;
  assign n44 = ~n31 & n42 ;
  assign n45 = ~n43 & ~n44 ;
  assign n46 = ~x1 & n45 ;
  assign n47 = x1 & ~n45 ;
  assign n48 = ~x3 & ~x4 ;
  assign n49 = x3 & x4 ;
  assign n50 = ~n48 & ~n49 ;
  assign n51 = x5 & n50 ;
  assign n52 = ~x5 & ~n50 ;
  assign n53 = ~n51 & ~n52 ;
  assign n54 = ~x6 & ~x7 ;
  assign n55 = x6 & x7 ;
  assign n56 = ~n54 & ~n55 ;
  assign n57 = x8 & n56 ;
  assign n58 = ~x8 & ~n56 ;
  assign n59 = ~n57 & ~n58 ;
  assign n60 = x2 & n59 ;
  assign n61 = ~x2 & ~n59 ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = n53 & n62 ;
  assign n64 = ~n53 & ~n62 ;
  assign n65 = ~n63 & ~n64 ;
  assign n66 = ~n47 & ~n65 ;
  assign n67 = ~n46 & ~n66 ;
  assign n68 = ~n41 & ~n67 ;
  assign n69 = n41 & n67 ;
  assign n70 = ~n49 & ~n51 ;
  assign n71 = ~n55 & ~n57 ;
  assign n72 = ~n60 & ~n63 ;
  assign n73 = n71 & n72 ;
  assign n74 = ~n71 & ~n72 ;
  assign n75 = ~n73 & ~n74 ;
  assign n76 = ~n70 & n75 ;
  assign n77 = n70 & ~n75 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = ~n69 & ~n78 ;
  assign n80 = ~n68 & ~n79 ;
  assign n81 = n39 & ~n80 ;
  assign n82 = ~n74 & ~n76 ;
  assign n83 = n81 & n82 ;
  assign n84 = ~n68 & ~n69 ;
  assign n85 = ~n78 & n84 ;
  assign n86 = n78 & ~n84 ;
  assign n87 = ~n85 & ~n86 ;
  assign n88 = ~n46 & ~n47 ;
  assign n89 = ~n65 & ~n88 ;
  assign n90 = n65 & n88 ;
  assign n91 = x0 & ~n90 ;
  assign n92 = ~n89 & n91 ;
  assign n93 = ~n87 & n92 ;
  assign n94 = ~n83 & n93 ;
  assign n95 = ~n39 & n80 ;
  assign n96 = n82 & ~n95 ;
  assign n97 = ~n81 & ~n96 ;
  assign n98 = ~n94 & ~n97 ;
  assign y0 = ~n98 ;
endmodule
