module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511;
output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129;
wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418, y127, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, y129, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y128;
assign n_0 = x0 & ~x128;
assign n_1 = x128 ^ x0;
assign n_2 = x129 ^ x1;
assign n_3 = x130 ^ x2;
assign n_4 = x131 ^ x3;
assign n_5 = x132 ^ x4;
assign n_6 = x133 ^ x5;
assign n_7 = x134 ^ x6;
assign n_8 = x135 ^ x7;
assign n_9 = x136 ^ x8;
assign n_10 = x137 ^ x9;
assign n_11 = x138 ^ x10;
assign n_12 = x139 ^ x11;
assign n_13 = x140 ^ x12;
assign n_14 = x141 ^ x13;
assign n_15 = x142 ^ x14;
assign n_16 = x143 ^ x15;
assign n_17 = x144 ^ x16;
assign n_18 = x145 ^ x17;
assign n_19 = x146 ^ x18;
assign n_20 = x147 ^ x19;
assign n_21 = x148 ^ x20;
assign n_22 = x149 ^ x21;
assign n_23 = x150 ^ x22;
assign n_24 = x151 ^ x23;
assign n_25 = x152 ^ x24;
assign n_26 = x153 ^ x25;
assign n_27 = x154 ^ x26;
assign n_28 = x155 ^ x27;
assign n_29 = x156 ^ x28;
assign n_30 = x157 ^ x29;
assign n_31 = x158 ^ x30;
assign n_32 = x159 ^ x31;
assign n_33 = x160 ^ x32;
assign n_34 = x161 ^ x33;
assign n_35 = x162 ^ x34;
assign n_36 = x163 ^ x35;
assign n_37 = x164 ^ x36;
assign n_38 = x165 ^ x37;
assign n_39 = x166 ^ x38;
assign n_40 = ~x39 & x167;
assign n_41 = x167 ^ x39;
assign n_42 = x40 & ~x168;
assign n_43 = x168 ^ x40;
assign n_44 = ~x41 ^ x169;
assign n_45 = x169 ^ x41;
assign n_46 = ~x42 ^ x170;
assign n_47 = x170 ^ x42;
assign n_48 = ~x43 & x171;
assign n_49 = x171 ^ x43;
assign n_50 = x44 & ~x172;
assign n_51 = x172 ^ x44;
assign n_52 = ~x45 ^ x173;
assign n_53 = x173 ^ x45;
assign n_54 = ~x46 ^ x174;
assign n_55 = x174 ^ x46;
assign n_56 = ~x47 & x175;
assign n_57 = x175 ^ x47;
assign n_58 = ~x48 & x176;
assign n_59 = x176 ^ x48;
assign n_60 = x177 ^ x49;
assign n_61 = x178 ^ x50;
assign n_62 = x179 ^ x51;
assign n_63 = x180 ^ x52;
assign n_64 = x181 ^ x53;
assign n_65 = x182 ^ x54;
assign n_66 = x183 ^ x55;
assign n_67 = x184 ^ x56;
assign n_68 = x185 ^ x57;
assign n_69 = x186 ^ x58;
assign n_70 = x59 & ~x187;
assign n_71 = x187 ^ x59;
assign n_72 = x60 & ~x188;
assign n_73 = x188 ^ x60;
assign n_74 = ~x61 ^ x189;
assign n_75 = x189 ^ x61;
assign n_76 = ~x62 ^ x190;
assign n_77 = x190 ^ x62;
assign n_78 = x63 & ~x191;
assign n_79 = x191 ^ x63;
assign n_80 = x192 ^ x64;
assign n_81 = x193 ^ x65;
assign n_82 = x194 ^ x66;
assign n_83 = x195 ^ x67;
assign n_84 = x68 & ~x196;
assign n_85 = x196 ^ x68;
assign n_86 = ~x69 ^ x197;
assign n_87 = x197 ^ x69;
assign n_88 = ~x70 ^ x198;
assign n_89 = x198 ^ x70;
assign n_90 = ~x71 & x199;
assign n_91 = x199 ^ x71;
assign n_92 = x72 & ~x200;
assign n_93 = x200 ^ x72;
assign n_94 = ~x73 & x201;
assign n_95 = x201 ^ x73;
assign n_96 = x74 & ~x202;
assign n_97 = x202 ^ x74;
assign n_98 = ~x75 & x203;
assign n_99 = x203 ^ x75;
assign n_100 = x76 & ~x204;
assign n_101 = x204 ^ x76;
assign n_102 = ~x77 & x205;
assign n_103 = x205 ^ x77;
assign n_104 = x78 & ~x206;
assign n_105 = x206 ^ x78;
assign n_106 = ~x79 & x207;
assign n_107 = x207 ^ x79;
assign n_108 = ~x80 & x208;
assign n_109 = x208 ^ x80;
assign n_110 = x209 ^ x81;
assign n_111 = x210 ^ x82;
assign n_112 = x211 ^ x83;
assign n_113 = x212 ^ x84;
assign n_114 = x213 ^ x85;
assign n_115 = x214 ^ x86;
assign n_116 = x215 ^ x87;
assign n_117 = x216 ^ x88;
assign n_118 = x217 ^ x89;
assign n_119 = x218 ^ x90;
assign n_120 = x219 ^ x91;
assign n_121 = x220 ^ x92;
assign n_122 = x221 ^ x93;
assign n_123 = x222 ^ x94;
assign n_124 = x223 ^ x95;
assign n_125 = x224 ^ x96;
assign n_126 = x225 ^ x97;
assign n_127 = x226 ^ x98;
assign n_128 = x227 ^ x99;
assign n_129 = x228 ^ x100;
assign n_130 = x229 ^ x101;
assign n_131 = x230 ^ x102;
assign n_132 = x231 ^ x103;
assign n_133 = x232 ^ x104;
assign n_134 = x233 ^ x105;
assign n_135 = x234 ^ x106;
assign n_136 = x235 ^ x107;
assign n_137 = x236 ^ x108;
assign n_138 = x237 ^ x109;
assign n_139 = x238 ^ x110;
assign n_140 = x239 ^ x111;
assign n_141 = x240 ^ x112;
assign n_142 = x241 ^ x113;
assign n_143 = x242 ^ x114;
assign n_144 = x243 ^ x115;
assign n_145 = x244 ^ x116;
assign n_146 = x245 ^ x117;
assign n_147 = x246 ^ x118;
assign n_148 = x247 ^ x119;
assign n_149 = x248 ^ x120;
assign n_150 = x249 ^ x121;
assign n_151 = x250 ^ x122;
assign n_152 = x123 & ~x251;
assign n_153 = x251 ^ x123;
assign n_154 = ~x124 & x252;
assign n_155 = x252 ^ x124;
assign n_156 = x253 ^ x125;
assign n_157 = ~x125 ^ x253;
assign n_158 = x254 ^ x126;
assign n_159 = ~x126 ^ x254;
assign n_160 = x127 & x255;
assign n_161 = x255 ^ x127;
assign n_162 = x256 & ~x384;
assign n_163 = x384 ^ x256;
assign n_164 = x385 ^ x257;
assign n_165 = x386 ^ x258;
assign n_166 = x387 ^ x259;
assign n_167 = x388 ^ x260;
assign n_168 = x389 ^ x261;
assign n_169 = x390 ^ x262;
assign n_170 = x391 ^ x263;
assign n_171 = x392 ^ x264;
assign n_172 = x393 ^ x265;
assign n_173 = x394 ^ x266;
assign n_174 = x395 ^ x267;
assign n_175 = x396 ^ x268;
assign n_176 = x397 ^ x269;
assign n_177 = x398 ^ x270;
assign n_178 = x399 ^ x271;
assign n_179 = x400 ^ x272;
assign n_180 = x401 ^ x273;
assign n_181 = x402 ^ x274;
assign n_182 = x403 ^ x275;
assign n_183 = x404 ^ x276;
assign n_184 = x405 ^ x277;
assign n_185 = x406 ^ x278;
assign n_186 = x407 ^ x279;
assign n_187 = x408 ^ x280;
assign n_188 = x409 ^ x281;
assign n_189 = x410 ^ x282;
assign n_190 = x411 ^ x283;
assign n_191 = x412 ^ x284;
assign n_192 = x413 ^ x285;
assign n_193 = x414 ^ x286;
assign n_194 = x415 ^ x287;
assign n_195 = x416 ^ x288;
assign n_196 = x417 ^ x289;
assign n_197 = x418 ^ x290;
assign n_198 = x419 ^ x291;
assign n_199 = x420 ^ x292;
assign n_200 = x421 ^ x293;
assign n_201 = x422 ^ x294;
assign n_202 = x295 & ~x423;
assign n_203 = x423 ^ x295;
assign n_204 = x296 & ~x424;
assign n_205 = x424 ^ x296;
assign n_206 = ~x297 ^ x425;
assign n_207 = x425 ^ x297;
assign n_208 = ~x298 ^ x426;
assign n_209 = x426 ^ x298;
assign n_210 = ~x299 & x427;
assign n_211 = x427 ^ x299;
assign n_212 = x300 & ~x428;
assign n_213 = x428 ^ x300;
assign n_214 = ~x301 ^ x429;
assign n_215 = x429 ^ x301;
assign n_216 = ~x302 ^ x430;
assign n_217 = x430 ^ x302;
assign n_218 = ~x303 & x431;
assign n_219 = x431 ^ x303;
assign n_220 = x304 & ~x432;
assign n_221 = x432 ^ x304;
assign n_222 = ~x305 & x433;
assign n_223 = x433 ^ x305;
assign n_224 = x306 & ~x434;
assign n_225 = x434 ^ x306;
assign n_226 = x307 & ~x435;
assign n_227 = x435 ^ x307;
assign n_228 = x436 ^ x308;
assign n_229 = x437 ^ x309;
assign n_230 = x438 ^ x310;
assign n_231 = x439 ^ x311;
assign n_232 = x440 ^ x312;
assign n_233 = x441 ^ x313;
assign n_234 = x442 ^ x314;
assign n_235 = ~x315 & x443;
assign n_236 = x443 ^ x315;
assign n_237 = x316 & ~x444;
assign n_238 = x444 ^ x316;
assign n_239 = x317 & ~x445;
assign n_240 = x445 ^ x317;
assign n_241 = x318 & ~x446;
assign n_242 = x446 ^ x318;
assign n_243 = ~x319 & x447;
assign n_244 = x447 ^ x319;
assign n_245 = x320 & ~x448;
assign n_246 = x448 ^ x320;
assign n_247 = x449 ^ x321;
assign n_248 = x450 ^ x322;
assign n_249 = x323 & ~x451;
assign n_250 = x451 ^ x323;
assign n_251 = x324 & ~x452;
assign n_252 = x452 ^ x324;
assign n_253 = ~x325 ^ x453;
assign n_254 = x453 ^ x325;
assign n_255 = ~x326 ^ x454;
assign n_256 = x454 ^ x326;
assign n_257 = x327 & ~x455;
assign n_258 = x455 ^ x327;
assign n_259 = x456 ^ x328;
assign n_260 = x457 ^ x329;
assign n_261 = x458 ^ x330;
assign n_262 = x459 ^ x331;
assign n_263 = x460 ^ x332;
assign n_264 = x461 ^ x333;
assign n_265 = x462 ^ x334;
assign n_266 = x463 ^ x335;
assign n_267 = x464 ^ x336;
assign n_268 = x465 ^ x337;
assign n_269 = x466 ^ x338;
assign n_270 = x467 ^ x339;
assign n_271 = x468 ^ x340;
assign n_272 = x469 ^ x341;
assign n_273 = x470 ^ x342;
assign n_274 = x471 ^ x343;
assign n_275 = x472 ^ x344;
assign n_276 = x473 ^ x345;
assign n_277 = x474 ^ x346;
assign n_278 = x475 ^ x347;
assign n_279 = x476 ^ x348;
assign n_280 = x477 ^ x349;
assign n_281 = x478 ^ x350;
assign n_282 = x479 ^ x351;
assign n_283 = x480 ^ x352;
assign n_284 = x481 ^ x353;
assign n_285 = x482 ^ x354;
assign n_286 = x483 ^ x355;
assign n_287 = x484 ^ x356;
assign n_288 = x485 ^ x357;
assign n_289 = x486 ^ x358;
assign n_290 = x487 ^ x359;
assign n_291 = x488 ^ x360;
assign n_292 = x489 ^ x361;
assign n_293 = x490 ^ x362;
assign n_294 = x491 ^ x363;
assign n_295 = x492 ^ x364;
assign n_296 = x493 ^ x365;
assign n_297 = x494 ^ x366;
assign n_298 = x495 ^ x367;
assign n_299 = x496 ^ x368;
assign n_300 = x497 ^ x369;
assign n_301 = x498 ^ x370;
assign n_302 = x499 ^ x371;
assign n_303 = x500 ^ x372;
assign n_304 = x501 ^ x373;
assign n_305 = x502 ^ x374;
assign n_306 = x503 ^ x375;
assign n_307 = x504 ^ x376;
assign n_308 = x505 ^ x377;
assign n_309 = x506 ^ x378;
assign n_310 = x379 & ~x507;
assign n_311 = x507 ^ x379;
assign n_312 = ~x380 & x508;
assign n_313 = x508 ^ x380;
assign n_314 = x509 ^ x381;
assign n_315 = ~x381 ^ x509;
assign n_316 = x510 ^ x382;
assign n_317 = ~x382 ^ x510;
assign n_318 = x383 & x511;
assign n_319 = x511 ^ x383;
assign n_320 = n_0 ^ x129;
assign n_321 = n_42 ^ x169;
assign n_322 = n_42 ^ n_43;
assign n_323 = n_44 & n_46;
assign n_324 = n_50 ^ x173;
assign n_325 = n_50 ^ n_51;
assign n_326 = n_54 & n_52;
assign n_327 = ~n_58 & ~n_56;
assign n_328 = n_58 ^ n_59;
assign n_329 = n_70 ^ n_71;
assign n_330 = n_72 ^ x189;
assign n_331 = n_72 ^ n_73;
assign n_332 = n_76 & n_74;
assign n_333 = n_78 ^ n_79;
assign n_334 = n_84 ^ x197;
assign n_335 = n_84 ^ n_85;
assign n_336 = n_88 & n_86;
assign n_337 = n_92 ^ n_93;
assign n_338 = n_94 ^ n_95;
assign n_339 = n_96 ^ n_97;
assign n_340 = n_98 ^ n_99;
assign n_341 = n_100 ^ n_101;
assign n_342 = n_102 ^ n_103;
assign n_343 = n_104 ^ n_105;
assign n_344 = n_106 ^ n_107;
assign n_345 = ~n_108 & ~n_106;
assign n_346 = n_108 ^ n_109;
assign n_347 = n_152 ^ n_153;
assign n_348 = n_154 ^ n_155;
assign n_349 = n_157 & n_159;
assign n_350 = n_162 ^ x385;
assign n_351 = n_202 ^ n_203;
assign n_352 = n_204 ^ x425;
assign n_353 = n_204 ^ n_205;
assign n_354 = n_206 & n_208;
assign n_355 = n_212 ^ x429;
assign n_356 = n_212 ^ n_213;
assign n_357 = n_216 & n_214;
assign n_358 = n_220 ^ n_221;
assign n_359 = n_222 ^ n_223;
assign n_360 = n_224 ^ n_225;
assign n_361 = ~n_226 & ~n_224;
assign n_362 = n_226 ^ n_227;
assign n_363 = n_237 ^ n_238;
assign n_364 = ~n_237 & ~n_239;
assign n_365 = n_239 ^ n_240;
assign n_366 = n_241 ^ x447;
assign n_367 = n_241 ^ n_242;
assign n_368 = n_245 ^ n_246;
assign n_369 = n_249 ^ n_250;
assign n_370 = n_251 ^ x453;
assign n_371 = n_251 ^ n_252;
assign n_372 = n_253 & n_255;
assign n_373 = n_257 ^ n_258;
assign n_374 = n_310 ^ n_311;
assign n_375 = n_312 ^ n_313;
assign n_376 = n_315 & n_317;
assign n_377 = n_318 ^ n_160;
assign n_378 = n_160 & n_318;
assign n_379 = ~n_2 & ~n_320;
assign n_380 = ~n_45 & ~n_321;
assign n_381 = ~n_40 & ~n_322;
assign n_382 = ~n_53 & ~n_324;
assign n_383 = ~n_48 & ~n_325;
assign n_384 = n_328 ^ x177;
assign n_385 = ~n_75 & ~n_330;
assign n_386 = ~n_329 & ~n_331;
assign n_387 = n_333 ^ x192;
assign n_388 = ~n_87 & ~n_334;
assign n_389 = n_336 & ~n_335;
assign n_390 = ~n_90 & ~n_337;
assign n_391 = ~n_92 & ~n_338;
assign n_392 = ~n_94 & ~n_339;
assign n_393 = ~n_96 & ~n_340;
assign n_394 = ~n_98 & ~n_341;
assign n_395 = ~n_100 & ~n_342;
assign n_396 = ~n_102 & ~n_343;
assign n_397 = ~n_104 & ~n_344;
assign n_398 = n_346 ^ x209;
assign n_399 = ~n_154 & ~n_347;
assign n_400 = n_348 ^ x253;
assign n_401 = ~n_164 & ~n_350;
assign n_402 = ~n_207 & ~n_352;
assign n_403 = ~n_351 & ~n_353;
assign n_404 = ~n_215 & ~n_355;
assign n_405 = ~n_210 & ~n_356;
assign n_406 = ~n_218 & ~n_358;
assign n_407 = ~n_220 & ~n_359;
assign n_408 = ~n_222 & ~n_360;
assign n_409 = n_362 ^ x436;
assign n_410 = ~n_235 & ~n_363;
assign n_411 = ~n_244 & n_366;
assign n_412 = ~n_367 & ~n_365;
assign n_413 = n_368 ^ x449;
assign n_414 = ~n_254 & ~n_370;
assign n_415 = ~n_369 & ~n_371;
assign n_416 = n_373 ^ x456;
assign n_417 = ~n_312 & ~n_374;
assign n_418 = n_375 ^ x509;
assign y127 = n_378;
assign n_419 = x129 ^ n_379;
assign n_420 = n_380 ^ x169;
assign n_421 = n_323 & n_381;
assign n_422 = n_382 ^ x173;
assign n_423 = n_326 & n_383;
assign n_424 = n_384 ^ x177;
assign n_425 = n_385 ^ x189;
assign n_426 = n_332 & n_386;
assign n_427 = n_387 ^ x192;
assign n_428 = n_388 ^ x197;
assign n_429 = n_398 ^ x209;
assign n_430 = n_349 & n_399;
assign n_431 = ~n_156 & ~n_400;
assign n_432 = x385 ^ n_401;
assign n_433 = n_402 ^ x425;
assign n_434 = n_354 & n_403;
assign n_435 = n_404 ^ x429;
assign n_436 = n_357 & n_405;
assign n_437 = n_409 ^ x436;
assign n_438 = n_411 ^ x319;
assign n_439 = n_412 & ~n_243;
assign n_440 = n_413 ^ x449;
assign n_441 = n_414 ^ x453;
assign n_442 = n_372 & n_415;
assign n_443 = n_416 ^ x456;
assign n_444 = n_376 & n_417;
assign n_445 = ~n_314 & ~n_418;
assign n_446 = n_419 ^ x130;
assign n_447 = n_420 ^ x170;
assign n_448 = n_422 ^ x174;
assign n_449 = n_425 ^ x190;
assign n_450 = n_428 ^ x198;
assign n_451 = n_431 ^ x253;
assign n_452 = n_432 ^ x386;
assign n_453 = n_433 ^ x426;
assign n_454 = n_435 ^ x430;
assign n_455 = ~n_245 & ~n_438;
assign n_456 = n_410 & n_439;
assign n_457 = ~n_364 & n_439;
assign n_458 = n_441 ^ x454;
assign n_459 = n_445 ^ x509;
assign n_460 = ~n_3 & n_446;
assign n_461 = ~n_47 & n_447;
assign n_462 = ~n_55 & n_448;
assign n_463 = ~n_77 & n_449;
assign n_464 = ~n_89 & n_450;
assign n_465 = n_451 ^ x254;
assign n_466 = ~n_165 & n_452;
assign n_467 = ~n_209 & n_453;
assign n_468 = ~n_217 & n_454;
assign n_469 = ~n_457 & n_455;
assign n_470 = ~n_256 & n_458;
assign n_471 = n_459 ^ x510;
assign n_472 = x130 ^ n_460;
assign n_473 = x170 ^ n_461;
assign n_474 = x174 ^ n_462;
assign n_475 = x190 ^ n_463;
assign n_476 = x198 ^ n_464;
assign n_477 = ~n_158 & n_465;
assign n_478 = x386 ^ n_466;
assign n_479 = x426 ^ n_467;
assign n_480 = x430 ^ n_468;
assign n_481 = x454 ^ n_470;
assign n_482 = ~n_316 & n_471;
assign n_483 = n_472 ^ x131;
assign n_484 = n_473 & ~n_49;
assign n_485 = n_474 & ~n_57;
assign n_486 = ~n_78 & n_475;
assign n_487 = n_476 & ~n_91;
assign n_488 = x254 ^ n_477;
assign n_489 = n_478 ^ x387;
assign n_490 = n_479 & ~n_211;
assign n_491 = n_480 & ~n_219;
assign n_492 = ~n_257 & n_481;
assign n_493 = x510 ^ n_482;
assign n_494 = ~n_4 & n_483;
assign n_495 = n_488 ^ x255;
assign n_496 = ~n_166 & ~n_489;
assign n_497 = n_493 ^ x511;
assign n_498 = x131 ^ n_494;
assign n_499 = n_495 ^ x255;
assign n_500 = x259 ^ n_496;
assign n_501 = n_497 ^ x511;
assign n_502 = n_498 ^ x132;
assign n_503 = n_500 ^ x388;
assign n_504 = ~n_5 & ~n_502;
assign n_505 = ~n_167 & n_503;
assign n_506 = x4 ^ n_504;
assign n_507 = x260 ^ n_505;
assign n_508 = n_506 ^ x133;
assign n_509 = n_507 ^ x389;
assign n_510 = ~n_6 & n_508;
assign n_511 = ~n_168 & ~n_509;
assign n_512 = x5 ^ n_510;
assign n_513 = x389 ^ n_511;
assign n_514 = n_512 ^ x134;
assign n_515 = n_513 ^ x390;
assign n_516 = ~n_7 & ~n_514;
assign n_517 = ~n_169 & n_515;
assign n_518 = x134 ^ n_516;
assign n_519 = x390 ^ n_517;
assign n_520 = n_518 ^ x135;
assign n_521 = n_519 ^ x391;
assign n_522 = ~n_8 & ~n_520;
assign n_523 = ~n_170 & n_521;
assign n_524 = x7 ^ n_522;
assign n_525 = x391 ^ n_523;
assign n_526 = n_524 ^ x136;
assign n_527 = n_525 ^ x392;
assign n_528 = ~n_9 & n_526;
assign n_529 = ~n_171 & n_527;
assign n_530 = x8 ^ n_528;
assign n_531 = x392 ^ n_529;
assign n_532 = n_530 ^ x137;
assign n_533 = n_531 ^ x393;
assign n_534 = ~n_10 & ~n_532;
assign n_535 = ~n_172 & n_533;
assign n_536 = x137 ^ n_534;
assign n_537 = x393 ^ n_535;
assign n_538 = n_536 ^ x138;
assign n_539 = n_537 ^ x394;
assign n_540 = ~n_11 & ~n_538;
assign n_541 = ~n_173 & ~n_539;
assign n_542 = x10 ^ n_540;
assign n_543 = x266 ^ n_541;
assign n_544 = n_542 ^ x139;
assign n_545 = n_543 ^ x395;
assign n_546 = ~n_12 & n_544;
assign n_547 = ~n_174 & n_545;
assign n_548 = x11 ^ n_546;
assign n_549 = x267 ^ n_547;
assign n_550 = n_548 ^ x140;
assign n_551 = n_549 ^ x396;
assign n_552 = ~n_13 & n_550;
assign n_553 = ~n_175 & n_551;
assign n_554 = x12 ^ n_552;
assign n_555 = x268 ^ n_553;
assign n_556 = n_554 ^ x141;
assign n_557 = n_555 ^ x397;
assign n_558 = ~n_14 & n_556;
assign n_559 = ~n_176 & n_557;
assign n_560 = x13 ^ n_558;
assign n_561 = x269 ^ n_559;
assign n_562 = n_560 ^ x142;
assign n_563 = n_561 ^ x398;
assign n_564 = ~n_15 & n_562;
assign n_565 = ~n_177 & n_563;
assign n_566 = x14 ^ n_564;
assign n_567 = x270 ^ n_565;
assign n_568 = n_566 ^ x143;
assign n_569 = n_567 ^ x399;
assign n_570 = ~n_16 & n_568;
assign n_571 = ~n_178 & n_569;
assign n_572 = x15 ^ n_570;
assign n_573 = x271 ^ n_571;
assign n_574 = n_572 ^ x144;
assign n_575 = n_573 ^ x400;
assign n_576 = ~n_17 & ~n_574;
assign n_577 = ~n_179 & n_575;
assign n_578 = x144 ^ n_576;
assign n_579 = x272 ^ n_577;
assign n_580 = n_578 ^ x145;
assign n_581 = n_579 ^ x401;
assign n_582 = ~n_18 & ~n_580;
assign n_583 = ~n_180 & n_581;
assign n_584 = x17 ^ n_582;
assign n_585 = x273 ^ n_583;
assign n_586 = n_584 ^ x146;
assign n_587 = n_585 ^ x402;
assign n_588 = ~n_19 & n_586;
assign n_589 = ~n_181 & ~n_587;
assign n_590 = x18 ^ n_588;
assign n_591 = x402 ^ n_589;
assign n_592 = n_590 ^ x147;
assign n_593 = n_591 ^ x403;
assign n_594 = ~n_20 & ~n_592;
assign n_595 = ~n_182 & ~n_593;
assign n_596 = x147 ^ n_594;
assign n_597 = x275 ^ n_595;
assign n_598 = n_596 ^ x148;
assign n_599 = n_597 ^ x404;
assign n_600 = ~n_21 & n_598;
assign n_601 = ~n_183 & n_599;
assign n_602 = x148 ^ n_600;
assign n_603 = x276 ^ n_601;
assign n_604 = n_602 ^ x149;
assign n_605 = n_603 ^ x405;
assign n_606 = ~n_22 & n_604;
assign n_607 = ~n_184 & ~n_605;
assign n_608 = x149 ^ n_606;
assign n_609 = x405 ^ n_607;
assign n_610 = n_608 ^ x150;
assign n_611 = n_609 ^ x406;
assign n_612 = ~n_23 & n_610;
assign n_613 = ~n_185 & n_611;
assign n_614 = x150 ^ n_612;
assign n_615 = x406 ^ n_613;
assign n_616 = n_614 ^ x151;
assign n_617 = n_615 ^ x407;
assign n_618 = ~n_24 & n_616;
assign n_619 = ~n_186 & n_617;
assign n_620 = x151 ^ n_618;
assign n_621 = x407 ^ n_619;
assign n_622 = n_620 ^ x152;
assign n_623 = n_621 ^ x408;
assign n_624 = ~n_25 & n_622;
assign n_625 = ~n_187 & n_623;
assign n_626 = x152 ^ n_624;
assign n_627 = x408 ^ n_625;
assign n_628 = n_626 ^ x153;
assign n_629 = n_627 ^ x409;
assign n_630 = ~n_26 & ~n_628;
assign n_631 = ~n_188 & ~n_629;
assign n_632 = x25 ^ n_630;
assign n_633 = x281 ^ n_631;
assign n_634 = n_632 ^ x154;
assign n_635 = n_633 ^ x410;
assign n_636 = ~n_27 & n_634;
assign n_637 = ~n_189 & n_635;
assign n_638 = x26 ^ n_636;
assign n_639 = x282 ^ n_637;
assign n_640 = n_638 ^ x155;
assign n_641 = n_639 ^ x411;
assign n_642 = ~n_28 & ~n_640;
assign n_643 = ~n_190 & ~n_641;
assign n_644 = x155 ^ n_642;
assign n_645 = x411 ^ n_643;
assign n_646 = n_644 ^ x156;
assign n_647 = n_645 ^ x412;
assign n_648 = ~n_29 & ~n_646;
assign n_649 = ~n_191 & n_647;
assign n_650 = x28 ^ n_648;
assign n_651 = x412 ^ n_649;
assign n_652 = n_650 ^ x157;
assign n_653 = n_651 ^ x413;
assign n_654 = ~n_30 & n_652;
assign n_655 = ~n_192 & ~n_653;
assign n_656 = x29 ^ n_654;
assign n_657 = x285 ^ n_655;
assign n_658 = n_656 ^ x158;
assign n_659 = n_657 ^ x414;
assign n_660 = ~n_31 & ~n_658;
assign n_661 = ~n_193 & n_659;
assign n_662 = x158 ^ n_660;
assign n_663 = x286 ^ n_661;
assign n_664 = n_662 ^ x159;
assign n_665 = n_663 ^ x415;
assign n_666 = ~n_32 & ~n_664;
assign n_667 = ~n_194 & ~n_665;
assign n_668 = x31 ^ n_666;
assign n_669 = x415 ^ n_667;
assign n_670 = n_668 ^ x160;
assign n_671 = n_669 ^ x416;
assign n_672 = ~n_33 & n_670;
assign n_673 = ~n_195 & n_671;
assign n_674 = x32 ^ n_672;
assign n_675 = x416 ^ n_673;
assign n_676 = n_674 ^ x161;
assign n_677 = n_675 ^ x417;
assign n_678 = ~n_34 & ~n_676;
assign n_679 = ~n_196 & n_677;
assign n_680 = x161 ^ n_678;
assign n_681 = x417 ^ n_679;
assign n_682 = n_680 ^ x162;
assign n_683 = n_681 ^ x418;
assign n_684 = ~n_35 & n_682;
assign n_685 = ~n_197 & ~n_683;
assign n_686 = x162 ^ n_684;
assign n_687 = x290 ^ n_685;
assign n_688 = n_686 ^ x163;
assign n_689 = n_687 ^ x419;
assign n_690 = ~n_36 & n_688;
assign n_691 = ~n_198 & n_689;
assign n_692 = x163 ^ n_690;
assign n_693 = x291 ^ n_691;
assign n_694 = n_692 ^ x164;
assign n_695 = n_693 ^ x420;
assign n_696 = ~n_37 & n_694;
assign n_697 = ~n_199 & n_695;
assign n_698 = x164 ^ n_696;
assign n_699 = x292 ^ n_697;
assign n_700 = n_698 ^ x165;
assign n_701 = n_699 ^ x421;
assign n_702 = ~n_38 & ~n_700;
assign n_703 = ~n_200 & n_701;
assign n_704 = x37 ^ n_702;
assign n_705 = x293 ^ n_703;
assign n_706 = n_704 ^ x166;
assign n_707 = n_705 ^ x422;
assign n_708 = ~n_39 & n_706;
assign n_709 = ~n_201 & ~n_707;
assign n_710 = x38 ^ n_708;
assign n_711 = x422 ^ n_709;
assign n_712 = ~n_710 & ~n_41;
assign n_713 = ~n_202 & n_711;
assign n_714 = ~n_712 & n_421;
assign n_715 = n_434 & ~n_713;
assign n_716 = ~n_714 & n_484;
assign n_717 = ~n_715 & n_490;
assign n_718 = ~n_716 & n_423;
assign n_719 = ~n_717 & n_436;
assign n_720 = ~n_718 & n_485;
assign n_721 = ~n_719 & n_491;
assign n_722 = n_327 & ~n_720;
assign n_723 = n_406 & ~n_721;
assign n_724 = x177 ^ n_722;
assign n_725 = n_407 & ~n_723;
assign n_726 = n_724 ^ x177;
assign n_727 = n_408 & ~n_725;
assign n_728 = ~n_424 & ~n_726;
assign n_729 = n_361 & ~n_727;
assign n_730 = x177 ^ n_728;
assign n_731 = x436 ^ n_729;
assign n_732 = ~n_60 & ~n_730;
assign n_733 = n_731 ^ x436;
assign n_734 = x49 ^ n_732;
assign n_735 = ~n_437 & ~n_733;
assign n_736 = n_734 ^ x178;
assign n_737 = x436 ^ n_735;
assign n_738 = ~n_61 & ~n_736;
assign n_739 = ~n_228 & n_737;
assign n_740 = x178 ^ n_738;
assign n_741 = x308 ^ n_739;
assign n_742 = n_740 ^ x179;
assign n_743 = n_741 ^ x437;
assign n_744 = ~n_62 & n_742;
assign n_745 = ~n_229 & ~n_743;
assign n_746 = x179 ^ n_744;
assign n_747 = x437 ^ n_745;
assign n_748 = n_746 ^ x180;
assign n_749 = n_747 ^ x438;
assign n_750 = ~n_63 & n_748;
assign n_751 = ~n_230 & n_749;
assign n_752 = x180 ^ n_750;
assign n_753 = x438 ^ n_751;
assign n_754 = n_752 ^ x181;
assign n_755 = n_753 ^ x439;
assign n_756 = ~n_64 & n_754;
assign n_757 = ~n_231 & n_755;
assign n_758 = x181 ^ n_756;
assign n_759 = x439 ^ n_757;
assign n_760 = n_758 ^ x182;
assign n_761 = n_759 ^ x440;
assign n_762 = ~n_65 & n_760;
assign n_763 = ~n_232 & n_761;
assign n_764 = x182 ^ n_762;
assign n_765 = x440 ^ n_763;
assign n_766 = n_764 ^ x183;
assign n_767 = n_765 ^ x441;
assign n_768 = ~n_66 & ~n_766;
assign n_769 = ~n_233 & ~n_767;
assign n_770 = x55 ^ n_768;
assign n_771 = x313 ^ n_769;
assign n_772 = n_770 ^ x184;
assign n_773 = n_771 ^ x442;
assign n_774 = ~n_67 & n_772;
assign n_775 = ~n_234 & n_773;
assign n_776 = x56 ^ n_774;
assign n_777 = x314 ^ n_775;
assign n_778 = n_776 ^ x185;
assign n_779 = ~n_777 & ~n_236;
assign n_780 = ~n_68 & ~n_778;
assign n_781 = ~n_779 & n_456;
assign n_782 = x185 ^ n_780;
assign n_783 = ~n_781 & n_469;
assign n_784 = n_782 ^ x186;
assign n_785 = x449 ^ n_783;
assign n_786 = ~n_69 & n_784;
assign n_787 = n_785 ^ x449;
assign n_788 = x186 ^ n_786;
assign n_789 = ~n_440 & ~n_787;
assign n_790 = ~n_70 & n_788;
assign n_791 = x449 ^ n_789;
assign n_792 = n_426 & ~n_790;
assign n_793 = ~n_247 & n_791;
assign n_794 = ~n_792 & n_486;
assign n_795 = x321 ^ n_793;
assign n_796 = x192 ^ n_794;
assign n_797 = n_795 ^ x450;
assign n_798 = n_796 ^ x192;
assign n_799 = ~n_248 & ~n_797;
assign n_800 = ~n_427 & ~n_798;
assign n_801 = x450 ^ n_799;
assign n_802 = x192 ^ n_800;
assign n_803 = ~n_249 & n_801;
assign n_804 = ~n_80 & n_802;
assign n_805 = n_442 & ~n_803;
assign n_806 = x64 ^ n_804;
assign n_807 = ~n_805 & n_492;
assign n_808 = n_806 ^ x193;
assign n_809 = x456 ^ n_807;
assign n_810 = ~n_81 & ~n_808;
assign n_811 = n_809 ^ x456;
assign n_812 = x193 ^ n_810;
assign n_813 = ~n_443 & ~n_811;
assign n_814 = n_812 ^ x194;
assign n_815 = x456 ^ n_813;
assign n_816 = ~n_82 & ~n_814;
assign n_817 = ~n_259 & n_815;
assign n_818 = x66 ^ n_816;
assign n_819 = x328 ^ n_817;
assign n_820 = n_818 ^ x195;
assign n_821 = n_819 ^ x457;
assign n_822 = ~n_83 & n_820;
assign n_823 = ~n_260 & ~n_821;
assign n_824 = x67 ^ n_822;
assign n_825 = x457 ^ n_823;
assign n_826 = n_824 & n_389;
assign n_827 = n_825 ^ x458;
assign n_828 = ~n_826 & n_487;
assign n_829 = ~n_261 & ~n_827;
assign n_830 = n_390 & ~n_828;
assign n_831 = x330 ^ n_829;
assign n_832 = n_391 & ~n_830;
assign n_833 = n_831 ^ x459;
assign n_834 = n_392 & ~n_832;
assign n_835 = ~n_262 & n_833;
assign n_836 = n_393 & ~n_834;
assign n_837 = x331 ^ n_835;
assign n_838 = n_394 & ~n_836;
assign n_839 = n_837 ^ x460;
assign n_840 = n_395 & ~n_838;
assign n_841 = ~n_263 & ~n_839;
assign n_842 = n_396 & ~n_840;
assign n_843 = x460 ^ n_841;
assign n_844 = n_397 & ~n_842;
assign n_845 = n_843 ^ x461;
assign n_846 = n_345 & ~n_844;
assign n_847 = ~n_264 & ~n_845;
assign n_848 = x209 ^ n_846;
assign n_849 = x333 ^ n_847;
assign n_850 = n_848 ^ x209;
assign n_851 = n_849 ^ x462;
assign n_852 = ~n_429 & ~n_850;
assign n_853 = ~n_265 & n_851;
assign n_854 = x209 ^ n_852;
assign n_855 = x334 ^ n_853;
assign n_856 = ~n_110 & ~n_854;
assign n_857 = n_855 ^ x463;
assign n_858 = x81 ^ n_856;
assign n_859 = ~n_266 & ~n_857;
assign n_860 = n_858 ^ x210;
assign n_861 = x463 ^ n_859;
assign n_862 = ~n_111 & ~n_860;
assign n_863 = n_861 ^ x464;
assign n_864 = x210 ^ n_862;
assign n_865 = ~n_267 & n_863;
assign n_866 = n_864 ^ x211;
assign n_867 = x464 ^ n_865;
assign n_868 = ~n_112 & n_866;
assign n_869 = n_867 ^ x465;
assign n_870 = x211 ^ n_868;
assign n_871 = ~n_268 & ~n_869;
assign n_872 = n_870 ^ x212;
assign n_873 = x337 ^ n_871;
assign n_874 = ~n_113 & n_872;
assign n_875 = n_873 ^ x466;
assign n_876 = x212 ^ n_874;
assign n_877 = ~n_269 & n_875;
assign n_878 = n_876 ^ x213;
assign n_879 = x338 ^ n_877;
assign n_880 = ~n_114 & n_878;
assign n_881 = n_879 ^ x467;
assign n_882 = x213 ^ n_880;
assign n_883 = ~n_270 & ~n_881;
assign n_884 = n_882 ^ x214;
assign n_885 = x467 ^ n_883;
assign n_886 = ~n_115 & n_884;
assign n_887 = n_885 ^ x468;
assign n_888 = x214 ^ n_886;
assign n_889 = ~n_271 & n_887;
assign n_890 = n_888 ^ x215;
assign n_891 = x468 ^ n_889;
assign n_892 = ~n_116 & n_890;
assign n_893 = n_891 ^ x469;
assign n_894 = x215 ^ n_892;
assign n_895 = ~n_272 & n_893;
assign n_896 = n_894 ^ x216;
assign n_897 = x469 ^ n_895;
assign n_898 = ~n_117 & n_896;
assign n_899 = n_897 ^ x470;
assign n_900 = x216 ^ n_898;
assign n_901 = ~n_273 & ~n_899;
assign n_902 = n_900 ^ x217;
assign n_903 = x342 ^ n_901;
assign n_904 = ~n_118 & ~n_902;
assign n_905 = n_903 ^ x471;
assign n_906 = x89 ^ n_904;
assign n_907 = ~n_274 & n_905;
assign n_908 = n_906 ^ x218;
assign n_909 = x343 ^ n_907;
assign n_910 = ~n_119 & n_908;
assign n_911 = n_909 ^ x472;
assign n_912 = x90 ^ n_910;
assign n_913 = ~n_275 & n_911;
assign n_914 = n_912 ^ x219;
assign n_915 = x344 ^ n_913;
assign n_916 = ~n_120 & n_914;
assign n_917 = n_915 ^ x473;
assign n_918 = x91 ^ n_916;
assign n_919 = ~n_276 & n_917;
assign n_920 = n_918 ^ x220;
assign n_921 = x345 ^ n_919;
assign n_922 = ~n_121 & n_920;
assign n_923 = n_921 ^ x474;
assign n_924 = x92 ^ n_922;
assign n_925 = ~n_277 & ~n_923;
assign n_926 = n_924 ^ x221;
assign n_927 = x474 ^ n_925;
assign n_928 = ~n_122 & n_926;
assign n_929 = n_927 ^ x475;
assign n_930 = x93 ^ n_928;
assign n_931 = ~n_278 & ~n_929;
assign n_932 = n_930 ^ x222;
assign n_933 = x347 ^ n_931;
assign n_934 = ~n_123 & n_932;
assign n_935 = n_933 ^ x476;
assign n_936 = x94 ^ n_934;
assign n_937 = ~n_279 & n_935;
assign n_938 = n_936 ^ x223;
assign n_939 = x348 ^ n_937;
assign n_940 = ~n_124 & ~n_938;
assign n_941 = n_939 ^ x477;
assign n_942 = x223 ^ n_940;
assign n_943 = ~n_280 & ~n_941;
assign n_944 = n_942 ^ x224;
assign n_945 = x477 ^ n_943;
assign n_946 = ~n_125 & ~n_944;
assign n_947 = n_945 ^ x478;
assign n_948 = x96 ^ n_946;
assign n_949 = ~n_281 & n_947;
assign n_950 = n_948 ^ x225;
assign n_951 = x478 ^ n_949;
assign n_952 = ~n_126 & n_950;
assign n_953 = n_951 ^ x479;
assign n_954 = x97 ^ n_952;
assign n_955 = ~n_282 & n_953;
assign n_956 = n_954 ^ x226;
assign n_957 = x479 ^ n_955;
assign n_958 = ~n_127 & ~n_956;
assign n_959 = n_957 ^ x480;
assign n_960 = x226 ^ n_958;
assign n_961 = ~n_283 & n_959;
assign n_962 = n_960 ^ x227;
assign n_963 = x480 ^ n_961;
assign n_964 = ~n_128 & n_962;
assign n_965 = n_963 ^ x481;
assign n_966 = x227 ^ n_964;
assign n_967 = ~n_284 & ~n_965;
assign n_968 = n_966 ^ x228;
assign n_969 = x353 ^ n_967;
assign n_970 = ~n_129 & ~n_968;
assign n_971 = n_969 ^ x482;
assign n_972 = x100 ^ n_970;
assign n_973 = ~n_285 & n_971;
assign n_974 = n_972 ^ x229;
assign n_975 = x354 ^ n_973;
assign n_976 = ~n_130 & n_974;
assign n_977 = n_975 ^ x483;
assign n_978 = x101 ^ n_976;
assign n_979 = ~n_286 & ~n_977;
assign n_980 = n_978 ^ x230;
assign n_981 = x483 ^ n_979;
assign n_982 = ~n_131 & ~n_980;
assign n_983 = n_981 ^ x484;
assign n_984 = x230 ^ n_982;
assign n_985 = ~n_287 & n_983;
assign n_986 = n_984 ^ x231;
assign n_987 = x484 ^ n_985;
assign n_988 = ~n_132 & n_986;
assign n_989 = n_987 ^ x485;
assign n_990 = x231 ^ n_988;
assign n_991 = ~n_288 & n_989;
assign n_992 = n_990 ^ x232;
assign n_993 = x485 ^ n_991;
assign n_994 = ~n_133 & ~n_992;
assign n_995 = n_993 ^ x486;
assign n_996 = x104 ^ n_994;
assign n_997 = ~n_289 & ~n_995;
assign n_998 = n_996 ^ x233;
assign n_999 = x358 ^ n_997;
assign n_1000 = ~n_134 & n_998;
assign n_1001 = n_999 ^ x487;
assign n_1002 = x105 ^ n_1000;
assign n_1003 = ~n_290 & n_1001;
assign n_1004 = n_1002 ^ x234;
assign n_1005 = x359 ^ n_1003;
assign n_1006 = ~n_135 & ~n_1004;
assign n_1007 = n_1005 ^ x488;
assign n_1008 = x234 ^ n_1006;
assign n_1009 = ~n_291 & n_1007;
assign n_1010 = n_1008 ^ x235;
assign n_1011 = x360 ^ n_1009;
assign n_1012 = ~n_136 & n_1010;
assign n_1013 = n_1011 ^ x489;
assign n_1014 = x235 ^ n_1012;
assign n_1015 = ~n_292 & n_1013;
assign n_1016 = n_1014 ^ x236;
assign n_1017 = x361 ^ n_1015;
assign n_1018 = ~n_137 & ~n_1016;
assign n_1019 = n_1017 ^ x490;
assign n_1020 = x108 ^ n_1018;
assign n_1021 = ~n_293 & n_1019;
assign n_1022 = n_1020 ^ x237;
assign n_1023 = x362 ^ n_1021;
assign n_1024 = ~n_138 & n_1022;
assign n_1025 = n_1023 ^ x491;
assign n_1026 = x109 ^ n_1024;
assign n_1027 = ~n_294 & n_1025;
assign n_1028 = n_1026 ^ x238;
assign n_1029 = x363 ^ n_1027;
assign n_1030 = ~n_139 & ~n_1028;
assign n_1031 = n_1029 ^ x492;
assign n_1032 = x238 ^ n_1030;
assign n_1033 = ~n_295 & ~n_1031;
assign n_1034 = n_1032 ^ x239;
assign n_1035 = x492 ^ n_1033;
assign n_1036 = ~n_140 & n_1034;
assign n_1037 = n_1035 ^ x493;
assign n_1038 = x239 ^ n_1036;
assign n_1039 = ~n_296 & ~n_1037;
assign n_1040 = n_1038 ^ x240;
assign n_1041 = x365 ^ n_1039;
assign n_1042 = ~n_141 & ~n_1040;
assign n_1043 = n_1041 ^ x494;
assign n_1044 = x112 ^ n_1042;
assign n_1045 = ~n_297 & n_1043;
assign n_1046 = n_1044 ^ x241;
assign n_1047 = x366 ^ n_1045;
assign n_1048 = ~n_142 & n_1046;
assign n_1049 = n_1047 ^ x495;
assign n_1050 = x113 ^ n_1048;
assign n_1051 = ~n_298 & ~n_1049;
assign n_1052 = n_1050 ^ x242;
assign n_1053 = x495 ^ n_1051;
assign n_1054 = ~n_143 & ~n_1052;
assign n_1055 = n_1053 ^ x496;
assign n_1056 = x242 ^ n_1054;
assign n_1057 = ~n_299 & n_1055;
assign n_1058 = n_1056 ^ x243;
assign n_1059 = x496 ^ n_1057;
assign n_1060 = ~n_144 & ~n_1058;
assign n_1061 = n_1059 ^ x497;
assign n_1062 = x115 ^ n_1060;
assign n_1063 = ~n_300 & n_1061;
assign n_1064 = n_1062 ^ x244;
assign n_1065 = x497 ^ n_1063;
assign n_1066 = ~n_145 & n_1064;
assign n_1067 = n_1065 ^ x498;
assign n_1068 = x116 ^ n_1066;
assign n_1069 = ~n_301 & n_1067;
assign n_1070 = n_1068 ^ x245;
assign n_1071 = x498 ^ n_1069;
assign n_1072 = ~n_146 & ~n_1070;
assign n_1073 = n_1071 ^ x499;
assign n_1074 = x245 ^ n_1072;
assign n_1075 = ~n_302 & ~n_1073;
assign n_1076 = n_1074 ^ x246;
assign n_1077 = x371 ^ n_1075;
assign n_1078 = ~n_147 & ~n_1076;
assign n_1079 = n_1077 ^ x500;
assign n_1080 = x118 ^ n_1078;
assign n_1081 = ~n_303 & n_1079;
assign n_1082 = n_1080 ^ x247;
assign n_1083 = x372 ^ n_1081;
assign n_1084 = ~n_148 & n_1082;
assign n_1085 = n_1083 ^ x501;
assign n_1086 = x119 ^ n_1084;
assign n_1087 = ~n_304 & ~n_1085;
assign n_1088 = n_1086 ^ x248;
assign n_1089 = x501 ^ n_1087;
assign n_1090 = ~n_149 & n_1088;
assign n_1091 = n_1089 ^ x502;
assign n_1092 = x120 ^ n_1090;
assign n_1093 = ~n_305 & ~n_1091;
assign n_1094 = n_1092 ^ x249;
assign n_1095 = x374 ^ n_1093;
assign n_1096 = ~n_150 & n_1094;
assign n_1097 = n_1095 ^ x503;
assign n_1098 = x121 ^ n_1096;
assign n_1099 = ~n_306 & n_1097;
assign n_1100 = n_1098 ^ x250;
assign n_1101 = x375 ^ n_1099;
assign n_1102 = ~n_151 & ~n_1100;
assign n_1103 = n_1101 ^ x504;
assign n_1104 = x250 ^ n_1102;
assign n_1105 = ~n_307 & ~n_1103;
assign n_1106 = ~n_152 & n_1104;
assign n_1107 = x504 ^ n_1105;
assign n_1108 = n_430 & ~n_1106;
assign n_1109 = n_1107 ^ x505;
assign n_1110 = x255 ^ n_1108;
assign n_1111 = ~n_308 & n_1109;
assign n_1112 = n_1110 ^ x255;
assign n_1113 = x505 ^ n_1111;
assign n_1114 = n_499 & ~n_1112;
assign n_1115 = n_1113 ^ x506;
assign n_1116 = x255 ^ n_1114;
assign n_1117 = ~n_309 & n_1115;
assign n_1118 = ~n_161 & n_1116;
assign n_1119 = x506 ^ n_1117;
assign n_1120 = x127 ^ n_1118;
assign n_1121 = ~n_310 & n_1119;
assign n_1122 = n_158 & n_1120;
assign n_1123 = n_156 & n_1120;
assign n_1124 = n_155 & n_1120;
assign n_1125 = n_153 & n_1120;
assign n_1126 = n_151 & n_1120;
assign n_1127 = n_150 & n_1120;
assign n_1128 = n_149 & n_1120;
assign n_1129 = n_148 & n_1120;
assign n_1130 = n_147 & n_1120;
assign n_1131 = n_146 & n_1120;
assign n_1132 = n_145 & n_1120;
assign n_1133 = n_144 & n_1120;
assign n_1134 = n_143 & n_1120;
assign n_1135 = n_142 & n_1120;
assign n_1136 = n_141 & n_1120;
assign n_1137 = n_140 & n_1120;
assign n_1138 = n_139 & n_1120;
assign n_1139 = n_138 & n_1120;
assign n_1140 = n_137 & n_1120;
assign n_1141 = n_136 & n_1120;
assign n_1142 = n_135 & n_1120;
assign n_1143 = n_134 & n_1120;
assign n_1144 = n_133 & n_1120;
assign n_1145 = n_132 & n_1120;
assign n_1146 = n_131 & n_1120;
assign n_1147 = n_130 & n_1120;
assign n_1148 = n_129 & n_1120;
assign n_1149 = n_128 & n_1120;
assign n_1150 = n_127 & n_1120;
assign n_1151 = n_126 & n_1120;
assign n_1152 = n_125 & n_1120;
assign n_1153 = n_124 & n_1120;
assign n_1154 = n_123 & n_1120;
assign n_1155 = n_122 & n_1120;
assign n_1156 = n_121 & n_1120;
assign n_1157 = n_120 & n_1120;
assign n_1158 = n_119 & n_1120;
assign n_1159 = n_118 & n_1120;
assign n_1160 = n_117 & n_1120;
assign n_1161 = n_116 & n_1120;
assign n_1162 = n_115 & n_1120;
assign n_1163 = n_114 & n_1120;
assign n_1164 = n_113 & n_1120;
assign n_1165 = n_112 & n_1120;
assign n_1166 = n_111 & n_1120;
assign n_1167 = n_110 & n_1120;
assign n_1168 = n_109 & n_1120;
assign n_1169 = n_107 & n_1120;
assign n_1170 = n_105 & n_1120;
assign n_1171 = n_103 & n_1120;
assign n_1172 = n_101 & n_1120;
assign n_1173 = n_99 & n_1120;
assign n_1174 = n_97 & n_1120;
assign n_1175 = n_95 & n_1120;
assign n_1176 = n_93 & n_1120;
assign n_1177 = n_91 & n_1120;
assign n_1178 = n_89 & n_1120;
assign n_1179 = n_87 & n_1120;
assign n_1180 = n_85 & n_1120;
assign n_1181 = n_83 & n_1120;
assign n_1182 = n_82 & n_1120;
assign n_1183 = n_81 & n_1120;
assign n_1184 = n_80 & n_1120;
assign n_1185 = n_79 & n_1120;
assign n_1186 = n_77 & n_1120;
assign n_1187 = n_75 & n_1120;
assign n_1188 = n_73 & n_1120;
assign n_1189 = n_71 & n_1120;
assign n_1190 = n_69 & n_1120;
assign n_1191 = n_68 & n_1120;
assign n_1192 = n_67 & n_1120;
assign n_1193 = n_66 & n_1120;
assign n_1194 = n_65 & n_1120;
assign n_1195 = n_64 & n_1120;
assign n_1196 = n_63 & n_1120;
assign n_1197 = n_62 & n_1120;
assign n_1198 = n_61 & n_1120;
assign n_1199 = n_60 & n_1120;
assign n_1200 = n_59 & n_1120;
assign n_1201 = n_57 & n_1120;
assign n_1202 = n_55 & n_1120;
assign n_1203 = n_53 & n_1120;
assign n_1204 = n_51 & n_1120;
assign n_1205 = n_49 & n_1120;
assign n_1206 = n_47 & n_1120;
assign n_1207 = n_45 & n_1120;
assign n_1208 = n_43 & n_1120;
assign n_1209 = n_41 & n_1120;
assign n_1210 = n_39 & n_1120;
assign n_1211 = n_38 & n_1120;
assign n_1212 = n_37 & n_1120;
assign n_1213 = n_36 & n_1120;
assign n_1214 = n_35 & n_1120;
assign n_1215 = n_34 & n_1120;
assign n_1216 = n_33 & n_1120;
assign n_1217 = n_32 & n_1120;
assign n_1218 = n_31 & n_1120;
assign n_1219 = n_30 & n_1120;
assign n_1220 = n_29 & n_1120;
assign n_1221 = n_28 & n_1120;
assign n_1222 = n_27 & n_1120;
assign n_1223 = n_26 & n_1120;
assign n_1224 = n_25 & n_1120;
assign n_1225 = n_24 & n_1120;
assign n_1226 = n_23 & n_1120;
assign n_1227 = n_22 & n_1120;
assign n_1228 = n_21 & n_1120;
assign n_1229 = n_20 & n_1120;
assign n_1230 = n_19 & n_1120;
assign n_1231 = n_18 & n_1120;
assign n_1232 = n_17 & n_1120;
assign n_1233 = n_16 & n_1120;
assign n_1234 = n_15 & n_1120;
assign n_1235 = n_14 & n_1120;
assign n_1236 = n_13 & n_1120;
assign n_1237 = n_12 & n_1120;
assign n_1238 = n_11 & n_1120;
assign n_1239 = n_10 & n_1120;
assign n_1240 = n_9 & n_1120;
assign n_1241 = n_8 & n_1120;
assign n_1242 = n_7 & n_1120;
assign n_1243 = n_6 & n_1120;
assign n_1244 = n_5 & n_1120;
assign n_1245 = n_4 & n_1120;
assign n_1246 = n_3 & n_1120;
assign n_1247 = n_2 & n_1120;
assign n_1248 = n_1120 & n_1;
assign n_1249 = n_444 & ~n_1121;
assign n_1250 = n_1122 ^ x126;
assign n_1251 = n_1123 ^ x125;
assign n_1252 = n_1124 ^ x124;
assign n_1253 = n_1125 ^ x123;
assign n_1254 = n_1126 ^ x122;
assign n_1255 = n_1127 ^ x121;
assign n_1256 = n_1128 ^ x120;
assign n_1257 = n_1129 ^ x119;
assign n_1258 = n_1130 ^ x118;
assign n_1259 = n_1131 ^ x117;
assign n_1260 = n_1132 ^ x116;
assign n_1261 = n_1133 ^ x115;
assign n_1262 = n_1134 ^ x114;
assign n_1263 = n_1135 ^ x113;
assign n_1264 = n_1136 ^ x112;
assign n_1265 = n_1137 ^ x111;
assign n_1266 = n_1138 ^ x110;
assign n_1267 = n_1139 ^ x109;
assign n_1268 = n_1140 ^ x108;
assign n_1269 = n_1141 ^ x107;
assign n_1270 = n_1142 ^ x106;
assign n_1271 = n_1143 ^ x105;
assign n_1272 = n_1144 ^ x104;
assign n_1273 = n_1145 ^ x103;
assign n_1274 = n_1146 ^ x102;
assign n_1275 = n_1147 ^ x101;
assign n_1276 = n_1148 ^ x100;
assign n_1277 = n_1149 ^ x99;
assign n_1278 = n_1150 ^ x98;
assign n_1279 = n_1151 ^ x97;
assign n_1280 = n_1152 ^ x96;
assign n_1281 = n_1153 ^ x95;
assign n_1282 = n_1154 ^ x94;
assign n_1283 = n_1155 ^ x93;
assign n_1284 = n_1156 ^ x92;
assign n_1285 = n_1157 ^ x91;
assign n_1286 = n_1158 ^ x90;
assign n_1287 = n_1159 ^ x89;
assign n_1288 = n_1160 ^ x88;
assign n_1289 = n_1161 ^ x87;
assign n_1290 = n_1162 ^ x86;
assign n_1291 = n_1163 ^ x85;
assign n_1292 = n_1164 ^ x84;
assign n_1293 = n_1165 ^ x83;
assign n_1294 = n_1166 ^ x82;
assign n_1295 = n_1167 ^ x81;
assign n_1296 = n_1168 ^ x80;
assign n_1297 = n_1169 ^ x79;
assign n_1298 = n_1170 ^ x78;
assign n_1299 = n_1171 ^ x77;
assign n_1300 = n_1172 ^ x76;
assign n_1301 = n_1173 ^ x75;
assign n_1302 = n_1174 ^ x74;
assign n_1303 = n_1175 ^ x73;
assign n_1304 = n_1176 ^ x72;
assign n_1305 = n_1177 ^ x71;
assign n_1306 = n_1178 ^ x70;
assign n_1307 = n_1179 ^ x69;
assign n_1308 = n_1180 ^ x68;
assign n_1309 = n_1181 ^ x67;
assign n_1310 = n_1182 ^ x66;
assign n_1311 = n_1183 ^ x65;
assign n_1312 = n_1184 ^ x64;
assign n_1313 = n_1185 ^ x63;
assign n_1314 = n_1186 ^ x62;
assign n_1315 = n_1187 ^ x61;
assign n_1316 = n_1188 ^ x60;
assign n_1317 = n_1189 ^ x59;
assign n_1318 = n_1190 ^ x58;
assign n_1319 = n_1191 ^ x57;
assign n_1320 = n_1192 ^ x56;
assign n_1321 = n_1193 ^ x55;
assign n_1322 = n_1194 ^ x54;
assign n_1323 = n_1195 ^ x53;
assign n_1324 = n_1196 ^ x52;
assign n_1325 = n_1197 ^ x51;
assign n_1326 = n_1198 ^ x50;
assign n_1327 = n_1199 ^ x49;
assign n_1328 = n_1200 ^ x48;
assign n_1329 = n_1201 ^ x47;
assign n_1330 = n_1202 ^ x46;
assign n_1331 = n_1203 ^ x45;
assign n_1332 = n_1204 ^ x44;
assign n_1333 = n_1205 ^ x43;
assign n_1334 = n_1206 ^ x42;
assign n_1335 = n_1207 ^ x41;
assign n_1336 = n_1208 ^ x40;
assign n_1337 = n_1209 ^ x39;
assign n_1338 = n_1210 ^ x38;
assign n_1339 = n_1211 ^ x37;
assign n_1340 = n_1212 ^ x36;
assign n_1341 = n_1213 ^ x35;
assign n_1342 = n_1214 ^ x34;
assign n_1343 = n_1215 ^ x33;
assign n_1344 = n_1216 ^ x32;
assign n_1345 = n_1217 ^ x31;
assign n_1346 = n_1218 ^ x30;
assign n_1347 = n_1219 ^ x29;
assign n_1348 = n_1220 ^ x28;
assign n_1349 = n_1221 ^ x27;
assign n_1350 = n_1222 ^ x26;
assign n_1351 = n_1223 ^ x25;
assign n_1352 = n_1224 ^ x24;
assign n_1353 = n_1225 ^ x23;
assign n_1354 = n_1226 ^ x22;
assign n_1355 = n_1227 ^ x21;
assign n_1356 = n_1228 ^ x20;
assign n_1357 = n_1229 ^ x19;
assign n_1358 = n_1230 ^ x18;
assign n_1359 = n_1231 ^ x17;
assign n_1360 = n_1232 ^ x16;
assign n_1361 = n_1233 ^ x15;
assign n_1362 = n_1234 ^ x14;
assign n_1363 = n_1235 ^ x13;
assign n_1364 = n_1236 ^ x12;
assign n_1365 = n_1237 ^ x11;
assign n_1366 = n_1238 ^ x10;
assign n_1367 = n_1239 ^ x9;
assign n_1368 = n_1240 ^ x8;
assign n_1369 = n_1241 ^ x7;
assign n_1370 = n_1242 ^ x6;
assign n_1371 = n_1243 ^ x5;
assign n_1372 = n_1244 ^ x4;
assign n_1373 = n_1245 ^ x3;
assign n_1374 = n_1246 ^ x2;
assign n_1375 = n_1247 ^ x1;
assign n_1376 = n_1248 ^ x0;
assign n_1377 = x511 ^ n_1249;
assign n_1378 = n_1377 ^ x511;
assign n_1379 = n_501 & ~n_1378;
assign n_1380 = x511 ^ n_1379;
assign n_1381 = ~n_319 & n_1380;
assign n_1382 = x383 ^ n_1381;
assign n_1383 = n_316 & n_1382;
assign n_1384 = n_314 & n_1382;
assign n_1385 = n_313 & n_1382;
assign n_1386 = n_311 & n_1382;
assign n_1387 = n_309 & n_1382;
assign n_1388 = n_308 & n_1382;
assign n_1389 = n_307 & n_1382;
assign n_1390 = n_306 & n_1382;
assign n_1391 = n_305 & n_1382;
assign n_1392 = n_304 & n_1382;
assign n_1393 = n_303 & n_1382;
assign n_1394 = n_302 & n_1382;
assign n_1395 = n_301 & n_1382;
assign n_1396 = n_300 & n_1382;
assign n_1397 = n_299 & n_1382;
assign n_1398 = n_298 & n_1382;
assign n_1399 = n_297 & n_1382;
assign n_1400 = n_296 & n_1382;
assign n_1401 = n_295 & n_1382;
assign n_1402 = n_294 & n_1382;
assign n_1403 = n_293 & n_1382;
assign n_1404 = n_292 & n_1382;
assign n_1405 = n_291 & n_1382;
assign n_1406 = n_290 & n_1382;
assign n_1407 = n_289 & n_1382;
assign n_1408 = n_288 & n_1382;
assign n_1409 = n_287 & n_1382;
assign n_1410 = n_286 & n_1382;
assign n_1411 = n_285 & n_1382;
assign n_1412 = n_284 & n_1382;
assign n_1413 = n_283 & n_1382;
assign n_1414 = n_282 & n_1382;
assign n_1415 = n_281 & n_1382;
assign n_1416 = n_280 & n_1382;
assign n_1417 = n_279 & n_1382;
assign n_1418 = n_278 & n_1382;
assign n_1419 = n_277 & n_1382;
assign n_1420 = n_276 & n_1382;
assign n_1421 = n_275 & n_1382;
assign n_1422 = n_274 & n_1382;
assign n_1423 = n_273 & n_1382;
assign n_1424 = n_272 & n_1382;
assign n_1425 = n_271 & n_1382;
assign n_1426 = n_270 & n_1382;
assign n_1427 = n_269 & n_1382;
assign n_1428 = n_268 & n_1382;
assign n_1429 = n_267 & n_1382;
assign n_1430 = n_266 & n_1382;
assign n_1431 = n_265 & n_1382;
assign n_1432 = n_264 & n_1382;
assign n_1433 = n_263 & n_1382;
assign n_1434 = n_262 & n_1382;
assign n_1435 = n_261 & n_1382;
assign n_1436 = n_260 & n_1382;
assign n_1437 = n_259 & n_1382;
assign n_1438 = n_258 & n_1382;
assign n_1439 = n_256 & n_1382;
assign n_1440 = n_254 & n_1382;
assign n_1441 = n_252 & n_1382;
assign n_1442 = n_250 & n_1382;
assign n_1443 = n_248 & n_1382;
assign n_1444 = n_247 & n_1382;
assign n_1445 = n_246 & n_1382;
assign n_1446 = n_244 & n_1382;
assign n_1447 = n_242 & n_1382;
assign n_1448 = n_240 & n_1382;
assign n_1449 = n_238 & n_1382;
assign n_1450 = n_236 & n_1382;
assign n_1451 = n_234 & n_1382;
assign n_1452 = n_233 & n_1382;
assign n_1453 = n_232 & n_1382;
assign n_1454 = n_231 & n_1382;
assign n_1455 = n_230 & n_1382;
assign n_1456 = n_229 & n_1382;
assign n_1457 = n_228 & n_1382;
assign n_1458 = n_227 & n_1382;
assign n_1459 = n_225 & n_1382;
assign n_1460 = n_223 & n_1382;
assign n_1461 = n_221 & n_1382;
assign n_1462 = n_219 & n_1382;
assign n_1463 = n_217 & n_1382;
assign n_1464 = n_215 & n_1382;
assign n_1465 = n_213 & n_1382;
assign n_1466 = n_211 & n_1382;
assign n_1467 = n_209 & n_1382;
assign n_1468 = n_207 & n_1382;
assign n_1469 = n_205 & n_1382;
assign n_1470 = n_203 & n_1382;
assign n_1471 = n_201 & n_1382;
assign n_1472 = n_200 & n_1382;
assign n_1473 = n_199 & n_1382;
assign n_1474 = n_198 & n_1382;
assign n_1475 = n_197 & n_1382;
assign n_1476 = n_196 & n_1382;
assign n_1477 = n_195 & n_1382;
assign n_1478 = n_194 & n_1382;
assign n_1479 = n_193 & n_1382;
assign n_1480 = n_192 & n_1382;
assign n_1481 = n_191 & n_1382;
assign n_1482 = n_190 & n_1382;
assign n_1483 = n_189 & n_1382;
assign n_1484 = n_188 & n_1382;
assign n_1485 = n_187 & n_1382;
assign n_1486 = n_186 & n_1382;
assign n_1487 = n_185 & n_1382;
assign n_1488 = n_184 & n_1382;
assign n_1489 = n_183 & n_1382;
assign n_1490 = n_182 & n_1382;
assign n_1491 = n_181 & n_1382;
assign n_1492 = n_180 & n_1382;
assign n_1493 = n_179 & n_1382;
assign n_1494 = n_178 & n_1382;
assign n_1495 = n_177 & n_1382;
assign n_1496 = n_176 & n_1382;
assign n_1497 = n_175 & n_1382;
assign n_1498 = n_174 & n_1382;
assign n_1499 = n_173 & n_1382;
assign n_1500 = n_172 & n_1382;
assign n_1501 = n_171 & n_1382;
assign n_1502 = n_170 & n_1382;
assign n_1503 = n_169 & n_1382;
assign n_1504 = n_168 & n_1382;
assign n_1505 = n_167 & n_1382;
assign n_1506 = n_166 & n_1382;
assign n_1507 = n_165 & n_1382;
assign n_1508 = n_164 & n_1382;
assign n_1509 = n_1382 & n_163;
assign n_1510 = n_1382 ^ n_1120;
assign n_1511 = n_1383 ^ x382;
assign n_1512 = n_1384 ^ x381;
assign n_1513 = n_1385 ^ x380;
assign n_1514 = n_1386 ^ x379;
assign n_1515 = n_1387 ^ x378;
assign n_1516 = n_1388 ^ x377;
assign n_1517 = n_1389 ^ x376;
assign n_1518 = n_1390 ^ x375;
assign n_1519 = n_1391 ^ x374;
assign n_1520 = n_1392 ^ x373;
assign n_1521 = n_1393 ^ x372;
assign n_1522 = n_1394 ^ x371;
assign n_1523 = n_1395 ^ x370;
assign n_1524 = n_1396 ^ x369;
assign n_1525 = n_1397 ^ x368;
assign n_1526 = n_1398 ^ x367;
assign n_1527 = n_1399 ^ x366;
assign n_1528 = n_1400 ^ x365;
assign n_1529 = n_1401 ^ x364;
assign n_1530 = n_1402 ^ x363;
assign n_1531 = n_1403 ^ x362;
assign n_1532 = n_1404 ^ x361;
assign n_1533 = n_1405 ^ x360;
assign n_1534 = n_1406 ^ x359;
assign n_1535 = n_1407 ^ x358;
assign n_1536 = n_1408 ^ x357;
assign n_1537 = n_1409 ^ x356;
assign n_1538 = n_1410 ^ x355;
assign n_1539 = n_1411 ^ x354;
assign n_1540 = n_1412 ^ x353;
assign n_1541 = n_1413 ^ x352;
assign n_1542 = n_1414 ^ x351;
assign n_1543 = n_1415 ^ x350;
assign n_1544 = n_1416 ^ x349;
assign n_1545 = n_1417 ^ x348;
assign n_1546 = n_1418 ^ x347;
assign n_1547 = n_1419 ^ x346;
assign n_1548 = n_1420 ^ x345;
assign n_1549 = n_1421 ^ x344;
assign n_1550 = n_1422 ^ x343;
assign n_1551 = n_1423 ^ x342;
assign n_1552 = n_1424 ^ x341;
assign n_1553 = n_1425 ^ x340;
assign n_1554 = n_1426 ^ x339;
assign n_1555 = n_1427 ^ x338;
assign n_1556 = n_1428 ^ x337;
assign n_1557 = n_1429 ^ x336;
assign n_1558 = n_1430 ^ x335;
assign n_1559 = n_1431 ^ x334;
assign n_1560 = n_1432 ^ x333;
assign n_1561 = n_1433 ^ x332;
assign n_1562 = n_1434 ^ x331;
assign n_1563 = n_1435 ^ x330;
assign n_1564 = n_1436 ^ x329;
assign n_1565 = n_1437 ^ x328;
assign n_1566 = n_1438 ^ x327;
assign n_1567 = n_1439 ^ x326;
assign n_1568 = n_1440 ^ x325;
assign n_1569 = n_1441 ^ x324;
assign n_1570 = n_1442 ^ x323;
assign n_1571 = n_1443 ^ x322;
assign n_1572 = n_1444 ^ x321;
assign n_1573 = n_1445 ^ x320;
assign n_1574 = n_1446 ^ x319;
assign n_1575 = n_1447 ^ x318;
assign n_1576 = n_1448 ^ x317;
assign n_1577 = n_1449 ^ x316;
assign n_1578 = n_1450 ^ x315;
assign n_1579 = n_1451 ^ x314;
assign n_1580 = n_1452 ^ x313;
assign n_1581 = n_1453 ^ x312;
assign n_1582 = n_1454 ^ x311;
assign n_1583 = n_1455 ^ x310;
assign n_1584 = n_1456 ^ x309;
assign n_1585 = n_1457 ^ x308;
assign n_1586 = n_1458 ^ x307;
assign n_1587 = n_1459 ^ x306;
assign n_1588 = n_1460 ^ x305;
assign n_1589 = n_1461 ^ x304;
assign n_1590 = n_1462 ^ x303;
assign n_1591 = n_1463 ^ x302;
assign n_1592 = n_1464 ^ x301;
assign n_1593 = n_1465 ^ x300;
assign n_1594 = n_1466 ^ x299;
assign n_1595 = n_1467 ^ x298;
assign n_1596 = n_1468 ^ x297;
assign n_1597 = n_1469 ^ x296;
assign n_1598 = n_1470 ^ x295;
assign n_1599 = n_1471 ^ x294;
assign n_1600 = n_1472 ^ x293;
assign n_1601 = n_1473 ^ x292;
assign n_1602 = n_1474 ^ x291;
assign n_1603 = n_1475 ^ x290;
assign n_1604 = n_1476 ^ x289;
assign n_1605 = n_1477 ^ x288;
assign n_1606 = n_1478 ^ x287;
assign n_1607 = n_1479 ^ x286;
assign n_1608 = n_1480 ^ x285;
assign n_1609 = n_1481 ^ x284;
assign n_1610 = n_1482 ^ x283;
assign n_1611 = n_1483 ^ x282;
assign n_1612 = n_1484 ^ x281;
assign n_1613 = n_1485 ^ x280;
assign n_1614 = n_1486 ^ x279;
assign n_1615 = n_1487 ^ x278;
assign n_1616 = n_1488 ^ x277;
assign n_1617 = n_1489 ^ x276;
assign n_1618 = n_1490 ^ x275;
assign n_1619 = n_1491 ^ x274;
assign n_1620 = n_1492 ^ x273;
assign n_1621 = n_1493 ^ x272;
assign n_1622 = n_1494 ^ x271;
assign n_1623 = n_1495 ^ x270;
assign n_1624 = n_1496 ^ x269;
assign n_1625 = n_1497 ^ x268;
assign n_1626 = n_1498 ^ x267;
assign n_1627 = n_1499 ^ x266;
assign n_1628 = n_1500 ^ x265;
assign n_1629 = n_1501 ^ x264;
assign n_1630 = n_1502 ^ x263;
assign n_1631 = n_1503 ^ x262;
assign n_1632 = n_1504 ^ x261;
assign n_1633 = n_1505 ^ x260;
assign n_1634 = n_1506 ^ x259;
assign n_1635 = n_1507 ^ x258;
assign n_1636 = n_1508 ^ x257;
assign n_1637 = n_1509 ^ x256;
assign n_1638 = n_1511 ^ n_318;
assign n_1639 = n_1511 ^ n_1250;
assign n_1640 = n_1251 ^ n_1512;
assign n_1641 = n_1252 ^ n_1513;
assign n_1642 = n_1253 ^ n_1514;
assign n_1643 = n_1254 ^ n_1515;
assign n_1644 = n_1255 ^ n_1516;
assign n_1645 = n_1517 ^ n_1256;
assign n_1646 = n_1257 ^ n_1518;
assign n_1647 = n_1258 ^ n_1519;
assign n_1648 = n_1259 ^ n_1520;
assign n_1649 = n_1521 ^ n_1260;
assign n_1650 = n_1522 ^ n_1261;
assign n_1651 = n_1262 ^ n_1523;
assign n_1652 = n_1263 ^ n_1524;
assign n_1653 = n_1264 ^ n_1525;
assign n_1654 = n_1265 ^ n_1526;
assign n_1655 = n_1527 ^ n_1266;
assign n_1656 = n_1528 ^ n_1267;
assign n_1657 = n_1529 ^ n_1268;
assign n_1658 = n_1269 ^ n_1530;
assign n_1659 = n_1270 ^ n_1531;
assign n_1660 = n_1271 ^ n_1532;
assign n_1661 = n_1533 ^ n_1272;
assign n_1662 = n_1534 ^ n_1273;
assign n_1663 = n_1274 ^ n_1535;
assign n_1664 = n_1536 ^ n_1275;
assign n_1665 = n_1537 ^ n_1276;
assign n_1666 = n_1277 ^ n_1538;
assign n_1667 = n_1278 ^ n_1539;
assign n_1668 = n_1540 ^ n_1279;
assign n_1669 = n_1280 ^ n_1541;
assign n_1670 = n_1281 ^ n_1542;
assign n_1671 = n_1282 ^ n_1543;
assign n_1672 = n_1283 ^ n_1544;
assign n_1673 = n_1545 ^ n_1284;
assign n_1674 = n_1546 ^ n_1285;
assign n_1675 = n_1547 ^ n_1286;
assign n_1676 = n_1287 ^ n_1548;
assign n_1677 = n_1549 ^ n_1288;
assign n_1678 = n_1550 ^ n_1289;
assign n_1679 = n_1551 ^ n_1290;
assign n_1680 = n_1552 ^ n_1291;
assign n_1681 = n_1292 ^ n_1553;
assign n_1682 = n_1554 ^ n_1293;
assign n_1683 = n_1294 ^ n_1555;
assign n_1684 = n_1556 ^ n_1295;
assign n_1685 = n_1557 ^ n_1296;
assign n_1686 = n_1558 ^ n_1297;
assign n_1687 = n_1298 ^ n_1559;
assign n_1688 = n_1560 ^ n_1299;
assign n_1689 = n_1300 ^ n_1561;
assign n_1690 = n_1301 ^ n_1562;
assign n_1691 = n_1302 ^ n_1563;
assign n_1692 = n_1303 ^ n_1564;
assign n_1693 = n_1565 ^ n_1304;
assign n_1694 = n_1566 ^ n_1305;
assign n_1695 = n_1306 ^ n_1567;
assign n_1696 = n_1568 ^ n_1307;
assign n_1697 = n_1308 ^ n_1569;
assign n_1698 = n_1570 ^ n_1309;
assign n_1699 = n_1571 ^ n_1310;
assign n_1700 = n_1311 ^ n_1572;
assign n_1701 = n_1573 ^ n_1312;
assign n_1702 = n_1313 ^ n_1574;
assign n_1703 = n_1575 ^ n_1314;
assign n_1704 = n_1576 ^ n_1315;
assign n_1705 = n_1577 ^ n_1316;
assign n_1706 = n_1578 ^ n_1317;
assign n_1707 = n_1318 ^ n_1579;
assign n_1708 = n_1319 ^ n_1580;
assign n_1709 = n_1581 ^ n_1320;
assign n_1710 = n_1582 ^ n_1321;
assign n_1711 = n_1583 ^ n_1322;
assign n_1712 = n_1323 ^ n_1584;
assign n_1713 = n_1585 ^ n_1324;
assign n_1714 = n_1325 ^ n_1586;
assign n_1715 = n_1587 ^ n_1326;
assign n_1716 = n_1588 ^ n_1327;
assign n_1717 = n_1328 ^ n_1589;
assign n_1718 = n_1590 ^ n_1329;
assign n_1719 = n_1591 ^ n_1330;
assign n_1720 = n_1592 ^ n_1331;
assign n_1721 = n_1593 ^ n_1332;
assign n_1722 = n_1333 ^ n_1594;
assign n_1723 = n_1595 ^ n_1334;
assign n_1724 = n_1596 ^ n_1335;
assign n_1725 = n_1597 ^ n_1336;
assign n_1726 = n_1598 ^ n_1337;
assign n_1727 = n_1599 ^ n_1338;
assign n_1728 = n_1339 ^ n_1600;
assign n_1729 = n_1601 ^ n_1340;
assign n_1730 = n_1341 ^ n_1602;
assign n_1731 = n_1342 ^ n_1603;
assign n_1732 = n_1604 ^ n_1343;
assign n_1733 = n_1605 ^ n_1344;
assign n_1734 = n_1606 ^ n_1345;
assign n_1735 = n_1346 ^ n_1607;
assign n_1736 = n_1608 ^ n_1347;
assign n_1737 = n_1609 ^ n_1348;
assign n_1738 = n_1349 ^ n_1610;
assign n_1739 = n_1611 ^ n_1350;
assign n_1740 = n_1612 ^ n_1351;
assign n_1741 = n_1613 ^ n_1352;
assign n_1742 = n_1614 ^ n_1353;
assign n_1743 = n_1354 ^ n_1615;
assign n_1744 = n_1355 ^ n_1616;
assign n_1745 = n_1617 ^ n_1356;
assign n_1746 = n_1357 ^ n_1618;
assign n_1747 = n_1619 ^ n_1358;
assign n_1748 = n_1620 ^ n_1359;
assign n_1749 = n_1360 ^ n_1621;
assign n_1750 = n_1622 ^ n_1361;
assign n_1751 = n_1623 ^ n_1362;
assign n_1752 = n_1363 ^ n_1624;
assign n_1753 = n_1364 ^ n_1625;
assign n_1754 = n_1626 ^ n_1365;
assign n_1755 = n_1366 ^ n_1627;
assign n_1756 = n_1367 ^ n_1628;
assign n_1757 = n_1368 ^ n_1629;
assign n_1758 = n_1630 ^ n_1369;
assign n_1759 = n_1370 ^ n_1631;
assign n_1760 = n_1632 ^ n_1371;
assign n_1761 = n_1633 ^ n_1372;
assign n_1762 = n_1634 ^ n_1373;
assign n_1763 = n_1374 ^ n_1635;
assign n_1764 = n_1375 ^ n_1636;
assign n_1765 = ~n_1637 & n_1376;
assign n_1766 = n_1376 ^ n_1637;
assign n_1767 = n_1765 ^ n_1375;
assign n_1768 = ~n_1764 & n_1767;
assign n_1769 = n_1375 ^ n_1768;
assign n_1770 = n_1769 ^ n_1374;
assign n_1771 = ~n_1763 & n_1770;
assign n_1772 = n_1374 ^ n_1771;
assign n_1773 = n_1772 ^ n_1373;
assign n_1774 = ~n_1762 & ~n_1773;
assign n_1775 = n_1634 ^ n_1774;
assign n_1776 = n_1775 ^ n_1633;
assign n_1777 = ~n_1761 & ~n_1776;
assign n_1778 = n_1372 ^ n_1777;
assign n_1779 = n_1778 ^ n_1632;
assign n_1780 = ~n_1760 & ~n_1779;
assign n_1781 = n_1632 ^ n_1780;
assign n_1782 = n_1781 ^ n_1370;
assign n_1783 = ~n_1759 & n_1782;
assign n_1784 = n_1631 ^ n_1783;
assign n_1785 = n_1784 ^ n_1630;
assign n_1786 = ~n_1758 & ~n_1785;
assign n_1787 = n_1369 ^ n_1786;
assign n_1788 = n_1787 ^ n_1368;
assign n_1789 = ~n_1757 & n_1788;
assign n_1790 = n_1368 ^ n_1789;
assign n_1791 = n_1790 ^ n_1367;
assign n_1792 = ~n_1756 & n_1791;
assign n_1793 = n_1367 ^ n_1792;
assign n_1794 = n_1793 ^ n_1627;
assign n_1795 = ~n_1755 & ~n_1794;
assign n_1796 = n_1627 ^ n_1795;
assign n_1797 = n_1796 ^ n_1626;
assign n_1798 = ~n_1754 & n_1797;
assign n_1799 = n_1626 ^ n_1798;
assign n_1800 = n_1799 ^ n_1625;
assign n_1801 = ~n_1753 & n_1800;
assign n_1802 = n_1625 ^ n_1801;
assign n_1803 = n_1802 ^ n_1363;
assign n_1804 = ~n_1752 & ~n_1803;
assign n_1805 = n_1363 ^ n_1804;
assign n_1806 = n_1805 ^ n_1362;
assign n_1807 = ~n_1751 & ~n_1806;
assign n_1808 = n_1623 ^ n_1807;
assign n_1809 = n_1808 ^ n_1622;
assign n_1810 = ~n_1750 & ~n_1809;
assign n_1811 = n_1361 ^ n_1810;
assign n_1812 = n_1811 ^ n_1360;
assign n_1813 = ~n_1749 & n_1812;
assign n_1814 = n_1360 ^ n_1813;
assign n_1815 = n_1814 ^ n_1620;
assign n_1816 = ~n_1748 & n_1815;
assign n_1817 = n_1359 ^ n_1816;
assign n_1818 = n_1817 ^ n_1619;
assign n_1819 = ~n_1747 & ~n_1818;
assign n_1820 = n_1619 ^ n_1819;
assign n_1821 = n_1820 ^ n_1357;
assign n_1822 = ~n_1746 & n_1821;
assign n_1823 = n_1618 ^ n_1822;
assign n_1824 = n_1823 ^ n_1617;
assign n_1825 = ~n_1745 & ~n_1824;
assign n_1826 = n_1356 ^ n_1825;
assign n_1827 = n_1826 ^ n_1355;
assign n_1828 = ~n_1744 & n_1827;
assign n_1829 = n_1355 ^ n_1828;
assign n_1830 = n_1829 ^ n_1354;
assign n_1831 = ~n_1743 & n_1830;
assign n_1832 = n_1354 ^ n_1831;
assign n_1833 = n_1832 ^ n_1353;
assign n_1834 = ~n_1742 & ~n_1833;
assign n_1835 = n_1614 ^ n_1834;
assign n_1836 = n_1835 ^ n_1613;
assign n_1837 = ~n_1741 & ~n_1836;
assign n_1838 = n_1352 ^ n_1837;
assign n_1839 = n_1838 ^ n_1612;
assign n_1840 = ~n_1740 & ~n_1839;
assign n_1841 = n_1612 ^ n_1840;
assign n_1842 = n_1841 ^ n_1611;
assign n_1843 = ~n_1739 & ~n_1842;
assign n_1844 = n_1350 ^ n_1843;
assign n_1845 = n_1844 ^ n_1349;
assign n_1846 = ~n_1738 & n_1845;
assign n_1847 = n_1349 ^ n_1846;
assign n_1848 = n_1847 ^ n_1609;
assign n_1849 = ~n_1737 & n_1848;
assign n_1850 = n_1348 ^ n_1849;
assign n_1851 = n_1850 ^ n_1608;
assign n_1852 = ~n_1736 & n_1851;
assign n_1853 = n_1347 ^ n_1852;
assign n_1854 = n_1853 ^ n_1346;
assign n_1855 = ~n_1735 & n_1854;
assign n_1856 = n_1346 ^ n_1855;
assign n_1857 = n_1856 ^ n_1606;
assign n_1858 = ~n_1734 & n_1857;
assign n_1859 = n_1345 ^ n_1858;
assign n_1860 = n_1859 ^ n_1605;
assign n_1861 = ~n_1733 & ~n_1860;
assign n_1862 = n_1605 ^ n_1861;
assign n_1863 = n_1862 ^ n_1604;
assign n_1864 = ~n_1732 & ~n_1863;
assign n_1865 = n_1343 ^ n_1864;
assign n_1866 = n_1865 ^ n_1342;
assign n_1867 = ~n_1731 & n_1866;
assign n_1868 = n_1342 ^ n_1867;
assign n_1869 = n_1868 ^ n_1602;
assign n_1870 = ~n_1730 & n_1869;
assign n_1871 = n_1341 ^ n_1870;
assign n_1872 = n_1871 ^ n_1601;
assign n_1873 = ~n_1729 & n_1872;
assign n_1874 = n_1340 ^ n_1873;
assign n_1875 = n_1874 ^ n_1339;
assign n_1876 = ~n_1728 & n_1875;
assign n_1877 = n_1339 ^ n_1876;
assign n_1878 = n_1877 ^ n_1599;
assign n_1879 = ~n_1727 & n_1878;
assign n_1880 = n_1338 ^ n_1879;
assign n_1881 = n_1880 ^ n_1598;
assign n_1882 = ~n_1726 & ~n_1881;
assign n_1883 = n_1598 ^ n_1882;
assign n_1884 = n_1883 ^ n_1597;
assign n_1885 = ~n_1725 & ~n_1884;
assign n_1886 = n_1336 ^ n_1885;
assign n_1887 = n_1886 ^ n_1596;
assign n_1888 = ~n_1724 & n_1887;
assign n_1889 = n_1335 ^ n_1888;
assign n_1890 = n_1889 ^ n_1595;
assign n_1891 = ~n_1723 & ~n_1890;
assign n_1892 = n_1595 ^ n_1891;
assign n_1893 = n_1892 ^ n_1333;
assign n_1894 = ~n_1722 & ~n_1893;
assign n_1895 = n_1333 ^ n_1894;
assign n_1896 = n_1895 ^ n_1332;
assign n_1897 = ~n_1721 & ~n_1896;
assign n_1898 = n_1593 ^ n_1897;
assign n_1899 = n_1898 ^ n_1592;
assign n_1900 = ~n_1720 & ~n_1899;
assign n_1901 = n_1331 ^ n_1900;
assign n_1902 = n_1901 ^ n_1591;
assign n_1903 = ~n_1719 & ~n_1902;
assign n_1904 = n_1591 ^ n_1903;
assign n_1905 = n_1904 ^ n_1590;
assign n_1906 = ~n_1718 & ~n_1905;
assign n_1907 = n_1329 ^ n_1906;
assign n_1908 = n_1907 ^ n_1328;
assign n_1909 = ~n_1717 & n_1908;
assign n_1910 = n_1328 ^ n_1909;
assign n_1911 = n_1910 ^ n_1588;
assign n_1912 = ~n_1716 & ~n_1911;
assign n_1913 = n_1588 ^ n_1912;
assign n_1914 = n_1913 ^ n_1326;
assign n_1915 = ~n_1715 & ~n_1914;
assign n_1916 = n_1326 ^ n_1915;
assign n_1917 = n_1916 ^ n_1325;
assign n_1918 = ~n_1714 & ~n_1917;
assign n_1919 = n_1586 ^ n_1918;
assign n_1920 = n_1919 ^ n_1585;
assign n_1921 = ~n_1713 & ~n_1920;
assign n_1922 = n_1324 ^ n_1921;
assign n_1923 = n_1922 ^ n_1323;
assign n_1924 = ~n_1712 & n_1923;
assign n_1925 = n_1323 ^ n_1924;
assign n_1926 = n_1925 ^ n_1583;
assign n_1927 = ~n_1711 & ~n_1926;
assign n_1928 = n_1583 ^ n_1927;
assign n_1929 = n_1928 ^ n_1321;
assign n_1930 = ~n_1710 & n_1929;
assign n_1931 = n_1582 ^ n_1930;
assign n_1932 = n_1931 ^ n_1581;
assign n_1933 = ~n_1709 & ~n_1932;
assign n_1934 = n_1320 ^ n_1933;
assign n_1935 = n_1934 ^ n_1319;
assign n_1936 = ~n_1708 & n_1935;
assign n_1937 = n_1319 ^ n_1936;
assign n_1938 = n_1937 ^ n_1318;
assign n_1939 = ~n_1707 & n_1938;
assign n_1940 = n_1318 ^ n_1939;
assign n_1941 = n_1940 ^ n_1317;
assign n_1942 = ~n_1706 & n_1941;
assign n_1943 = n_1317 ^ n_1942;
assign n_1944 = n_1943 ^ n_1577;
assign n_1945 = ~n_1705 & ~n_1944;
assign n_1946 = n_1577 ^ n_1945;
assign n_1947 = n_1946 ^ n_1315;
assign n_1948 = ~n_1704 & ~n_1947;
assign n_1949 = n_1315 ^ n_1948;
assign n_1950 = n_1949 ^ n_1575;
assign n_1951 = ~n_1703 & ~n_1950;
assign n_1952 = n_1575 ^ n_1951;
assign n_1953 = n_1952 ^ n_1574;
assign n_1954 = ~n_1702 & n_1953;
assign n_1955 = n_1574 ^ n_1954;
assign n_1956 = n_1955 ^ n_1573;
assign n_1957 = ~n_1701 & n_1956;
assign n_1958 = n_1573 ^ n_1957;
assign n_1959 = n_1958 ^ n_1572;
assign n_1960 = ~n_1700 & n_1959;
assign n_1961 = n_1572 ^ n_1960;
assign n_1962 = n_1961 ^ n_1571;
assign n_1963 = ~n_1699 & ~n_1962;
assign n_1964 = n_1310 ^ n_1963;
assign n_1965 = n_1964 ^ n_1570;
assign n_1966 = ~n_1698 & n_1965;
assign n_1967 = n_1309 ^ n_1966;
assign n_1968 = n_1967 ^ n_1308;
assign n_1969 = ~n_1697 & n_1968;
assign n_1970 = n_1308 ^ n_1969;
assign n_1971 = n_1970 ^ n_1568;
assign n_1972 = ~n_1696 & ~n_1971;
assign n_1973 = n_1568 ^ n_1972;
assign n_1974 = n_1973 ^ n_1567;
assign n_1975 = ~n_1695 & ~n_1974;
assign n_1976 = n_1306 ^ n_1975;
assign n_1977 = n_1976 ^ n_1566;
assign n_1978 = ~n_1694 & n_1977;
assign n_1979 = n_1305 ^ n_1978;
assign n_1980 = n_1979 ^ n_1565;
assign n_1981 = ~n_1693 & ~n_1980;
assign n_1982 = n_1565 ^ n_1981;
assign n_1983 = n_1982 ^ n_1303;
assign n_1984 = ~n_1692 & ~n_1983;
assign n_1985 = n_1303 ^ n_1984;
assign n_1986 = n_1985 ^ n_1302;
assign n_1987 = ~n_1691 & n_1986;
assign n_1988 = n_1302 ^ n_1987;
assign n_1989 = n_1988 ^ n_1562;
assign n_1990 = ~n_1690 & ~n_1989;
assign n_1991 = n_1562 ^ n_1990;
assign n_1992 = n_1991 ^ n_1300;
assign n_1993 = ~n_1689 & ~n_1992;
assign n_1994 = n_1300 ^ n_1993;
assign n_1995 = n_1994 ^ n_1299;
assign n_1996 = ~n_1688 & ~n_1995;
assign n_1997 = n_1560 ^ n_1996;
assign n_1998 = n_1997 ^ n_1298;
assign n_1999 = ~n_1687 & n_1998;
assign n_2000 = n_1559 ^ n_1999;
assign n_2001 = n_2000 ^ n_1297;
assign n_2002 = ~n_1686 & ~n_2001;
assign n_2003 = n_1297 ^ n_2002;
assign n_2004 = n_2003 ^ n_1557;
assign n_2005 = ~n_1685 & n_2004;
assign n_2006 = n_1296 ^ n_2005;
assign n_2007 = n_2006 ^ n_1556;
assign n_2008 = ~n_1684 & n_2007;
assign n_2009 = n_1295 ^ n_2008;
assign n_2010 = n_2009 ^ n_1555;
assign n_2011 = ~n_1683 & ~n_2010;
assign n_2012 = n_1555 ^ n_2011;
assign n_2013 = n_2012 ^ n_1293;
assign n_2014 = ~n_1682 & ~n_2013;
assign n_2015 = n_1293 ^ n_2014;
assign n_2016 = n_2015 ^ n_1292;
assign n_2017 = ~n_1681 & n_2016;
assign n_2018 = n_1292 ^ n_2017;
assign n_2019 = n_2018 ^ n_1291;
assign n_2020 = ~n_1680 & n_2019;
assign n_2021 = n_1291 ^ n_2020;
assign n_2022 = n_2021 ^ n_1290;
assign n_2023 = ~n_1679 & n_2022;
assign n_2024 = n_1290 ^ n_2023;
assign n_2025 = n_2024 ^ n_1289;
assign n_2026 = ~n_1678 & n_2025;
assign n_2027 = n_1289 ^ n_2026;
assign n_2028 = n_2027 ^ n_1549;
assign n_2029 = ~n_1677 & ~n_2028;
assign n_2030 = n_1549 ^ n_2029;
assign n_2031 = n_2030 ^ n_1548;
assign n_2032 = ~n_1676 & n_2031;
assign n_2033 = n_1548 ^ n_2032;
assign n_2034 = n_2033 ^ n_1547;
assign n_2035 = ~n_1675 & n_2034;
assign n_2036 = n_1547 ^ n_2035;
assign n_2037 = n_2036 ^ n_1285;
assign n_2038 = ~n_1674 & ~n_2037;
assign n_2039 = n_1285 ^ n_2038;
assign n_2040 = n_2039 ^ n_1284;
assign n_2041 = ~n_1673 & ~n_2040;
assign n_2042 = n_1545 ^ n_2041;
assign n_2043 = n_2042 ^ n_1283;
assign n_2044 = ~n_1672 & n_2043;
assign n_2045 = n_1544 ^ n_2044;
assign n_2046 = n_2045 ^ n_1543;
assign n_2047 = ~n_1671 & n_2046;
assign n_2048 = n_1543 ^ n_2047;
assign n_2049 = n_2048 ^ n_1542;
assign n_2050 = ~n_1670 & n_2049;
assign n_2051 = n_1542 ^ n_2050;
assign n_2052 = n_2051 ^ n_1541;
assign n_2053 = ~n_1669 & ~n_2052;
assign n_2054 = n_1280 ^ n_2053;
assign n_2055 = n_2054 ^ n_1540;
assign n_2056 = ~n_1668 & n_2055;
assign n_2057 = n_1279 ^ n_2056;
assign n_2058 = n_2057 ^ n_1539;
assign n_2059 = ~n_1667 & ~n_2058;
assign n_2060 = n_1539 ^ n_2059;
assign n_2061 = n_2060 ^ n_1538;
assign n_2062 = ~n_1666 & n_2061;
assign n_2063 = n_1538 ^ n_2062;
assign n_2064 = n_2063 ^ n_1537;
assign n_2065 = ~n_1665 & ~n_2064;
assign n_2066 = n_1276 ^ n_2065;
assign n_2067 = n_2066 ^ n_1536;
assign n_2068 = ~n_1664 & n_2067;
assign n_2069 = n_1275 ^ n_2068;
assign n_2070 = n_2069 ^ n_1535;
assign n_2071 = ~n_1663 & ~n_2070;
assign n_2072 = n_1535 ^ n_2071;
assign n_2073 = n_2072 ^ n_1273;
assign n_2074 = ~n_1662 & n_2073;
assign n_2075 = n_1534 ^ n_2074;
assign n_2076 = n_2075 ^ n_1533;
assign n_2077 = ~n_1661 & ~n_2076;
assign n_2078 = n_1272 ^ n_2077;
assign n_2079 = n_2078 ^ n_1532;
assign n_2080 = ~n_1660 & ~n_2079;
assign n_2081 = n_1532 ^ n_2080;
assign n_2082 = n_2081 ^ n_1270;
assign n_2083 = ~n_1659 & n_2082;
assign n_2084 = n_1531 ^ n_2083;
assign n_2085 = n_2084 ^ n_1269;
assign n_2086 = ~n_1658 & n_2085;
assign n_2087 = n_1530 ^ n_2086;
assign n_2088 = n_2087 ^ n_1529;
assign n_2089 = ~n_1657 & n_2088;
assign n_2090 = n_1529 ^ n_2089;
assign n_2091 = n_2090 ^ n_1528;
assign n_2092 = ~n_1656 & ~n_2091;
assign n_2093 = n_1267 ^ n_2092;
assign n_2094 = n_2093 ^ n_1527;
assign n_2095 = ~n_1655 & n_2094;
assign n_2096 = n_1266 ^ n_2095;
assign n_2097 = n_2096 ^ n_1526;
assign n_2098 = ~n_1654 & ~n_2097;
assign n_2099 = n_1526 ^ n_2098;
assign n_2100 = n_2099 ^ n_1525;
assign n_2101 = ~n_1653 & n_2100;
assign n_2102 = n_1525 ^ n_2101;
assign n_2103 = n_2102 ^ n_1263;
assign n_2104 = ~n_1652 & ~n_2103;
assign n_2105 = n_1263 ^ n_2104;
assign n_2106 = n_2105 ^ n_1523;
assign n_2107 = ~n_1651 & ~n_2106;
assign n_2108 = n_1523 ^ n_2107;
assign n_2109 = n_2108 ^ n_1522;
assign n_2110 = ~n_1650 & n_2109;
assign n_2111 = n_1522 ^ n_2110;
assign n_2112 = n_2111 ^ n_1260;
assign n_2113 = ~n_1649 & ~n_2112;
assign n_2114 = n_1260 ^ n_2113;
assign n_2115 = n_2114 ^ n_1259;
assign n_2116 = ~n_1648 & n_2115;
assign n_2117 = n_1259 ^ n_2116;
assign n_2118 = n_2117 ^ n_1258;
assign n_2119 = ~n_1647 & ~n_2118;
assign n_2120 = n_1519 ^ n_2119;
assign n_2121 = n_2120 ^ n_1257;
assign n_2122 = ~n_1646 & n_2121;
assign n_2123 = n_1518 ^ n_2122;
assign n_2124 = n_2123 ^ n_1517;
assign n_2125 = ~n_1645 & n_2124;
assign n_2126 = n_1517 ^ n_2125;
assign n_2127 = n_2126 ^ n_1516;
assign n_2128 = ~n_1644 & ~n_2127;
assign n_2129 = n_1255 ^ n_2128;
assign n_2130 = n_2129 ^ n_1254;
assign n_2131 = ~n_1643 & ~n_2130;
assign n_2132 = n_1515 ^ n_2131;
assign n_2133 = n_2132 ^ n_1514;
assign n_2134 = ~n_1642 & n_2133;
assign n_2135 = n_1514 ^ n_2134;
assign n_2136 = n_2135 ^ n_1513;
assign n_2137 = ~n_1641 & n_2136;
assign n_2138 = n_1513 ^ n_2137;
assign n_2139 = n_2138 ^ n_1251;
assign n_2140 = ~n_1640 & ~n_2139;
assign n_2141 = n_1251 ^ n_2140;
assign n_2142 = n_2141 ^ n_1250;
assign n_2143 = ~n_1639 & ~n_2142;
assign n_2144 = n_1638 ^ n_2143;
assign n_2145 = ~n_377 & n_2144;
assign n_2146 = n_160 ^ n_2145;
assign n_2147 = ~n_2146 & n_1766;
assign n_2148 = n_1764 & ~n_2146;
assign n_2149 = n_1763 & ~n_2146;
assign n_2150 = n_1762 & ~n_2146;
assign n_2151 = n_1761 & n_2146;
assign n_2152 = n_1760 & n_2146;
assign n_2153 = n_1759 & ~n_2146;
assign n_2154 = n_1758 & n_2146;
assign n_2155 = n_1757 & ~n_2146;
assign n_2156 = n_1756 & ~n_2146;
assign n_2157 = n_1755 & n_2146;
assign n_2158 = n_1754 & n_2146;
assign n_2159 = n_1753 & n_2146;
assign n_2160 = n_1752 & ~n_2146;
assign n_2161 = n_1751 & ~n_2146;
assign n_2162 = n_1750 & n_2146;
assign n_2163 = n_1749 & ~n_2146;
assign n_2164 = n_1748 & n_2146;
assign n_2165 = n_1747 & n_2146;
assign n_2166 = n_1746 & ~n_2146;
assign n_2167 = n_1745 & n_2146;
assign n_2168 = n_1744 & ~n_2146;
assign n_2169 = n_1743 & ~n_2146;
assign n_2170 = n_1742 & ~n_2146;
assign n_2171 = n_1741 & n_2146;
assign n_2172 = n_1740 & n_2146;
assign n_2173 = n_1739 & n_2146;
assign n_2174 = n_1738 & ~n_2146;
assign n_2175 = n_1737 & n_2146;
assign n_2176 = n_1736 & n_2146;
assign n_2177 = n_1735 & ~n_2146;
assign n_2178 = n_1734 & n_2146;
assign n_2179 = n_1733 & n_2146;
assign n_2180 = n_1732 & n_2146;
assign n_2181 = n_1731 & ~n_2146;
assign n_2182 = n_1730 & n_2146;
assign n_2183 = n_1729 & n_2146;
assign n_2184 = n_1728 & ~n_2146;
assign n_2185 = n_1727 & n_2146;
assign n_2186 = n_1726 & n_2146;
assign n_2187 = n_1725 & n_2146;
assign n_2188 = n_1724 & n_2146;
assign n_2189 = n_1723 & n_2146;
assign n_2190 = n_1722 & ~n_2146;
assign n_2191 = n_1721 & ~n_2146;
assign n_2192 = n_1720 & n_2146;
assign n_2193 = n_1719 & n_2146;
assign n_2194 = n_1718 & n_2146;
assign n_2195 = n_1717 & ~n_2146;
assign n_2196 = n_1716 & n_2146;
assign n_2197 = n_1715 & ~n_2146;
assign n_2198 = n_1714 & ~n_2146;
assign n_2199 = n_1713 & n_2146;
assign n_2200 = n_1712 & ~n_2146;
assign n_2201 = n_1711 & n_2146;
assign n_2202 = n_1710 & ~n_2146;
assign n_2203 = n_1709 & n_2146;
assign n_2204 = n_1708 & ~n_2146;
assign n_2205 = n_1707 & ~n_2146;
assign n_2206 = n_1706 & ~n_2146;
assign n_2207 = n_1705 & n_2146;
assign n_2208 = n_1704 & ~n_2146;
assign n_2209 = n_1703 & n_2146;
assign n_2210 = n_1702 & n_2146;
assign n_2211 = n_1701 & n_2146;
assign n_2212 = n_1700 & n_2146;
assign n_2213 = n_1699 & n_2146;
assign n_2214 = n_1698 & n_2146;
assign n_2215 = n_1697 & ~n_2146;
assign n_2216 = n_1696 & n_2146;
assign n_2217 = n_1695 & n_2146;
assign n_2218 = n_1694 & n_2146;
assign n_2219 = n_1693 & n_2146;
assign n_2220 = n_1692 & ~n_2146;
assign n_2221 = n_1691 & n_2146;
assign n_2222 = n_1690 & ~n_2146;
assign n_2223 = n_1689 & n_2146;
assign n_2224 = n_1688 & ~n_2146;
assign n_2225 = n_1687 & ~n_2146;
assign n_2226 = n_1686 & n_2146;
assign n_2227 = n_1685 & n_2146;
assign n_2228 = n_1684 & n_2146;
assign n_2229 = n_1683 & ~n_2146;
assign n_2230 = n_1682 & n_2146;
assign n_2231 = n_1681 & n_2146;
assign n_2232 = n_1680 & n_2146;
assign n_2233 = n_1679 & ~n_2146;
assign n_2234 = n_1678 & n_2146;
assign n_2235 = n_1677 & ~n_2146;
assign n_2236 = n_1676 & ~n_2146;
assign n_2237 = n_1675 & ~n_2146;
assign n_2238 = n_1674 & n_2146;
assign n_2239 = n_1673 & ~n_2146;
assign n_2240 = n_1672 & ~n_2146;
assign n_2241 = n_1671 & ~n_2146;
assign n_2242 = n_1670 & ~n_2146;
assign n_2243 = n_1669 & n_2146;
assign n_2244 = n_1668 & n_2146;
assign n_2245 = n_1667 & ~n_2146;
assign n_2246 = n_1666 & ~n_2146;
assign n_2247 = n_1665 & n_2146;
assign n_2248 = n_1664 & n_2146;
assign n_2249 = n_1663 & ~n_2146;
assign n_2250 = n_1662 & ~n_2146;
assign n_2251 = n_1661 & n_2146;
assign n_2252 = n_1660 & ~n_2146;
assign n_2253 = n_1659 & ~n_2146;
assign n_2254 = n_1658 & ~n_2146;
assign n_2255 = n_1657 & n_2146;
assign n_2256 = n_1656 & n_2146;
assign n_2257 = n_1655 & n_2146;
assign n_2258 = n_1654 & ~n_2146;
assign n_2259 = n_1653 & ~n_2146;
assign n_2260 = n_1652 & n_2146;
assign n_2261 = n_1651 & ~n_2146;
assign n_2262 = n_1650 & ~n_2146;
assign n_2263 = n_1649 & n_2146;
assign n_2264 = n_1648 & n_2146;
assign n_2265 = n_1647 & ~n_2146;
assign n_2266 = n_1646 & ~n_2146;
assign n_2267 = n_1645 & n_2146;
assign n_2268 = n_1644 & n_2146;
assign n_2269 = n_1643 & ~n_2146;
assign n_2270 = n_1642 & ~n_2146;
assign n_2271 = n_1641 & ~n_2146;
assign n_2272 = n_1640 & n_2146;
assign n_2273 = n_1639 & ~n_2146;
assign n_2274 = ~n_2146 & n_1510;
assign y129 = n_2146;
assign n_2275 = n_2147 ^ n_1637;
assign n_2276 = n_2148 ^ n_1636;
assign n_2277 = n_2149 ^ n_1635;
assign n_2278 = n_2150 ^ n_1634;
assign n_2279 = n_2151 ^ n_1372;
assign n_2280 = n_2152 ^ n_1371;
assign n_2281 = n_2153 ^ n_1631;
assign n_2282 = n_2154 ^ n_1369;
assign n_2283 = n_2155 ^ n_1629;
assign n_2284 = n_2156 ^ n_1628;
assign n_2285 = n_2157 ^ n_1366;
assign n_2286 = n_2158 ^ n_1365;
assign n_2287 = n_2159 ^ n_1364;
assign n_2288 = n_2160 ^ n_1624;
assign n_2289 = n_2161 ^ n_1623;
assign n_2290 = n_2162 ^ n_1361;
assign n_2291 = n_2163 ^ n_1621;
assign n_2292 = n_2164 ^ n_1359;
assign n_2293 = n_2165 ^ n_1358;
assign n_2294 = n_2166 ^ n_1618;
assign n_2295 = n_2167 ^ n_1356;
assign n_2296 = n_2168 ^ n_1616;
assign n_2297 = n_2169 ^ n_1615;
assign n_2298 = n_2170 ^ n_1614;
assign n_2299 = n_2171 ^ n_1352;
assign n_2300 = n_2172 ^ n_1351;
assign n_2301 = n_2173 ^ n_1350;
assign n_2302 = n_2174 ^ n_1610;
assign n_2303 = n_2175 ^ n_1348;
assign n_2304 = n_2176 ^ n_1347;
assign n_2305 = n_2177 ^ n_1607;
assign n_2306 = n_2178 ^ n_1345;
assign n_2307 = n_2179 ^ n_1344;
assign n_2308 = n_2180 ^ n_1343;
assign n_2309 = n_2181 ^ n_1603;
assign n_2310 = n_2182 ^ n_1341;
assign n_2311 = n_2183 ^ n_1340;
assign n_2312 = n_2184 ^ n_1600;
assign n_2313 = n_2185 ^ n_1338;
assign n_2314 = n_2186 ^ n_1337;
assign n_2315 = n_2187 ^ n_1336;
assign n_2316 = n_2188 ^ n_1335;
assign n_2317 = n_2189 ^ n_1334;
assign n_2318 = n_2190 ^ n_1594;
assign n_2319 = n_2191 ^ n_1593;
assign n_2320 = n_2192 ^ n_1331;
assign n_2321 = n_2193 ^ n_1330;
assign n_2322 = n_2194 ^ n_1329;
assign n_2323 = n_2195 ^ n_1589;
assign n_2324 = n_2196 ^ n_1327;
assign n_2325 = n_2197 ^ n_1587;
assign n_2326 = n_2198 ^ n_1586;
assign n_2327 = n_2199 ^ n_1324;
assign n_2328 = n_2200 ^ n_1584;
assign n_2329 = n_2201 ^ n_1322;
assign n_2330 = n_2202 ^ n_1582;
assign n_2331 = n_2203 ^ n_1320;
assign n_2332 = n_2204 ^ n_1580;
assign n_2333 = n_2205 ^ n_1579;
assign n_2334 = n_2206 ^ n_1578;
assign n_2335 = n_2207 ^ n_1316;
assign n_2336 = n_2208 ^ n_1576;
assign n_2337 = n_2209 ^ n_1314;
assign n_2338 = n_2210 ^ n_1313;
assign n_2339 = n_2211 ^ n_1312;
assign n_2340 = n_2212 ^ n_1311;
assign n_2341 = n_2213 ^ n_1310;
assign n_2342 = n_2214 ^ n_1309;
assign n_2343 = n_2215 ^ n_1569;
assign n_2344 = n_2216 ^ n_1307;
assign n_2345 = n_2217 ^ n_1306;
assign n_2346 = n_2218 ^ n_1305;
assign n_2347 = n_2219 ^ n_1304;
assign n_2348 = n_2220 ^ n_1564;
assign n_2349 = n_2221 ^ n_1302;
assign n_2350 = n_2222 ^ n_1562;
assign n_2351 = n_2223 ^ n_1300;
assign n_2352 = n_2224 ^ n_1560;
assign n_2353 = n_2225 ^ n_1559;
assign n_2354 = n_2226 ^ n_1297;
assign n_2355 = n_2227 ^ n_1296;
assign n_2356 = n_2228 ^ n_1295;
assign n_2357 = n_2229 ^ n_1555;
assign n_2358 = n_2230 ^ n_1293;
assign n_2359 = n_2231 ^ n_1292;
assign n_2360 = n_2232 ^ n_1291;
assign n_2361 = n_2233 ^ n_1551;
assign n_2362 = n_2234 ^ n_1289;
assign n_2363 = n_2235 ^ n_1549;
assign n_2364 = n_2236 ^ n_1548;
assign n_2365 = n_2237 ^ n_1547;
assign n_2366 = n_2238 ^ n_1285;
assign n_2367 = n_2239 ^ n_1545;
assign n_2368 = n_2240 ^ n_1544;
assign n_2369 = n_2241 ^ n_1543;
assign n_2370 = n_2242 ^ n_1542;
assign n_2371 = n_2243 ^ n_1280;
assign n_2372 = n_2244 ^ n_1279;
assign n_2373 = n_2245 ^ n_1539;
assign n_2374 = n_2246 ^ n_1538;
assign n_2375 = n_2247 ^ n_1276;
assign n_2376 = n_2248 ^ n_1275;
assign n_2377 = n_2249 ^ n_1535;
assign n_2378 = n_2250 ^ n_1534;
assign n_2379 = n_2251 ^ n_1272;
assign n_2380 = n_2252 ^ n_1532;
assign n_2381 = n_2253 ^ n_1531;
assign n_2382 = n_2254 ^ n_1530;
assign n_2383 = n_2255 ^ n_1268;
assign n_2384 = n_2256 ^ n_1267;
assign n_2385 = n_2257 ^ n_1266;
assign n_2386 = n_2258 ^ n_1526;
assign n_2387 = n_2259 ^ n_1525;
assign n_2388 = n_2260 ^ n_1263;
assign n_2389 = n_2261 ^ n_1523;
assign n_2390 = n_2262 ^ n_1522;
assign n_2391 = n_2263 ^ n_1260;
assign n_2392 = n_2264 ^ n_1259;
assign n_2393 = n_2265 ^ n_1519;
assign n_2394 = n_2266 ^ n_1518;
assign n_2395 = n_2267 ^ n_1256;
assign n_2396 = n_2268 ^ n_1255;
assign n_2397 = n_2269 ^ n_1515;
assign n_2398 = n_2270 ^ n_1514;
assign n_2399 = n_2271 ^ n_1513;
assign n_2400 = n_2272 ^ n_1251;
assign n_2401 = n_2273 ^ n_1511;
assign n_2402 = n_2274 ^ n_1382;
assign y0 = n_2275;
assign y1 = n_2276;
assign y2 = n_2277;
assign y3 = n_2278;
assign y4 = n_2279;
assign y5 = n_2280;
assign y6 = n_2281;
assign y7 = n_2282;
assign y8 = n_2283;
assign y9 = n_2284;
assign y10 = n_2285;
assign y11 = n_2286;
assign y12 = n_2287;
assign y13 = n_2288;
assign y14 = n_2289;
assign y15 = n_2290;
assign y16 = n_2291;
assign y17 = n_2292;
assign y18 = n_2293;
assign y19 = n_2294;
assign y20 = n_2295;
assign y21 = n_2296;
assign y22 = n_2297;
assign y23 = n_2298;
assign y24 = n_2299;
assign y25 = n_2300;
assign y26 = n_2301;
assign y27 = n_2302;
assign y28 = n_2303;
assign y29 = n_2304;
assign y30 = n_2305;
assign y31 = n_2306;
assign y32 = n_2307;
assign y33 = n_2308;
assign y34 = n_2309;
assign y35 = n_2310;
assign y36 = n_2311;
assign y37 = n_2312;
assign y38 = n_2313;
assign y39 = n_2314;
assign y40 = n_2315;
assign y41 = n_2316;
assign y42 = n_2317;
assign y43 = n_2318;
assign y44 = n_2319;
assign y45 = n_2320;
assign y46 = n_2321;
assign y47 = n_2322;
assign y48 = n_2323;
assign y49 = n_2324;
assign y50 = n_2325;
assign y51 = n_2326;
assign y52 = n_2327;
assign y53 = n_2328;
assign y54 = n_2329;
assign y55 = n_2330;
assign y56 = n_2331;
assign y57 = n_2332;
assign y58 = n_2333;
assign y59 = n_2334;
assign y60 = n_2335;
assign y61 = n_2336;
assign y62 = n_2337;
assign y63 = n_2338;
assign y64 = n_2339;
assign y65 = n_2340;
assign y66 = n_2341;
assign y67 = n_2342;
assign y68 = n_2343;
assign y69 = n_2344;
assign y70 = n_2345;
assign y71 = n_2346;
assign y72 = n_2347;
assign y73 = n_2348;
assign y74 = n_2349;
assign y75 = n_2350;
assign y76 = n_2351;
assign y77 = n_2352;
assign y78 = n_2353;
assign y79 = n_2354;
assign y80 = n_2355;
assign y81 = n_2356;
assign y82 = n_2357;
assign y83 = n_2358;
assign y84 = n_2359;
assign y85 = n_2360;
assign y86 = n_2361;
assign y87 = n_2362;
assign y88 = n_2363;
assign y89 = n_2364;
assign y90 = n_2365;
assign y91 = n_2366;
assign y92 = n_2367;
assign y93 = n_2368;
assign y94 = n_2369;
assign y95 = n_2370;
assign y96 = n_2371;
assign y97 = n_2372;
assign y98 = n_2373;
assign y99 = n_2374;
assign y100 = n_2375;
assign y101 = n_2376;
assign y102 = n_2377;
assign y103 = n_2378;
assign y104 = n_2379;
assign y105 = n_2380;
assign y106 = n_2381;
assign y107 = n_2382;
assign y108 = n_2383;
assign y109 = n_2384;
assign y110 = n_2385;
assign y111 = n_2386;
assign y112 = n_2387;
assign y113 = n_2388;
assign y114 = n_2389;
assign y115 = n_2390;
assign y116 = n_2391;
assign y117 = n_2392;
assign y118 = n_2393;
assign y119 = n_2394;
assign y120 = n_2395;
assign y121 = n_2396;
assign y122 = n_2397;
assign y123 = n_2398;
assign y124 = n_2399;
assign y125 = n_2400;
assign y126 = n_2401;
assign y128 = n_2402;
endmodule