module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 ;
  assign n344 = x40 ^ x32 ;
  assign n348 = x41 ^ x33 ;
  assign n349 = ~n344 & ~n348 ;
  assign n351 = x42 ^ x34 ;
  assign n357 = x43 ^ x35 ;
  assign n358 = ~n351 & ~n357 ;
  assign n359 = n349 & n358 ;
  assign n361 = x44 ^ x36 ;
  assign n365 = x45 ^ x37 ;
  assign n366 = ~n361 & ~n365 ;
  assign n368 = x46 ^ x38 ;
  assign n376 = x47 ^ x39 ;
  assign n377 = ~n368 & ~n376 ;
  assign n378 = n366 & n377 ;
  assign n379 = n359 & n378 ;
  assign n369 = x39 & ~x47 ;
  assign n370 = ~n368 & n369 ;
  assign n367 = x38 & ~x46 ;
  assign n371 = n370 ^ n367 ;
  assign n372 = n366 & n371 ;
  assign n362 = x37 & ~x45 ;
  assign n363 = ~n361 & n362 ;
  assign n360 = x36 & ~x44 ;
  assign n364 = n363 ^ n360 ;
  assign n373 = n372 ^ n364 ;
  assign n374 = n359 & n373 ;
  assign n352 = x35 & ~x43 ;
  assign n353 = ~n351 & n352 ;
  assign n350 = x34 & ~x42 ;
  assign n354 = n353 ^ n350 ;
  assign n355 = n349 & n354 ;
  assign n345 = x33 & ~x41 ;
  assign n346 = ~n344 & n345 ;
  assign n343 = x32 & ~x40 ;
  assign n347 = n346 ^ n343 ;
  assign n356 = n355 ^ n347 ;
  assign n375 = n374 ^ n356 ;
  assign n380 = n379 ^ n375 ;
  assign n382 = x40 & n380 ;
  assign n381 = x32 & ~n380 ;
  assign n383 = n382 ^ n381 ;
  assign n94 = x24 ^ x16 ;
  assign n98 = x25 ^ x17 ;
  assign n99 = ~n94 & ~n98 ;
  assign n101 = x26 ^ x18 ;
  assign n107 = x27 ^ x19 ;
  assign n108 = ~n101 & ~n107 ;
  assign n109 = n99 & n108 ;
  assign n111 = x28 ^ x20 ;
  assign n115 = x29 ^ x21 ;
  assign n116 = ~n111 & ~n115 ;
  assign n118 = x30 ^ x22 ;
  assign n126 = x31 ^ x23 ;
  assign n127 = ~n118 & ~n126 ;
  assign n128 = n116 & n127 ;
  assign n129 = n109 & n128 ;
  assign n119 = x23 & ~x31 ;
  assign n120 = ~n118 & n119 ;
  assign n117 = x22 & ~x30 ;
  assign n121 = n120 ^ n117 ;
  assign n122 = n116 & n121 ;
  assign n112 = x21 & ~x29 ;
  assign n113 = ~n111 & n112 ;
  assign n110 = x20 & ~x28 ;
  assign n114 = n113 ^ n110 ;
  assign n123 = n122 ^ n114 ;
  assign n124 = n109 & n123 ;
  assign n102 = x19 & ~x27 ;
  assign n103 = ~n101 & n102 ;
  assign n100 = x18 & ~x26 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = n99 & n104 ;
  assign n95 = x17 & ~x25 ;
  assign n96 = ~n94 & n95 ;
  assign n93 = x16 & ~x24 ;
  assign n97 = n96 ^ n93 ;
  assign n106 = n105 ^ n97 ;
  assign n125 = n124 ^ n106 ;
  assign n130 = n129 ^ n125 ;
  assign n341 = x16 & n130 ;
  assign n340 = x24 & ~n130 ;
  assign n342 = n341 ^ n340 ;
  assign n385 = n383 ^ n342 ;
  assign n390 = x41 & n380 ;
  assign n389 = x33 & ~n380 ;
  assign n391 = n390 ^ n389 ;
  assign n387 = x17 & n130 ;
  assign n386 = x25 & ~n130 ;
  assign n388 = n387 ^ n386 ;
  assign n395 = n391 ^ n388 ;
  assign n396 = ~n385 & ~n395 ;
  assign n401 = x42 & n380 ;
  assign n400 = x34 & ~n380 ;
  assign n402 = n401 ^ n400 ;
  assign n398 = x18 & n130 ;
  assign n397 = x26 & ~n130 ;
  assign n399 = n398 ^ n397 ;
  assign n404 = n402 ^ n399 ;
  assign n409 = x43 & n380 ;
  assign n408 = x35 & ~n380 ;
  assign n410 = n409 ^ n408 ;
  assign n406 = x19 & n130 ;
  assign n405 = x27 & ~n130 ;
  assign n407 = n406 ^ n405 ;
  assign n416 = n410 ^ n407 ;
  assign n417 = ~n404 & ~n416 ;
  assign n418 = n396 & n417 ;
  assign n423 = x44 & n380 ;
  assign n422 = x36 & ~n380 ;
  assign n424 = n423 ^ n422 ;
  assign n420 = x20 & n130 ;
  assign n419 = x28 & ~n130 ;
  assign n421 = n420 ^ n419 ;
  assign n426 = n424 ^ n421 ;
  assign n431 = x45 & n380 ;
  assign n430 = x37 & ~n380 ;
  assign n432 = n431 ^ n430 ;
  assign n428 = x21 & n130 ;
  assign n427 = x29 & ~n130 ;
  assign n429 = n428 ^ n427 ;
  assign n436 = n432 ^ n429 ;
  assign n437 = ~n426 & ~n436 ;
  assign n442 = x46 & n380 ;
  assign n441 = x38 & ~n380 ;
  assign n443 = n442 ^ n441 ;
  assign n439 = x22 & n130 ;
  assign n438 = x30 & ~n130 ;
  assign n440 = n439 ^ n438 ;
  assign n445 = n443 ^ n440 ;
  assign n462 = x47 & ~n356 ;
  assign n461 = x47 & ~n379 ;
  assign n463 = n462 ^ n461 ;
  assign n459 = x47 & n359 ;
  assign n460 = n373 & n459 ;
  assign n464 = n463 ^ n460 ;
  assign n456 = x39 & n356 ;
  assign n455 = x39 & ~n379 ;
  assign n457 = n456 ^ n455 ;
  assign n453 = x39 & n359 ;
  assign n454 = n373 & n453 ;
  assign n458 = n457 ^ n454 ;
  assign n465 = n464 ^ n458 ;
  assign n449 = x23 & ~n106 ;
  assign n197 = x23 & ~n129 ;
  assign n450 = n449 ^ n197 ;
  assign n199 = x23 & n109 ;
  assign n200 = n123 & n199 ;
  assign n451 = n450 ^ n200 ;
  assign n446 = x31 & n106 ;
  assign n203 = x31 & ~n129 ;
  assign n447 = n446 ^ n203 ;
  assign n205 = x31 & n109 ;
  assign n206 = n123 & n205 ;
  assign n448 = n447 ^ n206 ;
  assign n452 = n451 ^ n448 ;
  assign n473 = n465 ^ n452 ;
  assign n474 = ~n445 & ~n473 ;
  assign n475 = n437 & n474 ;
  assign n476 = n418 & n475 ;
  assign n466 = n452 & ~n465 ;
  assign n467 = ~n445 & n466 ;
  assign n444 = n440 & ~n443 ;
  assign n468 = n467 ^ n444 ;
  assign n469 = n437 & n468 ;
  assign n433 = n429 & ~n432 ;
  assign n434 = ~n426 & n433 ;
  assign n425 = n421 & ~n424 ;
  assign n435 = n434 ^ n425 ;
  assign n470 = n469 ^ n435 ;
  assign n471 = n418 & n470 ;
  assign n411 = n407 & ~n410 ;
  assign n412 = ~n404 & n411 ;
  assign n403 = n399 & ~n402 ;
  assign n413 = n412 ^ n403 ;
  assign n414 = n396 & n413 ;
  assign n392 = n388 & ~n391 ;
  assign n393 = ~n385 & n392 ;
  assign n384 = n342 & ~n383 ;
  assign n394 = n393 ^ n384 ;
  assign n415 = n414 ^ n394 ;
  assign n472 = n471 ^ n415 ;
  assign n477 = n476 ^ n472 ;
  assign n479 = n383 & n477 ;
  assign n478 = n342 & ~n477 ;
  assign n480 = n479 ^ n478 ;
  assign n50 = x8 ^ x0 ;
  assign n54 = x9 ^ x1 ;
  assign n55 = ~n50 & ~n54 ;
  assign n57 = x10 ^ x2 ;
  assign n63 = x11 ^ x3 ;
  assign n64 = ~n57 & ~n63 ;
  assign n65 = n55 & n64 ;
  assign n67 = x12 ^ x4 ;
  assign n71 = x13 ^ x5 ;
  assign n72 = ~n67 & ~n71 ;
  assign n74 = x14 ^ x6 ;
  assign n82 = x15 ^ x7 ;
  assign n83 = ~n74 & ~n82 ;
  assign n84 = n72 & n83 ;
  assign n85 = n65 & n84 ;
  assign n75 = x7 & ~x15 ;
  assign n76 = ~n74 & n75 ;
  assign n73 = x6 & ~x14 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = n72 & n77 ;
  assign n68 = x5 & ~x13 ;
  assign n69 = ~n67 & n68 ;
  assign n66 = x4 & ~x12 ;
  assign n70 = n69 ^ n66 ;
  assign n79 = n78 ^ n70 ;
  assign n80 = n65 & n79 ;
  assign n58 = x3 & ~x11 ;
  assign n59 = ~n57 & n58 ;
  assign n56 = x2 & ~x10 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n55 & n60 ;
  assign n51 = x1 & ~x9 ;
  assign n52 = ~n50 & n51 ;
  assign n49 = x0 & ~x8 ;
  assign n53 = n52 ^ n49 ;
  assign n62 = n61 ^ n53 ;
  assign n81 = n80 ^ n62 ;
  assign n86 = n85 ^ n81 ;
  assign n91 = x0 & n86 ;
  assign n90 = x8 & ~n86 ;
  assign n92 = n91 ^ n90 ;
  assign n132 = x24 & n130 ;
  assign n131 = x16 & ~n130 ;
  assign n133 = n132 ^ n131 ;
  assign n135 = n133 ^ n92 ;
  assign n140 = x1 & n86 ;
  assign n139 = x9 & ~n86 ;
  assign n141 = n140 ^ n139 ;
  assign n137 = x25 & n130 ;
  assign n136 = x17 & ~n130 ;
  assign n138 = n137 ^ n136 ;
  assign n145 = n141 ^ n138 ;
  assign n146 = ~n135 & ~n145 ;
  assign n151 = x26 & n130 ;
  assign n150 = x18 & ~n130 ;
  assign n152 = n151 ^ n150 ;
  assign n148 = x2 & n86 ;
  assign n147 = x10 & ~n86 ;
  assign n149 = n148 ^ n147 ;
  assign n154 = n152 ^ n149 ;
  assign n159 = x27 & n130 ;
  assign n158 = x19 & ~n130 ;
  assign n160 = n159 ^ n158 ;
  assign n156 = x3 & n86 ;
  assign n155 = x11 & ~n86 ;
  assign n157 = n156 ^ n155 ;
  assign n166 = n160 ^ n157 ;
  assign n167 = ~n154 & ~n166 ;
  assign n168 = n146 & n167 ;
  assign n173 = x28 & n130 ;
  assign n172 = x20 & ~n130 ;
  assign n174 = n173 ^ n172 ;
  assign n170 = x4 & n86 ;
  assign n169 = x12 & ~n86 ;
  assign n171 = n170 ^ n169 ;
  assign n176 = n174 ^ n171 ;
  assign n181 = x29 & n130 ;
  assign n180 = x21 & ~n130 ;
  assign n182 = n181 ^ n180 ;
  assign n178 = x5 & n86 ;
  assign n177 = x13 & ~n86 ;
  assign n179 = n178 ^ n177 ;
  assign n186 = n182 ^ n179 ;
  assign n187 = ~n176 & ~n186 ;
  assign n192 = x30 & n130 ;
  assign n191 = x22 & ~n130 ;
  assign n193 = n192 ^ n191 ;
  assign n189 = x6 & n86 ;
  assign n188 = x14 & ~n86 ;
  assign n190 = n189 ^ n188 ;
  assign n195 = n193 ^ n190 ;
  assign n218 = x7 & ~n62 ;
  assign n217 = x7 & ~n85 ;
  assign n219 = n218 ^ n217 ;
  assign n215 = x7 & n65 ;
  assign n216 = n79 & n215 ;
  assign n220 = n219 ^ n216 ;
  assign n212 = x15 & n62 ;
  assign n211 = x15 & ~n85 ;
  assign n213 = n212 ^ n211 ;
  assign n209 = x15 & n65 ;
  assign n210 = n79 & n209 ;
  assign n214 = n213 ^ n210 ;
  assign n221 = n220 ^ n214 ;
  assign n202 = x31 & ~n106 ;
  assign n204 = n203 ^ n202 ;
  assign n207 = n206 ^ n204 ;
  assign n196 = x23 & n106 ;
  assign n198 = n197 ^ n196 ;
  assign n201 = n200 ^ n198 ;
  assign n208 = n207 ^ n201 ;
  assign n229 = n221 ^ n208 ;
  assign n230 = ~n195 & ~n229 ;
  assign n231 = n187 & n230 ;
  assign n232 = n168 & n231 ;
  assign n222 = ~n208 & n221 ;
  assign n223 = ~n195 & n222 ;
  assign n194 = n190 & ~n193 ;
  assign n224 = n223 ^ n194 ;
  assign n225 = n187 & n224 ;
  assign n183 = n179 & ~n182 ;
  assign n184 = ~n176 & n183 ;
  assign n175 = n171 & ~n174 ;
  assign n185 = n184 ^ n175 ;
  assign n226 = n225 ^ n185 ;
  assign n227 = n168 & n226 ;
  assign n161 = n157 & ~n160 ;
  assign n162 = ~n154 & n161 ;
  assign n153 = n149 & ~n152 ;
  assign n163 = n162 ^ n153 ;
  assign n164 = n146 & n163 ;
  assign n142 = ~n138 & n141 ;
  assign n143 = ~n135 & n142 ;
  assign n134 = n92 & ~n133 ;
  assign n144 = n143 ^ n134 ;
  assign n165 = n164 ^ n144 ;
  assign n228 = n227 ^ n165 ;
  assign n233 = n232 ^ n228 ;
  assign n338 = n92 & n233 ;
  assign n337 = n133 & ~n233 ;
  assign n339 = n338 ^ n337 ;
  assign n482 = n480 ^ n339 ;
  assign n487 = n391 & n477 ;
  assign n486 = n388 & ~n477 ;
  assign n488 = n487 ^ n486 ;
  assign n484 = n141 & n233 ;
  assign n483 = n138 & ~n233 ;
  assign n485 = n484 ^ n483 ;
  assign n492 = n488 ^ n485 ;
  assign n493 = ~n482 & ~n492 ;
  assign n498 = n402 & n477 ;
  assign n497 = n399 & ~n477 ;
  assign n499 = n498 ^ n497 ;
  assign n495 = n149 & n233 ;
  assign n494 = n152 & ~n233 ;
  assign n496 = n495 ^ n494 ;
  assign n501 = n499 ^ n496 ;
  assign n506 = n410 & n477 ;
  assign n505 = n407 & ~n477 ;
  assign n507 = n506 ^ n505 ;
  assign n503 = n157 & n233 ;
  assign n502 = n160 & ~n233 ;
  assign n504 = n503 ^ n502 ;
  assign n513 = n507 ^ n504 ;
  assign n514 = ~n501 & ~n513 ;
  assign n515 = n493 & n514 ;
  assign n520 = n424 & n477 ;
  assign n519 = n421 & ~n477 ;
  assign n521 = n520 ^ n519 ;
  assign n517 = n171 & n233 ;
  assign n516 = n174 & ~n233 ;
  assign n518 = n517 ^ n516 ;
  assign n523 = n521 ^ n518 ;
  assign n528 = n432 & n477 ;
  assign n527 = n429 & ~n477 ;
  assign n529 = n528 ^ n527 ;
  assign n525 = n179 & n233 ;
  assign n524 = n182 & ~n233 ;
  assign n526 = n525 ^ n524 ;
  assign n533 = n529 ^ n526 ;
  assign n534 = ~n523 & ~n533 ;
  assign n539 = n443 & n477 ;
  assign n538 = n440 & ~n477 ;
  assign n540 = n539 ^ n538 ;
  assign n536 = n190 & n233 ;
  assign n535 = n193 & ~n233 ;
  assign n537 = n536 ^ n535 ;
  assign n542 = n540 ^ n537 ;
  assign n547 = n465 & n477 ;
  assign n546 = n452 & ~n477 ;
  assign n548 = n547 ^ n546 ;
  assign n544 = n221 & n233 ;
  assign n543 = n208 & ~n233 ;
  assign n545 = n544 ^ n543 ;
  assign n556 = n548 ^ n545 ;
  assign n557 = ~n542 & ~n556 ;
  assign n558 = n534 & n557 ;
  assign n559 = n515 & n558 ;
  assign n549 = n545 & ~n548 ;
  assign n550 = ~n542 & n549 ;
  assign n541 = n537 & ~n540 ;
  assign n551 = n550 ^ n541 ;
  assign n552 = n534 & n551 ;
  assign n530 = n526 & ~n529 ;
  assign n531 = ~n523 & n530 ;
  assign n522 = n518 & ~n521 ;
  assign n532 = n531 ^ n522 ;
  assign n553 = n552 ^ n532 ;
  assign n554 = n515 & n553 ;
  assign n508 = n504 & ~n507 ;
  assign n509 = ~n501 & n508 ;
  assign n500 = n496 & ~n499 ;
  assign n510 = n509 ^ n500 ;
  assign n511 = n493 & n510 ;
  assign n489 = n485 & ~n488 ;
  assign n490 = ~n482 & n489 ;
  assign n481 = n339 & ~n480 ;
  assign n491 = n490 ^ n481 ;
  assign n512 = n511 ^ n491 ;
  assign n555 = n554 ^ n512 ;
  assign n560 = n559 ^ n555 ;
  assign n562 = n480 & n560 ;
  assign n561 = n339 & ~n560 ;
  assign n563 = n562 ^ n561 ;
  assign n88 = x8 & n86 ;
  assign n87 = x0 & ~n86 ;
  assign n89 = n88 ^ n87 ;
  assign n235 = n133 & n233 ;
  assign n234 = n92 & ~n233 ;
  assign n236 = n235 ^ n234 ;
  assign n238 = n236 ^ n89 ;
  assign n243 = x9 & n86 ;
  assign n242 = x1 & ~n86 ;
  assign n244 = n243 ^ n242 ;
  assign n240 = n138 & n233 ;
  assign n239 = n141 & ~n233 ;
  assign n241 = n240 ^ n239 ;
  assign n248 = n244 ^ n241 ;
  assign n249 = ~n238 & ~n248 ;
  assign n254 = n152 & n233 ;
  assign n253 = n149 & ~n233 ;
  assign n255 = n254 ^ n253 ;
  assign n251 = x10 & n86 ;
  assign n250 = x2 & ~n86 ;
  assign n252 = n251 ^ n250 ;
  assign n257 = n255 ^ n252 ;
  assign n262 = n160 & n233 ;
  assign n261 = n157 & ~n233 ;
  assign n263 = n262 ^ n261 ;
  assign n259 = x11 & n86 ;
  assign n258 = x3 & ~n86 ;
  assign n260 = n259 ^ n258 ;
  assign n269 = n263 ^ n260 ;
  assign n270 = ~n257 & ~n269 ;
  assign n271 = n249 & n270 ;
  assign n276 = n174 & n233 ;
  assign n275 = n171 & ~n233 ;
  assign n277 = n276 ^ n275 ;
  assign n273 = x12 & n86 ;
  assign n272 = x4 & ~n86 ;
  assign n274 = n273 ^ n272 ;
  assign n279 = n277 ^ n274 ;
  assign n284 = n182 & n233 ;
  assign n283 = n179 & ~n233 ;
  assign n285 = n284 ^ n283 ;
  assign n281 = x13 & n86 ;
  assign n280 = x5 & ~n86 ;
  assign n282 = n281 ^ n280 ;
  assign n289 = n285 ^ n282 ;
  assign n290 = ~n279 & ~n289 ;
  assign n320 = n193 & n233 ;
  assign n319 = n190 & ~n233 ;
  assign n321 = n320 ^ n319 ;
  assign n292 = x14 & n86 ;
  assign n291 = x6 & ~n86 ;
  assign n293 = n292 ^ n291 ;
  assign n322 = n321 ^ n293 ;
  assign n324 = n208 & n233 ;
  assign n323 = n221 & ~n233 ;
  assign n325 = n324 ^ n323 ;
  assign n297 = x15 & n86 ;
  assign n296 = x7 & ~n86 ;
  assign n298 = n297 ^ n296 ;
  assign n326 = n325 ^ n298 ;
  assign n327 = ~n322 & ~n326 ;
  assign n328 = n290 & n327 ;
  assign n329 = n271 & n328 ;
  assign n311 = ~n193 & n293 ;
  assign n312 = n233 & n311 ;
  assign n301 = ~n221 & n298 ;
  assign n302 = ~n233 & n301 ;
  assign n299 = ~n208 & n298 ;
  assign n300 = n233 & n299 ;
  assign n303 = n302 ^ n300 ;
  assign n307 = ~n193 & n233 ;
  assign n308 = n303 & n307 ;
  assign n305 = ~n190 & ~n233 ;
  assign n306 = n303 & n305 ;
  assign n309 = n308 ^ n306 ;
  assign n304 = n293 & n303 ;
  assign n310 = n309 ^ n304 ;
  assign n313 = n312 ^ n310 ;
  assign n294 = ~n190 & n293 ;
  assign n295 = ~n233 & n294 ;
  assign n314 = n313 ^ n295 ;
  assign n315 = n290 & n314 ;
  assign n286 = n282 & ~n285 ;
  assign n287 = ~n279 & n286 ;
  assign n278 = n274 & ~n277 ;
  assign n288 = n287 ^ n278 ;
  assign n316 = n315 ^ n288 ;
  assign n317 = n271 & n316 ;
  assign n264 = n260 & ~n263 ;
  assign n265 = ~n257 & n264 ;
  assign n256 = n252 & ~n255 ;
  assign n266 = n265 ^ n256 ;
  assign n267 = n249 & n266 ;
  assign n245 = ~n241 & n244 ;
  assign n246 = ~n238 & n245 ;
  assign n237 = n89 & ~n236 ;
  assign n247 = n246 ^ n237 ;
  assign n268 = n267 ^ n247 ;
  assign n318 = n317 ^ n268 ;
  assign n330 = n329 ^ n318 ;
  assign n335 = n89 & n330 ;
  assign n334 = n236 & ~n330 ;
  assign n336 = n335 ^ n334 ;
  assign n565 = n563 ^ n336 ;
  assign n570 = n488 & n560 ;
  assign n569 = n485 & ~n560 ;
  assign n571 = n570 ^ n569 ;
  assign n567 = n244 & n330 ;
  assign n566 = n241 & ~n330 ;
  assign n568 = n567 ^ n566 ;
  assign n575 = n571 ^ n568 ;
  assign n576 = ~n565 & ~n575 ;
  assign n581 = n499 & n560 ;
  assign n580 = n496 & ~n560 ;
  assign n582 = n581 ^ n580 ;
  assign n578 = n252 & n330 ;
  assign n577 = n255 & ~n330 ;
  assign n579 = n578 ^ n577 ;
  assign n584 = n582 ^ n579 ;
  assign n589 = n507 & n560 ;
  assign n588 = n504 & ~n560 ;
  assign n590 = n589 ^ n588 ;
  assign n586 = n260 & n330 ;
  assign n585 = n263 & ~n330 ;
  assign n587 = n586 ^ n585 ;
  assign n596 = n590 ^ n587 ;
  assign n597 = ~n584 & ~n596 ;
  assign n598 = n576 & n597 ;
  assign n603 = n521 & n560 ;
  assign n602 = n518 & ~n560 ;
  assign n604 = n603 ^ n602 ;
  assign n600 = n274 & n330 ;
  assign n599 = n277 & ~n330 ;
  assign n601 = n600 ^ n599 ;
  assign n606 = n604 ^ n601 ;
  assign n611 = n529 & n560 ;
  assign n610 = n526 & ~n560 ;
  assign n612 = n611 ^ n610 ;
  assign n608 = n282 & n330 ;
  assign n607 = n285 & ~n330 ;
  assign n609 = n608 ^ n607 ;
  assign n616 = n612 ^ n609 ;
  assign n617 = ~n606 & ~n616 ;
  assign n622 = n540 & n560 ;
  assign n621 = n537 & ~n560 ;
  assign n623 = n622 ^ n621 ;
  assign n619 = n293 & n330 ;
  assign n618 = n321 & ~n330 ;
  assign n620 = n619 ^ n618 ;
  assign n625 = n623 ^ n620 ;
  assign n630 = n548 & n560 ;
  assign n629 = n545 & ~n560 ;
  assign n631 = n630 ^ n629 ;
  assign n627 = n298 & n330 ;
  assign n626 = n325 & ~n330 ;
  assign n628 = n627 ^ n626 ;
  assign n639 = n631 ^ n628 ;
  assign n640 = ~n625 & ~n639 ;
  assign n641 = n617 & n640 ;
  assign n642 = n598 & n641 ;
  assign n632 = n628 & ~n631 ;
  assign n633 = ~n625 & n632 ;
  assign n624 = n620 & ~n623 ;
  assign n634 = n633 ^ n624 ;
  assign n635 = n617 & n634 ;
  assign n613 = n609 & ~n612 ;
  assign n614 = ~n606 & n613 ;
  assign n605 = n601 & ~n604 ;
  assign n615 = n614 ^ n605 ;
  assign n636 = n635 ^ n615 ;
  assign n637 = n598 & n636 ;
  assign n591 = n587 & ~n590 ;
  assign n592 = ~n584 & n591 ;
  assign n583 = n579 & ~n582 ;
  assign n593 = n592 ^ n583 ;
  assign n594 = n576 & n593 ;
  assign n572 = n568 & ~n571 ;
  assign n573 = ~n565 & n572 ;
  assign n564 = n336 & ~n563 ;
  assign n574 = n573 ^ n564 ;
  assign n595 = n594 ^ n574 ;
  assign n638 = n637 ^ n595 ;
  assign n643 = n642 ^ n638 ;
  assign n645 = n563 & n643 ;
  assign n644 = n336 & ~n643 ;
  assign n646 = n645 ^ n644 ;
  assign n332 = n236 & n330 ;
  assign n331 = n89 & ~n330 ;
  assign n333 = n332 ^ n331 ;
  assign n648 = n646 ^ n333 ;
  assign n653 = n571 & n643 ;
  assign n652 = n568 & ~n643 ;
  assign n654 = n653 ^ n652 ;
  assign n650 = n241 & n330 ;
  assign n649 = n244 & ~n330 ;
  assign n651 = n650 ^ n649 ;
  assign n658 = n654 ^ n651 ;
  assign n659 = ~n648 & ~n658 ;
  assign n664 = n582 & n643 ;
  assign n663 = n579 & ~n643 ;
  assign n665 = n664 ^ n663 ;
  assign n661 = n255 & n330 ;
  assign n660 = n252 & ~n330 ;
  assign n662 = n661 ^ n660 ;
  assign n667 = n665 ^ n662 ;
  assign n672 = n590 & n643 ;
  assign n671 = n587 & ~n643 ;
  assign n673 = n672 ^ n671 ;
  assign n669 = n263 & n330 ;
  assign n668 = n260 & ~n330 ;
  assign n670 = n669 ^ n668 ;
  assign n679 = n673 ^ n670 ;
  assign n680 = ~n667 & ~n679 ;
  assign n681 = n659 & n680 ;
  assign n686 = n604 & n643 ;
  assign n685 = n601 & ~n643 ;
  assign n687 = n686 ^ n685 ;
  assign n683 = n277 & n330 ;
  assign n682 = n274 & ~n330 ;
  assign n684 = n683 ^ n682 ;
  assign n689 = n687 ^ n684 ;
  assign n694 = n612 & n643 ;
  assign n693 = n609 & ~n643 ;
  assign n695 = n694 ^ n693 ;
  assign n691 = n285 & n330 ;
  assign n690 = n282 & ~n330 ;
  assign n692 = n691 ^ n690 ;
  assign n699 = n695 ^ n692 ;
  assign n700 = ~n689 & ~n699 ;
  assign n730 = n623 & n643 ;
  assign n729 = n620 & ~n643 ;
  assign n731 = n730 ^ n729 ;
  assign n702 = n321 & n330 ;
  assign n701 = n293 & ~n330 ;
  assign n703 = n702 ^ n701 ;
  assign n732 = n731 ^ n703 ;
  assign n734 = n631 & n643 ;
  assign n733 = n628 & ~n643 ;
  assign n735 = n734 ^ n733 ;
  assign n707 = n325 & n330 ;
  assign n706 = n298 & ~n330 ;
  assign n708 = n707 ^ n706 ;
  assign n736 = n735 ^ n708 ;
  assign n737 = ~n732 & ~n736 ;
  assign n738 = n700 & n737 ;
  assign n739 = n681 & n738 ;
  assign n721 = ~n623 & n703 ;
  assign n722 = n643 & n721 ;
  assign n711 = ~n631 & n708 ;
  assign n712 = n643 & n711 ;
  assign n709 = ~n628 & n708 ;
  assign n710 = ~n643 & n709 ;
  assign n713 = n712 ^ n710 ;
  assign n717 = ~n623 & n643 ;
  assign n718 = n713 & n717 ;
  assign n715 = ~n620 & ~n643 ;
  assign n716 = n713 & n715 ;
  assign n719 = n718 ^ n716 ;
  assign n714 = n703 & n713 ;
  assign n720 = n719 ^ n714 ;
  assign n723 = n722 ^ n720 ;
  assign n704 = ~n620 & n703 ;
  assign n705 = ~n643 & n704 ;
  assign n724 = n723 ^ n705 ;
  assign n725 = n700 & n724 ;
  assign n696 = n692 & ~n695 ;
  assign n697 = ~n689 & n696 ;
  assign n688 = n684 & ~n687 ;
  assign n698 = n697 ^ n688 ;
  assign n726 = n725 ^ n698 ;
  assign n727 = n681 & n726 ;
  assign n674 = n670 & ~n673 ;
  assign n675 = ~n667 & n674 ;
  assign n666 = n662 & ~n665 ;
  assign n676 = n675 ^ n666 ;
  assign n677 = n659 & n676 ;
  assign n655 = n651 & ~n654 ;
  assign n656 = ~n648 & n655 ;
  assign n647 = n333 & ~n646 ;
  assign n657 = n656 ^ n647 ;
  assign n678 = n677 ^ n657 ;
  assign n728 = n727 ^ n678 ;
  assign n740 = n739 ^ n728 ;
  assign n742 = n646 & n740 ;
  assign n741 = n333 & ~n740 ;
  assign n743 = n742 ^ n741 ;
  assign n745 = n654 & n740 ;
  assign n744 = n651 & ~n740 ;
  assign n746 = n745 ^ n744 ;
  assign n748 = n665 & n740 ;
  assign n747 = n662 & ~n740 ;
  assign n749 = n748 ^ n747 ;
  assign n751 = n673 & n740 ;
  assign n750 = n670 & ~n740 ;
  assign n752 = n751 ^ n750 ;
  assign n754 = n687 & n740 ;
  assign n753 = n684 & ~n740 ;
  assign n755 = n754 ^ n753 ;
  assign n757 = n695 & n740 ;
  assign n756 = n692 & ~n740 ;
  assign n758 = n757 ^ n756 ;
  assign n760 = n731 & n740 ;
  assign n759 = n703 & ~n740 ;
  assign n761 = n760 ^ n759 ;
  assign n763 = n735 & n740 ;
  assign n762 = n708 & ~n740 ;
  assign n764 = n763 ^ n762 ;
  assign n766 = n333 & n740 ;
  assign n765 = n646 & ~n740 ;
  assign n767 = n766 ^ n765 ;
  assign n769 = n651 & n740 ;
  assign n768 = n654 & ~n740 ;
  assign n770 = n769 ^ n768 ;
  assign n772 = n662 & n740 ;
  assign n771 = n665 & ~n740 ;
  assign n773 = n772 ^ n771 ;
  assign n775 = n670 & n740 ;
  assign n774 = n673 & ~n740 ;
  assign n776 = n775 ^ n774 ;
  assign n778 = n684 & n740 ;
  assign n777 = n687 & ~n740 ;
  assign n779 = n778 ^ n777 ;
  assign n781 = n692 & n740 ;
  assign n780 = n695 & ~n740 ;
  assign n782 = n781 ^ n780 ;
  assign n784 = n703 & n740 ;
  assign n783 = n731 & ~n740 ;
  assign n785 = n784 ^ n783 ;
  assign n787 = n708 & n740 ;
  assign n786 = n735 & ~n740 ;
  assign n788 = n787 ^ n786 ;
  assign n799 = x32 & n380 ;
  assign n798 = x40 & ~n380 ;
  assign n800 = n799 ^ n798 ;
  assign n796 = n342 & n477 ;
  assign n795 = n383 & ~n477 ;
  assign n797 = n796 ^ n795 ;
  assign n802 = n800 ^ n797 ;
  assign n807 = x33 & n380 ;
  assign n806 = x41 & ~n380 ;
  assign n808 = n807 ^ n806 ;
  assign n804 = n388 & n477 ;
  assign n803 = n391 & ~n477 ;
  assign n805 = n804 ^ n803 ;
  assign n812 = n808 ^ n805 ;
  assign n813 = ~n802 & ~n812 ;
  assign n818 = x34 & n380 ;
  assign n817 = x42 & ~n380 ;
  assign n819 = n818 ^ n817 ;
  assign n815 = n399 & n477 ;
  assign n814 = n402 & ~n477 ;
  assign n816 = n815 ^ n814 ;
  assign n821 = n819 ^ n816 ;
  assign n826 = x35 & n380 ;
  assign n825 = x43 & ~n380 ;
  assign n827 = n826 ^ n825 ;
  assign n823 = n407 & n477 ;
  assign n822 = n410 & ~n477 ;
  assign n824 = n823 ^ n822 ;
  assign n833 = n827 ^ n824 ;
  assign n834 = ~n821 & ~n833 ;
  assign n835 = n813 & n834 ;
  assign n840 = x36 & n380 ;
  assign n839 = x44 & ~n380 ;
  assign n841 = n840 ^ n839 ;
  assign n837 = n421 & n477 ;
  assign n836 = n424 & ~n477 ;
  assign n838 = n837 ^ n836 ;
  assign n843 = n841 ^ n838 ;
  assign n848 = x37 & n380 ;
  assign n847 = x45 & ~n380 ;
  assign n849 = n848 ^ n847 ;
  assign n845 = n429 & n477 ;
  assign n844 = n432 & ~n477 ;
  assign n846 = n845 ^ n844 ;
  assign n853 = n849 ^ n846 ;
  assign n854 = ~n843 & ~n853 ;
  assign n859 = x38 & n380 ;
  assign n858 = x46 & ~n380 ;
  assign n860 = n859 ^ n858 ;
  assign n856 = n440 & n477 ;
  assign n855 = n443 & ~n477 ;
  assign n857 = n856 ^ n855 ;
  assign n880 = n860 ^ n857 ;
  assign n882 = n452 & n477 ;
  assign n881 = n465 & ~n477 ;
  assign n883 = n882 ^ n881 ;
  assign n863 = x39 & n380 ;
  assign n862 = x47 & ~n380 ;
  assign n864 = n863 ^ n862 ;
  assign n884 = n883 ^ n864 ;
  assign n885 = ~n880 & ~n884 ;
  assign n886 = n854 & n885 ;
  assign n887 = n835 & n886 ;
  assign n867 = n465 & ~n864 ;
  assign n868 = ~n477 & n867 ;
  assign n865 = n452 & ~n864 ;
  assign n866 = n477 & n865 ;
  assign n869 = n868 ^ n866 ;
  assign n872 = n856 & n869 ;
  assign n871 = n855 & n869 ;
  assign n873 = n872 ^ n871 ;
  assign n870 = ~n860 & n869 ;
  assign n874 = n873 ^ n870 ;
  assign n861 = n857 & ~n860 ;
  assign n875 = n874 ^ n861 ;
  assign n876 = n854 & n875 ;
  assign n850 = n846 & ~n849 ;
  assign n851 = ~n843 & n850 ;
  assign n842 = n838 & ~n841 ;
  assign n852 = n851 ^ n842 ;
  assign n877 = n876 ^ n852 ;
  assign n878 = n835 & n877 ;
  assign n828 = n824 & ~n827 ;
  assign n829 = ~n821 & n828 ;
  assign n820 = n816 & ~n819 ;
  assign n830 = n829 ^ n820 ;
  assign n831 = n813 & n830 ;
  assign n809 = n805 & ~n808 ;
  assign n810 = ~n802 & n809 ;
  assign n801 = n797 & ~n800 ;
  assign n811 = n810 ^ n801 ;
  assign n832 = n831 ^ n811 ;
  assign n879 = n878 ^ n832 ;
  assign n888 = n887 ^ n879 ;
  assign n890 = n800 & n888 ;
  assign n889 = n797 & ~n888 ;
  assign n891 = n890 ^ n889 ;
  assign n793 = n339 & n560 ;
  assign n792 = n480 & ~n560 ;
  assign n794 = n793 ^ n792 ;
  assign n893 = n891 ^ n794 ;
  assign n898 = n808 & n888 ;
  assign n897 = n805 & ~n888 ;
  assign n899 = n898 ^ n897 ;
  assign n895 = n485 & n560 ;
  assign n894 = n488 & ~n560 ;
  assign n896 = n895 ^ n894 ;
  assign n903 = n899 ^ n896 ;
  assign n904 = ~n893 & ~n903 ;
  assign n909 = n819 & n888 ;
  assign n908 = n816 & ~n888 ;
  assign n910 = n909 ^ n908 ;
  assign n906 = n496 & n560 ;
  assign n905 = n499 & ~n560 ;
  assign n907 = n906 ^ n905 ;
  assign n912 = n910 ^ n907 ;
  assign n917 = n827 & n888 ;
  assign n916 = n824 & ~n888 ;
  assign n918 = n917 ^ n916 ;
  assign n914 = n504 & n560 ;
  assign n913 = n507 & ~n560 ;
  assign n915 = n914 ^ n913 ;
  assign n924 = n918 ^ n915 ;
  assign n925 = ~n912 & ~n924 ;
  assign n926 = n904 & n925 ;
  assign n931 = n841 & n888 ;
  assign n930 = n838 & ~n888 ;
  assign n932 = n931 ^ n930 ;
  assign n928 = n518 & n560 ;
  assign n927 = n521 & ~n560 ;
  assign n929 = n928 ^ n927 ;
  assign n934 = n932 ^ n929 ;
  assign n939 = n849 & n888 ;
  assign n938 = n846 & ~n888 ;
  assign n940 = n939 ^ n938 ;
  assign n936 = n526 & n560 ;
  assign n935 = n529 & ~n560 ;
  assign n937 = n936 ^ n935 ;
  assign n944 = n940 ^ n937 ;
  assign n945 = ~n934 & ~n944 ;
  assign n950 = n860 & n888 ;
  assign n949 = n857 & ~n888 ;
  assign n951 = n950 ^ n949 ;
  assign n947 = n537 & n560 ;
  assign n946 = n540 & ~n560 ;
  assign n948 = n947 ^ n946 ;
  assign n953 = n951 ^ n948 ;
  assign n958 = n864 & n888 ;
  assign n957 = n883 & ~n888 ;
  assign n959 = n958 ^ n957 ;
  assign n955 = n545 & n560 ;
  assign n954 = n548 & ~n560 ;
  assign n956 = n955 ^ n954 ;
  assign n967 = n959 ^ n956 ;
  assign n968 = ~n953 & ~n967 ;
  assign n969 = n945 & n968 ;
  assign n970 = n926 & n969 ;
  assign n960 = n956 & ~n959 ;
  assign n961 = ~n953 & n960 ;
  assign n952 = n948 & ~n951 ;
  assign n962 = n961 ^ n952 ;
  assign n963 = n945 & n962 ;
  assign n941 = n937 & ~n940 ;
  assign n942 = ~n934 & n941 ;
  assign n933 = n929 & ~n932 ;
  assign n943 = n942 ^ n933 ;
  assign n964 = n963 ^ n943 ;
  assign n965 = n926 & n964 ;
  assign n919 = n915 & ~n918 ;
  assign n920 = ~n912 & n919 ;
  assign n911 = n907 & ~n910 ;
  assign n921 = n920 ^ n911 ;
  assign n922 = n904 & n921 ;
  assign n900 = n896 & ~n899 ;
  assign n901 = ~n893 & n900 ;
  assign n892 = n794 & ~n891 ;
  assign n902 = n901 ^ n892 ;
  assign n923 = n922 ^ n902 ;
  assign n966 = n965 ^ n923 ;
  assign n971 = n970 ^ n966 ;
  assign n973 = n891 & n971 ;
  assign n972 = n794 & ~n971 ;
  assign n974 = n973 ^ n972 ;
  assign n790 = n336 & n643 ;
  assign n789 = n563 & ~n643 ;
  assign n791 = n790 ^ n789 ;
  assign n976 = n974 ^ n791 ;
  assign n981 = n899 & n971 ;
  assign n980 = n896 & ~n971 ;
  assign n982 = n981 ^ n980 ;
  assign n978 = n568 & n643 ;
  assign n977 = n571 & ~n643 ;
  assign n979 = n978 ^ n977 ;
  assign n986 = n982 ^ n979 ;
  assign n987 = ~n976 & ~n986 ;
  assign n992 = n910 & n971 ;
  assign n991 = n907 & ~n971 ;
  assign n993 = n992 ^ n991 ;
  assign n989 = n579 & n643 ;
  assign n988 = n582 & ~n643 ;
  assign n990 = n989 ^ n988 ;
  assign n995 = n993 ^ n990 ;
  assign n1000 = n918 & n971 ;
  assign n999 = n915 & ~n971 ;
  assign n1001 = n1000 ^ n999 ;
  assign n997 = n587 & n643 ;
  assign n996 = n590 & ~n643 ;
  assign n998 = n997 ^ n996 ;
  assign n1007 = n1001 ^ n998 ;
  assign n1008 = ~n995 & ~n1007 ;
  assign n1009 = n987 & n1008 ;
  assign n1014 = n932 & n971 ;
  assign n1013 = n929 & ~n971 ;
  assign n1015 = n1014 ^ n1013 ;
  assign n1011 = n601 & n643 ;
  assign n1010 = n604 & ~n643 ;
  assign n1012 = n1011 ^ n1010 ;
  assign n1017 = n1015 ^ n1012 ;
  assign n1022 = n940 & n971 ;
  assign n1021 = n937 & ~n971 ;
  assign n1023 = n1022 ^ n1021 ;
  assign n1019 = n609 & n643 ;
  assign n1018 = n612 & ~n643 ;
  assign n1020 = n1019 ^ n1018 ;
  assign n1027 = n1023 ^ n1020 ;
  assign n1028 = ~n1017 & ~n1027 ;
  assign n1033 = n951 & n971 ;
  assign n1032 = n948 & ~n971 ;
  assign n1034 = n1033 ^ n1032 ;
  assign n1030 = n620 & n643 ;
  assign n1029 = n623 & ~n643 ;
  assign n1031 = n1030 ^ n1029 ;
  assign n1036 = n1034 ^ n1031 ;
  assign n1041 = n959 & n971 ;
  assign n1040 = n956 & ~n971 ;
  assign n1042 = n1041 ^ n1040 ;
  assign n1038 = n628 & n643 ;
  assign n1037 = n631 & ~n643 ;
  assign n1039 = n1038 ^ n1037 ;
  assign n1050 = n1042 ^ n1039 ;
  assign n1051 = ~n1036 & ~n1050 ;
  assign n1052 = n1028 & n1051 ;
  assign n1053 = n1009 & n1052 ;
  assign n1043 = n1039 & ~n1042 ;
  assign n1044 = ~n1036 & n1043 ;
  assign n1035 = n1031 & ~n1034 ;
  assign n1045 = n1044 ^ n1035 ;
  assign n1046 = n1028 & n1045 ;
  assign n1024 = n1020 & ~n1023 ;
  assign n1025 = ~n1017 & n1024 ;
  assign n1016 = n1012 & ~n1015 ;
  assign n1026 = n1025 ^ n1016 ;
  assign n1047 = n1046 ^ n1026 ;
  assign n1048 = n1009 & n1047 ;
  assign n1002 = n998 & ~n1001 ;
  assign n1003 = ~n995 & n1002 ;
  assign n994 = n990 & ~n993 ;
  assign n1004 = n1003 ^ n994 ;
  assign n1005 = n987 & n1004 ;
  assign n983 = n979 & ~n982 ;
  assign n984 = ~n976 & n983 ;
  assign n975 = n791 & ~n974 ;
  assign n985 = n984 ^ n975 ;
  assign n1006 = n1005 ^ n985 ;
  assign n1049 = n1048 ^ n1006 ;
  assign n1054 = n1053 ^ n1049 ;
  assign n1056 = n974 & n1054 ;
  assign n1055 = n791 & ~n1054 ;
  assign n1057 = n1056 ^ n1055 ;
  assign n1059 = n982 & n1054 ;
  assign n1058 = n979 & ~n1054 ;
  assign n1060 = n1059 ^ n1058 ;
  assign n1062 = n993 & n1054 ;
  assign n1061 = n990 & ~n1054 ;
  assign n1063 = n1062 ^ n1061 ;
  assign n1065 = n1001 & n1054 ;
  assign n1064 = n998 & ~n1054 ;
  assign n1066 = n1065 ^ n1064 ;
  assign n1068 = n1015 & n1054 ;
  assign n1067 = n1012 & ~n1054 ;
  assign n1069 = n1068 ^ n1067 ;
  assign n1071 = n1023 & n1054 ;
  assign n1070 = n1020 & ~n1054 ;
  assign n1072 = n1071 ^ n1070 ;
  assign n1074 = n1034 & n1054 ;
  assign n1073 = n1031 & ~n1054 ;
  assign n1075 = n1074 ^ n1073 ;
  assign n1077 = n1042 & n1054 ;
  assign n1076 = n1039 & ~n1054 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1080 = n791 & n1054 ;
  assign n1079 = n974 & ~n1054 ;
  assign n1081 = n1080 ^ n1079 ;
  assign n1083 = n979 & n1054 ;
  assign n1082 = n982 & ~n1054 ;
  assign n1084 = n1083 ^ n1082 ;
  assign n1086 = n990 & n1054 ;
  assign n1085 = n993 & ~n1054 ;
  assign n1087 = n1086 ^ n1085 ;
  assign n1089 = n998 & n1054 ;
  assign n1088 = n1001 & ~n1054 ;
  assign n1090 = n1089 ^ n1088 ;
  assign n1092 = n1012 & n1054 ;
  assign n1091 = n1015 & ~n1054 ;
  assign n1093 = n1092 ^ n1091 ;
  assign n1095 = n1020 & n1054 ;
  assign n1094 = n1023 & ~n1054 ;
  assign n1096 = n1095 ^ n1094 ;
  assign n1098 = n1031 & n1054 ;
  assign n1097 = n1034 & ~n1054 ;
  assign n1099 = n1098 ^ n1097 ;
  assign n1101 = n1039 & n1054 ;
  assign n1100 = n1042 & ~n1054 ;
  assign n1102 = n1101 ^ n1100 ;
  assign n1107 = n797 & n888 ;
  assign n1106 = n800 & ~n888 ;
  assign n1108 = n1107 ^ n1106 ;
  assign n1104 = n794 & n971 ;
  assign n1103 = n891 & ~n971 ;
  assign n1105 = n1104 ^ n1103 ;
  assign n1110 = n1108 ^ n1105 ;
  assign n1115 = n805 & n888 ;
  assign n1114 = n808 & ~n888 ;
  assign n1116 = n1115 ^ n1114 ;
  assign n1112 = n896 & n971 ;
  assign n1111 = n899 & ~n971 ;
  assign n1113 = n1112 ^ n1111 ;
  assign n1120 = n1116 ^ n1113 ;
  assign n1121 = ~n1110 & ~n1120 ;
  assign n1126 = n816 & n888 ;
  assign n1125 = n819 & ~n888 ;
  assign n1127 = n1126 ^ n1125 ;
  assign n1123 = n907 & n971 ;
  assign n1122 = n910 & ~n971 ;
  assign n1124 = n1123 ^ n1122 ;
  assign n1129 = n1127 ^ n1124 ;
  assign n1134 = n824 & n888 ;
  assign n1133 = n827 & ~n888 ;
  assign n1135 = n1134 ^ n1133 ;
  assign n1131 = n915 & n971 ;
  assign n1130 = n918 & ~n971 ;
  assign n1132 = n1131 ^ n1130 ;
  assign n1141 = n1135 ^ n1132 ;
  assign n1142 = ~n1129 & ~n1141 ;
  assign n1143 = n1121 & n1142 ;
  assign n1148 = n838 & n888 ;
  assign n1147 = n841 & ~n888 ;
  assign n1149 = n1148 ^ n1147 ;
  assign n1145 = n929 & n971 ;
  assign n1144 = n932 & ~n971 ;
  assign n1146 = n1145 ^ n1144 ;
  assign n1151 = n1149 ^ n1146 ;
  assign n1156 = n846 & n888 ;
  assign n1155 = n849 & ~n888 ;
  assign n1157 = n1156 ^ n1155 ;
  assign n1153 = n937 & n971 ;
  assign n1152 = n940 & ~n971 ;
  assign n1154 = n1153 ^ n1152 ;
  assign n1161 = n1157 ^ n1154 ;
  assign n1162 = ~n1151 & ~n1161 ;
  assign n1167 = n857 & n888 ;
  assign n1166 = n860 & ~n888 ;
  assign n1168 = n1167 ^ n1166 ;
  assign n1164 = n948 & n971 ;
  assign n1163 = n951 & ~n971 ;
  assign n1165 = n1164 ^ n1163 ;
  assign n1188 = n1168 ^ n1165 ;
  assign n1190 = n956 & n971 ;
  assign n1189 = n959 & ~n971 ;
  assign n1191 = n1190 ^ n1189 ;
  assign n1171 = n883 & n888 ;
  assign n1170 = n864 & ~n888 ;
  assign n1172 = n1171 ^ n1170 ;
  assign n1192 = n1191 ^ n1172 ;
  assign n1193 = ~n1188 & ~n1192 ;
  assign n1194 = n1162 & n1193 ;
  assign n1195 = n1143 & n1194 ;
  assign n1175 = n959 & ~n1172 ;
  assign n1176 = ~n971 & n1175 ;
  assign n1173 = n956 & ~n1172 ;
  assign n1174 = n971 & n1173 ;
  assign n1177 = n1176 ^ n1174 ;
  assign n1180 = n1164 & n1177 ;
  assign n1179 = n1163 & n1177 ;
  assign n1181 = n1180 ^ n1179 ;
  assign n1178 = ~n1168 & n1177 ;
  assign n1182 = n1181 ^ n1178 ;
  assign n1169 = n1165 & ~n1168 ;
  assign n1183 = n1182 ^ n1169 ;
  assign n1184 = n1162 & n1183 ;
  assign n1158 = n1154 & ~n1157 ;
  assign n1159 = ~n1151 & n1158 ;
  assign n1150 = n1146 & ~n1149 ;
  assign n1160 = n1159 ^ n1150 ;
  assign n1185 = n1184 ^ n1160 ;
  assign n1186 = n1143 & n1185 ;
  assign n1136 = n1132 & ~n1135 ;
  assign n1137 = ~n1129 & n1136 ;
  assign n1128 = n1124 & ~n1127 ;
  assign n1138 = n1137 ^ n1128 ;
  assign n1139 = n1121 & n1138 ;
  assign n1117 = n1113 & ~n1116 ;
  assign n1118 = ~n1110 & n1117 ;
  assign n1109 = n1105 & ~n1108 ;
  assign n1119 = n1118 ^ n1109 ;
  assign n1140 = n1139 ^ n1119 ;
  assign n1187 = n1186 ^ n1140 ;
  assign n1196 = n1195 ^ n1187 ;
  assign n1198 = n1108 & n1196 ;
  assign n1197 = n1105 & ~n1196 ;
  assign n1199 = n1198 ^ n1197 ;
  assign n1201 = n1116 & n1196 ;
  assign n1200 = n1113 & ~n1196 ;
  assign n1202 = n1201 ^ n1200 ;
  assign n1204 = n1127 & n1196 ;
  assign n1203 = n1124 & ~n1196 ;
  assign n1205 = n1204 ^ n1203 ;
  assign n1207 = n1135 & n1196 ;
  assign n1206 = n1132 & ~n1196 ;
  assign n1208 = n1207 ^ n1206 ;
  assign n1210 = n1149 & n1196 ;
  assign n1209 = n1146 & ~n1196 ;
  assign n1211 = n1210 ^ n1209 ;
  assign n1213 = n1157 & n1196 ;
  assign n1212 = n1154 & ~n1196 ;
  assign n1214 = n1213 ^ n1212 ;
  assign n1216 = n1168 & n1196 ;
  assign n1215 = n1165 & ~n1196 ;
  assign n1217 = n1216 ^ n1215 ;
  assign n1219 = n1172 & n1196 ;
  assign n1218 = n1191 & ~n1196 ;
  assign n1220 = n1219 ^ n1218 ;
  assign n1222 = n1105 & n1196 ;
  assign n1221 = n1108 & ~n1196 ;
  assign n1223 = n1222 ^ n1221 ;
  assign n1225 = n1113 & n1196 ;
  assign n1224 = n1116 & ~n1196 ;
  assign n1226 = n1225 ^ n1224 ;
  assign n1228 = n1124 & n1196 ;
  assign n1227 = n1127 & ~n1196 ;
  assign n1229 = n1228 ^ n1227 ;
  assign n1231 = n1132 & n1196 ;
  assign n1230 = n1135 & ~n1196 ;
  assign n1232 = n1231 ^ n1230 ;
  assign n1234 = n1146 & n1196 ;
  assign n1233 = n1149 & ~n1196 ;
  assign n1235 = n1234 ^ n1233 ;
  assign n1237 = n1154 & n1196 ;
  assign n1236 = n1157 & ~n1196 ;
  assign n1238 = n1237 ^ n1236 ;
  assign n1240 = n1165 & n1196 ;
  assign n1239 = n1168 & ~n1196 ;
  assign n1241 = n1240 ^ n1239 ;
  assign n1243 = n1191 & n1196 ;
  assign n1242 = n1172 & ~n1196 ;
  assign n1244 = n1243 ^ n1242 ;
  assign y0 = n743 ;
  assign y1 = n746 ;
  assign y2 = n749 ;
  assign y3 = n752 ;
  assign y4 = n755 ;
  assign y5 = n758 ;
  assign y6 = n761 ;
  assign y7 = n764 ;
  assign y8 = n767 ;
  assign y9 = n770 ;
  assign y10 = n773 ;
  assign y11 = n776 ;
  assign y12 = n779 ;
  assign y13 = n782 ;
  assign y14 = n785 ;
  assign y15 = n788 ;
  assign y16 = n1057 ;
  assign y17 = n1060 ;
  assign y18 = n1063 ;
  assign y19 = n1066 ;
  assign y20 = n1069 ;
  assign y21 = n1072 ;
  assign y22 = n1075 ;
  assign y23 = n1078 ;
  assign y24 = n1081 ;
  assign y25 = n1084 ;
  assign y26 = n1087 ;
  assign y27 = n1090 ;
  assign y28 = n1093 ;
  assign y29 = n1096 ;
  assign y30 = n1099 ;
  assign y31 = n1102 ;
  assign y32 = n1199 ;
  assign y33 = n1202 ;
  assign y34 = n1205 ;
  assign y35 = n1208 ;
  assign y36 = n1211 ;
  assign y37 = n1214 ;
  assign y38 = n1217 ;
  assign y39 = n1220 ;
  assign y40 = n1223 ;
  assign y41 = n1226 ;
  assign y42 = n1229 ;
  assign y43 = n1232 ;
  assign y44 = n1235 ;
  assign y45 = n1238 ;
  assign y46 = n1241 ;
  assign y47 = n1244 ;
endmodule
