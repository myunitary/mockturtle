module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 ;
  assign n185 = x132 & x133 ;
  assign n148 = ~x130 & ~x131 ;
  assign n386 = x80 & ~x128 ;
  assign n385 = x79 & x128 ;
  assign n387 = n386 ^ n385 ;
  assign n388 = ~x129 & n387 ;
  assign n382 = x78 & ~x128 ;
  assign n381 = x77 & x128 ;
  assign n383 = n382 ^ n381 ;
  assign n384 = x129 & n383 ;
  assign n389 = n388 ^ n384 ;
  assign n390 = n148 & n389 ;
  assign n137 = x130 & ~x131 ;
  assign n376 = x76 & ~x128 ;
  assign n375 = x75 & x128 ;
  assign n377 = n376 ^ n375 ;
  assign n378 = ~x129 & n377 ;
  assign n372 = x74 & ~x128 ;
  assign n371 = x73 & x128 ;
  assign n373 = n372 ^ n371 ;
  assign n374 = x129 & n373 ;
  assign n379 = n378 ^ n374 ;
  assign n380 = n137 & n379 ;
  assign n391 = n390 ^ n380 ;
  assign n171 = x130 & x131 ;
  assign n407 = x68 & ~x128 ;
  assign n406 = x67 & x128 ;
  assign n408 = n407 ^ n406 ;
  assign n409 = ~x129 & n408 ;
  assign n403 = x66 & ~x128 ;
  assign n402 = x65 & x128 ;
  assign n404 = n403 ^ n402 ;
  assign n405 = x129 & n404 ;
  assign n410 = n409 ^ n405 ;
  assign n411 = n171 & n410 ;
  assign n160 = ~x130 & x131 ;
  assign n397 = x72 & ~x128 ;
  assign n396 = x71 & x128 ;
  assign n398 = n397 ^ n396 ;
  assign n399 = ~x129 & n398 ;
  assign n393 = x70 & ~x128 ;
  assign n392 = x69 & x128 ;
  assign n394 = n393 ^ n392 ;
  assign n395 = x129 & n394 ;
  assign n400 = n399 ^ n395 ;
  assign n401 = n160 & n400 ;
  assign n412 = n411 ^ n401 ;
  assign n413 = ~n391 & ~n412 ;
  assign n414 = n185 & ~n413 ;
  assign n136 = ~x132 & x133 ;
  assign n342 = x96 & ~x128 ;
  assign n341 = x95 & x128 ;
  assign n343 = n342 ^ n341 ;
  assign n344 = ~x129 & n343 ;
  assign n338 = x94 & ~x128 ;
  assign n337 = x93 & x128 ;
  assign n339 = n338 ^ n337 ;
  assign n340 = x129 & n339 ;
  assign n345 = n344 ^ n340 ;
  assign n346 = n148 & n345 ;
  assign n332 = x92 & ~x128 ;
  assign n331 = x91 & x128 ;
  assign n333 = n332 ^ n331 ;
  assign n334 = ~x129 & n333 ;
  assign n328 = x90 & ~x128 ;
  assign n327 = x89 & x128 ;
  assign n329 = n328 ^ n327 ;
  assign n330 = x129 & n329 ;
  assign n335 = n334 ^ n330 ;
  assign n336 = n137 & n335 ;
  assign n347 = n346 ^ n336 ;
  assign n363 = x84 & ~x128 ;
  assign n362 = x83 & x128 ;
  assign n364 = n363 ^ n362 ;
  assign n365 = ~x129 & n364 ;
  assign n359 = x82 & ~x128 ;
  assign n358 = x81 & x128 ;
  assign n360 = n359 ^ n358 ;
  assign n361 = x129 & n360 ;
  assign n366 = n365 ^ n361 ;
  assign n367 = n171 & n366 ;
  assign n353 = x88 & ~x128 ;
  assign n352 = x87 & x128 ;
  assign n354 = n353 ^ n352 ;
  assign n355 = ~x129 & n354 ;
  assign n349 = x86 & ~x128 ;
  assign n348 = x85 & x128 ;
  assign n350 = n349 ^ n348 ;
  assign n351 = x129 & n350 ;
  assign n356 = n355 ^ n351 ;
  assign n357 = n160 & n356 ;
  assign n368 = n367 ^ n357 ;
  assign n369 = ~n347 & ~n368 ;
  assign n370 = n136 & ~n369 ;
  assign n415 = n414 ^ n370 ;
  assign n279 = ~x132 & ~x133 ;
  assign n475 = x127 & x128 ;
  assign n474 = x0 & ~x128 ;
  assign n476 = n475 ^ n474 ;
  assign n477 = ~x129 & n476 ;
  assign n471 = x126 & ~x128 ;
  assign n470 = x125 & x128 ;
  assign n472 = n471 ^ n470 ;
  assign n473 = x129 & n472 ;
  assign n478 = n477 ^ n473 ;
  assign n479 = n148 & n478 ;
  assign n465 = x124 & ~x128 ;
  assign n464 = x123 & x128 ;
  assign n466 = n465 ^ n464 ;
  assign n467 = ~x129 & n466 ;
  assign n461 = x122 & ~x128 ;
  assign n460 = x121 & x128 ;
  assign n462 = n461 ^ n460 ;
  assign n463 = x129 & n462 ;
  assign n468 = n467 ^ n463 ;
  assign n469 = n137 & n468 ;
  assign n480 = n479 ^ n469 ;
  assign n496 = x116 & ~x128 ;
  assign n495 = x115 & x128 ;
  assign n497 = n496 ^ n495 ;
  assign n498 = ~x129 & n497 ;
  assign n492 = x114 & ~x128 ;
  assign n491 = x113 & x128 ;
  assign n493 = n492 ^ n491 ;
  assign n494 = x129 & n493 ;
  assign n499 = n498 ^ n494 ;
  assign n500 = n171 & n499 ;
  assign n486 = x120 & ~x128 ;
  assign n485 = x119 & x128 ;
  assign n487 = n486 ^ n485 ;
  assign n488 = ~x129 & n487 ;
  assign n482 = x118 & ~x128 ;
  assign n481 = x117 & x128 ;
  assign n483 = n482 ^ n481 ;
  assign n484 = x129 & n483 ;
  assign n489 = n488 ^ n484 ;
  assign n490 = n160 & n489 ;
  assign n501 = n500 ^ n490 ;
  assign n502 = ~n480 & ~n501 ;
  assign n503 = n279 & ~n502 ;
  assign n254 = x132 & ~x133 ;
  assign n431 = x112 & ~x128 ;
  assign n430 = x111 & x128 ;
  assign n432 = n431 ^ n430 ;
  assign n433 = ~x129 & n432 ;
  assign n427 = x110 & ~x128 ;
  assign n426 = x109 & x128 ;
  assign n428 = n427 ^ n426 ;
  assign n429 = x129 & n428 ;
  assign n434 = n433 ^ n429 ;
  assign n435 = n148 & n434 ;
  assign n421 = x108 & ~x128 ;
  assign n420 = x107 & x128 ;
  assign n422 = n421 ^ n420 ;
  assign n423 = ~x129 & n422 ;
  assign n417 = x106 & ~x128 ;
  assign n416 = x105 & x128 ;
  assign n418 = n417 ^ n416 ;
  assign n419 = x129 & n418 ;
  assign n424 = n423 ^ n419 ;
  assign n425 = n137 & n424 ;
  assign n436 = n435 ^ n425 ;
  assign n452 = x100 & ~x128 ;
  assign n451 = x99 & x128 ;
  assign n453 = n452 ^ n451 ;
  assign n454 = ~x129 & n453 ;
  assign n448 = x98 & ~x128 ;
  assign n447 = x97 & x128 ;
  assign n449 = n448 ^ n447 ;
  assign n450 = x129 & n449 ;
  assign n455 = n454 ^ n450 ;
  assign n456 = n171 & n455 ;
  assign n442 = x104 & ~x128 ;
  assign n441 = x103 & x128 ;
  assign n443 = n442 ^ n441 ;
  assign n444 = ~x129 & n443 ;
  assign n438 = x102 & ~x128 ;
  assign n437 = x101 & x128 ;
  assign n439 = n438 ^ n437 ;
  assign n440 = x129 & n439 ;
  assign n445 = n444 ^ n440 ;
  assign n446 = n160 & n445 ;
  assign n457 = n456 ^ n446 ;
  assign n458 = ~n436 & ~n457 ;
  assign n459 = n254 & ~n458 ;
  assign n504 = n503 ^ n459 ;
  assign n505 = ~n415 & ~n504 ;
  assign n506 = ~x134 & n505 ;
  assign n201 = x16 & ~x128 ;
  assign n200 = x15 & x128 ;
  assign n202 = n201 ^ n200 ;
  assign n203 = ~x129 & n202 ;
  assign n197 = x14 & ~x128 ;
  assign n196 = x13 & x128 ;
  assign n198 = n197 ^ n196 ;
  assign n199 = x129 & n198 ;
  assign n204 = n203 ^ n199 ;
  assign n205 = n148 & n204 ;
  assign n191 = x12 & ~x128 ;
  assign n190 = x11 & x128 ;
  assign n192 = n191 ^ n190 ;
  assign n193 = ~x129 & n192 ;
  assign n187 = x10 & ~x128 ;
  assign n186 = x9 & x128 ;
  assign n188 = n187 ^ n186 ;
  assign n189 = x129 & n188 ;
  assign n194 = n193 ^ n189 ;
  assign n195 = n137 & n194 ;
  assign n206 = n205 ^ n195 ;
  assign n222 = x4 & ~x128 ;
  assign n221 = x3 & x128 ;
  assign n223 = n222 ^ n221 ;
  assign n224 = ~x129 & n223 ;
  assign n218 = x2 & ~x128 ;
  assign n217 = x1 & x128 ;
  assign n219 = n218 ^ n217 ;
  assign n220 = x129 & n219 ;
  assign n225 = n224 ^ n220 ;
  assign n226 = n171 & n225 ;
  assign n212 = x8 & ~x128 ;
  assign n211 = x7 & x128 ;
  assign n213 = n212 ^ n211 ;
  assign n214 = ~x129 & n213 ;
  assign n208 = x6 & ~x128 ;
  assign n207 = x5 & x128 ;
  assign n209 = n208 ^ n207 ;
  assign n210 = x129 & n209 ;
  assign n215 = n214 ^ n210 ;
  assign n216 = n160 & n215 ;
  assign n227 = n226 ^ n216 ;
  assign n228 = ~n206 & ~n227 ;
  assign n229 = n185 & ~n228 ;
  assign n154 = x32 & ~x128 ;
  assign n153 = x31 & x128 ;
  assign n155 = n154 ^ n153 ;
  assign n156 = ~x129 & n155 ;
  assign n150 = x30 & ~x128 ;
  assign n149 = x29 & x128 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = x129 & n151 ;
  assign n157 = n156 ^ n152 ;
  assign n158 = n148 & n157 ;
  assign n143 = x28 & ~x128 ;
  assign n142 = x27 & x128 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = ~x129 & n144 ;
  assign n139 = x26 & ~x128 ;
  assign n138 = x25 & x128 ;
  assign n140 = n139 ^ n138 ;
  assign n141 = x129 & n140 ;
  assign n146 = n145 ^ n141 ;
  assign n147 = n137 & n146 ;
  assign n159 = n158 ^ n147 ;
  assign n177 = x20 & ~x128 ;
  assign n176 = x19 & x128 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = ~x129 & n178 ;
  assign n173 = x18 & ~x128 ;
  assign n172 = x17 & x128 ;
  assign n174 = n173 ^ n172 ;
  assign n175 = x129 & n174 ;
  assign n180 = n179 ^ n175 ;
  assign n181 = n171 & n180 ;
  assign n166 = x24 & ~x128 ;
  assign n165 = x23 & x128 ;
  assign n167 = n166 ^ n165 ;
  assign n168 = ~x129 & n167 ;
  assign n162 = x22 & ~x128 ;
  assign n161 = x21 & x128 ;
  assign n163 = n162 ^ n161 ;
  assign n164 = x129 & n163 ;
  assign n169 = n168 ^ n164 ;
  assign n170 = n160 & n169 ;
  assign n182 = n181 ^ n170 ;
  assign n183 = ~n159 & ~n182 ;
  assign n184 = n136 & ~n183 ;
  assign n230 = n229 ^ n184 ;
  assign n295 = x64 & ~x128 ;
  assign n294 = x63 & x128 ;
  assign n296 = n295 ^ n294 ;
  assign n297 = ~x129 & n296 ;
  assign n291 = x62 & ~x128 ;
  assign n290 = x61 & x128 ;
  assign n292 = n291 ^ n290 ;
  assign n293 = x129 & n292 ;
  assign n298 = n297 ^ n293 ;
  assign n299 = n148 & n298 ;
  assign n285 = x60 & ~x128 ;
  assign n284 = x59 & x128 ;
  assign n286 = n285 ^ n284 ;
  assign n287 = ~x129 & n286 ;
  assign n281 = x58 & ~x128 ;
  assign n280 = x57 & x128 ;
  assign n282 = n281 ^ n280 ;
  assign n283 = x129 & n282 ;
  assign n288 = n287 ^ n283 ;
  assign n289 = n137 & n288 ;
  assign n300 = n299 ^ n289 ;
  assign n316 = x52 & ~x128 ;
  assign n315 = x51 & x128 ;
  assign n317 = n316 ^ n315 ;
  assign n318 = ~x129 & n317 ;
  assign n312 = x50 & ~x128 ;
  assign n311 = x49 & x128 ;
  assign n313 = n312 ^ n311 ;
  assign n314 = x129 & n313 ;
  assign n319 = n318 ^ n314 ;
  assign n320 = n171 & n319 ;
  assign n306 = x56 & ~x128 ;
  assign n305 = x55 & x128 ;
  assign n307 = n306 ^ n305 ;
  assign n308 = ~x129 & n307 ;
  assign n302 = x54 & ~x128 ;
  assign n301 = x53 & x128 ;
  assign n303 = n302 ^ n301 ;
  assign n304 = x129 & n303 ;
  assign n309 = n308 ^ n304 ;
  assign n310 = n160 & n309 ;
  assign n321 = n320 ^ n310 ;
  assign n322 = ~n300 & ~n321 ;
  assign n323 = n279 & n322 ;
  assign n248 = x36 & ~x128 ;
  assign n247 = x35 & x128 ;
  assign n249 = n248 ^ n247 ;
  assign n250 = ~x129 & n249 ;
  assign n244 = x34 & ~x128 ;
  assign n243 = x33 & x128 ;
  assign n245 = n244 ^ n243 ;
  assign n246 = x129 & n245 ;
  assign n251 = n250 ^ n246 ;
  assign n252 = n171 & n251 ;
  assign n233 = x39 & x128 ;
  assign n234 = ~x129 & n233 ;
  assign n231 = x38 & ~x128 ;
  assign n232 = x129 & n231 ;
  assign n235 = n234 ^ n232 ;
  assign n238 = x40 & ~x128 ;
  assign n239 = ~x129 & ~n238 ;
  assign n236 = x37 & x128 ;
  assign n237 = x129 & ~n236 ;
  assign n240 = n239 ^ n237 ;
  assign n241 = ~n235 & n240 ;
  assign n242 = n160 & ~n241 ;
  assign n253 = n252 ^ n242 ;
  assign n270 = x48 & ~x128 ;
  assign n269 = x47 & x128 ;
  assign n271 = n270 ^ n269 ;
  assign n272 = ~x129 & n271 ;
  assign n266 = x46 & ~x128 ;
  assign n265 = x45 & x128 ;
  assign n267 = n266 ^ n265 ;
  assign n268 = x129 & n267 ;
  assign n273 = n272 ^ n268 ;
  assign n274 = n148 & n273 ;
  assign n260 = x44 & ~x128 ;
  assign n259 = x43 & x128 ;
  assign n261 = n260 ^ n259 ;
  assign n262 = ~x129 & n261 ;
  assign n256 = x42 & ~x128 ;
  assign n255 = x41 & x128 ;
  assign n257 = n256 ^ n255 ;
  assign n258 = x129 & n257 ;
  assign n263 = n262 ^ n258 ;
  assign n264 = n137 & n263 ;
  assign n275 = n274 ^ n264 ;
  assign n276 = n254 & ~n275 ;
  assign n277 = ~n253 & n276 ;
  assign n278 = n277 ^ x133 ;
  assign n324 = n323 ^ n278 ;
  assign n325 = ~n230 & n324 ;
  assign n326 = x134 & n325 ;
  assign n507 = n506 ^ n326 ;
  assign n782 = x80 & x128 ;
  assign n783 = ~x129 & n782 ;
  assign n780 = x79 & ~x128 ;
  assign n781 = x129 & n780 ;
  assign n784 = n783 ^ n781 ;
  assign n787 = x81 & ~x128 ;
  assign n788 = ~x129 & ~n787 ;
  assign n785 = x78 & x128 ;
  assign n786 = x129 & ~n785 ;
  assign n789 = n788 ^ n786 ;
  assign n790 = ~n784 & n789 ;
  assign n791 = n148 & ~n790 ;
  assign n770 = x76 & x128 ;
  assign n771 = ~x129 & n770 ;
  assign n768 = x75 & ~x128 ;
  assign n769 = x129 & n768 ;
  assign n772 = n771 ^ n769 ;
  assign n775 = x77 & ~x128 ;
  assign n776 = ~x129 & ~n775 ;
  assign n773 = x74 & x128 ;
  assign n774 = x129 & ~n773 ;
  assign n777 = n776 ^ n774 ;
  assign n778 = ~n772 & n777 ;
  assign n779 = n137 & ~n778 ;
  assign n792 = n791 ^ n779 ;
  assign n807 = x68 & x128 ;
  assign n808 = ~x129 & n807 ;
  assign n805 = x67 & ~x128 ;
  assign n806 = x129 & n805 ;
  assign n809 = n808 ^ n806 ;
  assign n812 = x69 & ~x128 ;
  assign n813 = ~x129 & ~n812 ;
  assign n810 = x66 & x128 ;
  assign n811 = x129 & ~n810 ;
  assign n814 = n813 ^ n811 ;
  assign n815 = ~n809 & n814 ;
  assign n816 = n171 & ~n815 ;
  assign n795 = x72 & x128 ;
  assign n796 = ~x129 & n795 ;
  assign n793 = x71 & ~x128 ;
  assign n794 = x129 & n793 ;
  assign n797 = n796 ^ n794 ;
  assign n800 = x73 & ~x128 ;
  assign n801 = ~x129 & ~n800 ;
  assign n798 = x70 & x128 ;
  assign n799 = x129 & ~n798 ;
  assign n802 = n801 ^ n799 ;
  assign n803 = ~n797 & n802 ;
  assign n804 = n160 & ~n803 ;
  assign n817 = n816 ^ n804 ;
  assign n818 = ~n792 & ~n817 ;
  assign n819 = n185 & ~n818 ;
  assign n730 = x96 & x128 ;
  assign n731 = ~x129 & n730 ;
  assign n728 = x95 & ~x128 ;
  assign n729 = x129 & n728 ;
  assign n732 = n731 ^ n729 ;
  assign n735 = x97 & ~x128 ;
  assign n736 = ~x129 & ~n735 ;
  assign n733 = x94 & x128 ;
  assign n734 = x129 & ~n733 ;
  assign n737 = n736 ^ n734 ;
  assign n738 = ~n732 & n737 ;
  assign n739 = n148 & ~n738 ;
  assign n718 = x92 & x128 ;
  assign n719 = ~x129 & n718 ;
  assign n716 = x91 & ~x128 ;
  assign n717 = x129 & n716 ;
  assign n720 = n719 ^ n717 ;
  assign n723 = x93 & ~x128 ;
  assign n724 = ~x129 & ~n723 ;
  assign n721 = x90 & x128 ;
  assign n722 = x129 & ~n721 ;
  assign n725 = n724 ^ n722 ;
  assign n726 = ~n720 & n725 ;
  assign n727 = n137 & ~n726 ;
  assign n740 = n739 ^ n727 ;
  assign n755 = x84 & x128 ;
  assign n756 = ~x129 & n755 ;
  assign n753 = x83 & ~x128 ;
  assign n754 = x129 & n753 ;
  assign n757 = n756 ^ n754 ;
  assign n760 = x85 & ~x128 ;
  assign n761 = ~x129 & ~n760 ;
  assign n758 = x82 & x128 ;
  assign n759 = x129 & ~n758 ;
  assign n762 = n761 ^ n759 ;
  assign n763 = ~n757 & n762 ;
  assign n764 = n171 & ~n763 ;
  assign n743 = x88 & x128 ;
  assign n744 = ~x129 & n743 ;
  assign n741 = x87 & ~x128 ;
  assign n742 = x129 & n741 ;
  assign n745 = n744 ^ n742 ;
  assign n748 = x89 & ~x128 ;
  assign n749 = ~x129 & ~n748 ;
  assign n746 = x86 & x128 ;
  assign n747 = x129 & ~n746 ;
  assign n750 = n749 ^ n747 ;
  assign n751 = ~n745 & n750 ;
  assign n752 = n160 & ~n751 ;
  assign n765 = n764 ^ n752 ;
  assign n766 = ~n740 & ~n765 ;
  assign n767 = n136 & ~n766 ;
  assign n820 = n819 ^ n767 ;
  assign n887 = x0 & x128 ;
  assign n888 = ~x129 & n887 ;
  assign n885 = x127 & ~x128 ;
  assign n886 = x129 & n885 ;
  assign n889 = n888 ^ n886 ;
  assign n892 = x1 & ~x128 ;
  assign n893 = ~x129 & ~n892 ;
  assign n890 = x126 & x128 ;
  assign n891 = x129 & ~n890 ;
  assign n894 = n893 ^ n891 ;
  assign n895 = ~n889 & n894 ;
  assign n896 = n148 & ~n895 ;
  assign n875 = x124 & x128 ;
  assign n876 = ~x129 & n875 ;
  assign n873 = x123 & ~x128 ;
  assign n874 = x129 & n873 ;
  assign n877 = n876 ^ n874 ;
  assign n880 = x125 & ~x128 ;
  assign n881 = ~x129 & ~n880 ;
  assign n878 = x122 & x128 ;
  assign n879 = x129 & ~n878 ;
  assign n882 = n881 ^ n879 ;
  assign n883 = ~n877 & n882 ;
  assign n884 = n137 & ~n883 ;
  assign n897 = n896 ^ n884 ;
  assign n912 = x116 & x128 ;
  assign n913 = ~x129 & n912 ;
  assign n910 = x115 & ~x128 ;
  assign n911 = x129 & n910 ;
  assign n914 = n913 ^ n911 ;
  assign n917 = x117 & ~x128 ;
  assign n918 = ~x129 & ~n917 ;
  assign n915 = x114 & x128 ;
  assign n916 = x129 & ~n915 ;
  assign n919 = n918 ^ n916 ;
  assign n920 = ~n914 & n919 ;
  assign n921 = n171 & ~n920 ;
  assign n900 = x120 & x128 ;
  assign n901 = ~x129 & n900 ;
  assign n898 = x119 & ~x128 ;
  assign n899 = x129 & n898 ;
  assign n902 = n901 ^ n899 ;
  assign n905 = x121 & ~x128 ;
  assign n906 = ~x129 & ~n905 ;
  assign n903 = x118 & x128 ;
  assign n904 = x129 & ~n903 ;
  assign n907 = n906 ^ n904 ;
  assign n908 = ~n902 & n907 ;
  assign n909 = n160 & ~n908 ;
  assign n922 = n921 ^ n909 ;
  assign n923 = ~n897 & ~n922 ;
  assign n924 = n279 & ~n923 ;
  assign n835 = x112 & x128 ;
  assign n836 = ~x129 & n835 ;
  assign n833 = x111 & ~x128 ;
  assign n834 = x129 & n833 ;
  assign n837 = n836 ^ n834 ;
  assign n840 = x113 & ~x128 ;
  assign n841 = ~x129 & ~n840 ;
  assign n838 = x110 & x128 ;
  assign n839 = x129 & ~n838 ;
  assign n842 = n841 ^ n839 ;
  assign n843 = ~n837 & n842 ;
  assign n844 = n148 & ~n843 ;
  assign n823 = x108 & x128 ;
  assign n824 = ~x129 & n823 ;
  assign n821 = x107 & ~x128 ;
  assign n822 = x129 & n821 ;
  assign n825 = n824 ^ n822 ;
  assign n828 = x109 & ~x128 ;
  assign n829 = ~x129 & ~n828 ;
  assign n826 = x106 & x128 ;
  assign n827 = x129 & ~n826 ;
  assign n830 = n829 ^ n827 ;
  assign n831 = ~n825 & n830 ;
  assign n832 = n137 & ~n831 ;
  assign n845 = n844 ^ n832 ;
  assign n860 = x100 & x128 ;
  assign n861 = ~x129 & n860 ;
  assign n858 = x99 & ~x128 ;
  assign n859 = x129 & n858 ;
  assign n862 = n861 ^ n859 ;
  assign n865 = x101 & ~x128 ;
  assign n866 = ~x129 & ~n865 ;
  assign n863 = x98 & x128 ;
  assign n864 = x129 & ~n863 ;
  assign n867 = n866 ^ n864 ;
  assign n868 = ~n862 & n867 ;
  assign n869 = n171 & ~n868 ;
  assign n848 = x104 & x128 ;
  assign n849 = ~x129 & n848 ;
  assign n846 = x103 & ~x128 ;
  assign n847 = x129 & n846 ;
  assign n850 = n849 ^ n847 ;
  assign n853 = x105 & ~x128 ;
  assign n854 = ~x129 & ~n853 ;
  assign n851 = x102 & x128 ;
  assign n852 = x129 & ~n851 ;
  assign n855 = n854 ^ n852 ;
  assign n856 = ~n850 & n855 ;
  assign n857 = n160 & ~n856 ;
  assign n870 = n869 ^ n857 ;
  assign n871 = ~n845 & ~n870 ;
  assign n872 = n254 & ~n871 ;
  assign n925 = n924 ^ n872 ;
  assign n926 = ~n820 & ~n925 ;
  assign n927 = ~x134 & n926 ;
  assign n574 = x64 & x128 ;
  assign n575 = ~x129 & n574 ;
  assign n572 = x63 & ~x128 ;
  assign n573 = x129 & n572 ;
  assign n576 = n575 ^ n573 ;
  assign n579 = x65 & ~x128 ;
  assign n580 = ~x129 & ~n579 ;
  assign n577 = x62 & x128 ;
  assign n578 = x129 & ~n577 ;
  assign n581 = n580 ^ n578 ;
  assign n582 = ~n576 & n581 ;
  assign n583 = n148 & ~n582 ;
  assign n562 = x60 & x128 ;
  assign n563 = ~x129 & n562 ;
  assign n560 = x59 & ~x128 ;
  assign n561 = x129 & n560 ;
  assign n564 = n563 ^ n561 ;
  assign n567 = x61 & ~x128 ;
  assign n568 = ~x129 & ~n567 ;
  assign n565 = x58 & x128 ;
  assign n566 = x129 & ~n565 ;
  assign n569 = n568 ^ n566 ;
  assign n570 = ~n564 & n569 ;
  assign n571 = n137 & ~n570 ;
  assign n584 = n583 ^ n571 ;
  assign n599 = x52 & x128 ;
  assign n600 = ~x129 & n599 ;
  assign n597 = x51 & ~x128 ;
  assign n598 = x129 & n597 ;
  assign n601 = n600 ^ n598 ;
  assign n604 = x53 & ~x128 ;
  assign n605 = ~x129 & ~n604 ;
  assign n602 = x50 & x128 ;
  assign n603 = x129 & ~n602 ;
  assign n606 = n605 ^ n603 ;
  assign n607 = ~n601 & n606 ;
  assign n608 = n171 & ~n607 ;
  assign n587 = x56 & x128 ;
  assign n588 = ~x129 & n587 ;
  assign n585 = x55 & ~x128 ;
  assign n586 = x129 & n585 ;
  assign n589 = n588 ^ n586 ;
  assign n592 = x57 & ~x128 ;
  assign n593 = ~x129 & ~n592 ;
  assign n590 = x54 & x128 ;
  assign n591 = x129 & ~n590 ;
  assign n594 = n593 ^ n591 ;
  assign n595 = ~n589 & n594 ;
  assign n596 = n160 & ~n595 ;
  assign n609 = n608 ^ n596 ;
  assign n610 = ~n584 & ~n609 ;
  assign n611 = n279 & ~n610 ;
  assign n522 = x16 & x128 ;
  assign n523 = ~x129 & n522 ;
  assign n520 = x15 & ~x128 ;
  assign n521 = x129 & n520 ;
  assign n524 = n523 ^ n521 ;
  assign n527 = x17 & ~x128 ;
  assign n528 = ~x129 & ~n527 ;
  assign n525 = x14 & x128 ;
  assign n526 = x129 & ~n525 ;
  assign n529 = n528 ^ n526 ;
  assign n530 = ~n524 & n529 ;
  assign n531 = n148 & ~n530 ;
  assign n510 = x12 & x128 ;
  assign n511 = ~x129 & n510 ;
  assign n508 = x11 & ~x128 ;
  assign n509 = x129 & n508 ;
  assign n512 = n511 ^ n509 ;
  assign n515 = x13 & ~x128 ;
  assign n516 = ~x129 & ~n515 ;
  assign n513 = x10 & x128 ;
  assign n514 = x129 & ~n513 ;
  assign n517 = n516 ^ n514 ;
  assign n518 = ~n512 & n517 ;
  assign n519 = n137 & ~n518 ;
  assign n532 = n531 ^ n519 ;
  assign n547 = x4 & x128 ;
  assign n548 = ~x129 & n547 ;
  assign n545 = x3 & ~x128 ;
  assign n546 = x129 & n545 ;
  assign n549 = n548 ^ n546 ;
  assign n552 = x5 & ~x128 ;
  assign n553 = ~x129 & ~n552 ;
  assign n550 = x2 & x128 ;
  assign n551 = x129 & ~n550 ;
  assign n554 = n553 ^ n551 ;
  assign n555 = ~n549 & n554 ;
  assign n556 = n171 & ~n555 ;
  assign n535 = x8 & x128 ;
  assign n536 = ~x129 & n535 ;
  assign n533 = x7 & ~x128 ;
  assign n534 = x129 & n533 ;
  assign n537 = n536 ^ n534 ;
  assign n540 = x9 & ~x128 ;
  assign n541 = ~x129 & ~n540 ;
  assign n538 = x6 & x128 ;
  assign n539 = x129 & ~n538 ;
  assign n542 = n541 ^ n539 ;
  assign n543 = ~n537 & n542 ;
  assign n544 = n160 & ~n543 ;
  assign n557 = n556 ^ n544 ;
  assign n558 = ~n532 & ~n557 ;
  assign n559 = n185 & ~n558 ;
  assign n612 = n611 ^ n559 ;
  assign n677 = x48 & x128 ;
  assign n678 = ~x129 & n677 ;
  assign n675 = x47 & ~x128 ;
  assign n676 = x129 & n675 ;
  assign n679 = n678 ^ n676 ;
  assign n682 = x49 & ~x128 ;
  assign n683 = ~x129 & ~n682 ;
  assign n680 = x46 & x128 ;
  assign n681 = x129 & ~n680 ;
  assign n684 = n683 ^ n681 ;
  assign n685 = ~n679 & n684 ;
  assign n686 = n148 & ~n685 ;
  assign n670 = x45 & ~x128 ;
  assign n669 = x44 & x128 ;
  assign n671 = n670 ^ n669 ;
  assign n672 = ~x129 & ~n671 ;
  assign n666 = ~x43 & ~x128 ;
  assign n665 = ~x42 & x128 ;
  assign n667 = n666 ^ n665 ;
  assign n668 = x129 & n667 ;
  assign n673 = n672 ^ n668 ;
  assign n674 = n137 & ~n673 ;
  assign n687 = n686 ^ n674 ;
  assign n700 = x36 & x128 ;
  assign n701 = ~x129 & n700 ;
  assign n698 = x35 & ~x128 ;
  assign n699 = x129 & n698 ;
  assign n702 = n701 ^ n699 ;
  assign n705 = x37 & ~x128 ;
  assign n706 = ~x129 & ~n705 ;
  assign n703 = x34 & x128 ;
  assign n704 = x129 & ~n703 ;
  assign n707 = n706 ^ n704 ;
  assign n708 = ~n702 & n707 ;
  assign n709 = n171 & ~n708 ;
  assign n693 = ~x41 & ~x128 ;
  assign n692 = ~x40 & x128 ;
  assign n694 = n693 ^ n692 ;
  assign n695 = ~x129 & n694 ;
  assign n689 = ~x39 & ~x128 ;
  assign n688 = ~x38 & x128 ;
  assign n690 = n689 ^ n688 ;
  assign n691 = x129 & n690 ;
  assign n696 = n695 ^ n691 ;
  assign n697 = n160 & ~n696 ;
  assign n710 = n709 ^ n697 ;
  assign n711 = ~n687 & ~n710 ;
  assign n712 = n254 & ~n711 ;
  assign n627 = x32 & x128 ;
  assign n628 = ~x129 & n627 ;
  assign n625 = x31 & ~x128 ;
  assign n626 = x129 & n625 ;
  assign n629 = n628 ^ n626 ;
  assign n632 = x33 & ~x128 ;
  assign n633 = ~x129 & ~n632 ;
  assign n630 = x30 & x128 ;
  assign n631 = x129 & ~n630 ;
  assign n634 = n633 ^ n631 ;
  assign n635 = ~n629 & n634 ;
  assign n636 = n148 & ~n635 ;
  assign n615 = x28 & x128 ;
  assign n616 = ~x129 & n615 ;
  assign n613 = x27 & ~x128 ;
  assign n614 = x129 & n613 ;
  assign n617 = n616 ^ n614 ;
  assign n620 = x29 & ~x128 ;
  assign n621 = ~x129 & ~n620 ;
  assign n618 = x26 & x128 ;
  assign n619 = x129 & ~n618 ;
  assign n622 = n621 ^ n619 ;
  assign n623 = ~n617 & n622 ;
  assign n624 = n137 & ~n623 ;
  assign n637 = n636 ^ n624 ;
  assign n652 = x20 & x128 ;
  assign n653 = ~x129 & n652 ;
  assign n650 = x19 & ~x128 ;
  assign n651 = x129 & n650 ;
  assign n654 = n653 ^ n651 ;
  assign n657 = x21 & ~x128 ;
  assign n658 = ~x129 & ~n657 ;
  assign n655 = x18 & x128 ;
  assign n656 = x129 & ~n655 ;
  assign n659 = n658 ^ n656 ;
  assign n660 = ~n654 & n659 ;
  assign n661 = n171 & ~n660 ;
  assign n640 = x24 & x128 ;
  assign n641 = ~x129 & n640 ;
  assign n638 = x23 & ~x128 ;
  assign n639 = x129 & n638 ;
  assign n642 = n641 ^ n639 ;
  assign n645 = x25 & ~x128 ;
  assign n646 = ~x129 & ~n645 ;
  assign n643 = x22 & x128 ;
  assign n644 = x129 & ~n643 ;
  assign n647 = n646 ^ n644 ;
  assign n648 = ~n642 & n647 ;
  assign n649 = n160 & ~n648 ;
  assign n662 = n661 ^ n649 ;
  assign n663 = ~n637 & ~n662 ;
  assign n664 = n136 & ~n663 ;
  assign n713 = n712 ^ n664 ;
  assign n714 = ~n612 & ~n713 ;
  assign n715 = x134 & n714 ;
  assign n928 = n927 ^ n715 ;
  assign n1044 = ~x129 & n360 ;
  assign n1043 = x129 & n387 ;
  assign n1045 = n1044 ^ n1043 ;
  assign n1046 = n148 & n1045 ;
  assign n1040 = ~x129 & n383 ;
  assign n1039 = x129 & n377 ;
  assign n1041 = n1040 ^ n1039 ;
  assign n1042 = n137 & n1041 ;
  assign n1047 = n1046 ^ n1042 ;
  assign n1053 = ~x129 & n394 ;
  assign n1052 = x129 & n408 ;
  assign n1054 = n1053 ^ n1052 ;
  assign n1055 = n171 & n1054 ;
  assign n1049 = ~x129 & n373 ;
  assign n1048 = x129 & n398 ;
  assign n1050 = n1049 ^ n1048 ;
  assign n1051 = n160 & n1050 ;
  assign n1056 = n1055 ^ n1051 ;
  assign n1057 = ~n1047 & ~n1056 ;
  assign n1058 = n185 & ~n1057 ;
  assign n1024 = ~x129 & n449 ;
  assign n1023 = x129 & n343 ;
  assign n1025 = n1024 ^ n1023 ;
  assign n1026 = n148 & n1025 ;
  assign n1020 = ~x129 & n339 ;
  assign n1019 = x129 & n333 ;
  assign n1021 = n1020 ^ n1019 ;
  assign n1022 = n137 & n1021 ;
  assign n1027 = n1026 ^ n1022 ;
  assign n1033 = ~x129 & n350 ;
  assign n1032 = x129 & n364 ;
  assign n1034 = n1033 ^ n1032 ;
  assign n1035 = n171 & n1034 ;
  assign n1029 = ~x129 & n329 ;
  assign n1028 = x129 & n354 ;
  assign n1030 = n1029 ^ n1028 ;
  assign n1031 = n160 & n1030 ;
  assign n1036 = n1035 ^ n1031 ;
  assign n1037 = ~n1027 & ~n1036 ;
  assign n1038 = n136 & ~n1037 ;
  assign n1059 = n1058 ^ n1038 ;
  assign n1085 = ~x129 & n219 ;
  assign n1084 = x129 & n476 ;
  assign n1086 = n1085 ^ n1084 ;
  assign n1087 = n148 & n1086 ;
  assign n1081 = ~x129 & n472 ;
  assign n1080 = x129 & n466 ;
  assign n1082 = n1081 ^ n1080 ;
  assign n1083 = n137 & n1082 ;
  assign n1088 = n1087 ^ n1083 ;
  assign n1094 = ~x129 & n483 ;
  assign n1093 = x129 & n497 ;
  assign n1095 = n1094 ^ n1093 ;
  assign n1096 = n171 & n1095 ;
  assign n1090 = ~x129 & n462 ;
  assign n1089 = x129 & n487 ;
  assign n1091 = n1090 ^ n1089 ;
  assign n1092 = n160 & n1091 ;
  assign n1097 = n1096 ^ n1092 ;
  assign n1098 = ~n1088 & ~n1097 ;
  assign n1099 = n279 & ~n1098 ;
  assign n1065 = ~x129 & n493 ;
  assign n1064 = x129 & n432 ;
  assign n1066 = n1065 ^ n1064 ;
  assign n1067 = n148 & n1066 ;
  assign n1061 = ~x129 & n428 ;
  assign n1060 = x129 & n422 ;
  assign n1062 = n1061 ^ n1060 ;
  assign n1063 = n137 & n1062 ;
  assign n1068 = n1067 ^ n1063 ;
  assign n1074 = ~x129 & n439 ;
  assign n1073 = x129 & n453 ;
  assign n1075 = n1074 ^ n1073 ;
  assign n1076 = n171 & n1075 ;
  assign n1070 = ~x129 & n418 ;
  assign n1069 = x129 & n443 ;
  assign n1071 = n1070 ^ n1069 ;
  assign n1072 = n160 & n1071 ;
  assign n1077 = n1076 ^ n1072 ;
  assign n1078 = ~n1068 & ~n1077 ;
  assign n1079 = n254 & ~n1078 ;
  assign n1100 = n1099 ^ n1079 ;
  assign n1101 = ~n1059 & ~n1100 ;
  assign n1102 = ~x134 & n1101 ;
  assign n954 = ~x129 & n404 ;
  assign n953 = x129 & n296 ;
  assign n955 = n954 ^ n953 ;
  assign n956 = n148 & n955 ;
  assign n950 = ~x129 & n292 ;
  assign n949 = x129 & n286 ;
  assign n951 = n950 ^ n949 ;
  assign n952 = n137 & n951 ;
  assign n957 = n956 ^ n952 ;
  assign n963 = ~x129 & n303 ;
  assign n962 = x129 & n317 ;
  assign n964 = n963 ^ n962 ;
  assign n965 = n171 & n964 ;
  assign n959 = ~x129 & n282 ;
  assign n958 = x129 & n307 ;
  assign n960 = n959 ^ n958 ;
  assign n961 = n160 & n960 ;
  assign n966 = n965 ^ n961 ;
  assign n967 = ~n957 & ~n966 ;
  assign n968 = n279 & ~n967 ;
  assign n934 = ~x129 & n174 ;
  assign n933 = x129 & n202 ;
  assign n935 = n934 ^ n933 ;
  assign n936 = n148 & n935 ;
  assign n930 = ~x129 & n198 ;
  assign n929 = x129 & n192 ;
  assign n931 = n930 ^ n929 ;
  assign n932 = n137 & n931 ;
  assign n937 = n936 ^ n932 ;
  assign n943 = ~x129 & n209 ;
  assign n942 = x129 & n223 ;
  assign n944 = n943 ^ n942 ;
  assign n945 = n171 & n944 ;
  assign n939 = ~x129 & n188 ;
  assign n938 = x129 & n213 ;
  assign n940 = n939 ^ n938 ;
  assign n941 = n160 & n940 ;
  assign n946 = n945 ^ n941 ;
  assign n947 = ~n937 & ~n946 ;
  assign n948 = n185 & ~n947 ;
  assign n969 = n968 ^ n948 ;
  assign n995 = ~x129 & n313 ;
  assign n994 = x129 & n271 ;
  assign n996 = n995 ^ n994 ;
  assign n997 = n148 & n996 ;
  assign n991 = ~x129 & n267 ;
  assign n990 = x129 & n261 ;
  assign n992 = n991 ^ n990 ;
  assign n993 = n137 & n992 ;
  assign n998 = n997 ^ n993 ;
  assign n1008 = ~x38 & ~x128 ;
  assign n1007 = ~x37 & x128 ;
  assign n1009 = n1008 ^ n1007 ;
  assign n1010 = ~x129 & n1009 ;
  assign n1006 = x129 & ~n249 ;
  assign n1011 = n1010 ^ n1006 ;
  assign n1012 = n171 & ~n1011 ;
  assign n1003 = ~x129 & ~n257 ;
  assign n1000 = ~x40 & ~x128 ;
  assign n999 = ~x39 & x128 ;
  assign n1001 = n1000 ^ n999 ;
  assign n1002 = x129 & n1001 ;
  assign n1004 = n1003 ^ n1002 ;
  assign n1005 = n160 & ~n1004 ;
  assign n1013 = n1012 ^ n1005 ;
  assign n1014 = ~n998 & ~n1013 ;
  assign n1015 = n254 & ~n1014 ;
  assign n975 = ~x129 & n245 ;
  assign n974 = x129 & n155 ;
  assign n976 = n975 ^ n974 ;
  assign n977 = n148 & n976 ;
  assign n971 = ~x129 & n151 ;
  assign n970 = x129 & n144 ;
  assign n972 = n971 ^ n970 ;
  assign n973 = n137 & n972 ;
  assign n978 = n977 ^ n973 ;
  assign n984 = ~x129 & n163 ;
  assign n983 = x129 & n178 ;
  assign n985 = n984 ^ n983 ;
  assign n986 = n171 & n985 ;
  assign n980 = ~x129 & n140 ;
  assign n979 = x129 & n167 ;
  assign n981 = n980 ^ n979 ;
  assign n982 = n160 & n981 ;
  assign n987 = n986 ^ n982 ;
  assign n988 = ~n978 & ~n987 ;
  assign n989 = n136 & ~n988 ;
  assign n1016 = n1015 ^ n989 ;
  assign n1017 = ~n969 & ~n1016 ;
  assign n1018 = x134 & n1017 ;
  assign n1103 = n1102 ^ n1018 ;
  assign n1302 = ~x129 & n910 ;
  assign n1301 = x129 & n835 ;
  assign n1303 = n1302 ^ n1301 ;
  assign n1305 = ~x129 & ~n915 ;
  assign n1304 = x129 & ~n840 ;
  assign n1306 = n1305 ^ n1304 ;
  assign n1307 = ~n1303 & n1306 ;
  assign n1308 = n148 & ~n1307 ;
  assign n1294 = ~x129 & n833 ;
  assign n1293 = x129 & n823 ;
  assign n1295 = n1294 ^ n1293 ;
  assign n1297 = ~x129 & ~n838 ;
  assign n1296 = x129 & ~n828 ;
  assign n1298 = n1297 ^ n1296 ;
  assign n1299 = ~n1295 & n1298 ;
  assign n1300 = n137 & ~n1299 ;
  assign n1309 = n1308 ^ n1300 ;
  assign n1319 = ~x129 & n846 ;
  assign n1318 = x129 & n860 ;
  assign n1320 = n1319 ^ n1318 ;
  assign n1322 = ~x129 & ~n851 ;
  assign n1321 = x129 & ~n865 ;
  assign n1323 = n1322 ^ n1321 ;
  assign n1324 = ~n1320 & n1323 ;
  assign n1325 = n171 & ~n1324 ;
  assign n1311 = ~x129 & n821 ;
  assign n1310 = x129 & n848 ;
  assign n1312 = n1311 ^ n1310 ;
  assign n1314 = ~x129 & ~n826 ;
  assign n1313 = x129 & ~n853 ;
  assign n1315 = n1314 ^ n1313 ;
  assign n1316 = ~n1312 & n1315 ;
  assign n1317 = n160 & ~n1316 ;
  assign n1326 = n1325 ^ n1317 ;
  assign n1327 = ~n1309 & ~n1326 ;
  assign n1328 = n254 & ~n1327 ;
  assign n1266 = ~x129 & n858 ;
  assign n1265 = x129 & n730 ;
  assign n1267 = n1266 ^ n1265 ;
  assign n1269 = ~x129 & ~n863 ;
  assign n1268 = x129 & ~n735 ;
  assign n1270 = n1269 ^ n1268 ;
  assign n1271 = ~n1267 & n1270 ;
  assign n1272 = n148 & ~n1271 ;
  assign n1258 = ~x129 & n728 ;
  assign n1257 = x129 & n718 ;
  assign n1259 = n1258 ^ n1257 ;
  assign n1261 = ~x129 & ~n733 ;
  assign n1260 = x129 & ~n723 ;
  assign n1262 = n1261 ^ n1260 ;
  assign n1263 = ~n1259 & n1262 ;
  assign n1264 = n137 & ~n1263 ;
  assign n1273 = n1272 ^ n1264 ;
  assign n1283 = ~x129 & n741 ;
  assign n1282 = x129 & n755 ;
  assign n1284 = n1283 ^ n1282 ;
  assign n1286 = ~x129 & ~n746 ;
  assign n1285 = x129 & ~n760 ;
  assign n1287 = n1286 ^ n1285 ;
  assign n1288 = ~n1284 & n1287 ;
  assign n1289 = n171 & ~n1288 ;
  assign n1275 = ~x129 & n716 ;
  assign n1274 = x129 & n743 ;
  assign n1276 = n1275 ^ n1274 ;
  assign n1278 = ~x129 & ~n721 ;
  assign n1277 = x129 & ~n748 ;
  assign n1279 = n1278 ^ n1277 ;
  assign n1280 = ~n1276 & n1279 ;
  assign n1281 = n160 & ~n1280 ;
  assign n1290 = n1289 ^ n1281 ;
  assign n1291 = ~n1273 & ~n1290 ;
  assign n1292 = n136 & ~n1291 ;
  assign n1329 = n1328 ^ n1292 ;
  assign n1375 = ~x129 & n545 ;
  assign n1374 = x129 & n887 ;
  assign n1376 = n1375 ^ n1374 ;
  assign n1378 = ~x129 & ~n550 ;
  assign n1377 = x129 & ~n892 ;
  assign n1379 = n1378 ^ n1377 ;
  assign n1380 = ~n1376 & n1379 ;
  assign n1381 = n148 & ~n1380 ;
  assign n1367 = ~x129 & n885 ;
  assign n1366 = x129 & n875 ;
  assign n1368 = n1367 ^ n1366 ;
  assign n1370 = ~x129 & ~n890 ;
  assign n1369 = x129 & ~n880 ;
  assign n1371 = n1370 ^ n1369 ;
  assign n1372 = ~n1368 & n1371 ;
  assign n1373 = n137 & ~n1372 ;
  assign n1382 = n1381 ^ n1373 ;
  assign n1392 = ~x129 & n898 ;
  assign n1391 = x129 & n912 ;
  assign n1393 = n1392 ^ n1391 ;
  assign n1395 = ~x129 & ~n903 ;
  assign n1394 = x129 & ~n917 ;
  assign n1396 = n1395 ^ n1394 ;
  assign n1397 = ~n1393 & n1396 ;
  assign n1398 = n171 & ~n1397 ;
  assign n1384 = ~x129 & n873 ;
  assign n1383 = x129 & n900 ;
  assign n1385 = n1384 ^ n1383 ;
  assign n1387 = ~x129 & ~n878 ;
  assign n1386 = x129 & ~n905 ;
  assign n1388 = n1387 ^ n1386 ;
  assign n1389 = ~n1385 & n1388 ;
  assign n1390 = n160 & ~n1389 ;
  assign n1399 = n1398 ^ n1390 ;
  assign n1400 = ~n1382 & ~n1399 ;
  assign n1401 = n279 & ~n1400 ;
  assign n1339 = ~x129 & n753 ;
  assign n1338 = x129 & n782 ;
  assign n1340 = n1339 ^ n1338 ;
  assign n1342 = ~x129 & ~n758 ;
  assign n1341 = x129 & ~n787 ;
  assign n1343 = n1342 ^ n1341 ;
  assign n1344 = ~n1340 & n1343 ;
  assign n1345 = n148 & ~n1344 ;
  assign n1331 = ~x129 & n780 ;
  assign n1330 = x129 & n770 ;
  assign n1332 = n1331 ^ n1330 ;
  assign n1334 = ~x129 & ~n785 ;
  assign n1333 = x129 & ~n775 ;
  assign n1335 = n1334 ^ n1333 ;
  assign n1336 = ~n1332 & n1335 ;
  assign n1337 = n137 & ~n1336 ;
  assign n1346 = n1345 ^ n1337 ;
  assign n1356 = ~x129 & n793 ;
  assign n1355 = x129 & n807 ;
  assign n1357 = n1356 ^ n1355 ;
  assign n1359 = ~x129 & ~n798 ;
  assign n1358 = x129 & ~n812 ;
  assign n1360 = n1359 ^ n1358 ;
  assign n1361 = ~n1357 & n1360 ;
  assign n1362 = n171 & ~n1361 ;
  assign n1348 = ~x129 & n768 ;
  assign n1347 = x129 & n795 ;
  assign n1349 = n1348 ^ n1347 ;
  assign n1351 = ~x129 & ~n773 ;
  assign n1350 = x129 & ~n800 ;
  assign n1352 = n1351 ^ n1350 ;
  assign n1353 = ~n1349 & n1352 ;
  assign n1354 = n160 & ~n1353 ;
  assign n1363 = n1362 ^ n1354 ;
  assign n1364 = ~n1346 & ~n1363 ;
  assign n1365 = n185 & ~n1364 ;
  assign n1402 = n1401 ^ n1365 ;
  assign n1403 = ~n1329 & ~n1402 ;
  assign n1404 = ~x134 & n1403 ;
  assign n1154 = ~x129 & n805 ;
  assign n1153 = x129 & n574 ;
  assign n1155 = n1154 ^ n1153 ;
  assign n1157 = ~x129 & ~n810 ;
  assign n1156 = x129 & ~n579 ;
  assign n1158 = n1157 ^ n1156 ;
  assign n1159 = ~n1155 & n1158 ;
  assign n1160 = n148 & ~n1159 ;
  assign n1146 = ~x129 & n572 ;
  assign n1145 = x129 & n562 ;
  assign n1147 = n1146 ^ n1145 ;
  assign n1149 = ~x129 & ~n577 ;
  assign n1148 = x129 & ~n567 ;
  assign n1150 = n1149 ^ n1148 ;
  assign n1151 = ~n1147 & n1150 ;
  assign n1152 = n137 & ~n1151 ;
  assign n1161 = n1160 ^ n1152 ;
  assign n1171 = ~x129 & n585 ;
  assign n1170 = x129 & n599 ;
  assign n1172 = n1171 ^ n1170 ;
  assign n1174 = ~x129 & ~n590 ;
  assign n1173 = x129 & ~n604 ;
  assign n1175 = n1174 ^ n1173 ;
  assign n1176 = ~n1172 & n1175 ;
  assign n1177 = n171 & ~n1176 ;
  assign n1163 = ~x129 & n560 ;
  assign n1162 = x129 & n587 ;
  assign n1164 = n1163 ^ n1162 ;
  assign n1166 = ~x129 & ~n565 ;
  assign n1165 = x129 & ~n592 ;
  assign n1167 = n1166 ^ n1165 ;
  assign n1168 = ~n1164 & n1167 ;
  assign n1169 = n160 & ~n1168 ;
  assign n1178 = n1177 ^ n1169 ;
  assign n1179 = ~n1161 & ~n1178 ;
  assign n1180 = n279 & ~n1179 ;
  assign n1112 = ~x129 & n597 ;
  assign n1111 = x129 & n677 ;
  assign n1113 = n1112 ^ n1111 ;
  assign n1115 = ~x129 & ~n602 ;
  assign n1114 = x129 & ~n682 ;
  assign n1116 = n1115 ^ n1114 ;
  assign n1117 = ~n1113 & n1116 ;
  assign n1118 = n148 & ~n1117 ;
  assign n1106 = ~x47 & ~x128 ;
  assign n1105 = ~x46 & x128 ;
  assign n1107 = n1106 ^ n1105 ;
  assign n1108 = ~x129 & n1107 ;
  assign n1104 = x129 & ~n671 ;
  assign n1109 = n1108 ^ n1104 ;
  assign n1110 = n137 & ~n1109 ;
  assign n1119 = n1118 ^ n1110 ;
  assign n1133 = x39 & ~x128 ;
  assign n1134 = ~x129 & n1133 ;
  assign n1132 = x129 & n700 ;
  assign n1135 = n1134 ^ n1132 ;
  assign n1137 = x38 & x128 ;
  assign n1138 = ~x129 & ~n1137 ;
  assign n1136 = x129 & ~n705 ;
  assign n1139 = n1138 ^ n1136 ;
  assign n1140 = ~n1135 & n1139 ;
  assign n1141 = n171 & ~n1140 ;
  assign n1122 = x43 & ~x128 ;
  assign n1123 = ~x129 & n1122 ;
  assign n1120 = x40 & x128 ;
  assign n1121 = x129 & n1120 ;
  assign n1124 = n1123 ^ n1121 ;
  assign n1127 = x42 & x128 ;
  assign n1128 = ~x129 & ~n1127 ;
  assign n1125 = x41 & ~x128 ;
  assign n1126 = x129 & ~n1125 ;
  assign n1129 = n1128 ^ n1126 ;
  assign n1130 = ~n1124 & n1129 ;
  assign n1131 = n160 & ~n1130 ;
  assign n1142 = n1141 ^ n1131 ;
  assign n1143 = ~n1119 & ~n1142 ;
  assign n1144 = n254 & ~n1143 ;
  assign n1181 = n1180 ^ n1144 ;
  assign n1227 = ~x129 & n650 ;
  assign n1226 = x129 & n522 ;
  assign n1228 = n1227 ^ n1226 ;
  assign n1230 = ~x129 & ~n655 ;
  assign n1229 = x129 & ~n527 ;
  assign n1231 = n1230 ^ n1229 ;
  assign n1232 = ~n1228 & n1231 ;
  assign n1233 = n148 & ~n1232 ;
  assign n1219 = ~x129 & n520 ;
  assign n1218 = x129 & n510 ;
  assign n1220 = n1219 ^ n1218 ;
  assign n1222 = ~x129 & ~n525 ;
  assign n1221 = x129 & ~n515 ;
  assign n1223 = n1222 ^ n1221 ;
  assign n1224 = ~n1220 & n1223 ;
  assign n1225 = n137 & ~n1224 ;
  assign n1234 = n1233 ^ n1225 ;
  assign n1244 = ~x129 & n533 ;
  assign n1243 = x129 & n547 ;
  assign n1245 = n1244 ^ n1243 ;
  assign n1247 = ~x129 & ~n538 ;
  assign n1246 = x129 & ~n552 ;
  assign n1248 = n1247 ^ n1246 ;
  assign n1249 = ~n1245 & n1248 ;
  assign n1250 = n171 & ~n1249 ;
  assign n1236 = ~x129 & n508 ;
  assign n1235 = x129 & n535 ;
  assign n1237 = n1236 ^ n1235 ;
  assign n1239 = ~x129 & ~n513 ;
  assign n1238 = x129 & ~n540 ;
  assign n1240 = n1239 ^ n1238 ;
  assign n1241 = ~n1237 & n1240 ;
  assign n1242 = n160 & ~n1241 ;
  assign n1251 = n1250 ^ n1242 ;
  assign n1252 = ~n1234 & ~n1251 ;
  assign n1253 = n185 & ~n1252 ;
  assign n1191 = ~x129 & n698 ;
  assign n1190 = x129 & n627 ;
  assign n1192 = n1191 ^ n1190 ;
  assign n1194 = ~x129 & ~n703 ;
  assign n1193 = x129 & ~n632 ;
  assign n1195 = n1194 ^ n1193 ;
  assign n1196 = ~n1192 & n1195 ;
  assign n1197 = n148 & ~n1196 ;
  assign n1183 = ~x129 & n625 ;
  assign n1182 = x129 & n615 ;
  assign n1184 = n1183 ^ n1182 ;
  assign n1186 = ~x129 & ~n630 ;
  assign n1185 = x129 & ~n620 ;
  assign n1187 = n1186 ^ n1185 ;
  assign n1188 = ~n1184 & n1187 ;
  assign n1189 = n137 & ~n1188 ;
  assign n1198 = n1197 ^ n1189 ;
  assign n1208 = ~x129 & n638 ;
  assign n1207 = x129 & n652 ;
  assign n1209 = n1208 ^ n1207 ;
  assign n1211 = ~x129 & ~n643 ;
  assign n1210 = x129 & ~n657 ;
  assign n1212 = n1211 ^ n1210 ;
  assign n1213 = ~n1209 & n1212 ;
  assign n1214 = n171 & ~n1213 ;
  assign n1200 = ~x129 & n613 ;
  assign n1199 = x129 & n640 ;
  assign n1201 = n1200 ^ n1199 ;
  assign n1203 = ~x129 & ~n618 ;
  assign n1202 = x129 & ~n645 ;
  assign n1204 = n1203 ^ n1202 ;
  assign n1205 = ~n1201 & n1204 ;
  assign n1206 = n160 & ~n1205 ;
  assign n1215 = n1214 ^ n1206 ;
  assign n1216 = ~n1198 & ~n1215 ;
  assign n1217 = n136 & ~n1216 ;
  assign n1254 = n1253 ^ n1217 ;
  assign n1255 = ~n1181 & ~n1254 ;
  assign n1256 = x134 & n1255 ;
  assign n1405 = n1404 ^ n1256 ;
  assign n1452 = n148 & n366 ;
  assign n1451 = n137 & n389 ;
  assign n1453 = n1452 ^ n1451 ;
  assign n1455 = n171 & n400 ;
  assign n1454 = n160 & n379 ;
  assign n1456 = n1455 ^ n1454 ;
  assign n1457 = ~n1453 & ~n1456 ;
  assign n1458 = n185 & ~n1457 ;
  assign n1444 = n148 & n455 ;
  assign n1443 = n137 & n345 ;
  assign n1445 = n1444 ^ n1443 ;
  assign n1447 = n171 & n356 ;
  assign n1446 = n160 & n335 ;
  assign n1448 = n1447 ^ n1446 ;
  assign n1449 = ~n1445 & ~n1448 ;
  assign n1450 = n136 & ~n1449 ;
  assign n1459 = n1458 ^ n1450 ;
  assign n1469 = n148 & n225 ;
  assign n1468 = n137 & n478 ;
  assign n1470 = n1469 ^ n1468 ;
  assign n1472 = n171 & n489 ;
  assign n1471 = n160 & n468 ;
  assign n1473 = n1472 ^ n1471 ;
  assign n1474 = ~n1470 & ~n1473 ;
  assign n1475 = n279 & ~n1474 ;
  assign n1461 = n148 & n499 ;
  assign n1460 = n137 & n434 ;
  assign n1462 = n1461 ^ n1460 ;
  assign n1464 = n171 & n445 ;
  assign n1463 = n160 & n424 ;
  assign n1465 = n1464 ^ n1463 ;
  assign n1466 = ~n1462 & ~n1465 ;
  assign n1467 = n254 & ~n1466 ;
  assign n1476 = n1475 ^ n1467 ;
  assign n1477 = ~n1459 & ~n1476 ;
  assign n1478 = ~x134 & n1477 ;
  assign n1415 = n171 & ~n241 ;
  assign n1414 = n160 & n263 ;
  assign n1416 = n1415 ^ n1414 ;
  assign n1418 = n148 & n319 ;
  assign n1417 = n137 & n273 ;
  assign n1419 = n1418 ^ n1417 ;
  assign n1420 = n254 & ~n1419 ;
  assign n1421 = ~n1416 & n1420 ;
  assign n1407 = n148 & n410 ;
  assign n1406 = n137 & n298 ;
  assign n1408 = n1407 ^ n1406 ;
  assign n1410 = n171 & n309 ;
  assign n1409 = n160 & n288 ;
  assign n1411 = n1410 ^ n1409 ;
  assign n1412 = ~n1408 & ~n1411 ;
  assign n1413 = n279 & n1412 ;
  assign n1422 = n1421 ^ n1413 ;
  assign n1423 = n1422 ^ x133 ;
  assign n1433 = n148 & n251 ;
  assign n1432 = n137 & n157 ;
  assign n1434 = n1433 ^ n1432 ;
  assign n1436 = n169 & n171 ;
  assign n1435 = n146 & n160 ;
  assign n1437 = n1436 ^ n1435 ;
  assign n1438 = ~n1434 & ~n1437 ;
  assign n1439 = n136 & ~n1438 ;
  assign n1425 = n148 & n180 ;
  assign n1424 = n137 & n204 ;
  assign n1426 = n1425 ^ n1424 ;
  assign n1428 = n171 & n215 ;
  assign n1427 = n160 & n194 ;
  assign n1429 = n1428 ^ n1427 ;
  assign n1430 = ~n1426 & ~n1429 ;
  assign n1431 = n185 & ~n1430 ;
  assign n1440 = n1439 ^ n1431 ;
  assign n1441 = n1423 & ~n1440 ;
  assign n1442 = x134 & n1441 ;
  assign n1479 = n1478 ^ n1442 ;
  assign n1525 = n148 & ~n763 ;
  assign n1524 = n137 & ~n790 ;
  assign n1526 = n1525 ^ n1524 ;
  assign n1528 = n171 & ~n803 ;
  assign n1527 = n160 & ~n778 ;
  assign n1529 = n1528 ^ n1527 ;
  assign n1530 = ~n1526 & ~n1529 ;
  assign n1531 = n185 & ~n1530 ;
  assign n1517 = n148 & ~n868 ;
  assign n1516 = n137 & ~n738 ;
  assign n1518 = n1517 ^ n1516 ;
  assign n1520 = n171 & ~n751 ;
  assign n1519 = n160 & ~n726 ;
  assign n1521 = n1520 ^ n1519 ;
  assign n1522 = ~n1518 & ~n1521 ;
  assign n1523 = n136 & ~n1522 ;
  assign n1532 = n1531 ^ n1523 ;
  assign n1542 = n148 & ~n555 ;
  assign n1541 = n137 & ~n895 ;
  assign n1543 = n1542 ^ n1541 ;
  assign n1545 = n171 & ~n908 ;
  assign n1544 = n160 & ~n883 ;
  assign n1546 = n1545 ^ n1544 ;
  assign n1547 = ~n1543 & ~n1546 ;
  assign n1548 = n279 & ~n1547 ;
  assign n1534 = n148 & ~n920 ;
  assign n1533 = n137 & ~n843 ;
  assign n1535 = n1534 ^ n1533 ;
  assign n1537 = n171 & ~n856 ;
  assign n1536 = n160 & ~n831 ;
  assign n1538 = n1537 ^ n1536 ;
  assign n1539 = ~n1535 & ~n1538 ;
  assign n1540 = n254 & ~n1539 ;
  assign n1549 = n1548 ^ n1540 ;
  assign n1550 = ~n1532 & ~n1549 ;
  assign n1551 = ~x134 & n1550 ;
  assign n1489 = n148 & ~n607 ;
  assign n1488 = n137 & ~n685 ;
  assign n1490 = n1489 ^ n1488 ;
  assign n1492 = n171 & ~n696 ;
  assign n1491 = n160 & ~n673 ;
  assign n1493 = n1492 ^ n1491 ;
  assign n1494 = ~n1490 & ~n1493 ;
  assign n1495 = n254 & ~n1494 ;
  assign n1481 = n148 & ~n815 ;
  assign n1480 = n137 & ~n582 ;
  assign n1482 = n1481 ^ n1480 ;
  assign n1484 = n171 & ~n595 ;
  assign n1483 = n160 & ~n570 ;
  assign n1485 = n1484 ^ n1483 ;
  assign n1486 = ~n1482 & ~n1485 ;
  assign n1487 = n279 & ~n1486 ;
  assign n1496 = n1495 ^ n1487 ;
  assign n1506 = n148 & ~n708 ;
  assign n1505 = n137 & ~n635 ;
  assign n1507 = n1506 ^ n1505 ;
  assign n1509 = n171 & ~n648 ;
  assign n1508 = n160 & ~n623 ;
  assign n1510 = n1509 ^ n1508 ;
  assign n1511 = ~n1507 & ~n1510 ;
  assign n1512 = n136 & ~n1511 ;
  assign n1498 = n148 & ~n660 ;
  assign n1497 = n137 & ~n530 ;
  assign n1499 = n1498 ^ n1497 ;
  assign n1501 = n171 & ~n543 ;
  assign n1500 = n160 & ~n518 ;
  assign n1502 = n1501 ^ n1500 ;
  assign n1503 = ~n1499 & ~n1502 ;
  assign n1504 = n185 & ~n1503 ;
  assign n1513 = n1512 ^ n1504 ;
  assign n1514 = ~n1496 & ~n1513 ;
  assign n1515 = x134 & n1514 ;
  assign n1552 = n1551 ^ n1515 ;
  assign n1598 = n148 & n1034 ;
  assign n1597 = n137 & n1045 ;
  assign n1599 = n1598 ^ n1597 ;
  assign n1601 = n171 & n1050 ;
  assign n1600 = n160 & n1041 ;
  assign n1602 = n1601 ^ n1600 ;
  assign n1603 = ~n1599 & ~n1602 ;
  assign n1604 = n185 & ~n1603 ;
  assign n1590 = n148 & n1075 ;
  assign n1589 = n137 & n1025 ;
  assign n1591 = n1590 ^ n1589 ;
  assign n1593 = n171 & n1030 ;
  assign n1592 = n160 & n1021 ;
  assign n1594 = n1593 ^ n1592 ;
  assign n1595 = ~n1591 & ~n1594 ;
  assign n1596 = n136 & ~n1595 ;
  assign n1605 = n1604 ^ n1596 ;
  assign n1615 = n148 & n944 ;
  assign n1614 = n137 & n1086 ;
  assign n1616 = n1615 ^ n1614 ;
  assign n1618 = n171 & n1091 ;
  assign n1617 = n160 & n1082 ;
  assign n1619 = n1618 ^ n1617 ;
  assign n1620 = ~n1616 & ~n1619 ;
  assign n1621 = n279 & ~n1620 ;
  assign n1607 = n148 & n1095 ;
  assign n1606 = n137 & n1066 ;
  assign n1608 = n1607 ^ n1606 ;
  assign n1610 = n171 & n1071 ;
  assign n1609 = n160 & n1062 ;
  assign n1611 = n1610 ^ n1609 ;
  assign n1612 = ~n1608 & ~n1611 ;
  assign n1613 = n254 & ~n1612 ;
  assign n1622 = n1621 ^ n1613 ;
  assign n1623 = ~n1605 & ~n1622 ;
  assign n1624 = ~x134 & n1623 ;
  assign n1562 = n148 & n964 ;
  assign n1561 = n137 & n996 ;
  assign n1563 = n1562 ^ n1561 ;
  assign n1565 = n171 & ~n1004 ;
  assign n1564 = n160 & n992 ;
  assign n1566 = n1565 ^ n1564 ;
  assign n1567 = ~n1563 & ~n1566 ;
  assign n1568 = n254 & ~n1567 ;
  assign n1554 = n148 & n1054 ;
  assign n1553 = n137 & n955 ;
  assign n1555 = n1554 ^ n1553 ;
  assign n1557 = n171 & n960 ;
  assign n1556 = n160 & n951 ;
  assign n1558 = n1557 ^ n1556 ;
  assign n1559 = ~n1555 & ~n1558 ;
  assign n1560 = n279 & ~n1559 ;
  assign n1569 = n1568 ^ n1560 ;
  assign n1579 = n148 & ~n1011 ;
  assign n1578 = n137 & n976 ;
  assign n1580 = n1579 ^ n1578 ;
  assign n1582 = n171 & n981 ;
  assign n1581 = n160 & n972 ;
  assign n1583 = n1582 ^ n1581 ;
  assign n1584 = ~n1580 & ~n1583 ;
  assign n1585 = n136 & ~n1584 ;
  assign n1571 = n148 & n985 ;
  assign n1570 = n137 & n935 ;
  assign n1572 = n1571 ^ n1570 ;
  assign n1574 = n171 & n940 ;
  assign n1573 = n160 & n931 ;
  assign n1575 = n1574 ^ n1573 ;
  assign n1576 = ~n1572 & ~n1575 ;
  assign n1577 = n185 & ~n1576 ;
  assign n1586 = n1585 ^ n1577 ;
  assign n1587 = ~n1569 & ~n1586 ;
  assign n1588 = x134 & n1587 ;
  assign n1625 = n1624 ^ n1588 ;
  assign n1671 = n148 & ~n1288 ;
  assign n1670 = n137 & ~n1344 ;
  assign n1672 = n1671 ^ n1670 ;
  assign n1674 = n171 & ~n1353 ;
  assign n1673 = n160 & ~n1336 ;
  assign n1675 = n1674 ^ n1673 ;
  assign n1676 = ~n1672 & ~n1675 ;
  assign n1677 = n185 & ~n1676 ;
  assign n1663 = n148 & ~n1324 ;
  assign n1662 = n137 & ~n1271 ;
  assign n1664 = n1663 ^ n1662 ;
  assign n1666 = n171 & ~n1280 ;
  assign n1665 = n160 & ~n1263 ;
  assign n1667 = n1666 ^ n1665 ;
  assign n1668 = ~n1664 & ~n1667 ;
  assign n1669 = n136 & ~n1668 ;
  assign n1678 = n1677 ^ n1669 ;
  assign n1688 = n148 & ~n1249 ;
  assign n1687 = n137 & ~n1380 ;
  assign n1689 = n1688 ^ n1687 ;
  assign n1691 = n171 & ~n1389 ;
  assign n1690 = n160 & ~n1372 ;
  assign n1692 = n1691 ^ n1690 ;
  assign n1693 = ~n1689 & ~n1692 ;
  assign n1694 = n279 & ~n1693 ;
  assign n1680 = n148 & ~n1397 ;
  assign n1679 = n137 & ~n1307 ;
  assign n1681 = n1680 ^ n1679 ;
  assign n1683 = n171 & ~n1316 ;
  assign n1682 = n160 & ~n1299 ;
  assign n1684 = n1683 ^ n1682 ;
  assign n1685 = ~n1681 & ~n1684 ;
  assign n1686 = n254 & ~n1685 ;
  assign n1695 = n1694 ^ n1686 ;
  assign n1696 = ~n1678 & ~n1695 ;
  assign n1697 = ~x134 & n1696 ;
  assign n1635 = n137 & ~n1117 ;
  assign n1634 = n160 & ~n1109 ;
  assign n1636 = n1635 ^ n1634 ;
  assign n1638 = n171 & ~n1130 ;
  assign n1637 = n148 & ~n1176 ;
  assign n1639 = n1638 ^ n1637 ;
  assign n1640 = ~n1636 & ~n1639 ;
  assign n1641 = n254 & ~n1640 ;
  assign n1627 = n148 & ~n1361 ;
  assign n1626 = n137 & ~n1159 ;
  assign n1628 = n1627 ^ n1626 ;
  assign n1630 = n171 & ~n1168 ;
  assign n1629 = n160 & ~n1151 ;
  assign n1631 = n1630 ^ n1629 ;
  assign n1632 = ~n1628 & ~n1631 ;
  assign n1633 = n279 & ~n1632 ;
  assign n1642 = n1641 ^ n1633 ;
  assign n1652 = n148 & ~n1140 ;
  assign n1651 = n137 & ~n1196 ;
  assign n1653 = n1652 ^ n1651 ;
  assign n1655 = n171 & ~n1205 ;
  assign n1654 = n160 & ~n1188 ;
  assign n1656 = n1655 ^ n1654 ;
  assign n1657 = ~n1653 & ~n1656 ;
  assign n1658 = n136 & ~n1657 ;
  assign n1644 = n148 & ~n1213 ;
  assign n1643 = n137 & ~n1232 ;
  assign n1645 = n1644 ^ n1643 ;
  assign n1647 = n171 & ~n1241 ;
  assign n1646 = n160 & ~n1224 ;
  assign n1648 = n1647 ^ n1646 ;
  assign n1649 = ~n1645 & ~n1648 ;
  assign n1650 = n185 & ~n1649 ;
  assign n1659 = n1658 ^ n1650 ;
  assign n1660 = ~n1642 & ~n1659 ;
  assign n1661 = x134 & n1660 ;
  assign n1698 = n1697 ^ n1661 ;
  assign n1745 = n148 & n356 ;
  assign n1744 = n137 & n366 ;
  assign n1746 = n1745 ^ n1744 ;
  assign n1748 = n171 & n379 ;
  assign n1747 = n160 & n389 ;
  assign n1749 = n1748 ^ n1747 ;
  assign n1750 = ~n1746 & ~n1749 ;
  assign n1751 = n185 & ~n1750 ;
  assign n1737 = n148 & n445 ;
  assign n1736 = n137 & n455 ;
  assign n1738 = n1737 ^ n1736 ;
  assign n1740 = n171 & n335 ;
  assign n1739 = n160 & n345 ;
  assign n1741 = n1740 ^ n1739 ;
  assign n1742 = ~n1738 & ~n1741 ;
  assign n1743 = n136 & ~n1742 ;
  assign n1752 = n1751 ^ n1743 ;
  assign n1762 = n148 & n215 ;
  assign n1761 = n137 & n225 ;
  assign n1763 = n1762 ^ n1761 ;
  assign n1765 = n171 & n468 ;
  assign n1764 = n160 & n478 ;
  assign n1766 = n1765 ^ n1764 ;
  assign n1767 = ~n1763 & ~n1766 ;
  assign n1768 = n279 & ~n1767 ;
  assign n1754 = n148 & n489 ;
  assign n1753 = n137 & n499 ;
  assign n1755 = n1754 ^ n1753 ;
  assign n1757 = n171 & n424 ;
  assign n1756 = n160 & n434 ;
  assign n1758 = n1757 ^ n1756 ;
  assign n1759 = ~n1755 & ~n1758 ;
  assign n1760 = n254 & ~n1759 ;
  assign n1769 = n1768 ^ n1760 ;
  assign n1770 = ~n1752 & ~n1769 ;
  assign n1771 = ~x134 & n1770 ;
  assign n1708 = n148 & n309 ;
  assign n1707 = n137 & n319 ;
  assign n1709 = n1708 ^ n1707 ;
  assign n1711 = n171 & n263 ;
  assign n1710 = n160 & n273 ;
  assign n1712 = n1711 ^ n1710 ;
  assign n1713 = ~n1709 & ~n1712 ;
  assign n1714 = n254 & ~n1713 ;
  assign n1700 = n148 & n400 ;
  assign n1699 = n137 & n410 ;
  assign n1701 = n1700 ^ n1699 ;
  assign n1703 = n171 & n288 ;
  assign n1702 = n160 & n298 ;
  assign n1704 = n1703 ^ n1702 ;
  assign n1705 = ~n1701 & ~n1704 ;
  assign n1706 = n279 & ~n1705 ;
  assign n1715 = n1714 ^ n1706 ;
  assign n1726 = n148 & n169 ;
  assign n1725 = n137 & n180 ;
  assign n1727 = n1726 ^ n1725 ;
  assign n1729 = n171 & n194 ;
  assign n1728 = n160 & n204 ;
  assign n1730 = n1729 ^ n1728 ;
  assign n1731 = ~n1727 & ~n1730 ;
  assign n1732 = n185 & n1731 ;
  assign n1717 = n148 & ~n241 ;
  assign n1716 = n137 & n251 ;
  assign n1718 = n1717 ^ n1716 ;
  assign n1720 = n146 & n171 ;
  assign n1719 = n157 & n160 ;
  assign n1721 = n1720 ^ n1719 ;
  assign n1722 = n136 & ~n1721 ;
  assign n1723 = ~n1718 & n1722 ;
  assign n1724 = n1723 ^ x133 ;
  assign n1733 = n1732 ^ n1724 ;
  assign n1734 = ~n1715 & ~n1733 ;
  assign n1735 = x134 & n1734 ;
  assign n1772 = n1771 ^ n1735 ;
  assign n1818 = n148 & ~n751 ;
  assign n1817 = n137 & ~n763 ;
  assign n1819 = n1818 ^ n1817 ;
  assign n1821 = n171 & ~n778 ;
  assign n1820 = n160 & ~n790 ;
  assign n1822 = n1821 ^ n1820 ;
  assign n1823 = ~n1819 & ~n1822 ;
  assign n1824 = n185 & ~n1823 ;
  assign n1810 = n148 & ~n856 ;
  assign n1809 = n137 & ~n868 ;
  assign n1811 = n1810 ^ n1809 ;
  assign n1813 = n171 & ~n726 ;
  assign n1812 = n160 & ~n738 ;
  assign n1814 = n1813 ^ n1812 ;
  assign n1815 = ~n1811 & ~n1814 ;
  assign n1816 = n136 & ~n1815 ;
  assign n1825 = n1824 ^ n1816 ;
  assign n1835 = n148 & ~n543 ;
  assign n1834 = n137 & ~n555 ;
  assign n1836 = n1835 ^ n1834 ;
  assign n1838 = n171 & ~n883 ;
  assign n1837 = n160 & ~n895 ;
  assign n1839 = n1838 ^ n1837 ;
  assign n1840 = ~n1836 & ~n1839 ;
  assign n1841 = n279 & ~n1840 ;
  assign n1827 = n148 & ~n908 ;
  assign n1826 = n137 & ~n920 ;
  assign n1828 = n1827 ^ n1826 ;
  assign n1830 = n171 & ~n831 ;
  assign n1829 = n160 & ~n843 ;
  assign n1831 = n1830 ^ n1829 ;
  assign n1832 = ~n1828 & ~n1831 ;
  assign n1833 = n254 & ~n1832 ;
  assign n1842 = n1841 ^ n1833 ;
  assign n1843 = ~n1825 & ~n1842 ;
  assign n1844 = ~x134 & n1843 ;
  assign n1782 = n148 & ~n595 ;
  assign n1781 = n137 & ~n607 ;
  assign n1783 = n1782 ^ n1781 ;
  assign n1785 = n171 & ~n673 ;
  assign n1784 = n160 & ~n685 ;
  assign n1786 = n1785 ^ n1784 ;
  assign n1787 = ~n1783 & ~n1786 ;
  assign n1788 = n254 & ~n1787 ;
  assign n1774 = n148 & ~n803 ;
  assign n1773 = n137 & ~n815 ;
  assign n1775 = n1774 ^ n1773 ;
  assign n1777 = n171 & ~n570 ;
  assign n1776 = n160 & ~n582 ;
  assign n1778 = n1777 ^ n1776 ;
  assign n1779 = ~n1775 & ~n1778 ;
  assign n1780 = n279 & ~n1779 ;
  assign n1789 = n1788 ^ n1780 ;
  assign n1799 = n148 & ~n696 ;
  assign n1798 = n137 & ~n708 ;
  assign n1800 = n1799 ^ n1798 ;
  assign n1802 = n171 & ~n623 ;
  assign n1801 = n160 & ~n635 ;
  assign n1803 = n1802 ^ n1801 ;
  assign n1804 = ~n1800 & ~n1803 ;
  assign n1805 = n136 & ~n1804 ;
  assign n1791 = n148 & ~n648 ;
  assign n1790 = n137 & ~n660 ;
  assign n1792 = n1791 ^ n1790 ;
  assign n1794 = n171 & ~n518 ;
  assign n1793 = n160 & ~n530 ;
  assign n1795 = n1794 ^ n1793 ;
  assign n1796 = ~n1792 & ~n1795 ;
  assign n1797 = n185 & ~n1796 ;
  assign n1806 = n1805 ^ n1797 ;
  assign n1807 = ~n1789 & ~n1806 ;
  assign n1808 = x134 & n1807 ;
  assign n1845 = n1844 ^ n1808 ;
  assign n1891 = n148 & n1030 ;
  assign n1890 = n137 & n1034 ;
  assign n1892 = n1891 ^ n1890 ;
  assign n1894 = n171 & n1041 ;
  assign n1893 = n160 & n1045 ;
  assign n1895 = n1894 ^ n1893 ;
  assign n1896 = ~n1892 & ~n1895 ;
  assign n1897 = n185 & ~n1896 ;
  assign n1883 = n148 & n1071 ;
  assign n1882 = n137 & n1075 ;
  assign n1884 = n1883 ^ n1882 ;
  assign n1886 = n171 & n1021 ;
  assign n1885 = n160 & n1025 ;
  assign n1887 = n1886 ^ n1885 ;
  assign n1888 = ~n1884 & ~n1887 ;
  assign n1889 = n136 & ~n1888 ;
  assign n1898 = n1897 ^ n1889 ;
  assign n1908 = n148 & n940 ;
  assign n1907 = n137 & n944 ;
  assign n1909 = n1908 ^ n1907 ;
  assign n1911 = n171 & n1082 ;
  assign n1910 = n160 & n1086 ;
  assign n1912 = n1911 ^ n1910 ;
  assign n1913 = ~n1909 & ~n1912 ;
  assign n1914 = n279 & ~n1913 ;
  assign n1900 = n148 & n1091 ;
  assign n1899 = n137 & n1095 ;
  assign n1901 = n1900 ^ n1899 ;
  assign n1903 = n171 & n1062 ;
  assign n1902 = n160 & n1066 ;
  assign n1904 = n1903 ^ n1902 ;
  assign n1905 = ~n1901 & ~n1904 ;
  assign n1906 = n254 & ~n1905 ;
  assign n1915 = n1914 ^ n1906 ;
  assign n1916 = ~n1898 & ~n1915 ;
  assign n1917 = ~x134 & n1916 ;
  assign n1855 = n148 & n960 ;
  assign n1854 = n137 & n964 ;
  assign n1856 = n1855 ^ n1854 ;
  assign n1858 = n171 & n992 ;
  assign n1857 = n160 & n996 ;
  assign n1859 = n1858 ^ n1857 ;
  assign n1860 = ~n1856 & ~n1859 ;
  assign n1861 = n254 & ~n1860 ;
  assign n1847 = n148 & n1050 ;
  assign n1846 = n137 & n1054 ;
  assign n1848 = n1847 ^ n1846 ;
  assign n1850 = n171 & n951 ;
  assign n1849 = n160 & n955 ;
  assign n1851 = n1850 ^ n1849 ;
  assign n1852 = ~n1848 & ~n1851 ;
  assign n1853 = n279 & ~n1852 ;
  assign n1862 = n1861 ^ n1853 ;
  assign n1872 = n148 & ~n1004 ;
  assign n1871 = n137 & ~n1011 ;
  assign n1873 = n1872 ^ n1871 ;
  assign n1875 = n171 & n972 ;
  assign n1874 = n160 & n976 ;
  assign n1876 = n1875 ^ n1874 ;
  assign n1877 = ~n1873 & ~n1876 ;
  assign n1878 = n136 & ~n1877 ;
  assign n1864 = n148 & n981 ;
  assign n1863 = n137 & n985 ;
  assign n1865 = n1864 ^ n1863 ;
  assign n1867 = n171 & n931 ;
  assign n1866 = n160 & n935 ;
  assign n1868 = n1867 ^ n1866 ;
  assign n1869 = ~n1865 & ~n1868 ;
  assign n1870 = n185 & ~n1869 ;
  assign n1879 = n1878 ^ n1870 ;
  assign n1880 = ~n1862 & ~n1879 ;
  assign n1881 = x134 & n1880 ;
  assign n1918 = n1917 ^ n1881 ;
  assign n1964 = n148 & ~n1280 ;
  assign n1963 = n137 & ~n1288 ;
  assign n1965 = n1964 ^ n1963 ;
  assign n1967 = n171 & ~n1336 ;
  assign n1966 = n160 & ~n1344 ;
  assign n1968 = n1967 ^ n1966 ;
  assign n1969 = ~n1965 & ~n1968 ;
  assign n1970 = n185 & ~n1969 ;
  assign n1956 = n148 & ~n1316 ;
  assign n1955 = n137 & ~n1324 ;
  assign n1957 = n1956 ^ n1955 ;
  assign n1959 = n171 & ~n1263 ;
  assign n1958 = n160 & ~n1271 ;
  assign n1960 = n1959 ^ n1958 ;
  assign n1961 = ~n1957 & ~n1960 ;
  assign n1962 = n136 & ~n1961 ;
  assign n1971 = n1970 ^ n1962 ;
  assign n1981 = n148 & ~n1241 ;
  assign n1980 = n137 & ~n1249 ;
  assign n1982 = n1981 ^ n1980 ;
  assign n1984 = n171 & ~n1372 ;
  assign n1983 = n160 & ~n1380 ;
  assign n1985 = n1984 ^ n1983 ;
  assign n1986 = ~n1982 & ~n1985 ;
  assign n1987 = n279 & ~n1986 ;
  assign n1973 = n148 & ~n1389 ;
  assign n1972 = n137 & ~n1397 ;
  assign n1974 = n1973 ^ n1972 ;
  assign n1976 = n171 & ~n1299 ;
  assign n1975 = n160 & ~n1307 ;
  assign n1977 = n1976 ^ n1975 ;
  assign n1978 = ~n1974 & ~n1977 ;
  assign n1979 = n254 & ~n1978 ;
  assign n1988 = n1987 ^ n1979 ;
  assign n1989 = ~n1971 & ~n1988 ;
  assign n1990 = ~x134 & n1989 ;
  assign n1928 = n148 & ~n1168 ;
  assign n1927 = n160 & ~n1117 ;
  assign n1929 = n1928 ^ n1927 ;
  assign n1931 = n171 & ~n1109 ;
  assign n1930 = n137 & ~n1176 ;
  assign n1932 = n1931 ^ n1930 ;
  assign n1933 = ~n1929 & ~n1932 ;
  assign n1934 = n254 & ~n1933 ;
  assign n1920 = n148 & ~n1353 ;
  assign n1919 = n137 & ~n1361 ;
  assign n1921 = n1920 ^ n1919 ;
  assign n1923 = n171 & ~n1151 ;
  assign n1922 = n160 & ~n1159 ;
  assign n1924 = n1923 ^ n1922 ;
  assign n1925 = ~n1921 & ~n1924 ;
  assign n1926 = n279 & ~n1925 ;
  assign n1935 = n1934 ^ n1926 ;
  assign n1945 = n148 & ~n1130 ;
  assign n1944 = n137 & ~n1140 ;
  assign n1946 = n1945 ^ n1944 ;
  assign n1948 = n171 & ~n1188 ;
  assign n1947 = n160 & ~n1196 ;
  assign n1949 = n1948 ^ n1947 ;
  assign n1950 = ~n1946 & ~n1949 ;
  assign n1951 = n136 & ~n1950 ;
  assign n1937 = n148 & ~n1205 ;
  assign n1936 = n137 & ~n1213 ;
  assign n1938 = n1937 ^ n1936 ;
  assign n1940 = n171 & ~n1224 ;
  assign n1939 = n160 & ~n1232 ;
  assign n1941 = n1940 ^ n1939 ;
  assign n1942 = ~n1938 & ~n1941 ;
  assign n1943 = n185 & ~n1942 ;
  assign n1952 = n1951 ^ n1943 ;
  assign n1953 = ~n1935 & ~n1952 ;
  assign n1954 = x134 & n1953 ;
  assign n1991 = n1990 ^ n1954 ;
  assign n2038 = n148 & n335 ;
  assign n2037 = n137 & n356 ;
  assign n2039 = n2038 ^ n2037 ;
  assign n2041 = n171 & n389 ;
  assign n2040 = n160 & n366 ;
  assign n2042 = n2041 ^ n2040 ;
  assign n2043 = ~n2039 & ~n2042 ;
  assign n2044 = n185 & ~n2043 ;
  assign n2030 = n148 & n424 ;
  assign n2029 = n137 & n445 ;
  assign n2031 = n2030 ^ n2029 ;
  assign n2033 = n171 & n345 ;
  assign n2032 = n160 & n455 ;
  assign n2034 = n2033 ^ n2032 ;
  assign n2035 = ~n2031 & ~n2034 ;
  assign n2036 = n136 & ~n2035 ;
  assign n2045 = n2044 ^ n2036 ;
  assign n2055 = n148 & n194 ;
  assign n2054 = n137 & n215 ;
  assign n2056 = n2055 ^ n2054 ;
  assign n2058 = n171 & n478 ;
  assign n2057 = n160 & n225 ;
  assign n2059 = n2058 ^ n2057 ;
  assign n2060 = ~n2056 & ~n2059 ;
  assign n2061 = n279 & ~n2060 ;
  assign n2047 = n148 & n468 ;
  assign n2046 = n137 & n489 ;
  assign n2048 = n2047 ^ n2046 ;
  assign n2050 = n171 & n434 ;
  assign n2049 = n160 & n499 ;
  assign n2051 = n2050 ^ n2049 ;
  assign n2052 = ~n2048 & ~n2051 ;
  assign n2053 = n254 & ~n2052 ;
  assign n2062 = n2061 ^ n2053 ;
  assign n2063 = ~n2045 & ~n2062 ;
  assign n2064 = ~x134 & n2063 ;
  assign n2001 = n148 & n288 ;
  assign n2000 = n137 & n309 ;
  assign n2002 = n2001 ^ n2000 ;
  assign n2004 = n171 & n273 ;
  assign n2003 = n160 & n319 ;
  assign n2005 = n2004 ^ n2003 ;
  assign n2006 = ~n2002 & ~n2005 ;
  assign n2007 = n254 & ~n2006 ;
  assign n1993 = n148 & n379 ;
  assign n1992 = n137 & n400 ;
  assign n1994 = n1993 ^ n1992 ;
  assign n1996 = n171 & n298 ;
  assign n1995 = n160 & n410 ;
  assign n1997 = n1996 ^ n1995 ;
  assign n1998 = ~n1994 & ~n1997 ;
  assign n1999 = n279 & ~n1998 ;
  assign n2008 = n2007 ^ n1999 ;
  assign n2019 = n146 & n148 ;
  assign n2018 = n137 & n169 ;
  assign n2020 = n2019 ^ n2018 ;
  assign n2022 = n171 & n204 ;
  assign n2021 = n160 & n180 ;
  assign n2023 = n2022 ^ n2021 ;
  assign n2024 = ~n2020 & ~n2023 ;
  assign n2025 = n185 & n2024 ;
  assign n2010 = n148 & n263 ;
  assign n2009 = n137 & ~n241 ;
  assign n2011 = n2010 ^ n2009 ;
  assign n2013 = n157 & n171 ;
  assign n2012 = n160 & n251 ;
  assign n2014 = n2013 ^ n2012 ;
  assign n2015 = n136 & ~n2014 ;
  assign n2016 = ~n2011 & n2015 ;
  assign n2017 = n2016 ^ x133 ;
  assign n2026 = n2025 ^ n2017 ;
  assign n2027 = ~n2008 & ~n2026 ;
  assign n2028 = x134 & n2027 ;
  assign n2065 = n2064 ^ n2028 ;
  assign n2111 = n148 & ~n726 ;
  assign n2110 = n137 & ~n751 ;
  assign n2112 = n2111 ^ n2110 ;
  assign n2114 = n171 & ~n790 ;
  assign n2113 = n160 & ~n763 ;
  assign n2115 = n2114 ^ n2113 ;
  assign n2116 = ~n2112 & ~n2115 ;
  assign n2117 = n185 & ~n2116 ;
  assign n2103 = n148 & ~n831 ;
  assign n2102 = n137 & ~n856 ;
  assign n2104 = n2103 ^ n2102 ;
  assign n2106 = n171 & ~n738 ;
  assign n2105 = n160 & ~n868 ;
  assign n2107 = n2106 ^ n2105 ;
  assign n2108 = ~n2104 & ~n2107 ;
  assign n2109 = n136 & ~n2108 ;
  assign n2118 = n2117 ^ n2109 ;
  assign n2128 = n148 & ~n518 ;
  assign n2127 = n137 & ~n543 ;
  assign n2129 = n2128 ^ n2127 ;
  assign n2131 = n171 & ~n895 ;
  assign n2130 = n160 & ~n555 ;
  assign n2132 = n2131 ^ n2130 ;
  assign n2133 = ~n2129 & ~n2132 ;
  assign n2134 = n279 & ~n2133 ;
  assign n2120 = n148 & ~n883 ;
  assign n2119 = n137 & ~n908 ;
  assign n2121 = n2120 ^ n2119 ;
  assign n2123 = n171 & ~n843 ;
  assign n2122 = n160 & ~n920 ;
  assign n2124 = n2123 ^ n2122 ;
  assign n2125 = ~n2121 & ~n2124 ;
  assign n2126 = n254 & ~n2125 ;
  assign n2135 = n2134 ^ n2126 ;
  assign n2136 = ~n2118 & ~n2135 ;
  assign n2137 = ~x134 & n2136 ;
  assign n2075 = n148 & ~n570 ;
  assign n2074 = n137 & ~n595 ;
  assign n2076 = n2075 ^ n2074 ;
  assign n2078 = n171 & ~n685 ;
  assign n2077 = n160 & ~n607 ;
  assign n2079 = n2078 ^ n2077 ;
  assign n2080 = ~n2076 & ~n2079 ;
  assign n2081 = n254 & ~n2080 ;
  assign n2067 = n148 & ~n778 ;
  assign n2066 = n137 & ~n803 ;
  assign n2068 = n2067 ^ n2066 ;
  assign n2070 = n171 & ~n582 ;
  assign n2069 = n160 & ~n815 ;
  assign n2071 = n2070 ^ n2069 ;
  assign n2072 = ~n2068 & ~n2071 ;
  assign n2073 = n279 & ~n2072 ;
  assign n2082 = n2081 ^ n2073 ;
  assign n2092 = n148 & ~n673 ;
  assign n2091 = n137 & ~n696 ;
  assign n2093 = n2092 ^ n2091 ;
  assign n2095 = n171 & ~n635 ;
  assign n2094 = n160 & ~n708 ;
  assign n2096 = n2095 ^ n2094 ;
  assign n2097 = ~n2093 & ~n2096 ;
  assign n2098 = n136 & ~n2097 ;
  assign n2084 = n148 & ~n623 ;
  assign n2083 = n137 & ~n648 ;
  assign n2085 = n2084 ^ n2083 ;
  assign n2087 = n171 & ~n530 ;
  assign n2086 = n160 & ~n660 ;
  assign n2088 = n2087 ^ n2086 ;
  assign n2089 = ~n2085 & ~n2088 ;
  assign n2090 = n185 & ~n2089 ;
  assign n2099 = n2098 ^ n2090 ;
  assign n2100 = ~n2082 & ~n2099 ;
  assign n2101 = x134 & n2100 ;
  assign n2138 = n2137 ^ n2101 ;
  assign n2184 = n148 & n1021 ;
  assign n2183 = n137 & n1030 ;
  assign n2185 = n2184 ^ n2183 ;
  assign n2187 = n171 & n1045 ;
  assign n2186 = n160 & n1034 ;
  assign n2188 = n2187 ^ n2186 ;
  assign n2189 = ~n2185 & ~n2188 ;
  assign n2190 = n185 & ~n2189 ;
  assign n2176 = n148 & n1062 ;
  assign n2175 = n137 & n1071 ;
  assign n2177 = n2176 ^ n2175 ;
  assign n2179 = n171 & n1025 ;
  assign n2178 = n160 & n1075 ;
  assign n2180 = n2179 ^ n2178 ;
  assign n2181 = ~n2177 & ~n2180 ;
  assign n2182 = n136 & ~n2181 ;
  assign n2191 = n2190 ^ n2182 ;
  assign n2201 = n148 & n931 ;
  assign n2200 = n137 & n940 ;
  assign n2202 = n2201 ^ n2200 ;
  assign n2204 = n171 & n1086 ;
  assign n2203 = n160 & n944 ;
  assign n2205 = n2204 ^ n2203 ;
  assign n2206 = ~n2202 & ~n2205 ;
  assign n2207 = n279 & ~n2206 ;
  assign n2193 = n148 & n1082 ;
  assign n2192 = n137 & n1091 ;
  assign n2194 = n2193 ^ n2192 ;
  assign n2196 = n171 & n1066 ;
  assign n2195 = n160 & n1095 ;
  assign n2197 = n2196 ^ n2195 ;
  assign n2198 = ~n2194 & ~n2197 ;
  assign n2199 = n254 & ~n2198 ;
  assign n2208 = n2207 ^ n2199 ;
  assign n2209 = ~n2191 & ~n2208 ;
  assign n2210 = ~x134 & n2209 ;
  assign n2148 = n148 & n951 ;
  assign n2147 = n137 & n960 ;
  assign n2149 = n2148 ^ n2147 ;
  assign n2151 = n171 & n996 ;
  assign n2150 = n160 & n964 ;
  assign n2152 = n2151 ^ n2150 ;
  assign n2153 = ~n2149 & ~n2152 ;
  assign n2154 = n254 & ~n2153 ;
  assign n2140 = n148 & n1041 ;
  assign n2139 = n137 & n1050 ;
  assign n2141 = n2140 ^ n2139 ;
  assign n2143 = n171 & n955 ;
  assign n2142 = n160 & n1054 ;
  assign n2144 = n2143 ^ n2142 ;
  assign n2145 = ~n2141 & ~n2144 ;
  assign n2146 = n279 & ~n2145 ;
  assign n2155 = n2154 ^ n2146 ;
  assign n2165 = n148 & n992 ;
  assign n2164 = n137 & ~n1004 ;
  assign n2166 = n2165 ^ n2164 ;
  assign n2168 = n171 & n976 ;
  assign n2167 = n160 & ~n1011 ;
  assign n2169 = n2168 ^ n2167 ;
  assign n2170 = ~n2166 & ~n2169 ;
  assign n2171 = n136 & ~n2170 ;
  assign n2157 = n148 & n972 ;
  assign n2156 = n137 & n981 ;
  assign n2158 = n2157 ^ n2156 ;
  assign n2160 = n171 & n935 ;
  assign n2159 = n160 & n985 ;
  assign n2161 = n2160 ^ n2159 ;
  assign n2162 = ~n2158 & ~n2161 ;
  assign n2163 = n185 & ~n2162 ;
  assign n2172 = n2171 ^ n2163 ;
  assign n2173 = ~n2155 & ~n2172 ;
  assign n2174 = x134 & n2173 ;
  assign n2211 = n2210 ^ n2174 ;
  assign n2257 = n148 & ~n1263 ;
  assign n2256 = n137 & ~n1280 ;
  assign n2258 = n2257 ^ n2256 ;
  assign n2260 = n171 & ~n1344 ;
  assign n2259 = n160 & ~n1288 ;
  assign n2261 = n2260 ^ n2259 ;
  assign n2262 = ~n2258 & ~n2261 ;
  assign n2263 = n185 & ~n2262 ;
  assign n2249 = n148 & ~n1299 ;
  assign n2248 = n137 & ~n1316 ;
  assign n2250 = n2249 ^ n2248 ;
  assign n2252 = n171 & ~n1271 ;
  assign n2251 = n160 & ~n1324 ;
  assign n2253 = n2252 ^ n2251 ;
  assign n2254 = ~n2250 & ~n2253 ;
  assign n2255 = n136 & ~n2254 ;
  assign n2264 = n2263 ^ n2255 ;
  assign n2274 = n148 & ~n1224 ;
  assign n2273 = n137 & ~n1241 ;
  assign n2275 = n2274 ^ n2273 ;
  assign n2277 = n171 & ~n1380 ;
  assign n2276 = n160 & ~n1249 ;
  assign n2278 = n2277 ^ n2276 ;
  assign n2279 = ~n2275 & ~n2278 ;
  assign n2280 = n279 & ~n2279 ;
  assign n2266 = n148 & ~n1372 ;
  assign n2265 = n137 & ~n1389 ;
  assign n2267 = n2266 ^ n2265 ;
  assign n2269 = n171 & ~n1307 ;
  assign n2268 = n160 & ~n1397 ;
  assign n2270 = n2269 ^ n2268 ;
  assign n2271 = ~n2267 & ~n2270 ;
  assign n2272 = n254 & ~n2271 ;
  assign n2281 = n2280 ^ n2272 ;
  assign n2282 = ~n2264 & ~n2281 ;
  assign n2283 = ~x134 & n2282 ;
  assign n2221 = n148 & ~n1151 ;
  assign n2220 = n137 & ~n1168 ;
  assign n2222 = n2221 ^ n2220 ;
  assign n2224 = n171 & ~n1117 ;
  assign n2223 = n160 & ~n1176 ;
  assign n2225 = n2224 ^ n2223 ;
  assign n2226 = ~n2222 & ~n2225 ;
  assign n2227 = n254 & ~n2226 ;
  assign n2213 = n148 & ~n1336 ;
  assign n2212 = n137 & ~n1353 ;
  assign n2214 = n2213 ^ n2212 ;
  assign n2216 = n171 & ~n1159 ;
  assign n2215 = n160 & ~n1361 ;
  assign n2217 = n2216 ^ n2215 ;
  assign n2218 = ~n2214 & ~n2217 ;
  assign n2219 = n279 & ~n2218 ;
  assign n2228 = n2227 ^ n2219 ;
  assign n2238 = n148 & ~n1109 ;
  assign n2237 = n137 & ~n1130 ;
  assign n2239 = n2238 ^ n2237 ;
  assign n2241 = n171 & ~n1196 ;
  assign n2240 = n160 & ~n1140 ;
  assign n2242 = n2241 ^ n2240 ;
  assign n2243 = ~n2239 & ~n2242 ;
  assign n2244 = n136 & ~n2243 ;
  assign n2230 = n148 & ~n1188 ;
  assign n2229 = n137 & ~n1205 ;
  assign n2231 = n2230 ^ n2229 ;
  assign n2233 = n171 & ~n1232 ;
  assign n2232 = n160 & ~n1213 ;
  assign n2234 = n2233 ^ n2232 ;
  assign n2235 = ~n2231 & ~n2234 ;
  assign n2236 = n185 & ~n2235 ;
  assign n2245 = n2244 ^ n2236 ;
  assign n2246 = ~n2228 & ~n2245 ;
  assign n2247 = x134 & n2246 ;
  assign n2284 = n2283 ^ n2247 ;
  assign n2297 = n185 & ~n369 ;
  assign n2296 = n136 & ~n458 ;
  assign n2298 = n2297 ^ n2296 ;
  assign n2300 = ~n228 & n279 ;
  assign n2299 = n254 & ~n502 ;
  assign n2301 = n2300 ^ n2299 ;
  assign n2302 = ~n2298 & ~n2301 ;
  assign n2303 = ~x134 & n2302 ;
  assign n2286 = n279 & ~n413 ;
  assign n2285 = ~n183 & n185 ;
  assign n2287 = n2286 ^ n2285 ;
  assign n2291 = n254 & n322 ;
  assign n2292 = n2291 ^ x133 ;
  assign n2288 = n136 & ~n275 ;
  assign n2289 = ~n253 & n2288 ;
  assign n2290 = n2289 ^ x132 ;
  assign n2293 = n2292 ^ n2290 ;
  assign n2294 = ~n2287 & ~n2293 ;
  assign n2295 = x134 & n2294 ;
  assign n2304 = n2303 ^ n2295 ;
  assign n2314 = n185 & ~n766 ;
  assign n2313 = n136 & ~n871 ;
  assign n2315 = n2314 ^ n2313 ;
  assign n2317 = n279 & ~n558 ;
  assign n2316 = n254 & ~n923 ;
  assign n2318 = n2317 ^ n2316 ;
  assign n2319 = ~n2315 & ~n2318 ;
  assign n2320 = ~x134 & n2319 ;
  assign n2306 = n254 & ~n610 ;
  assign n2305 = n279 & ~n818 ;
  assign n2307 = n2306 ^ n2305 ;
  assign n2309 = n136 & ~n711 ;
  assign n2308 = n185 & ~n663 ;
  assign n2310 = n2309 ^ n2308 ;
  assign n2311 = ~n2307 & ~n2310 ;
  assign n2312 = x134 & n2311 ;
  assign n2321 = n2320 ^ n2312 ;
  assign n2331 = n185 & ~n1037 ;
  assign n2330 = n136 & ~n1078 ;
  assign n2332 = n2331 ^ n2330 ;
  assign n2334 = n279 & ~n947 ;
  assign n2333 = n254 & ~n1098 ;
  assign n2335 = n2334 ^ n2333 ;
  assign n2336 = ~n2332 & ~n2335 ;
  assign n2337 = ~x134 & n2336 ;
  assign n2323 = n254 & ~n967 ;
  assign n2322 = n279 & ~n1057 ;
  assign n2324 = n2323 ^ n2322 ;
  assign n2326 = n136 & ~n1014 ;
  assign n2325 = n185 & ~n988 ;
  assign n2327 = n2326 ^ n2325 ;
  assign n2328 = ~n2324 & ~n2327 ;
  assign n2329 = x134 & n2328 ;
  assign n2338 = n2337 ^ n2329 ;
  assign n2348 = n136 & ~n1327 ;
  assign n2347 = n185 & ~n1291 ;
  assign n2349 = n2348 ^ n2347 ;
  assign n2351 = n254 & ~n1400 ;
  assign n2350 = n279 & ~n1252 ;
  assign n2352 = n2351 ^ n2350 ;
  assign n2353 = ~n2349 & ~n2352 ;
  assign n2354 = ~x134 & n2353 ;
  assign n2340 = n254 & ~n1179 ;
  assign n2339 = n279 & ~n1364 ;
  assign n2341 = n2340 ^ n2339 ;
  assign n2343 = n185 & ~n1216 ;
  assign n2342 = n136 & ~n1143 ;
  assign n2344 = n2343 ^ n2342 ;
  assign n2345 = ~n2341 & ~n2344 ;
  assign n2346 = x134 & n2345 ;
  assign n2355 = n2354 ^ n2346 ;
  assign n2367 = n185 & ~n1449 ;
  assign n2366 = n136 & ~n1466 ;
  assign n2368 = n2367 ^ n2366 ;
  assign n2370 = n279 & ~n1430 ;
  assign n2369 = n254 & ~n1474 ;
  assign n2371 = n2370 ^ n2369 ;
  assign n2372 = ~n2368 & ~n2371 ;
  assign n2373 = ~x134 & n2372 ;
  assign n2359 = n279 & n1457 ;
  assign n2356 = n136 & ~n1419 ;
  assign n2357 = ~n1416 & n2356 ;
  assign n2358 = n2357 ^ x132 ;
  assign n2360 = n2359 ^ n2358 ;
  assign n2362 = n185 & ~n1438 ;
  assign n2361 = n254 & ~n1412 ;
  assign n2363 = n2362 ^ n2361 ;
  assign n2364 = n2360 & ~n2363 ;
  assign n2365 = x134 & n2364 ;
  assign n2374 = n2373 ^ n2365 ;
  assign n2384 = n185 & ~n1522 ;
  assign n2383 = n136 & ~n1539 ;
  assign n2385 = n2384 ^ n2383 ;
  assign n2387 = n279 & ~n1503 ;
  assign n2386 = n254 & ~n1547 ;
  assign n2388 = n2387 ^ n2386 ;
  assign n2389 = ~n2385 & ~n2388 ;
  assign n2390 = ~x134 & n2389 ;
  assign n2376 = n279 & ~n1530 ;
  assign n2375 = n136 & ~n1494 ;
  assign n2377 = n2376 ^ n2375 ;
  assign n2379 = n185 & ~n1511 ;
  assign n2378 = n254 & ~n1486 ;
  assign n2380 = n2379 ^ n2378 ;
  assign n2381 = ~n2377 & ~n2380 ;
  assign n2382 = x134 & n2381 ;
  assign n2391 = n2390 ^ n2382 ;
  assign n2401 = n185 & ~n1595 ;
  assign n2400 = n136 & ~n1612 ;
  assign n2402 = n2401 ^ n2400 ;
  assign n2404 = n279 & ~n1576 ;
  assign n2403 = n254 & ~n1620 ;
  assign n2405 = n2404 ^ n2403 ;
  assign n2406 = ~n2402 & ~n2405 ;
  assign n2407 = ~x134 & n2406 ;
  assign n2393 = n279 & ~n1603 ;
  assign n2392 = n136 & ~n1567 ;
  assign n2394 = n2393 ^ n2392 ;
  assign n2396 = n185 & ~n1584 ;
  assign n2395 = n254 & ~n1559 ;
  assign n2397 = n2396 ^ n2395 ;
  assign n2398 = ~n2394 & ~n2397 ;
  assign n2399 = x134 & n2398 ;
  assign n2408 = n2407 ^ n2399 ;
  assign n2418 = n185 & ~n1668 ;
  assign n2417 = n279 & ~n1649 ;
  assign n2419 = n2418 ^ n2417 ;
  assign n2421 = n254 & ~n1693 ;
  assign n2420 = n136 & ~n1685 ;
  assign n2422 = n2421 ^ n2420 ;
  assign n2423 = ~n2419 & ~n2422 ;
  assign n2424 = ~x134 & n2423 ;
  assign n2410 = n136 & ~n1640 ;
  assign n2409 = n254 & ~n1632 ;
  assign n2411 = n2410 ^ n2409 ;
  assign n2413 = n185 & ~n1657 ;
  assign n2412 = n279 & ~n1676 ;
  assign n2414 = n2413 ^ n2412 ;
  assign n2415 = ~n2411 & ~n2414 ;
  assign n2416 = x134 & n2415 ;
  assign n2425 = n2424 ^ n2416 ;
  assign n2438 = n185 & ~n1742 ;
  assign n2437 = n279 & ~n1731 ;
  assign n2439 = n2438 ^ n2437 ;
  assign n2441 = n254 & ~n1767 ;
  assign n2440 = n136 & ~n1759 ;
  assign n2442 = n2441 ^ n2440 ;
  assign n2443 = ~n2439 & ~n2442 ;
  assign n2444 = ~x134 & n2443 ;
  assign n2427 = n136 & ~n1713 ;
  assign n2426 = n254 & ~n1705 ;
  assign n2428 = n2427 ^ n2426 ;
  assign n2432 = n279 & n1750 ;
  assign n2433 = n2432 ^ x133 ;
  assign n2429 = n185 & ~n1721 ;
  assign n2430 = ~n1718 & n2429 ;
  assign n2431 = n2430 ^ x132 ;
  assign n2434 = n2433 ^ n2431 ;
  assign n2435 = ~n2428 & n2434 ;
  assign n2436 = x134 & n2435 ;
  assign n2445 = n2444 ^ n2436 ;
  assign n2455 = n185 & ~n1815 ;
  assign n2454 = n279 & ~n1796 ;
  assign n2456 = n2455 ^ n2454 ;
  assign n2458 = n254 & ~n1840 ;
  assign n2457 = n136 & ~n1832 ;
  assign n2459 = n2458 ^ n2457 ;
  assign n2460 = ~n2456 & ~n2459 ;
  assign n2461 = ~x134 & n2460 ;
  assign n2447 = n136 & ~n1787 ;
  assign n2446 = n254 & ~n1779 ;
  assign n2448 = n2447 ^ n2446 ;
  assign n2450 = n185 & ~n1804 ;
  assign n2449 = n279 & ~n1823 ;
  assign n2451 = n2450 ^ n2449 ;
  assign n2452 = ~n2448 & ~n2451 ;
  assign n2453 = x134 & n2452 ;
  assign n2462 = n2461 ^ n2453 ;
  assign n2472 = n185 & ~n1888 ;
  assign n2471 = n136 & ~n1905 ;
  assign n2473 = n2472 ^ n2471 ;
  assign n2475 = n279 & ~n1869 ;
  assign n2474 = n254 & ~n1913 ;
  assign n2476 = n2475 ^ n2474 ;
  assign n2477 = ~n2473 & ~n2476 ;
  assign n2478 = ~x134 & n2477 ;
  assign n2464 = n136 & ~n1860 ;
  assign n2463 = n254 & ~n1852 ;
  assign n2465 = n2464 ^ n2463 ;
  assign n2467 = n185 & ~n1877 ;
  assign n2466 = n279 & ~n1896 ;
  assign n2468 = n2467 ^ n2466 ;
  assign n2469 = ~n2465 & ~n2468 ;
  assign n2470 = x134 & n2469 ;
  assign n2479 = n2478 ^ n2470 ;
  assign n2489 = n185 & ~n1961 ;
  assign n2488 = n136 & ~n1978 ;
  assign n2490 = n2489 ^ n2488 ;
  assign n2492 = n279 & ~n1942 ;
  assign n2491 = n254 & ~n1986 ;
  assign n2493 = n2492 ^ n2491 ;
  assign n2494 = ~n2490 & ~n2493 ;
  assign n2495 = ~x134 & n2494 ;
  assign n2481 = n136 & ~n1933 ;
  assign n2480 = n254 & ~n1925 ;
  assign n2482 = n2481 ^ n2480 ;
  assign n2484 = n185 & ~n1950 ;
  assign n2483 = n279 & ~n1969 ;
  assign n2485 = n2484 ^ n2483 ;
  assign n2486 = ~n2482 & ~n2485 ;
  assign n2487 = x134 & n2486 ;
  assign n2496 = n2495 ^ n2487 ;
  assign n2509 = n185 & ~n2035 ;
  assign n2508 = n136 & ~n2052 ;
  assign n2510 = n2509 ^ n2508 ;
  assign n2512 = n279 & ~n2024 ;
  assign n2511 = n254 & ~n2060 ;
  assign n2513 = n2512 ^ n2511 ;
  assign n2514 = ~n2510 & ~n2513 ;
  assign n2515 = ~x134 & n2514 ;
  assign n2498 = n136 & ~n2006 ;
  assign n2497 = n254 & ~n1998 ;
  assign n2499 = n2498 ^ n2497 ;
  assign n2503 = n279 & n2043 ;
  assign n2504 = n2503 ^ x133 ;
  assign n2500 = n185 & ~n2014 ;
  assign n2501 = ~n2011 & n2500 ;
  assign n2502 = n2501 ^ x132 ;
  assign n2505 = n2504 ^ n2502 ;
  assign n2506 = ~n2499 & n2505 ;
  assign n2507 = x134 & n2506 ;
  assign n2516 = n2515 ^ n2507 ;
  assign n2526 = n185 & ~n2108 ;
  assign n2525 = n136 & ~n2125 ;
  assign n2527 = n2526 ^ n2525 ;
  assign n2529 = n279 & ~n2089 ;
  assign n2528 = n254 & ~n2133 ;
  assign n2530 = n2529 ^ n2528 ;
  assign n2531 = ~n2527 & ~n2530 ;
  assign n2532 = ~x134 & n2531 ;
  assign n2518 = n136 & ~n2080 ;
  assign n2517 = n254 & ~n2072 ;
  assign n2519 = n2518 ^ n2517 ;
  assign n2521 = n185 & ~n2097 ;
  assign n2520 = n279 & ~n2116 ;
  assign n2522 = n2521 ^ n2520 ;
  assign n2523 = ~n2519 & ~n2522 ;
  assign n2524 = x134 & n2523 ;
  assign n2533 = n2532 ^ n2524 ;
  assign n2543 = n185 & ~n2181 ;
  assign n2542 = n136 & ~n2198 ;
  assign n2544 = n2543 ^ n2542 ;
  assign n2546 = n279 & ~n2162 ;
  assign n2545 = n254 & ~n2206 ;
  assign n2547 = n2546 ^ n2545 ;
  assign n2548 = ~n2544 & ~n2547 ;
  assign n2549 = ~x134 & n2548 ;
  assign n2535 = n136 & ~n2153 ;
  assign n2534 = n254 & ~n2145 ;
  assign n2536 = n2535 ^ n2534 ;
  assign n2538 = n185 & ~n2170 ;
  assign n2537 = n279 & ~n2189 ;
  assign n2539 = n2538 ^ n2537 ;
  assign n2540 = ~n2536 & ~n2539 ;
  assign n2541 = x134 & n2540 ;
  assign n2550 = n2549 ^ n2541 ;
  assign n2560 = n185 & ~n2254 ;
  assign n2559 = n136 & ~n2271 ;
  assign n2561 = n2560 ^ n2559 ;
  assign n2563 = n279 & ~n2235 ;
  assign n2562 = n254 & ~n2279 ;
  assign n2564 = n2563 ^ n2562 ;
  assign n2565 = ~n2561 & ~n2564 ;
  assign n2566 = ~x134 & n2565 ;
  assign n2552 = n136 & ~n2226 ;
  assign n2551 = n254 & ~n2218 ;
  assign n2553 = n2552 ^ n2551 ;
  assign n2555 = n185 & ~n2243 ;
  assign n2554 = n279 & ~n2262 ;
  assign n2556 = n2555 ^ n2554 ;
  assign n2557 = ~n2553 & ~n2556 ;
  assign n2558 = x134 & n2557 ;
  assign n2567 = n2566 ^ n2558 ;
  assign n2579 = n185 & ~n458 ;
  assign n2578 = n136 & ~n502 ;
  assign n2580 = n2579 ^ n2578 ;
  assign n2582 = ~n183 & n279 ;
  assign n2581 = ~n228 & n254 ;
  assign n2583 = n2582 ^ n2581 ;
  assign n2584 = ~n2580 & ~n2583 ;
  assign n2585 = ~x134 & n2584 ;
  assign n2569 = n254 & ~n413 ;
  assign n2568 = n279 & ~n369 ;
  assign n2570 = n2569 ^ n2568 ;
  assign n2572 = n185 & ~n275 ;
  assign n2573 = ~n253 & n2572 ;
  assign n2571 = n136 & n322 ;
  assign n2574 = n2573 ^ n2571 ;
  assign n2575 = n2574 ^ x133 ;
  assign n2576 = ~n2570 & ~n2575 ;
  assign n2577 = x134 & n2576 ;
  assign n2586 = n2585 ^ n2577 ;
  assign n2596 = n185 & ~n871 ;
  assign n2595 = n136 & ~n923 ;
  assign n2597 = n2596 ^ n2595 ;
  assign n2599 = n279 & ~n663 ;
  assign n2598 = n254 & ~n558 ;
  assign n2600 = n2599 ^ n2598 ;
  assign n2601 = ~n2597 & ~n2600 ;
  assign n2602 = ~x134 & n2601 ;
  assign n2588 = n136 & ~n610 ;
  assign n2587 = n254 & ~n818 ;
  assign n2589 = n2588 ^ n2587 ;
  assign n2591 = n185 & ~n711 ;
  assign n2590 = n279 & ~n766 ;
  assign n2592 = n2591 ^ n2590 ;
  assign n2593 = ~n2589 & ~n2592 ;
  assign n2594 = x134 & n2593 ;
  assign n2603 = n2602 ^ n2594 ;
  assign n2613 = n185 & ~n1078 ;
  assign n2612 = n136 & ~n1098 ;
  assign n2614 = n2613 ^ n2612 ;
  assign n2616 = n279 & ~n988 ;
  assign n2615 = n254 & ~n947 ;
  assign n2617 = n2616 ^ n2615 ;
  assign n2618 = ~n2614 & ~n2617 ;
  assign n2619 = ~x134 & n2618 ;
  assign n2605 = n136 & ~n967 ;
  assign n2604 = n254 & ~n1057 ;
  assign n2606 = n2605 ^ n2604 ;
  assign n2608 = n185 & ~n1014 ;
  assign n2607 = n279 & ~n1037 ;
  assign n2609 = n2608 ^ n2607 ;
  assign n2610 = ~n2606 & ~n2609 ;
  assign n2611 = x134 & n2610 ;
  assign n2620 = n2619 ^ n2611 ;
  assign n2630 = n185 & ~n1327 ;
  assign n2629 = n279 & ~n1216 ;
  assign n2631 = n2630 ^ n2629 ;
  assign n2633 = n136 & ~n1400 ;
  assign n2632 = n254 & ~n1252 ;
  assign n2634 = n2633 ^ n2632 ;
  assign n2635 = ~n2631 & ~n2634 ;
  assign n2636 = ~x134 & n2635 ;
  assign n2622 = n136 & ~n1179 ;
  assign n2621 = n279 & ~n1291 ;
  assign n2623 = n2622 ^ n2621 ;
  assign n2625 = n185 & ~n1143 ;
  assign n2624 = n254 & ~n1364 ;
  assign n2626 = n2625 ^ n2624 ;
  assign n2627 = ~n2623 & ~n2626 ;
  assign n2628 = x134 & n2627 ;
  assign n2637 = n2636 ^ n2628 ;
  assign n2649 = n185 & ~n1466 ;
  assign n2648 = n136 & ~n1474 ;
  assign n2650 = n2649 ^ n2648 ;
  assign n2652 = n279 & ~n1438 ;
  assign n2651 = n254 & ~n1430 ;
  assign n2653 = n2652 ^ n2651 ;
  assign n2654 = ~n2650 & ~n2653 ;
  assign n2655 = ~x134 & n2654 ;
  assign n2639 = n254 & ~n1457 ;
  assign n2638 = n279 & ~n1449 ;
  assign n2640 = n2639 ^ n2638 ;
  assign n2644 = n136 & n1412 ;
  assign n2641 = n185 & ~n1419 ;
  assign n2642 = ~n1416 & n2641 ;
  assign n2643 = n2642 ^ x133 ;
  assign n2645 = n2644 ^ n2643 ;
  assign n2646 = ~n2640 & ~n2645 ;
  assign n2647 = x134 & n2646 ;
  assign n2656 = n2655 ^ n2647 ;
  assign n2666 = n185 & ~n1539 ;
  assign n2665 = n136 & ~n1547 ;
  assign n2667 = n2666 ^ n2665 ;
  assign n2669 = n279 & ~n1511 ;
  assign n2668 = n254 & ~n1503 ;
  assign n2670 = n2669 ^ n2668 ;
  assign n2671 = ~n2667 & ~n2670 ;
  assign n2672 = ~x134 & n2671 ;
  assign n2658 = n254 & ~n1530 ;
  assign n2657 = n279 & ~n1522 ;
  assign n2659 = n2658 ^ n2657 ;
  assign n2661 = n136 & ~n1486 ;
  assign n2660 = n185 & ~n1494 ;
  assign n2662 = n2661 ^ n2660 ;
  assign n2663 = ~n2659 & ~n2662 ;
  assign n2664 = x134 & n2663 ;
  assign n2673 = n2672 ^ n2664 ;
  assign n2683 = n185 & ~n1612 ;
  assign n2682 = n136 & ~n1620 ;
  assign n2684 = n2683 ^ n2682 ;
  assign n2686 = n279 & ~n1584 ;
  assign n2685 = n254 & ~n1576 ;
  assign n2687 = n2686 ^ n2685 ;
  assign n2688 = ~n2684 & ~n2687 ;
  assign n2689 = ~x134 & n2688 ;
  assign n2675 = n254 & ~n1603 ;
  assign n2674 = n279 & ~n1595 ;
  assign n2676 = n2675 ^ n2674 ;
  assign n2678 = n136 & ~n1559 ;
  assign n2677 = n185 & ~n1567 ;
  assign n2679 = n2678 ^ n2677 ;
  assign n2680 = ~n2676 & ~n2679 ;
  assign n2681 = x134 & n2680 ;
  assign n2690 = n2689 ^ n2681 ;
  assign n2700 = n254 & ~n1649 ;
  assign n2699 = n279 & ~n1657 ;
  assign n2701 = n2700 ^ n2699 ;
  assign n2703 = n136 & ~n1693 ;
  assign n2702 = n185 & ~n1685 ;
  assign n2704 = n2703 ^ n2702 ;
  assign n2705 = ~n2701 & ~n2704 ;
  assign n2706 = ~x134 & n2705 ;
  assign n2692 = n185 & ~n1640 ;
  assign n2691 = n136 & ~n1632 ;
  assign n2693 = n2692 ^ n2691 ;
  assign n2695 = n279 & ~n1668 ;
  assign n2694 = n254 & ~n1676 ;
  assign n2696 = n2695 ^ n2694 ;
  assign n2697 = ~n2693 & ~n2696 ;
  assign n2698 = x134 & n2697 ;
  assign n2707 = n2706 ^ n2698 ;
  assign n2719 = n254 & n1731 ;
  assign n2716 = n279 & ~n1721 ;
  assign n2717 = ~n1718 & n2716 ;
  assign n2718 = n2717 ^ x133 ;
  assign n2720 = n2719 ^ n2718 ;
  assign n2722 = n136 & ~n1767 ;
  assign n2721 = n185 & ~n1759 ;
  assign n2723 = n2722 ^ n2721 ;
  assign n2724 = n2720 & ~n2723 ;
  assign n2725 = ~x134 & n2724 ;
  assign n2709 = n185 & ~n1713 ;
  assign n2708 = n136 & ~n1705 ;
  assign n2710 = n2709 ^ n2708 ;
  assign n2712 = n279 & ~n1742 ;
  assign n2711 = n254 & ~n1750 ;
  assign n2713 = n2712 ^ n2711 ;
  assign n2714 = ~n2710 & ~n2713 ;
  assign n2715 = x134 & n2714 ;
  assign n2726 = n2725 ^ n2715 ;
  assign n2736 = n254 & ~n1796 ;
  assign n2735 = n279 & ~n1804 ;
  assign n2737 = n2736 ^ n2735 ;
  assign n2739 = n136 & ~n1840 ;
  assign n2738 = n185 & ~n1832 ;
  assign n2740 = n2739 ^ n2738 ;
  assign n2741 = ~n2737 & ~n2740 ;
  assign n2742 = ~x134 & n2741 ;
  assign n2728 = n185 & ~n1787 ;
  assign n2727 = n136 & ~n1779 ;
  assign n2729 = n2728 ^ n2727 ;
  assign n2731 = n279 & ~n1815 ;
  assign n2730 = n254 & ~n1823 ;
  assign n2732 = n2731 ^ n2730 ;
  assign n2733 = ~n2729 & ~n2732 ;
  assign n2734 = x134 & n2733 ;
  assign n2743 = n2742 ^ n2734 ;
  assign n2753 = n185 & ~n1905 ;
  assign n2752 = n136 & ~n1913 ;
  assign n2754 = n2753 ^ n2752 ;
  assign n2756 = n279 & ~n1877 ;
  assign n2755 = n254 & ~n1869 ;
  assign n2757 = n2756 ^ n2755 ;
  assign n2758 = ~n2754 & ~n2757 ;
  assign n2759 = ~x134 & n2758 ;
  assign n2745 = n185 & ~n1860 ;
  assign n2744 = n136 & ~n1852 ;
  assign n2746 = n2745 ^ n2744 ;
  assign n2748 = n279 & ~n1888 ;
  assign n2747 = n254 & ~n1896 ;
  assign n2749 = n2748 ^ n2747 ;
  assign n2750 = ~n2746 & ~n2749 ;
  assign n2751 = x134 & n2750 ;
  assign n2760 = n2759 ^ n2751 ;
  assign n2770 = n185 & ~n1978 ;
  assign n2769 = n136 & ~n1986 ;
  assign n2771 = n2770 ^ n2769 ;
  assign n2773 = n279 & ~n1950 ;
  assign n2772 = n254 & ~n1942 ;
  assign n2774 = n2773 ^ n2772 ;
  assign n2775 = ~n2771 & ~n2774 ;
  assign n2776 = ~x134 & n2775 ;
  assign n2762 = n185 & ~n1933 ;
  assign n2761 = n136 & ~n1925 ;
  assign n2763 = n2762 ^ n2761 ;
  assign n2765 = n279 & ~n1961 ;
  assign n2764 = n254 & ~n1969 ;
  assign n2766 = n2765 ^ n2764 ;
  assign n2767 = ~n2763 & ~n2766 ;
  assign n2768 = x134 & n2767 ;
  assign n2777 = n2776 ^ n2768 ;
  assign n2787 = n185 & ~n2052 ;
  assign n2786 = n136 & ~n2060 ;
  assign n2788 = n2787 ^ n2786 ;
  assign n2792 = n254 & n2024 ;
  assign n2789 = n279 & ~n2014 ;
  assign n2790 = ~n2011 & n2789 ;
  assign n2791 = n2790 ^ x133 ;
  assign n2793 = n2792 ^ n2791 ;
  assign n2794 = ~n2788 & n2793 ;
  assign n2795 = ~x134 & n2794 ;
  assign n2779 = n185 & ~n2006 ;
  assign n2778 = n136 & ~n1998 ;
  assign n2780 = n2779 ^ n2778 ;
  assign n2782 = n279 & ~n2035 ;
  assign n2781 = n254 & ~n2043 ;
  assign n2783 = n2782 ^ n2781 ;
  assign n2784 = ~n2780 & ~n2783 ;
  assign n2785 = x134 & n2784 ;
  assign n2796 = n2795 ^ n2785 ;
  assign n2806 = n185 & ~n2125 ;
  assign n2805 = n136 & ~n2133 ;
  assign n2807 = n2806 ^ n2805 ;
  assign n2809 = n279 & ~n2097 ;
  assign n2808 = n254 & ~n2089 ;
  assign n2810 = n2809 ^ n2808 ;
  assign n2811 = ~n2807 & ~n2810 ;
  assign n2812 = ~x134 & n2811 ;
  assign n2798 = n185 & ~n2080 ;
  assign n2797 = n136 & ~n2072 ;
  assign n2799 = n2798 ^ n2797 ;
  assign n2801 = n279 & ~n2108 ;
  assign n2800 = n254 & ~n2116 ;
  assign n2802 = n2801 ^ n2800 ;
  assign n2803 = ~n2799 & ~n2802 ;
  assign n2804 = x134 & n2803 ;
  assign n2813 = n2812 ^ n2804 ;
  assign n2823 = n185 & ~n2198 ;
  assign n2822 = n136 & ~n2206 ;
  assign n2824 = n2823 ^ n2822 ;
  assign n2826 = n279 & ~n2170 ;
  assign n2825 = n254 & ~n2162 ;
  assign n2827 = n2826 ^ n2825 ;
  assign n2828 = ~n2824 & ~n2827 ;
  assign n2829 = ~x134 & n2828 ;
  assign n2815 = n185 & ~n2153 ;
  assign n2814 = n136 & ~n2145 ;
  assign n2816 = n2815 ^ n2814 ;
  assign n2818 = n279 & ~n2181 ;
  assign n2817 = n254 & ~n2189 ;
  assign n2819 = n2818 ^ n2817 ;
  assign n2820 = ~n2816 & ~n2819 ;
  assign n2821 = x134 & n2820 ;
  assign n2830 = n2829 ^ n2821 ;
  assign n2840 = n185 & ~n2271 ;
  assign n2839 = n136 & ~n2279 ;
  assign n2841 = n2840 ^ n2839 ;
  assign n2843 = n279 & ~n2243 ;
  assign n2842 = n254 & ~n2235 ;
  assign n2844 = n2843 ^ n2842 ;
  assign n2845 = ~n2841 & ~n2844 ;
  assign n2846 = ~x134 & n2845 ;
  assign n2832 = n185 & ~n2226 ;
  assign n2831 = n136 & ~n2218 ;
  assign n2833 = n2832 ^ n2831 ;
  assign n2835 = n279 & ~n2254 ;
  assign n2834 = n254 & ~n2262 ;
  assign n2836 = n2835 ^ n2834 ;
  assign n2837 = ~n2833 & ~n2836 ;
  assign n2838 = x134 & n2837 ;
  assign n2847 = n2846 ^ n2838 ;
  assign n2857 = n185 & ~n502 ;
  assign n2856 = n136 & ~n228 ;
  assign n2858 = n2857 ^ n2856 ;
  assign n2860 = ~n275 & n279 ;
  assign n2861 = ~n253 & n2860 ;
  assign n2859 = n183 & n254 ;
  assign n2862 = n2861 ^ n2859 ;
  assign n2863 = n2862 ^ x133 ;
  assign n2864 = ~n2858 & n2863 ;
  assign n2865 = ~x134 & n2864 ;
  assign n2849 = n136 & ~n413 ;
  assign n2848 = n254 & ~n369 ;
  assign n2850 = n2849 ^ n2848 ;
  assign n2852 = n185 & ~n322 ;
  assign n2851 = n279 & ~n458 ;
  assign n2853 = n2852 ^ n2851 ;
  assign n2854 = ~n2850 & ~n2853 ;
  assign n2855 = x134 & n2854 ;
  assign n2866 = n2865 ^ n2855 ;
  assign n2876 = n185 & ~n923 ;
  assign n2875 = n136 & ~n558 ;
  assign n2877 = n2876 ^ n2875 ;
  assign n2879 = n279 & ~n711 ;
  assign n2878 = n254 & ~n663 ;
  assign n2880 = n2879 ^ n2878 ;
  assign n2881 = ~n2877 & ~n2880 ;
  assign n2882 = ~x134 & n2881 ;
  assign n2868 = n185 & ~n610 ;
  assign n2867 = n136 & ~n818 ;
  assign n2869 = n2868 ^ n2867 ;
  assign n2871 = n279 & ~n871 ;
  assign n2870 = n254 & ~n766 ;
  assign n2872 = n2871 ^ n2870 ;
  assign n2873 = ~n2869 & ~n2872 ;
  assign n2874 = x134 & n2873 ;
  assign n2883 = n2882 ^ n2874 ;
  assign n2893 = n185 & ~n1098 ;
  assign n2892 = n136 & ~n947 ;
  assign n2894 = n2893 ^ n2892 ;
  assign n2896 = n279 & ~n1014 ;
  assign n2895 = n254 & ~n988 ;
  assign n2897 = n2896 ^ n2895 ;
  assign n2898 = ~n2894 & ~n2897 ;
  assign n2899 = ~x134 & n2898 ;
  assign n2885 = n185 & ~n967 ;
  assign n2884 = n136 & ~n1057 ;
  assign n2886 = n2885 ^ n2884 ;
  assign n2888 = n279 & ~n1078 ;
  assign n2887 = n254 & ~n1037 ;
  assign n2889 = n2888 ^ n2887 ;
  assign n2890 = ~n2886 & ~n2889 ;
  assign n2891 = x134 & n2890 ;
  assign n2900 = n2899 ^ n2891 ;
  assign n2910 = n279 & ~n1143 ;
  assign n2909 = n254 & ~n1216 ;
  assign n2911 = n2910 ^ n2909 ;
  assign n2913 = n185 & ~n1400 ;
  assign n2912 = n136 & ~n1252 ;
  assign n2914 = n2913 ^ n2912 ;
  assign n2915 = ~n2911 & ~n2914 ;
  assign n2916 = ~x134 & n2915 ;
  assign n2902 = n185 & ~n1179 ;
  assign n2901 = n279 & ~n1327 ;
  assign n2903 = n2902 ^ n2901 ;
  assign n2905 = n136 & ~n1364 ;
  assign n2904 = n254 & ~n1291 ;
  assign n2906 = n2905 ^ n2904 ;
  assign n2907 = ~n2903 & ~n2906 ;
  assign n2908 = x134 & n2907 ;
  assign n2917 = n2916 ^ n2908 ;
  assign n2929 = n185 & n1474 ;
  assign n2930 = n2929 ^ x133 ;
  assign n2926 = n279 & ~n1419 ;
  assign n2927 = ~n1416 & n2926 ;
  assign n2928 = n2927 ^ x132 ;
  assign n2931 = n2930 ^ n2928 ;
  assign n2933 = n254 & ~n1438 ;
  assign n2932 = n136 & ~n1430 ;
  assign n2934 = n2933 ^ n2932 ;
  assign n2935 = n2931 & ~n2934 ;
  assign n2936 = ~x134 & n2935 ;
  assign n2919 = n136 & ~n1457 ;
  assign n2918 = n254 & ~n1449 ;
  assign n2920 = n2919 ^ n2918 ;
  assign n2922 = n279 & ~n1466 ;
  assign n2921 = n185 & ~n1412 ;
  assign n2923 = n2922 ^ n2921 ;
  assign n2924 = ~n2920 & ~n2923 ;
  assign n2925 = x134 & n2924 ;
  assign n2937 = n2936 ^ n2925 ;
  assign n2947 = n279 & ~n1494 ;
  assign n2946 = n185 & ~n1547 ;
  assign n2948 = n2947 ^ n2946 ;
  assign n2950 = n254 & ~n1511 ;
  assign n2949 = n136 & ~n1503 ;
  assign n2951 = n2950 ^ n2949 ;
  assign n2952 = ~n2948 & ~n2951 ;
  assign n2953 = ~x134 & n2952 ;
  assign n2939 = n136 & ~n1530 ;
  assign n2938 = n254 & ~n1522 ;
  assign n2940 = n2939 ^ n2938 ;
  assign n2942 = n279 & ~n1539 ;
  assign n2941 = n185 & ~n1486 ;
  assign n2943 = n2942 ^ n2941 ;
  assign n2944 = ~n2940 & ~n2943 ;
  assign n2945 = x134 & n2944 ;
  assign n2954 = n2953 ^ n2945 ;
  assign n2964 = n279 & ~n1567 ;
  assign n2963 = n185 & ~n1620 ;
  assign n2965 = n2964 ^ n2963 ;
  assign n2967 = n254 & ~n1584 ;
  assign n2966 = n136 & ~n1576 ;
  assign n2968 = n2967 ^ n2966 ;
  assign n2969 = ~n2965 & ~n2968 ;
  assign n2970 = ~x134 & n2969 ;
  assign n2956 = n136 & ~n1603 ;
  assign n2955 = n254 & ~n1595 ;
  assign n2957 = n2956 ^ n2955 ;
  assign n2959 = n279 & ~n1612 ;
  assign n2958 = n185 & ~n1559 ;
  assign n2960 = n2959 ^ n2958 ;
  assign n2961 = ~n2957 & ~n2960 ;
  assign n2962 = x134 & n2961 ;
  assign n2971 = n2970 ^ n2962 ;
  assign n2981 = n279 & ~n1640 ;
  assign n2980 = n136 & ~n1649 ;
  assign n2982 = n2981 ^ n2980 ;
  assign n2984 = n185 & ~n1693 ;
  assign n2983 = n254 & ~n1657 ;
  assign n2985 = n2984 ^ n2983 ;
  assign n2986 = ~n2982 & ~n2985 ;
  assign n2987 = ~x134 & n2986 ;
  assign n2973 = n185 & ~n1632 ;
  assign n2972 = n136 & ~n1676 ;
  assign n2974 = n2973 ^ n2972 ;
  assign n2976 = n279 & ~n1685 ;
  assign n2975 = n254 & ~n1668 ;
  assign n2977 = n2976 ^ n2975 ;
  assign n2978 = ~n2974 & ~n2977 ;
  assign n2979 = x134 & n2978 ;
  assign n2988 = n2987 ^ n2979 ;
  assign n2998 = n279 & ~n1713 ;
  assign n2997 = n136 & ~n1731 ;
  assign n2999 = n2998 ^ n2997 ;
  assign n3001 = n254 & ~n1721 ;
  assign n3002 = ~n1718 & n3001 ;
  assign n3000 = n185 & n1767 ;
  assign n3003 = n3002 ^ n3000 ;
  assign n3004 = n3003 ^ x132 ;
  assign n3005 = ~n2999 & ~n3004 ;
  assign n3006 = ~x134 & n3005 ;
  assign n2990 = n185 & ~n1705 ;
  assign n2989 = n136 & ~n1750 ;
  assign n2991 = n2990 ^ n2989 ;
  assign n2993 = n279 & ~n1759 ;
  assign n2992 = n254 & ~n1742 ;
  assign n2994 = n2993 ^ n2992 ;
  assign n2995 = ~n2991 & ~n2994 ;
  assign n2996 = x134 & n2995 ;
  assign n3007 = n3006 ^ n2996 ;
  assign n3017 = n279 & ~n1787 ;
  assign n3016 = n136 & ~n1796 ;
  assign n3018 = n3017 ^ n3016 ;
  assign n3020 = n185 & ~n1840 ;
  assign n3019 = n254 & ~n1804 ;
  assign n3021 = n3020 ^ n3019 ;
  assign n3022 = ~n3018 & ~n3021 ;
  assign n3023 = ~x134 & n3022 ;
  assign n3009 = n185 & ~n1779 ;
  assign n3008 = n136 & ~n1823 ;
  assign n3010 = n3009 ^ n3008 ;
  assign n3012 = n279 & ~n1832 ;
  assign n3011 = n254 & ~n1815 ;
  assign n3013 = n3012 ^ n3011 ;
  assign n3014 = ~n3010 & ~n3013 ;
  assign n3015 = x134 & n3014 ;
  assign n3024 = n3023 ^ n3015 ;
  assign n3034 = n279 & ~n1860 ;
  assign n3033 = n185 & ~n1913 ;
  assign n3035 = n3034 ^ n3033 ;
  assign n3037 = n254 & ~n1877 ;
  assign n3036 = n136 & ~n1869 ;
  assign n3038 = n3037 ^ n3036 ;
  assign n3039 = ~n3035 & ~n3038 ;
  assign n3040 = ~x134 & n3039 ;
  assign n3026 = n185 & ~n1852 ;
  assign n3025 = n136 & ~n1896 ;
  assign n3027 = n3026 ^ n3025 ;
  assign n3029 = n279 & ~n1905 ;
  assign n3028 = n254 & ~n1888 ;
  assign n3030 = n3029 ^ n3028 ;
  assign n3031 = ~n3027 & ~n3030 ;
  assign n3032 = x134 & n3031 ;
  assign n3041 = n3040 ^ n3032 ;
  assign n3051 = n279 & ~n1933 ;
  assign n3050 = n185 & ~n1986 ;
  assign n3052 = n3051 ^ n3050 ;
  assign n3054 = n254 & ~n1950 ;
  assign n3053 = n136 & ~n1942 ;
  assign n3055 = n3054 ^ n3053 ;
  assign n3056 = ~n3052 & ~n3055 ;
  assign n3057 = ~x134 & n3056 ;
  assign n3043 = n185 & ~n1925 ;
  assign n3042 = n136 & ~n1969 ;
  assign n3044 = n3043 ^ n3042 ;
  assign n3046 = n279 & ~n1978 ;
  assign n3045 = n254 & ~n1961 ;
  assign n3047 = n3046 ^ n3045 ;
  assign n3048 = ~n3044 & ~n3047 ;
  assign n3049 = x134 & n3048 ;
  assign n3058 = n3057 ^ n3049 ;
  assign n3068 = n279 & ~n2006 ;
  assign n3067 = n185 & ~n2060 ;
  assign n3069 = n3068 ^ n3067 ;
  assign n3073 = n136 & n2024 ;
  assign n3074 = n3073 ^ x133 ;
  assign n3070 = n254 & ~n2014 ;
  assign n3071 = ~n2011 & n3070 ;
  assign n3072 = n3071 ^ x132 ;
  assign n3075 = n3074 ^ n3072 ;
  assign n3076 = ~n3069 & ~n3075 ;
  assign n3077 = ~x134 & n3076 ;
  assign n3060 = n185 & ~n1998 ;
  assign n3059 = n136 & ~n2043 ;
  assign n3061 = n3060 ^ n3059 ;
  assign n3063 = n279 & ~n2052 ;
  assign n3062 = n254 & ~n2035 ;
  assign n3064 = n3063 ^ n3062 ;
  assign n3065 = ~n3061 & ~n3064 ;
  assign n3066 = x134 & n3065 ;
  assign n3078 = n3077 ^ n3066 ;
  assign n3088 = n279 & ~n2080 ;
  assign n3087 = n185 & ~n2133 ;
  assign n3089 = n3088 ^ n3087 ;
  assign n3091 = n254 & ~n2097 ;
  assign n3090 = n136 & ~n2089 ;
  assign n3092 = n3091 ^ n3090 ;
  assign n3093 = ~n3089 & ~n3092 ;
  assign n3094 = ~x134 & n3093 ;
  assign n3080 = n185 & ~n2072 ;
  assign n3079 = n136 & ~n2116 ;
  assign n3081 = n3080 ^ n3079 ;
  assign n3083 = n279 & ~n2125 ;
  assign n3082 = n254 & ~n2108 ;
  assign n3084 = n3083 ^ n3082 ;
  assign n3085 = ~n3081 & ~n3084 ;
  assign n3086 = x134 & n3085 ;
  assign n3095 = n3094 ^ n3086 ;
  assign n3105 = n279 & ~n2153 ;
  assign n3104 = n185 & ~n2206 ;
  assign n3106 = n3105 ^ n3104 ;
  assign n3108 = n254 & ~n2170 ;
  assign n3107 = n136 & ~n2162 ;
  assign n3109 = n3108 ^ n3107 ;
  assign n3110 = ~n3106 & ~n3109 ;
  assign n3111 = ~x134 & n3110 ;
  assign n3097 = n185 & ~n2145 ;
  assign n3096 = n136 & ~n2189 ;
  assign n3098 = n3097 ^ n3096 ;
  assign n3100 = n279 & ~n2198 ;
  assign n3099 = n254 & ~n2181 ;
  assign n3101 = n3100 ^ n3099 ;
  assign n3102 = ~n3098 & ~n3101 ;
  assign n3103 = x134 & n3102 ;
  assign n3112 = n3111 ^ n3103 ;
  assign n3122 = n279 & ~n2226 ;
  assign n3121 = n185 & ~n2279 ;
  assign n3123 = n3122 ^ n3121 ;
  assign n3125 = n254 & ~n2243 ;
  assign n3124 = n136 & ~n2235 ;
  assign n3126 = n3125 ^ n3124 ;
  assign n3127 = ~n3123 & ~n3126 ;
  assign n3128 = ~x134 & n3127 ;
  assign n3114 = n185 & ~n2218 ;
  assign n3113 = n136 & ~n2262 ;
  assign n3115 = n3114 ^ n3113 ;
  assign n3117 = n279 & ~n2271 ;
  assign n3116 = n254 & ~n2254 ;
  assign n3118 = n3117 ^ n3116 ;
  assign n3119 = ~n3115 & ~n3118 ;
  assign n3120 = x134 & n3119 ;
  assign n3129 = n3128 ^ n3120 ;
  assign n3131 = ~x134 & n325 ;
  assign n3130 = x134 & n505 ;
  assign n3132 = n3131 ^ n3130 ;
  assign n3134 = ~x134 & n714 ;
  assign n3133 = x134 & n926 ;
  assign n3135 = n3134 ^ n3133 ;
  assign n3137 = ~x134 & n1017 ;
  assign n3136 = x134 & n1101 ;
  assign n3138 = n3137 ^ n3136 ;
  assign n3140 = ~x134 & n1255 ;
  assign n3139 = x134 & n1403 ;
  assign n3141 = n3140 ^ n3139 ;
  assign n3143 = ~x134 & n1441 ;
  assign n3142 = x134 & n1477 ;
  assign n3144 = n3143 ^ n3142 ;
  assign n3146 = ~x134 & n1514 ;
  assign n3145 = x134 & n1550 ;
  assign n3147 = n3146 ^ n3145 ;
  assign n3149 = ~x134 & n1587 ;
  assign n3148 = x134 & n1623 ;
  assign n3150 = n3149 ^ n3148 ;
  assign n3152 = ~x134 & n1660 ;
  assign n3151 = x134 & n1696 ;
  assign n3153 = n3152 ^ n3151 ;
  assign n3155 = ~x134 & n1734 ;
  assign n3154 = x134 & n1770 ;
  assign n3156 = n3155 ^ n3154 ;
  assign n3158 = ~x134 & n1807 ;
  assign n3157 = x134 & n1843 ;
  assign n3159 = n3158 ^ n3157 ;
  assign n3161 = ~x134 & n1880 ;
  assign n3160 = x134 & n1916 ;
  assign n3162 = n3161 ^ n3160 ;
  assign n3164 = ~x134 & n1953 ;
  assign n3163 = x134 & n1989 ;
  assign n3165 = n3164 ^ n3163 ;
  assign n3167 = ~x134 & n2027 ;
  assign n3166 = x134 & n2063 ;
  assign n3168 = n3167 ^ n3166 ;
  assign n3170 = ~x134 & n2100 ;
  assign n3169 = x134 & n2136 ;
  assign n3171 = n3170 ^ n3169 ;
  assign n3173 = ~x134 & n2173 ;
  assign n3172 = x134 & n2209 ;
  assign n3174 = n3173 ^ n3172 ;
  assign n3176 = ~x134 & n2246 ;
  assign n3175 = x134 & n2282 ;
  assign n3177 = n3176 ^ n3175 ;
  assign n3179 = ~x134 & n2294 ;
  assign n3178 = x134 & n2302 ;
  assign n3180 = n3179 ^ n3178 ;
  assign n3182 = ~x134 & n2311 ;
  assign n3181 = x134 & n2319 ;
  assign n3183 = n3182 ^ n3181 ;
  assign n3185 = ~x134 & n2328 ;
  assign n3184 = x134 & n2336 ;
  assign n3186 = n3185 ^ n3184 ;
  assign n3188 = ~x134 & n2345 ;
  assign n3187 = x134 & n2353 ;
  assign n3189 = n3188 ^ n3187 ;
  assign n3191 = ~x134 & n2364 ;
  assign n3190 = x134 & n2372 ;
  assign n3192 = n3191 ^ n3190 ;
  assign n3194 = ~x134 & n2381 ;
  assign n3193 = x134 & n2389 ;
  assign n3195 = n3194 ^ n3193 ;
  assign n3197 = ~x134 & n2398 ;
  assign n3196 = x134 & n2406 ;
  assign n3198 = n3197 ^ n3196 ;
  assign n3200 = ~x134 & n2415 ;
  assign n3199 = x134 & n2423 ;
  assign n3201 = n3200 ^ n3199 ;
  assign n3203 = ~x134 & n2435 ;
  assign n3202 = x134 & n2443 ;
  assign n3204 = n3203 ^ n3202 ;
  assign n3206 = ~x134 & n2452 ;
  assign n3205 = x134 & n2460 ;
  assign n3207 = n3206 ^ n3205 ;
  assign n3209 = ~x134 & n2469 ;
  assign n3208 = x134 & n2477 ;
  assign n3210 = n3209 ^ n3208 ;
  assign n3212 = ~x134 & n2486 ;
  assign n3211 = x134 & n2494 ;
  assign n3213 = n3212 ^ n3211 ;
  assign n3215 = ~x134 & n2506 ;
  assign n3214 = x134 & n2514 ;
  assign n3216 = n3215 ^ n3214 ;
  assign n3218 = ~x134 & n2523 ;
  assign n3217 = x134 & n2531 ;
  assign n3219 = n3218 ^ n3217 ;
  assign n3221 = ~x134 & n2540 ;
  assign n3220 = x134 & n2548 ;
  assign n3222 = n3221 ^ n3220 ;
  assign n3224 = ~x134 & n2557 ;
  assign n3223 = x134 & n2565 ;
  assign n3225 = n3224 ^ n3223 ;
  assign n3227 = ~x134 & n2576 ;
  assign n3226 = x134 & n2584 ;
  assign n3228 = n3227 ^ n3226 ;
  assign n3230 = ~x134 & n2593 ;
  assign n3229 = x134 & n2601 ;
  assign n3231 = n3230 ^ n3229 ;
  assign n3233 = ~x134 & n2610 ;
  assign n3232 = x134 & n2618 ;
  assign n3234 = n3233 ^ n3232 ;
  assign n3236 = ~x134 & n2627 ;
  assign n3235 = x134 & n2635 ;
  assign n3237 = n3236 ^ n3235 ;
  assign n3239 = ~x134 & n2646 ;
  assign n3238 = x134 & n2654 ;
  assign n3240 = n3239 ^ n3238 ;
  assign n3242 = ~x134 & n2663 ;
  assign n3241 = x134 & n2671 ;
  assign n3243 = n3242 ^ n3241 ;
  assign n3245 = ~x134 & n2680 ;
  assign n3244 = x134 & n2688 ;
  assign n3246 = n3245 ^ n3244 ;
  assign n3248 = ~x134 & n2697 ;
  assign n3247 = x134 & n2705 ;
  assign n3249 = n3248 ^ n3247 ;
  assign n3251 = ~x134 & n2714 ;
  assign n3250 = x134 & n2724 ;
  assign n3252 = n3251 ^ n3250 ;
  assign n3254 = ~x134 & n2733 ;
  assign n3253 = x134 & n2741 ;
  assign n3255 = n3254 ^ n3253 ;
  assign n3257 = ~x134 & n2750 ;
  assign n3256 = x134 & n2758 ;
  assign n3258 = n3257 ^ n3256 ;
  assign n3260 = ~x134 & n2767 ;
  assign n3259 = x134 & n2775 ;
  assign n3261 = n3260 ^ n3259 ;
  assign n3263 = ~x134 & n2784 ;
  assign n3262 = x134 & n2794 ;
  assign n3264 = n3263 ^ n3262 ;
  assign n3266 = ~x134 & n2803 ;
  assign n3265 = x134 & n2811 ;
  assign n3267 = n3266 ^ n3265 ;
  assign n3269 = ~x134 & n2820 ;
  assign n3268 = x134 & n2828 ;
  assign n3270 = n3269 ^ n3268 ;
  assign n3272 = ~x134 & n2837 ;
  assign n3271 = x134 & n2845 ;
  assign n3273 = n3272 ^ n3271 ;
  assign n3275 = ~x134 & n2854 ;
  assign n3274 = x134 & n2864 ;
  assign n3276 = n3275 ^ n3274 ;
  assign n3278 = ~x134 & n2873 ;
  assign n3277 = x134 & n2881 ;
  assign n3279 = n3278 ^ n3277 ;
  assign n3281 = ~x134 & n2890 ;
  assign n3280 = x134 & n2898 ;
  assign n3282 = n3281 ^ n3280 ;
  assign n3284 = ~x134 & n2907 ;
  assign n3283 = x134 & n2915 ;
  assign n3285 = n3284 ^ n3283 ;
  assign n3287 = ~x134 & n2924 ;
  assign n3286 = x134 & n2935 ;
  assign n3288 = n3287 ^ n3286 ;
  assign n3290 = ~x134 & n2944 ;
  assign n3289 = x134 & n2952 ;
  assign n3291 = n3290 ^ n3289 ;
  assign n3293 = ~x134 & n2961 ;
  assign n3292 = x134 & n2969 ;
  assign n3294 = n3293 ^ n3292 ;
  assign n3296 = ~x134 & n2978 ;
  assign n3295 = x134 & n2986 ;
  assign n3297 = n3296 ^ n3295 ;
  assign n3299 = ~x134 & n2995 ;
  assign n3298 = x134 & n3005 ;
  assign n3300 = n3299 ^ n3298 ;
  assign n3302 = ~x134 & n3014 ;
  assign n3301 = x134 & n3022 ;
  assign n3303 = n3302 ^ n3301 ;
  assign n3305 = ~x134 & n3031 ;
  assign n3304 = x134 & n3039 ;
  assign n3306 = n3305 ^ n3304 ;
  assign n3308 = ~x134 & n3048 ;
  assign n3307 = x134 & n3056 ;
  assign n3309 = n3308 ^ n3307 ;
  assign n3311 = ~x134 & n3065 ;
  assign n3310 = x134 & n3076 ;
  assign n3312 = n3311 ^ n3310 ;
  assign n3314 = ~x134 & n3085 ;
  assign n3313 = x134 & n3093 ;
  assign n3315 = n3314 ^ n3313 ;
  assign n3317 = ~x134 & n3102 ;
  assign n3316 = x134 & n3110 ;
  assign n3318 = n3317 ^ n3316 ;
  assign n3320 = ~x134 & n3119 ;
  assign n3319 = x134 & n3127 ;
  assign n3321 = n3320 ^ n3319 ;
  assign y0 = ~n507 ;
  assign y1 = ~n928 ;
  assign y2 = ~n1103 ;
  assign y3 = ~n1405 ;
  assign y4 = ~n1479 ;
  assign y5 = ~n1552 ;
  assign y6 = ~n1625 ;
  assign y7 = ~n1698 ;
  assign y8 = ~n1772 ;
  assign y9 = ~n1845 ;
  assign y10 = ~n1918 ;
  assign y11 = ~n1991 ;
  assign y12 = ~n2065 ;
  assign y13 = ~n2138 ;
  assign y14 = ~n2211 ;
  assign y15 = ~n2284 ;
  assign y16 = ~n2304 ;
  assign y17 = ~n2321 ;
  assign y18 = ~n2338 ;
  assign y19 = ~n2355 ;
  assign y20 = ~n2374 ;
  assign y21 = ~n2391 ;
  assign y22 = ~n2408 ;
  assign y23 = ~n2425 ;
  assign y24 = ~n2445 ;
  assign y25 = ~n2462 ;
  assign y26 = ~n2479 ;
  assign y27 = ~n2496 ;
  assign y28 = ~n2516 ;
  assign y29 = ~n2533 ;
  assign y30 = ~n2550 ;
  assign y31 = ~n2567 ;
  assign y32 = ~n2586 ;
  assign y33 = ~n2603 ;
  assign y34 = ~n2620 ;
  assign y35 = ~n2637 ;
  assign y36 = ~n2656 ;
  assign y37 = ~n2673 ;
  assign y38 = ~n2690 ;
  assign y39 = ~n2707 ;
  assign y40 = ~n2726 ;
  assign y41 = ~n2743 ;
  assign y42 = ~n2760 ;
  assign y43 = ~n2777 ;
  assign y44 = ~n2796 ;
  assign y45 = ~n2813 ;
  assign y46 = ~n2830 ;
  assign y47 = ~n2847 ;
  assign y48 = ~n2866 ;
  assign y49 = ~n2883 ;
  assign y50 = ~n2900 ;
  assign y51 = ~n2917 ;
  assign y52 = ~n2937 ;
  assign y53 = ~n2954 ;
  assign y54 = ~n2971 ;
  assign y55 = ~n2988 ;
  assign y56 = ~n3007 ;
  assign y57 = ~n3024 ;
  assign y58 = ~n3041 ;
  assign y59 = ~n3058 ;
  assign y60 = ~n3078 ;
  assign y61 = ~n3095 ;
  assign y62 = ~n3112 ;
  assign y63 = ~n3129 ;
  assign y64 = ~n3132 ;
  assign y65 = ~n3135 ;
  assign y66 = ~n3138 ;
  assign y67 = ~n3141 ;
  assign y68 = ~n3144 ;
  assign y69 = ~n3147 ;
  assign y70 = ~n3150 ;
  assign y71 = ~n3153 ;
  assign y72 = ~n3156 ;
  assign y73 = ~n3159 ;
  assign y74 = ~n3162 ;
  assign y75 = ~n3165 ;
  assign y76 = ~n3168 ;
  assign y77 = ~n3171 ;
  assign y78 = ~n3174 ;
  assign y79 = ~n3177 ;
  assign y80 = ~n3180 ;
  assign y81 = ~n3183 ;
  assign y82 = ~n3186 ;
  assign y83 = ~n3189 ;
  assign y84 = ~n3192 ;
  assign y85 = ~n3195 ;
  assign y86 = ~n3198 ;
  assign y87 = ~n3201 ;
  assign y88 = ~n3204 ;
  assign y89 = ~n3207 ;
  assign y90 = ~n3210 ;
  assign y91 = ~n3213 ;
  assign y92 = ~n3216 ;
  assign y93 = ~n3219 ;
  assign y94 = ~n3222 ;
  assign y95 = ~n3225 ;
  assign y96 = ~n3228 ;
  assign y97 = ~n3231 ;
  assign y98 = ~n3234 ;
  assign y99 = ~n3237 ;
  assign y100 = ~n3240 ;
  assign y101 = ~n3243 ;
  assign y102 = ~n3246 ;
  assign y103 = ~n3249 ;
  assign y104 = ~n3252 ;
  assign y105 = ~n3255 ;
  assign y106 = ~n3258 ;
  assign y107 = ~n3261 ;
  assign y108 = ~n3264 ;
  assign y109 = ~n3267 ;
  assign y110 = ~n3270 ;
  assign y111 = ~n3273 ;
  assign y112 = ~n3276 ;
  assign y113 = ~n3279 ;
  assign y114 = ~n3282 ;
  assign y115 = ~n3285 ;
  assign y116 = ~n3288 ;
  assign y117 = ~n3291 ;
  assign y118 = ~n3294 ;
  assign y119 = ~n3297 ;
  assign y120 = ~n3300 ;
  assign y121 = ~n3303 ;
  assign y122 = ~n3306 ;
  assign y123 = ~n3309 ;
  assign y124 = ~n3312 ;
  assign y125 = ~n3315 ;
  assign y126 = ~n3318 ;
  assign y127 = ~n3321 ;
endmodule
