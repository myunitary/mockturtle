module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 ;
  assign n9 = x4 & x5 ;
  assign n10 = n9 ^ x4 ;
  assign n11 = n10 ^ x5 ;
  assign n12 = x6 & x7 ;
  assign n13 = n12 ^ x7 ;
  assign n14 = ~n11 & n13 ;
  assign n15 = x0 & x2 ;
  assign n16 = n15 ^ x0 ;
  assign n17 = n16 ^ x2 ;
  assign n18 = x1 & x3 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = ~n17 & ~n20 ;
  assign n22 = n14 & n21 ;
  assign n23 = n16 & ~n20 ;
  assign n24 = n14 & n23 ;
  assign n25 = ~n17 & n19 ;
  assign n26 = n14 & n25 ;
  assign n27 = n16 & n19 ;
  assign n28 = n14 & n27 ;
  assign n29 = n15 ^ x2 ;
  assign n30 = ~n20 & n29 ;
  assign n31 = n14 & n30 ;
  assign n32 = n15 & ~n20 ;
  assign n33 = n14 & n32 ;
  assign n34 = n19 & n29 ;
  assign n35 = n14 & n34 ;
  assign n36 = n15 & n19 ;
  assign n37 = n14 & n36 ;
  assign n38 = n18 ^ x3 ;
  assign n39 = ~n17 & n38 ;
  assign n40 = n14 & n39 ;
  assign n41 = n16 & n38 ;
  assign n42 = n14 & n41 ;
  assign n43 = ~n17 & n18 ;
  assign n44 = n14 & n43 ;
  assign n45 = n16 & n18 ;
  assign n46 = n14 & n45 ;
  assign n47 = n29 & n38 ;
  assign n48 = n14 & n47 ;
  assign n49 = n15 & n38 ;
  assign n50 = n14 & n49 ;
  assign n51 = n18 & n29 ;
  assign n52 = n14 & n51 ;
  assign n53 = n15 & n18 ;
  assign n54 = n14 & n53 ;
  assign n55 = n10 & n13 ;
  assign n56 = n21 & n55 ;
  assign n57 = n23 & n55 ;
  assign n58 = n25 & n55 ;
  assign n59 = n27 & n55 ;
  assign n60 = n30 & n55 ;
  assign n61 = n32 & n55 ;
  assign n62 = n34 & n55 ;
  assign n63 = n36 & n55 ;
  assign n64 = n39 & n55 ;
  assign n65 = n41 & n55 ;
  assign n66 = n43 & n55 ;
  assign n67 = n45 & n55 ;
  assign n68 = n47 & n55 ;
  assign n69 = n49 & n55 ;
  assign n70 = n51 & n55 ;
  assign n71 = n53 & n55 ;
  assign n72 = n9 ^ x5 ;
  assign n73 = n13 & n72 ;
  assign n74 = n21 & n73 ;
  assign n75 = n23 & n73 ;
  assign n76 = n25 & n73 ;
  assign n77 = n27 & n73 ;
  assign n78 = n30 & n73 ;
  assign n79 = n32 & n73 ;
  assign n80 = n34 & n73 ;
  assign n81 = n36 & n73 ;
  assign n82 = n39 & n73 ;
  assign n83 = n41 & n73 ;
  assign n84 = n43 & n73 ;
  assign n85 = n45 & n73 ;
  assign n86 = n47 & n73 ;
  assign n87 = n49 & n73 ;
  assign n88 = n51 & n73 ;
  assign n89 = n53 & n73 ;
  assign n90 = n9 & n13 ;
  assign n91 = n21 & n90 ;
  assign n92 = n23 & n90 ;
  assign n93 = n25 & n90 ;
  assign n94 = n27 & n90 ;
  assign n95 = n30 & n90 ;
  assign n96 = n32 & n90 ;
  assign n97 = n34 & n90 ;
  assign n98 = n36 & n90 ;
  assign n99 = n39 & n90 ;
  assign n100 = n41 & n90 ;
  assign n101 = n43 & n90 ;
  assign n102 = n45 & n90 ;
  assign n103 = n47 & n90 ;
  assign n104 = n49 & n90 ;
  assign n105 = n51 & n90 ;
  assign n106 = n53 & n90 ;
  assign n107 = ~n11 & n12 ;
  assign n108 = n21 & n107 ;
  assign n109 = n23 & n107 ;
  assign n110 = n25 & n107 ;
  assign n111 = n27 & n107 ;
  assign n112 = n30 & n107 ;
  assign n113 = n32 & n107 ;
  assign n114 = n34 & n107 ;
  assign n115 = n36 & n107 ;
  assign n116 = n39 & n107 ;
  assign n117 = n41 & n107 ;
  assign n118 = n43 & n107 ;
  assign n119 = n45 & n107 ;
  assign n120 = n47 & n107 ;
  assign n121 = n49 & n107 ;
  assign n122 = n51 & n107 ;
  assign n123 = n53 & n107 ;
  assign n124 = n10 & n12 ;
  assign n125 = n21 & n124 ;
  assign n126 = n23 & n124 ;
  assign n127 = n25 & n124 ;
  assign n128 = n27 & n124 ;
  assign n129 = n30 & n124 ;
  assign n130 = n32 & n124 ;
  assign n131 = n34 & n124 ;
  assign n132 = n36 & n124 ;
  assign n133 = n39 & n124 ;
  assign n134 = n41 & n124 ;
  assign n135 = n43 & n124 ;
  assign n136 = n45 & n124 ;
  assign n137 = n47 & n124 ;
  assign n138 = n49 & n124 ;
  assign n139 = n51 & n124 ;
  assign n140 = n53 & n124 ;
  assign n141 = n12 & n72 ;
  assign n142 = n21 & n141 ;
  assign n143 = n23 & n141 ;
  assign n144 = n25 & n141 ;
  assign n145 = n27 & n141 ;
  assign n146 = n30 & n141 ;
  assign n147 = n32 & n141 ;
  assign n148 = n34 & n141 ;
  assign n149 = n36 & n141 ;
  assign n150 = n39 & n141 ;
  assign n151 = n41 & n141 ;
  assign n152 = n43 & n141 ;
  assign n153 = n45 & n141 ;
  assign n154 = n47 & n141 ;
  assign n155 = n49 & n141 ;
  assign n156 = n51 & n141 ;
  assign n157 = n53 & n141 ;
  assign n158 = n9 & n12 ;
  assign n159 = n21 & n158 ;
  assign n160 = n23 & n158 ;
  assign n161 = n25 & n158 ;
  assign n162 = n27 & n158 ;
  assign n163 = n30 & n158 ;
  assign n164 = n32 & n158 ;
  assign n165 = n34 & n158 ;
  assign n166 = n36 & n158 ;
  assign n167 = n39 & n158 ;
  assign n168 = n41 & n158 ;
  assign n169 = n43 & n158 ;
  assign n170 = n45 & n158 ;
  assign n171 = n47 & n158 ;
  assign n172 = n49 & n158 ;
  assign n173 = n51 & n158 ;
  assign n174 = n53 & n158 ;
  assign n175 = n12 ^ x6 ;
  assign n176 = n175 ^ x7 ;
  assign n177 = ~n11 & ~n176 ;
  assign n178 = n21 & n177 ;
  assign n179 = n23 & n177 ;
  assign n180 = n25 & n177 ;
  assign n181 = n27 & n177 ;
  assign n182 = n30 & n177 ;
  assign n183 = n32 & n177 ;
  assign n184 = n34 & n177 ;
  assign n185 = n36 & n177 ;
  assign n186 = n39 & n177 ;
  assign n187 = n41 & n177 ;
  assign n188 = n43 & n177 ;
  assign n189 = n45 & n177 ;
  assign n190 = n47 & n177 ;
  assign n191 = n49 & n177 ;
  assign n192 = n51 & n177 ;
  assign n193 = n53 & n177 ;
  assign n194 = n10 & ~n176 ;
  assign n195 = n21 & n194 ;
  assign n196 = n23 & n194 ;
  assign n197 = n25 & n194 ;
  assign n198 = n27 & n194 ;
  assign n199 = n30 & n194 ;
  assign n200 = n32 & n194 ;
  assign n201 = n34 & n194 ;
  assign n202 = n36 & n194 ;
  assign n203 = n39 & n194 ;
  assign n204 = n41 & n194 ;
  assign n205 = n43 & n194 ;
  assign n206 = n45 & n194 ;
  assign n207 = n47 & n194 ;
  assign n208 = n49 & n194 ;
  assign n209 = n51 & n194 ;
  assign n210 = n53 & n194 ;
  assign n211 = n72 & ~n176 ;
  assign n212 = n21 & n211 ;
  assign n213 = n23 & n211 ;
  assign n214 = n25 & n211 ;
  assign n215 = n27 & n211 ;
  assign n216 = n30 & n211 ;
  assign n217 = n32 & n211 ;
  assign n218 = n34 & n211 ;
  assign n219 = n36 & n211 ;
  assign n220 = n39 & n211 ;
  assign n221 = n41 & n211 ;
  assign n222 = n43 & n211 ;
  assign n223 = n45 & n211 ;
  assign n224 = n47 & n211 ;
  assign n225 = n49 & n211 ;
  assign n226 = n51 & n211 ;
  assign n227 = n53 & n211 ;
  assign n228 = n9 & ~n176 ;
  assign n229 = n21 & n228 ;
  assign n230 = n23 & n228 ;
  assign n231 = n25 & n228 ;
  assign n232 = n27 & n228 ;
  assign n233 = n30 & n228 ;
  assign n234 = n32 & n228 ;
  assign n235 = n34 & n228 ;
  assign n236 = n36 & n228 ;
  assign n237 = n39 & n228 ;
  assign n238 = n41 & n228 ;
  assign n239 = n43 & n228 ;
  assign n240 = n45 & n228 ;
  assign n241 = n47 & n228 ;
  assign n242 = n49 & n228 ;
  assign n243 = n51 & n228 ;
  assign n244 = n53 & n228 ;
  assign n245 = ~n11 & n175 ;
  assign n246 = n21 & n245 ;
  assign n247 = n23 & n245 ;
  assign n248 = n25 & n245 ;
  assign n249 = n27 & n245 ;
  assign n250 = n30 & n245 ;
  assign n251 = n32 & n245 ;
  assign n252 = n34 & n245 ;
  assign n253 = n36 & n245 ;
  assign n254 = n39 & n245 ;
  assign n255 = n41 & n245 ;
  assign n256 = n43 & n245 ;
  assign n257 = n45 & n245 ;
  assign n258 = n47 & n245 ;
  assign n259 = n49 & n245 ;
  assign n260 = n51 & n245 ;
  assign n261 = n53 & n245 ;
  assign n262 = n10 & n175 ;
  assign n263 = n21 & n262 ;
  assign n264 = n23 & n262 ;
  assign n265 = n25 & n262 ;
  assign n266 = n27 & n262 ;
  assign n267 = n30 & n262 ;
  assign n268 = n32 & n262 ;
  assign n269 = n34 & n262 ;
  assign n270 = n36 & n262 ;
  assign n271 = n39 & n262 ;
  assign n272 = n41 & n262 ;
  assign n273 = n43 & n262 ;
  assign n274 = n45 & n262 ;
  assign n275 = n47 & n262 ;
  assign n276 = n49 & n262 ;
  assign n277 = n51 & n262 ;
  assign n278 = n53 & n262 ;
  assign n279 = n72 & n175 ;
  assign n280 = n21 & n279 ;
  assign n281 = n23 & n279 ;
  assign n282 = n25 & n279 ;
  assign n283 = n27 & n279 ;
  assign n284 = n30 & n279 ;
  assign n285 = n32 & n279 ;
  assign n286 = n34 & n279 ;
  assign n287 = n36 & n279 ;
  assign n288 = n39 & n279 ;
  assign n289 = n41 & n279 ;
  assign n290 = n43 & n279 ;
  assign n291 = n45 & n279 ;
  assign n292 = n47 & n279 ;
  assign n293 = n49 & n279 ;
  assign n294 = n51 & n279 ;
  assign n295 = n53 & n279 ;
  assign n296 = n9 & n175 ;
  assign n297 = n21 & n296 ;
  assign n298 = n23 & n296 ;
  assign n299 = n25 & n296 ;
  assign n300 = n27 & n296 ;
  assign n301 = n30 & n296 ;
  assign n302 = n32 & n296 ;
  assign n303 = n34 & n296 ;
  assign n304 = n36 & n296 ;
  assign n305 = n39 & n296 ;
  assign n306 = n41 & n296 ;
  assign n307 = n43 & n296 ;
  assign n308 = n45 & n296 ;
  assign n309 = n47 & n296 ;
  assign n310 = n49 & n296 ;
  assign n311 = n51 & n296 ;
  assign n312 = n53 & n296 ;
  assign y0 = n22 ;
  assign y1 = n24 ;
  assign y2 = n26 ;
  assign y3 = n28 ;
  assign y4 = n31 ;
  assign y5 = n33 ;
  assign y6 = n35 ;
  assign y7 = n37 ;
  assign y8 = n40 ;
  assign y9 = n42 ;
  assign y10 = n44 ;
  assign y11 = n46 ;
  assign y12 = n48 ;
  assign y13 = n50 ;
  assign y14 = n52 ;
  assign y15 = n54 ;
  assign y16 = n56 ;
  assign y17 = n57 ;
  assign y18 = n58 ;
  assign y19 = n59 ;
  assign y20 = n60 ;
  assign y21 = n61 ;
  assign y22 = n62 ;
  assign y23 = n63 ;
  assign y24 = n64 ;
  assign y25 = n65 ;
  assign y26 = n66 ;
  assign y27 = n67 ;
  assign y28 = n68 ;
  assign y29 = n69 ;
  assign y30 = n70 ;
  assign y31 = n71 ;
  assign y32 = n74 ;
  assign y33 = n75 ;
  assign y34 = n76 ;
  assign y35 = n77 ;
  assign y36 = n78 ;
  assign y37 = n79 ;
  assign y38 = n80 ;
  assign y39 = n81 ;
  assign y40 = n82 ;
  assign y41 = n83 ;
  assign y42 = n84 ;
  assign y43 = n85 ;
  assign y44 = n86 ;
  assign y45 = n87 ;
  assign y46 = n88 ;
  assign y47 = n89 ;
  assign y48 = n91 ;
  assign y49 = n92 ;
  assign y50 = n93 ;
  assign y51 = n94 ;
  assign y52 = n95 ;
  assign y53 = n96 ;
  assign y54 = n97 ;
  assign y55 = n98 ;
  assign y56 = n99 ;
  assign y57 = n100 ;
  assign y58 = n101 ;
  assign y59 = n102 ;
  assign y60 = n103 ;
  assign y61 = n104 ;
  assign y62 = n105 ;
  assign y63 = n106 ;
  assign y64 = n108 ;
  assign y65 = n109 ;
  assign y66 = n110 ;
  assign y67 = n111 ;
  assign y68 = n112 ;
  assign y69 = n113 ;
  assign y70 = n114 ;
  assign y71 = n115 ;
  assign y72 = n116 ;
  assign y73 = n117 ;
  assign y74 = n118 ;
  assign y75 = n119 ;
  assign y76 = n120 ;
  assign y77 = n121 ;
  assign y78 = n122 ;
  assign y79 = n123 ;
  assign y80 = n125 ;
  assign y81 = n126 ;
  assign y82 = n127 ;
  assign y83 = n128 ;
  assign y84 = n129 ;
  assign y85 = n130 ;
  assign y86 = n131 ;
  assign y87 = n132 ;
  assign y88 = n133 ;
  assign y89 = n134 ;
  assign y90 = n135 ;
  assign y91 = n136 ;
  assign y92 = n137 ;
  assign y93 = n138 ;
  assign y94 = n139 ;
  assign y95 = n140 ;
  assign y96 = n142 ;
  assign y97 = n143 ;
  assign y98 = n144 ;
  assign y99 = n145 ;
  assign y100 = n146 ;
  assign y101 = n147 ;
  assign y102 = n148 ;
  assign y103 = n149 ;
  assign y104 = n150 ;
  assign y105 = n151 ;
  assign y106 = n152 ;
  assign y107 = n153 ;
  assign y108 = n154 ;
  assign y109 = n155 ;
  assign y110 = n156 ;
  assign y111 = n157 ;
  assign y112 = n159 ;
  assign y113 = n160 ;
  assign y114 = n161 ;
  assign y115 = n162 ;
  assign y116 = n163 ;
  assign y117 = n164 ;
  assign y118 = n165 ;
  assign y119 = n166 ;
  assign y120 = n167 ;
  assign y121 = n168 ;
  assign y122 = n169 ;
  assign y123 = n170 ;
  assign y124 = n171 ;
  assign y125 = n172 ;
  assign y126 = n173 ;
  assign y127 = n174 ;
  assign y128 = n178 ;
  assign y129 = n179 ;
  assign y130 = n180 ;
  assign y131 = n181 ;
  assign y132 = n182 ;
  assign y133 = n183 ;
  assign y134 = n184 ;
  assign y135 = n185 ;
  assign y136 = n186 ;
  assign y137 = n187 ;
  assign y138 = n188 ;
  assign y139 = n189 ;
  assign y140 = n190 ;
  assign y141 = n191 ;
  assign y142 = n192 ;
  assign y143 = n193 ;
  assign y144 = n195 ;
  assign y145 = n196 ;
  assign y146 = n197 ;
  assign y147 = n198 ;
  assign y148 = n199 ;
  assign y149 = n200 ;
  assign y150 = n201 ;
  assign y151 = n202 ;
  assign y152 = n203 ;
  assign y153 = n204 ;
  assign y154 = n205 ;
  assign y155 = n206 ;
  assign y156 = n207 ;
  assign y157 = n208 ;
  assign y158 = n209 ;
  assign y159 = n210 ;
  assign y160 = n212 ;
  assign y161 = n213 ;
  assign y162 = n214 ;
  assign y163 = n215 ;
  assign y164 = n216 ;
  assign y165 = n217 ;
  assign y166 = n218 ;
  assign y167 = n219 ;
  assign y168 = n220 ;
  assign y169 = n221 ;
  assign y170 = n222 ;
  assign y171 = n223 ;
  assign y172 = n224 ;
  assign y173 = n225 ;
  assign y174 = n226 ;
  assign y175 = n227 ;
  assign y176 = n229 ;
  assign y177 = n230 ;
  assign y178 = n231 ;
  assign y179 = n232 ;
  assign y180 = n233 ;
  assign y181 = n234 ;
  assign y182 = n235 ;
  assign y183 = n236 ;
  assign y184 = n237 ;
  assign y185 = n238 ;
  assign y186 = n239 ;
  assign y187 = n240 ;
  assign y188 = n241 ;
  assign y189 = n242 ;
  assign y190 = n243 ;
  assign y191 = n244 ;
  assign y192 = n246 ;
  assign y193 = n247 ;
  assign y194 = n248 ;
  assign y195 = n249 ;
  assign y196 = n250 ;
  assign y197 = n251 ;
  assign y198 = n252 ;
  assign y199 = n253 ;
  assign y200 = n254 ;
  assign y201 = n255 ;
  assign y202 = n256 ;
  assign y203 = n257 ;
  assign y204 = n258 ;
  assign y205 = n259 ;
  assign y206 = n260 ;
  assign y207 = n261 ;
  assign y208 = n263 ;
  assign y209 = n264 ;
  assign y210 = n265 ;
  assign y211 = n266 ;
  assign y212 = n267 ;
  assign y213 = n268 ;
  assign y214 = n269 ;
  assign y215 = n270 ;
  assign y216 = n271 ;
  assign y217 = n272 ;
  assign y218 = n273 ;
  assign y219 = n274 ;
  assign y220 = n275 ;
  assign y221 = n276 ;
  assign y222 = n277 ;
  assign y223 = n278 ;
  assign y224 = n280 ;
  assign y225 = n281 ;
  assign y226 = n282 ;
  assign y227 = n283 ;
  assign y228 = n284 ;
  assign y229 = n285 ;
  assign y230 = n286 ;
  assign y231 = n287 ;
  assign y232 = n288 ;
  assign y233 = n289 ;
  assign y234 = n290 ;
  assign y235 = n291 ;
  assign y236 = n292 ;
  assign y237 = n293 ;
  assign y238 = n294 ;
  assign y239 = n295 ;
  assign y240 = n297 ;
  assign y241 = n298 ;
  assign y242 = n299 ;
  assign y243 = n300 ;
  assign y244 = n301 ;
  assign y245 = n302 ;
  assign y246 = n303 ;
  assign y247 = n304 ;
  assign y248 = n305 ;
  assign y249 = n306 ;
  assign y250 = n307 ;
  assign y251 = n308 ;
  assign y252 = n309 ;
  assign y253 = n310 ;
  assign y254 = n311 ;
  assign y255 = n312 ;
endmodule
