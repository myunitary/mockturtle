module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , y0 , y1 , y2 , y3 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 ;
  output y0 , y1 , y2 , y3 ;
  wire n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 ;
  assign n282 = x61 ^ x5 ;
  assign n322 = x62 ^ x6 ;
  assign n113 = x63 ^ x7 ;
  assign n297 = x70 ^ x14 ;
  assign n298 = x71 ^ x15 ;
  assign n315 = ~n297 & n298 ;
  assign n316 = n315 ^ n297 ;
  assign n283 = x67 ^ x11 ;
  assign n284 = x66 ^ x10 ;
  assign n285 = n283 & n284 ;
  assign n286 = x65 ^ x9 ;
  assign n287 = x64 ^ x8 ;
  assign n288 = n286 & n287 ;
  assign n289 = n288 ^ n286 ;
  assign n290 = n289 ^ n287 ;
  assign n291 = n285 & ~n290 ;
  assign n292 = x69 ^ x13 ;
  assign n293 = x68 ^ x12 ;
  assign n294 = n292 & n293 ;
  assign n317 = n291 & n294 ;
  assign n318 = n316 & n317 ;
  assign n305 = n286 & ~n287 ;
  assign n306 = n305 ^ n287 ;
  assign n319 = n318 ^ n306 ;
  assign n320 = ~n113 & n319 ;
  assign n301 = n292 & ~n293 ;
  assign n302 = n301 ^ n293 ;
  assign n295 = n294 ^ n292 ;
  assign n296 = n295 ^ n293 ;
  assign n299 = n297 & n298 ;
  assign n300 = ~n296 & n299 ;
  assign n303 = n302 ^ n300 ;
  assign n304 = n291 & n303 ;
  assign n307 = n306 ^ n304 ;
  assign n308 = n306 ^ n113 ;
  assign n309 = ~n113 & n308 ;
  assign n310 = n309 ^ n113 ;
  assign n311 = n310 ^ n304 ;
  assign n312 = n307 & n311 ;
  assign n313 = n312 ^ n309 ;
  assign n314 = n313 ^ n304 ;
  assign n321 = n320 ^ n314 ;
  assign n323 = n322 ^ n321 ;
  assign n342 = n282 & n323 ;
  assign n344 = n314 & n320 ;
  assign n343 = n321 & n322 ;
  assign n345 = n344 ^ n343 ;
  assign n363 = n342 & n345 ;
  assign n364 = n343 & n344 ;
  assign n379 = n363 & n364 ;
  assign n281 = x60 ^ x4 ;
  assign n324 = n323 ^ n282 ;
  assign n341 = n281 & n324 ;
  assign n346 = n345 ^ n342 ;
  assign n362 = n341 & n346 ;
  assign n365 = n364 ^ n363 ;
  assign n378 = n362 & n365 ;
  assign n380 = n379 ^ n378 ;
  assign n280 = x59 ^ x3 ;
  assign n325 = n324 ^ n281 ;
  assign n340 = n280 & n325 ;
  assign n347 = n346 ^ n341 ;
  assign n361 = n340 & n347 ;
  assign n366 = n365 ^ n362 ;
  assign n377 = n361 & n366 ;
  assign n381 = n380 ^ n377 ;
  assign n252 = x73 ^ x17 ;
  assign n253 = x72 ^ x16 ;
  assign n275 = n252 & ~n253 ;
  assign n276 = n275 ^ n253 ;
  assign n254 = ~n252 & ~n253 ;
  assign n255 = x75 ^ x19 ;
  assign n256 = x74 ^ x18 ;
  assign n273 = n255 & n256 ;
  assign n274 = n254 & n273 ;
  assign n277 = n276 ^ n274 ;
  assign n257 = ~n255 & n256 ;
  assign n258 = n254 & n257 ;
  assign n259 = x77 ^ x21 ;
  assign n260 = x76 ^ x20 ;
  assign n270 = n259 & n260 ;
  assign n261 = ~n259 & n260 ;
  assign n262 = x79 ^ x23 ;
  assign n263 = x78 ^ x22 ;
  assign n267 = n262 & ~n263 ;
  assign n268 = n267 ^ n263 ;
  assign n269 = n261 & n268 ;
  assign n271 = n270 ^ n269 ;
  assign n272 = n258 & n271 ;
  assign n278 = n277 ^ n272 ;
  assign n264 = ~n262 & ~n263 ;
  assign n265 = n261 & n264 ;
  assign n266 = n258 & n265 ;
  assign n279 = n278 ^ n266 ;
  assign n326 = n325 ^ n280 ;
  assign n338 = n279 & n326 ;
  assign n339 = n338 ^ n326 ;
  assign n348 = n347 ^ n340 ;
  assign n360 = n339 & n348 ;
  assign n367 = n366 ^ n361 ;
  assign n376 = n360 & n367 ;
  assign n382 = n381 ^ n376 ;
  assign n167 = x80 ^ x24 ;
  assign n195 = x88 ^ x32 ;
  assign n169 = x92 ^ x36 ;
  assign n173 = x94 ^ x38 ;
  assign n174 = x93 ^ x37 ;
  assign n175 = n173 & n174 ;
  assign n176 = n175 ^ n174 ;
  assign n177 = n176 ^ n173 ;
  assign n183 = n169 & n177 ;
  assign n184 = n183 ^ n177 ;
  assign n185 = n184 ^ n177 ;
  assign n168 = x91 ^ x35 ;
  assign n170 = n169 ^ n168 ;
  assign n171 = ~n168 & ~n170 ;
  assign n172 = n171 ^ n168 ;
  assign n178 = n177 ^ n172 ;
  assign n179 = n177 ^ n169 ;
  assign n180 = ~n178 & n179 ;
  assign n181 = n180 ^ n171 ;
  assign n182 = n181 ^ n177 ;
  assign n186 = n185 ^ n182 ;
  assign n187 = x90 ^ x34 ;
  assign n191 = ~n186 & n187 ;
  assign n192 = n191 ^ n187 ;
  assign n193 = n192 ^ n186 ;
  assign n188 = x89 ^ x33 ;
  assign n189 = ~n187 & n188 ;
  assign n190 = n186 & n189 ;
  assign n194 = n193 ^ n190 ;
  assign n196 = n195 ^ n194 ;
  assign n248 = ~n167 & n196 ;
  assign n197 = n196 ^ n167 ;
  assign n198 = x81 ^ x25 ;
  assign n245 = n193 ^ n188 ;
  assign n246 = ~n198 & n245 ;
  assign n247 = ~n197 & n246 ;
  assign n249 = n248 ^ n247 ;
  assign n199 = n198 ^ n188 ;
  assign n200 = n199 ^ n193 ;
  assign n201 = ~n197 & ~n200 ;
  assign n231 = x82 ^ x26 ;
  assign n232 = n187 ^ n186 ;
  assign n242 = ~n231 & n232 ;
  assign n233 = n232 ^ n231 ;
  assign n234 = n185 ^ n168 ;
  assign n235 = x83 ^ x27 ;
  assign n240 = ~n234 & ~n235 ;
  assign n241 = ~n233 & n240 ;
  assign n243 = n242 ^ n241 ;
  assign n244 = n201 & n243 ;
  assign n250 = n249 ^ n244 ;
  assign n211 = x84 ^ x28 ;
  assign n228 = n179 & ~n211 ;
  assign n212 = n211 ^ n179 ;
  assign n214 = n174 ^ n173 ;
  assign n215 = x85 ^ x29 ;
  assign n226 = ~n214 & ~n215 ;
  assign n227 = ~n212 & n226 ;
  assign n229 = n228 ^ n227 ;
  assign n202 = x86 ^ x30 ;
  assign n209 = ~n173 & ~n202 ;
  assign n203 = n202 ^ n173 ;
  assign n204 = x87 ^ x31 ;
  assign n205 = x95 ^ x39 ;
  assign n206 = n204 & n205 ;
  assign n207 = n206 ^ n205 ;
  assign n208 = n203 & n207 ;
  assign n210 = n209 ^ n208 ;
  assign n213 = n212 ^ n210 ;
  assign n216 = n215 ^ n214 ;
  assign n217 = n216 ^ n212 ;
  assign n218 = n216 & n217 ;
  assign n219 = n218 ^ n216 ;
  assign n220 = n219 ^ n217 ;
  assign n221 = n220 ^ n212 ;
  assign n222 = n213 & ~n221 ;
  assign n223 = n222 ^ n221 ;
  assign n224 = n223 ^ n220 ;
  assign n225 = n224 ^ n210 ;
  assign n230 = n229 ^ n225 ;
  assign n236 = n235 ^ n234 ;
  assign n237 = ~n233 & n236 ;
  assign n238 = n230 & n237 ;
  assign n239 = n201 & n238 ;
  assign n251 = n250 ^ n239 ;
  assign n327 = n326 ^ n279 ;
  assign n336 = n251 & n327 ;
  assign n337 = n336 ^ n251 ;
  assign n349 = n348 ^ n339 ;
  assign n359 = n337 & n349 ;
  assign n368 = n367 ^ n360 ;
  assign n375 = n359 & n368 ;
  assign n383 = n382 ^ n375 ;
  assign n143 = x97 ^ x41 ;
  assign n144 = x96 ^ x40 ;
  assign n162 = n143 & ~n144 ;
  assign n163 = n162 ^ n144 ;
  assign n145 = ~n143 & ~n144 ;
  assign n146 = x98 ^ x42 ;
  assign n161 = n145 & n146 ;
  assign n164 = n163 ^ n161 ;
  assign n147 = x99 ^ x43 ;
  assign n148 = ~n146 & n147 ;
  assign n149 = n145 & n148 ;
  assign n150 = x101 ^ x45 ;
  assign n151 = x100 ^ x44 ;
  assign n152 = n150 & n151 ;
  assign n153 = x103 ^ x47 ;
  assign n154 = x102 ^ x46 ;
  assign n158 = n153 & n154 ;
  assign n159 = n152 & n158 ;
  assign n160 = n149 & n159 ;
  assign n165 = n164 ^ n160 ;
  assign n155 = ~n153 & n154 ;
  assign n156 = n152 & n155 ;
  assign n157 = n149 & n156 ;
  assign n166 = n165 ^ n157 ;
  assign n328 = n327 ^ n251 ;
  assign n333 = n166 & n328 ;
  assign n334 = n333 ^ n166 ;
  assign n335 = n334 ^ n328 ;
  assign n350 = n349 ^ n337 ;
  assign n357 = n335 & n350 ;
  assign n358 = n357 ^ n350 ;
  assign n369 = n368 ^ n359 ;
  assign n374 = n358 & n369 ;
  assign n384 = n383 ^ n374 ;
  assign n114 = x105 ^ x49 ;
  assign n115 = x104 ^ x48 ;
  assign n116 = ~n114 & ~n115 ;
  assign n117 = x107 ^ x51 ;
  assign n118 = x106 ^ x50 ;
  assign n119 = ~n117 & ~n118 ;
  assign n120 = n116 & n119 ;
  assign n124 = x109 ^ x53 ;
  assign n125 = x108 ^ x52 ;
  assign n128 = n124 & ~n125 ;
  assign n129 = n128 ^ n125 ;
  assign n140 = n120 & n129 ;
  assign n135 = n114 & ~n115 ;
  assign n136 = n135 ^ n115 ;
  assign n132 = n117 & ~n118 ;
  assign n133 = n132 ^ n118 ;
  assign n134 = n116 & n133 ;
  assign n137 = n136 ^ n134 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n113 & n141 ;
  assign n329 = n328 ^ n166 ;
  assign n332 = n142 & n329 ;
  assign n351 = n350 ^ n335 ;
  assign n355 = n332 & n351 ;
  assign n356 = n355 ^ n332 ;
  assign n370 = n369 ^ n358 ;
  assign n373 = n356 & n370 ;
  assign n385 = n384 ^ n373 ;
  assign n121 = x111 ^ x55 ;
  assign n122 = x110 ^ x54 ;
  assign n123 = n121 & n122 ;
  assign n126 = ~n124 & ~n125 ;
  assign n127 = n123 & n126 ;
  assign n130 = n129 ^ n127 ;
  assign n131 = n120 & n130 ;
  assign n138 = n137 ^ n131 ;
  assign n139 = ~n113 & n138 ;
  assign n330 = n329 ^ n142 ;
  assign n331 = n139 & n330 ;
  assign n352 = n351 ^ n332 ;
  assign n353 = n331 & n352 ;
  assign n354 = n353 ^ n331 ;
  assign n371 = n370 ^ n356 ;
  assign n372 = n354 & n371 ;
  assign n386 = n385 ^ n372 ;
  assign n387 = n371 ^ n354 ;
  assign n388 = n352 ^ n331 ;
  assign n389 = n330 ^ n139 ;
  assign y0 = n386 ;
  assign y1 = n387 ;
  assign y2 = ~n388 ;
  assign y3 = n389 ;
endmodule
