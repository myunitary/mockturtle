module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 ;
  assign n257 = x0 & ~x8 ;
  assign n222 = x8 ^ x0 ;
  assign n255 = x1 & ~x9 ;
  assign n256 = ~n222 & n255 ;
  assign n258 = n257 ^ n256 ;
  assign n223 = x9 ^ x1 ;
  assign n224 = ~n222 & ~n223 ;
  assign n252 = x2 & ~x10 ;
  assign n225 = x10 ^ x2 ;
  assign n250 = x3 & ~x11 ;
  assign n251 = ~n225 & n250 ;
  assign n253 = n252 ^ n251 ;
  assign n254 = n224 & n253 ;
  assign n259 = n258 ^ n254 ;
  assign n226 = x11 ^ x3 ;
  assign n227 = ~n225 & ~n226 ;
  assign n228 = n224 & n227 ;
  assign n246 = x4 & ~x12 ;
  assign n229 = x12 ^ x4 ;
  assign n244 = x5 & ~x13 ;
  assign n245 = ~n229 & n244 ;
  assign n247 = n246 ^ n245 ;
  assign n230 = x13 ^ x5 ;
  assign n231 = ~n229 & ~n230 ;
  assign n241 = x6 & ~x14 ;
  assign n232 = x14 ^ x6 ;
  assign n237 = x7 & x15 ;
  assign n238 = n237 ^ x7 ;
  assign n239 = n232 & n238 ;
  assign n240 = n239 ^ n238 ;
  assign n242 = n241 ^ n240 ;
  assign n243 = n231 & n242 ;
  assign n248 = n247 ^ n243 ;
  assign n249 = n228 & n248 ;
  assign n260 = n259 ^ n249 ;
  assign n233 = x15 ^ x7 ;
  assign n234 = ~n232 & ~n233 ;
  assign n235 = n231 & n234 ;
  assign n236 = n228 & n235 ;
  assign n261 = n260 ^ n236 ;
  assign n441 = x0 & ~n261 ;
  assign n440 = x8 & n261 ;
  assign n442 = n441 ^ n440 ;
  assign n263 = x8 & ~n261 ;
  assign n262 = x0 & n261 ;
  assign n264 = n263 ^ n262 ;
  assign n127 = x16 & ~x24 ;
  assign n92 = x24 ^ x16 ;
  assign n125 = x17 & ~x25 ;
  assign n126 = ~n92 & n125 ;
  assign n128 = n127 ^ n126 ;
  assign n93 = x25 ^ x17 ;
  assign n94 = ~n92 & ~n93 ;
  assign n122 = x18 & ~x26 ;
  assign n95 = x26 ^ x18 ;
  assign n120 = x19 & ~x27 ;
  assign n121 = ~n95 & n120 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = n94 & n123 ;
  assign n129 = n128 ^ n124 ;
  assign n96 = x27 ^ x19 ;
  assign n97 = ~n95 & ~n96 ;
  assign n98 = n94 & n97 ;
  assign n116 = x20 & ~x28 ;
  assign n99 = x28 ^ x20 ;
  assign n114 = x21 & ~x29 ;
  assign n115 = ~n99 & n114 ;
  assign n117 = n116 ^ n115 ;
  assign n100 = x29 ^ x21 ;
  assign n101 = ~n99 & ~n100 ;
  assign n111 = x22 & ~x30 ;
  assign n102 = x30 ^ x22 ;
  assign n107 = x23 & x31 ;
  assign n108 = n107 ^ x23 ;
  assign n109 = n102 & n108 ;
  assign n110 = n109 ^ n108 ;
  assign n112 = n111 ^ n110 ;
  assign n113 = n101 & n112 ;
  assign n118 = n117 ^ n113 ;
  assign n119 = n98 & n118 ;
  assign n130 = n129 ^ n119 ;
  assign n103 = x31 ^ x23 ;
  assign n104 = ~n102 & ~n103 ;
  assign n105 = n101 & n104 ;
  assign n106 = n98 & n105 ;
  assign n131 = n130 ^ n106 ;
  assign n266 = x16 & ~n131 ;
  assign n265 = x24 & n131 ;
  assign n267 = n266 ^ n265 ;
  assign n345 = n264 & ~n267 ;
  assign n268 = n267 ^ n264 ;
  assign n270 = x17 & ~n131 ;
  assign n269 = x25 & n131 ;
  assign n271 = n270 ^ n269 ;
  assign n273 = x9 & ~n261 ;
  assign n272 = x1 & n261 ;
  assign n274 = n273 ^ n272 ;
  assign n343 = ~n271 & n274 ;
  assign n344 = ~n268 & n343 ;
  assign n346 = n345 ^ n344 ;
  assign n275 = n274 ^ n271 ;
  assign n276 = ~n268 & ~n275 ;
  assign n278 = x10 & ~n261 ;
  assign n277 = x2 & n261 ;
  assign n279 = n278 ^ n277 ;
  assign n281 = x18 & ~n131 ;
  assign n280 = x26 & n131 ;
  assign n282 = n281 ^ n280 ;
  assign n340 = n279 & ~n282 ;
  assign n283 = n282 ^ n279 ;
  assign n285 = x11 & ~n261 ;
  assign n284 = x3 & n261 ;
  assign n286 = n285 ^ n284 ;
  assign n288 = x19 & ~n131 ;
  assign n287 = x27 & n131 ;
  assign n289 = n288 ^ n287 ;
  assign n338 = n286 & ~n289 ;
  assign n339 = ~n283 & n338 ;
  assign n341 = n340 ^ n339 ;
  assign n342 = n276 & n341 ;
  assign n347 = n346 ^ n342 ;
  assign n290 = n289 ^ n286 ;
  assign n291 = ~n283 & ~n290 ;
  assign n292 = n276 & n291 ;
  assign n294 = x12 & ~n261 ;
  assign n293 = x4 & n261 ;
  assign n295 = n294 ^ n293 ;
  assign n297 = x20 & ~n131 ;
  assign n296 = x28 & n131 ;
  assign n298 = n297 ^ n296 ;
  assign n334 = n295 & ~n298 ;
  assign n299 = n298 ^ n295 ;
  assign n301 = x13 & ~n261 ;
  assign n300 = x5 & n261 ;
  assign n302 = n301 ^ n300 ;
  assign n304 = x21 & ~n131 ;
  assign n303 = x29 & n131 ;
  assign n305 = n304 ^ n303 ;
  assign n332 = n302 & ~n305 ;
  assign n333 = ~n299 & n332 ;
  assign n335 = n334 ^ n333 ;
  assign n306 = n305 ^ n302 ;
  assign n307 = ~n299 & ~n306 ;
  assign n309 = x14 & ~n261 ;
  assign n308 = x6 & n261 ;
  assign n310 = n309 ^ n308 ;
  assign n312 = x22 & ~n131 ;
  assign n311 = x30 & n131 ;
  assign n313 = n312 ^ n311 ;
  assign n329 = n310 & ~n313 ;
  assign n314 = n313 ^ n310 ;
  assign n184 = x23 & n131 ;
  assign n315 = n184 ^ x23 ;
  assign n182 = x31 & n131 ;
  assign n316 = n315 ^ n182 ;
  assign n318 = x15 & n261 ;
  assign n319 = n318 ^ x15 ;
  assign n317 = x7 & n261 ;
  assign n320 = n319 ^ n317 ;
  assign n325 = n316 & n320 ;
  assign n326 = n325 ^ n320 ;
  assign n327 = n314 & n326 ;
  assign n328 = n327 ^ n326 ;
  assign n330 = n329 ^ n328 ;
  assign n331 = n307 & n330 ;
  assign n336 = n335 ^ n331 ;
  assign n337 = n292 & n336 ;
  assign n348 = n347 ^ n337 ;
  assign n321 = n320 ^ n316 ;
  assign n322 = ~n314 & ~n321 ;
  assign n323 = n307 & n322 ;
  assign n324 = n292 & n323 ;
  assign n349 = n348 ^ n324 ;
  assign n444 = n264 & ~n349 ;
  assign n443 = n267 & n349 ;
  assign n445 = n444 ^ n443 ;
  assign n521 = n442 & ~n445 ;
  assign n446 = n445 ^ n442 ;
  assign n448 = n274 & ~n349 ;
  assign n447 = n271 & n349 ;
  assign n449 = n448 ^ n447 ;
  assign n451 = x1 & ~n261 ;
  assign n450 = x9 & n261 ;
  assign n452 = n451 ^ n450 ;
  assign n519 = ~n449 & n452 ;
  assign n520 = ~n446 & n519 ;
  assign n522 = n521 ^ n520 ;
  assign n453 = n452 ^ n449 ;
  assign n454 = ~n446 & ~n453 ;
  assign n456 = x2 & ~n261 ;
  assign n455 = x10 & n261 ;
  assign n457 = n456 ^ n455 ;
  assign n459 = n279 & ~n349 ;
  assign n458 = n282 & n349 ;
  assign n460 = n459 ^ n458 ;
  assign n516 = n457 & ~n460 ;
  assign n461 = n460 ^ n457 ;
  assign n463 = x3 & ~n261 ;
  assign n462 = x11 & n261 ;
  assign n464 = n463 ^ n462 ;
  assign n466 = n286 & ~n349 ;
  assign n465 = n289 & n349 ;
  assign n467 = n466 ^ n465 ;
  assign n514 = n464 & ~n467 ;
  assign n515 = ~n461 & n514 ;
  assign n517 = n516 ^ n515 ;
  assign n518 = n454 & n517 ;
  assign n523 = n522 ^ n518 ;
  assign n468 = n467 ^ n464 ;
  assign n469 = ~n461 & ~n468 ;
  assign n470 = n454 & n469 ;
  assign n472 = x4 & ~n261 ;
  assign n471 = x12 & n261 ;
  assign n473 = n472 ^ n471 ;
  assign n475 = n295 & ~n349 ;
  assign n474 = n298 & n349 ;
  assign n476 = n475 ^ n474 ;
  assign n510 = n473 & ~n476 ;
  assign n477 = n476 ^ n473 ;
  assign n479 = x5 & ~n261 ;
  assign n478 = x13 & n261 ;
  assign n480 = n479 ^ n478 ;
  assign n482 = n302 & ~n349 ;
  assign n481 = n305 & n349 ;
  assign n483 = n482 ^ n481 ;
  assign n508 = n480 & ~n483 ;
  assign n509 = ~n477 & n508 ;
  assign n511 = n510 ^ n509 ;
  assign n484 = n483 ^ n480 ;
  assign n485 = ~n477 & ~n484 ;
  assign n487 = x6 & ~n261 ;
  assign n486 = x14 & n261 ;
  assign n488 = n487 ^ n486 ;
  assign n490 = n310 & ~n349 ;
  assign n489 = n313 & n349 ;
  assign n491 = n490 ^ n489 ;
  assign n505 = n488 & ~n491 ;
  assign n492 = n491 ^ n488 ;
  assign n402 = n320 & n349 ;
  assign n493 = n402 ^ n320 ;
  assign n400 = n316 & n349 ;
  assign n494 = n493 ^ n400 ;
  assign n495 = x7 & ~n261 ;
  assign n496 = n495 ^ n318 ;
  assign n501 = n494 & n496 ;
  assign n502 = n501 ^ n496 ;
  assign n503 = n492 & n502 ;
  assign n504 = n503 ^ n502 ;
  assign n506 = n505 ^ n504 ;
  assign n507 = n485 & n506 ;
  assign n512 = n511 ^ n507 ;
  assign n513 = n470 & n512 ;
  assign n524 = n523 ^ n513 ;
  assign n497 = n496 ^ n494 ;
  assign n498 = ~n492 & ~n497 ;
  assign n499 = n485 & n498 ;
  assign n500 = n470 & n499 ;
  assign n525 = n524 ^ n500 ;
  assign n617 = n442 & ~n525 ;
  assign n616 = n445 & n525 ;
  assign n618 = n617 ^ n616 ;
  assign n527 = n445 & ~n525 ;
  assign n526 = n442 & n525 ;
  assign n528 = n527 ^ n526 ;
  assign n351 = n267 & ~n349 ;
  assign n350 = n264 & n349 ;
  assign n352 = n351 ^ n350 ;
  assign n133 = x24 & ~n131 ;
  assign n132 = x16 & n131 ;
  assign n134 = n133 ^ n132 ;
  assign n84 = x32 & ~x40 ;
  assign n49 = x40 ^ x32 ;
  assign n82 = x33 & ~x41 ;
  assign n83 = ~n49 & n82 ;
  assign n85 = n84 ^ n83 ;
  assign n50 = x41 ^ x33 ;
  assign n51 = ~n49 & ~n50 ;
  assign n79 = x34 & ~x42 ;
  assign n52 = x42 ^ x34 ;
  assign n77 = x35 & ~x43 ;
  assign n78 = ~n52 & n77 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n51 & n80 ;
  assign n86 = n85 ^ n81 ;
  assign n53 = x43 ^ x35 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n51 & n54 ;
  assign n73 = x36 & ~x44 ;
  assign n56 = x44 ^ x36 ;
  assign n71 = x37 & ~x45 ;
  assign n72 = ~n56 & n71 ;
  assign n74 = n73 ^ n72 ;
  assign n57 = x45 ^ x37 ;
  assign n58 = ~n56 & ~n57 ;
  assign n68 = x38 & ~x46 ;
  assign n59 = x46 ^ x38 ;
  assign n64 = x39 & x47 ;
  assign n65 = n64 ^ x39 ;
  assign n66 = n59 & n65 ;
  assign n67 = n66 ^ n65 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n58 & n69 ;
  assign n75 = n74 ^ n70 ;
  assign n76 = n55 & n75 ;
  assign n87 = n86 ^ n76 ;
  assign n60 = x47 ^ x39 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = n58 & n61 ;
  assign n63 = n55 & n62 ;
  assign n88 = n87 ^ n63 ;
  assign n90 = x32 & ~n88 ;
  assign n89 = x40 & n88 ;
  assign n91 = n90 ^ n89 ;
  assign n214 = ~n91 & n134 ;
  assign n135 = n134 ^ n91 ;
  assign n137 = x25 & ~n131 ;
  assign n136 = x17 & n131 ;
  assign n138 = n137 ^ n136 ;
  assign n140 = x33 & ~n88 ;
  assign n139 = x41 & n88 ;
  assign n141 = n140 ^ n139 ;
  assign n212 = n138 & ~n141 ;
  assign n213 = ~n135 & n212 ;
  assign n215 = n214 ^ n213 ;
  assign n142 = n141 ^ n138 ;
  assign n143 = ~n135 & ~n142 ;
  assign n145 = x26 & ~n131 ;
  assign n144 = x18 & n131 ;
  assign n146 = n145 ^ n144 ;
  assign n148 = x34 & ~n88 ;
  assign n147 = x42 & n88 ;
  assign n149 = n148 ^ n147 ;
  assign n209 = n146 & ~n149 ;
  assign n150 = n149 ^ n146 ;
  assign n152 = x27 & ~n131 ;
  assign n151 = x19 & n131 ;
  assign n153 = n152 ^ n151 ;
  assign n155 = x35 & ~n88 ;
  assign n154 = x43 & n88 ;
  assign n156 = n155 ^ n154 ;
  assign n207 = n153 & ~n156 ;
  assign n208 = ~n150 & n207 ;
  assign n210 = n209 ^ n208 ;
  assign n211 = n143 & n210 ;
  assign n216 = n215 ^ n211 ;
  assign n157 = n156 ^ n153 ;
  assign n158 = ~n150 & ~n157 ;
  assign n159 = n143 & n158 ;
  assign n161 = x28 & ~n131 ;
  assign n160 = x20 & n131 ;
  assign n162 = n161 ^ n160 ;
  assign n164 = x36 & ~n88 ;
  assign n163 = x44 & n88 ;
  assign n165 = n164 ^ n163 ;
  assign n203 = n162 & ~n165 ;
  assign n166 = n165 ^ n162 ;
  assign n168 = x29 & ~n131 ;
  assign n167 = x21 & n131 ;
  assign n169 = n168 ^ n167 ;
  assign n171 = x37 & ~n88 ;
  assign n170 = x45 & n88 ;
  assign n172 = n171 ^ n170 ;
  assign n201 = n169 & ~n172 ;
  assign n202 = ~n166 & n201 ;
  assign n204 = n203 ^ n202 ;
  assign n173 = n172 ^ n169 ;
  assign n174 = ~n166 & ~n173 ;
  assign n176 = x30 & ~n131 ;
  assign n175 = x22 & n131 ;
  assign n177 = n176 ^ n175 ;
  assign n179 = x38 & ~n88 ;
  assign n178 = x46 & n88 ;
  assign n180 = n179 ^ n178 ;
  assign n198 = n177 & ~n180 ;
  assign n181 = n180 ^ n177 ;
  assign n183 = n182 ^ x31 ;
  assign n185 = n184 ^ n183 ;
  assign n187 = x39 & n88 ;
  assign n188 = n187 ^ x39 ;
  assign n186 = x47 & n88 ;
  assign n189 = n188 ^ n186 ;
  assign n194 = n185 & n189 ;
  assign n195 = n194 ^ n185 ;
  assign n196 = n181 & n195 ;
  assign n197 = n196 ^ n195 ;
  assign n199 = n198 ^ n197 ;
  assign n200 = n174 & n199 ;
  assign n205 = n204 ^ n200 ;
  assign n206 = n159 & n205 ;
  assign n217 = n216 ^ n206 ;
  assign n190 = n189 ^ n185 ;
  assign n191 = ~n181 & ~n190 ;
  assign n192 = n174 & n191 ;
  assign n193 = n159 & n192 ;
  assign n218 = n217 ^ n193 ;
  assign n220 = n134 & ~n218 ;
  assign n219 = n91 & n218 ;
  assign n221 = n220 ^ n219 ;
  assign n432 = ~n221 & n352 ;
  assign n353 = n352 ^ n221 ;
  assign n355 = n271 & ~n349 ;
  assign n354 = n274 & n349 ;
  assign n356 = n355 ^ n354 ;
  assign n358 = n138 & ~n218 ;
  assign n357 = n141 & n218 ;
  assign n359 = n358 ^ n357 ;
  assign n430 = n356 & ~n359 ;
  assign n431 = ~n353 & n430 ;
  assign n433 = n432 ^ n431 ;
  assign n360 = n359 ^ n356 ;
  assign n361 = ~n353 & ~n360 ;
  assign n363 = n282 & ~n349 ;
  assign n362 = n279 & n349 ;
  assign n364 = n363 ^ n362 ;
  assign n366 = n146 & ~n218 ;
  assign n365 = n149 & n218 ;
  assign n367 = n366 ^ n365 ;
  assign n427 = n364 & ~n367 ;
  assign n368 = n367 ^ n364 ;
  assign n370 = n289 & ~n349 ;
  assign n369 = n286 & n349 ;
  assign n371 = n370 ^ n369 ;
  assign n373 = n153 & ~n218 ;
  assign n372 = n156 & n218 ;
  assign n374 = n373 ^ n372 ;
  assign n425 = n371 & ~n374 ;
  assign n426 = ~n368 & n425 ;
  assign n428 = n427 ^ n426 ;
  assign n429 = n361 & n428 ;
  assign n434 = n433 ^ n429 ;
  assign n375 = n374 ^ n371 ;
  assign n376 = ~n368 & ~n375 ;
  assign n377 = n361 & n376 ;
  assign n379 = n298 & ~n349 ;
  assign n378 = n295 & n349 ;
  assign n380 = n379 ^ n378 ;
  assign n382 = n162 & ~n218 ;
  assign n381 = n165 & n218 ;
  assign n383 = n382 ^ n381 ;
  assign n421 = n380 & ~n383 ;
  assign n384 = n383 ^ n380 ;
  assign n386 = n305 & ~n349 ;
  assign n385 = n302 & n349 ;
  assign n387 = n386 ^ n385 ;
  assign n389 = n169 & ~n218 ;
  assign n388 = n172 & n218 ;
  assign n390 = n389 ^ n388 ;
  assign n419 = n387 & ~n390 ;
  assign n420 = ~n384 & n419 ;
  assign n422 = n421 ^ n420 ;
  assign n391 = n390 ^ n387 ;
  assign n392 = ~n384 & ~n391 ;
  assign n394 = n313 & ~n349 ;
  assign n393 = n310 & n349 ;
  assign n395 = n394 ^ n393 ;
  assign n397 = n177 & ~n218 ;
  assign n396 = n180 & n218 ;
  assign n398 = n397 ^ n396 ;
  assign n416 = n395 & ~n398 ;
  assign n399 = n398 ^ n395 ;
  assign n401 = n400 ^ n316 ;
  assign n403 = n402 ^ n401 ;
  assign n405 = n185 & n218 ;
  assign n406 = n405 ^ n185 ;
  assign n404 = n189 & n218 ;
  assign n407 = n406 ^ n404 ;
  assign n412 = n403 & n407 ;
  assign n413 = n412 ^ n403 ;
  assign n414 = n399 & n413 ;
  assign n415 = n414 ^ n413 ;
  assign n417 = n416 ^ n415 ;
  assign n418 = n392 & n417 ;
  assign n423 = n422 ^ n418 ;
  assign n424 = n377 & n423 ;
  assign n435 = n434 ^ n424 ;
  assign n408 = n407 ^ n403 ;
  assign n409 = ~n399 & ~n408 ;
  assign n410 = n392 & n409 ;
  assign n411 = n377 & n410 ;
  assign n436 = n435 ^ n411 ;
  assign n438 = n352 & ~n436 ;
  assign n437 = n221 & n436 ;
  assign n439 = n438 ^ n437 ;
  assign n608 = ~n439 & n528 ;
  assign n529 = n528 ^ n439 ;
  assign n531 = n449 & ~n525 ;
  assign n530 = n452 & n525 ;
  assign n532 = n531 ^ n530 ;
  assign n534 = n356 & ~n436 ;
  assign n533 = n359 & n436 ;
  assign n535 = n534 ^ n533 ;
  assign n606 = n532 & ~n535 ;
  assign n607 = ~n529 & n606 ;
  assign n609 = n608 ^ n607 ;
  assign n536 = n535 ^ n532 ;
  assign n537 = ~n529 & ~n536 ;
  assign n539 = n460 & ~n525 ;
  assign n538 = n457 & n525 ;
  assign n540 = n539 ^ n538 ;
  assign n542 = n364 & ~n436 ;
  assign n541 = n367 & n436 ;
  assign n543 = n542 ^ n541 ;
  assign n603 = n540 & ~n543 ;
  assign n544 = n543 ^ n540 ;
  assign n546 = n467 & ~n525 ;
  assign n545 = n464 & n525 ;
  assign n547 = n546 ^ n545 ;
  assign n549 = n371 & ~n436 ;
  assign n548 = n374 & n436 ;
  assign n550 = n549 ^ n548 ;
  assign n601 = n547 & ~n550 ;
  assign n602 = ~n544 & n601 ;
  assign n604 = n603 ^ n602 ;
  assign n605 = n537 & n604 ;
  assign n610 = n609 ^ n605 ;
  assign n551 = n550 ^ n547 ;
  assign n552 = ~n544 & ~n551 ;
  assign n553 = n537 & n552 ;
  assign n555 = n476 & ~n525 ;
  assign n554 = n473 & n525 ;
  assign n556 = n555 ^ n554 ;
  assign n558 = n380 & ~n436 ;
  assign n557 = n383 & n436 ;
  assign n559 = n558 ^ n557 ;
  assign n597 = n556 & ~n559 ;
  assign n560 = n559 ^ n556 ;
  assign n562 = n483 & ~n525 ;
  assign n561 = n480 & n525 ;
  assign n563 = n562 ^ n561 ;
  assign n565 = n387 & ~n436 ;
  assign n564 = n390 & n436 ;
  assign n566 = n565 ^ n564 ;
  assign n595 = n563 & ~n566 ;
  assign n596 = ~n560 & n595 ;
  assign n598 = n597 ^ n596 ;
  assign n567 = n566 ^ n563 ;
  assign n568 = ~n560 & ~n567 ;
  assign n570 = n491 & ~n525 ;
  assign n569 = n488 & n525 ;
  assign n571 = n570 ^ n569 ;
  assign n573 = n395 & ~n436 ;
  assign n572 = n398 & n436 ;
  assign n574 = n573 ^ n572 ;
  assign n592 = n571 & ~n574 ;
  assign n575 = n574 ^ n571 ;
  assign n577 = n494 & n525 ;
  assign n578 = n577 ^ n494 ;
  assign n576 = n496 & n525 ;
  assign n579 = n578 ^ n576 ;
  assign n581 = n403 & n436 ;
  assign n582 = n581 ^ n403 ;
  assign n580 = n407 & n436 ;
  assign n583 = n582 ^ n580 ;
  assign n588 = n579 & n583 ;
  assign n589 = n588 ^ n579 ;
  assign n590 = n575 & n589 ;
  assign n591 = n590 ^ n589 ;
  assign n593 = n592 ^ n591 ;
  assign n594 = n568 & n593 ;
  assign n599 = n598 ^ n594 ;
  assign n600 = n553 & n599 ;
  assign n611 = n610 ^ n600 ;
  assign n584 = n583 ^ n579 ;
  assign n585 = ~n575 & ~n584 ;
  assign n586 = n568 & n585 ;
  assign n587 = n553 & n586 ;
  assign n612 = n611 ^ n587 ;
  assign n614 = n528 & ~n612 ;
  assign n613 = n439 & n612 ;
  assign n615 = n614 ^ n613 ;
  assign n696 = ~n615 & n618 ;
  assign n619 = n618 ^ n615 ;
  assign n621 = n452 & ~n525 ;
  assign n620 = n449 & n525 ;
  assign n622 = n621 ^ n620 ;
  assign n624 = n532 & ~n612 ;
  assign n623 = n535 & n612 ;
  assign n625 = n624 ^ n623 ;
  assign n694 = n622 & ~n625 ;
  assign n695 = ~n619 & n694 ;
  assign n697 = n696 ^ n695 ;
  assign n626 = n625 ^ n622 ;
  assign n627 = ~n619 & ~n626 ;
  assign n629 = n457 & ~n525 ;
  assign n628 = n460 & n525 ;
  assign n630 = n629 ^ n628 ;
  assign n632 = n540 & ~n612 ;
  assign n631 = n543 & n612 ;
  assign n633 = n632 ^ n631 ;
  assign n691 = n630 & ~n633 ;
  assign n634 = n633 ^ n630 ;
  assign n636 = n464 & ~n525 ;
  assign n635 = n467 & n525 ;
  assign n637 = n636 ^ n635 ;
  assign n639 = n547 & ~n612 ;
  assign n638 = n550 & n612 ;
  assign n640 = n639 ^ n638 ;
  assign n689 = n637 & ~n640 ;
  assign n690 = ~n634 & n689 ;
  assign n692 = n691 ^ n690 ;
  assign n693 = n627 & n692 ;
  assign n698 = n697 ^ n693 ;
  assign n641 = n640 ^ n637 ;
  assign n642 = ~n634 & ~n641 ;
  assign n643 = n627 & n642 ;
  assign n645 = n473 & ~n525 ;
  assign n644 = n476 & n525 ;
  assign n646 = n645 ^ n644 ;
  assign n648 = n556 & ~n612 ;
  assign n647 = n559 & n612 ;
  assign n649 = n648 ^ n647 ;
  assign n685 = n646 & ~n649 ;
  assign n650 = n649 ^ n646 ;
  assign n652 = n480 & ~n525 ;
  assign n651 = n483 & n525 ;
  assign n653 = n652 ^ n651 ;
  assign n655 = n563 & ~n612 ;
  assign n654 = n566 & n612 ;
  assign n656 = n655 ^ n654 ;
  assign n683 = n653 & ~n656 ;
  assign n684 = ~n650 & n683 ;
  assign n686 = n685 ^ n684 ;
  assign n657 = n656 ^ n653 ;
  assign n658 = ~n650 & ~n657 ;
  assign n660 = n488 & ~n525 ;
  assign n659 = n491 & n525 ;
  assign n661 = n660 ^ n659 ;
  assign n663 = n571 & ~n612 ;
  assign n662 = n574 & n612 ;
  assign n664 = n663 ^ n662 ;
  assign n680 = n661 & ~n664 ;
  assign n665 = n664 ^ n661 ;
  assign n666 = n496 & ~n525 ;
  assign n667 = n666 ^ n577 ;
  assign n669 = n579 & n612 ;
  assign n670 = n669 ^ n579 ;
  assign n668 = n583 & n612 ;
  assign n671 = n670 ^ n668 ;
  assign n676 = n667 & n671 ;
  assign n677 = n676 ^ n667 ;
  assign n678 = n665 & n677 ;
  assign n679 = n678 ^ n677 ;
  assign n681 = n680 ^ n679 ;
  assign n682 = n658 & n681 ;
  assign n687 = n686 ^ n682 ;
  assign n688 = n643 & n687 ;
  assign n699 = n698 ^ n688 ;
  assign n672 = n671 ^ n667 ;
  assign n673 = ~n665 & ~n672 ;
  assign n674 = n658 & n673 ;
  assign n675 = n643 & n674 ;
  assign n700 = n699 ^ n675 ;
  assign n702 = n618 & n700 ;
  assign n703 = n702 ^ n618 ;
  assign n701 = n615 & n700 ;
  assign n704 = n703 ^ n701 ;
  assign n706 = n622 & n700 ;
  assign n707 = n706 ^ n622 ;
  assign n705 = n625 & n700 ;
  assign n708 = n707 ^ n705 ;
  assign n710 = n630 & n700 ;
  assign n711 = n710 ^ n630 ;
  assign n709 = n633 & n700 ;
  assign n712 = n711 ^ n709 ;
  assign n714 = n637 & n700 ;
  assign n715 = n714 ^ n637 ;
  assign n713 = n640 & n700 ;
  assign n716 = n715 ^ n713 ;
  assign n718 = n646 & n700 ;
  assign n719 = n718 ^ n646 ;
  assign n717 = n649 & n700 ;
  assign n720 = n719 ^ n717 ;
  assign n722 = n653 & n700 ;
  assign n723 = n722 ^ n653 ;
  assign n721 = n656 & n700 ;
  assign n724 = n723 ^ n721 ;
  assign n726 = n661 & n700 ;
  assign n727 = n726 ^ n661 ;
  assign n725 = n664 & n700 ;
  assign n728 = n727 ^ n725 ;
  assign n730 = n667 & n700 ;
  assign n731 = n730 ^ n667 ;
  assign n729 = n671 & n700 ;
  assign n732 = n731 ^ n729 ;
  assign n733 = n701 ^ n615 ;
  assign n734 = n733 ^ n702 ;
  assign n735 = n705 ^ n625 ;
  assign n736 = n735 ^ n706 ;
  assign n737 = n709 ^ n633 ;
  assign n738 = n737 ^ n710 ;
  assign n739 = n713 ^ n640 ;
  assign n740 = n739 ^ n714 ;
  assign n741 = n717 ^ n649 ;
  assign n742 = n741 ^ n718 ;
  assign n743 = n721 ^ n656 ;
  assign n744 = n743 ^ n722 ;
  assign n745 = n725 ^ n664 ;
  assign n746 = n745 ^ n726 ;
  assign n747 = n729 ^ n671 ;
  assign n748 = n747 ^ n730 ;
  assign n927 = n439 & ~n612 ;
  assign n926 = n528 & n612 ;
  assign n928 = n927 ^ n926 ;
  assign n839 = n221 & ~n436 ;
  assign n838 = n352 & n436 ;
  assign n840 = n839 ^ n838 ;
  assign n753 = n91 & ~n218 ;
  assign n752 = n134 & n218 ;
  assign n754 = n753 ^ n752 ;
  assign n750 = x40 & ~n88 ;
  assign n749 = x32 & n88 ;
  assign n751 = n750 ^ n749 ;
  assign n830 = ~n751 & n754 ;
  assign n755 = n754 ^ n751 ;
  assign n757 = n141 & ~n218 ;
  assign n756 = n138 & n218 ;
  assign n758 = n757 ^ n756 ;
  assign n760 = x41 & ~n88 ;
  assign n759 = x33 & n88 ;
  assign n761 = n760 ^ n759 ;
  assign n828 = n758 & ~n761 ;
  assign n829 = ~n755 & n828 ;
  assign n831 = n830 ^ n829 ;
  assign n762 = n761 ^ n758 ;
  assign n763 = ~n755 & ~n762 ;
  assign n765 = n149 & ~n218 ;
  assign n764 = n146 & n218 ;
  assign n766 = n765 ^ n764 ;
  assign n768 = x42 & ~n88 ;
  assign n767 = x34 & n88 ;
  assign n769 = n768 ^ n767 ;
  assign n825 = n766 & ~n769 ;
  assign n770 = n769 ^ n766 ;
  assign n772 = n156 & ~n218 ;
  assign n771 = n153 & n218 ;
  assign n773 = n772 ^ n771 ;
  assign n775 = x43 & ~n88 ;
  assign n774 = x35 & n88 ;
  assign n776 = n775 ^ n774 ;
  assign n823 = n773 & ~n776 ;
  assign n824 = ~n770 & n823 ;
  assign n826 = n825 ^ n824 ;
  assign n827 = n763 & n826 ;
  assign n832 = n831 ^ n827 ;
  assign n777 = n776 ^ n773 ;
  assign n778 = ~n770 & ~n777 ;
  assign n779 = n763 & n778 ;
  assign n781 = n165 & ~n218 ;
  assign n780 = n162 & n218 ;
  assign n782 = n781 ^ n780 ;
  assign n784 = x44 & ~n88 ;
  assign n783 = x36 & n88 ;
  assign n785 = n784 ^ n783 ;
  assign n819 = n782 & ~n785 ;
  assign n786 = n785 ^ n782 ;
  assign n788 = n172 & ~n218 ;
  assign n787 = n169 & n218 ;
  assign n789 = n788 ^ n787 ;
  assign n791 = x45 & ~n88 ;
  assign n790 = x37 & n88 ;
  assign n792 = n791 ^ n790 ;
  assign n817 = n789 & ~n792 ;
  assign n818 = ~n786 & n817 ;
  assign n820 = n819 ^ n818 ;
  assign n793 = n792 ^ n789 ;
  assign n794 = ~n786 & ~n793 ;
  assign n796 = n180 & ~n218 ;
  assign n795 = n177 & n218 ;
  assign n797 = n796 ^ n795 ;
  assign n799 = x46 & ~n88 ;
  assign n798 = x38 & n88 ;
  assign n800 = n799 ^ n798 ;
  assign n814 = n797 & ~n800 ;
  assign n801 = n800 ^ n797 ;
  assign n802 = n404 ^ n189 ;
  assign n803 = n802 ^ n405 ;
  assign n804 = x47 & ~n88 ;
  assign n805 = n804 ^ n187 ;
  assign n810 = n803 & n805 ;
  assign n811 = n810 ^ n803 ;
  assign n812 = n801 & n811 ;
  assign n813 = n812 ^ n811 ;
  assign n815 = n814 ^ n813 ;
  assign n816 = n794 & n815 ;
  assign n821 = n820 ^ n816 ;
  assign n822 = n779 & n821 ;
  assign n833 = n832 ^ n822 ;
  assign n806 = n805 ^ n803 ;
  assign n807 = ~n801 & ~n806 ;
  assign n808 = n794 & n807 ;
  assign n809 = n779 & n808 ;
  assign n834 = n833 ^ n809 ;
  assign n836 = n754 & ~n834 ;
  assign n835 = n751 & n834 ;
  assign n837 = n836 ^ n835 ;
  assign n918 = ~n837 & n840 ;
  assign n841 = n840 ^ n837 ;
  assign n843 = n359 & ~n436 ;
  assign n842 = n356 & n436 ;
  assign n844 = n843 ^ n842 ;
  assign n846 = n758 & ~n834 ;
  assign n845 = n761 & n834 ;
  assign n847 = n846 ^ n845 ;
  assign n916 = n844 & ~n847 ;
  assign n917 = ~n841 & n916 ;
  assign n919 = n918 ^ n917 ;
  assign n848 = n847 ^ n844 ;
  assign n849 = ~n841 & ~n848 ;
  assign n851 = n367 & ~n436 ;
  assign n850 = n364 & n436 ;
  assign n852 = n851 ^ n850 ;
  assign n854 = n766 & ~n834 ;
  assign n853 = n769 & n834 ;
  assign n855 = n854 ^ n853 ;
  assign n913 = n852 & ~n855 ;
  assign n856 = n855 ^ n852 ;
  assign n858 = n374 & ~n436 ;
  assign n857 = n371 & n436 ;
  assign n859 = n858 ^ n857 ;
  assign n861 = n773 & ~n834 ;
  assign n860 = n776 & n834 ;
  assign n862 = n861 ^ n860 ;
  assign n911 = n859 & ~n862 ;
  assign n912 = ~n856 & n911 ;
  assign n914 = n913 ^ n912 ;
  assign n915 = n849 & n914 ;
  assign n920 = n919 ^ n915 ;
  assign n863 = n862 ^ n859 ;
  assign n864 = ~n856 & ~n863 ;
  assign n865 = n849 & n864 ;
  assign n867 = n383 & ~n436 ;
  assign n866 = n380 & n436 ;
  assign n868 = n867 ^ n866 ;
  assign n870 = n782 & ~n834 ;
  assign n869 = n785 & n834 ;
  assign n871 = n870 ^ n869 ;
  assign n907 = n868 & ~n871 ;
  assign n872 = n871 ^ n868 ;
  assign n874 = n390 & ~n436 ;
  assign n873 = n387 & n436 ;
  assign n875 = n874 ^ n873 ;
  assign n877 = n789 & ~n834 ;
  assign n876 = n792 & n834 ;
  assign n878 = n877 ^ n876 ;
  assign n905 = n875 & ~n878 ;
  assign n906 = ~n872 & n905 ;
  assign n908 = n907 ^ n906 ;
  assign n879 = n878 ^ n875 ;
  assign n880 = ~n872 & ~n879 ;
  assign n882 = n398 & ~n436 ;
  assign n881 = n395 & n436 ;
  assign n883 = n882 ^ n881 ;
  assign n885 = n797 & ~n834 ;
  assign n884 = n800 & n834 ;
  assign n886 = n885 ^ n884 ;
  assign n902 = n883 & ~n886 ;
  assign n887 = n886 ^ n883 ;
  assign n888 = n580 ^ n407 ;
  assign n889 = n888 ^ n581 ;
  assign n891 = n803 & n834 ;
  assign n892 = n891 ^ n803 ;
  assign n890 = n805 & n834 ;
  assign n893 = n892 ^ n890 ;
  assign n898 = n889 & n893 ;
  assign n899 = n898 ^ n889 ;
  assign n900 = n887 & n899 ;
  assign n901 = n900 ^ n899 ;
  assign n903 = n902 ^ n901 ;
  assign n904 = n880 & n903 ;
  assign n909 = n908 ^ n904 ;
  assign n910 = n865 & n909 ;
  assign n921 = n920 ^ n910 ;
  assign n894 = n893 ^ n889 ;
  assign n895 = ~n887 & ~n894 ;
  assign n896 = n880 & n895 ;
  assign n897 = n865 & n896 ;
  assign n922 = n921 ^ n897 ;
  assign n924 = n840 & ~n922 ;
  assign n923 = n837 & n922 ;
  assign n925 = n924 ^ n923 ;
  assign n1006 = ~n925 & n928 ;
  assign n929 = n928 ^ n925 ;
  assign n931 = n535 & ~n612 ;
  assign n930 = n532 & n612 ;
  assign n932 = n931 ^ n930 ;
  assign n934 = n844 & ~n922 ;
  assign n933 = n847 & n922 ;
  assign n935 = n934 ^ n933 ;
  assign n1004 = n932 & ~n935 ;
  assign n1005 = ~n929 & n1004 ;
  assign n1007 = n1006 ^ n1005 ;
  assign n936 = n935 ^ n932 ;
  assign n937 = ~n929 & ~n936 ;
  assign n939 = n543 & ~n612 ;
  assign n938 = n540 & n612 ;
  assign n940 = n939 ^ n938 ;
  assign n942 = n852 & ~n922 ;
  assign n941 = n855 & n922 ;
  assign n943 = n942 ^ n941 ;
  assign n1001 = n940 & ~n943 ;
  assign n944 = n943 ^ n940 ;
  assign n946 = n550 & ~n612 ;
  assign n945 = n547 & n612 ;
  assign n947 = n946 ^ n945 ;
  assign n949 = n859 & ~n922 ;
  assign n948 = n862 & n922 ;
  assign n950 = n949 ^ n948 ;
  assign n999 = n947 & ~n950 ;
  assign n1000 = ~n944 & n999 ;
  assign n1002 = n1001 ^ n1000 ;
  assign n1003 = n937 & n1002 ;
  assign n1008 = n1007 ^ n1003 ;
  assign n951 = n950 ^ n947 ;
  assign n952 = ~n944 & ~n951 ;
  assign n953 = n937 & n952 ;
  assign n955 = n559 & ~n612 ;
  assign n954 = n556 & n612 ;
  assign n956 = n955 ^ n954 ;
  assign n958 = n868 & ~n922 ;
  assign n957 = n871 & n922 ;
  assign n959 = n958 ^ n957 ;
  assign n995 = n956 & ~n959 ;
  assign n960 = n959 ^ n956 ;
  assign n962 = n566 & ~n612 ;
  assign n961 = n563 & n612 ;
  assign n963 = n962 ^ n961 ;
  assign n965 = n875 & ~n922 ;
  assign n964 = n878 & n922 ;
  assign n966 = n965 ^ n964 ;
  assign n993 = n963 & ~n966 ;
  assign n994 = ~n960 & n993 ;
  assign n996 = n995 ^ n994 ;
  assign n967 = n966 ^ n963 ;
  assign n968 = ~n960 & ~n967 ;
  assign n970 = n574 & ~n612 ;
  assign n969 = n571 & n612 ;
  assign n971 = n970 ^ n969 ;
  assign n973 = n883 & ~n922 ;
  assign n972 = n886 & n922 ;
  assign n974 = n973 ^ n972 ;
  assign n990 = n971 & ~n974 ;
  assign n975 = n974 ^ n971 ;
  assign n976 = n668 ^ n583 ;
  assign n977 = n976 ^ n669 ;
  assign n979 = n889 & n922 ;
  assign n980 = n979 ^ n889 ;
  assign n978 = n893 & n922 ;
  assign n981 = n980 ^ n978 ;
  assign n986 = n977 & n981 ;
  assign n987 = n986 ^ n977 ;
  assign n988 = n975 & n987 ;
  assign n989 = n988 ^ n987 ;
  assign n991 = n990 ^ n989 ;
  assign n992 = n968 & n991 ;
  assign n997 = n996 ^ n992 ;
  assign n998 = n953 & n997 ;
  assign n1009 = n1008 ^ n998 ;
  assign n982 = n981 ^ n977 ;
  assign n983 = ~n975 & ~n982 ;
  assign n984 = n968 & n983 ;
  assign n985 = n953 & n984 ;
  assign n1010 = n1009 ^ n985 ;
  assign n1012 = n928 & n1010 ;
  assign n1013 = n1012 ^ n928 ;
  assign n1011 = n925 & n1010 ;
  assign n1014 = n1013 ^ n1011 ;
  assign n1016 = n932 & n1010 ;
  assign n1017 = n1016 ^ n932 ;
  assign n1015 = n935 & n1010 ;
  assign n1018 = n1017 ^ n1015 ;
  assign n1020 = n940 & n1010 ;
  assign n1021 = n1020 ^ n940 ;
  assign n1019 = n943 & n1010 ;
  assign n1022 = n1021 ^ n1019 ;
  assign n1024 = n947 & n1010 ;
  assign n1025 = n1024 ^ n947 ;
  assign n1023 = n950 & n1010 ;
  assign n1026 = n1025 ^ n1023 ;
  assign n1028 = n956 & n1010 ;
  assign n1029 = n1028 ^ n956 ;
  assign n1027 = n959 & n1010 ;
  assign n1030 = n1029 ^ n1027 ;
  assign n1032 = n963 & n1010 ;
  assign n1033 = n1032 ^ n963 ;
  assign n1031 = n966 & n1010 ;
  assign n1034 = n1033 ^ n1031 ;
  assign n1036 = n971 & n1010 ;
  assign n1037 = n1036 ^ n971 ;
  assign n1035 = n974 & n1010 ;
  assign n1038 = n1037 ^ n1035 ;
  assign n1040 = n977 & n1010 ;
  assign n1041 = n1040 ^ n977 ;
  assign n1039 = n981 & n1010 ;
  assign n1042 = n1041 ^ n1039 ;
  assign n1043 = n1011 ^ n925 ;
  assign n1044 = n1043 ^ n1012 ;
  assign n1045 = n1015 ^ n935 ;
  assign n1046 = n1045 ^ n1016 ;
  assign n1047 = n1019 ^ n943 ;
  assign n1048 = n1047 ^ n1020 ;
  assign n1049 = n1023 ^ n950 ;
  assign n1050 = n1049 ^ n1024 ;
  assign n1051 = n1027 ^ n959 ;
  assign n1052 = n1051 ^ n1028 ;
  assign n1053 = n1031 ^ n966 ;
  assign n1054 = n1053 ^ n1032 ;
  assign n1055 = n1035 ^ n974 ;
  assign n1056 = n1055 ^ n1036 ;
  assign n1057 = n1039 ^ n981 ;
  assign n1058 = n1057 ^ n1040 ;
  assign n1063 = n837 & ~n922 ;
  assign n1062 = n840 & n922 ;
  assign n1064 = n1063 ^ n1062 ;
  assign n1060 = n751 & ~n834 ;
  assign n1059 = n754 & n834 ;
  assign n1061 = n1060 ^ n1059 ;
  assign n1140 = ~n1061 & n1064 ;
  assign n1065 = n1064 ^ n1061 ;
  assign n1067 = n847 & ~n922 ;
  assign n1066 = n844 & n922 ;
  assign n1068 = n1067 ^ n1066 ;
  assign n1070 = n761 & ~n834 ;
  assign n1069 = n758 & n834 ;
  assign n1071 = n1070 ^ n1069 ;
  assign n1138 = n1068 & ~n1071 ;
  assign n1139 = ~n1065 & n1138 ;
  assign n1141 = n1140 ^ n1139 ;
  assign n1072 = n1071 ^ n1068 ;
  assign n1073 = ~n1065 & ~n1072 ;
  assign n1075 = n855 & ~n922 ;
  assign n1074 = n852 & n922 ;
  assign n1076 = n1075 ^ n1074 ;
  assign n1078 = n769 & ~n834 ;
  assign n1077 = n766 & n834 ;
  assign n1079 = n1078 ^ n1077 ;
  assign n1135 = n1076 & ~n1079 ;
  assign n1080 = n1079 ^ n1076 ;
  assign n1082 = n862 & ~n922 ;
  assign n1081 = n859 & n922 ;
  assign n1083 = n1082 ^ n1081 ;
  assign n1085 = n776 & ~n834 ;
  assign n1084 = n773 & n834 ;
  assign n1086 = n1085 ^ n1084 ;
  assign n1133 = n1083 & ~n1086 ;
  assign n1134 = ~n1080 & n1133 ;
  assign n1136 = n1135 ^ n1134 ;
  assign n1137 = n1073 & n1136 ;
  assign n1142 = n1141 ^ n1137 ;
  assign n1087 = n1086 ^ n1083 ;
  assign n1088 = ~n1080 & ~n1087 ;
  assign n1089 = n1073 & n1088 ;
  assign n1091 = n871 & ~n922 ;
  assign n1090 = n868 & n922 ;
  assign n1092 = n1091 ^ n1090 ;
  assign n1094 = n785 & ~n834 ;
  assign n1093 = n782 & n834 ;
  assign n1095 = n1094 ^ n1093 ;
  assign n1129 = n1092 & ~n1095 ;
  assign n1096 = n1095 ^ n1092 ;
  assign n1098 = n878 & ~n922 ;
  assign n1097 = n875 & n922 ;
  assign n1099 = n1098 ^ n1097 ;
  assign n1101 = n792 & ~n834 ;
  assign n1100 = n789 & n834 ;
  assign n1102 = n1101 ^ n1100 ;
  assign n1127 = n1099 & ~n1102 ;
  assign n1128 = ~n1096 & n1127 ;
  assign n1130 = n1129 ^ n1128 ;
  assign n1103 = n1102 ^ n1099 ;
  assign n1104 = ~n1096 & ~n1103 ;
  assign n1106 = n886 & ~n922 ;
  assign n1105 = n883 & n922 ;
  assign n1107 = n1106 ^ n1105 ;
  assign n1109 = n800 & ~n834 ;
  assign n1108 = n797 & n834 ;
  assign n1110 = n1109 ^ n1108 ;
  assign n1124 = n1107 & ~n1110 ;
  assign n1111 = n1110 ^ n1107 ;
  assign n1112 = n978 ^ n893 ;
  assign n1113 = n1112 ^ n979 ;
  assign n1114 = n805 & ~n834 ;
  assign n1115 = n1114 ^ n891 ;
  assign n1120 = n1113 & n1115 ;
  assign n1121 = n1120 ^ n1113 ;
  assign n1122 = n1111 & n1121 ;
  assign n1123 = n1122 ^ n1121 ;
  assign n1125 = n1124 ^ n1123 ;
  assign n1126 = n1104 & n1125 ;
  assign n1131 = n1130 ^ n1126 ;
  assign n1132 = n1089 & n1131 ;
  assign n1143 = n1142 ^ n1132 ;
  assign n1116 = n1115 ^ n1113 ;
  assign n1117 = ~n1111 & ~n1116 ;
  assign n1118 = n1104 & n1117 ;
  assign n1119 = n1089 & n1118 ;
  assign n1144 = n1143 ^ n1119 ;
  assign n1146 = n1064 & n1144 ;
  assign n1147 = n1146 ^ n1064 ;
  assign n1145 = n1061 & n1144 ;
  assign n1148 = n1147 ^ n1145 ;
  assign n1150 = n1068 & n1144 ;
  assign n1151 = n1150 ^ n1068 ;
  assign n1149 = n1071 & n1144 ;
  assign n1152 = n1151 ^ n1149 ;
  assign n1154 = n1076 & n1144 ;
  assign n1155 = n1154 ^ n1076 ;
  assign n1153 = n1079 & n1144 ;
  assign n1156 = n1155 ^ n1153 ;
  assign n1158 = n1083 & n1144 ;
  assign n1159 = n1158 ^ n1083 ;
  assign n1157 = n1086 & n1144 ;
  assign n1160 = n1159 ^ n1157 ;
  assign n1162 = n1092 & n1144 ;
  assign n1163 = n1162 ^ n1092 ;
  assign n1161 = n1095 & n1144 ;
  assign n1164 = n1163 ^ n1161 ;
  assign n1166 = n1099 & n1144 ;
  assign n1167 = n1166 ^ n1099 ;
  assign n1165 = n1102 & n1144 ;
  assign n1168 = n1167 ^ n1165 ;
  assign n1170 = n1107 & n1144 ;
  assign n1171 = n1170 ^ n1107 ;
  assign n1169 = n1110 & n1144 ;
  assign n1172 = n1171 ^ n1169 ;
  assign n1174 = n1113 & n1144 ;
  assign n1175 = n1174 ^ n1113 ;
  assign n1173 = n1115 & n1144 ;
  assign n1176 = n1175 ^ n1173 ;
  assign n1177 = n1145 ^ n1061 ;
  assign n1178 = n1177 ^ n1146 ;
  assign n1179 = n1149 ^ n1071 ;
  assign n1180 = n1179 ^ n1150 ;
  assign n1181 = n1153 ^ n1079 ;
  assign n1182 = n1181 ^ n1154 ;
  assign n1183 = n1157 ^ n1086 ;
  assign n1184 = n1183 ^ n1158 ;
  assign n1185 = n1161 ^ n1095 ;
  assign n1186 = n1185 ^ n1162 ;
  assign n1187 = n1165 ^ n1102 ;
  assign n1188 = n1187 ^ n1166 ;
  assign n1189 = n1169 ^ n1110 ;
  assign n1190 = n1189 ^ n1170 ;
  assign n1191 = n1173 ^ n1115 ;
  assign n1192 = n1191 ^ n1174 ;
  assign y0 = n704 ;
  assign y1 = n708 ;
  assign y2 = n712 ;
  assign y3 = n716 ;
  assign y4 = n720 ;
  assign y5 = n724 ;
  assign y6 = n728 ;
  assign y7 = n732 ;
  assign y8 = n734 ;
  assign y9 = n736 ;
  assign y10 = n738 ;
  assign y11 = n740 ;
  assign y12 = n742 ;
  assign y13 = n744 ;
  assign y14 = n746 ;
  assign y15 = n748 ;
  assign y16 = n1014 ;
  assign y17 = n1018 ;
  assign y18 = n1022 ;
  assign y19 = n1026 ;
  assign y20 = n1030 ;
  assign y21 = n1034 ;
  assign y22 = n1038 ;
  assign y23 = n1042 ;
  assign y24 = n1044 ;
  assign y25 = n1046 ;
  assign y26 = n1048 ;
  assign y27 = n1050 ;
  assign y28 = n1052 ;
  assign y29 = n1054 ;
  assign y30 = n1056 ;
  assign y31 = n1058 ;
  assign y32 = n1148 ;
  assign y33 = n1152 ;
  assign y34 = n1156 ;
  assign y35 = n1160 ;
  assign y36 = n1164 ;
  assign y37 = n1168 ;
  assign y38 = n1172 ;
  assign y39 = n1176 ;
  assign y40 = n1178 ;
  assign y41 = n1180 ;
  assign y42 = n1182 ;
  assign y43 = n1184 ;
  assign y44 = n1186 ;
  assign y45 = n1188 ;
  assign y46 = n1190 ;
  assign y47 = n1192 ;
endmodule
