module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 ;
  assign n27 = x10 ^ x2 ;
  assign n28 = ~x3 & ~x11 ;
  assign n32 = ~n27 & n28 ;
  assign n17 = x5 & x13 ;
  assign n18 = x6 & x14 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = ~x5 & ~x13 ;
  assign n21 = ~x4 & ~x12 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = ~n19 & n22 ;
  assign n24 = x3 & x11 ;
  assign n25 = x4 & x12 ;
  assign n26 = ~n24 & ~n25 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = n26 & n29 ;
  assign n31 = ~n23 & n30 ;
  assign n33 = n32 ^ n31 ;
  assign n39 = x1 & x9 ;
  assign n40 = ~x8 & n39 ;
  assign n47 = ~n33 & n40 ;
  assign n34 = x14 ^ x6 ;
  assign n35 = x7 & x15 ;
  assign n36 = n34 & n35 ;
  assign n37 = x13 ^ x5 ;
  assign n38 = n36 & n37 ;
  assign n41 = x12 ^ x4 ;
  assign n42 = x11 ^ x3 ;
  assign n43 = n41 & n42 ;
  assign n44 = ~n40 & n43 ;
  assign n45 = n38 & n44 ;
  assign n46 = ~n33 & n45 ;
  assign n48 = n47 ^ n46 ;
  assign n50 = x9 ^ x1 ;
  assign n51 = x2 & x10 ;
  assign n52 = ~n50 & ~n51 ;
  assign n59 = n48 & ~n52 ;
  assign n49 = n38 & n43 ;
  assign n53 = x0 & x8 ;
  assign n54 = ~n39 & n53 ;
  assign n55 = ~n40 & ~n54 ;
  assign n56 = ~n52 & ~n55 ;
  assign n57 = n49 & n56 ;
  assign n58 = n48 & n57 ;
  assign n60 = n59 ^ n58 ;
  assign n61 = ~x2 & ~x10 ;
  assign n62 = ~n28 & ~n61 ;
  assign n63 = n26 & n62 ;
  assign n64 = ~n23 & n63 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = ~x0 & ~x8 ;
  assign n67 = ~n39 & ~n51 ;
  assign n68 = ~n66 & n67 ;
  assign n69 = ~n65 & n68 ;
  assign n70 = x2 & ~n28 ;
  assign n71 = n26 & n70 ;
  assign n72 = ~n23 & n71 ;
  assign n73 = n72 ^ n70 ;
  assign n74 = ~x0 & x10 ;
  assign n75 = n40 & n74 ;
  assign n76 = ~x1 & ~x9 ;
  assign n77 = ~n53 & ~n76 ;
  assign n78 = ~n66 & ~n77 ;
  assign n79 = n75 & ~n78 ;
  assign n80 = n73 & n79 ;
  assign n81 = n80 ^ n78 ;
  assign n82 = ~n69 & ~n81 ;
  assign n83 = ~n60 & ~n82 ;
  assign n84 = n73 ^ n50 ;
  assign n85 = n26 & ~n28 ;
  assign n86 = ~n23 & n85 ;
  assign n87 = n86 ^ n28 ;
  assign n88 = n87 ^ n27 ;
  assign n89 = n84 & ~n88 ;
  assign n90 = x8 ^ x0 ;
  assign n91 = n90 ^ n39 ;
  assign n92 = n91 ^ n49 ;
  assign n93 = n89 & ~n92 ;
  assign n94 = n50 & n61 ;
  assign n95 = ~n76 & ~n94 ;
  assign n96 = n95 ^ n90 ;
  assign n97 = ~n89 & ~n96 ;
  assign n98 = ~n93 & ~n97 ;
  assign n102 = ~n84 & ~n88 ;
  assign n101 = ~n49 & ~n88 ;
  assign n103 = n102 ^ n101 ;
  assign n99 = n61 ^ n50 ;
  assign n100 = n88 & ~n99 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = n88 ^ n49 ;
  assign n106 = n19 & ~n36 ;
  assign n107 = ~n20 & ~n106 ;
  assign n108 = ~n25 & ~n107 ;
  assign n109 = ~n21 & ~n108 ;
  assign n110 = n109 ^ n42 ;
  assign n111 = ~n18 & ~n38 ;
  assign n112 = n37 & ~n111 ;
  assign n113 = ~n17 & ~n112 ;
  assign n114 = n113 ^ n41 ;
  assign n115 = ~n18 & ~n36 ;
  assign n116 = n115 ^ n37 ;
  assign n117 = n35 ^ n34 ;
  assign y0 = n83 ;
  assign y1 = n98 ;
  assign y2 = n104 ;
  assign y3 = ~n105 ;
  assign y4 = n110 ;
  assign y5 = ~n114 ;
  assign y6 = ~n116 ;
  assign y7 = n117 ;
endmodule
