module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 ;
  assign n148 = ~x5 & ~x22 ;
  assign n191 = ~x56 & ~n148 ;
  assign n149 = ~x9 & ~x11 ;
  assign n213 = n191 ^ n149 ;
  assign n150 = ~x56 & ~n149 ;
  assign n151 = n148 & n150 ;
  assign n201 = n151 ^ x54 ;
  assign n214 = n213 ^ n201 ;
  assign n152 = n151 ^ n149 ;
  assign n192 = n191 ^ n151 ;
  assign n193 = ~n152 & n192 ;
  assign n194 = n193 ^ n191 ;
  assign n168 = x14 ^ x10 ;
  assign n169 = n168 ^ x14 ;
  assign n156 = x21 ^ x7 ;
  assign n155 = x21 ^ x8 ;
  assign n157 = n156 ^ n155 ;
  assign n154 = x21 ^ x13 ;
  assign n158 = n157 ^ n154 ;
  assign n159 = n155 ^ x21 ;
  assign n160 = n159 ^ x21 ;
  assign n161 = n154 ^ x21 ;
  assign n162 = n161 ^ n159 ;
  assign n163 = n160 & n162 ;
  assign n164 = n163 ^ n159 ;
  assign n165 = n158 & n164 ;
  assign n166 = n165 ^ n158 ;
  assign n170 = n169 ^ n166 ;
  assign n167 = n166 ^ x14 ;
  assign n171 = n170 ^ n167 ;
  assign n177 = n158 & ~n169 ;
  assign n178 = ~n164 & n177 ;
  assign n172 = ~x7 & ~x13 ;
  assign n173 = x8 & x21 ;
  assign n174 = n173 ^ x8 ;
  assign n175 = n174 ^ x21 ;
  assign n176 = n172 & ~n175 ;
  assign n179 = n178 ^ n176 ;
  assign n180 = n171 & n179 ;
  assign n181 = n180 ^ n178 ;
  assign n182 = ~x4 & ~x19 ;
  assign n183 = ~x16 & ~x18 ;
  assign n184 = n182 & n183 ;
  assign n185 = ~x6 & ~x12 ;
  assign n186 = ~x17 & n185 ;
  assign n187 = n148 & n186 ;
  assign n188 = n184 & n187 ;
  assign n189 = ~n181 & n188 ;
  assign n190 = n189 ^ n188 ;
  assign n195 = n194 ^ n190 ;
  assign n200 = n194 ^ n149 ;
  assign n202 = n201 ^ n200 ;
  assign n203 = n195 & n202 ;
  assign n211 = n203 ^ n193 ;
  assign n153 = n152 ^ x54 ;
  assign n196 = n195 ^ n153 ;
  assign n197 = n190 ^ n149 ;
  assign n198 = n197 ^ n194 ;
  assign n199 = ~n196 & n198 ;
  assign n204 = n203 ^ n199 ;
  assign n205 = n204 ^ n194 ;
  assign n206 = n205 ^ n153 ;
  assign n207 = n203 ^ n190 ;
  assign n208 = n207 ^ x54 ;
  assign n209 = n206 & ~n208 ;
  assign n210 = n209 ^ n199 ;
  assign n212 = n211 ^ n210 ;
  assign n215 = n214 ^ n212 ;
  assign n216 = n215 ^ x54 ;
  assign n218 = ~x14 & ~x22 ;
  assign n219 = n172 & n218 ;
  assign n220 = n149 & n219 ;
  assign n221 = ~x17 & ~x21 ;
  assign n222 = ~x8 & n221 ;
  assign n223 = ~x5 & n185 ;
  assign n224 = n222 & n223 ;
  assign n225 = n220 & n224 ;
  assign n226 = ~x0 & x54 ;
  assign n227 = n184 & n226 ;
  assign n228 = n225 & n227 ;
  assign n217 = ~x0 & ~x54 ;
  assign n229 = n228 ^ n217 ;
  assign n230 = ~x3 & ~x129 ;
  assign n231 = ~n229 & n230 ;
  assign n232 = ~n216 & n231 ;
  assign n233 = n232 ^ n230 ;
  assign n234 = ~x5 & ~x6 ;
  assign n235 = ~x7 & ~x12 ;
  assign n236 = ~n234 & ~n235 ;
  assign n237 = ~x13 & ~n236 ;
  assign n238 = ~x5 & ~x7 ;
  assign n239 = n238 ^ n185 ;
  assign n240 = n237 & n239 ;
  assign n241 = x13 & n185 ;
  assign n242 = n238 & n241 ;
  assign n243 = ~x9 & ~n242 ;
  assign n244 = ~n240 & n243 ;
  assign n245 = n172 & n223 ;
  assign n246 = x9 & ~n245 ;
  assign n247 = ~x10 & x54 ;
  assign n248 = n218 & n247 ;
  assign n249 = ~x8 & ~x11 ;
  assign n250 = n221 & n249 ;
  assign n251 = n248 & n250 ;
  assign n252 = n184 & n251 ;
  assign n253 = ~n246 & n252 ;
  assign n254 = ~n244 & n253 ;
  assign n255 = n172 & n234 ;
  assign n256 = n184 & n255 ;
  assign n257 = ~x14 & ~n175 ;
  assign n258 = ~x11 & ~x12 ;
  assign n259 = ~x10 & ~x22 ;
  assign n260 = n258 & n259 ;
  assign n261 = n257 & n260 ;
  assign n262 = n256 & n261 ;
  assign n263 = ~x17 & x54 ;
  assign n264 = ~x1 & n263 ;
  assign n265 = ~n262 & n264 ;
  assign n266 = n265 ^ x1 ;
  assign n267 = n230 & n266 ;
  assign n268 = ~n254 & n267 ;
  assign n269 = n268 ^ n230 ;
  assign n270 = ~x38 & ~x50 ;
  assign n271 = ~x40 & ~x46 ;
  assign n272 = n270 & n271 ;
  assign n273 = ~x41 & ~x43 ;
  assign n274 = ~x42 & ~x44 ;
  assign n275 = n273 & n274 ;
  assign n276 = n272 & n275 ;
  assign n277 = ~x47 & ~x48 ;
  assign n278 = n276 & n277 ;
  assign n279 = ~x15 & ~x20 ;
  assign n280 = ~x45 & n279 ;
  assign n281 = ~x24 & ~x49 ;
  assign n282 = x82 & n281 ;
  assign n283 = n280 & n282 ;
  assign n284 = x122 & x127 ;
  assign n285 = ~x82 & ~n284 ;
  assign n286 = x2 & ~n285 ;
  assign n287 = n283 & n286 ;
  assign n288 = n278 & n287 ;
  assign n289 = n288 ^ n286 ;
  assign n299 = ~x65 & ~n284 ;
  assign n304 = ~x82 & n299 ;
  assign n305 = ~n289 & n304 ;
  assign n306 = n305 ^ n289 ;
  assign n290 = n280 & n281 ;
  assign n291 = ~x41 & ~x46 ;
  assign n292 = n270 & n291 ;
  assign n293 = ~x43 & ~x47 ;
  assign n294 = ~x2 & ~x48 ;
  assign n295 = n293 & n294 ;
  assign n296 = n292 & n295 ;
  assign n297 = n290 & n296 ;
  assign n298 = ~x40 & n274 ;
  assign n300 = x82 & n299 ;
  assign n301 = n298 & n300 ;
  assign n302 = n297 & n301 ;
  assign n303 = ~n289 & n302 ;
  assign n307 = n306 ^ n303 ;
  assign n308 = ~x129 & n307 ;
  assign n309 = x0 & ~x113 ;
  assign n310 = ~x123 & n309 ;
  assign n311 = ~x9 & ~x14 ;
  assign n312 = n259 & n311 ;
  assign n313 = ~x12 & n250 ;
  assign n314 = n312 & n313 ;
  assign n315 = n256 & n314 ;
  assign n316 = ~x61 & ~x118 ;
  assign n317 = ~n315 & n316 ;
  assign n318 = ~n310 & ~n317 ;
  assign n319 = ~x129 & ~n318 ;
  assign n320 = x4 & ~x54 ;
  assign n321 = n245 & n311 ;
  assign n322 = ~x18 & n182 ;
  assign n323 = ~x16 & x54 ;
  assign n324 = n221 & n323 ;
  assign n325 = n322 & n324 ;
  assign n326 = n249 & n325 ;
  assign n327 = x10 & ~x22 ;
  assign n328 = n326 & n327 ;
  assign n329 = n321 & n328 ;
  assign n330 = ~n320 & ~n329 ;
  assign n331 = n230 & ~n330 ;
  assign n332 = x5 & ~x54 ;
  assign n333 = ~x13 & n312 ;
  assign n334 = ~x59 & n250 ;
  assign n335 = n333 & n334 ;
  assign n336 = n185 & n238 ;
  assign n337 = n323 & n336 ;
  assign n338 = ~x25 & x28 ;
  assign n339 = ~x29 & n338 ;
  assign n340 = n322 & n339 ;
  assign n341 = n337 & n340 ;
  assign n342 = n335 & n341 ;
  assign n343 = ~n332 & ~n342 ;
  assign n344 = n230 & ~n343 ;
  assign n345 = x6 & ~x54 ;
  assign n346 = ~x28 & ~x29 ;
  assign n347 = x25 & n346 ;
  assign n348 = n322 & n347 ;
  assign n349 = n337 & n348 ;
  assign n350 = n335 & n349 ;
  assign n351 = ~n345 & ~n350 ;
  assign n352 = n230 & ~n351 ;
  assign n353 = x7 & ~x54 ;
  assign n354 = x8 & n325 ;
  assign n355 = ~x11 & n336 ;
  assign n356 = n333 & n355 ;
  assign n357 = n354 & n356 ;
  assign n358 = ~n353 & ~n357 ;
  assign n359 = n230 & ~n358 ;
  assign n360 = x8 & ~x54 ;
  assign n361 = ~x12 & n312 ;
  assign n362 = n255 & n361 ;
  assign n363 = n182 & n323 ;
  assign n364 = ~x17 & ~x18 ;
  assign n365 = n249 & n364 ;
  assign n366 = x21 & n365 ;
  assign n367 = n363 & n366 ;
  assign n368 = n362 & n367 ;
  assign n369 = ~n360 & ~n368 ;
  assign n370 = n230 & ~n369 ;
  assign n371 = x9 & ~x54 ;
  assign n372 = ~x8 & n325 ;
  assign n373 = x11 & n336 ;
  assign n374 = n333 & n373 ;
  assign n375 = n372 & n374 ;
  assign n376 = ~n371 & ~n375 ;
  assign n377 = n230 & ~n376 ;
  assign n378 = x10 & ~x54 ;
  assign n379 = ~x9 & ~x18 ;
  assign n380 = n222 & n379 ;
  assign n381 = n259 & n380 ;
  assign n382 = ~x13 & x14 ;
  assign n383 = n363 & n382 ;
  assign n384 = n355 & n383 ;
  assign n385 = n381 & n384 ;
  assign n386 = ~n378 & ~n385 ;
  assign n387 = n230 & ~n386 ;
  assign n388 = x11 & ~x54 ;
  assign n389 = ~x10 & ~x11 ;
  assign n390 = x22 & n389 ;
  assign n391 = n321 & n390 ;
  assign n392 = n372 & n391 ;
  assign n393 = ~n388 & ~n392 ;
  assign n394 = n230 & ~n393 ;
  assign n395 = x12 & ~x54 ;
  assign n396 = x18 & n255 ;
  assign n397 = n312 & n363 ;
  assign n398 = n396 & n397 ;
  assign n399 = n313 & n398 ;
  assign n400 = ~n395 & ~n399 ;
  assign n401 = n230 & ~n400 ;
  assign n402 = x13 & ~x54 ;
  assign n403 = ~x25 & ~x28 ;
  assign n404 = x29 & n403 ;
  assign n405 = ~x59 & n259 ;
  assign n406 = n404 & n405 ;
  assign n407 = n326 & n406 ;
  assign n408 = n321 & n407 ;
  assign n409 = ~n402 & ~n408 ;
  assign n410 = n230 & ~n409 ;
  assign n411 = x14 & ~x54 ;
  assign n412 = x13 & ~x16 ;
  assign n413 = n182 & n412 ;
  assign n414 = n248 & n413 ;
  assign n415 = n355 & n414 ;
  assign n416 = n380 & n415 ;
  assign n417 = ~n411 & ~n416 ;
  assign n418 = n230 & ~n417 ;
  assign n432 = n277 & n281 ;
  assign n433 = ~x15 & ~x45 ;
  assign n434 = n273 & n433 ;
  assign n435 = n432 & n434 ;
  assign n436 = x82 & n274 ;
  assign n437 = n272 & n436 ;
  assign n438 = n435 & n437 ;
  assign n439 = n438 ^ x82 ;
  assign n440 = ~x82 & n284 ;
  assign n441 = x15 & n440 ;
  assign n442 = ~x70 & ~n284 ;
  assign n443 = ~n441 & n442 ;
  assign n444 = ~n439 & n443 ;
  assign n445 = n444 ^ n441 ;
  assign n449 = ~x129 & n445 ;
  assign n419 = n292 & n298 ;
  assign n420 = ~x45 & n281 ;
  assign n421 = ~x48 & n293 ;
  assign n422 = n420 & n421 ;
  assign n423 = n419 & n422 ;
  assign n424 = x15 & ~n423 ;
  assign n425 = ~x15 & n281 ;
  assign n426 = ~x45 & n277 ;
  assign n427 = ~x2 & ~x20 ;
  assign n428 = n426 & ~n427 ;
  assign n429 = n425 & n428 ;
  assign n430 = n276 & n429 ;
  assign n431 = ~n424 & ~n430 ;
  assign n446 = x82 & ~x129 ;
  assign n447 = ~n445 & n446 ;
  assign n448 = ~n431 & n447 ;
  assign n450 = n449 ^ n448 ;
  assign n451 = x16 & ~x54 ;
  assign n452 = x6 & ~x13 ;
  assign n453 = n238 & n452 ;
  assign n454 = n361 & n453 ;
  assign n455 = n326 & n454 ;
  assign n456 = ~n451 & ~n455 ;
  assign n457 = n230 & ~n456 ;
  assign n458 = x17 & ~x54 ;
  assign n459 = ~x25 & x59 ;
  assign n460 = ~n175 & n459 ;
  assign n461 = n263 & n346 ;
  assign n462 = n460 & n461 ;
  assign n463 = n184 & n462 ;
  assign n464 = n356 & n463 ;
  assign n465 = ~n458 & ~n464 ;
  assign n466 = n230 & ~n465 ;
  assign n467 = x18 & ~x54 ;
  assign n468 = n322 & n362 ;
  assign n469 = x16 & x54 ;
  assign n470 = n250 & n469 ;
  assign n471 = n468 & n470 ;
  assign n472 = ~n467 & ~n471 ;
  assign n473 = n230 & ~n472 ;
  assign n474 = x19 & ~x54 ;
  assign n475 = x17 & ~x21 ;
  assign n476 = n249 & n475 ;
  assign n477 = n323 & n476 ;
  assign n478 = n468 & n477 ;
  assign n479 = ~n474 & ~n478 ;
  assign n480 = n230 & ~n479 ;
  assign n482 = ~x46 & ~x50 ;
  assign n483 = ~x38 & ~x40 ;
  assign n484 = n274 & n483 ;
  assign n485 = n482 & n484 ;
  assign n486 = n273 & n281 ;
  assign n487 = n426 & n486 ;
  assign n488 = n485 & n487 ;
  assign n491 = ~x2 & ~x15 ;
  assign n492 = ~x20 & x82 ;
  assign n493 = n491 & n492 ;
  assign n494 = n488 & n493 ;
  assign n489 = ~x15 & x82 ;
  assign n490 = n488 & n489 ;
  assign n495 = n494 ^ n490 ;
  assign n481 = x20 & x82 ;
  assign n496 = n495 ^ n481 ;
  assign n497 = x20 & n440 ;
  assign n498 = ~x71 & ~n284 ;
  assign n503 = ~x82 & n498 ;
  assign n504 = ~n497 & n503 ;
  assign n505 = n504 ^ n497 ;
  assign n499 = x82 & n279 ;
  assign n500 = n498 & n499 ;
  assign n501 = ~n497 & n500 ;
  assign n502 = n488 & n501 ;
  assign n506 = n505 ^ n502 ;
  assign n507 = ~n496 & ~n506 ;
  assign n508 = ~x129 & ~n507 ;
  assign n509 = x21 & ~x54 ;
  assign n510 = ~x4 & x19 ;
  assign n511 = ~x21 & n510 ;
  assign n512 = n323 & n511 ;
  assign n513 = n365 & n512 ;
  assign n514 = n362 & n513 ;
  assign n515 = ~n509 & ~n514 ;
  assign n516 = n230 & ~n515 ;
  assign n517 = x22 & ~x54 ;
  assign n518 = x5 & ~x6 ;
  assign n519 = ~x14 & n518 ;
  assign n520 = n172 & n258 ;
  assign n521 = n519 & n520 ;
  assign n522 = n363 & n521 ;
  assign n523 = n381 & n522 ;
  assign n524 = ~n517 & ~n523 ;
  assign n525 = n230 & ~n524 ;
  assign n526 = ~x23 & x55 ;
  assign n527 = x61 & ~x129 ;
  assign n528 = ~n526 & n527 ;
  assign n534 = ~x2 & n279 ;
  assign n544 = ~x49 & n534 ;
  assign n545 = x82 & ~n544 ;
  assign n546 = n284 & ~n545 ;
  assign n529 = n273 & n426 ;
  assign n547 = n272 & n274 ;
  assign n548 = n529 & n547 ;
  assign n549 = x82 & ~n548 ;
  assign n550 = ~n546 & ~n549 ;
  assign n530 = n485 & n529 ;
  assign n531 = x24 & x82 ;
  assign n532 = n530 & n531 ;
  assign n533 = ~x129 & ~n532 ;
  assign n535 = ~x45 & ~x49 ;
  assign n536 = n277 & n535 ;
  assign n537 = n534 & n536 ;
  assign n538 = n276 & n537 ;
  assign n539 = x63 & ~n284 ;
  assign n540 = x82 & n539 ;
  assign n541 = ~n538 & n540 ;
  assign n542 = n541 ^ n539 ;
  assign n551 = ~x24 & ~n542 ;
  assign n552 = n533 & n551 ;
  assign n553 = ~n550 & n552 ;
  assign n543 = n533 & ~n542 ;
  assign n554 = n553 ^ n543 ;
  assign n587 = ~x39 & ~x52 ;
  assign n588 = ~x51 & x116 ;
  assign n589 = n587 & n588 ;
  assign n590 = ~x85 & ~n589 ;
  assign n591 = ~x25 & ~x116 ;
  assign n592 = x26 & ~x27 ;
  assign n593 = ~n591 & n592 ;
  assign n594 = n590 & n593 ;
  assign n578 = ~x85 & ~x96 ;
  assign n579 = x100 & ~x110 ;
  assign n580 = n578 & n579 ;
  assign n576 = x85 & x100 ;
  assign n577 = x116 & n576 ;
  assign n581 = n580 ^ n577 ;
  assign n582 = x85 & ~x116 ;
  assign n583 = x25 & n582 ;
  assign n584 = ~n581 & ~n583 ;
  assign n585 = ~x26 & ~x27 ;
  assign n586 = ~n584 & n585 ;
  assign n595 = n594 ^ n586 ;
  assign n564 = ~x51 & ~x52 ;
  assign n565 = ~x39 & n564 ;
  assign n566 = x27 & ~n565 ;
  assign n567 = ~x95 & ~x100 ;
  assign n568 = ~x97 & ~x110 ;
  assign n569 = n567 & n568 ;
  assign n570 = n569 ^ x110 ;
  assign n571 = x25 & n570 ;
  assign n572 = ~n566 & n571 ;
  assign n573 = ~x26 & ~x85 ;
  assign n599 = n572 & n573 ;
  assign n600 = ~n595 & n599 ;
  assign n601 = n600 ^ n595 ;
  assign n574 = x27 & n573 ;
  assign n575 = ~n572 & n574 ;
  assign n557 = x25 & ~x116 ;
  assign n596 = ~n557 & ~n589 ;
  assign n597 = ~n595 & ~n596 ;
  assign n598 = n575 & n597 ;
  assign n602 = n601 ^ n598 ;
  assign n555 = ~x53 & ~x58 ;
  assign n556 = ~x27 & ~x85 ;
  assign n558 = ~x26 & n557 ;
  assign n559 = n556 & n558 ;
  assign n560 = ~n555 & ~n559 ;
  assign n561 = n230 & ~n560 ;
  assign n562 = x58 ^ x53 ;
  assign n603 = ~x53 & ~n562 ;
  assign n604 = n561 & n603 ;
  assign n605 = n602 & n604 ;
  assign n563 = n561 & n562 ;
  assign n606 = n605 ^ n563 ;
  assign n607 = x26 & ~x85 ;
  assign n608 = ~n589 & n607 ;
  assign n609 = x26 & x116 ;
  assign n610 = n581 & ~n609 ;
  assign n611 = ~n608 & ~n610 ;
  assign n612 = ~x27 & ~x53 ;
  assign n613 = ~x58 & n612 ;
  assign n614 = n230 & n613 ;
  assign n615 = ~n611 & n614 ;
  assign n616 = x27 & n590 ;
  assign n617 = x85 & x116 ;
  assign n618 = ~x85 & ~x110 ;
  assign n619 = x95 & ~x96 ;
  assign n620 = n618 & n619 ;
  assign n621 = ~n617 & ~n620 ;
  assign n622 = ~x27 & ~x100 ;
  assign n623 = ~n621 & n622 ;
  assign n624 = ~n616 & ~n623 ;
  assign n625 = ~x26 & n230 ;
  assign n626 = n555 & n625 ;
  assign n627 = ~n624 & n626 ;
  assign n668 = ~x26 & ~x53 ;
  assign n669 = ~x85 & n668 ;
  assign n670 = ~x27 & x28 ;
  assign n671 = ~x116 & n670 ;
  assign n672 = x58 & n671 ;
  assign n673 = n669 & n672 ;
  assign n680 = x58 & n230 ;
  assign n681 = ~n673 & n680 ;
  assign n682 = n681 ^ n230 ;
  assign n628 = ~x51 & n587 ;
  assign n629 = n609 & n628 ;
  assign n635 = n556 & n629 ;
  assign n636 = n635 ^ x85 ;
  assign n630 = ~x26 & ~x100 ;
  assign n631 = ~x110 & n630 ;
  assign n632 = n556 & n619 ;
  assign n633 = n631 & n632 ;
  assign n634 = ~n629 & n633 ;
  assign n637 = n636 ^ n634 ;
  assign n638 = ~x26 & x116 ;
  assign n639 = n566 & n638 ;
  assign n640 = ~n637 & n639 ;
  assign n641 = n640 ^ n637 ;
  assign n644 = ~x27 & ~x39 ;
  assign n645 = n564 & n644 ;
  assign n646 = n645 ^ x26 ;
  assign n642 = ~x26 & ~x39 ;
  assign n643 = n564 & n642 ;
  assign n647 = n646 ^ n643 ;
  assign n648 = n570 & ~n647 ;
  assign n649 = x27 ^ x26 ;
  assign n650 = ~x116 & n649 ;
  assign n651 = x28 & ~n650 ;
  assign n652 = ~n648 & n651 ;
  assign n653 = n652 ^ x28 ;
  assign n654 = x100 & x116 ;
  assign n655 = ~x28 & ~x116 ;
  assign n656 = n585 & ~n655 ;
  assign n657 = ~n654 & n656 ;
  assign n663 = ~x53 & n657 ;
  assign n664 = ~n653 & n663 ;
  assign n665 = ~n641 & n664 ;
  assign n666 = n665 ^ n663 ;
  assign n658 = ~x53 & ~x85 ;
  assign n659 = ~n657 & n658 ;
  assign n660 = ~n653 & n659 ;
  assign n661 = ~n641 & n660 ;
  assign n662 = n661 ^ n659 ;
  assign n667 = n666 ^ n662 ;
  assign n674 = ~x58 & n230 ;
  assign n675 = x53 & n573 ;
  assign n676 = n671 & n675 ;
  assign n677 = n674 & ~n676 ;
  assign n678 = ~n673 & n677 ;
  assign n679 = ~n667 & n678 ;
  assign n683 = n682 ^ n679 ;
  assign n684 = x29 & ~x116 ;
  assign n685 = ~x85 & n555 ;
  assign n686 = n592 & n685 ;
  assign n687 = n684 & n686 ;
  assign n777 = n687 ^ x26 ;
  assign n755 = x129 ^ x3 ;
  assign n778 = n777 ^ n755 ;
  assign n694 = x27 & n555 ;
  assign n695 = n684 & n694 ;
  assign n749 = n695 ^ x27 ;
  assign n692 = x85 & n684 ;
  assign n693 = n613 & n692 ;
  assign n737 = n693 ^ x85 ;
  assign n750 = n749 ^ n737 ;
  assign n696 = n695 ^ n693 ;
  assign n728 = n693 ^ x27 ;
  assign n729 = n696 & n728 ;
  assign n730 = n729 ^ x27 ;
  assign n700 = x96 & x110 ;
  assign n701 = n700 ^ x96 ;
  assign n702 = n701 ^ x110 ;
  assign n703 = x97 & ~n702 ;
  assign n704 = n703 ^ x97 ;
  assign n705 = x29 & ~x110 ;
  assign n706 = n567 & n705 ;
  assign n707 = ~n704 & n706 ;
  assign n708 = n707 ^ n705 ;
  assign n709 = n708 ^ x29 ;
  assign n710 = ~x58 & x97 ;
  assign n711 = n567 & ~n702 ;
  assign n712 = n710 & n711 ;
  assign n713 = n712 ^ x58 ;
  assign n714 = n709 & ~n713 ;
  assign n715 = n714 ^ n713 ;
  assign n719 = ~x29 & ~x53 ;
  assign n720 = x58 & ~x116 ;
  assign n721 = n719 & n720 ;
  assign n722 = n721 ^ x53 ;
  assign n716 = ~x53 & x58 ;
  assign n717 = ~x97 & x116 ;
  assign n718 = n716 & n717 ;
  assign n723 = n722 ^ n718 ;
  assign n724 = n723 ^ n715 ;
  assign n725 = n715 & ~n724 ;
  assign n698 = x53 & ~x58 ;
  assign n699 = n684 & n698 ;
  assign n726 = n725 ^ n699 ;
  assign n727 = n726 ^ n715 ;
  assign n731 = n730 ^ n727 ;
  assign n736 = n730 ^ n695 ;
  assign n738 = n737 ^ n736 ;
  assign n739 = ~n731 & n738 ;
  assign n747 = n739 ^ n729 ;
  assign n697 = n696 ^ x85 ;
  assign n732 = n731 ^ n697 ;
  assign n733 = n727 ^ n695 ;
  assign n734 = n733 ^ n730 ;
  assign n735 = n732 & n734 ;
  assign n740 = n739 ^ n735 ;
  assign n741 = n740 ^ n730 ;
  assign n742 = n741 ^ n697 ;
  assign n743 = n739 ^ n727 ;
  assign n744 = n743 ^ x85 ;
  assign n745 = n742 & ~n744 ;
  assign n746 = n745 ^ n735 ;
  assign n748 = n747 ^ n746 ;
  assign n751 = n750 ^ n748 ;
  assign n752 = n751 ^ n693 ;
  assign n768 = x3 & ~x26 ;
  assign n769 = ~x129 & n768 ;
  assign n770 = ~n687 & n769 ;
  assign n771 = n752 & n770 ;
  assign n766 = x3 & x129 ;
  assign n767 = n687 & n766 ;
  assign n772 = n771 ^ n767 ;
  assign n763 = x26 & x129 ;
  assign n764 = n687 & n763 ;
  assign n765 = ~n752 & n764 ;
  assign n773 = n772 ^ n765 ;
  assign n688 = n687 ^ x129 ;
  assign n758 = n688 ^ x3 ;
  assign n689 = x129 ^ x26 ;
  assign n690 = n688 & n689 ;
  assign n691 = n690 ^ x26 ;
  assign n753 = n752 ^ n691 ;
  assign n759 = n758 ^ n753 ;
  assign n760 = n752 ^ n687 ;
  assign n761 = n760 ^ n691 ;
  assign n762 = n759 & n761 ;
  assign n774 = n773 ^ n762 ;
  assign n754 = n691 ^ n687 ;
  assign n756 = n755 ^ n754 ;
  assign n757 = ~n753 & n756 ;
  assign n775 = n774 ^ n757 ;
  assign n776 = n775 ^ n690 ;
  assign n779 = n778 ^ n776 ;
  assign n780 = ~x30 & ~x109 ;
  assign n781 = ~x60 & x109 ;
  assign n782 = ~n780 & ~n781 ;
  assign n783 = ~x106 & ~n782 ;
  assign n784 = ~x88 & x106 ;
  assign n785 = ~x129 & ~n784 ;
  assign n786 = ~n783 & n785 ;
  assign n787 = ~x31 & ~x109 ;
  assign n788 = ~x30 & x109 ;
  assign n789 = ~n787 & ~n788 ;
  assign n790 = ~x106 & ~n789 ;
  assign n791 = ~x89 & x106 ;
  assign n792 = ~x129 & ~n791 ;
  assign n793 = ~n790 & n792 ;
  assign n794 = ~x32 & ~x109 ;
  assign n795 = ~x31 & x109 ;
  assign n796 = ~n794 & ~n795 ;
  assign n797 = ~x106 & ~n796 ;
  assign n798 = ~x99 & x106 ;
  assign n799 = ~x129 & ~n798 ;
  assign n800 = ~n797 & n799 ;
  assign n801 = ~x33 & ~x109 ;
  assign n802 = ~x32 & x109 ;
  assign n803 = ~n801 & ~n802 ;
  assign n804 = ~x106 & ~n803 ;
  assign n805 = ~x90 & x106 ;
  assign n806 = ~x129 & ~n805 ;
  assign n807 = ~n804 & n806 ;
  assign n808 = ~x34 & ~x109 ;
  assign n809 = ~x33 & x109 ;
  assign n810 = ~n808 & ~n809 ;
  assign n811 = ~x106 & ~n810 ;
  assign n812 = ~x91 & x106 ;
  assign n813 = ~x129 & ~n812 ;
  assign n814 = ~n811 & n813 ;
  assign n815 = ~x35 & ~x109 ;
  assign n816 = ~x34 & x109 ;
  assign n817 = ~n815 & ~n816 ;
  assign n818 = ~x106 & ~n817 ;
  assign n819 = ~x92 & x106 ;
  assign n820 = ~x129 & ~n819 ;
  assign n821 = ~n818 & n820 ;
  assign n822 = ~x36 & ~x109 ;
  assign n823 = ~x35 & x109 ;
  assign n824 = ~n822 & ~n823 ;
  assign n825 = ~x106 & ~n824 ;
  assign n826 = ~x98 & x106 ;
  assign n827 = ~x129 & ~n826 ;
  assign n828 = ~n825 & n827 ;
  assign n829 = ~x37 & ~x109 ;
  assign n830 = ~x36 & x109 ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = ~x106 & ~n831 ;
  assign n833 = ~x93 & x106 ;
  assign n834 = ~x129 & ~n833 ;
  assign n835 = ~n832 & n834 ;
  assign n843 = x82 & ~n298 ;
  assign n847 = ~x38 & n843 ;
  assign n836 = ~x45 & ~x50 ;
  assign n837 = n281 & n836 ;
  assign n838 = n534 & n837 ;
  assign n839 = x82 & n291 ;
  assign n840 = n421 & n839 ;
  assign n841 = n838 & n840 ;
  assign n842 = n841 ^ x82 ;
  assign n844 = ~x38 & n284 ;
  assign n845 = ~n843 & n844 ;
  assign n846 = ~n842 & n845 ;
  assign n848 = n847 ^ n846 ;
  assign n856 = ~x45 & ~x48 ;
  assign n857 = n281 & n856 ;
  assign n858 = n534 & n857 ;
  assign n859 = n291 & n293 ;
  assign n860 = ~x40 & ~x50 ;
  assign n861 = n274 & n860 ;
  assign n862 = n859 & n861 ;
  assign n863 = n858 & n862 ;
  assign n849 = ~x44 & x82 ;
  assign n850 = ~x40 & ~x42 ;
  assign n851 = x38 & n850 ;
  assign n852 = n849 & n851 ;
  assign n853 = x74 & ~n284 ;
  assign n864 = n446 & n853 ;
  assign n865 = ~n852 & n864 ;
  assign n866 = ~n863 & n865 ;
  assign n854 = ~x129 & ~n853 ;
  assign n855 = ~n852 & n854 ;
  assign n867 = n866 ^ n855 ;
  assign n868 = ~n848 & n867 ;
  assign n869 = x109 & n564 ;
  assign n870 = x39 & ~n869 ;
  assign n871 = ~x51 & x109 ;
  assign n872 = n587 & n871 ;
  assign n873 = ~x106 & ~n872 ;
  assign n874 = ~n870 & n873 ;
  assign n875 = ~x129 & ~n874 ;
  assign n878 = x82 & ~n274 ;
  assign n882 = ~x40 & n878 ;
  assign n876 = n283 & n296 ;
  assign n877 = n876 ^ x82 ;
  assign n879 = ~x40 & n284 ;
  assign n880 = ~n878 & n879 ;
  assign n881 = ~n877 & n880 ;
  assign n883 = n882 ^ n881 ;
  assign n884 = ~x42 & n849 ;
  assign n885 = x40 & n884 ;
  assign n886 = ~x129 & ~n885 ;
  assign n887 = ~n883 & n886 ;
  assign n896 = x73 & ~n284 ;
  assign n900 = n887 & ~n896 ;
  assign n888 = ~x46 & n270 ;
  assign n889 = n273 & n888 ;
  assign n890 = ~x2 & ~x45 ;
  assign n891 = n281 & n890 ;
  assign n892 = n277 & n279 ;
  assign n893 = n891 & n892 ;
  assign n894 = n889 & n893 ;
  assign n895 = n274 & n894 ;
  assign n897 = x82 & n896 ;
  assign n898 = ~n895 & n897 ;
  assign n899 = n887 & n898 ;
  assign n901 = n900 ^ n899 ;
  assign n902 = x82 & n284 ;
  assign n903 = n295 & n902 ;
  assign n904 = n290 & n903 ;
  assign n905 = n904 ^ n440 ;
  assign n909 = ~x41 & n905 ;
  assign n906 = ~x41 & x82 ;
  assign n907 = ~n547 & n906 ;
  assign n908 = ~n905 & n907 ;
  assign n910 = n909 ^ n908 ;
  assign n911 = x41 & n884 ;
  assign n912 = n272 & n911 ;
  assign n913 = ~x129 & ~n912 ;
  assign n914 = ~n910 & n913 ;
  assign n917 = x76 & ~n284 ;
  assign n921 = n914 & ~n917 ;
  assign n915 = n290 & n295 ;
  assign n916 = n485 & n915 ;
  assign n918 = x82 & n917 ;
  assign n919 = ~n916 & n918 ;
  assign n920 = n914 & n919 ;
  assign n922 = n921 ^ n920 ;
  assign n938 = n850 & n894 ;
  assign n928 = x44 & x82 ;
  assign n932 = ~x42 & n928 ;
  assign n923 = ~x40 & x82 ;
  assign n924 = n273 & n923 ;
  assign n925 = n888 & n924 ;
  assign n926 = n893 & n925 ;
  assign n927 = n926 ^ x82 ;
  assign n929 = ~x42 & n284 ;
  assign n930 = ~n928 & n929 ;
  assign n931 = ~n927 & n930 ;
  assign n933 = n932 ^ n931 ;
  assign n934 = x42 & n849 ;
  assign n935 = ~x129 & ~n934 ;
  assign n939 = x72 & ~n285 ;
  assign n940 = n935 & n939 ;
  assign n941 = ~n933 & n940 ;
  assign n942 = ~n938 & n941 ;
  assign n936 = ~x72 & n935 ;
  assign n937 = ~n933 & n936 ;
  assign n943 = n942 ^ n937 ;
  assign n944 = n419 & n893 ;
  assign n945 = x82 & ~n944 ;
  assign n946 = x77 & ~n284 ;
  assign n947 = ~n945 & n946 ;
  assign n948 = n281 & n427 ;
  assign n949 = n277 & n433 ;
  assign n950 = n948 & n949 ;
  assign n952 = n284 & n950 ;
  assign n951 = n440 & ~n950 ;
  assign n953 = n952 ^ n951 ;
  assign n957 = ~x43 & n953 ;
  assign n954 = ~x43 & x82 ;
  assign n955 = ~n419 & n954 ;
  assign n956 = ~n953 & n955 ;
  assign n958 = n957 ^ n956 ;
  assign n959 = n849 & n850 ;
  assign n960 = n292 & n959 ;
  assign n961 = x43 & n960 ;
  assign n962 = ~x129 & ~n961 ;
  assign n963 = ~n958 & n962 ;
  assign n964 = ~n947 & n963 ;
  assign n965 = x82 & ~n938 ;
  assign n966 = ~x67 & ~n284 ;
  assign n967 = x44 & n284 ;
  assign n968 = ~n966 & ~n967 ;
  assign n969 = ~n965 & n968 ;
  assign n970 = ~x129 & ~n928 ;
  assign n971 = ~n969 & n970 ;
  assign n972 = n425 & n427 ;
  assign n973 = x82 & ~n972 ;
  assign n974 = n284 & ~n973 ;
  assign n975 = n291 & n421 ;
  assign n976 = ~x50 & n484 ;
  assign n977 = n975 & n976 ;
  assign n978 = x82 & ~n977 ;
  assign n979 = ~n974 & ~n978 ;
  assign n980 = ~x45 & ~n979 ;
  assign n981 = n277 & n427 ;
  assign n982 = n425 & n981 ;
  assign n983 = n276 & n982 ;
  assign n984 = x68 & ~n284 ;
  assign n985 = x82 & n984 ;
  assign n986 = ~n983 & n985 ;
  assign n987 = n986 ^ n984 ;
  assign n988 = x45 & x82 ;
  assign n989 = n977 & n988 ;
  assign n990 = ~x129 & ~n989 ;
  assign n991 = ~n987 & n990 ;
  assign n992 = ~n980 & n991 ;
  assign n993 = ~x75 & ~n284 ;
  assign n995 = x82 & n273 ;
  assign n996 = ~n993 & n995 ;
  assign n997 = n893 & n996 ;
  assign n994 = ~x82 & ~n993 ;
  assign n998 = n997 ^ n994 ;
  assign n999 = n485 & ~n998 ;
  assign n1002 = x82 & n976 ;
  assign n1000 = ~x75 & n285 ;
  assign n1003 = x46 & ~n285 ;
  assign n1004 = ~n1000 & n1003 ;
  assign n1005 = ~n1002 & n1004 ;
  assign n1006 = ~n999 & n1005 ;
  assign n1001 = ~n999 & ~n1000 ;
  assign n1007 = n1006 ^ n1001 ;
  assign n1008 = ~x129 & ~n1007 ;
  assign n1010 = n284 & n858 ;
  assign n1009 = n440 & ~n858 ;
  assign n1011 = n1010 ^ n1009 ;
  assign n1015 = ~x47 & n1011 ;
  assign n1012 = ~x47 & x82 ;
  assign n1013 = ~n276 & n1012 ;
  assign n1014 = ~n1011 & n1013 ;
  assign n1016 = n1015 ^ n1014 ;
  assign n1017 = ~x43 & x47 ;
  assign n1018 = n960 & n1017 ;
  assign n1019 = ~x129 & ~n1018 ;
  assign n1020 = ~n1016 & n1019 ;
  assign n1022 = x64 & ~n284 ;
  assign n1026 = n1020 & ~n1022 ;
  assign n1021 = n276 & n858 ;
  assign n1023 = x82 & n1022 ;
  assign n1024 = ~n1021 & n1023 ;
  assign n1025 = n1020 & n1024 ;
  assign n1027 = n1026 ^ n1025 ;
  assign n1028 = x82 & n859 ;
  assign n1029 = n976 & n1028 ;
  assign n1030 = n1029 ^ x82 ;
  assign n1038 = ~x48 & n1030 ;
  assign n1031 = ~x45 & x82 ;
  assign n1032 = n281 & n1031 ;
  assign n1033 = n534 & n1032 ;
  assign n1034 = n1033 ^ x82 ;
  assign n1035 = ~x48 & n284 ;
  assign n1036 = ~n1034 & n1035 ;
  assign n1037 = ~n1030 & n1036 ;
  assign n1039 = n1038 ^ n1037 ;
  assign n1040 = x48 & n293 ;
  assign n1041 = n960 & n1040 ;
  assign n1042 = ~x129 & ~n1041 ;
  assign n1043 = ~n1039 & n1042 ;
  assign n1047 = x62 & ~n284 ;
  assign n1051 = n1043 & ~n1047 ;
  assign n1044 = n420 & n534 ;
  assign n1045 = ~x47 & n276 ;
  assign n1046 = n1044 & n1045 ;
  assign n1048 = x82 & n1047 ;
  assign n1049 = ~n1046 & n1048 ;
  assign n1050 = n1043 & n1049 ;
  assign n1052 = n1051 ^ n1050 ;
  assign n1053 = n488 & ~n534 ;
  assign n1054 = ~x24 & ~x40 ;
  assign n1055 = n274 & n1054 ;
  assign n1056 = n888 & n1055 ;
  assign n1057 = x49 & n273 ;
  assign n1058 = n426 & n1057 ;
  assign n1059 = n1056 & n1058 ;
  assign n1060 = n1059 ^ x49 ;
  assign n1061 = x82 & ~n1060 ;
  assign n1062 = ~n1053 & n1061 ;
  assign n1063 = n1062 ^ x82 ;
  assign n1064 = x82 & n482 ;
  assign n1065 = n484 & n1064 ;
  assign n1066 = n487 & n1065 ;
  assign n1067 = n1066 ^ x82 ;
  assign n1068 = x49 & n440 ;
  assign n1069 = ~x69 & ~n284 ;
  assign n1070 = ~n1068 & n1069 ;
  assign n1071 = ~n1067 & n1070 ;
  assign n1072 = n1071 ^ n1068 ;
  assign n1073 = ~x129 & ~n1072 ;
  assign n1074 = ~n1063 & n1073 ;
  assign n1075 = n1074 ^ x129 ;
  assign n1089 = ~x50 & n859 ;
  assign n1090 = n858 & n1089 ;
  assign n1091 = x82 & ~n1090 ;
  assign n1079 = x82 & ~n484 ;
  assign n1083 = ~x50 & n1079 ;
  assign n1076 = n295 & n839 ;
  assign n1077 = n290 & n1076 ;
  assign n1078 = n1077 ^ x82 ;
  assign n1080 = ~x50 & n284 ;
  assign n1081 = ~n1079 & n1080 ;
  assign n1082 = ~n1078 & n1081 ;
  assign n1084 = n1083 ^ n1082 ;
  assign n1085 = x50 & x82 ;
  assign n1086 = n484 & n1085 ;
  assign n1087 = ~x129 & ~n1086 ;
  assign n1092 = x66 & ~n284 ;
  assign n1093 = n1087 & n1092 ;
  assign n1094 = ~n1084 & n1093 ;
  assign n1095 = ~n1091 & n1094 ;
  assign n1088 = ~n1084 & n1087 ;
  assign n1096 = n1095 ^ n1088 ;
  assign n1097 = x51 & ~x109 ;
  assign n1098 = ~x106 & ~n871 ;
  assign n1099 = ~n1097 & n1098 ;
  assign n1100 = ~x129 & ~n1099 ;
  assign n1101 = x52 & ~n871 ;
  assign n1102 = ~x106 & ~n869 ;
  assign n1103 = ~n1101 & n1102 ;
  assign n1104 = ~x129 & ~n1103 ;
  assign n1105 = ~x116 & n698 ;
  assign n1106 = ~x53 & x97 ;
  assign n1107 = x58 & x116 ;
  assign n1108 = ~x58 & n567 ;
  assign n1109 = ~n702 & n1108 ;
  assign n1110 = ~n1107 & ~n1109 ;
  assign n1111 = n1106 & ~n1110 ;
  assign n1112 = ~n1105 & ~n1111 ;
  assign n1113 = n556 & n625 ;
  assign n1114 = ~n1112 & n1113 ;
  assign n1115 = ~n284 & n972 ;
  assign n1116 = n548 & n1115 ;
  assign n1117 = ~x129 & ~n285 ;
  assign n1118 = ~n1116 & n1117 ;
  assign n1119 = ~x123 & ~x129 ;
  assign n1120 = x114 & ~x122 ;
  assign n1121 = n1119 & n1120 ;
  assign n1131 = x37 & ~x58 ;
  assign n1132 = ~x116 & n1131 ;
  assign n1128 = x26 & ~x58 ;
  assign n1129 = x94 & x116 ;
  assign n1130 = n1128 & n1129 ;
  assign n1133 = n1132 ^ n1130 ;
  assign n1124 = ~x26 & x58 ;
  assign n1125 = ~x94 & ~x116 ;
  assign n1126 = n1124 & n1125 ;
  assign n1127 = n1126 ^ n1124 ;
  assign n1134 = n1133 ^ n1127 ;
  assign n1122 = ~x26 & x37 ;
  assign n1137 = n555 & n1122 ;
  assign n1138 = n1134 & n1137 ;
  assign n1136 = ~x58 & n1122 ;
  assign n1139 = n1138 ^ n1136 ;
  assign n1135 = ~x53 & n1134 ;
  assign n1140 = n1139 ^ n1135 ;
  assign n1147 = n556 & n1140 ;
  assign n1145 = x85 & n555 ;
  assign n1146 = n1122 & n1145 ;
  assign n1148 = n1147 ^ n1146 ;
  assign n1141 = n556 & n1122 ;
  assign n1142 = n555 & n1141 ;
  assign n1143 = ~n1140 & n1142 ;
  assign n1123 = n694 & n1122 ;
  assign n1144 = n1143 ^ n1123 ;
  assign n1149 = n1148 ^ n1144 ;
  assign n1150 = n230 & n1149 ;
  assign n1169 = x57 & ~x58 ;
  assign n1170 = n669 & n1169 ;
  assign n1174 = n230 & n1170 ;
  assign n1153 = ~x26 & ~x58 ;
  assign n1154 = ~x85 & n1153 ;
  assign n1151 = x26 & ~x53 ;
  assign n1152 = ~x58 & n1151 ;
  assign n1155 = n1154 ^ n1152 ;
  assign n1156 = n1155 ^ n1145 ;
  assign n1163 = x57 & x116 ;
  assign n1164 = ~n1156 & n1163 ;
  assign n1160 = x60 & n1107 ;
  assign n1165 = n669 & ~n1160 ;
  assign n1166 = n1164 & n1165 ;
  assign n1161 = ~x57 & n669 ;
  assign n1162 = ~n1160 & n1161 ;
  assign n1167 = n1166 ^ n1162 ;
  assign n1157 = x57 & ~n669 ;
  assign n1158 = n1156 & n1157 ;
  assign n1159 = n1158 ^ n669 ;
  assign n1168 = n1167 ^ n1159 ;
  assign n1171 = ~x27 & n230 ;
  assign n1172 = ~n1170 & n1171 ;
  assign n1173 = n1168 & n1172 ;
  assign n1175 = n1174 ^ n1173 ;
  assign n1176 = n585 & n720 ;
  assign n1177 = ~x58 & n649 ;
  assign n1178 = n589 & n1177 ;
  assign n1179 = ~n1176 & ~n1178 ;
  assign n1180 = n230 & n658 ;
  assign n1181 = ~n1179 & n1180 ;
  assign n1182 = x59 & ~x116 ;
  assign n1197 = x26 & n1182 ;
  assign n1198 = n685 & n1197 ;
  assign n1193 = n1145 & n1182 ;
  assign n1194 = n1193 ^ x85 ;
  assign n1187 = x59 & n555 ;
  assign n1188 = n570 & n1187 ;
  assign n1185 = x96 & n555 ;
  assign n1186 = ~n570 & n1185 ;
  assign n1189 = n1188 ^ n1186 ;
  assign n1190 = n562 & n1182 ;
  assign n1191 = ~x85 & ~n1190 ;
  assign n1192 = ~n1189 & n1191 ;
  assign n1195 = n1194 ^ n1192 ;
  assign n1196 = n585 & ~n1195 ;
  assign n1199 = n1198 ^ n1196 ;
  assign n1183 = x27 & n1182 ;
  assign n1184 = n685 & n1183 ;
  assign n1200 = n1199 ^ n1184 ;
  assign n1201 = n230 & n1200 ;
  assign n1202 = ~x117 & ~x122 ;
  assign n1203 = x60 & ~n1202 ;
  assign n1204 = x123 & n1202 ;
  assign n1205 = ~n1203 & ~n1204 ;
  assign n1206 = ~x114 & ~x122 ;
  assign n1207 = x123 & ~x129 ;
  assign n1208 = n1206 & n1207 ;
  assign n1209 = x136 & ~x137 ;
  assign n1210 = x131 & x132 ;
  assign n1211 = x133 & n1210 ;
  assign n1212 = ~x138 & n1211 ;
  assign n1213 = n1209 & n1212 ;
  assign n1214 = x140 & n1213 ;
  assign n1215 = ~x62 & ~n1213 ;
  assign n1216 = ~x129 & ~n1215 ;
  assign n1217 = ~n1214 & n1216 ;
  assign n1218 = x142 & n1213 ;
  assign n1219 = ~x63 & ~n1213 ;
  assign n1220 = ~x129 & ~n1219 ;
  assign n1221 = ~n1218 & n1220 ;
  assign n1222 = x139 & n1213 ;
  assign n1223 = ~x64 & ~n1213 ;
  assign n1224 = ~x129 & ~n1223 ;
  assign n1225 = ~n1222 & n1224 ;
  assign n1226 = x146 & n1213 ;
  assign n1227 = ~x65 & ~n1213 ;
  assign n1228 = ~x129 & ~n1227 ;
  assign n1229 = ~n1226 & n1228 ;
  assign n1230 = ~x136 & ~x137 ;
  assign n1231 = n1212 & n1230 ;
  assign n1232 = x143 & n1231 ;
  assign n1233 = ~x66 & ~n1231 ;
  assign n1234 = ~x129 & ~n1233 ;
  assign n1235 = ~n1232 & n1234 ;
  assign n1236 = x139 & n1231 ;
  assign n1237 = ~x67 & ~n1231 ;
  assign n1238 = ~x129 & ~n1237 ;
  assign n1239 = ~n1236 & n1238 ;
  assign n1240 = x141 & n1213 ;
  assign n1241 = ~x68 & ~n1213 ;
  assign n1242 = ~x129 & ~n1241 ;
  assign n1243 = ~n1240 & n1242 ;
  assign n1244 = x143 & n1213 ;
  assign n1245 = ~x69 & ~n1213 ;
  assign n1246 = ~x129 & ~n1245 ;
  assign n1247 = ~n1244 & n1246 ;
  assign n1248 = x144 & n1213 ;
  assign n1249 = ~x70 & ~n1213 ;
  assign n1250 = ~x129 & ~n1249 ;
  assign n1251 = ~n1248 & n1250 ;
  assign n1252 = x145 & n1213 ;
  assign n1253 = ~x71 & ~n1213 ;
  assign n1254 = ~x129 & ~n1253 ;
  assign n1255 = ~n1252 & n1254 ;
  assign n1256 = x140 & n1231 ;
  assign n1257 = ~x72 & ~n1231 ;
  assign n1258 = ~x129 & ~n1257 ;
  assign n1259 = ~n1256 & n1258 ;
  assign n1260 = x141 & n1231 ;
  assign n1261 = ~x73 & ~n1231 ;
  assign n1262 = ~x129 & ~n1261 ;
  assign n1263 = ~n1260 & n1262 ;
  assign n1264 = x142 & n1231 ;
  assign n1265 = ~x74 & ~n1231 ;
  assign n1266 = ~x129 & ~n1265 ;
  assign n1267 = ~n1264 & n1266 ;
  assign n1268 = x144 & n1231 ;
  assign n1269 = ~x75 & ~n1231 ;
  assign n1270 = ~x129 & ~n1269 ;
  assign n1271 = ~n1268 & n1270 ;
  assign n1272 = x145 & n1231 ;
  assign n1273 = ~x76 & ~n1231 ;
  assign n1274 = ~x129 & ~n1273 ;
  assign n1275 = ~n1272 & n1274 ;
  assign n1276 = x146 & n1231 ;
  assign n1277 = ~x77 & ~n1231 ;
  assign n1278 = ~x129 & ~n1277 ;
  assign n1279 = ~n1276 & n1278 ;
  assign n1280 = ~x136 & x137 ;
  assign n1281 = n1212 & n1280 ;
  assign n1282 = ~x142 & n1281 ;
  assign n1283 = ~x78 & ~n1281 ;
  assign n1284 = ~x129 & ~n1283 ;
  assign n1285 = ~n1282 & n1284 ;
  assign n1286 = ~x143 & n1281 ;
  assign n1287 = ~x79 & ~n1281 ;
  assign n1288 = ~x129 & ~n1287 ;
  assign n1289 = ~n1286 & n1288 ;
  assign n1290 = ~x144 & n1281 ;
  assign n1291 = ~x80 & ~n1281 ;
  assign n1292 = ~x129 & ~n1291 ;
  assign n1293 = ~n1290 & n1292 ;
  assign n1294 = ~x145 & n1281 ;
  assign n1295 = ~x81 & ~n1281 ;
  assign n1296 = ~x129 & ~n1295 ;
  assign n1297 = ~n1294 & n1296 ;
  assign n1298 = ~x146 & n1281 ;
  assign n1299 = ~x82 & ~n1281 ;
  assign n1300 = ~x129 & ~n1299 ;
  assign n1301 = ~n1298 & n1300 ;
  assign n1302 = x136 & ~x138 ;
  assign n1303 = x31 & n1302 ;
  assign n1304 = x115 & x138 ;
  assign n1305 = ~x87 & ~x138 ;
  assign n1306 = ~x136 & ~n1305 ;
  assign n1307 = ~n1304 & n1306 ;
  assign n1308 = ~n1303 & ~n1307 ;
  assign n1309 = x137 & ~n1308 ;
  assign n1310 = x62 & ~x138 ;
  assign n1311 = ~x89 & x138 ;
  assign n1312 = x136 & ~n1311 ;
  assign n1313 = ~n1310 & n1312 ;
  assign n1314 = x72 & ~x138 ;
  assign n1315 = ~x119 & x138 ;
  assign n1316 = ~x136 & ~n1315 ;
  assign n1317 = ~n1314 & n1316 ;
  assign n1318 = ~n1313 & ~n1317 ;
  assign n1319 = ~x137 & ~n1318 ;
  assign n1320 = ~n1309 & ~n1319 ;
  assign n1321 = ~x141 & n1281 ;
  assign n1322 = ~x84 & ~n1281 ;
  assign n1323 = ~x129 & ~n1322 ;
  assign n1324 = ~n1321 & n1323 ;
  assign n1325 = ~x97 & n567 ;
  assign n1326 = n618 & ~n1325 ;
  assign n1327 = x96 & n1326 ;
  assign n1328 = ~n582 & ~n1327 ;
  assign n1329 = n613 & n625 ;
  assign n1330 = ~n1328 & n1329 ;
  assign n1331 = ~x139 & n1281 ;
  assign n1332 = ~x86 & ~n1281 ;
  assign n1333 = ~x129 & ~n1332 ;
  assign n1334 = ~n1331 & n1333 ;
  assign n1335 = ~x140 & n1281 ;
  assign n1336 = ~x87 & ~n1281 ;
  assign n1337 = ~x129 & ~n1336 ;
  assign n1338 = ~n1335 & n1337 ;
  assign n1339 = x137 & n1302 ;
  assign n1340 = n1211 & n1339 ;
  assign n1341 = ~x139 & n1340 ;
  assign n1342 = ~x88 & ~n1340 ;
  assign n1343 = ~x129 & ~n1342 ;
  assign n1344 = ~n1341 & n1343 ;
  assign n1345 = ~x140 & n1340 ;
  assign n1346 = ~x89 & ~n1340 ;
  assign n1347 = ~x129 & ~n1346 ;
  assign n1348 = ~n1345 & n1347 ;
  assign n1349 = ~x142 & n1340 ;
  assign n1350 = ~x90 & ~n1340 ;
  assign n1351 = ~x129 & ~n1350 ;
  assign n1352 = ~n1349 & n1351 ;
  assign n1353 = ~x143 & n1340 ;
  assign n1354 = ~x91 & ~n1340 ;
  assign n1355 = ~x129 & ~n1354 ;
  assign n1356 = ~n1353 & n1355 ;
  assign n1357 = ~x144 & n1340 ;
  assign n1358 = ~x92 & ~n1340 ;
  assign n1359 = ~x129 & ~n1358 ;
  assign n1360 = ~n1357 & n1359 ;
  assign n1361 = ~x146 & n1340 ;
  assign n1362 = ~x93 & ~n1340 ;
  assign n1363 = ~x129 & ~n1362 ;
  assign n1364 = ~n1361 & n1363 ;
  assign n1365 = x82 & x138 ;
  assign n1366 = n1230 & n1365 ;
  assign n1367 = n1211 & n1366 ;
  assign n1368 = ~x142 & n1367 ;
  assign n1369 = ~x94 & ~n1367 ;
  assign n1370 = ~x129 & ~n1369 ;
  assign n1371 = ~n1368 & n1370 ;
  assign n1372 = ~x3 & ~x110 ;
  assign n1373 = ~n1211 & ~n1372 ;
  assign n1374 = ~n1367 & ~n1373 ;
  assign n1375 = x95 & n1374 ;
  assign n1376 = x143 & n1367 ;
  assign n1377 = ~n1375 & ~n1376 ;
  assign n1378 = ~x129 & ~n1377 ;
  assign n1379 = x96 & n1374 ;
  assign n1380 = x146 & n1367 ;
  assign n1381 = ~n1379 & ~n1380 ;
  assign n1382 = ~x129 & ~n1381 ;
  assign n1383 = x97 & n1374 ;
  assign n1384 = x145 & n1367 ;
  assign n1385 = ~n1383 & ~n1384 ;
  assign n1386 = ~x129 & ~n1385 ;
  assign n1387 = ~x145 & n1340 ;
  assign n1388 = ~x98 & ~n1340 ;
  assign n1389 = ~x129 & ~n1388 ;
  assign n1390 = ~n1387 & n1389 ;
  assign n1391 = ~x141 & n1340 ;
  assign n1392 = ~x99 & ~n1340 ;
  assign n1393 = ~x129 & ~n1392 ;
  assign n1394 = ~n1391 & n1393 ;
  assign n1395 = x100 & n1374 ;
  assign n1396 = x144 & n1367 ;
  assign n1397 = ~n1395 & ~n1396 ;
  assign n1398 = ~x129 & ~n1397 ;
  assign n1399 = x37 & n1302 ;
  assign n1400 = ~x96 & x138 ;
  assign n1401 = ~x82 & ~x138 ;
  assign n1402 = ~x136 & ~n1401 ;
  assign n1403 = ~n1400 & n1402 ;
  assign n1404 = ~n1399 & ~n1403 ;
  assign n1405 = x137 & ~n1404 ;
  assign n1406 = x65 & ~x138 ;
  assign n1407 = ~x93 & x138 ;
  assign n1408 = x136 & ~n1407 ;
  assign n1409 = ~n1406 & n1408 ;
  assign n1410 = x77 & ~x138 ;
  assign n1411 = ~x124 & x138 ;
  assign n1412 = ~x136 & ~n1411 ;
  assign n1413 = ~n1410 & n1412 ;
  assign n1414 = ~n1409 & ~n1413 ;
  assign n1415 = ~x137 & ~n1414 ;
  assign n1416 = ~n1405 & ~n1415 ;
  assign n1417 = x91 & n1209 ;
  assign n1418 = x95 & n1280 ;
  assign n1419 = ~n1417 & ~n1418 ;
  assign n1420 = x138 & ~n1419 ;
  assign n1421 = ~x34 & x136 ;
  assign n1422 = ~x79 & ~x136 ;
  assign n1423 = x137 & ~n1422 ;
  assign n1424 = ~n1421 & n1423 ;
  assign n1425 = x69 & x136 ;
  assign n1426 = x66 & ~x136 ;
  assign n1427 = ~x137 & ~n1426 ;
  assign n1428 = ~n1425 & n1427 ;
  assign n1429 = ~n1424 & ~n1428 ;
  assign n1430 = ~x138 & ~n1429 ;
  assign n1431 = ~n1420 & ~n1430 ;
  assign n1432 = x90 & n1209 ;
  assign n1433 = x94 & n1280 ;
  assign n1434 = ~n1432 & ~n1433 ;
  assign n1435 = x138 & ~n1434 ;
  assign n1436 = ~x33 & x136 ;
  assign n1437 = ~x78 & ~x136 ;
  assign n1438 = x137 & ~n1437 ;
  assign n1439 = ~n1436 & n1438 ;
  assign n1440 = x63 & x136 ;
  assign n1441 = x74 & ~x136 ;
  assign n1442 = ~x137 & ~n1441 ;
  assign n1443 = ~n1440 & n1442 ;
  assign n1444 = ~n1439 & ~n1443 ;
  assign n1445 = ~x138 & ~n1444 ;
  assign n1446 = ~n1435 & ~n1445 ;
  assign n1447 = x99 & n1209 ;
  assign n1448 = ~x112 & n1280 ;
  assign n1449 = ~n1447 & ~n1448 ;
  assign n1450 = x138 & ~n1449 ;
  assign n1451 = ~x32 & x136 ;
  assign n1452 = ~x84 & ~x136 ;
  assign n1453 = x137 & ~n1452 ;
  assign n1454 = ~n1451 & n1453 ;
  assign n1455 = x68 & x136 ;
  assign n1456 = x73 & ~x136 ;
  assign n1457 = ~x137 & ~n1456 ;
  assign n1458 = ~n1455 & n1457 ;
  assign n1459 = ~n1454 & ~n1458 ;
  assign n1460 = ~x138 & ~n1459 ;
  assign n1461 = ~n1450 & ~n1460 ;
  assign n1462 = x35 & n1302 ;
  assign n1463 = ~x100 & x138 ;
  assign n1464 = ~x80 & ~x138 ;
  assign n1465 = ~x136 & ~n1464 ;
  assign n1466 = ~n1463 & n1465 ;
  assign n1467 = ~n1462 & ~n1466 ;
  assign n1468 = x137 & ~n1467 ;
  assign n1469 = x70 & ~x138 ;
  assign n1470 = ~x92 & x138 ;
  assign n1471 = x136 & ~n1470 ;
  assign n1472 = ~n1469 & n1471 ;
  assign n1473 = x75 & ~x138 ;
  assign n1474 = ~x125 & x138 ;
  assign n1475 = ~x136 & ~n1474 ;
  assign n1476 = ~n1473 & n1475 ;
  assign n1477 = ~n1472 & ~n1476 ;
  assign n1478 = ~x137 & ~n1477 ;
  assign n1479 = ~n1468 & ~n1478 ;
  assign n1480 = ~x26 & n613 ;
  assign n1481 = n1326 & n1480 ;
  assign n1482 = ~n617 & ~n1481 ;
  assign n1483 = n230 & ~n1482 ;
  assign n1484 = x36 & n1302 ;
  assign n1485 = ~x97 & x138 ;
  assign n1486 = ~x81 & ~x138 ;
  assign n1487 = ~x136 & ~n1486 ;
  assign n1488 = ~n1485 & n1487 ;
  assign n1489 = ~n1484 & ~n1488 ;
  assign n1490 = x137 & ~n1489 ;
  assign n1491 = x71 & ~x138 ;
  assign n1492 = ~x98 & x138 ;
  assign n1493 = x136 & ~n1492 ;
  assign n1494 = ~n1491 & n1493 ;
  assign n1495 = x76 & ~x138 ;
  assign n1496 = ~x23 & x138 ;
  assign n1497 = ~x136 & ~n1496 ;
  assign n1498 = ~n1495 & n1497 ;
  assign n1499 = ~n1494 & ~n1498 ;
  assign n1500 = ~x137 & ~n1499 ;
  assign n1501 = ~n1490 & ~n1500 ;
  assign n1502 = x30 & n1302 ;
  assign n1503 = ~x111 & x138 ;
  assign n1504 = ~x86 & ~x138 ;
  assign n1505 = ~x136 & ~n1504 ;
  assign n1506 = ~n1503 & n1505 ;
  assign n1507 = ~n1502 & ~n1506 ;
  assign n1508 = x137 & ~n1507 ;
  assign n1509 = x64 & ~x138 ;
  assign n1510 = ~x88 & x138 ;
  assign n1511 = x136 & ~n1510 ;
  assign n1512 = ~n1509 & n1511 ;
  assign n1513 = x67 & ~x138 ;
  assign n1514 = ~x120 & x138 ;
  assign n1515 = ~x136 & ~n1514 ;
  assign n1516 = ~n1513 & n1515 ;
  assign n1517 = ~n1512 & ~n1516 ;
  assign n1518 = ~x137 & ~n1517 ;
  assign n1519 = ~n1508 & ~n1518 ;
  assign n1520 = ~x26 & n566 ;
  assign n1521 = ~n592 & ~n1520 ;
  assign n1522 = x116 & n230 ;
  assign n1523 = ~n1521 & n1522 ;
  assign n1524 = ~x97 & n716 ;
  assign n1525 = ~n698 & ~n1524 ;
  assign n1526 = n1522 & ~n1525 ;
  assign n1527 = ~x139 & n1366 ;
  assign n1528 = ~x129 & n1211 ;
  assign n1529 = ~x111 & ~n1366 ;
  assign n1530 = n1528 & ~n1529 ;
  assign n1531 = ~n1527 & n1530 ;
  assign n1532 = x112 & ~n1366 ;
  assign n1533 = ~x141 & n1366 ;
  assign n1534 = n1528 & ~n1533 ;
  assign n1535 = ~n1532 & n1534 ;
  assign n1536 = ~x11 & ~x22 ;
  assign n1537 = x54 & n1536 ;
  assign n1538 = ~x54 & x113 ;
  assign n1539 = n230 & ~n1538 ;
  assign n1540 = ~n1537 & n1539 ;
  assign n1541 = x115 & ~n1366 ;
  assign n1542 = ~x140 & n1366 ;
  assign n1543 = n1528 & ~n1542 ;
  assign n1544 = ~n1541 & n1543 ;
  assign n1545 = x54 & n230 ;
  assign n1546 = ~x4 & ~x9 ;
  assign n1547 = n235 & n1546 ;
  assign n1548 = n1545 & ~n1547 ;
  assign n1549 = x122 & ~x129 ;
  assign n1550 = ~x54 & x118 ;
  assign n1551 = x54 & ~x59 ;
  assign n1552 = n404 & n1551 ;
  assign n1553 = ~n1550 & ~n1552 ;
  assign n1554 = ~x129 & ~n1553 ;
  assign n1555 = ~x129 & ~n567 ;
  assign n1556 = ~x120 & n1372 ;
  assign n1557 = ~x111 & ~x129 ;
  assign n1558 = ~n1556 & n1557 ;
  assign n1559 = x81 & x120 ;
  assign n1560 = ~x129 & n1559 ;
  assign n1561 = ~x129 & ~x134 ;
  assign n1562 = ~x129 & ~x135 ;
  assign n1563 = x57 & ~x129 ;
  assign n1564 = ~x96 & x125 ;
  assign n1565 = ~x3 & ~n1564 ;
  assign n1566 = ~x129 & ~n1565 ;
  assign n1567 = ~x126 & x132 ;
  assign n1568 = x133 & n1567 ;
  assign y0 = x108 ;
  assign y1 = x83 ;
  assign y2 = x104 ;
  assign y3 = x103 ;
  assign y4 = x102 ;
  assign y5 = x105 ;
  assign y6 = x107 ;
  assign y7 = x101 ;
  assign y8 = x126 ;
  assign y9 = x121 ;
  assign y10 = x1 ;
  assign y11 = x0 ;
  assign y12 = ~1'b0 ;
  assign y13 = x130 ;
  assign y14 = x128 ;
  assign y15 = ~n233 ;
  assign y16 = ~n269 ;
  assign y17 = n308 ;
  assign y18 = n319 ;
  assign y19 = n331 ;
  assign y20 = n344 ;
  assign y21 = n352 ;
  assign y22 = n359 ;
  assign y23 = n370 ;
  assign y24 = n377 ;
  assign y25 = n387 ;
  assign y26 = n394 ;
  assign y27 = n401 ;
  assign y28 = n410 ;
  assign y29 = n418 ;
  assign y30 = n450 ;
  assign y31 = n457 ;
  assign y32 = n466 ;
  assign y33 = n473 ;
  assign y34 = n480 ;
  assign y35 = n508 ;
  assign y36 = n516 ;
  assign y37 = n525 ;
  assign y38 = n528 ;
  assign y39 = n554 ;
  assign y40 = n606 ;
  assign y41 = n615 ;
  assign y42 = n627 ;
  assign y43 = n683 ;
  assign y44 = n779 ;
  assign y45 = n786 ;
  assign y46 = n793 ;
  assign y47 = n800 ;
  assign y48 = n807 ;
  assign y49 = n814 ;
  assign y50 = n821 ;
  assign y51 = n828 ;
  assign y52 = n835 ;
  assign y53 = n868 ;
  assign y54 = n875 ;
  assign y55 = n901 ;
  assign y56 = n922 ;
  assign y57 = n943 ;
  assign y58 = n964 ;
  assign y59 = n971 ;
  assign y60 = n992 ;
  assign y61 = n1008 ;
  assign y62 = n1027 ;
  assign y63 = n1052 ;
  assign y64 = ~n1075 ;
  assign y65 = n1096 ;
  assign y66 = n1100 ;
  assign y67 = n1104 ;
  assign y68 = n1114 ;
  assign y69 = ~n1118 ;
  assign y70 = n1121 ;
  assign y71 = n1150 ;
  assign y72 = n1175 ;
  assign y73 = n1181 ;
  assign y74 = n1201 ;
  assign y75 = ~n1205 ;
  assign y76 = n1208 ;
  assign y77 = ~n1217 ;
  assign y78 = ~n1221 ;
  assign y79 = ~n1225 ;
  assign y80 = ~n1229 ;
  assign y81 = ~n1235 ;
  assign y82 = ~n1239 ;
  assign y83 = ~n1243 ;
  assign y84 = ~n1247 ;
  assign y85 = ~n1251 ;
  assign y86 = ~n1255 ;
  assign y87 = ~n1259 ;
  assign y88 = ~n1263 ;
  assign y89 = ~n1267 ;
  assign y90 = ~n1271 ;
  assign y91 = ~n1275 ;
  assign y92 = ~n1279 ;
  assign y93 = n1285 ;
  assign y94 = n1289 ;
  assign y95 = n1293 ;
  assign y96 = n1297 ;
  assign y97 = n1301 ;
  assign y98 = ~n1320 ;
  assign y99 = n1324 ;
  assign y100 = n1330 ;
  assign y101 = n1334 ;
  assign y102 = n1338 ;
  assign y103 = n1344 ;
  assign y104 = n1348 ;
  assign y105 = n1352 ;
  assign y106 = n1356 ;
  assign y107 = n1360 ;
  assign y108 = n1364 ;
  assign y109 = n1371 ;
  assign y110 = n1378 ;
  assign y111 = n1382 ;
  assign y112 = n1386 ;
  assign y113 = n1390 ;
  assign y114 = n1394 ;
  assign y115 = n1398 ;
  assign y116 = ~n1416 ;
  assign y117 = ~n1431 ;
  assign y118 = ~n1446 ;
  assign y119 = ~n1461 ;
  assign y120 = ~n1479 ;
  assign y121 = n1483 ;
  assign y122 = ~n1501 ;
  assign y123 = ~n1519 ;
  assign y124 = n1523 ;
  assign y125 = n1526 ;
  assign y126 = n1531 ;
  assign y127 = n1535 ;
  assign y128 = n1540 ;
  assign y129 = ~n1119 ;
  assign y130 = n1544 ;
  assign y131 = n1548 ;
  assign y132 = ~n1549 ;
  assign y133 = n1554 ;
  assign y134 = n1555 ;
  assign y135 = n1558 ;
  assign y136 = n1560 ;
  assign y137 = ~n1561 ;
  assign y138 = ~n1562 ;
  assign y139 = n1563 ;
  assign y140 = n1566 ;
  assign y141 = n1568 ;
endmodule
