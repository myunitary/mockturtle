module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 ;
  assign n50 = x8 ^ x0 ;
  assign n54 = x9 ^ x1 ;
  assign n55 = ~n50 & ~n54 ;
  assign n57 = x10 ^ x2 ;
  assign n63 = x11 ^ x3 ;
  assign n64 = ~n57 & ~n63 ;
  assign n65 = n55 & n64 ;
  assign n67 = x12 ^ x4 ;
  assign n71 = x13 ^ x5 ;
  assign n72 = ~n67 & ~n71 ;
  assign n74 = x14 ^ x6 ;
  assign n84 = x15 ^ x7 ;
  assign n85 = ~n74 & ~n84 ;
  assign n86 = n72 & n85 ;
  assign n87 = n65 & n86 ;
  assign n75 = x7 & x15 ;
  assign n76 = n75 ^ x7 ;
  assign n77 = n74 & n76 ;
  assign n78 = n77 ^ n76 ;
  assign n73 = x6 & ~x14 ;
  assign n79 = n78 ^ n73 ;
  assign n80 = n72 & n79 ;
  assign n68 = x5 & ~x13 ;
  assign n69 = ~n67 & n68 ;
  assign n66 = x4 & ~x12 ;
  assign n70 = n69 ^ n66 ;
  assign n81 = n80 ^ n70 ;
  assign n82 = n65 & n81 ;
  assign n58 = x3 & ~x11 ;
  assign n59 = ~n57 & n58 ;
  assign n56 = x2 & ~x10 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n55 & n60 ;
  assign n51 = x1 & ~x9 ;
  assign n52 = ~n50 & n51 ;
  assign n49 = x0 & ~x8 ;
  assign n53 = n52 ^ n49 ;
  assign n62 = n61 ^ n53 ;
  assign n83 = n82 ^ n62 ;
  assign n88 = n87 ^ n83 ;
  assign n93 = x0 & n88 ;
  assign n92 = x8 & ~n88 ;
  assign n94 = n93 ^ n92 ;
  assign n96 = n94 ^ x16 ;
  assign n98 = x1 & n88 ;
  assign n97 = x9 & ~n88 ;
  assign n99 = n98 ^ n97 ;
  assign n103 = n99 ^ x17 ;
  assign n104 = ~n96 & ~n103 ;
  assign n106 = x2 & n88 ;
  assign n105 = x10 & ~n88 ;
  assign n107 = n106 ^ n105 ;
  assign n109 = n107 ^ x18 ;
  assign n111 = x3 & n88 ;
  assign n110 = x11 & ~n88 ;
  assign n112 = n111 ^ n110 ;
  assign n118 = n112 ^ x19 ;
  assign n119 = ~n109 & ~n118 ;
  assign n120 = n104 & n119 ;
  assign n122 = x4 & n88 ;
  assign n121 = x12 & ~n88 ;
  assign n123 = n122 ^ n121 ;
  assign n125 = n123 ^ x20 ;
  assign n127 = x5 & n88 ;
  assign n126 = x13 & ~n88 ;
  assign n128 = n127 ^ n126 ;
  assign n132 = n128 ^ x21 ;
  assign n133 = ~n125 & ~n132 ;
  assign n135 = x6 & n88 ;
  assign n134 = x14 & ~n88 ;
  assign n136 = n135 ^ n134 ;
  assign n138 = n136 ^ x22 ;
  assign n149 = x7 & ~n62 ;
  assign n148 = x7 & ~n87 ;
  assign n150 = n149 ^ n148 ;
  assign n146 = x7 & n65 ;
  assign n147 = n81 & n146 ;
  assign n151 = n150 ^ n147 ;
  assign n142 = x15 & ~n62 ;
  assign n141 = x15 & ~n87 ;
  assign n143 = n142 ^ n141 ;
  assign n139 = x15 & n65 ;
  assign n140 = n81 & n139 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = n144 ^ x15 ;
  assign n152 = n151 ^ n145 ;
  assign n162 = n152 ^ x23 ;
  assign n163 = ~n138 & ~n162 ;
  assign n164 = n133 & n163 ;
  assign n165 = n120 & n164 ;
  assign n153 = x23 & n152 ;
  assign n154 = n153 ^ n152 ;
  assign n155 = n138 & n154 ;
  assign n156 = n155 ^ n154 ;
  assign n137 = ~x22 & n136 ;
  assign n157 = n156 ^ n137 ;
  assign n158 = n133 & n157 ;
  assign n129 = ~x21 & n128 ;
  assign n130 = ~n125 & n129 ;
  assign n124 = ~x20 & n123 ;
  assign n131 = n130 ^ n124 ;
  assign n159 = n158 ^ n131 ;
  assign n160 = n120 & n159 ;
  assign n113 = ~x19 & n112 ;
  assign n114 = ~n109 & n113 ;
  assign n108 = ~x18 & n107 ;
  assign n115 = n114 ^ n108 ;
  assign n116 = n104 & n115 ;
  assign n100 = ~x17 & n99 ;
  assign n101 = ~n96 & n100 ;
  assign n95 = ~x16 & n94 ;
  assign n102 = n101 ^ n95 ;
  assign n117 = n116 ^ n102 ;
  assign n161 = n160 ^ n117 ;
  assign n166 = n165 ^ n161 ;
  assign n263 = n94 & n166 ;
  assign n262 = x16 & ~n166 ;
  assign n264 = n263 ^ n262 ;
  assign n266 = n264 ^ x24 ;
  assign n268 = n99 & n166 ;
  assign n267 = x17 & ~n166 ;
  assign n269 = n268 ^ n267 ;
  assign n273 = n269 ^ x25 ;
  assign n274 = ~n266 & ~n273 ;
  assign n276 = n107 & n166 ;
  assign n275 = x18 & ~n166 ;
  assign n277 = n276 ^ n275 ;
  assign n279 = n277 ^ x26 ;
  assign n281 = n112 & n166 ;
  assign n280 = x19 & ~n166 ;
  assign n282 = n281 ^ n280 ;
  assign n288 = n282 ^ x27 ;
  assign n289 = ~n279 & ~n288 ;
  assign n290 = n274 & n289 ;
  assign n292 = n123 & n166 ;
  assign n291 = x20 & ~n166 ;
  assign n293 = n292 ^ n291 ;
  assign n295 = n293 ^ x28 ;
  assign n297 = n128 & n166 ;
  assign n296 = x21 & ~n166 ;
  assign n298 = n297 ^ n296 ;
  assign n302 = n298 ^ x29 ;
  assign n303 = ~n295 & ~n302 ;
  assign n317 = x22 & ~n166 ;
  assign n315 = n136 & n166 ;
  assign n330 = n317 ^ n315 ;
  assign n331 = n330 ^ x30 ;
  assign n249 = x23 & n166 ;
  assign n311 = n249 ^ x23 ;
  assign n247 = n152 & n166 ;
  assign n312 = n311 ^ n247 ;
  assign n332 = n312 ^ x31 ;
  assign n333 = ~n331 & ~n332 ;
  assign n334 = n303 & n333 ;
  assign n335 = n290 & n334 ;
  assign n322 = x22 & ~x30 ;
  assign n323 = ~n166 & n322 ;
  assign n308 = x23 & x31 ;
  assign n309 = ~n166 & n308 ;
  assign n306 = x31 & n152 ;
  assign n307 = n166 & n306 ;
  assign n310 = n309 ^ n307 ;
  assign n313 = n312 ^ n310 ;
  assign n318 = n313 & n317 ;
  assign n316 = n313 & n315 ;
  assign n319 = n318 ^ n316 ;
  assign n314 = x30 & n313 ;
  assign n320 = n319 ^ n314 ;
  assign n321 = n320 ^ n313 ;
  assign n324 = n323 ^ n321 ;
  assign n304 = ~x30 & n136 ;
  assign n305 = n166 & n304 ;
  assign n325 = n324 ^ n305 ;
  assign n326 = n303 & n325 ;
  assign n299 = ~x29 & n298 ;
  assign n300 = ~n295 & n299 ;
  assign n294 = ~x28 & n293 ;
  assign n301 = n300 ^ n294 ;
  assign n327 = n326 ^ n301 ;
  assign n328 = n290 & n327 ;
  assign n283 = ~x27 & n282 ;
  assign n284 = ~n279 & n283 ;
  assign n278 = ~x26 & n277 ;
  assign n285 = n284 ^ n278 ;
  assign n286 = n274 & n285 ;
  assign n270 = ~x25 & n269 ;
  assign n271 = ~n266 & n270 ;
  assign n265 = ~x24 & n264 ;
  assign n272 = n271 ^ n265 ;
  assign n287 = n286 ^ n272 ;
  assign n329 = n328 ^ n287 ;
  assign n336 = n335 ^ n329 ;
  assign n523 = n264 & n336 ;
  assign n522 = x24 & ~n336 ;
  assign n524 = n523 ^ n522 ;
  assign n526 = n524 ^ x32 ;
  assign n528 = n269 & n336 ;
  assign n527 = x25 & ~n336 ;
  assign n529 = n528 ^ n527 ;
  assign n533 = n529 ^ x33 ;
  assign n534 = ~n526 & ~n533 ;
  assign n536 = n277 & n336 ;
  assign n535 = x26 & ~n336 ;
  assign n537 = n536 ^ n535 ;
  assign n539 = n537 ^ x34 ;
  assign n541 = n282 & n336 ;
  assign n540 = x27 & ~n336 ;
  assign n542 = n541 ^ n540 ;
  assign n548 = n542 ^ x35 ;
  assign n549 = ~n539 & ~n548 ;
  assign n550 = n534 & n549 ;
  assign n552 = n293 & n336 ;
  assign n551 = x28 & ~n336 ;
  assign n553 = n552 ^ n551 ;
  assign n555 = n553 ^ x36 ;
  assign n557 = n298 & n336 ;
  assign n556 = x29 & ~n336 ;
  assign n558 = n557 ^ n556 ;
  assign n562 = n558 ^ x37 ;
  assign n563 = ~n555 & ~n562 ;
  assign n577 = x30 & ~n336 ;
  assign n575 = n330 & n336 ;
  assign n590 = n577 ^ n575 ;
  assign n591 = n590 ^ x38 ;
  assign n408 = x31 & n336 ;
  assign n571 = n408 ^ x31 ;
  assign n406 = n312 & n336 ;
  assign n572 = n571 ^ n406 ;
  assign n592 = n572 ^ x39 ;
  assign n593 = ~n591 & ~n592 ;
  assign n594 = n563 & n593 ;
  assign n595 = n550 & n594 ;
  assign n582 = x30 & ~x38 ;
  assign n583 = ~n336 & n582 ;
  assign n568 = x31 & x39 ;
  assign n569 = ~n336 & n568 ;
  assign n566 = x39 & n312 ;
  assign n567 = n336 & n566 ;
  assign n570 = n569 ^ n567 ;
  assign n573 = n572 ^ n570 ;
  assign n578 = n573 & n577 ;
  assign n576 = n573 & n575 ;
  assign n579 = n578 ^ n576 ;
  assign n574 = x38 & n573 ;
  assign n580 = n579 ^ n574 ;
  assign n581 = n580 ^ n573 ;
  assign n584 = n583 ^ n581 ;
  assign n564 = ~x38 & n330 ;
  assign n565 = n336 & n564 ;
  assign n585 = n584 ^ n565 ;
  assign n586 = n563 & n585 ;
  assign n559 = ~x37 & n558 ;
  assign n560 = ~n555 & n559 ;
  assign n554 = ~x36 & n553 ;
  assign n561 = n560 ^ n554 ;
  assign n587 = n586 ^ n561 ;
  assign n588 = n550 & n587 ;
  assign n543 = ~x35 & n542 ;
  assign n544 = ~n539 & n543 ;
  assign n538 = ~x34 & n537 ;
  assign n545 = n544 ^ n538 ;
  assign n546 = n534 & n545 ;
  assign n530 = ~x33 & n529 ;
  assign n531 = ~n526 & n530 ;
  assign n525 = ~x32 & n524 ;
  assign n532 = n531 ^ n525 ;
  assign n547 = n546 ^ n532 ;
  assign n589 = n588 ^ n547 ;
  assign n596 = n595 ^ n589 ;
  assign n871 = n524 & n596 ;
  assign n870 = x32 & ~n596 ;
  assign n872 = n871 ^ n870 ;
  assign n874 = n872 ^ x40 ;
  assign n876 = n529 & n596 ;
  assign n875 = x33 & ~n596 ;
  assign n877 = n876 ^ n875 ;
  assign n881 = n877 ^ x41 ;
  assign n882 = ~n874 & ~n881 ;
  assign n884 = n537 & n596 ;
  assign n883 = x34 & ~n596 ;
  assign n885 = n884 ^ n883 ;
  assign n887 = n885 ^ x42 ;
  assign n889 = n542 & n596 ;
  assign n888 = x35 & ~n596 ;
  assign n890 = n889 ^ n888 ;
  assign n896 = n890 ^ x43 ;
  assign n897 = ~n887 & ~n896 ;
  assign n898 = n882 & n897 ;
  assign n900 = n553 & n596 ;
  assign n899 = x36 & ~n596 ;
  assign n901 = n900 ^ n899 ;
  assign n903 = n901 ^ x44 ;
  assign n905 = n558 & n596 ;
  assign n904 = x37 & ~n596 ;
  assign n906 = n905 ^ n904 ;
  assign n910 = n906 ^ x45 ;
  assign n911 = ~n903 & ~n910 ;
  assign n925 = x38 & ~n596 ;
  assign n923 = n590 & n596 ;
  assign n938 = n925 ^ n923 ;
  assign n939 = n938 ^ x46 ;
  assign n666 = x39 & n596 ;
  assign n919 = n666 ^ x39 ;
  assign n664 = n572 & n596 ;
  assign n920 = n919 ^ n664 ;
  assign n940 = n920 ^ x47 ;
  assign n941 = ~n939 & ~n940 ;
  assign n942 = n911 & n941 ;
  assign n943 = n898 & n942 ;
  assign n930 = x38 & ~x46 ;
  assign n931 = ~n596 & n930 ;
  assign n916 = x39 & x47 ;
  assign n917 = ~n596 & n916 ;
  assign n914 = x47 & n572 ;
  assign n915 = n596 & n914 ;
  assign n918 = n917 ^ n915 ;
  assign n921 = n920 ^ n918 ;
  assign n926 = n921 & n925 ;
  assign n924 = n921 & n923 ;
  assign n927 = n926 ^ n924 ;
  assign n922 = x46 & n921 ;
  assign n928 = n927 ^ n922 ;
  assign n929 = n928 ^ n921 ;
  assign n932 = n931 ^ n929 ;
  assign n912 = ~x46 & n590 ;
  assign n913 = n596 & n912 ;
  assign n933 = n932 ^ n913 ;
  assign n934 = n911 & n933 ;
  assign n907 = ~x45 & n906 ;
  assign n908 = ~n903 & n907 ;
  assign n902 = ~x44 & n901 ;
  assign n909 = n908 ^ n902 ;
  assign n935 = n934 ^ n909 ;
  assign n936 = n898 & n935 ;
  assign n891 = ~x43 & n890 ;
  assign n892 = ~n887 & n891 ;
  assign n886 = ~x42 & n885 ;
  assign n893 = n892 ^ n886 ;
  assign n894 = n882 & n893 ;
  assign n878 = ~x41 & n877 ;
  assign n879 = ~n874 & n878 ;
  assign n873 = ~x40 & n872 ;
  assign n880 = n879 ^ n873 ;
  assign n895 = n894 ^ n880 ;
  assign n937 = n936 ^ n895 ;
  assign n944 = n943 ^ n937 ;
  assign n946 = x40 & n944 ;
  assign n945 = n872 & ~n944 ;
  assign n947 = n946 ^ n945 ;
  assign n90 = x8 & n88 ;
  assign n89 = x0 & ~n88 ;
  assign n91 = n90 ^ n89 ;
  assign n168 = x16 & n166 ;
  assign n167 = n94 & ~n166 ;
  assign n169 = n168 ^ n167 ;
  assign n171 = n169 ^ n91 ;
  assign n176 = x17 & n166 ;
  assign n175 = n99 & ~n166 ;
  assign n177 = n176 ^ n175 ;
  assign n173 = x9 & n88 ;
  assign n172 = x1 & ~n88 ;
  assign n174 = n173 ^ n172 ;
  assign n181 = n177 ^ n174 ;
  assign n182 = ~n171 & ~n181 ;
  assign n187 = x10 & n88 ;
  assign n186 = x2 & ~n88 ;
  assign n188 = n187 ^ n186 ;
  assign n184 = x18 & n166 ;
  assign n183 = n107 & ~n166 ;
  assign n185 = n184 ^ n183 ;
  assign n190 = n188 ^ n185 ;
  assign n195 = x11 & n88 ;
  assign n194 = x3 & ~n88 ;
  assign n196 = n195 ^ n194 ;
  assign n192 = x19 & n166 ;
  assign n191 = n112 & ~n166 ;
  assign n193 = n192 ^ n191 ;
  assign n202 = n196 ^ n193 ;
  assign n203 = ~n190 & ~n202 ;
  assign n204 = n182 & n203 ;
  assign n209 = x12 & n88 ;
  assign n208 = x4 & ~n88 ;
  assign n210 = n209 ^ n208 ;
  assign n206 = x20 & n166 ;
  assign n205 = n123 & ~n166 ;
  assign n207 = n206 ^ n205 ;
  assign n212 = n210 ^ n207 ;
  assign n217 = x13 & n88 ;
  assign n216 = x5 & ~n88 ;
  assign n218 = n217 ^ n216 ;
  assign n214 = x21 & n166 ;
  assign n213 = n128 & ~n166 ;
  assign n215 = n214 ^ n213 ;
  assign n222 = n218 ^ n215 ;
  assign n223 = ~n212 & ~n222 ;
  assign n228 = x14 & n88 ;
  assign n227 = x6 & ~n88 ;
  assign n229 = n228 ^ n227 ;
  assign n225 = x22 & n166 ;
  assign n224 = n136 & ~n166 ;
  assign n226 = n225 ^ n224 ;
  assign n231 = n229 ^ n226 ;
  assign n248 = n247 ^ n152 ;
  assign n250 = n249 ^ n248 ;
  assign n232 = x7 & ~n88 ;
  assign n233 = n232 ^ n144 ;
  assign n251 = n250 ^ n233 ;
  assign n252 = ~n231 & ~n251 ;
  assign n253 = n223 & n252 ;
  assign n254 = n204 & n253 ;
  assign n236 = x23 & n233 ;
  assign n237 = n166 & n236 ;
  assign n234 = n152 & n233 ;
  assign n235 = ~n166 & n234 ;
  assign n238 = n237 ^ n235 ;
  assign n239 = n238 ^ n233 ;
  assign n240 = n231 & n239 ;
  assign n241 = n240 ^ n239 ;
  assign n230 = ~n226 & n229 ;
  assign n242 = n241 ^ n230 ;
  assign n243 = n223 & n242 ;
  assign n219 = ~n215 & n218 ;
  assign n220 = ~n212 & n219 ;
  assign n211 = ~n207 & n210 ;
  assign n221 = n220 ^ n211 ;
  assign n244 = n243 ^ n221 ;
  assign n245 = n204 & n244 ;
  assign n197 = ~n193 & n196 ;
  assign n198 = ~n190 & n197 ;
  assign n189 = ~n185 & n188 ;
  assign n199 = n198 ^ n189 ;
  assign n200 = n182 & n199 ;
  assign n178 = n174 & ~n177 ;
  assign n179 = ~n171 & n178 ;
  assign n170 = n91 & ~n169 ;
  assign n180 = n179 ^ n170 ;
  assign n201 = n200 ^ n180 ;
  assign n246 = n245 ^ n201 ;
  assign n255 = n254 ^ n246 ;
  assign n260 = n91 & n255 ;
  assign n259 = n169 & ~n255 ;
  assign n261 = n260 ^ n259 ;
  assign n338 = x24 & n336 ;
  assign n337 = n264 & ~n336 ;
  assign n339 = n338 ^ n337 ;
  assign n341 = n339 ^ n261 ;
  assign n346 = x25 & n336 ;
  assign n345 = n269 & ~n336 ;
  assign n347 = n346 ^ n345 ;
  assign n343 = n174 & n255 ;
  assign n342 = n177 & ~n255 ;
  assign n344 = n343 ^ n342 ;
  assign n351 = n347 ^ n344 ;
  assign n352 = ~n341 & ~n351 ;
  assign n357 = n188 & n255 ;
  assign n356 = n185 & ~n255 ;
  assign n358 = n357 ^ n356 ;
  assign n354 = x26 & n336 ;
  assign n353 = n277 & ~n336 ;
  assign n355 = n354 ^ n353 ;
  assign n360 = n358 ^ n355 ;
  assign n365 = n196 & n255 ;
  assign n364 = n193 & ~n255 ;
  assign n366 = n365 ^ n364 ;
  assign n362 = x27 & n336 ;
  assign n361 = n282 & ~n336 ;
  assign n363 = n362 ^ n361 ;
  assign n372 = n366 ^ n363 ;
  assign n373 = ~n360 & ~n372 ;
  assign n374 = n352 & n373 ;
  assign n379 = n210 & n255 ;
  assign n378 = n207 & ~n255 ;
  assign n380 = n379 ^ n378 ;
  assign n376 = x28 & n336 ;
  assign n375 = n293 & ~n336 ;
  assign n377 = n376 ^ n375 ;
  assign n382 = n380 ^ n377 ;
  assign n387 = n218 & n255 ;
  assign n386 = n215 & ~n255 ;
  assign n388 = n387 ^ n386 ;
  assign n384 = x29 & n336 ;
  assign n383 = n298 & ~n336 ;
  assign n385 = n384 ^ n383 ;
  assign n392 = n388 ^ n385 ;
  assign n393 = ~n382 & ~n392 ;
  assign n398 = n229 & n255 ;
  assign n397 = n226 & ~n255 ;
  assign n399 = n398 ^ n397 ;
  assign n395 = x30 & n336 ;
  assign n394 = n330 & ~n336 ;
  assign n396 = n395 ^ n394 ;
  assign n401 = n399 ^ n396 ;
  assign n407 = n406 ^ n312 ;
  assign n409 = n408 ^ n407 ;
  assign n404 = n233 & n255 ;
  assign n402 = n250 & n255 ;
  assign n403 = n402 ^ n250 ;
  assign n405 = n404 ^ n403 ;
  assign n419 = n409 ^ n405 ;
  assign n420 = ~n401 & ~n419 ;
  assign n421 = n393 & n420 ;
  assign n422 = n374 & n421 ;
  assign n410 = n405 & n409 ;
  assign n411 = n410 ^ n405 ;
  assign n412 = n401 & n411 ;
  assign n413 = n412 ^ n411 ;
  assign n400 = ~n396 & n399 ;
  assign n414 = n413 ^ n400 ;
  assign n415 = n393 & n414 ;
  assign n389 = ~n385 & n388 ;
  assign n390 = ~n382 & n389 ;
  assign n381 = ~n377 & n380 ;
  assign n391 = n390 ^ n381 ;
  assign n416 = n415 ^ n391 ;
  assign n417 = n374 & n416 ;
  assign n367 = ~n363 & n366 ;
  assign n368 = ~n360 & n367 ;
  assign n359 = ~n355 & n358 ;
  assign n369 = n368 ^ n359 ;
  assign n370 = n352 & n369 ;
  assign n348 = n344 & ~n347 ;
  assign n349 = ~n341 & n348 ;
  assign n340 = n261 & ~n339 ;
  assign n350 = n349 ^ n340 ;
  assign n371 = n370 ^ n350 ;
  assign n418 = n417 ^ n371 ;
  assign n423 = n422 ^ n418 ;
  assign n520 = n261 & n423 ;
  assign n519 = n339 & ~n423 ;
  assign n521 = n520 ^ n519 ;
  assign n598 = x32 & n596 ;
  assign n597 = n524 & ~n596 ;
  assign n599 = n598 ^ n597 ;
  assign n601 = n599 ^ n521 ;
  assign n606 = x33 & n596 ;
  assign n605 = n529 & ~n596 ;
  assign n607 = n606 ^ n605 ;
  assign n603 = n344 & n423 ;
  assign n602 = n347 & ~n423 ;
  assign n604 = n603 ^ n602 ;
  assign n611 = n607 ^ n604 ;
  assign n612 = ~n601 & ~n611 ;
  assign n617 = n358 & n423 ;
  assign n616 = n355 & ~n423 ;
  assign n618 = n617 ^ n616 ;
  assign n614 = x34 & n596 ;
  assign n613 = n537 & ~n596 ;
  assign n615 = n614 ^ n613 ;
  assign n620 = n618 ^ n615 ;
  assign n625 = n366 & n423 ;
  assign n624 = n363 & ~n423 ;
  assign n626 = n625 ^ n624 ;
  assign n622 = x35 & n596 ;
  assign n621 = n542 & ~n596 ;
  assign n623 = n622 ^ n621 ;
  assign n632 = n626 ^ n623 ;
  assign n633 = ~n620 & ~n632 ;
  assign n634 = n612 & n633 ;
  assign n639 = n380 & n423 ;
  assign n638 = n377 & ~n423 ;
  assign n640 = n639 ^ n638 ;
  assign n636 = x36 & n596 ;
  assign n635 = n553 & ~n596 ;
  assign n637 = n636 ^ n635 ;
  assign n642 = n640 ^ n637 ;
  assign n647 = n388 & n423 ;
  assign n646 = n385 & ~n423 ;
  assign n648 = n647 ^ n646 ;
  assign n644 = x37 & n596 ;
  assign n643 = n558 & ~n596 ;
  assign n645 = n644 ^ n643 ;
  assign n652 = n648 ^ n645 ;
  assign n653 = ~n642 & ~n652 ;
  assign n658 = n399 & n423 ;
  assign n657 = n396 & ~n423 ;
  assign n659 = n658 ^ n657 ;
  assign n655 = x38 & n596 ;
  assign n654 = n590 & ~n596 ;
  assign n656 = n655 ^ n654 ;
  assign n661 = n659 ^ n656 ;
  assign n665 = n664 ^ n572 ;
  assign n667 = n666 ^ n665 ;
  assign n506 = n409 & n423 ;
  assign n662 = n506 ^ n409 ;
  assign n504 = n405 & n423 ;
  assign n663 = n662 ^ n504 ;
  assign n677 = n667 ^ n663 ;
  assign n678 = ~n661 & ~n677 ;
  assign n679 = n653 & n678 ;
  assign n680 = n634 & n679 ;
  assign n668 = n663 & n667 ;
  assign n669 = n668 ^ n663 ;
  assign n670 = n661 & n669 ;
  assign n671 = n670 ^ n669 ;
  assign n660 = ~n656 & n659 ;
  assign n672 = n671 ^ n660 ;
  assign n673 = n653 & n672 ;
  assign n649 = ~n645 & n648 ;
  assign n650 = ~n642 & n649 ;
  assign n641 = ~n637 & n640 ;
  assign n651 = n650 ^ n641 ;
  assign n674 = n673 ^ n651 ;
  assign n675 = n634 & n674 ;
  assign n627 = ~n623 & n626 ;
  assign n628 = ~n620 & n627 ;
  assign n619 = ~n615 & n618 ;
  assign n629 = n628 ^ n619 ;
  assign n630 = n612 & n629 ;
  assign n608 = n604 & ~n607 ;
  assign n609 = ~n601 & n608 ;
  assign n600 = n521 & ~n599 ;
  assign n610 = n609 ^ n600 ;
  assign n631 = n630 ^ n610 ;
  assign n676 = n675 ^ n631 ;
  assign n681 = n680 ^ n676 ;
  assign n868 = n521 & n681 ;
  assign n867 = n599 & ~n681 ;
  assign n869 = n868 ^ n867 ;
  assign n949 = n947 ^ n869 ;
  assign n954 = n604 & n681 ;
  assign n953 = n607 & ~n681 ;
  assign n955 = n954 ^ n953 ;
  assign n951 = x41 & n944 ;
  assign n950 = n877 & ~n944 ;
  assign n952 = n951 ^ n950 ;
  assign n959 = n955 ^ n952 ;
  assign n960 = ~n949 & ~n959 ;
  assign n965 = n618 & n681 ;
  assign n964 = n615 & ~n681 ;
  assign n966 = n965 ^ n964 ;
  assign n962 = x42 & n944 ;
  assign n961 = n885 & ~n944 ;
  assign n963 = n962 ^ n961 ;
  assign n968 = n966 ^ n963 ;
  assign n973 = n626 & n681 ;
  assign n972 = n623 & ~n681 ;
  assign n974 = n973 ^ n972 ;
  assign n970 = x43 & n944 ;
  assign n969 = n890 & ~n944 ;
  assign n971 = n970 ^ n969 ;
  assign n980 = n974 ^ n971 ;
  assign n981 = ~n968 & ~n980 ;
  assign n982 = n960 & n981 ;
  assign n987 = n640 & n681 ;
  assign n986 = n637 & ~n681 ;
  assign n988 = n987 ^ n986 ;
  assign n984 = x44 & n944 ;
  assign n983 = n901 & ~n944 ;
  assign n985 = n984 ^ n983 ;
  assign n990 = n988 ^ n985 ;
  assign n995 = n648 & n681 ;
  assign n994 = n645 & ~n681 ;
  assign n996 = n995 ^ n994 ;
  assign n992 = x45 & n944 ;
  assign n991 = n906 & ~n944 ;
  assign n993 = n992 ^ n991 ;
  assign n1000 = n996 ^ n993 ;
  assign n1001 = ~n990 & ~n1000 ;
  assign n1006 = n659 & n681 ;
  assign n1005 = n656 & ~n681 ;
  assign n1007 = n1006 ^ n1005 ;
  assign n1003 = x46 & n944 ;
  assign n1002 = n938 & ~n944 ;
  assign n1004 = n1003 ^ n1002 ;
  assign n1009 = n1007 ^ n1004 ;
  assign n753 = n667 & n681 ;
  assign n1014 = n753 ^ n667 ;
  assign n751 = n663 & n681 ;
  assign n1015 = n1014 ^ n751 ;
  assign n1012 = x47 & n944 ;
  assign n1010 = n920 & n944 ;
  assign n1011 = n1010 ^ n920 ;
  assign n1013 = n1012 ^ n1011 ;
  assign n1025 = n1015 ^ n1013 ;
  assign n1026 = ~n1009 & ~n1025 ;
  assign n1027 = n1001 & n1026 ;
  assign n1028 = n982 & n1027 ;
  assign n1016 = n1013 & n1015 ;
  assign n1017 = n1016 ^ n1015 ;
  assign n1018 = n1009 & n1017 ;
  assign n1019 = n1018 ^ n1017 ;
  assign n1008 = ~n1004 & n1007 ;
  assign n1020 = n1019 ^ n1008 ;
  assign n1021 = n1001 & n1020 ;
  assign n997 = ~n993 & n996 ;
  assign n998 = ~n990 & n997 ;
  assign n989 = ~n985 & n988 ;
  assign n999 = n998 ^ n989 ;
  assign n1022 = n1021 ^ n999 ;
  assign n1023 = n982 & n1022 ;
  assign n975 = ~n971 & n974 ;
  assign n976 = ~n968 & n975 ;
  assign n967 = ~n963 & n966 ;
  assign n977 = n976 ^ n967 ;
  assign n978 = n960 & n977 ;
  assign n956 = ~n952 & n955 ;
  assign n957 = ~n949 & n956 ;
  assign n948 = n869 & ~n947 ;
  assign n958 = n957 ^ n948 ;
  assign n979 = n978 ^ n958 ;
  assign n1024 = n1023 ^ n979 ;
  assign n1029 = n1028 ^ n1024 ;
  assign n1031 = n947 & n1029 ;
  assign n1030 = n869 & ~n1029 ;
  assign n1032 = n1031 ^ n1030 ;
  assign n257 = n169 & n255 ;
  assign n256 = n91 & ~n255 ;
  assign n258 = n257 ^ n256 ;
  assign n425 = n339 & n423 ;
  assign n424 = n261 & ~n423 ;
  assign n426 = n425 ^ n424 ;
  assign n428 = n426 ^ n258 ;
  assign n433 = n347 & n423 ;
  assign n432 = n344 & ~n423 ;
  assign n434 = n433 ^ n432 ;
  assign n430 = n177 & n255 ;
  assign n429 = n174 & ~n255 ;
  assign n431 = n430 ^ n429 ;
  assign n438 = n434 ^ n431 ;
  assign n439 = ~n428 & ~n438 ;
  assign n444 = n185 & n255 ;
  assign n443 = n188 & ~n255 ;
  assign n445 = n444 ^ n443 ;
  assign n441 = n355 & n423 ;
  assign n440 = n358 & ~n423 ;
  assign n442 = n441 ^ n440 ;
  assign n447 = n445 ^ n442 ;
  assign n452 = n193 & n255 ;
  assign n451 = n196 & ~n255 ;
  assign n453 = n452 ^ n451 ;
  assign n449 = n363 & n423 ;
  assign n448 = n366 & ~n423 ;
  assign n450 = n449 ^ n448 ;
  assign n459 = n453 ^ n450 ;
  assign n460 = ~n447 & ~n459 ;
  assign n461 = n439 & n460 ;
  assign n466 = n207 & n255 ;
  assign n465 = n210 & ~n255 ;
  assign n467 = n466 ^ n465 ;
  assign n463 = n377 & n423 ;
  assign n462 = n380 & ~n423 ;
  assign n464 = n463 ^ n462 ;
  assign n469 = n467 ^ n464 ;
  assign n474 = n215 & n255 ;
  assign n473 = n218 & ~n255 ;
  assign n475 = n474 ^ n473 ;
  assign n471 = n385 & n423 ;
  assign n470 = n388 & ~n423 ;
  assign n472 = n471 ^ n470 ;
  assign n479 = n475 ^ n472 ;
  assign n480 = ~n469 & ~n479 ;
  assign n485 = n226 & n255 ;
  assign n484 = n229 & ~n255 ;
  assign n486 = n485 ^ n484 ;
  assign n482 = n396 & n423 ;
  assign n481 = n399 & ~n423 ;
  assign n483 = n482 ^ n481 ;
  assign n488 = n486 ^ n483 ;
  assign n505 = n504 ^ n405 ;
  assign n507 = n506 ^ n505 ;
  assign n489 = n233 & ~n255 ;
  assign n490 = n489 ^ n402 ;
  assign n508 = n507 ^ n490 ;
  assign n509 = ~n488 & ~n508 ;
  assign n510 = n480 & n509 ;
  assign n511 = n461 & n510 ;
  assign n493 = n409 & n490 ;
  assign n494 = n423 & n493 ;
  assign n491 = n405 & n490 ;
  assign n492 = ~n423 & n491 ;
  assign n495 = n494 ^ n492 ;
  assign n496 = n495 ^ n490 ;
  assign n497 = n488 & n496 ;
  assign n498 = n497 ^ n496 ;
  assign n487 = ~n483 & n486 ;
  assign n499 = n498 ^ n487 ;
  assign n500 = n480 & n499 ;
  assign n476 = ~n472 & n475 ;
  assign n477 = ~n469 & n476 ;
  assign n468 = ~n464 & n467 ;
  assign n478 = n477 ^ n468 ;
  assign n501 = n500 ^ n478 ;
  assign n502 = n461 & n501 ;
  assign n454 = ~n450 & n453 ;
  assign n455 = ~n447 & n454 ;
  assign n446 = ~n442 & n445 ;
  assign n456 = n455 ^ n446 ;
  assign n457 = n439 & n456 ;
  assign n435 = n431 & ~n434 ;
  assign n436 = ~n428 & n435 ;
  assign n427 = n258 & ~n426 ;
  assign n437 = n436 ^ n427 ;
  assign n458 = n457 ^ n437 ;
  assign n503 = n502 ^ n458 ;
  assign n512 = n511 ^ n503 ;
  assign n517 = n258 & n512 ;
  assign n516 = n426 & ~n512 ;
  assign n518 = n517 ^ n516 ;
  assign n683 = n599 & n681 ;
  assign n682 = n521 & ~n681 ;
  assign n684 = n683 ^ n682 ;
  assign n686 = n684 ^ n518 ;
  assign n691 = n607 & n681 ;
  assign n690 = n604 & ~n681 ;
  assign n692 = n691 ^ n690 ;
  assign n688 = n431 & n512 ;
  assign n687 = n434 & ~n512 ;
  assign n689 = n688 ^ n687 ;
  assign n696 = n692 ^ n689 ;
  assign n697 = ~n686 & ~n696 ;
  assign n702 = n445 & n512 ;
  assign n701 = n442 & ~n512 ;
  assign n703 = n702 ^ n701 ;
  assign n699 = n615 & n681 ;
  assign n698 = n618 & ~n681 ;
  assign n700 = n699 ^ n698 ;
  assign n705 = n703 ^ n700 ;
  assign n710 = n453 & n512 ;
  assign n709 = n450 & ~n512 ;
  assign n711 = n710 ^ n709 ;
  assign n707 = n623 & n681 ;
  assign n706 = n626 & ~n681 ;
  assign n708 = n707 ^ n706 ;
  assign n717 = n711 ^ n708 ;
  assign n718 = ~n705 & ~n717 ;
  assign n719 = n697 & n718 ;
  assign n724 = n467 & n512 ;
  assign n723 = n464 & ~n512 ;
  assign n725 = n724 ^ n723 ;
  assign n721 = n637 & n681 ;
  assign n720 = n640 & ~n681 ;
  assign n722 = n721 ^ n720 ;
  assign n727 = n725 ^ n722 ;
  assign n732 = n475 & n512 ;
  assign n731 = n472 & ~n512 ;
  assign n733 = n732 ^ n731 ;
  assign n729 = n645 & n681 ;
  assign n728 = n648 & ~n681 ;
  assign n730 = n729 ^ n728 ;
  assign n737 = n733 ^ n730 ;
  assign n738 = ~n727 & ~n737 ;
  assign n743 = n486 & n512 ;
  assign n742 = n483 & ~n512 ;
  assign n744 = n743 ^ n742 ;
  assign n740 = n656 & n681 ;
  assign n739 = n659 & ~n681 ;
  assign n741 = n740 ^ n739 ;
  assign n746 = n744 ^ n741 ;
  assign n752 = n751 ^ n663 ;
  assign n754 = n753 ^ n752 ;
  assign n749 = n490 & n512 ;
  assign n747 = n507 & n512 ;
  assign n748 = n747 ^ n507 ;
  assign n750 = n749 ^ n748 ;
  assign n764 = n754 ^ n750 ;
  assign n765 = ~n746 & ~n764 ;
  assign n766 = n738 & n765 ;
  assign n767 = n719 & n766 ;
  assign n755 = n750 & n754 ;
  assign n756 = n755 ^ n750 ;
  assign n757 = n746 & n756 ;
  assign n758 = n757 ^ n756 ;
  assign n745 = ~n741 & n744 ;
  assign n759 = n758 ^ n745 ;
  assign n760 = n738 & n759 ;
  assign n734 = ~n730 & n733 ;
  assign n735 = ~n727 & n734 ;
  assign n726 = ~n722 & n725 ;
  assign n736 = n735 ^ n726 ;
  assign n761 = n760 ^ n736 ;
  assign n762 = n719 & n761 ;
  assign n712 = ~n708 & n711 ;
  assign n713 = ~n705 & n712 ;
  assign n704 = ~n700 & n703 ;
  assign n714 = n713 ^ n704 ;
  assign n715 = n697 & n714 ;
  assign n693 = n689 & ~n692 ;
  assign n694 = ~n686 & n693 ;
  assign n685 = n518 & ~n684 ;
  assign n695 = n694 ^ n685 ;
  assign n716 = n715 ^ n695 ;
  assign n763 = n762 ^ n716 ;
  assign n768 = n767 ^ n763 ;
  assign n865 = n518 & n768 ;
  assign n864 = n684 & ~n768 ;
  assign n866 = n865 ^ n864 ;
  assign n1034 = n1032 ^ n866 ;
  assign n1039 = n689 & n768 ;
  assign n1038 = n692 & ~n768 ;
  assign n1040 = n1039 ^ n1038 ;
  assign n1036 = n952 & n1029 ;
  assign n1035 = n955 & ~n1029 ;
  assign n1037 = n1036 ^ n1035 ;
  assign n1044 = n1040 ^ n1037 ;
  assign n1045 = ~n1034 & ~n1044 ;
  assign n1050 = n703 & n768 ;
  assign n1049 = n700 & ~n768 ;
  assign n1051 = n1050 ^ n1049 ;
  assign n1047 = n963 & n1029 ;
  assign n1046 = n966 & ~n1029 ;
  assign n1048 = n1047 ^ n1046 ;
  assign n1053 = n1051 ^ n1048 ;
  assign n1058 = n711 & n768 ;
  assign n1057 = n708 & ~n768 ;
  assign n1059 = n1058 ^ n1057 ;
  assign n1055 = n971 & n1029 ;
  assign n1054 = n974 & ~n1029 ;
  assign n1056 = n1055 ^ n1054 ;
  assign n1065 = n1059 ^ n1056 ;
  assign n1066 = ~n1053 & ~n1065 ;
  assign n1067 = n1045 & n1066 ;
  assign n1072 = n725 & n768 ;
  assign n1071 = n722 & ~n768 ;
  assign n1073 = n1072 ^ n1071 ;
  assign n1069 = n985 & n1029 ;
  assign n1068 = n988 & ~n1029 ;
  assign n1070 = n1069 ^ n1068 ;
  assign n1075 = n1073 ^ n1070 ;
  assign n1080 = n733 & n768 ;
  assign n1079 = n730 & ~n768 ;
  assign n1081 = n1080 ^ n1079 ;
  assign n1077 = n993 & n1029 ;
  assign n1076 = n996 & ~n1029 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1085 = n1081 ^ n1078 ;
  assign n1086 = ~n1075 & ~n1085 ;
  assign n1091 = n744 & n768 ;
  assign n1090 = n741 & ~n768 ;
  assign n1092 = n1091 ^ n1090 ;
  assign n1088 = n1004 & n1029 ;
  assign n1087 = n1007 & ~n1029 ;
  assign n1089 = n1088 ^ n1087 ;
  assign n1094 = n1092 ^ n1089 ;
  assign n851 = n754 & n768 ;
  assign n1099 = n851 ^ n754 ;
  assign n849 = n750 & n768 ;
  assign n1100 = n1099 ^ n849 ;
  assign n1097 = n1013 & n1029 ;
  assign n1095 = n1015 & n1029 ;
  assign n1096 = n1095 ^ n1015 ;
  assign n1098 = n1097 ^ n1096 ;
  assign n1110 = n1100 ^ n1098 ;
  assign n1111 = ~n1094 & ~n1110 ;
  assign n1112 = n1086 & n1111 ;
  assign n1113 = n1067 & n1112 ;
  assign n1101 = n1098 & n1100 ;
  assign n1102 = n1101 ^ n1100 ;
  assign n1103 = n1094 & n1102 ;
  assign n1104 = n1103 ^ n1102 ;
  assign n1093 = ~n1089 & n1092 ;
  assign n1105 = n1104 ^ n1093 ;
  assign n1106 = n1086 & n1105 ;
  assign n1082 = ~n1078 & n1081 ;
  assign n1083 = ~n1075 & n1082 ;
  assign n1074 = ~n1070 & n1073 ;
  assign n1084 = n1083 ^ n1074 ;
  assign n1107 = n1106 ^ n1084 ;
  assign n1108 = n1067 & n1107 ;
  assign n1060 = ~n1056 & n1059 ;
  assign n1061 = ~n1053 & n1060 ;
  assign n1052 = ~n1048 & n1051 ;
  assign n1062 = n1061 ^ n1052 ;
  assign n1063 = n1045 & n1062 ;
  assign n1041 = ~n1037 & n1040 ;
  assign n1042 = ~n1034 & n1041 ;
  assign n1033 = n866 & ~n1032 ;
  assign n1043 = n1042 ^ n1033 ;
  assign n1064 = n1063 ^ n1043 ;
  assign n1109 = n1108 ^ n1064 ;
  assign n1114 = n1113 ^ n1109 ;
  assign n1116 = n1032 & n1114 ;
  assign n1115 = n866 & ~n1114 ;
  assign n1117 = n1116 ^ n1115 ;
  assign n514 = n426 & n512 ;
  assign n513 = n258 & ~n512 ;
  assign n515 = n514 ^ n513 ;
  assign n770 = n684 & n768 ;
  assign n769 = n518 & ~n768 ;
  assign n771 = n770 ^ n769 ;
  assign n773 = n771 ^ n515 ;
  assign n778 = n692 & n768 ;
  assign n777 = n689 & ~n768 ;
  assign n779 = n778 ^ n777 ;
  assign n775 = n434 & n512 ;
  assign n774 = n431 & ~n512 ;
  assign n776 = n775 ^ n774 ;
  assign n783 = n779 ^ n776 ;
  assign n784 = ~n773 & ~n783 ;
  assign n789 = n442 & n512 ;
  assign n788 = n445 & ~n512 ;
  assign n790 = n789 ^ n788 ;
  assign n786 = n700 & n768 ;
  assign n785 = n703 & ~n768 ;
  assign n787 = n786 ^ n785 ;
  assign n792 = n790 ^ n787 ;
  assign n797 = n450 & n512 ;
  assign n796 = n453 & ~n512 ;
  assign n798 = n797 ^ n796 ;
  assign n794 = n708 & n768 ;
  assign n793 = n711 & ~n768 ;
  assign n795 = n794 ^ n793 ;
  assign n804 = n798 ^ n795 ;
  assign n805 = ~n792 & ~n804 ;
  assign n806 = n784 & n805 ;
  assign n811 = n464 & n512 ;
  assign n810 = n467 & ~n512 ;
  assign n812 = n811 ^ n810 ;
  assign n808 = n722 & n768 ;
  assign n807 = n725 & ~n768 ;
  assign n809 = n808 ^ n807 ;
  assign n814 = n812 ^ n809 ;
  assign n819 = n472 & n512 ;
  assign n818 = n475 & ~n512 ;
  assign n820 = n819 ^ n818 ;
  assign n816 = n730 & n768 ;
  assign n815 = n733 & ~n768 ;
  assign n817 = n816 ^ n815 ;
  assign n824 = n820 ^ n817 ;
  assign n825 = ~n814 & ~n824 ;
  assign n830 = n483 & n512 ;
  assign n829 = n486 & ~n512 ;
  assign n831 = n830 ^ n829 ;
  assign n827 = n741 & n768 ;
  assign n826 = n744 & ~n768 ;
  assign n828 = n827 ^ n826 ;
  assign n833 = n831 ^ n828 ;
  assign n850 = n849 ^ n750 ;
  assign n852 = n851 ^ n850 ;
  assign n834 = n490 & ~n512 ;
  assign n835 = n834 ^ n747 ;
  assign n853 = n852 ^ n835 ;
  assign n854 = ~n833 & ~n853 ;
  assign n855 = n825 & n854 ;
  assign n856 = n806 & n855 ;
  assign n838 = n754 & n835 ;
  assign n839 = n768 & n838 ;
  assign n836 = n750 & n835 ;
  assign n837 = ~n768 & n836 ;
  assign n840 = n839 ^ n837 ;
  assign n841 = n840 ^ n835 ;
  assign n842 = n833 & n841 ;
  assign n843 = n842 ^ n841 ;
  assign n832 = ~n828 & n831 ;
  assign n844 = n843 ^ n832 ;
  assign n845 = n825 & n844 ;
  assign n821 = ~n817 & n820 ;
  assign n822 = ~n814 & n821 ;
  assign n813 = ~n809 & n812 ;
  assign n823 = n822 ^ n813 ;
  assign n846 = n845 ^ n823 ;
  assign n847 = n806 & n846 ;
  assign n799 = ~n795 & n798 ;
  assign n800 = ~n792 & n799 ;
  assign n791 = ~n787 & n790 ;
  assign n801 = n800 ^ n791 ;
  assign n802 = n784 & n801 ;
  assign n780 = n776 & ~n779 ;
  assign n781 = ~n773 & n780 ;
  assign n772 = n515 & ~n771 ;
  assign n782 = n781 ^ n772 ;
  assign n803 = n802 ^ n782 ;
  assign n848 = n847 ^ n803 ;
  assign n857 = n856 ^ n848 ;
  assign n862 = n515 & n857 ;
  assign n861 = n771 & ~n857 ;
  assign n863 = n862 ^ n861 ;
  assign n1119 = n1117 ^ n863 ;
  assign n1124 = n776 & n857 ;
  assign n1123 = n779 & ~n857 ;
  assign n1125 = n1124 ^ n1123 ;
  assign n1121 = n1037 & n1114 ;
  assign n1120 = n1040 & ~n1114 ;
  assign n1122 = n1121 ^ n1120 ;
  assign n1129 = n1125 ^ n1122 ;
  assign n1130 = ~n1119 & ~n1129 ;
  assign n1135 = n790 & n857 ;
  assign n1134 = n787 & ~n857 ;
  assign n1136 = n1135 ^ n1134 ;
  assign n1132 = n1048 & n1114 ;
  assign n1131 = n1051 & ~n1114 ;
  assign n1133 = n1132 ^ n1131 ;
  assign n1138 = n1136 ^ n1133 ;
  assign n1143 = n798 & n857 ;
  assign n1142 = n795 & ~n857 ;
  assign n1144 = n1143 ^ n1142 ;
  assign n1140 = n1056 & n1114 ;
  assign n1139 = n1059 & ~n1114 ;
  assign n1141 = n1140 ^ n1139 ;
  assign n1150 = n1144 ^ n1141 ;
  assign n1151 = ~n1138 & ~n1150 ;
  assign n1152 = n1130 & n1151 ;
  assign n1157 = n812 & n857 ;
  assign n1156 = n809 & ~n857 ;
  assign n1158 = n1157 ^ n1156 ;
  assign n1154 = n1070 & n1114 ;
  assign n1153 = n1073 & ~n1114 ;
  assign n1155 = n1154 ^ n1153 ;
  assign n1160 = n1158 ^ n1155 ;
  assign n1165 = n820 & n857 ;
  assign n1164 = n817 & ~n857 ;
  assign n1166 = n1165 ^ n1164 ;
  assign n1162 = n1078 & n1114 ;
  assign n1161 = n1081 & ~n1114 ;
  assign n1163 = n1162 ^ n1161 ;
  assign n1170 = n1166 ^ n1163 ;
  assign n1171 = ~n1160 & ~n1170 ;
  assign n1176 = n831 & n857 ;
  assign n1175 = n828 & ~n857 ;
  assign n1177 = n1176 ^ n1175 ;
  assign n1173 = n1089 & n1114 ;
  assign n1172 = n1092 & ~n1114 ;
  assign n1174 = n1173 ^ n1172 ;
  assign n1179 = n1177 ^ n1174 ;
  assign n1186 = n835 & n857 ;
  assign n1184 = n852 & n857 ;
  assign n1185 = n1184 ^ n852 ;
  assign n1187 = n1186 ^ n1185 ;
  assign n1182 = n1098 & n1114 ;
  assign n1180 = n1100 & n1114 ;
  assign n1181 = n1180 ^ n1100 ;
  assign n1183 = n1182 ^ n1181 ;
  assign n1197 = n1187 ^ n1183 ;
  assign n1198 = ~n1179 & ~n1197 ;
  assign n1199 = n1171 & n1198 ;
  assign n1200 = n1152 & n1199 ;
  assign n1188 = n1183 & n1187 ;
  assign n1189 = n1188 ^ n1187 ;
  assign n1190 = n1179 & n1189 ;
  assign n1191 = n1190 ^ n1189 ;
  assign n1178 = ~n1174 & n1177 ;
  assign n1192 = n1191 ^ n1178 ;
  assign n1193 = n1171 & n1192 ;
  assign n1167 = ~n1163 & n1166 ;
  assign n1168 = ~n1160 & n1167 ;
  assign n1159 = ~n1155 & n1158 ;
  assign n1169 = n1168 ^ n1159 ;
  assign n1194 = n1193 ^ n1169 ;
  assign n1195 = n1152 & n1194 ;
  assign n1145 = ~n1141 & n1144 ;
  assign n1146 = ~n1138 & n1145 ;
  assign n1137 = ~n1133 & n1136 ;
  assign n1147 = n1146 ^ n1137 ;
  assign n1148 = n1130 & n1147 ;
  assign n1126 = ~n1122 & n1125 ;
  assign n1127 = ~n1119 & n1126 ;
  assign n1118 = n863 & ~n1117 ;
  assign n1128 = n1127 ^ n1118 ;
  assign n1149 = n1148 ^ n1128 ;
  assign n1196 = n1195 ^ n1149 ;
  assign n1201 = n1200 ^ n1196 ;
  assign n1203 = n1117 & n1201 ;
  assign n1202 = n863 & ~n1201 ;
  assign n1204 = n1203 ^ n1202 ;
  assign n859 = n771 & n857 ;
  assign n858 = n515 & ~n857 ;
  assign n860 = n859 ^ n858 ;
  assign n1206 = n1204 ^ n860 ;
  assign n1211 = n779 & n857 ;
  assign n1210 = n776 & ~n857 ;
  assign n1212 = n1211 ^ n1210 ;
  assign n1208 = n1122 & n1201 ;
  assign n1207 = n1125 & ~n1201 ;
  assign n1209 = n1208 ^ n1207 ;
  assign n1216 = n1212 ^ n1209 ;
  assign n1217 = ~n1206 & ~n1216 ;
  assign n1222 = n787 & n857 ;
  assign n1221 = n790 & ~n857 ;
  assign n1223 = n1222 ^ n1221 ;
  assign n1219 = n1133 & n1201 ;
  assign n1218 = n1136 & ~n1201 ;
  assign n1220 = n1219 ^ n1218 ;
  assign n1225 = n1223 ^ n1220 ;
  assign n1230 = n795 & n857 ;
  assign n1229 = n798 & ~n857 ;
  assign n1231 = n1230 ^ n1229 ;
  assign n1227 = n1141 & n1201 ;
  assign n1226 = n1144 & ~n1201 ;
  assign n1228 = n1227 ^ n1226 ;
  assign n1237 = n1231 ^ n1228 ;
  assign n1238 = ~n1225 & ~n1237 ;
  assign n1239 = n1217 & n1238 ;
  assign n1244 = n809 & n857 ;
  assign n1243 = n812 & ~n857 ;
  assign n1245 = n1244 ^ n1243 ;
  assign n1241 = n1155 & n1201 ;
  assign n1240 = n1158 & ~n1201 ;
  assign n1242 = n1241 ^ n1240 ;
  assign n1247 = n1245 ^ n1242 ;
  assign n1252 = n817 & n857 ;
  assign n1251 = n820 & ~n857 ;
  assign n1253 = n1252 ^ n1251 ;
  assign n1249 = n1163 & n1201 ;
  assign n1248 = n1166 & ~n1201 ;
  assign n1250 = n1249 ^ n1248 ;
  assign n1257 = n1253 ^ n1250 ;
  assign n1258 = ~n1247 & ~n1257 ;
  assign n1263 = n828 & n857 ;
  assign n1262 = n831 & ~n857 ;
  assign n1264 = n1263 ^ n1262 ;
  assign n1260 = n1174 & n1201 ;
  assign n1259 = n1177 & ~n1201 ;
  assign n1261 = n1260 ^ n1259 ;
  assign n1266 = n1264 ^ n1261 ;
  assign n1284 = n1183 & n1201 ;
  assign n1282 = n1187 & n1201 ;
  assign n1283 = n1282 ^ n1187 ;
  assign n1285 = n1284 ^ n1283 ;
  assign n1267 = n835 & ~n857 ;
  assign n1268 = n1267 ^ n1184 ;
  assign n1286 = n1285 ^ n1268 ;
  assign n1287 = ~n1266 & ~n1286 ;
  assign n1288 = n1258 & n1287 ;
  assign n1289 = n1239 & n1288 ;
  assign n1271 = n1187 & n1268 ;
  assign n1272 = ~n1201 & n1271 ;
  assign n1269 = n1183 & n1268 ;
  assign n1270 = n1201 & n1269 ;
  assign n1273 = n1272 ^ n1270 ;
  assign n1274 = n1273 ^ n1268 ;
  assign n1275 = n1266 & n1274 ;
  assign n1276 = n1275 ^ n1274 ;
  assign n1265 = ~n1261 & n1264 ;
  assign n1277 = n1276 ^ n1265 ;
  assign n1278 = n1258 & n1277 ;
  assign n1254 = ~n1250 & n1253 ;
  assign n1255 = ~n1247 & n1254 ;
  assign n1246 = ~n1242 & n1245 ;
  assign n1256 = n1255 ^ n1246 ;
  assign n1279 = n1278 ^ n1256 ;
  assign n1280 = n1239 & n1279 ;
  assign n1232 = ~n1228 & n1231 ;
  assign n1233 = ~n1225 & n1232 ;
  assign n1224 = ~n1220 & n1223 ;
  assign n1234 = n1233 ^ n1224 ;
  assign n1235 = n1217 & n1234 ;
  assign n1213 = ~n1209 & n1212 ;
  assign n1214 = ~n1206 & n1213 ;
  assign n1205 = n860 & ~n1204 ;
  assign n1215 = n1214 ^ n1205 ;
  assign n1236 = n1235 ^ n1215 ;
  assign n1281 = n1280 ^ n1236 ;
  assign n1290 = n1289 ^ n1281 ;
  assign n1293 = n1204 & n1290 ;
  assign n1291 = n860 & n1290 ;
  assign n1292 = n1291 ^ n860 ;
  assign n1294 = n1293 ^ n1292 ;
  assign n1297 = n1209 & n1290 ;
  assign n1295 = n1212 & n1290 ;
  assign n1296 = n1295 ^ n1212 ;
  assign n1298 = n1297 ^ n1296 ;
  assign n1301 = n1220 & n1290 ;
  assign n1299 = n1223 & n1290 ;
  assign n1300 = n1299 ^ n1223 ;
  assign n1302 = n1301 ^ n1300 ;
  assign n1305 = n1228 & n1290 ;
  assign n1303 = n1231 & n1290 ;
  assign n1304 = n1303 ^ n1231 ;
  assign n1306 = n1305 ^ n1304 ;
  assign n1309 = n1242 & n1290 ;
  assign n1307 = n1245 & n1290 ;
  assign n1308 = n1307 ^ n1245 ;
  assign n1310 = n1309 ^ n1308 ;
  assign n1313 = n1250 & n1290 ;
  assign n1311 = n1253 & n1290 ;
  assign n1312 = n1311 ^ n1253 ;
  assign n1314 = n1313 ^ n1312 ;
  assign n1317 = n1261 & n1290 ;
  assign n1315 = n1264 & n1290 ;
  assign n1316 = n1315 ^ n1264 ;
  assign n1318 = n1317 ^ n1316 ;
  assign n1321 = n1285 & n1290 ;
  assign n1319 = n1268 & n1290 ;
  assign n1320 = n1319 ^ n1268 ;
  assign n1322 = n1321 ^ n1320 ;
  assign n1323 = n1293 ^ n1204 ;
  assign n1324 = n1323 ^ n1291 ;
  assign n1325 = n1297 ^ n1209 ;
  assign n1326 = n1325 ^ n1295 ;
  assign n1327 = n1301 ^ n1220 ;
  assign n1328 = n1327 ^ n1299 ;
  assign n1329 = n1305 ^ n1228 ;
  assign n1330 = n1329 ^ n1303 ;
  assign n1331 = n1309 ^ n1242 ;
  assign n1332 = n1331 ^ n1307 ;
  assign n1333 = n1313 ^ n1250 ;
  assign n1334 = n1333 ^ n1311 ;
  assign n1335 = n1317 ^ n1261 ;
  assign n1336 = n1335 ^ n1315 ;
  assign n1337 = n1321 ^ n1285 ;
  assign n1338 = n1337 ^ n1319 ;
  assign n1340 = n863 & n1201 ;
  assign n1339 = n1117 & ~n1201 ;
  assign n1341 = n1340 ^ n1339 ;
  assign n1343 = n1125 & n1201 ;
  assign n1342 = n1122 & ~n1201 ;
  assign n1344 = n1343 ^ n1342 ;
  assign n1346 = n1136 & n1201 ;
  assign n1345 = n1133 & ~n1201 ;
  assign n1347 = n1346 ^ n1345 ;
  assign n1349 = n1144 & n1201 ;
  assign n1348 = n1141 & ~n1201 ;
  assign n1350 = n1349 ^ n1348 ;
  assign n1352 = n1158 & n1201 ;
  assign n1351 = n1155 & ~n1201 ;
  assign n1353 = n1352 ^ n1351 ;
  assign n1355 = n1166 & n1201 ;
  assign n1354 = n1163 & ~n1201 ;
  assign n1356 = n1355 ^ n1354 ;
  assign n1358 = n1177 & n1201 ;
  assign n1357 = n1174 & ~n1201 ;
  assign n1359 = n1358 ^ n1357 ;
  assign n1360 = n1183 & ~n1201 ;
  assign n1361 = n1360 ^ n1282 ;
  assign n1363 = n866 & n1114 ;
  assign n1362 = n1032 & ~n1114 ;
  assign n1364 = n1363 ^ n1362 ;
  assign n1366 = n1040 & n1114 ;
  assign n1365 = n1037 & ~n1114 ;
  assign n1367 = n1366 ^ n1365 ;
  assign n1369 = n1051 & n1114 ;
  assign n1368 = n1048 & ~n1114 ;
  assign n1370 = n1369 ^ n1368 ;
  assign n1372 = n1059 & n1114 ;
  assign n1371 = n1056 & ~n1114 ;
  assign n1373 = n1372 ^ n1371 ;
  assign n1375 = n1073 & n1114 ;
  assign n1374 = n1070 & ~n1114 ;
  assign n1376 = n1375 ^ n1374 ;
  assign n1378 = n1081 & n1114 ;
  assign n1377 = n1078 & ~n1114 ;
  assign n1379 = n1378 ^ n1377 ;
  assign n1381 = n1092 & n1114 ;
  assign n1380 = n1089 & ~n1114 ;
  assign n1382 = n1381 ^ n1380 ;
  assign n1383 = n1098 & ~n1114 ;
  assign n1384 = n1383 ^ n1180 ;
  assign n1386 = n869 & n1029 ;
  assign n1385 = n947 & ~n1029 ;
  assign n1387 = n1386 ^ n1385 ;
  assign n1389 = n955 & n1029 ;
  assign n1388 = n952 & ~n1029 ;
  assign n1390 = n1389 ^ n1388 ;
  assign n1392 = n966 & n1029 ;
  assign n1391 = n963 & ~n1029 ;
  assign n1393 = n1392 ^ n1391 ;
  assign n1395 = n974 & n1029 ;
  assign n1394 = n971 & ~n1029 ;
  assign n1396 = n1395 ^ n1394 ;
  assign n1398 = n988 & n1029 ;
  assign n1397 = n985 & ~n1029 ;
  assign n1399 = n1398 ^ n1397 ;
  assign n1401 = n996 & n1029 ;
  assign n1400 = n993 & ~n1029 ;
  assign n1402 = n1401 ^ n1400 ;
  assign n1404 = n1007 & n1029 ;
  assign n1403 = n1004 & ~n1029 ;
  assign n1405 = n1404 ^ n1403 ;
  assign n1406 = n1013 & ~n1029 ;
  assign n1407 = n1406 ^ n1095 ;
  assign n1409 = n872 & n944 ;
  assign n1408 = x40 & ~n944 ;
  assign n1410 = n1409 ^ n1408 ;
  assign n1412 = n877 & n944 ;
  assign n1411 = x41 & ~n944 ;
  assign n1413 = n1412 ^ n1411 ;
  assign n1415 = n885 & n944 ;
  assign n1414 = x42 & ~n944 ;
  assign n1416 = n1415 ^ n1414 ;
  assign n1418 = n890 & n944 ;
  assign n1417 = x43 & ~n944 ;
  assign n1419 = n1418 ^ n1417 ;
  assign n1421 = n901 & n944 ;
  assign n1420 = x44 & ~n944 ;
  assign n1422 = n1421 ^ n1420 ;
  assign n1424 = n906 & n944 ;
  assign n1423 = x45 & ~n944 ;
  assign n1425 = n1424 ^ n1423 ;
  assign n1427 = n938 & n944 ;
  assign n1426 = x46 & ~n944 ;
  assign n1428 = n1427 ^ n1426 ;
  assign n1429 = x47 & ~n944 ;
  assign n1430 = n1429 ^ n1010 ;
  assign y0 = n1294 ;
  assign y1 = n1298 ;
  assign y2 = n1302 ;
  assign y3 = n1306 ;
  assign y4 = n1310 ;
  assign y5 = n1314 ;
  assign y6 = n1318 ;
  assign y7 = n1322 ;
  assign y8 = n1324 ;
  assign y9 = n1326 ;
  assign y10 = n1328 ;
  assign y11 = n1330 ;
  assign y12 = n1332 ;
  assign y13 = n1334 ;
  assign y14 = n1336 ;
  assign y15 = n1338 ;
  assign y16 = n1341 ;
  assign y17 = n1344 ;
  assign y18 = n1347 ;
  assign y19 = n1350 ;
  assign y20 = n1353 ;
  assign y21 = n1356 ;
  assign y22 = n1359 ;
  assign y23 = n1361 ;
  assign y24 = n1364 ;
  assign y25 = n1367 ;
  assign y26 = n1370 ;
  assign y27 = n1373 ;
  assign y28 = n1376 ;
  assign y29 = n1379 ;
  assign y30 = n1382 ;
  assign y31 = n1384 ;
  assign y32 = n1387 ;
  assign y33 = n1390 ;
  assign y34 = n1393 ;
  assign y35 = n1396 ;
  assign y36 = n1399 ;
  assign y37 = n1402 ;
  assign y38 = n1405 ;
  assign y39 = n1407 ;
  assign y40 = n1410 ;
  assign y41 = n1413 ;
  assign y42 = n1416 ;
  assign y43 = n1419 ;
  assign y44 = n1422 ;
  assign y45 = n1425 ;
  assign y46 = n1428 ;
  assign y47 = n1430 ;
endmodule
