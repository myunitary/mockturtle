module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 ;
  assign n61 = x27 & x28 ;
  assign n62 = x29 & n61 ;
  assign n68 = x15 & x16 ;
  assign n69 = n68 ^ x15 ;
  assign n70 = x12 & x13 ;
  assign n71 = n70 ^ x12 ;
  assign n72 = n71 ^ x13 ;
  assign n164 = n69 & ~n72 ;
  assign n165 = x19 & x25 ;
  assign n166 = ~x26 & n165 ;
  assign n167 = n164 & n166 ;
  assign n168 = n62 & n167 ;
  assign n120 = x20 & ~x21 ;
  assign n121 = x22 & x23 ;
  assign n122 = n121 ^ x23 ;
  assign n169 = n120 & n122 ;
  assign n76 = x9 & x10 ;
  assign n77 = n76 ^ x9 ;
  assign n78 = n77 ^ x10 ;
  assign n170 = x0 & x1 ;
  assign n171 = ~n78 & n170 ;
  assign n172 = n169 & n171 ;
  assign n173 = x6 & x7 ;
  assign n174 = x8 & x11 ;
  assign n175 = n173 & n174 ;
  assign n176 = x2 & x3 ;
  assign n177 = x4 & x5 ;
  assign n178 = n176 & n177 ;
  assign n179 = n175 & n178 ;
  assign n180 = n172 & n179 ;
  assign n181 = n168 & n180 ;
  assign n140 = x11 & n78 ;
  assign n141 = n140 ^ x11 ;
  assign n142 = n141 ^ x11 ;
  assign n182 = ~n72 & ~n142 ;
  assign n183 = n182 ^ x14 ;
  assign n79 = n69 & n78 ;
  assign n80 = x11 & x14 ;
  assign n81 = ~n72 & n80 ;
  assign n82 = n79 & n81 ;
  assign n73 = x14 & ~n72 ;
  assign n74 = n73 ^ x14 ;
  assign n75 = n69 & n74 ;
  assign n83 = n82 ^ n75 ;
  assign n84 = n83 ^ x16 ;
  assign n187 = ~x18 & ~n84 ;
  assign n188 = ~n183 & n187 ;
  assign n189 = n181 & n188 ;
  assign n184 = ~x17 & ~x18 ;
  assign n185 = ~n183 & n184 ;
  assign n186 = n181 & n185 ;
  assign n190 = n189 ^ n186 ;
  assign n65 = x19 & x20 ;
  assign n64 = ~x21 & ~x22 ;
  assign n85 = x17 & ~x18 ;
  assign n86 = n64 & n85 ;
  assign n87 = n65 & n86 ;
  assign n88 = n84 & n87 ;
  assign n66 = x18 & n65 ;
  assign n67 = n64 & n66 ;
  assign n89 = n88 ^ n67 ;
  assign n90 = n89 ^ n64 ;
  assign n91 = x23 & x24 ;
  assign n92 = x25 & ~x26 ;
  assign n93 = n91 & n92 ;
  assign n94 = n62 & n93 ;
  assign n95 = ~n90 & n94 ;
  assign n63 = ~x26 & n62 ;
  assign n96 = n95 ^ n63 ;
  assign n97 = n96 ^ n62 ;
  assign n223 = n65 ^ x18 ;
  assign n197 = n64 ^ x23 ;
  assign n224 = n223 ^ n197 ;
  assign n137 = x17 & n84 ;
  assign n138 = n137 ^ x17 ;
  assign n139 = n138 ^ x17 ;
  assign n214 = n64 & n65 ;
  assign n215 = ~x18 & ~x23 ;
  assign n216 = n214 & n215 ;
  assign n217 = ~n139 & n216 ;
  assign n212 = ~x23 & ~n65 ;
  assign n213 = ~n64 & n212 ;
  assign n218 = n217 ^ n213 ;
  assign n209 = x18 & ~n64 ;
  assign n210 = ~n65 & n209 ;
  assign n211 = n139 & n210 ;
  assign n219 = n218 ^ n211 ;
  assign n192 = n65 ^ n64 ;
  assign n193 = n64 ^ x18 ;
  assign n194 = n192 & ~n193 ;
  assign n195 = n194 ^ x18 ;
  assign n204 = n195 ^ n139 ;
  assign n203 = n192 ^ x23 ;
  assign n205 = n204 ^ n203 ;
  assign n206 = n139 ^ n65 ;
  assign n207 = n206 ^ n195 ;
  assign n208 = n205 & n207 ;
  assign n220 = n219 ^ n208 ;
  assign n196 = n195 ^ n65 ;
  assign n198 = n197 ^ n196 ;
  assign n200 = x17 & ~n198 ;
  assign n201 = n84 & n200 ;
  assign n199 = n195 & ~n198 ;
  assign n202 = n201 ^ n199 ;
  assign n221 = n220 ^ n202 ;
  assign n222 = n221 ^ n194 ;
  assign n225 = n224 ^ n222 ;
  assign n226 = n225 ^ x23 ;
  assign n227 = ~n97 & n226 ;
  assign n191 = ~x24 & ~n97 ;
  assign n228 = n227 ^ n191 ;
  assign n229 = n190 & n228 ;
  assign n230 = n229 ^ n97 ;
  assign n98 = x7 & x8 ;
  assign n99 = n98 ^ x7 ;
  assign n100 = n99 ^ x8 ;
  assign n101 = n77 & ~n100 ;
  assign n102 = x3 & x4 ;
  assign n103 = n102 ^ x3 ;
  assign n104 = n103 ^ x4 ;
  assign n105 = x5 & x6 ;
  assign n106 = n105 ^ x5 ;
  assign n107 = n106 ^ x6 ;
  assign n108 = ~n104 & ~n107 ;
  assign n109 = n101 & n108 ;
  assign n110 = x24 & x25 ;
  assign n111 = x26 & n110 ;
  assign n112 = n111 ^ n110 ;
  assign n113 = x13 & x14 ;
  assign n114 = n113 ^ x14 ;
  assign n115 = x18 & x19 ;
  assign n116 = n115 ^ x19 ;
  assign n117 = n114 & n116 ;
  assign n118 = n112 & n117 ;
  assign n119 = n109 & n118 ;
  assign n123 = x1 & x2 ;
  assign n124 = n123 ^ x1 ;
  assign n125 = n124 ^ x2 ;
  assign n126 = n122 & ~n125 ;
  assign n127 = n120 & n126 ;
  assign n132 = x11 & ~x12 ;
  assign n133 = n78 & n132 ;
  assign n134 = n127 & n133 ;
  assign n135 = n119 & n134 ;
  assign n128 = ~x11 & x12 ;
  assign n129 = ~n78 & n128 ;
  assign n130 = n127 & n129 ;
  assign n131 = n119 & n130 ;
  assign n136 = n135 ^ n131 ;
  assign n143 = n142 ^ n72 ;
  assign n144 = n72 ^ x14 ;
  assign n145 = x14 & ~n144 ;
  assign n146 = n145 ^ x14 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = n147 ^ x14 ;
  assign n149 = n148 ^ n142 ;
  assign n150 = ~n143 & n149 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = n151 ^ n147 ;
  assign n153 = n152 ^ n142 ;
  assign n159 = n69 & n153 ;
  assign n160 = n139 & n159 ;
  assign n161 = n136 & n160 ;
  assign n154 = x15 & n153 ;
  assign n155 = n154 ^ x15 ;
  assign n156 = n155 ^ n153 ;
  assign n157 = n139 & ~n156 ;
  assign n158 = n136 & n157 ;
  assign n162 = n161 ^ n158 ;
  assign n163 = n97 & ~n162 ;
  assign n231 = n230 ^ n163 ;
  assign n232 = x36 & x37 ;
  assign n233 = x38 & x41 ;
  assign n234 = n232 & n233 ;
  assign n235 = x32 & x33 ;
  assign n236 = x34 & x35 ;
  assign n237 = n235 & n236 ;
  assign n238 = n234 & n237 ;
  assign n239 = x57 & x58 ;
  assign n240 = x59 & n239 ;
  assign n241 = x46 & x47 ;
  assign n242 = n241 ^ x47 ;
  assign n243 = x50 & x56 ;
  assign n244 = n243 ^ x50 ;
  assign n245 = n242 & n244 ;
  assign n246 = n240 & n245 ;
  assign n247 = n238 & n246 ;
  assign n248 = x39 & x40 ;
  assign n249 = n248 ^ x39 ;
  assign n250 = n249 ^ x40 ;
  assign n251 = x41 & x42 ;
  assign n261 = n250 & n251 ;
  assign n262 = x43 & n261 ;
  assign n263 = x44 & x45 ;
  assign n264 = n263 ^ x45 ;
  assign n265 = n262 & n264 ;
  assign n266 = n265 ^ n264 ;
  assign n252 = n251 ^ x41 ;
  assign n253 = n250 & n252 ;
  assign n254 = n253 ^ x42 ;
  assign n255 = x43 & x44 ;
  assign n256 = n255 ^ x44 ;
  assign n257 = n254 & n256 ;
  assign n258 = n257 ^ n256 ;
  assign n259 = n258 ^ x44 ;
  assign n260 = x45 & ~n259 ;
  assign n267 = n266 ^ n260 ;
  assign n268 = n247 & n267 ;
  assign n269 = x45 & x46 ;
  assign n270 = n269 ^ x45 ;
  assign n272 = n256 & n270 ;
  assign n273 = n254 & n272 ;
  assign n274 = n273 ^ n272 ;
  assign n271 = x44 & n270 ;
  assign n275 = n274 ^ n271 ;
  assign n276 = n275 ^ x46 ;
  assign n277 = x49 ^ x48 ;
  assign n278 = x47 & n277 ;
  assign n279 = n276 & n278 ;
  assign n280 = n279 ^ n277 ;
  assign n281 = n280 ^ x49 ;
  assign n282 = x54 & x55 ;
  assign n283 = x30 & x31 ;
  assign n284 = n282 & n283 ;
  assign n285 = ~x48 & ~x49 ;
  assign n286 = ~n250 & ~n285 ;
  assign n287 = n284 & n286 ;
  assign n288 = ~n281 & n287 ;
  assign n289 = n268 & n288 ;
  assign n290 = x47 & ~x48 ;
  assign n291 = n276 & n290 ;
  assign n292 = n291 ^ x48 ;
  assign n293 = x49 & x50 ;
  assign n294 = x52 & x53 ;
  assign n295 = n294 ^ x53 ;
  assign n296 = n293 & ~n295 ;
  assign n297 = n292 & n296 ;
  assign n298 = n297 ^ n295 ;
  assign n307 = x53 & n282 ;
  assign n300 = x51 & x52 ;
  assign n301 = n300 ^ x51 ;
  assign n302 = n301 ^ x52 ;
  assign n316 = n307 ^ n302 ;
  assign n317 = n307 & ~n316 ;
  assign n308 = n307 ^ x49 ;
  assign n299 = x50 ^ x49 ;
  assign n303 = n302 ^ n299 ;
  assign n304 = n302 ^ x49 ;
  assign n305 = ~n303 & ~n304 ;
  assign n306 = n305 ^ x50 ;
  assign n309 = n308 ^ n306 ;
  assign n313 = ~x49 & n309 ;
  assign n312 = ~x48 & n309 ;
  assign n314 = n313 ^ n312 ;
  assign n310 = n290 & n309 ;
  assign n311 = n276 & n310 ;
  assign n315 = n314 ^ n311 ;
  assign n318 = n317 ^ n315 ;
  assign n319 = n318 ^ n305 ;
  assign n320 = n319 ^ n303 ;
  assign n327 = x53 & ~x56 ;
  assign n328 = n282 & n327 ;
  assign n329 = n328 ^ x56 ;
  assign n330 = n240 & ~n329 ;
  assign n331 = ~n320 & n330 ;
  assign n321 = ~x56 & x59 ;
  assign n322 = n239 & n321 ;
  assign n323 = n317 & n322 ;
  assign n324 = n323 ^ n322 ;
  assign n325 = ~n320 & n324 ;
  assign n326 = n325 ^ n324 ;
  assign n332 = n331 ^ n326 ;
  assign n333 = n332 ^ n240 ;
  assign n334 = x52 & ~x53 ;
  assign n335 = n293 & ~n334 ;
  assign n337 = n290 & n335 ;
  assign n338 = n276 & n337 ;
  assign n336 = x48 & n335 ;
  assign n339 = n338 ^ n336 ;
  assign n340 = n333 & n339 ;
  assign n341 = n340 ^ n333 ;
  assign n342 = ~n298 & n341 ;
  assign n343 = n342 ^ n341 ;
  assign n344 = n289 & n343 ;
  assign n345 = n344 ^ n333 ;
  assign n351 = ~x56 & x57 ;
  assign n352 = ~x46 & ~x51 ;
  assign n353 = n351 & n352 ;
  assign n354 = x41 & ~x43 ;
  assign n355 = n263 & n354 ;
  assign n356 = x39 & ~x40 ;
  assign n357 = ~x37 & ~x38 ;
  assign n358 = n356 & n357 ;
  assign n359 = n355 & n358 ;
  assign n360 = n353 & n359 ;
  assign n361 = x41 & n250 ;
  assign n362 = n361 ^ x41 ;
  assign n363 = n362 ^ x41 ;
  assign n364 = n363 ^ x42 ;
  assign n365 = x47 & x48 ;
  assign n366 = n293 & n295 ;
  assign n367 = n365 & n366 ;
  assign n368 = n367 ^ n366 ;
  assign n369 = x33 & x34 ;
  assign n370 = n369 ^ x33 ;
  assign n371 = n370 ^ x34 ;
  assign n372 = x35 & x36 ;
  assign n373 = n372 ^ x35 ;
  assign n374 = n373 ^ x36 ;
  assign n375 = ~n371 & ~n374 ;
  assign n376 = x31 & x32 ;
  assign n377 = n376 ^ x31 ;
  assign n378 = n377 ^ x32 ;
  assign n379 = n282 & ~n378 ;
  assign n380 = n375 & n379 ;
  assign n381 = n368 & n380 ;
  assign n382 = ~n364 & n381 ;
  assign n383 = n382 ^ n381 ;
  assign n384 = n360 & n383 ;
  assign n346 = x47 & n276 ;
  assign n347 = n346 ^ x47 ;
  assign n348 = n347 ^ x47 ;
  assign n349 = x48 & ~n276 ;
  assign n350 = ~n348 & ~n349 ;
  assign n385 = n384 ^ n350 ;
  assign n386 = ~x0 & ~x30 ;
  assign n387 = n386 ^ n350 ;
  assign n388 = ~n386 & ~n387 ;
  assign n389 = n388 ^ n350 ;
  assign n390 = ~n385 & n389 ;
  assign n391 = n390 ^ n388 ;
  assign n392 = n391 ^ n384 ;
  assign n416 = n190 & n226 ;
  assign n415 = ~x24 & n190 ;
  assign n417 = n416 ^ n415 ;
  assign n420 = ~n392 & n417 ;
  assign n421 = n345 & n420 ;
  assign n395 = ~x0 & ~x51 ;
  assign n396 = n333 & n395 ;
  assign n397 = n396 ^ n333 ;
  assign n398 = n397 ^ n395 ;
  assign n399 = n298 & ~n339 ;
  assign n400 = n398 & n399 ;
  assign n401 = n289 & n400 ;
  assign n419 = n401 & n417 ;
  assign n422 = n421 ^ n419 ;
  assign n418 = n97 & n417 ;
  assign n423 = n422 ^ n418 ;
  assign n406 = ~x24 & n97 ;
  assign n407 = n190 & n406 ;
  assign n404 = n97 & n226 ;
  assign n405 = n190 & n404 ;
  assign n408 = n407 ^ n405 ;
  assign n403 = n97 & n162 ;
  assign n409 = n408 ^ n403 ;
  assign n411 = ~n392 & n409 ;
  assign n412 = n345 & n411 ;
  assign n410 = n401 & n409 ;
  assign n413 = n412 ^ n410 ;
  assign n414 = n413 ^ n409 ;
  assign n424 = n423 ^ n414 ;
  assign n393 = n345 & n392 ;
  assign n394 = n393 ^ n345 ;
  assign n402 = n401 ^ n394 ;
  assign n425 = n424 ^ n402 ;
  assign n426 = n425 ^ n97 ;
  assign n427 = n426 ^ n402 ;
  assign n428 = n403 ^ n97 ;
  assign n429 = n428 ^ n230 ;
  assign n430 = x0 & x30 ;
  assign n431 = n430 ^ n350 ;
  assign n432 = n430 & n431 ;
  assign n433 = n432 ^ n350 ;
  assign n434 = ~n385 & n433 ;
  assign n435 = n434 ^ n432 ;
  assign n436 = n435 ^ n384 ;
  assign n437 = n162 ^ n97 ;
  assign n438 = n333 ^ n97 ;
  assign n439 = ~n333 & ~n438 ;
  assign n440 = n439 ^ n333 ;
  assign n441 = n440 ^ n162 ;
  assign n442 = ~n437 & n441 ;
  assign n443 = n442 ^ n439 ;
  assign n444 = n443 ^ n162 ;
  assign n445 = n436 & n444 ;
  assign n446 = n445 ^ n444 ;
  assign n447 = n446 ^ n428 ;
  assign n448 = n447 ^ n428 ;
  assign n449 = n429 & n448 ;
  assign n450 = n449 ^ n429 ;
  assign n451 = n450 ^ n448 ;
  assign n452 = n451 ^ n447 ;
  assign n453 = n452 ^ n230 ;
  assign y0 = ~n231 ;
  assign y1 = ~n427 ;
  assign y2 = n453 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
