module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 ;
  assign n33 = x29 & x30 ;
  assign n34 = x27 & x28 ;
  assign n35 = n33 & n34 ;
  assign n36 = x26 & x27 ;
  assign n37 = n35 & n36 ;
  assign n38 = x22 & x23 ;
  assign n39 = x23 & x24 ;
  assign n40 = n38 & n39 ;
  assign n41 = x25 & x26 ;
  assign n42 = x24 & x25 ;
  assign n43 = n41 & n42 ;
  assign n44 = n40 & n43 ;
  assign n45 = ~n37 & ~n44 ;
  assign n46 = n34 & n36 ;
  assign n47 = n43 & n46 ;
  assign n48 = ~n45 & n47 ;
  assign n49 = x28 & x29 ;
  assign n50 = x30 & x31 ;
  assign n51 = n33 & n50 ;
  assign n52 = n49 & n51 ;
  assign n53 = n34 & n52 ;
  assign n54 = n36 & n41 ;
  assign n55 = n39 & n42 ;
  assign n56 = n54 & n55 ;
  assign n57 = ~n53 & ~n56 ;
  assign n58 = n34 & n49 ;
  assign n59 = n54 & n58 ;
  assign n60 = ~n57 & n59 ;
  assign n61 = n48 & n60 ;
  assign n62 = x10 & x11 ;
  assign n63 = x17 & x18 ;
  assign n64 = ~n62 & ~n63 ;
  assign n65 = x12 & x13 ;
  assign n66 = x13 & x14 ;
  assign n67 = n65 & n66 ;
  assign n68 = x14 & x15 ;
  assign n69 = x15 & x16 ;
  assign n70 = n68 & n69 ;
  assign n71 = n67 & n70 ;
  assign n72 = ~n64 & n71 ;
  assign n73 = x19 & x20 ;
  assign n74 = x18 & x19 ;
  assign n75 = n73 & n74 ;
  assign n76 = n63 & n74 ;
  assign n77 = x16 & x17 ;
  assign n78 = n69 & n77 ;
  assign n79 = n76 & n78 ;
  assign n80 = n75 & n79 ;
  assign n81 = ~n72 & ~n80 ;
  assign n82 = x11 & x12 ;
  assign n83 = ~n74 & ~n82 ;
  assign n84 = n66 & n68 ;
  assign n85 = n78 & n84 ;
  assign n86 = ~n83 & n85 ;
  assign n87 = ~n81 & n86 ;
  assign n88 = x21 & x22 ;
  assign n89 = ~n68 & ~n88 ;
  assign n90 = n63 & n77 ;
  assign n91 = n75 & n90 ;
  assign n92 = ~n89 & n91 ;
  assign n93 = x20 & x21 ;
  assign n94 = n74 & n93 ;
  assign n95 = n90 & n94 ;
  assign n96 = n79 & n95 ;
  assign n97 = n92 & n96 ;
  assign n98 = ~n87 & ~n97 ;
  assign n99 = ~n61 & n98 ;
  assign n100 = n73 & n88 ;
  assign n101 = n75 & n100 ;
  assign n102 = n38 & n93 ;
  assign n103 = n101 & n102 ;
  assign n104 = n63 & n94 ;
  assign n105 = n103 & n104 ;
  assign n106 = ~n39 & ~n77 ;
  assign n107 = n105 & ~n106 ;
  assign n108 = ~n41 & ~n74 ;
  assign n109 = n39 & n88 ;
  assign n110 = n93 & n109 ;
  assign n111 = ~n108 & n110 ;
  assign n112 = n46 & n56 ;
  assign n113 = ~n111 & ~n112 ;
  assign n114 = ~n36 & ~n73 ;
  assign n115 = n38 & n88 ;
  assign n116 = n55 & n115 ;
  assign n117 = ~n114 & n116 ;
  assign n118 = ~n113 & n117 ;
  assign n119 = ~n107 & ~n118 ;
  assign n120 = n99 & n119 ;
  assign n121 = x8 & x9 ;
  assign n122 = x7 & n121 ;
  assign n123 = x9 & x10 ;
  assign n124 = n62 & n123 ;
  assign n125 = n122 & n124 ;
  assign n126 = n62 & n82 ;
  assign n127 = n125 & n126 ;
  assign n128 = x7 & x8 ;
  assign n129 = x6 & x7 ;
  assign n130 = n128 & n129 ;
  assign n131 = n123 & n128 ;
  assign n132 = n130 & n131 ;
  assign n133 = n127 & n132 ;
  assign n134 = n65 & n82 ;
  assign n135 = n124 & n134 ;
  assign n136 = n67 & n135 ;
  assign n137 = n121 & n123 ;
  assign n138 = n126 & n137 ;
  assign n139 = n136 & n138 ;
  assign n140 = ~n133 & ~n139 ;
  assign n141 = n84 & n134 ;
  assign n142 = n70 & n141 ;
  assign n143 = n140 & ~n142 ;
  assign n144 = ~n68 & ~n128 ;
  assign n145 = n135 & ~n144 ;
  assign n146 = ~n143 & n145 ;
  assign n147 = x5 & x6 ;
  assign n148 = n129 & n147 ;
  assign n149 = x4 & x5 ;
  assign n150 = x3 & x4 ;
  assign n151 = n149 & n150 ;
  assign n152 = n148 & n151 ;
  assign n153 = n130 & n152 ;
  assign n154 = n147 & n149 ;
  assign n155 = x2 & x3 ;
  assign n156 = n150 & n155 ;
  assign n157 = n154 & n156 ;
  assign n158 = n153 & n157 ;
  assign n159 = n121 & n129 ;
  assign n160 = n147 & n159 ;
  assign n161 = n131 & n160 ;
  assign n162 = x1 & x2 ;
  assign n163 = n150 & n162 ;
  assign n164 = x0 & x1 ;
  assign n165 = n163 & n164 ;
  assign n166 = n149 & n155 ;
  assign n167 = n165 & n166 ;
  assign n168 = ~n161 & ~n167 ;
  assign n169 = ~n158 & n168 ;
  assign n170 = n154 & n159 ;
  assign n171 = n152 & n170 ;
  assign n172 = n148 & n157 ;
  assign n173 = n155 & n162 ;
  assign n174 = n151 & n173 ;
  assign n175 = n172 & n174 ;
  assign n176 = ~n171 & ~n175 ;
  assign n177 = ~n169 & ~n176 ;
  assign n178 = n130 & n154 ;
  assign n179 = n161 & n178 ;
  assign n180 = ~n133 & ~n179 ;
  assign n181 = n62 & n121 ;
  assign n182 = n132 & n181 ;
  assign n183 = n160 & n182 ;
  assign n184 = ~n180 & n183 ;
  assign n185 = ~n177 & ~n184 ;
  assign n186 = ~n146 & n185 ;
  assign n187 = n120 & n186 ;
  assign n386 = ~n69 & ~n155 ;
  assign n387 = ~n33 & ~n49 ;
  assign n388 = n386 & n387 ;
  assign n389 = ~n62 & ~n82 ;
  assign n390 = ~n65 & ~n66 ;
  assign n391 = n389 & n390 ;
  assign n392 = n388 & n391 ;
  assign n393 = ~n50 & ~n88 ;
  assign n394 = ~n42 & n393 ;
  assign n395 = ~n34 & ~n36 ;
  assign n396 = n108 & n395 ;
  assign n397 = n394 & n396 ;
  assign n398 = n392 & n397 ;
  assign n399 = ~n129 & ~n147 ;
  assign n400 = n106 & n399 ;
  assign n333 = ~n38 & ~n93 ;
  assign n401 = ~n63 & ~n73 ;
  assign n402 = n333 & n401 ;
  assign n403 = n400 & n402 ;
  assign n404 = ~n121 & ~n123 ;
  assign n405 = ~n162 & ~n164 ;
  assign n406 = n404 & n405 ;
  assign n407 = ~n149 & ~n150 ;
  assign n408 = n144 & n407 ;
  assign n409 = n406 & n408 ;
  assign n410 = n403 & n409 ;
  assign n411 = n398 & n410 ;
  assign n357 = ~x18 & ~x19 ;
  assign n358 = ~x21 & ~x22 ;
  assign n359 = n357 & n358 ;
  assign n360 = ~x14 & ~x15 ;
  assign n361 = ~x16 & ~x17 ;
  assign n362 = n360 & n361 ;
  assign n363 = n359 & n362 ;
  assign n364 = ~x28 & ~x29 ;
  assign n365 = ~x30 & ~x31 ;
  assign n366 = n364 & n365 ;
  assign n367 = ~x23 & ~x24 ;
  assign n368 = ~x25 & ~x27 ;
  assign n369 = n367 & n368 ;
  assign n370 = n366 & n369 ;
  assign n371 = n363 & n370 ;
  assign n372 = ~x1 & ~x2 ;
  assign n373 = ~x4 & ~x5 ;
  assign n374 = n372 & n373 ;
  assign n215 = ~x20 & ~x26 ;
  assign n321 = ~x0 & ~x3 ;
  assign n375 = n215 & n321 ;
  assign n376 = n374 & n375 ;
  assign n377 = ~x10 & ~x11 ;
  assign n378 = ~x12 & ~x13 ;
  assign n379 = n377 & n378 ;
  assign n380 = ~x6 & ~x7 ;
  assign n381 = ~x8 & ~x9 ;
  assign n382 = n380 & n381 ;
  assign n383 = n379 & n382 ;
  assign n384 = n376 & n383 ;
  assign n385 = n371 & n384 ;
  assign n412 = n411 ^ n385 ;
  assign n314 = ~n40 & ~n43 ;
  assign n315 = ~n46 & ~n51 ;
  assign n316 = n314 & n315 ;
  assign n317 = ~n84 & ~n137 ;
  assign n224 = n33 & n49 ;
  assign n318 = ~n70 & ~n224 ;
  assign n319 = n317 & n318 ;
  assign n320 = n316 & n319 ;
  assign n322 = n162 & ~n321 ;
  assign n323 = ~x15 & x16 ;
  assign n324 = x17 & ~x18 ;
  assign n325 = n323 & n324 ;
  assign n326 = n325 ^ n77 ;
  assign n327 = ~n322 & ~n326 ;
  assign n328 = ~n54 & ~n55 ;
  assign n221 = x19 & n93 ;
  assign n329 = ~n58 & ~n221 ;
  assign n330 = n328 & n329 ;
  assign n331 = n327 & n330 ;
  assign n332 = n320 & n331 ;
  assign n334 = n88 & ~n333 ;
  assign n335 = ~x17 & x18 ;
  assign n336 = x19 & ~x20 ;
  assign n337 = n335 & n336 ;
  assign n338 = n337 ^ n74 ;
  assign n339 = ~n148 & ~n151 ;
  assign n340 = ~n338 & n339 ;
  assign n341 = ~n334 & n340 ;
  assign n342 = ~x9 & x10 ;
  assign n343 = x11 & ~x12 ;
  assign n344 = n342 & n343 ;
  assign n345 = n344 ^ n62 ;
  assign n346 = ~x11 & x12 ;
  assign n347 = x13 & ~x14 ;
  assign n348 = n346 & n347 ;
  assign n349 = n348 ^ n65 ;
  assign n350 = ~n345 & ~n349 ;
  assign n351 = ~n130 & ~n154 ;
  assign n352 = ~n122 & ~n156 ;
  assign n353 = n351 & n352 ;
  assign n354 = n350 & n353 ;
  assign n355 = n341 & n354 ;
  assign n356 = n332 & n355 ;
  assign n413 = n412 ^ n356 ;
  assign n272 = n38 & n42 ;
  assign n273 = n155 & n164 ;
  assign n274 = ~n272 & ~n273 ;
  assign n275 = n62 & n65 ;
  assign n276 = n63 & n69 ;
  assign n277 = ~n275 & ~n276 ;
  assign n278 = n274 & n277 ;
  assign n279 = n147 & n150 ;
  assign n280 = n66 & n82 ;
  assign n281 = ~n279 & ~n280 ;
  assign n282 = n128 & n147 ;
  assign n283 = n34 & n41 ;
  assign n284 = ~n282 & ~n283 ;
  assign n285 = n281 & n284 ;
  assign n286 = n278 & n285 ;
  assign n287 = n63 & n75 ;
  assign n288 = n129 & n149 ;
  assign n289 = n74 & n77 ;
  assign n290 = ~n288 & ~n289 ;
  assign n291 = ~n287 & n290 ;
  assign n292 = n66 & n69 ;
  assign n293 = n82 & n123 ;
  assign n294 = ~n292 & ~n293 ;
  assign n295 = n39 & n41 ;
  assign n296 = n65 & n68 ;
  assign n297 = ~n295 & ~n296 ;
  assign n298 = n294 & n297 ;
  assign n299 = n291 & n298 ;
  assign n300 = n286 & n299 ;
  assign n231 = n42 & n54 ;
  assign n232 = ~n52 & ~n231 ;
  assign n301 = ~n131 & ~n159 ;
  assign n302 = ~n163 & ~n166 ;
  assign n303 = n301 & n302 ;
  assign n304 = n232 & n303 ;
  assign n305 = ~n94 & ~n109 ;
  assign n233 = n36 & n49 ;
  assign n235 = n68 & n77 ;
  assign n306 = ~n233 & ~n235 ;
  assign n307 = n305 & n306 ;
  assign n308 = ~n35 & ~n181 ;
  assign n309 = ~n100 & ~n102 ;
  assign n310 = n308 & n309 ;
  assign n311 = n307 & n310 ;
  assign n312 = n304 & n311 ;
  assign n313 = n300 & n312 ;
  assign n414 = n413 ^ n313 ;
  assign n207 = n67 & n126 ;
  assign n247 = ~n116 & ~n207 ;
  assign n217 = n70 & n90 ;
  assign n222 = n115 & n221 ;
  assign n248 = ~n217 & ~n222 ;
  assign n249 = n247 & n248 ;
  assign n250 = ~n71 & ~n79 ;
  assign n251 = ~n85 & ~n91 ;
  assign n252 = n250 & n251 ;
  assign n253 = n249 & n252 ;
  assign n254 = n45 & n57 ;
  assign n255 = n253 & n254 ;
  assign n256 = ~n101 & ~n104 ;
  assign n257 = ~n110 & n256 ;
  assign n258 = ~n152 & ~n157 ;
  assign n259 = ~n160 & n258 ;
  assign n260 = ~n132 & ~n165 ;
  assign n261 = n259 & n260 ;
  assign n262 = ~n138 & ~n141 ;
  assign n263 = ~n47 & ~n59 ;
  assign n264 = n262 & n263 ;
  assign n265 = ~n125 & ~n174 ;
  assign n266 = ~n135 & ~n178 ;
  assign n267 = n265 & n266 ;
  assign n268 = n264 & n267 ;
  assign n269 = n261 & n268 ;
  assign n270 = n257 & n269 ;
  assign n271 = n255 & n270 ;
  assign n415 = n414 ^ n271 ;
  assign n193 = n154 & n174 ;
  assign n205 = ~n112 & ~n193 ;
  assign n206 = n44 & n54 ;
  assign n208 = n84 & n207 ;
  assign n209 = ~n206 & ~n208 ;
  assign n210 = n205 & n209 ;
  assign n211 = ~n136 & ~n142 ;
  assign n212 = ~n80 & ~n95 ;
  assign n213 = n211 & n212 ;
  assign n214 = n210 & n213 ;
  assign n216 = n116 & ~n215 ;
  assign n218 = ~x13 & ~x19 ;
  assign n219 = n217 & ~n218 ;
  assign n220 = ~n216 & ~n219 ;
  assign n223 = n40 & n222 ;
  assign n225 = n59 & n224 ;
  assign n226 = ~n223 & ~n225 ;
  assign n227 = n220 & n226 ;
  assign n228 = n168 & n227 ;
  assign n229 = n214 & n228 ;
  assign n230 = n100 & n104 ;
  assign n234 = ~n232 & n233 ;
  assign n236 = ~n138 & ~n235 ;
  assign n237 = n65 & ~n236 ;
  assign n238 = ~n234 & ~n237 ;
  assign n239 = ~n230 & n238 ;
  assign n240 = ~n153 & ~n170 ;
  assign n241 = ~n127 & ~n172 ;
  assign n242 = n240 & n241 ;
  assign n243 = ~n103 & ~n182 ;
  assign n244 = n242 & n243 ;
  assign n245 = n239 & n244 ;
  assign n246 = n229 & n245 ;
  assign n416 = n415 ^ n246 ;
  assign n188 = ~n48 & ~n60 ;
  assign n189 = ~n105 & n188 ;
  assign n190 = n176 & ~n179 ;
  assign n191 = n140 & ~n183 ;
  assign n192 = n190 & n191 ;
  assign n194 = n165 & n193 ;
  assign n195 = ~n96 & ~n111 ;
  assign n196 = ~n194 & n195 ;
  assign n197 = ~n86 & ~n92 ;
  assign n198 = ~n117 & n197 ;
  assign n199 = ~n72 & ~n145 ;
  assign n200 = ~n158 & n199 ;
  assign n201 = n198 & n200 ;
  assign n202 = n196 & n201 ;
  assign n203 = n192 & n202 ;
  assign n204 = n189 & n203 ;
  assign n417 = n416 ^ n204 ;
  assign n418 = ~n187 & ~n417 ;
  assign n431 = ~n313 & ~n385 ;
  assign n430 = n313 & ~n411 ;
  assign n432 = n431 ^ n430 ;
  assign n427 = ~n385 & n411 ;
  assign n428 = ~n356 & n427 ;
  assign n425 = ~n313 & ~n356 ;
  assign n423 = n385 & ~n411 ;
  assign n424 = n356 & n423 ;
  assign n426 = n425 ^ n424 ;
  assign n429 = n428 ^ n426 ;
  assign n433 = n432 ^ n429 ;
  assign n422 = n271 & ~n414 ;
  assign n434 = n433 ^ n422 ;
  assign n420 = n246 & n414 ;
  assign n419 = n246 & ~n271 ;
  assign n421 = n420 ^ n419 ;
  assign n435 = n434 ^ n421 ;
  assign n436 = n418 & ~n435 ;
  assign n447 = n433 ^ n413 ;
  assign n443 = n255 & n313 ;
  assign n444 = n270 & n443 ;
  assign n441 = n255 & n413 ;
  assign n442 = n270 & n441 ;
  assign n445 = n444 ^ n442 ;
  assign n446 = n445 ^ n313 ;
  assign n448 = n447 ^ n446 ;
  assign n451 = ~n246 & n448 ;
  assign n452 = ~n204 & n451 ;
  assign n449 = ~n415 & n448 ;
  assign n450 = ~n204 & n449 ;
  assign n453 = n452 ^ n450 ;
  assign n455 = ~n271 & n414 ;
  assign n438 = ~n356 & n385 ;
  assign n437 = n356 & n411 ;
  assign n439 = n438 ^ n437 ;
  assign n440 = n439 ^ n423 ;
  assign n456 = n433 & ~n440 ;
  assign n457 = ~n455 & n456 ;
  assign n458 = ~n453 & n457 ;
  assign n454 = n440 & ~n453 ;
  assign n459 = n458 ^ n454 ;
  assign n460 = n436 & ~n459 ;
  assign n461 = ~n246 & ~n415 ;
  assign n462 = n433 & n461 ;
  assign n466 = n459 & ~n462 ;
  assign n463 = ~n448 & ~n461 ;
  assign n464 = ~n462 & ~n463 ;
  assign n465 = n418 & n464 ;
  assign n467 = n466 ^ n465 ;
  assign n468 = ~n204 & n416 ;
  assign n469 = ~n418 & ~n468 ;
  assign n470 = n469 ^ n435 ;
  assign n471 = n417 ^ n187 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = 1'b0 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = n460 ;
  assign y29 = ~n467 ;
  assign y30 = n470 ;
  assign y31 = n471 ;
endmodule
