module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 ;
  assign n22 = x5 & x13 ;
  assign n23 = x6 & x14 ;
  assign n24 = n22 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n22 ^ x5 ;
  assign n28 = n27 ^ x13 ;
  assign n29 = x4 & x12 ;
  assign n30 = n29 ^ x4 ;
  assign n31 = n30 ^ x12 ;
  assign n32 = ~n28 & ~n31 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = ~n26 & ~n34 ;
  assign n36 = n35 ^ n34 ;
  assign n17 = x10 ^ x2 ;
  assign n37 = x11 ^ x3 ;
  assign n38 = ~n17 & n37 ;
  assign n39 = ~n29 & n38 ;
  assign n40 = ~n36 & n39 ;
  assign n41 = n40 ^ n39 ;
  assign n18 = x3 & x11 ;
  assign n19 = n18 ^ x3 ;
  assign n20 = n19 ^ x11 ;
  assign n21 = ~n17 & ~n20 ;
  assign n42 = n41 ^ n21 ;
  assign n49 = x14 ^ x6 ;
  assign n48 = x7 & x15 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = x13 ^ x5 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = ~n51 & n52 ;
  assign n54 = n53 ^ n49 ;
  assign n55 = n50 & ~n54 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = n56 ^ n48 ;
  assign n43 = x1 & x9 ;
  assign n44 = x8 & n43 ;
  assign n45 = n44 ^ n43 ;
  assign n58 = x12 ^ x4 ;
  assign n59 = n37 & n58 ;
  assign n60 = n45 & n59 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = n57 & n61 ;
  assign n63 = n42 & n62 ;
  assign n64 = n63 ^ n62 ;
  assign n46 = n42 & n45 ;
  assign n47 = n46 ^ n45 ;
  assign n65 = n64 ^ n47 ;
  assign n71 = n57 & n59 ;
  assign n66 = x9 ^ x1 ;
  assign n67 = x2 & x10 ;
  assign n68 = ~n66 & ~n67 ;
  assign n72 = ~x0 & x8 ;
  assign n73 = ~n43 & n72 ;
  assign n74 = n73 ^ x8 ;
  assign n75 = n74 ^ n43 ;
  assign n76 = n68 & ~n75 ;
  assign n77 = n76 ^ n68 ;
  assign n78 = n77 ^ n75 ;
  assign n79 = n71 & n78 ;
  assign n80 = n65 & n79 ;
  assign n69 = n65 & n68 ;
  assign n70 = n69 ^ n65 ;
  assign n81 = n80 ^ n70 ;
  assign n82 = n18 & n29 ;
  assign n83 = n82 ^ n18 ;
  assign n84 = n83 ^ n29 ;
  assign n85 = n67 ^ x2 ;
  assign n86 = n85 ^ x10 ;
  assign n87 = ~n20 & ~n86 ;
  assign n88 = n87 ^ n20 ;
  assign n89 = n88 ^ n86 ;
  assign n90 = ~n84 & ~n89 ;
  assign n91 = ~n36 & n90 ;
  assign n92 = n91 ^ n90 ;
  assign n93 = n92 ^ n89 ;
  assign n94 = ~x0 & ~x8 ;
  assign n95 = ~n43 & ~n67 ;
  assign n96 = ~n94 & n95 ;
  assign n97 = ~n93 & n96 ;
  assign n98 = n97 ^ n96 ;
  assign n111 = n43 ^ x1 ;
  assign n112 = n111 ^ x9 ;
  assign n113 = n112 ^ x8 ;
  assign n114 = n112 ^ x0 ;
  assign n115 = ~n113 & ~n114 ;
  assign n116 = n115 ^ n112 ;
  assign n103 = x2 & ~n20 ;
  assign n104 = n103 ^ x2 ;
  assign n99 = x2 & n37 ;
  assign n100 = ~n29 & n99 ;
  assign n101 = ~n36 & n100 ;
  assign n102 = n101 ^ n100 ;
  assign n105 = n104 ^ n102 ;
  assign n106 = ~x0 & x1 ;
  assign n107 = ~x8 & x9 ;
  assign n108 = n106 & n107 ;
  assign n109 = x10 & n108 ;
  assign n110 = n105 & n109 ;
  assign n117 = n116 ^ n110 ;
  assign n118 = n98 & ~n117 ;
  assign n119 = n118 ^ n98 ;
  assign n120 = n119 ^ n117 ;
  assign n121 = n81 & n120 ;
  assign n122 = n121 ^ n81 ;
  assign n123 = n122 ^ n120 ;
  assign n124 = n105 ^ n66 ;
  assign n125 = n29 & n37 ;
  assign n126 = n125 ^ n37 ;
  assign n127 = ~n36 & n126 ;
  assign n128 = n127 ^ n126 ;
  assign n129 = n128 ^ n20 ;
  assign n130 = n129 ^ n17 ;
  assign n131 = n124 & ~n130 ;
  assign n132 = n131 ^ n124 ;
  assign n135 = x8 ^ x0 ;
  assign n137 = n135 ^ n43 ;
  assign n138 = n137 ^ n71 ;
  assign n133 = n66 & ~n86 ;
  assign n134 = n112 & ~n133 ;
  assign n136 = n135 ^ n134 ;
  assign n139 = n138 ^ n136 ;
  assign n140 = n132 & n139 ;
  assign n141 = n140 ^ n136 ;
  assign n145 = n86 ^ n66 ;
  assign n146 = ~n130 & n145 ;
  assign n143 = ~n71 & n130 ;
  assign n142 = ~n124 & n130 ;
  assign n144 = n143 ^ n142 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = n130 ^ n71 ;
  assign n149 = n48 & n49 ;
  assign n150 = ~n26 & ~n149 ;
  assign n151 = n28 & ~n150 ;
  assign n152 = ~n29 & ~n151 ;
  assign n153 = n31 & ~n152 ;
  assign n154 = n153 ^ n37 ;
  assign n155 = ~n23 & ~n57 ;
  assign n156 = n51 & ~n155 ;
  assign n157 = ~n22 & ~n156 ;
  assign n158 = n157 ^ n58 ;
  assign n159 = ~n23 & ~n149 ;
  assign n160 = n159 ^ n51 ;
  assign y0 = ~n123 ;
  assign y1 = n141 ;
  assign y2 = n147 ;
  assign y3 = n148 ;
  assign y4 = n154 ;
  assign y5 = ~n158 ;
  assign y6 = ~n160 ;
  assign y7 = n50 ;
endmodule
