module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 ;
  assign n437 = x40 ^ x16 ;
  assign n441 = x41 ^ x17 ;
  assign n442 = ~n437 & ~n441 ;
  assign n444 = x42 ^ x18 ;
  assign n450 = x43 ^ x19 ;
  assign n451 = ~n444 & ~n450 ;
  assign n452 = n442 & n451 ;
  assign n454 = x44 ^ x20 ;
  assign n458 = x45 ^ x21 ;
  assign n459 = ~n454 & ~n458 ;
  assign n461 = x46 ^ x22 ;
  assign n469 = x47 ^ x23 ;
  assign n470 = ~n461 & ~n469 ;
  assign n471 = n459 & n470 ;
  assign n472 = n452 & n471 ;
  assign n462 = x23 & ~x47 ;
  assign n463 = ~n461 & n462 ;
  assign n460 = x22 & ~x46 ;
  assign n464 = n463 ^ n460 ;
  assign n465 = n459 & n464 ;
  assign n455 = x21 & ~x45 ;
  assign n456 = ~n454 & n455 ;
  assign n453 = x20 & ~x44 ;
  assign n457 = n456 ^ n453 ;
  assign n466 = n465 ^ n457 ;
  assign n467 = n452 & n466 ;
  assign n445 = x19 & ~x43 ;
  assign n446 = ~n444 & n445 ;
  assign n443 = x18 & ~x42 ;
  assign n447 = n446 ^ n443 ;
  assign n448 = n442 & n447 ;
  assign n438 = x17 & ~x41 ;
  assign n439 = ~n437 & n438 ;
  assign n436 = x16 & ~x40 ;
  assign n440 = n439 ^ n436 ;
  assign n449 = n448 ^ n440 ;
  assign n468 = n467 ^ n449 ;
  assign n473 = n472 ^ n468 ;
  assign n262 = x40 ^ x8 ;
  assign n266 = x41 ^ x9 ;
  assign n267 = ~n262 & ~n266 ;
  assign n269 = x42 ^ x10 ;
  assign n275 = x43 ^ x11 ;
  assign n276 = ~n269 & ~n275 ;
  assign n277 = n267 & n276 ;
  assign n279 = x44 ^ x12 ;
  assign n283 = x45 ^ x13 ;
  assign n284 = ~n279 & ~n283 ;
  assign n286 = x46 ^ x14 ;
  assign n294 = x47 ^ x15 ;
  assign n295 = ~n286 & ~n294 ;
  assign n296 = n284 & n295 ;
  assign n297 = n277 & n296 ;
  assign n287 = x15 & ~x47 ;
  assign n288 = ~n286 & n287 ;
  assign n285 = x14 & ~x46 ;
  assign n289 = n288 ^ n285 ;
  assign n290 = n284 & n289 ;
  assign n280 = x13 & ~x45 ;
  assign n281 = ~n279 & n280 ;
  assign n278 = x12 & ~x44 ;
  assign n282 = n281 ^ n278 ;
  assign n291 = n290 ^ n282 ;
  assign n292 = n277 & n291 ;
  assign n270 = x11 & ~x43 ;
  assign n271 = ~n269 & n270 ;
  assign n268 = x10 & ~x42 ;
  assign n272 = n271 ^ n268 ;
  assign n273 = n267 & n272 ;
  assign n263 = x9 & ~x41 ;
  assign n264 = ~n262 & n263 ;
  assign n261 = x8 & ~x40 ;
  assign n265 = n264 ^ n261 ;
  assign n274 = n273 ^ n265 ;
  assign n293 = n292 ^ n274 ;
  assign n298 = n297 ^ n293 ;
  assign n736 = n473 ^ n298 ;
  assign n50 = x40 ^ x0 ;
  assign n54 = x41 ^ x1 ;
  assign n55 = ~n50 & ~n54 ;
  assign n57 = x42 ^ x2 ;
  assign n63 = x43 ^ x3 ;
  assign n64 = ~n57 & ~n63 ;
  assign n65 = n55 & n64 ;
  assign n67 = x44 ^ x4 ;
  assign n71 = x45 ^ x5 ;
  assign n72 = ~n67 & ~n71 ;
  assign n74 = x46 ^ x6 ;
  assign n82 = x47 ^ x7 ;
  assign n83 = ~n74 & ~n82 ;
  assign n84 = n72 & n83 ;
  assign n85 = n65 & n84 ;
  assign n75 = x7 & ~x47 ;
  assign n76 = ~n74 & n75 ;
  assign n73 = x6 & ~x46 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = n72 & n77 ;
  assign n68 = x5 & ~x45 ;
  assign n69 = ~n67 & n68 ;
  assign n66 = x4 & ~x44 ;
  assign n70 = n69 ^ n66 ;
  assign n79 = n78 ^ n70 ;
  assign n80 = n65 & n79 ;
  assign n58 = x3 & ~x43 ;
  assign n59 = ~n57 & n58 ;
  assign n56 = x2 & ~x42 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n55 & n60 ;
  assign n51 = x1 & ~x41 ;
  assign n52 = ~n50 & n51 ;
  assign n49 = x0 & ~x40 ;
  assign n53 = n52 ^ n49 ;
  assign n62 = n61 ^ n53 ;
  assign n81 = n80 ^ n62 ;
  assign n86 = n85 ^ n81 ;
  assign n741 = n736 ^ n86 ;
  assign n682 = x40 ^ x32 ;
  assign n686 = x41 ^ x33 ;
  assign n687 = ~n682 & ~n686 ;
  assign n689 = x42 ^ x34 ;
  assign n695 = x43 ^ x35 ;
  assign n696 = ~n689 & ~n695 ;
  assign n697 = n687 & n696 ;
  assign n699 = x44 ^ x36 ;
  assign n703 = x45 ^ x37 ;
  assign n704 = ~n699 & ~n703 ;
  assign n706 = x46 ^ x38 ;
  assign n714 = x47 ^ x39 ;
  assign n715 = ~n706 & ~n714 ;
  assign n716 = n704 & n715 ;
  assign n717 = n697 & n716 ;
  assign n707 = x39 & ~x47 ;
  assign n708 = ~n706 & n707 ;
  assign n705 = x38 & ~x46 ;
  assign n709 = n708 ^ n705 ;
  assign n710 = n704 & n709 ;
  assign n700 = x37 & ~x45 ;
  assign n701 = ~n699 & n700 ;
  assign n698 = x36 & ~x44 ;
  assign n702 = n701 ^ n698 ;
  assign n711 = n710 ^ n702 ;
  assign n712 = n697 & n711 ;
  assign n690 = x35 & ~x43 ;
  assign n691 = ~n689 & n690 ;
  assign n688 = x34 & ~x42 ;
  assign n692 = n691 ^ n688 ;
  assign n693 = n687 & n692 ;
  assign n683 = x33 & ~x41 ;
  assign n684 = ~n682 & n683 ;
  assign n681 = x32 & ~x40 ;
  assign n685 = n684 ^ n681 ;
  assign n694 = n693 ^ n685 ;
  assign n713 = n712 ^ n694 ;
  assign n718 = n717 ^ n713 ;
  assign n620 = x40 ^ x24 ;
  assign n624 = x41 ^ x25 ;
  assign n625 = ~n620 & ~n624 ;
  assign n627 = x42 ^ x26 ;
  assign n633 = x43 ^ x27 ;
  assign n634 = ~n627 & ~n633 ;
  assign n635 = n625 & n634 ;
  assign n637 = x44 ^ x28 ;
  assign n641 = x45 ^ x29 ;
  assign n642 = ~n637 & ~n641 ;
  assign n644 = x46 ^ x30 ;
  assign n652 = x47 ^ x31 ;
  assign n653 = ~n644 & ~n652 ;
  assign n654 = n642 & n653 ;
  assign n655 = n635 & n654 ;
  assign n645 = x31 & ~x47 ;
  assign n646 = ~n644 & n645 ;
  assign n643 = x30 & ~x46 ;
  assign n647 = n646 ^ n643 ;
  assign n648 = n642 & n647 ;
  assign n638 = x29 & ~x45 ;
  assign n639 = ~n637 & n638 ;
  assign n636 = x28 & ~x44 ;
  assign n640 = n639 ^ n636 ;
  assign n649 = n648 ^ n640 ;
  assign n650 = n635 & n649 ;
  assign n628 = x27 & ~x43 ;
  assign n629 = ~n627 & n628 ;
  assign n626 = x26 & ~x42 ;
  assign n630 = n629 ^ n626 ;
  assign n631 = n625 & n630 ;
  assign n621 = x25 & ~x41 ;
  assign n622 = ~n620 & n621 ;
  assign n619 = x24 & ~x40 ;
  assign n623 = n622 ^ n619 ;
  assign n632 = n631 ^ n623 ;
  assign n651 = n650 ^ n632 ;
  assign n656 = n655 ^ n651 ;
  assign n742 = n718 ^ n656 ;
  assign n743 = ~n741 & n742 ;
  assign n739 = ~n298 & ~n473 ;
  assign n737 = ~n86 & n736 ;
  assign n740 = n739 ^ n737 ;
  assign n744 = n743 ^ n740 ;
  assign n745 = ~n656 & ~n718 ;
  assign n746 = n745 ^ n743 ;
  assign n747 = n744 & n746 ;
  assign n748 = n747 ^ n743 ;
  assign n734 = ~n86 & ~n298 ;
  assign n733 = ~n86 & ~n473 ;
  assign n735 = n734 ^ n733 ;
  assign n738 = n737 ^ n735 ;
  assign n749 = n748 ^ n738 ;
  assign n750 = n745 ^ n744 ;
  assign n751 = n742 ^ n741 ;
  assign n752 = x40 & n751 ;
  assign n753 = ~n750 & n752 ;
  assign n754 = ~n749 & n753 ;
  assign n514 = x32 ^ x16 ;
  assign n518 = x33 ^ x17 ;
  assign n519 = ~n514 & ~n518 ;
  assign n521 = x34 ^ x18 ;
  assign n527 = x35 ^ x19 ;
  assign n528 = ~n521 & ~n527 ;
  assign n529 = n519 & n528 ;
  assign n531 = x36 ^ x20 ;
  assign n535 = x37 ^ x21 ;
  assign n536 = ~n531 & ~n535 ;
  assign n538 = x38 ^ x22 ;
  assign n546 = x39 ^ x23 ;
  assign n547 = ~n538 & ~n546 ;
  assign n548 = n536 & n547 ;
  assign n549 = n529 & n548 ;
  assign n539 = x23 & ~x39 ;
  assign n540 = ~n538 & n539 ;
  assign n537 = x22 & ~x38 ;
  assign n541 = n540 ^ n537 ;
  assign n542 = n536 & n541 ;
  assign n532 = x21 & ~x37 ;
  assign n533 = ~n531 & n532 ;
  assign n530 = x20 & ~x36 ;
  assign n534 = n533 ^ n530 ;
  assign n543 = n542 ^ n534 ;
  assign n544 = n529 & n543 ;
  assign n522 = x19 & ~x35 ;
  assign n523 = ~n521 & n522 ;
  assign n520 = x18 & ~x34 ;
  assign n524 = n523 ^ n520 ;
  assign n525 = n519 & n524 ;
  assign n515 = x17 & ~x33 ;
  assign n516 = ~n514 & n515 ;
  assign n513 = x16 & ~x32 ;
  assign n517 = n516 ^ n513 ;
  assign n526 = n525 ^ n517 ;
  assign n545 = n544 ^ n526 ;
  assign n550 = n549 ^ n545 ;
  assign n339 = x32 ^ x8 ;
  assign n343 = x33 ^ x9 ;
  assign n344 = ~n339 & ~n343 ;
  assign n346 = x34 ^ x10 ;
  assign n352 = x35 ^ x11 ;
  assign n353 = ~n346 & ~n352 ;
  assign n354 = n344 & n353 ;
  assign n356 = x36 ^ x12 ;
  assign n360 = x37 ^ x13 ;
  assign n361 = ~n356 & ~n360 ;
  assign n363 = x38 ^ x14 ;
  assign n371 = x39 ^ x15 ;
  assign n372 = ~n363 & ~n371 ;
  assign n373 = n361 & n372 ;
  assign n374 = n354 & n373 ;
  assign n364 = x15 & ~x39 ;
  assign n365 = ~n363 & n364 ;
  assign n362 = x14 & ~x38 ;
  assign n366 = n365 ^ n362 ;
  assign n367 = n361 & n366 ;
  assign n357 = x13 & ~x37 ;
  assign n358 = ~n356 & n357 ;
  assign n355 = x12 & ~x36 ;
  assign n359 = n358 ^ n355 ;
  assign n368 = n367 ^ n359 ;
  assign n369 = n354 & n368 ;
  assign n347 = x11 & ~x35 ;
  assign n348 = ~n346 & n347 ;
  assign n345 = x10 & ~x34 ;
  assign n349 = n348 ^ n345 ;
  assign n350 = n344 & n349 ;
  assign n340 = x9 & ~x33 ;
  assign n341 = ~n339 & n340 ;
  assign n338 = x8 & ~x32 ;
  assign n342 = n341 ^ n338 ;
  assign n351 = n350 ^ n342 ;
  assign n370 = n369 ^ n351 ;
  assign n375 = n374 ^ n370 ;
  assign n675 = n550 ^ n375 ;
  assign n127 = x32 ^ x0 ;
  assign n131 = x33 ^ x1 ;
  assign n132 = ~n127 & ~n131 ;
  assign n134 = x34 ^ x2 ;
  assign n140 = x35 ^ x3 ;
  assign n141 = ~n134 & ~n140 ;
  assign n142 = n132 & n141 ;
  assign n144 = x36 ^ x4 ;
  assign n148 = x37 ^ x5 ;
  assign n149 = ~n144 & ~n148 ;
  assign n151 = x38 ^ x6 ;
  assign n159 = x39 ^ x7 ;
  assign n160 = ~n151 & ~n159 ;
  assign n161 = n149 & n160 ;
  assign n162 = n142 & n161 ;
  assign n152 = x7 & ~x39 ;
  assign n153 = ~n151 & n152 ;
  assign n150 = x6 & ~x38 ;
  assign n154 = n153 ^ n150 ;
  assign n155 = n149 & n154 ;
  assign n145 = x5 & ~x37 ;
  assign n146 = ~n144 & n145 ;
  assign n143 = x4 & ~x36 ;
  assign n147 = n146 ^ n143 ;
  assign n156 = n155 ^ n147 ;
  assign n157 = n142 & n156 ;
  assign n135 = x3 & ~x35 ;
  assign n136 = ~n134 & n135 ;
  assign n133 = x2 & ~x34 ;
  assign n137 = n136 ^ n133 ;
  assign n138 = n132 & n137 ;
  assign n128 = x1 & ~x33 ;
  assign n129 = ~n127 & n128 ;
  assign n126 = x0 & ~x32 ;
  assign n130 = n129 ^ n126 ;
  assign n139 = n138 ^ n130 ;
  assign n158 = n157 ^ n139 ;
  assign n163 = n162 ^ n158 ;
  assign n680 = n675 ^ n163 ;
  assign n582 = x32 ^ x24 ;
  assign n586 = x33 ^ x25 ;
  assign n587 = ~n582 & ~n586 ;
  assign n589 = x34 ^ x26 ;
  assign n595 = x35 ^ x27 ;
  assign n596 = ~n589 & ~n595 ;
  assign n597 = n587 & n596 ;
  assign n599 = x36 ^ x28 ;
  assign n603 = x37 ^ x29 ;
  assign n604 = ~n599 & ~n603 ;
  assign n606 = x38 ^ x30 ;
  assign n614 = x39 ^ x31 ;
  assign n615 = ~n606 & ~n614 ;
  assign n616 = n604 & n615 ;
  assign n617 = n597 & n616 ;
  assign n607 = x31 & ~x39 ;
  assign n608 = ~n606 & n607 ;
  assign n605 = x30 & ~x38 ;
  assign n609 = n608 ^ n605 ;
  assign n610 = n604 & n609 ;
  assign n600 = x29 & ~x37 ;
  assign n601 = ~n599 & n600 ;
  assign n598 = x28 & ~x36 ;
  assign n602 = n601 ^ n598 ;
  assign n611 = n610 ^ n602 ;
  assign n612 = n597 & n611 ;
  assign n590 = x27 & ~x35 ;
  assign n591 = ~n589 & n590 ;
  assign n588 = x26 & ~x34 ;
  assign n592 = n591 ^ n588 ;
  assign n593 = n587 & n592 ;
  assign n583 = x25 & ~x33 ;
  assign n584 = ~n582 & n583 ;
  assign n581 = x24 & ~x32 ;
  assign n585 = n584 ^ n581 ;
  assign n594 = n593 ^ n585 ;
  assign n613 = n612 ^ n594 ;
  assign n618 = n617 ^ n613 ;
  assign n719 = n718 ^ n618 ;
  assign n720 = ~n680 & ~n719 ;
  assign n678 = ~n375 & ~n550 ;
  assign n676 = ~n163 & n675 ;
  assign n679 = n678 ^ n676 ;
  assign n721 = n720 ^ n679 ;
  assign n722 = ~n618 & n718 ;
  assign n723 = n722 ^ n720 ;
  assign n724 = n721 & n723 ;
  assign n725 = n724 ^ n720 ;
  assign n673 = ~n163 & ~n375 ;
  assign n672 = ~n163 & ~n550 ;
  assign n674 = n673 ^ n672 ;
  assign n677 = n676 ^ n674 ;
  assign n726 = n725 ^ n677 ;
  assign n727 = n722 ^ n721 ;
  assign n728 = n719 ^ n680 ;
  assign n729 = x32 & ~n728 ;
  assign n730 = ~n727 & n729 ;
  assign n731 = ~n726 & n730 ;
  assign n657 = n656 ^ n618 ;
  assign n475 = x24 ^ x16 ;
  assign n479 = x25 ^ x17 ;
  assign n480 = ~n475 & ~n479 ;
  assign n482 = x26 ^ x18 ;
  assign n488 = x27 ^ x19 ;
  assign n489 = ~n482 & ~n488 ;
  assign n490 = n480 & n489 ;
  assign n492 = x28 ^ x20 ;
  assign n496 = x29 ^ x21 ;
  assign n497 = ~n492 & ~n496 ;
  assign n499 = x30 ^ x22 ;
  assign n507 = x31 ^ x23 ;
  assign n508 = ~n499 & ~n507 ;
  assign n509 = n497 & n508 ;
  assign n510 = n490 & n509 ;
  assign n500 = x23 & ~x31 ;
  assign n501 = ~n499 & n500 ;
  assign n498 = x22 & ~x30 ;
  assign n502 = n501 ^ n498 ;
  assign n503 = n497 & n502 ;
  assign n493 = x21 & ~x29 ;
  assign n494 = ~n492 & n493 ;
  assign n491 = x20 & ~x28 ;
  assign n495 = n494 ^ n491 ;
  assign n504 = n503 ^ n495 ;
  assign n505 = n490 & n504 ;
  assign n483 = x19 & ~x27 ;
  assign n484 = ~n482 & n483 ;
  assign n481 = x18 & ~x26 ;
  assign n485 = n484 ^ n481 ;
  assign n486 = n480 & n485 ;
  assign n476 = x17 & ~x25 ;
  assign n477 = ~n475 & n476 ;
  assign n474 = x16 & ~x24 ;
  assign n478 = n477 ^ n474 ;
  assign n487 = n486 ^ n478 ;
  assign n506 = n505 ^ n487 ;
  assign n511 = n510 ^ n506 ;
  assign n300 = x24 ^ x8 ;
  assign n304 = x25 ^ x9 ;
  assign n305 = ~n300 & ~n304 ;
  assign n307 = x26 ^ x10 ;
  assign n313 = x27 ^ x11 ;
  assign n314 = ~n307 & ~n313 ;
  assign n315 = n305 & n314 ;
  assign n317 = x28 ^ x12 ;
  assign n321 = x29 ^ x13 ;
  assign n322 = ~n317 & ~n321 ;
  assign n324 = x30 ^ x14 ;
  assign n332 = x31 ^ x15 ;
  assign n333 = ~n324 & ~n332 ;
  assign n334 = n322 & n333 ;
  assign n335 = n315 & n334 ;
  assign n325 = x15 & ~x31 ;
  assign n326 = ~n324 & n325 ;
  assign n323 = x14 & ~x30 ;
  assign n327 = n326 ^ n323 ;
  assign n328 = n322 & n327 ;
  assign n318 = x13 & ~x29 ;
  assign n319 = ~n317 & n318 ;
  assign n316 = x12 & ~x28 ;
  assign n320 = n319 ^ n316 ;
  assign n329 = n328 ^ n320 ;
  assign n330 = n315 & n329 ;
  assign n308 = x11 & ~x27 ;
  assign n309 = ~n307 & n308 ;
  assign n306 = x10 & ~x26 ;
  assign n310 = n309 ^ n306 ;
  assign n311 = n305 & n310 ;
  assign n301 = x9 & ~x25 ;
  assign n302 = ~n300 & n301 ;
  assign n299 = x8 & ~x24 ;
  assign n303 = n302 ^ n299 ;
  assign n312 = n311 ^ n303 ;
  assign n331 = n330 ^ n312 ;
  assign n336 = n335 ^ n331 ;
  assign n576 = n511 ^ n336 ;
  assign n88 = x24 ^ x0 ;
  assign n92 = x25 ^ x1 ;
  assign n93 = ~n88 & ~n92 ;
  assign n95 = x26 ^ x2 ;
  assign n101 = x27 ^ x3 ;
  assign n102 = ~n95 & ~n101 ;
  assign n103 = n93 & n102 ;
  assign n105 = x28 ^ x4 ;
  assign n109 = x29 ^ x5 ;
  assign n110 = ~n105 & ~n109 ;
  assign n112 = x30 ^ x6 ;
  assign n120 = x31 ^ x7 ;
  assign n121 = ~n112 & ~n120 ;
  assign n122 = n110 & n121 ;
  assign n123 = n103 & n122 ;
  assign n113 = x7 & ~x31 ;
  assign n114 = ~n112 & n113 ;
  assign n111 = x6 & ~x30 ;
  assign n115 = n114 ^ n111 ;
  assign n116 = n110 & n115 ;
  assign n106 = x5 & ~x29 ;
  assign n107 = ~n105 & n106 ;
  assign n104 = x4 & ~x28 ;
  assign n108 = n107 ^ n104 ;
  assign n117 = n116 ^ n108 ;
  assign n118 = n103 & n117 ;
  assign n96 = x3 & ~x27 ;
  assign n97 = ~n95 & n96 ;
  assign n94 = x2 & ~x26 ;
  assign n98 = n97 ^ n94 ;
  assign n99 = n93 & n98 ;
  assign n89 = x1 & ~x25 ;
  assign n90 = ~n88 & n89 ;
  assign n87 = x0 & ~x24 ;
  assign n91 = n90 ^ n87 ;
  assign n100 = n99 ^ n91 ;
  assign n119 = n118 ^ n100 ;
  assign n124 = n123 ^ n119 ;
  assign n658 = n576 ^ n124 ;
  assign n659 = n657 & ~n658 ;
  assign n579 = ~n336 & ~n511 ;
  assign n577 = ~n124 & n576 ;
  assign n580 = n579 ^ n577 ;
  assign n660 = n659 ^ n580 ;
  assign n661 = n618 & n656 ;
  assign n662 = n661 ^ n659 ;
  assign n663 = n660 & n662 ;
  assign n664 = n663 ^ n659 ;
  assign n574 = ~n124 & ~n336 ;
  assign n573 = ~n124 & ~n511 ;
  assign n575 = n574 ^ n573 ;
  assign n578 = n577 ^ n575 ;
  assign n665 = n664 ^ n578 ;
  assign n666 = n661 ^ n660 ;
  assign n667 = n658 ^ n657 ;
  assign n668 = x24 & n667 ;
  assign n669 = ~n666 & n668 ;
  assign n670 = ~n665 & n669 ;
  assign n208 = x16 ^ x0 ;
  assign n212 = x17 ^ x1 ;
  assign n213 = ~n208 & ~n212 ;
  assign n215 = x18 ^ x2 ;
  assign n221 = x19 ^ x3 ;
  assign n222 = ~n215 & ~n221 ;
  assign n223 = n213 & n222 ;
  assign n225 = x20 ^ x4 ;
  assign n229 = x21 ^ x5 ;
  assign n230 = ~n225 & ~n229 ;
  assign n232 = x22 ^ x6 ;
  assign n240 = x23 ^ x7 ;
  assign n241 = ~n232 & ~n240 ;
  assign n242 = n230 & n241 ;
  assign n243 = n223 & n242 ;
  assign n233 = x7 & ~x23 ;
  assign n234 = ~n232 & n233 ;
  assign n231 = x6 & ~x22 ;
  assign n235 = n234 ^ n231 ;
  assign n236 = n230 & n235 ;
  assign n226 = x5 & ~x21 ;
  assign n227 = ~n225 & n226 ;
  assign n224 = x4 & ~x20 ;
  assign n228 = n227 ^ n224 ;
  assign n237 = n236 ^ n228 ;
  assign n238 = n223 & n237 ;
  assign n216 = x3 & ~x19 ;
  assign n217 = ~n215 & n216 ;
  assign n214 = x2 & ~x18 ;
  assign n218 = n217 ^ n214 ;
  assign n219 = n213 & n218 ;
  assign n209 = x1 & ~x17 ;
  assign n210 = ~n208 & n209 ;
  assign n207 = x0 & ~x16 ;
  assign n211 = n210 ^ n207 ;
  assign n220 = n219 ^ n211 ;
  assign n239 = n238 ^ n220 ;
  assign n244 = n243 ^ n239 ;
  assign n382 = x16 ^ x8 ;
  assign n386 = x17 ^ x9 ;
  assign n387 = ~n382 & ~n386 ;
  assign n389 = x18 ^ x10 ;
  assign n395 = x19 ^ x11 ;
  assign n396 = ~n389 & ~n395 ;
  assign n397 = n387 & n396 ;
  assign n399 = x20 ^ x12 ;
  assign n403 = x21 ^ x13 ;
  assign n404 = ~n399 & ~n403 ;
  assign n406 = x22 ^ x14 ;
  assign n414 = x23 ^ x15 ;
  assign n415 = ~n406 & ~n414 ;
  assign n416 = n404 & n415 ;
  assign n417 = n397 & n416 ;
  assign n407 = x15 & ~x23 ;
  assign n408 = ~n406 & n407 ;
  assign n405 = x14 & ~x22 ;
  assign n409 = n408 ^ n405 ;
  assign n410 = n404 & n409 ;
  assign n400 = x13 & ~x21 ;
  assign n401 = ~n399 & n400 ;
  assign n398 = x12 & ~x20 ;
  assign n402 = n401 ^ n398 ;
  assign n411 = n410 ^ n402 ;
  assign n412 = n397 & n411 ;
  assign n390 = x11 & ~x19 ;
  assign n391 = ~n389 & n390 ;
  assign n388 = x10 & ~x18 ;
  assign n392 = n391 ^ n388 ;
  assign n393 = n387 & n392 ;
  assign n383 = x9 & ~x17 ;
  assign n384 = ~n382 & n383 ;
  assign n381 = x8 & ~x16 ;
  assign n385 = n384 ^ n381 ;
  assign n394 = n393 ^ n385 ;
  assign n413 = n412 ^ n394 ;
  assign n418 = n417 ^ n413 ;
  assign n559 = ~n244 & ~n418 ;
  assign n556 = n418 ^ n244 ;
  assign n553 = n550 ^ n473 ;
  assign n557 = n553 ^ n511 ;
  assign n558 = n556 & n557 ;
  assign n560 = n559 ^ n558 ;
  assign n561 = n473 & n550 ;
  assign n554 = n511 & n553 ;
  assign n562 = n561 ^ n554 ;
  assign n563 = n562 ^ n558 ;
  assign n564 = n560 & n563 ;
  assign n565 = n564 ^ n558 ;
  assign n551 = n511 & ~n550 ;
  assign n512 = ~n473 & n511 ;
  assign n552 = n551 ^ n512 ;
  assign n555 = n554 ^ n552 ;
  assign n566 = n565 ^ n555 ;
  assign n567 = n562 ^ n560 ;
  assign n568 = n557 ^ n556 ;
  assign n569 = x16 & ~n568 ;
  assign n570 = ~n567 & n569 ;
  assign n571 = ~n566 & n570 ;
  assign n170 = x8 ^ x0 ;
  assign n174 = x9 ^ x1 ;
  assign n175 = ~n170 & ~n174 ;
  assign n177 = x10 ^ x2 ;
  assign n183 = x11 ^ x3 ;
  assign n184 = ~n177 & ~n183 ;
  assign n185 = n175 & n184 ;
  assign n187 = x12 ^ x4 ;
  assign n191 = x13 ^ x5 ;
  assign n192 = ~n187 & ~n191 ;
  assign n194 = x14 ^ x6 ;
  assign n202 = x15 ^ x7 ;
  assign n203 = ~n194 & ~n202 ;
  assign n204 = n192 & n203 ;
  assign n205 = n185 & n204 ;
  assign n195 = x7 & ~x15 ;
  assign n196 = ~n194 & n195 ;
  assign n193 = x6 & ~x14 ;
  assign n197 = n196 ^ n193 ;
  assign n198 = n192 & n197 ;
  assign n188 = x5 & ~x13 ;
  assign n189 = ~n187 & n188 ;
  assign n186 = x4 & ~x12 ;
  assign n190 = n189 ^ n186 ;
  assign n199 = n198 ^ n190 ;
  assign n200 = n185 & n199 ;
  assign n178 = x3 & ~x11 ;
  assign n179 = ~n177 & n178 ;
  assign n176 = x2 & ~x10 ;
  assign n180 = n179 ^ n176 ;
  assign n181 = n175 & n180 ;
  assign n171 = x1 & ~x9 ;
  assign n172 = ~n170 & n171 ;
  assign n169 = x0 & ~x8 ;
  assign n173 = n172 ^ n169 ;
  assign n182 = n181 ^ n173 ;
  assign n201 = n200 ^ n182 ;
  assign n206 = n205 ^ n201 ;
  assign n422 = ~n206 & n418 ;
  assign n419 = n418 ^ n206 ;
  assign n378 = n375 ^ n298 ;
  assign n420 = n378 ^ n336 ;
  assign n421 = ~n419 & n420 ;
  assign n423 = n422 ^ n421 ;
  assign n424 = n298 & n375 ;
  assign n379 = n336 & n378 ;
  assign n425 = n424 ^ n379 ;
  assign n426 = n425 ^ n421 ;
  assign n427 = n423 & n426 ;
  assign n428 = n427 ^ n421 ;
  assign n376 = n336 & ~n375 ;
  assign n337 = ~n298 & n336 ;
  assign n377 = n376 ^ n337 ;
  assign n380 = n379 ^ n377 ;
  assign n429 = n428 ^ n380 ;
  assign n430 = n425 ^ n423 ;
  assign n431 = n420 ^ n419 ;
  assign n432 = x8 & n431 ;
  assign n433 = ~n430 & n432 ;
  assign n434 = ~n429 & n433 ;
  assign n248 = n206 & n244 ;
  assign n245 = n244 ^ n206 ;
  assign n166 = n163 ^ n86 ;
  assign n246 = n166 ^ n124 ;
  assign n247 = n245 & n246 ;
  assign n249 = n248 ^ n247 ;
  assign n250 = n86 & n163 ;
  assign n167 = n124 & n166 ;
  assign n251 = n250 ^ n167 ;
  assign n252 = n251 ^ n247 ;
  assign n253 = n249 & n252 ;
  assign n254 = n253 ^ n247 ;
  assign n164 = n124 & ~n163 ;
  assign n125 = ~n86 & n124 ;
  assign n165 = n164 ^ n125 ;
  assign n168 = n167 ^ n165 ;
  assign n255 = n254 ^ n168 ;
  assign n256 = n251 ^ n249 ;
  assign n257 = n246 ^ n245 ;
  assign n258 = x0 & ~n257 ;
  assign n259 = ~n256 & n258 ;
  assign n260 = ~n255 & n259 ;
  assign n435 = n434 ^ n260 ;
  assign n572 = n571 ^ n435 ;
  assign n671 = n670 ^ n572 ;
  assign n732 = n731 ^ n671 ;
  assign n755 = n754 ^ n732 ;
  assign n775 = x41 & n751 ;
  assign n776 = ~n750 & n775 ;
  assign n777 = ~n749 & n776 ;
  assign n771 = x33 & ~n728 ;
  assign n772 = ~n727 & n771 ;
  assign n773 = ~n726 & n772 ;
  assign n767 = x25 & n667 ;
  assign n768 = ~n666 & n767 ;
  assign n769 = ~n665 & n768 ;
  assign n763 = x17 & ~n568 ;
  assign n764 = ~n567 & n763 ;
  assign n765 = ~n566 & n764 ;
  assign n759 = x9 & n431 ;
  assign n760 = ~n430 & n759 ;
  assign n761 = ~n429 & n760 ;
  assign n756 = x1 & ~n257 ;
  assign n757 = ~n256 & n756 ;
  assign n758 = ~n255 & n757 ;
  assign n762 = n761 ^ n758 ;
  assign n766 = n765 ^ n762 ;
  assign n770 = n769 ^ n766 ;
  assign n774 = n773 ^ n770 ;
  assign n778 = n777 ^ n774 ;
  assign n798 = x42 & n751 ;
  assign n799 = ~n750 & n798 ;
  assign n800 = ~n749 & n799 ;
  assign n794 = x34 & ~n728 ;
  assign n795 = ~n727 & n794 ;
  assign n796 = ~n726 & n795 ;
  assign n790 = x26 & n667 ;
  assign n791 = ~n666 & n790 ;
  assign n792 = ~n665 & n791 ;
  assign n786 = x18 & ~n568 ;
  assign n787 = ~n567 & n786 ;
  assign n788 = ~n566 & n787 ;
  assign n782 = x10 & n431 ;
  assign n783 = ~n430 & n782 ;
  assign n784 = ~n429 & n783 ;
  assign n779 = x2 & ~n257 ;
  assign n780 = ~n256 & n779 ;
  assign n781 = ~n255 & n780 ;
  assign n785 = n784 ^ n781 ;
  assign n789 = n788 ^ n785 ;
  assign n793 = n792 ^ n789 ;
  assign n797 = n796 ^ n793 ;
  assign n801 = n800 ^ n797 ;
  assign n821 = x43 & n751 ;
  assign n822 = ~n750 & n821 ;
  assign n823 = ~n749 & n822 ;
  assign n817 = x35 & ~n728 ;
  assign n818 = ~n727 & n817 ;
  assign n819 = ~n726 & n818 ;
  assign n813 = x27 & n667 ;
  assign n814 = ~n666 & n813 ;
  assign n815 = ~n665 & n814 ;
  assign n809 = x19 & ~n568 ;
  assign n810 = ~n567 & n809 ;
  assign n811 = ~n566 & n810 ;
  assign n805 = x11 & n431 ;
  assign n806 = ~n430 & n805 ;
  assign n807 = ~n429 & n806 ;
  assign n802 = x3 & ~n257 ;
  assign n803 = ~n256 & n802 ;
  assign n804 = ~n255 & n803 ;
  assign n808 = n807 ^ n804 ;
  assign n812 = n811 ^ n808 ;
  assign n816 = n815 ^ n812 ;
  assign n820 = n819 ^ n816 ;
  assign n824 = n823 ^ n820 ;
  assign n844 = x44 & n751 ;
  assign n845 = ~n750 & n844 ;
  assign n846 = ~n749 & n845 ;
  assign n840 = x36 & ~n728 ;
  assign n841 = ~n727 & n840 ;
  assign n842 = ~n726 & n841 ;
  assign n836 = x28 & n667 ;
  assign n837 = ~n666 & n836 ;
  assign n838 = ~n665 & n837 ;
  assign n832 = x20 & ~n568 ;
  assign n833 = ~n567 & n832 ;
  assign n834 = ~n566 & n833 ;
  assign n828 = x12 & n431 ;
  assign n829 = ~n430 & n828 ;
  assign n830 = ~n429 & n829 ;
  assign n825 = x4 & ~n257 ;
  assign n826 = ~n256 & n825 ;
  assign n827 = ~n255 & n826 ;
  assign n831 = n830 ^ n827 ;
  assign n835 = n834 ^ n831 ;
  assign n839 = n838 ^ n835 ;
  assign n843 = n842 ^ n839 ;
  assign n847 = n846 ^ n843 ;
  assign n867 = x45 & n751 ;
  assign n868 = ~n750 & n867 ;
  assign n869 = ~n749 & n868 ;
  assign n863 = x37 & ~n728 ;
  assign n864 = ~n727 & n863 ;
  assign n865 = ~n726 & n864 ;
  assign n859 = x29 & n667 ;
  assign n860 = ~n666 & n859 ;
  assign n861 = ~n665 & n860 ;
  assign n855 = x21 & ~n568 ;
  assign n856 = ~n567 & n855 ;
  assign n857 = ~n566 & n856 ;
  assign n851 = x13 & n431 ;
  assign n852 = ~n430 & n851 ;
  assign n853 = ~n429 & n852 ;
  assign n848 = x5 & ~n257 ;
  assign n849 = ~n256 & n848 ;
  assign n850 = ~n255 & n849 ;
  assign n854 = n853 ^ n850 ;
  assign n858 = n857 ^ n854 ;
  assign n862 = n861 ^ n858 ;
  assign n866 = n865 ^ n862 ;
  assign n870 = n869 ^ n866 ;
  assign n890 = x46 & n751 ;
  assign n891 = ~n750 & n890 ;
  assign n892 = ~n749 & n891 ;
  assign n886 = x38 & ~n728 ;
  assign n887 = ~n727 & n886 ;
  assign n888 = ~n726 & n887 ;
  assign n882 = x30 & n667 ;
  assign n883 = ~n666 & n882 ;
  assign n884 = ~n665 & n883 ;
  assign n878 = x22 & ~n568 ;
  assign n879 = ~n567 & n878 ;
  assign n880 = ~n566 & n879 ;
  assign n874 = x14 & n431 ;
  assign n875 = ~n430 & n874 ;
  assign n876 = ~n429 & n875 ;
  assign n871 = x6 & ~n257 ;
  assign n872 = ~n256 & n871 ;
  assign n873 = ~n255 & n872 ;
  assign n877 = n876 ^ n873 ;
  assign n881 = n880 ^ n877 ;
  assign n885 = n884 ^ n881 ;
  assign n889 = n888 ^ n885 ;
  assign n893 = n892 ^ n889 ;
  assign n913 = x47 & n751 ;
  assign n914 = ~n750 & n913 ;
  assign n915 = ~n749 & n914 ;
  assign n909 = x39 & ~n728 ;
  assign n910 = ~n727 & n909 ;
  assign n911 = ~n726 & n910 ;
  assign n905 = x31 & n667 ;
  assign n906 = ~n666 & n905 ;
  assign n907 = ~n665 & n906 ;
  assign n901 = x23 & ~n568 ;
  assign n902 = ~n567 & n901 ;
  assign n903 = ~n566 & n902 ;
  assign n897 = x15 & n431 ;
  assign n898 = ~n430 & n897 ;
  assign n899 = ~n429 & n898 ;
  assign n894 = x7 & ~n257 ;
  assign n895 = ~n256 & n894 ;
  assign n896 = ~n255 & n895 ;
  assign n900 = n899 ^ n896 ;
  assign n904 = n903 ^ n900 ;
  assign n908 = n907 ^ n904 ;
  assign n912 = n911 ^ n908 ;
  assign n916 = n915 ^ n912 ;
  assign n936 = x40 & ~n751 ;
  assign n937 = ~n750 & n936 ;
  assign n938 = ~n749 & n937 ;
  assign n932 = x32 & n728 ;
  assign n933 = ~n727 & n932 ;
  assign n934 = ~n726 & n933 ;
  assign n928 = x24 & ~n667 ;
  assign n929 = ~n666 & n928 ;
  assign n930 = ~n665 & n929 ;
  assign n924 = x16 & n568 ;
  assign n925 = ~n567 & n924 ;
  assign n926 = ~n566 & n925 ;
  assign n920 = x8 & ~n431 ;
  assign n921 = ~n430 & n920 ;
  assign n922 = ~n429 & n921 ;
  assign n917 = x0 & n257 ;
  assign n918 = ~n256 & n917 ;
  assign n919 = ~n255 & n918 ;
  assign n923 = n922 ^ n919 ;
  assign n927 = n926 ^ n923 ;
  assign n931 = n930 ^ n927 ;
  assign n935 = n934 ^ n931 ;
  assign n939 = n938 ^ n935 ;
  assign n959 = x41 & ~n751 ;
  assign n960 = ~n750 & n959 ;
  assign n961 = ~n749 & n960 ;
  assign n955 = x33 & n728 ;
  assign n956 = ~n727 & n955 ;
  assign n957 = ~n726 & n956 ;
  assign n951 = x25 & ~n667 ;
  assign n952 = ~n666 & n951 ;
  assign n953 = ~n665 & n952 ;
  assign n947 = x17 & n568 ;
  assign n948 = ~n567 & n947 ;
  assign n949 = ~n566 & n948 ;
  assign n943 = x9 & ~n431 ;
  assign n944 = ~n430 & n943 ;
  assign n945 = ~n429 & n944 ;
  assign n940 = x1 & n257 ;
  assign n941 = ~n256 & n940 ;
  assign n942 = ~n255 & n941 ;
  assign n946 = n945 ^ n942 ;
  assign n950 = n949 ^ n946 ;
  assign n954 = n953 ^ n950 ;
  assign n958 = n957 ^ n954 ;
  assign n962 = n961 ^ n958 ;
  assign n982 = x42 & ~n751 ;
  assign n983 = ~n750 & n982 ;
  assign n984 = ~n749 & n983 ;
  assign n978 = x34 & n728 ;
  assign n979 = ~n727 & n978 ;
  assign n980 = ~n726 & n979 ;
  assign n974 = x26 & ~n667 ;
  assign n975 = ~n666 & n974 ;
  assign n976 = ~n665 & n975 ;
  assign n970 = x18 & n568 ;
  assign n971 = ~n567 & n970 ;
  assign n972 = ~n566 & n971 ;
  assign n966 = x10 & ~n431 ;
  assign n967 = ~n430 & n966 ;
  assign n968 = ~n429 & n967 ;
  assign n963 = x2 & n257 ;
  assign n964 = ~n256 & n963 ;
  assign n965 = ~n255 & n964 ;
  assign n969 = n968 ^ n965 ;
  assign n973 = n972 ^ n969 ;
  assign n977 = n976 ^ n973 ;
  assign n981 = n980 ^ n977 ;
  assign n985 = n984 ^ n981 ;
  assign n1005 = x43 & ~n751 ;
  assign n1006 = ~n750 & n1005 ;
  assign n1007 = ~n749 & n1006 ;
  assign n1001 = x35 & n728 ;
  assign n1002 = ~n727 & n1001 ;
  assign n1003 = ~n726 & n1002 ;
  assign n997 = x27 & ~n667 ;
  assign n998 = ~n666 & n997 ;
  assign n999 = ~n665 & n998 ;
  assign n993 = x19 & n568 ;
  assign n994 = ~n567 & n993 ;
  assign n995 = ~n566 & n994 ;
  assign n989 = x11 & ~n431 ;
  assign n990 = ~n430 & n989 ;
  assign n991 = ~n429 & n990 ;
  assign n986 = x3 & n257 ;
  assign n987 = ~n256 & n986 ;
  assign n988 = ~n255 & n987 ;
  assign n992 = n991 ^ n988 ;
  assign n996 = n995 ^ n992 ;
  assign n1000 = n999 ^ n996 ;
  assign n1004 = n1003 ^ n1000 ;
  assign n1008 = n1007 ^ n1004 ;
  assign n1028 = x44 & ~n751 ;
  assign n1029 = ~n750 & n1028 ;
  assign n1030 = ~n749 & n1029 ;
  assign n1024 = x36 & n728 ;
  assign n1025 = ~n727 & n1024 ;
  assign n1026 = ~n726 & n1025 ;
  assign n1020 = x28 & ~n667 ;
  assign n1021 = ~n666 & n1020 ;
  assign n1022 = ~n665 & n1021 ;
  assign n1016 = x20 & n568 ;
  assign n1017 = ~n567 & n1016 ;
  assign n1018 = ~n566 & n1017 ;
  assign n1012 = x12 & ~n431 ;
  assign n1013 = ~n430 & n1012 ;
  assign n1014 = ~n429 & n1013 ;
  assign n1009 = x4 & n257 ;
  assign n1010 = ~n256 & n1009 ;
  assign n1011 = ~n255 & n1010 ;
  assign n1015 = n1014 ^ n1011 ;
  assign n1019 = n1018 ^ n1015 ;
  assign n1023 = n1022 ^ n1019 ;
  assign n1027 = n1026 ^ n1023 ;
  assign n1031 = n1030 ^ n1027 ;
  assign n1051 = x45 & ~n751 ;
  assign n1052 = ~n750 & n1051 ;
  assign n1053 = ~n749 & n1052 ;
  assign n1047 = x37 & n728 ;
  assign n1048 = ~n727 & n1047 ;
  assign n1049 = ~n726 & n1048 ;
  assign n1043 = x29 & ~n667 ;
  assign n1044 = ~n666 & n1043 ;
  assign n1045 = ~n665 & n1044 ;
  assign n1039 = x21 & n568 ;
  assign n1040 = ~n567 & n1039 ;
  assign n1041 = ~n566 & n1040 ;
  assign n1035 = x13 & ~n431 ;
  assign n1036 = ~n430 & n1035 ;
  assign n1037 = ~n429 & n1036 ;
  assign n1032 = x5 & n257 ;
  assign n1033 = ~n256 & n1032 ;
  assign n1034 = ~n255 & n1033 ;
  assign n1038 = n1037 ^ n1034 ;
  assign n1042 = n1041 ^ n1038 ;
  assign n1046 = n1045 ^ n1042 ;
  assign n1050 = n1049 ^ n1046 ;
  assign n1054 = n1053 ^ n1050 ;
  assign n1074 = x46 & ~n751 ;
  assign n1075 = ~n750 & n1074 ;
  assign n1076 = ~n749 & n1075 ;
  assign n1070 = x38 & n728 ;
  assign n1071 = ~n727 & n1070 ;
  assign n1072 = ~n726 & n1071 ;
  assign n1066 = x30 & ~n667 ;
  assign n1067 = ~n666 & n1066 ;
  assign n1068 = ~n665 & n1067 ;
  assign n1062 = x22 & n568 ;
  assign n1063 = ~n567 & n1062 ;
  assign n1064 = ~n566 & n1063 ;
  assign n1058 = x14 & ~n431 ;
  assign n1059 = ~n430 & n1058 ;
  assign n1060 = ~n429 & n1059 ;
  assign n1055 = x6 & n257 ;
  assign n1056 = ~n256 & n1055 ;
  assign n1057 = ~n255 & n1056 ;
  assign n1061 = n1060 ^ n1057 ;
  assign n1065 = n1064 ^ n1061 ;
  assign n1069 = n1068 ^ n1065 ;
  assign n1073 = n1072 ^ n1069 ;
  assign n1077 = n1076 ^ n1073 ;
  assign n1097 = x47 & ~n751 ;
  assign n1098 = ~n750 & n1097 ;
  assign n1099 = ~n749 & n1098 ;
  assign n1093 = x39 & n728 ;
  assign n1094 = ~n727 & n1093 ;
  assign n1095 = ~n726 & n1094 ;
  assign n1089 = x31 & ~n667 ;
  assign n1090 = ~n666 & n1089 ;
  assign n1091 = ~n665 & n1090 ;
  assign n1085 = x23 & n568 ;
  assign n1086 = ~n567 & n1085 ;
  assign n1087 = ~n566 & n1086 ;
  assign n1081 = x15 & ~n431 ;
  assign n1082 = ~n430 & n1081 ;
  assign n1083 = ~n429 & n1082 ;
  assign n1078 = x7 & n257 ;
  assign n1079 = ~n256 & n1078 ;
  assign n1080 = ~n255 & n1079 ;
  assign n1084 = n1083 ^ n1080 ;
  assign n1088 = n1087 ^ n1084 ;
  assign n1092 = n1091 ^ n1088 ;
  assign n1096 = n1095 ^ n1092 ;
  assign n1100 = n1099 ^ n1096 ;
  assign n1115 = n750 & n752 ;
  assign n1116 = ~n749 & n1115 ;
  assign n1112 = n727 & n729 ;
  assign n1113 = ~n726 & n1112 ;
  assign n1109 = n666 & n668 ;
  assign n1110 = ~n665 & n1109 ;
  assign n1106 = n567 & n569 ;
  assign n1107 = ~n566 & n1106 ;
  assign n1103 = n430 & n432 ;
  assign n1104 = ~n429 & n1103 ;
  assign n1101 = n256 & n258 ;
  assign n1102 = ~n255 & n1101 ;
  assign n1105 = n1104 ^ n1102 ;
  assign n1108 = n1107 ^ n1105 ;
  assign n1111 = n1110 ^ n1108 ;
  assign n1114 = n1113 ^ n1111 ;
  assign n1117 = n1116 ^ n1114 ;
  assign n1132 = n750 & n775 ;
  assign n1133 = ~n749 & n1132 ;
  assign n1129 = n727 & n771 ;
  assign n1130 = ~n726 & n1129 ;
  assign n1126 = n666 & n767 ;
  assign n1127 = ~n665 & n1126 ;
  assign n1123 = n567 & n763 ;
  assign n1124 = ~n566 & n1123 ;
  assign n1120 = n430 & n759 ;
  assign n1121 = ~n429 & n1120 ;
  assign n1118 = n256 & n756 ;
  assign n1119 = ~n255 & n1118 ;
  assign n1122 = n1121 ^ n1119 ;
  assign n1125 = n1124 ^ n1122 ;
  assign n1128 = n1127 ^ n1125 ;
  assign n1131 = n1130 ^ n1128 ;
  assign n1134 = n1133 ^ n1131 ;
  assign n1149 = n750 & n798 ;
  assign n1150 = ~n749 & n1149 ;
  assign n1146 = n727 & n794 ;
  assign n1147 = ~n726 & n1146 ;
  assign n1143 = n666 & n790 ;
  assign n1144 = ~n665 & n1143 ;
  assign n1140 = n567 & n786 ;
  assign n1141 = ~n566 & n1140 ;
  assign n1137 = n430 & n782 ;
  assign n1138 = ~n429 & n1137 ;
  assign n1135 = n256 & n779 ;
  assign n1136 = ~n255 & n1135 ;
  assign n1139 = n1138 ^ n1136 ;
  assign n1142 = n1141 ^ n1139 ;
  assign n1145 = n1144 ^ n1142 ;
  assign n1148 = n1147 ^ n1145 ;
  assign n1151 = n1150 ^ n1148 ;
  assign n1166 = n750 & n821 ;
  assign n1167 = ~n749 & n1166 ;
  assign n1163 = n727 & n817 ;
  assign n1164 = ~n726 & n1163 ;
  assign n1160 = n666 & n813 ;
  assign n1161 = ~n665 & n1160 ;
  assign n1157 = n567 & n809 ;
  assign n1158 = ~n566 & n1157 ;
  assign n1154 = n430 & n805 ;
  assign n1155 = ~n429 & n1154 ;
  assign n1152 = n256 & n802 ;
  assign n1153 = ~n255 & n1152 ;
  assign n1156 = n1155 ^ n1153 ;
  assign n1159 = n1158 ^ n1156 ;
  assign n1162 = n1161 ^ n1159 ;
  assign n1165 = n1164 ^ n1162 ;
  assign n1168 = n1167 ^ n1165 ;
  assign n1183 = n750 & n844 ;
  assign n1184 = ~n749 & n1183 ;
  assign n1180 = n727 & n840 ;
  assign n1181 = ~n726 & n1180 ;
  assign n1177 = n666 & n836 ;
  assign n1178 = ~n665 & n1177 ;
  assign n1174 = n567 & n832 ;
  assign n1175 = ~n566 & n1174 ;
  assign n1171 = n430 & n828 ;
  assign n1172 = ~n429 & n1171 ;
  assign n1169 = n256 & n825 ;
  assign n1170 = ~n255 & n1169 ;
  assign n1173 = n1172 ^ n1170 ;
  assign n1176 = n1175 ^ n1173 ;
  assign n1179 = n1178 ^ n1176 ;
  assign n1182 = n1181 ^ n1179 ;
  assign n1185 = n1184 ^ n1182 ;
  assign n1200 = n750 & n867 ;
  assign n1201 = ~n749 & n1200 ;
  assign n1197 = n727 & n863 ;
  assign n1198 = ~n726 & n1197 ;
  assign n1194 = n666 & n859 ;
  assign n1195 = ~n665 & n1194 ;
  assign n1191 = n567 & n855 ;
  assign n1192 = ~n566 & n1191 ;
  assign n1188 = n430 & n851 ;
  assign n1189 = ~n429 & n1188 ;
  assign n1186 = n256 & n848 ;
  assign n1187 = ~n255 & n1186 ;
  assign n1190 = n1189 ^ n1187 ;
  assign n1193 = n1192 ^ n1190 ;
  assign n1196 = n1195 ^ n1193 ;
  assign n1199 = n1198 ^ n1196 ;
  assign n1202 = n1201 ^ n1199 ;
  assign n1217 = n750 & n890 ;
  assign n1218 = ~n749 & n1217 ;
  assign n1214 = n727 & n886 ;
  assign n1215 = ~n726 & n1214 ;
  assign n1211 = n666 & n882 ;
  assign n1212 = ~n665 & n1211 ;
  assign n1208 = n567 & n878 ;
  assign n1209 = ~n566 & n1208 ;
  assign n1205 = n430 & n874 ;
  assign n1206 = ~n429 & n1205 ;
  assign n1203 = n256 & n871 ;
  assign n1204 = ~n255 & n1203 ;
  assign n1207 = n1206 ^ n1204 ;
  assign n1210 = n1209 ^ n1207 ;
  assign n1213 = n1212 ^ n1210 ;
  assign n1216 = n1215 ^ n1213 ;
  assign n1219 = n1218 ^ n1216 ;
  assign n1234 = n750 & n913 ;
  assign n1235 = ~n749 & n1234 ;
  assign n1231 = n727 & n909 ;
  assign n1232 = ~n726 & n1231 ;
  assign n1228 = n666 & n905 ;
  assign n1229 = ~n665 & n1228 ;
  assign n1225 = n567 & n901 ;
  assign n1226 = ~n566 & n1225 ;
  assign n1222 = n430 & n897 ;
  assign n1223 = ~n429 & n1222 ;
  assign n1220 = n256 & n894 ;
  assign n1221 = ~n255 & n1220 ;
  assign n1224 = n1223 ^ n1221 ;
  assign n1227 = n1226 ^ n1224 ;
  assign n1230 = n1229 ^ n1227 ;
  assign n1233 = n1232 ^ n1230 ;
  assign n1236 = n1235 ^ n1233 ;
  assign n1251 = n750 & n936 ;
  assign n1252 = ~n749 & n1251 ;
  assign n1248 = n727 & n932 ;
  assign n1249 = ~n726 & n1248 ;
  assign n1245 = n666 & n928 ;
  assign n1246 = ~n665 & n1245 ;
  assign n1242 = n567 & n924 ;
  assign n1243 = ~n566 & n1242 ;
  assign n1239 = n430 & n920 ;
  assign n1240 = ~n429 & n1239 ;
  assign n1237 = n256 & n917 ;
  assign n1238 = ~n255 & n1237 ;
  assign n1241 = n1240 ^ n1238 ;
  assign n1244 = n1243 ^ n1241 ;
  assign n1247 = n1246 ^ n1244 ;
  assign n1250 = n1249 ^ n1247 ;
  assign n1253 = n1252 ^ n1250 ;
  assign n1268 = n750 & n959 ;
  assign n1269 = ~n749 & n1268 ;
  assign n1265 = n727 & n955 ;
  assign n1266 = ~n726 & n1265 ;
  assign n1262 = n666 & n951 ;
  assign n1263 = ~n665 & n1262 ;
  assign n1259 = n567 & n947 ;
  assign n1260 = ~n566 & n1259 ;
  assign n1256 = n430 & n943 ;
  assign n1257 = ~n429 & n1256 ;
  assign n1254 = n256 & n940 ;
  assign n1255 = ~n255 & n1254 ;
  assign n1258 = n1257 ^ n1255 ;
  assign n1261 = n1260 ^ n1258 ;
  assign n1264 = n1263 ^ n1261 ;
  assign n1267 = n1266 ^ n1264 ;
  assign n1270 = n1269 ^ n1267 ;
  assign n1285 = n750 & n982 ;
  assign n1286 = ~n749 & n1285 ;
  assign n1282 = n727 & n978 ;
  assign n1283 = ~n726 & n1282 ;
  assign n1279 = n666 & n974 ;
  assign n1280 = ~n665 & n1279 ;
  assign n1276 = n567 & n970 ;
  assign n1277 = ~n566 & n1276 ;
  assign n1273 = n430 & n966 ;
  assign n1274 = ~n429 & n1273 ;
  assign n1271 = n256 & n963 ;
  assign n1272 = ~n255 & n1271 ;
  assign n1275 = n1274 ^ n1272 ;
  assign n1278 = n1277 ^ n1275 ;
  assign n1281 = n1280 ^ n1278 ;
  assign n1284 = n1283 ^ n1281 ;
  assign n1287 = n1286 ^ n1284 ;
  assign n1302 = n750 & n1005 ;
  assign n1303 = ~n749 & n1302 ;
  assign n1299 = n727 & n1001 ;
  assign n1300 = ~n726 & n1299 ;
  assign n1296 = n666 & n997 ;
  assign n1297 = ~n665 & n1296 ;
  assign n1293 = n567 & n993 ;
  assign n1294 = ~n566 & n1293 ;
  assign n1290 = n430 & n989 ;
  assign n1291 = ~n429 & n1290 ;
  assign n1288 = n256 & n986 ;
  assign n1289 = ~n255 & n1288 ;
  assign n1292 = n1291 ^ n1289 ;
  assign n1295 = n1294 ^ n1292 ;
  assign n1298 = n1297 ^ n1295 ;
  assign n1301 = n1300 ^ n1298 ;
  assign n1304 = n1303 ^ n1301 ;
  assign n1319 = n750 & n1028 ;
  assign n1320 = ~n749 & n1319 ;
  assign n1316 = n727 & n1024 ;
  assign n1317 = ~n726 & n1316 ;
  assign n1313 = n666 & n1020 ;
  assign n1314 = ~n665 & n1313 ;
  assign n1310 = n567 & n1016 ;
  assign n1311 = ~n566 & n1310 ;
  assign n1307 = n430 & n1012 ;
  assign n1308 = ~n429 & n1307 ;
  assign n1305 = n256 & n1009 ;
  assign n1306 = ~n255 & n1305 ;
  assign n1309 = n1308 ^ n1306 ;
  assign n1312 = n1311 ^ n1309 ;
  assign n1315 = n1314 ^ n1312 ;
  assign n1318 = n1317 ^ n1315 ;
  assign n1321 = n1320 ^ n1318 ;
  assign n1336 = n750 & n1051 ;
  assign n1337 = ~n749 & n1336 ;
  assign n1333 = n727 & n1047 ;
  assign n1334 = ~n726 & n1333 ;
  assign n1330 = n666 & n1043 ;
  assign n1331 = ~n665 & n1330 ;
  assign n1327 = n567 & n1039 ;
  assign n1328 = ~n566 & n1327 ;
  assign n1324 = n430 & n1035 ;
  assign n1325 = ~n429 & n1324 ;
  assign n1322 = n256 & n1032 ;
  assign n1323 = ~n255 & n1322 ;
  assign n1326 = n1325 ^ n1323 ;
  assign n1329 = n1328 ^ n1326 ;
  assign n1332 = n1331 ^ n1329 ;
  assign n1335 = n1334 ^ n1332 ;
  assign n1338 = n1337 ^ n1335 ;
  assign n1353 = n750 & n1074 ;
  assign n1354 = ~n749 & n1353 ;
  assign n1350 = n727 & n1070 ;
  assign n1351 = ~n726 & n1350 ;
  assign n1347 = n666 & n1066 ;
  assign n1348 = ~n665 & n1347 ;
  assign n1344 = n567 & n1062 ;
  assign n1345 = ~n566 & n1344 ;
  assign n1341 = n430 & n1058 ;
  assign n1342 = ~n429 & n1341 ;
  assign n1339 = n256 & n1055 ;
  assign n1340 = ~n255 & n1339 ;
  assign n1343 = n1342 ^ n1340 ;
  assign n1346 = n1345 ^ n1343 ;
  assign n1349 = n1348 ^ n1346 ;
  assign n1352 = n1351 ^ n1349 ;
  assign n1355 = n1354 ^ n1352 ;
  assign n1370 = n750 & n1097 ;
  assign n1371 = ~n749 & n1370 ;
  assign n1367 = n727 & n1093 ;
  assign n1368 = ~n726 & n1367 ;
  assign n1364 = n666 & n1089 ;
  assign n1365 = ~n665 & n1364 ;
  assign n1361 = n567 & n1085 ;
  assign n1362 = ~n566 & n1361 ;
  assign n1358 = n430 & n1081 ;
  assign n1359 = ~n429 & n1358 ;
  assign n1356 = n256 & n1078 ;
  assign n1357 = ~n255 & n1356 ;
  assign n1360 = n1359 ^ n1357 ;
  assign n1363 = n1362 ^ n1360 ;
  assign n1366 = n1365 ^ n1363 ;
  assign n1369 = n1368 ^ n1366 ;
  assign n1372 = n1371 ^ n1369 ;
  assign n1382 = n749 & n753 ;
  assign n1380 = n726 & n730 ;
  assign n1378 = n665 & n669 ;
  assign n1376 = n566 & n570 ;
  assign n1374 = n429 & n433 ;
  assign n1373 = n255 & n259 ;
  assign n1375 = n1374 ^ n1373 ;
  assign n1377 = n1376 ^ n1375 ;
  assign n1379 = n1378 ^ n1377 ;
  assign n1381 = n1380 ^ n1379 ;
  assign n1383 = n1382 ^ n1381 ;
  assign n1393 = n749 & n776 ;
  assign n1391 = n726 & n772 ;
  assign n1389 = n665 & n768 ;
  assign n1387 = n566 & n764 ;
  assign n1385 = n429 & n760 ;
  assign n1384 = n255 & n757 ;
  assign n1386 = n1385 ^ n1384 ;
  assign n1388 = n1387 ^ n1386 ;
  assign n1390 = n1389 ^ n1388 ;
  assign n1392 = n1391 ^ n1390 ;
  assign n1394 = n1393 ^ n1392 ;
  assign n1404 = n749 & n799 ;
  assign n1402 = n726 & n795 ;
  assign n1400 = n665 & n791 ;
  assign n1398 = n566 & n787 ;
  assign n1396 = n429 & n783 ;
  assign n1395 = n255 & n780 ;
  assign n1397 = n1396 ^ n1395 ;
  assign n1399 = n1398 ^ n1397 ;
  assign n1401 = n1400 ^ n1399 ;
  assign n1403 = n1402 ^ n1401 ;
  assign n1405 = n1404 ^ n1403 ;
  assign n1415 = n749 & n822 ;
  assign n1413 = n726 & n818 ;
  assign n1411 = n665 & n814 ;
  assign n1409 = n566 & n810 ;
  assign n1407 = n429 & n806 ;
  assign n1406 = n255 & n803 ;
  assign n1408 = n1407 ^ n1406 ;
  assign n1410 = n1409 ^ n1408 ;
  assign n1412 = n1411 ^ n1410 ;
  assign n1414 = n1413 ^ n1412 ;
  assign n1416 = n1415 ^ n1414 ;
  assign n1426 = n749 & n845 ;
  assign n1424 = n726 & n841 ;
  assign n1422 = n665 & n837 ;
  assign n1420 = n566 & n833 ;
  assign n1418 = n429 & n829 ;
  assign n1417 = n255 & n826 ;
  assign n1419 = n1418 ^ n1417 ;
  assign n1421 = n1420 ^ n1419 ;
  assign n1423 = n1422 ^ n1421 ;
  assign n1425 = n1424 ^ n1423 ;
  assign n1427 = n1426 ^ n1425 ;
  assign n1437 = n749 & n868 ;
  assign n1435 = n726 & n864 ;
  assign n1433 = n665 & n860 ;
  assign n1431 = n566 & n856 ;
  assign n1429 = n429 & n852 ;
  assign n1428 = n255 & n849 ;
  assign n1430 = n1429 ^ n1428 ;
  assign n1432 = n1431 ^ n1430 ;
  assign n1434 = n1433 ^ n1432 ;
  assign n1436 = n1435 ^ n1434 ;
  assign n1438 = n1437 ^ n1436 ;
  assign n1448 = n749 & n891 ;
  assign n1446 = n726 & n887 ;
  assign n1444 = n665 & n883 ;
  assign n1442 = n566 & n879 ;
  assign n1440 = n429 & n875 ;
  assign n1439 = n255 & n872 ;
  assign n1441 = n1440 ^ n1439 ;
  assign n1443 = n1442 ^ n1441 ;
  assign n1445 = n1444 ^ n1443 ;
  assign n1447 = n1446 ^ n1445 ;
  assign n1449 = n1448 ^ n1447 ;
  assign n1459 = n749 & n914 ;
  assign n1457 = n726 & n910 ;
  assign n1455 = n665 & n906 ;
  assign n1453 = n566 & n902 ;
  assign n1451 = n429 & n898 ;
  assign n1450 = n255 & n895 ;
  assign n1452 = n1451 ^ n1450 ;
  assign n1454 = n1453 ^ n1452 ;
  assign n1456 = n1455 ^ n1454 ;
  assign n1458 = n1457 ^ n1456 ;
  assign n1460 = n1459 ^ n1458 ;
  assign n1470 = n749 & n937 ;
  assign n1468 = n726 & n933 ;
  assign n1466 = n665 & n929 ;
  assign n1464 = n566 & n925 ;
  assign n1462 = n429 & n921 ;
  assign n1461 = n255 & n918 ;
  assign n1463 = n1462 ^ n1461 ;
  assign n1465 = n1464 ^ n1463 ;
  assign n1467 = n1466 ^ n1465 ;
  assign n1469 = n1468 ^ n1467 ;
  assign n1471 = n1470 ^ n1469 ;
  assign n1481 = n749 & n960 ;
  assign n1479 = n726 & n956 ;
  assign n1477 = n665 & n952 ;
  assign n1475 = n566 & n948 ;
  assign n1473 = n429 & n944 ;
  assign n1472 = n255 & n941 ;
  assign n1474 = n1473 ^ n1472 ;
  assign n1476 = n1475 ^ n1474 ;
  assign n1478 = n1477 ^ n1476 ;
  assign n1480 = n1479 ^ n1478 ;
  assign n1482 = n1481 ^ n1480 ;
  assign n1492 = n749 & n983 ;
  assign n1490 = n726 & n979 ;
  assign n1488 = n665 & n975 ;
  assign n1486 = n566 & n971 ;
  assign n1484 = n429 & n967 ;
  assign n1483 = n255 & n964 ;
  assign n1485 = n1484 ^ n1483 ;
  assign n1487 = n1486 ^ n1485 ;
  assign n1489 = n1488 ^ n1487 ;
  assign n1491 = n1490 ^ n1489 ;
  assign n1493 = n1492 ^ n1491 ;
  assign n1503 = n749 & n1006 ;
  assign n1501 = n726 & n1002 ;
  assign n1499 = n665 & n998 ;
  assign n1497 = n566 & n994 ;
  assign n1495 = n429 & n990 ;
  assign n1494 = n255 & n987 ;
  assign n1496 = n1495 ^ n1494 ;
  assign n1498 = n1497 ^ n1496 ;
  assign n1500 = n1499 ^ n1498 ;
  assign n1502 = n1501 ^ n1500 ;
  assign n1504 = n1503 ^ n1502 ;
  assign n1514 = n749 & n1029 ;
  assign n1512 = n726 & n1025 ;
  assign n1510 = n665 & n1021 ;
  assign n1508 = n566 & n1017 ;
  assign n1506 = n429 & n1013 ;
  assign n1505 = n255 & n1010 ;
  assign n1507 = n1506 ^ n1505 ;
  assign n1509 = n1508 ^ n1507 ;
  assign n1511 = n1510 ^ n1509 ;
  assign n1513 = n1512 ^ n1511 ;
  assign n1515 = n1514 ^ n1513 ;
  assign n1525 = n749 & n1052 ;
  assign n1523 = n726 & n1048 ;
  assign n1521 = n665 & n1044 ;
  assign n1519 = n566 & n1040 ;
  assign n1517 = n429 & n1036 ;
  assign n1516 = n255 & n1033 ;
  assign n1518 = n1517 ^ n1516 ;
  assign n1520 = n1519 ^ n1518 ;
  assign n1522 = n1521 ^ n1520 ;
  assign n1524 = n1523 ^ n1522 ;
  assign n1526 = n1525 ^ n1524 ;
  assign n1536 = n749 & n1075 ;
  assign n1534 = n726 & n1071 ;
  assign n1532 = n665 & n1067 ;
  assign n1530 = n566 & n1063 ;
  assign n1528 = n429 & n1059 ;
  assign n1527 = n255 & n1056 ;
  assign n1529 = n1528 ^ n1527 ;
  assign n1531 = n1530 ^ n1529 ;
  assign n1533 = n1532 ^ n1531 ;
  assign n1535 = n1534 ^ n1533 ;
  assign n1537 = n1536 ^ n1535 ;
  assign n1547 = n749 & n1098 ;
  assign n1545 = n726 & n1094 ;
  assign n1543 = n665 & n1090 ;
  assign n1541 = n566 & n1086 ;
  assign n1539 = n429 & n1082 ;
  assign n1538 = n255 & n1079 ;
  assign n1540 = n1539 ^ n1538 ;
  assign n1542 = n1541 ^ n1540 ;
  assign n1544 = n1543 ^ n1542 ;
  assign n1546 = n1545 ^ n1544 ;
  assign n1548 = n1547 ^ n1546 ;
  assign y0 = n755 ;
  assign y1 = n778 ;
  assign y2 = n801 ;
  assign y3 = n824 ;
  assign y4 = n847 ;
  assign y5 = n870 ;
  assign y6 = n893 ;
  assign y7 = n916 ;
  assign y8 = n939 ;
  assign y9 = n962 ;
  assign y10 = n985 ;
  assign y11 = n1008 ;
  assign y12 = n1031 ;
  assign y13 = n1054 ;
  assign y14 = n1077 ;
  assign y15 = n1100 ;
  assign y16 = n1117 ;
  assign y17 = n1134 ;
  assign y18 = n1151 ;
  assign y19 = n1168 ;
  assign y20 = n1185 ;
  assign y21 = n1202 ;
  assign y22 = n1219 ;
  assign y23 = n1236 ;
  assign y24 = n1253 ;
  assign y25 = n1270 ;
  assign y26 = n1287 ;
  assign y27 = n1304 ;
  assign y28 = n1321 ;
  assign y29 = n1338 ;
  assign y30 = n1355 ;
  assign y31 = n1372 ;
  assign y32 = n1383 ;
  assign y33 = n1394 ;
  assign y34 = n1405 ;
  assign y35 = n1416 ;
  assign y36 = n1427 ;
  assign y37 = n1438 ;
  assign y38 = n1449 ;
  assign y39 = n1460 ;
  assign y40 = n1471 ;
  assign y41 = n1482 ;
  assign y42 = n1493 ;
  assign y43 = n1504 ;
  assign y44 = n1515 ;
  assign y45 = n1526 ;
  assign y46 = n1537 ;
  assign y47 = n1548 ;
endmodule
