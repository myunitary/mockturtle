module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , y0 , y1 , y2 , y3 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 ;
  output y0 , y1 , y2 , y3 ;
  wire n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 ;
  assign n115 = x63 ^ x7 ;
  assign n342 = x105 ^ x49 ;
  assign n343 = x104 ^ x48 ;
  assign n344 = ~n342 & ~n343 ;
  assign n345 = x107 ^ x51 ;
  assign n346 = x106 ^ x50 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = n344 & n347 ;
  assign n370 = x111 ^ x55 ;
  assign n371 = x110 ^ x54 ;
  assign n372 = n370 & n371 ;
  assign n349 = x109 ^ x53 ;
  assign n350 = x108 ^ x52 ;
  assign n373 = ~n349 & ~n350 ;
  assign n374 = n372 & n373 ;
  assign n351 = n349 & ~n350 ;
  assign n352 = n351 ^ n350 ;
  assign n375 = n374 ^ n352 ;
  assign n376 = n348 & n375 ;
  assign n356 = n345 & ~n346 ;
  assign n357 = n356 ^ n346 ;
  assign n358 = n344 & n357 ;
  assign n354 = n342 & ~n343 ;
  assign n355 = n354 ^ n343 ;
  assign n359 = n358 ^ n355 ;
  assign n377 = n376 ^ n359 ;
  assign n378 = ~n115 & n377 ;
  assign n120 = x67 ^ x11 ;
  assign n121 = x66 ^ x10 ;
  assign n122 = n120 & n121 ;
  assign n123 = x65 ^ x9 ;
  assign n124 = x64 ^ x8 ;
  assign n125 = n123 & n124 ;
  assign n126 = n125 ^ n123 ;
  assign n127 = n126 ^ n124 ;
  assign n128 = n122 & ~n127 ;
  assign n129 = x69 ^ x13 ;
  assign n130 = x68 ^ x12 ;
  assign n131 = n129 & n130 ;
  assign n140 = n131 ^ n129 ;
  assign n141 = n140 ^ n130 ;
  assign n116 = x70 ^ x14 ;
  assign n117 = x71 ^ x15 ;
  assign n142 = n116 & n117 ;
  assign n143 = ~n141 & n142 ;
  assign n138 = n129 & ~n130 ;
  assign n139 = n138 ^ n130 ;
  assign n144 = n143 ^ n139 ;
  assign n145 = n128 & n144 ;
  assign n134 = n123 & ~n124 ;
  assign n135 = n134 ^ n124 ;
  assign n146 = n145 ^ n135 ;
  assign n147 = n135 ^ n115 ;
  assign n148 = ~n115 & n147 ;
  assign n149 = n148 ^ n115 ;
  assign n150 = n149 ^ n145 ;
  assign n151 = n146 & n150 ;
  assign n152 = n151 ^ n148 ;
  assign n153 = n152 ^ n145 ;
  assign n118 = ~n116 & n117 ;
  assign n119 = n118 ^ n116 ;
  assign n132 = n128 & n131 ;
  assign n133 = n119 & n132 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = ~n115 & n136 ;
  assign n154 = n153 ^ n137 ;
  assign n114 = x62 ^ x6 ;
  assign n155 = n154 ^ n114 ;
  assign n113 = x61 ^ x5 ;
  assign n164 = n155 ^ n113 ;
  assign n163 = x60 ^ x4 ;
  assign n172 = n164 ^ n163 ;
  assign n171 = x59 ^ x3 ;
  assign n207 = n172 ^ n171 ;
  assign n179 = x73 ^ x17 ;
  assign n180 = x72 ^ x16 ;
  assign n183 = ~n179 & ~n180 ;
  assign n184 = x75 ^ x19 ;
  assign n185 = x74 ^ x18 ;
  assign n189 = ~n184 & n185 ;
  assign n190 = n183 & n189 ;
  assign n191 = x77 ^ x21 ;
  assign n192 = x76 ^ x20 ;
  assign n194 = ~n191 & n192 ;
  assign n195 = x79 ^ x23 ;
  assign n196 = x78 ^ x22 ;
  assign n203 = ~n195 & ~n196 ;
  assign n204 = n194 & n203 ;
  assign n205 = n190 & n204 ;
  assign n197 = n195 & ~n196 ;
  assign n198 = n197 ^ n196 ;
  assign n199 = n194 & n198 ;
  assign n193 = n191 & n192 ;
  assign n200 = n199 ^ n193 ;
  assign n201 = n190 & n200 ;
  assign n186 = n184 & n185 ;
  assign n187 = n183 & n186 ;
  assign n181 = n179 & ~n180 ;
  assign n182 = n181 ^ n180 ;
  assign n188 = n187 ^ n182 ;
  assign n202 = n201 ^ n188 ;
  assign n206 = n205 ^ n202 ;
  assign n300 = n207 ^ n206 ;
  assign n226 = x91 ^ x35 ;
  assign n217 = x92 ^ x36 ;
  assign n227 = n226 ^ n217 ;
  assign n228 = ~n226 & ~n227 ;
  assign n229 = n228 ^ n226 ;
  assign n218 = x94 ^ x38 ;
  assign n219 = x93 ^ x37 ;
  assign n220 = n218 & n219 ;
  assign n221 = n220 ^ n219 ;
  assign n222 = n221 ^ n218 ;
  assign n230 = n229 ^ n222 ;
  assign n231 = n222 ^ n217 ;
  assign n232 = ~n230 & n231 ;
  assign n233 = n232 ^ n228 ;
  assign n234 = n233 ^ n222 ;
  assign n223 = n217 & n222 ;
  assign n224 = n223 ^ n222 ;
  assign n225 = n224 ^ n222 ;
  assign n235 = n234 ^ n225 ;
  assign n236 = x90 ^ x34 ;
  assign n240 = x89 ^ x33 ;
  assign n241 = ~n236 & n240 ;
  assign n242 = n235 & n241 ;
  assign n237 = ~n235 & n236 ;
  assign n238 = n237 ^ n236 ;
  assign n239 = n238 ^ n235 ;
  assign n243 = n242 ^ n239 ;
  assign n216 = x88 ^ x32 ;
  assign n244 = n243 ^ n216 ;
  assign n215 = x80 ^ x24 ;
  assign n246 = n244 ^ n215 ;
  assign n247 = x81 ^ x25 ;
  assign n252 = n247 ^ n240 ;
  assign n253 = n252 ^ n239 ;
  assign n254 = ~n246 & ~n253 ;
  assign n274 = x86 ^ x30 ;
  assign n276 = n274 ^ n218 ;
  assign n277 = x87 ^ x31 ;
  assign n278 = x95 ^ x39 ;
  assign n279 = n277 & n278 ;
  assign n280 = n279 ^ n278 ;
  assign n281 = n276 & n280 ;
  assign n275 = ~n218 & ~n274 ;
  assign n282 = n281 ^ n275 ;
  assign n266 = x84 ^ x28 ;
  assign n268 = n266 ^ n231 ;
  assign n283 = n282 ^ n268 ;
  assign n270 = x85 ^ x29 ;
  assign n269 = n219 ^ n218 ;
  assign n284 = n270 ^ n269 ;
  assign n285 = n284 ^ n268 ;
  assign n286 = n284 & n285 ;
  assign n287 = n286 ^ n284 ;
  assign n288 = n287 ^ n285 ;
  assign n289 = n288 ^ n268 ;
  assign n290 = n283 & ~n289 ;
  assign n291 = n290 ^ n289 ;
  assign n292 = n291 ^ n288 ;
  assign n293 = n292 ^ n282 ;
  assign n271 = ~n269 & ~n270 ;
  assign n272 = ~n268 & n271 ;
  assign n267 = n231 & ~n266 ;
  assign n273 = n272 ^ n267 ;
  assign n294 = n293 ^ n273 ;
  assign n256 = n236 ^ n235 ;
  assign n255 = x82 ^ x26 ;
  assign n258 = n256 ^ n255 ;
  assign n260 = x83 ^ x27 ;
  assign n259 = n226 ^ n225 ;
  assign n295 = n260 ^ n259 ;
  assign n296 = ~n258 & n295 ;
  assign n297 = n294 & n296 ;
  assign n298 = n254 & n297 ;
  assign n261 = ~n259 & ~n260 ;
  assign n262 = ~n258 & n261 ;
  assign n257 = ~n255 & n256 ;
  assign n263 = n262 ^ n257 ;
  assign n264 = n254 & n263 ;
  assign n248 = n240 ^ n239 ;
  assign n249 = ~n247 & n248 ;
  assign n250 = ~n246 & n249 ;
  assign n245 = ~n215 & n244 ;
  assign n251 = n250 ^ n245 ;
  assign n265 = n264 ^ n251 ;
  assign n299 = n298 ^ n265 ;
  assign n332 = n300 ^ n299 ;
  assign n308 = x97 ^ x41 ;
  assign n309 = x96 ^ x40 ;
  assign n312 = ~n308 & ~n309 ;
  assign n313 = x98 ^ x42 ;
  assign n316 = x99 ^ x43 ;
  assign n317 = ~n313 & n316 ;
  assign n318 = n312 & n317 ;
  assign n319 = x101 ^ x45 ;
  assign n320 = x100 ^ x44 ;
  assign n321 = n319 & n320 ;
  assign n322 = x103 ^ x47 ;
  assign n323 = x102 ^ x46 ;
  assign n328 = ~n322 & n323 ;
  assign n329 = n321 & n328 ;
  assign n330 = n318 & n329 ;
  assign n324 = n322 & n323 ;
  assign n325 = n321 & n324 ;
  assign n326 = n318 & n325 ;
  assign n314 = n312 & n313 ;
  assign n310 = n308 & ~n309 ;
  assign n311 = n310 ^ n309 ;
  assign n315 = n314 ^ n311 ;
  assign n327 = n326 ^ n315 ;
  assign n331 = n330 ^ n327 ;
  assign n362 = n332 ^ n331 ;
  assign n353 = n348 & n352 ;
  assign n360 = n359 ^ n353 ;
  assign n361 = n115 & n360 ;
  assign n379 = n362 ^ n361 ;
  assign n380 = n378 & n379 ;
  assign n158 = n114 & n154 ;
  assign n157 = n137 & n153 ;
  assign n159 = n158 ^ n157 ;
  assign n156 = n113 & n155 ;
  assign n166 = n159 ^ n156 ;
  assign n165 = n163 & n164 ;
  assign n174 = n166 ^ n165 ;
  assign n173 = n171 & n172 ;
  assign n210 = n174 ^ n173 ;
  assign n208 = n206 & n207 ;
  assign n209 = n208 ^ n207 ;
  assign n303 = n210 ^ n209 ;
  assign n301 = n299 & n300 ;
  assign n302 = n301 ^ n299 ;
  assign n336 = n303 ^ n302 ;
  assign n333 = n331 & n332 ;
  assign n334 = n333 ^ n331 ;
  assign n335 = n334 ^ n332 ;
  assign n364 = n336 ^ n335 ;
  assign n363 = n361 & n362 ;
  assign n381 = n364 ^ n363 ;
  assign n382 = n380 & n381 ;
  assign n383 = n382 ^ n380 ;
  assign n161 = n157 & n158 ;
  assign n160 = n156 & n159 ;
  assign n168 = n161 ^ n160 ;
  assign n167 = n165 & n166 ;
  assign n176 = n168 ^ n167 ;
  assign n175 = n173 & n174 ;
  assign n212 = n176 ^ n175 ;
  assign n211 = n209 & n210 ;
  assign n305 = n212 ^ n211 ;
  assign n304 = n302 & n303 ;
  assign n339 = n305 ^ n304 ;
  assign n337 = n335 & n336 ;
  assign n338 = n337 ^ n336 ;
  assign n367 = n339 ^ n338 ;
  assign n365 = n363 & n364 ;
  assign n366 = n365 ^ n363 ;
  assign n384 = n367 ^ n366 ;
  assign n385 = n383 & n384 ;
  assign n368 = n366 & n367 ;
  assign n340 = n338 & n339 ;
  assign n306 = n304 & n305 ;
  assign n213 = n211 & n212 ;
  assign n177 = n175 & n176 ;
  assign n169 = n167 & n168 ;
  assign n162 = n160 & n161 ;
  assign n170 = n169 ^ n162 ;
  assign n178 = n177 ^ n170 ;
  assign n214 = n213 ^ n178 ;
  assign n307 = n306 ^ n214 ;
  assign n341 = n340 ^ n307 ;
  assign n369 = n368 ^ n341 ;
  assign n386 = n385 ^ n369 ;
  assign n387 = n384 ^ n383 ;
  assign n388 = n381 ^ n380 ;
  assign n389 = n379 ^ n378 ;
  assign y0 = n386 ;
  assign y1 = n387 ;
  assign y2 = ~n388 ;
  assign y3 = n389 ;
endmodule
