// nine parties (one provide the reference data), each holding a 32-bit data, finding the three closest to the reference
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 ;
  wire n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 ;
  assign n387 = x258 ^ x162 ;
  assign n384 = x266 ^ x170 ;
  assign n382 = x272 ^ x176 ;
  assign n380 = x270 ^ x174 ;
  assign n379 = x271 ^ x175 ;
  assign n381 = n380 ^ n379 ;
  assign n383 = n382 ^ n381 ;
  assign n385 = n384 ^ n383 ;
  assign n377 = x269 ^ x173 ;
  assign n375 = x267 ^ x171 ;
  assign n374 = x268 ^ x172 ;
  assign n376 = n375 ^ n374 ;
  assign n378 = n377 ^ n376 ;
  assign n386 = n385 ^ n378 ;
  assign n388 = n387 ^ n386 ;
  assign n371 = x259 ^ x163 ;
  assign n369 = x265 ^ x169 ;
  assign n367 = x263 ^ x167 ;
  assign n366 = x264 ^ x168 ;
  assign n368 = n367 ^ n366 ;
  assign n370 = n369 ^ n368 ;
  assign n372 = n371 ^ n370 ;
  assign n364 = x262 ^ x166 ;
  assign n362 = x260 ^ x164 ;
  assign n361 = x261 ^ x165 ;
  assign n363 = n362 ^ n361 ;
  assign n365 = n364 ^ n363 ;
  assign n373 = n372 ^ n365 ;
  assign n416 = n387 ^ n373 ;
  assign n417 = n388 & ~n416 ;
  assign n418 = n417 ^ n386 ;
  assign n412 = n377 ^ n375 ;
  assign n413 = n376 & ~n412 ;
  assign n414 = n413 ^ n374 ;
  assign n408 = n382 ^ n380 ;
  assign n409 = n381 & ~n408 ;
  assign n410 = n409 ^ n379 ;
  assign n405 = n383 ^ n378 ;
  assign n406 = ~n385 & n405 ;
  assign n407 = n406 ^ n378 ;
  assign n411 = n410 ^ n407 ;
  assign n415 = n414 ^ n411 ;
  assign n419 = n418 ^ n415 ;
  assign n401 = n364 ^ n362 ;
  assign n402 = n363 & ~n401 ;
  assign n403 = n402 ^ n361 ;
  assign n397 = n370 ^ n365 ;
  assign n398 = ~n372 & n397 ;
  assign n399 = n398 ^ n365 ;
  assign n394 = n369 ^ n367 ;
  assign n395 = n368 & ~n394 ;
  assign n396 = n395 ^ n366 ;
  assign n400 = n399 ^ n396 ;
  assign n404 = n403 ^ n400 ;
  assign n431 = n418 ^ n404 ;
  assign n432 = n419 & ~n431 ;
  assign n433 = n432 ^ n415 ;
  assign n428 = n414 ^ n410 ;
  assign n429 = n411 & ~n428 ;
  assign n430 = n429 ^ n407 ;
  assign n434 = n433 ^ n430 ;
  assign n425 = n403 ^ n399 ;
  assign n426 = n400 & ~n425 ;
  assign n427 = n426 ^ n396 ;
  assign n440 = n430 ^ n427 ;
  assign n441 = ~n434 & n440 ;
  assign n442 = n441 ^ n427 ;
  assign n359 = x257 ^ x161 ;
  assign n325 = x277 ^ x181 ;
  assign n323 = x275 ^ x179 ;
  assign n322 = x276 ^ x180 ;
  assign n324 = n323 ^ n322 ;
  assign n326 = n325 ^ n324 ;
  assign n320 = x274 ^ x178 ;
  assign n318 = x280 ^ x184 ;
  assign n316 = x278 ^ x182 ;
  assign n315 = x279 ^ x183 ;
  assign n317 = n316 ^ n315 ;
  assign n319 = n318 ^ n317 ;
  assign n321 = n320 ^ n319 ;
  assign n327 = n326 ^ n321 ;
  assign n298 = x282 ^ x186 ;
  assign n297 = x283 ^ x187 ;
  assign n299 = n298 ^ n297 ;
  assign n296 = x284 ^ x188 ;
  assign n300 = n299 ^ n296 ;
  assign n294 = x281 ^ x185 ;
  assign n291 = x285 ^ x189 ;
  assign n290 = x286 ^ x190 ;
  assign n292 = n291 ^ n290 ;
  assign n289 = x287 ^ x191 ;
  assign n293 = n292 ^ n289 ;
  assign n295 = n294 ^ n293 ;
  assign n313 = n300 ^ n295 ;
  assign n312 = x273 ^ x177 ;
  assign n314 = n313 ^ n312 ;
  assign n358 = n327 ^ n314 ;
  assign n360 = n359 ^ n358 ;
  assign n389 = n388 ^ n373 ;
  assign n390 = n389 ^ n359 ;
  assign n391 = n360 & ~n390 ;
  assign n392 = n391 ^ n358 ;
  assign n339 = n325 ^ n323 ;
  assign n340 = n324 & ~n339 ;
  assign n341 = n340 ^ n322 ;
  assign n335 = n318 ^ n316 ;
  assign n336 = n317 & ~n335 ;
  assign n337 = n336 ^ n315 ;
  assign n332 = n326 ^ n320 ;
  assign n333 = n321 & ~n332 ;
  assign n334 = n333 ^ n319 ;
  assign n338 = n337 ^ n334 ;
  assign n342 = n341 ^ n338 ;
  assign n328 = n327 ^ n313 ;
  assign n329 = n314 & ~n328 ;
  assign n330 = n329 ^ n312 ;
  assign n308 = n297 ^ n296 ;
  assign n309 = ~n299 & n308 ;
  assign n310 = n309 ^ n296 ;
  assign n304 = n290 ^ n289 ;
  assign n305 = ~n292 & n304 ;
  assign n306 = n305 ^ n289 ;
  assign n301 = n300 ^ n294 ;
  assign n302 = n295 & ~n301 ;
  assign n303 = n302 ^ n293 ;
  assign n307 = n306 ^ n303 ;
  assign n311 = n310 ^ n307 ;
  assign n331 = n330 ^ n311 ;
  assign n357 = n342 ^ n331 ;
  assign n393 = n392 ^ n357 ;
  assign n420 = n419 ^ n404 ;
  assign n421 = n420 ^ n357 ;
  assign n422 = n393 & ~n421 ;
  assign n423 = n422 ^ n392 ;
  assign n350 = n341 ^ n337 ;
  assign n351 = n338 & ~n350 ;
  assign n352 = n351 ^ n334 ;
  assign n346 = n310 ^ n306 ;
  assign n347 = n307 & ~n346 ;
  assign n348 = n347 ^ n303 ;
  assign n343 = n342 ^ n330 ;
  assign n344 = n331 & ~n343 ;
  assign n345 = n344 ^ n311 ;
  assign n349 = n348 ^ n345 ;
  assign n356 = n352 ^ n349 ;
  assign n424 = n423 ^ n356 ;
  assign n435 = n434 ^ n427 ;
  assign n436 = n435 ^ n423 ;
  assign n437 = n424 & ~n436 ;
  assign n438 = n437 ^ n356 ;
  assign n353 = n352 ^ n348 ;
  assign n354 = n349 & ~n353 ;
  assign n355 = n354 ^ n345 ;
  assign n439 = n438 ^ n355 ;
  assign n443 = n442 ^ n439 ;
  assign n444 = n420 ^ n393 ;
  assign n445 = n389 ^ n360 ;
  assign n446 = x256 ^ x160 ;
  assign n447 = n445 & n446 ;
  assign n448 = n444 & n447 ;
  assign n449 = n435 ^ n424 ;
  assign n450 = n448 & n449 ;
  assign n451 = n443 & n450 ;
  assign n452 = n442 ^ n438 ;
  assign n453 = n439 & ~n452 ;
  assign n454 = n453 ^ n355 ;
  assign n455 = n451 & n454 ;
  assign n557 = x277 ^ x245 ;
  assign n555 = x275 ^ x243 ;
  assign n554 = x276 ^ x244 ;
  assign n556 = n555 ^ n554 ;
  assign n558 = n557 ^ n556 ;
  assign n550 = x279 ^ x247 ;
  assign n549 = x278 ^ x246 ;
  assign n551 = n550 ^ n549 ;
  assign n548 = x280 ^ x248 ;
  assign n552 = n551 ^ n548 ;
  assign n547 = x274 ^ x242 ;
  assign n553 = n552 ^ n547 ;
  assign n559 = n558 ^ n553 ;
  assign n534 = x284 ^ x252 ;
  assign n532 = x282 ^ x250 ;
  assign n531 = x283 ^ x251 ;
  assign n533 = n532 ^ n531 ;
  assign n535 = n534 ^ n533 ;
  assign n524 = x287 ^ x255 ;
  assign n522 = x286 ^ x254 ;
  assign n521 = x285 ^ x253 ;
  assign n523 = n522 ^ n521 ;
  assign n529 = n524 ^ n523 ;
  assign n528 = x281 ^ x249 ;
  assign n530 = n529 ^ n528 ;
  assign n545 = n535 ^ n530 ;
  assign n544 = x273 ^ x241 ;
  assign n546 = n545 ^ n544 ;
  assign n588 = n559 ^ n546 ;
  assign n587 = x257 ^ x225 ;
  assign n589 = n588 ^ n587 ;
  assign n492 = x262 ^ x230 ;
  assign n490 = x260 ^ x228 ;
  assign n489 = x261 ^ x229 ;
  assign n491 = n490 ^ n489 ;
  assign n493 = n492 ^ n491 ;
  assign n487 = x259 ^ x227 ;
  assign n482 = x265 ^ x233 ;
  assign n480 = x263 ^ x231 ;
  assign n479 = x264 ^ x232 ;
  assign n481 = n480 ^ n479 ;
  assign n486 = n482 ^ n481 ;
  assign n488 = n487 ^ n486 ;
  assign n506 = n493 ^ n488 ;
  assign n466 = x269 ^ x237 ;
  assign n464 = x267 ^ x235 ;
  assign n463 = x268 ^ x236 ;
  assign n465 = n464 ^ n463 ;
  assign n467 = n466 ^ n465 ;
  assign n461 = x266 ^ x234 ;
  assign n459 = x272 ^ x240 ;
  assign n457 = x270 ^ x238 ;
  assign n456 = x271 ^ x239 ;
  assign n458 = n457 ^ n456 ;
  assign n460 = n459 ^ n458 ;
  assign n462 = n461 ^ n460 ;
  assign n504 = n467 ^ n462 ;
  assign n503 = x258 ^ x226 ;
  assign n505 = n504 ^ n503 ;
  assign n590 = n506 ^ n505 ;
  assign n591 = n590 ^ n588 ;
  assign n592 = n589 & ~n591 ;
  assign n593 = n592 ^ n587 ;
  assign n571 = n557 ^ n555 ;
  assign n572 = n556 & ~n571 ;
  assign n573 = n572 ^ n554 ;
  assign n567 = n558 ^ n552 ;
  assign n568 = n553 & ~n567 ;
  assign n569 = n568 ^ n547 ;
  assign n564 = n550 ^ n548 ;
  assign n565 = n551 & ~n564 ;
  assign n566 = n565 ^ n549 ;
  assign n570 = n569 ^ n566 ;
  assign n574 = n573 ^ n570 ;
  assign n560 = n559 ^ n544 ;
  assign n561 = ~n546 & n560 ;
  assign n562 = n561 ^ n559 ;
  assign n540 = n534 ^ n532 ;
  assign n541 = n533 & ~n540 ;
  assign n542 = n541 ^ n531 ;
  assign n536 = n535 ^ n528 ;
  assign n537 = ~n530 & n536 ;
  assign n538 = n537 ^ n535 ;
  assign n525 = n524 ^ n522 ;
  assign n526 = n523 & ~n525 ;
  assign n527 = n526 ^ n521 ;
  assign n539 = n538 ^ n527 ;
  assign n543 = n542 ^ n539 ;
  assign n563 = n562 ^ n543 ;
  assign n586 = n574 ^ n563 ;
  assign n594 = n593 ^ n586 ;
  assign n507 = n506 ^ n504 ;
  assign n508 = n505 & ~n507 ;
  assign n509 = n508 ^ n503 ;
  assign n498 = n492 ^ n490 ;
  assign n499 = n491 & ~n498 ;
  assign n500 = n499 ^ n489 ;
  assign n494 = n493 ^ n486 ;
  assign n495 = ~n488 & n494 ;
  assign n496 = n495 ^ n493 ;
  assign n483 = n482 ^ n480 ;
  assign n484 = n481 & ~n483 ;
  assign n485 = n484 ^ n479 ;
  assign n497 = n496 ^ n485 ;
  assign n501 = n500 ^ n497 ;
  assign n475 = n466 ^ n464 ;
  assign n476 = n465 & ~n475 ;
  assign n477 = n476 ^ n463 ;
  assign n471 = n459 ^ n457 ;
  assign n472 = n458 & ~n471 ;
  assign n473 = n472 ^ n456 ;
  assign n468 = n467 ^ n460 ;
  assign n469 = ~n462 & n468 ;
  assign n470 = n469 ^ n467 ;
  assign n474 = n473 ^ n470 ;
  assign n478 = n477 ^ n474 ;
  assign n502 = n501 ^ n478 ;
  assign n595 = n509 ^ n502 ;
  assign n596 = n595 ^ n586 ;
  assign n597 = n594 & ~n596 ;
  assign n598 = n597 ^ n593 ;
  assign n582 = n573 ^ n569 ;
  assign n583 = n570 & n582 ;
  assign n584 = n583 ^ n569 ;
  assign n578 = n542 ^ n527 ;
  assign n579 = n539 & n578 ;
  assign n580 = n579 ^ n527 ;
  assign n575 = n574 ^ n543 ;
  assign n576 = ~n563 & n575 ;
  assign n577 = n576 ^ n574 ;
  assign n581 = n580 ^ n577 ;
  assign n585 = n584 ^ n581 ;
  assign n599 = n598 ^ n585 ;
  assign n517 = n500 ^ n496 ;
  assign n518 = n497 & n517 ;
  assign n519 = n518 ^ n496 ;
  assign n513 = n477 ^ n473 ;
  assign n514 = n474 & ~n513 ;
  assign n515 = n514 ^ n470 ;
  assign n510 = n509 ^ n478 ;
  assign n511 = ~n502 & n510 ;
  assign n512 = n511 ^ n509 ;
  assign n516 = n515 ^ n512 ;
  assign n520 = n519 ^ n516 ;
  assign n600 = n599 ^ n520 ;
  assign n601 = n595 ^ n594 ;
  assign n602 = x256 ^ x224 ;
  assign n603 = n590 ^ n589 ;
  assign n604 = n602 & n603 ;
  assign n605 = n601 & n604 ;
  assign n606 = n600 & n605 ;
  assign n614 = n519 ^ n515 ;
  assign n615 = n516 & ~n614 ;
  assign n616 = n615 ^ n512 ;
  assign n610 = n584 ^ n580 ;
  assign n611 = n581 & ~n610 ;
  assign n612 = n611 ^ n577 ;
  assign n607 = n585 ^ n520 ;
  assign n608 = ~n599 & n607 ;
  assign n609 = n608 ^ n520 ;
  assign n613 = n612 ^ n609 ;
  assign n617 = n616 ^ n613 ;
  assign n618 = n606 & n617 ;
  assign n619 = n616 ^ n612 ;
  assign n620 = n613 & ~n619 ;
  assign n621 = n620 ^ n609 ;
  assign n622 = n618 & n621 ;
  assign n661 = x280 ^ x216 ;
  assign n659 = x279 ^ x215 ;
  assign n658 = x278 ^ x214 ;
  assign n660 = n659 ^ n658 ;
  assign n662 = n661 ^ n660 ;
  assign n657 = x274 ^ x210 ;
  assign n663 = n662 ^ n657 ;
  assign n655 = x277 ^ x213 ;
  assign n653 = x275 ^ x211 ;
  assign n652 = x276 ^ x212 ;
  assign n654 = n653 ^ n652 ;
  assign n656 = n655 ^ n654 ;
  assign n675 = n662 ^ n656 ;
  assign n676 = n663 & ~n675 ;
  assign n677 = n676 ^ n657 ;
  assign n672 = n661 ^ n659 ;
  assign n673 = n660 & ~n672 ;
  assign n674 = n673 ^ n658 ;
  assign n678 = n677 ^ n674 ;
  assign n669 = n655 ^ n653 ;
  assign n670 = n654 & ~n669 ;
  assign n671 = n670 ^ n652 ;
  assign n684 = n677 ^ n671 ;
  assign n685 = n678 & n684 ;
  assign n686 = n685 ^ n677 ;
  assign n635 = x283 ^ x219 ;
  assign n634 = x282 ^ x218 ;
  assign n636 = n635 ^ n634 ;
  assign n633 = x284 ^ x220 ;
  assign n637 = n636 ^ n633 ;
  assign n626 = x287 ^ x223 ;
  assign n624 = x286 ^ x222 ;
  assign n623 = x285 ^ x221 ;
  assign n625 = n624 ^ n623 ;
  assign n631 = n626 ^ n625 ;
  assign n630 = x281 ^ x217 ;
  assign n632 = n631 ^ n630 ;
  assign n650 = n637 ^ n632 ;
  assign n649 = x273 ^ x209 ;
  assign n651 = n650 ^ n649 ;
  assign n664 = n663 ^ n656 ;
  assign n665 = n664 ^ n649 ;
  assign n666 = ~n651 & n665 ;
  assign n667 = n666 ^ n664 ;
  assign n642 = n635 ^ n633 ;
  assign n643 = n636 & ~n642 ;
  assign n644 = n643 ^ n634 ;
  assign n638 = n637 ^ n630 ;
  assign n639 = ~n632 & n638 ;
  assign n640 = n639 ^ n637 ;
  assign n627 = n626 ^ n624 ;
  assign n628 = n625 & ~n627 ;
  assign n629 = n628 ^ n623 ;
  assign n641 = n640 ^ n629 ;
  assign n648 = n644 ^ n641 ;
  assign n668 = n667 ^ n648 ;
  assign n679 = n678 ^ n671 ;
  assign n680 = n679 ^ n648 ;
  assign n681 = ~n668 & n680 ;
  assign n682 = n681 ^ n679 ;
  assign n645 = n644 ^ n629 ;
  assign n646 = ~n641 & n645 ;
  assign n647 = n646 ^ n644 ;
  assign n683 = n682 ^ n647 ;
  assign n757 = n686 ^ n683 ;
  assign n692 = n664 ^ n651 ;
  assign n691 = x257 ^ x193 ;
  assign n693 = n692 ^ n691 ;
  assign n719 = x262 ^ x198 ;
  assign n717 = x260 ^ x196 ;
  assign n716 = x261 ^ x197 ;
  assign n718 = n717 ^ n716 ;
  assign n720 = n719 ^ n718 ;
  assign n714 = x259 ^ x195 ;
  assign n712 = x265 ^ x201 ;
  assign n710 = x263 ^ x199 ;
  assign n709 = x264 ^ x200 ;
  assign n711 = n710 ^ n709 ;
  assign n713 = n712 ^ n711 ;
  assign n715 = n714 ^ n713 ;
  assign n721 = n720 ^ n715 ;
  assign n705 = x269 ^ x205 ;
  assign n703 = x267 ^ x203 ;
  assign n702 = x268 ^ x204 ;
  assign n704 = n703 ^ n702 ;
  assign n706 = n705 ^ n704 ;
  assign n700 = x266 ^ x202 ;
  assign n698 = x272 ^ x208 ;
  assign n696 = x270 ^ x206 ;
  assign n695 = x271 ^ x207 ;
  assign n697 = n696 ^ n695 ;
  assign n699 = n698 ^ n697 ;
  assign n701 = n700 ^ n699 ;
  assign n707 = n706 ^ n701 ;
  assign n694 = x258 ^ x194 ;
  assign n708 = n707 ^ n694 ;
  assign n722 = n721 ^ n708 ;
  assign n723 = n722 ^ n692 ;
  assign n724 = n693 & ~n723 ;
  assign n725 = n724 ^ n691 ;
  assign n690 = n679 ^ n668 ;
  assign n726 = n725 ^ n690 ;
  assign n750 = n721 ^ n707 ;
  assign n751 = n708 & ~n750 ;
  assign n752 = n751 ^ n694 ;
  assign n745 = n719 ^ n717 ;
  assign n746 = n718 & ~n745 ;
  assign n747 = n746 ^ n716 ;
  assign n741 = n720 ^ n713 ;
  assign n742 = ~n715 & n741 ;
  assign n743 = n742 ^ n720 ;
  assign n738 = n712 ^ n710 ;
  assign n739 = n711 & ~n738 ;
  assign n740 = n739 ^ n709 ;
  assign n744 = n743 ^ n740 ;
  assign n748 = n747 ^ n744 ;
  assign n734 = n705 ^ n703 ;
  assign n735 = n704 & ~n734 ;
  assign n736 = n735 ^ n702 ;
  assign n730 = n698 ^ n696 ;
  assign n731 = n697 & ~n730 ;
  assign n732 = n731 ^ n695 ;
  assign n727 = n706 ^ n699 ;
  assign n728 = ~n701 & n727 ;
  assign n729 = n728 ^ n706 ;
  assign n733 = n732 ^ n729 ;
  assign n737 = n736 ^ n733 ;
  assign n749 = n748 ^ n737 ;
  assign n753 = n752 ^ n749 ;
  assign n754 = n753 ^ n690 ;
  assign n755 = n726 & ~n754 ;
  assign n756 = n755 ^ n725 ;
  assign n758 = n757 ^ n756 ;
  assign n766 = n747 ^ n743 ;
  assign n767 = n744 & n766 ;
  assign n768 = n767 ^ n743 ;
  assign n762 = n736 ^ n732 ;
  assign n763 = n733 & ~n762 ;
  assign n764 = n763 ^ n729 ;
  assign n759 = n752 ^ n737 ;
  assign n760 = ~n749 & n759 ;
  assign n761 = n760 ^ n752 ;
  assign n765 = n764 ^ n761 ;
  assign n769 = n768 ^ n765 ;
  assign n770 = n769 ^ n756 ;
  assign n771 = ~n758 & n770 ;
  assign n772 = n771 ^ n769 ;
  assign n687 = n686 ^ n682 ;
  assign n688 = n683 & ~n687 ;
  assign n689 = n688 ^ n647 ;
  assign n773 = n772 ^ n689 ;
  assign n774 = n768 ^ n764 ;
  assign n775 = n765 & ~n774 ;
  assign n776 = n775 ^ n761 ;
  assign n777 = n776 ^ n772 ;
  assign n778 = n773 & ~n777 ;
  assign n779 = n778 ^ n689 ;
  assign n780 = n769 ^ n758 ;
  assign n781 = n753 ^ n726 ;
  assign n782 = x256 ^ x192 ;
  assign n783 = n722 ^ n693 ;
  assign n784 = n782 & n783 ;
  assign n785 = n781 & n784 ;
  assign n786 = n780 & n785 ;
  assign n787 = n776 ^ n773 ;
  assign n788 = n786 & n787 ;
  assign n790 = ~n779 & ~n788 ;
  assign n789 = n788 ^ n779 ;
  assign n791 = n790 ^ n789 ;
  assign n792 = ~n622 & ~n791 ;
  assign n793 = n792 ^ n622 ;
  assign n794 = n455 & n793 ;
  assign n795 = n793 ^ n791 ;
  assign n796 = n795 ^ n622 ;
  assign n797 = n794 & n796 ;
  assign n798 = n797 ^ n794 ;
  assign n799 = n798 ^ n796 ;
  assign n800 = n799 ^ n794 ;
  assign n801 = n793 ^ n455 ;
  assign n802 = n801 ^ n794 ;
  assign n901 = x258 ^ x130 ;
  assign n898 = x266 ^ x138 ;
  assign n896 = x272 ^ x144 ;
  assign n894 = x270 ^ x142 ;
  assign n893 = x271 ^ x143 ;
  assign n895 = n894 ^ n893 ;
  assign n897 = n896 ^ n895 ;
  assign n899 = n898 ^ n897 ;
  assign n891 = x269 ^ x141 ;
  assign n889 = x267 ^ x139 ;
  assign n888 = x268 ^ x140 ;
  assign n890 = n889 ^ n888 ;
  assign n892 = n891 ^ n890 ;
  assign n900 = n899 ^ n892 ;
  assign n902 = n901 ^ n900 ;
  assign n885 = x259 ^ x131 ;
  assign n883 = x265 ^ x137 ;
  assign n881 = x263 ^ x135 ;
  assign n880 = x264 ^ x136 ;
  assign n882 = n881 ^ n880 ;
  assign n884 = n883 ^ n882 ;
  assign n886 = n885 ^ n884 ;
  assign n878 = x262 ^ x134 ;
  assign n876 = x260 ^ x132 ;
  assign n875 = x261 ^ x133 ;
  assign n877 = n876 ^ n875 ;
  assign n879 = n878 ^ n877 ;
  assign n887 = n886 ^ n879 ;
  assign n930 = n901 ^ n887 ;
  assign n931 = n902 & ~n930 ;
  assign n932 = n931 ^ n900 ;
  assign n926 = n891 ^ n889 ;
  assign n927 = n890 & ~n926 ;
  assign n928 = n927 ^ n888 ;
  assign n922 = n896 ^ n894 ;
  assign n923 = n895 & ~n922 ;
  assign n924 = n923 ^ n893 ;
  assign n919 = n897 ^ n892 ;
  assign n920 = ~n899 & n919 ;
  assign n921 = n920 ^ n892 ;
  assign n925 = n924 ^ n921 ;
  assign n929 = n928 ^ n925 ;
  assign n933 = n932 ^ n929 ;
  assign n915 = n878 ^ n876 ;
  assign n916 = n877 & ~n915 ;
  assign n917 = n916 ^ n875 ;
  assign n911 = n884 ^ n879 ;
  assign n912 = ~n886 & n911 ;
  assign n913 = n912 ^ n879 ;
  assign n908 = n883 ^ n881 ;
  assign n909 = n882 & ~n908 ;
  assign n910 = n909 ^ n880 ;
  assign n914 = n913 ^ n910 ;
  assign n918 = n917 ^ n914 ;
  assign n945 = n932 ^ n918 ;
  assign n946 = n933 & ~n945 ;
  assign n947 = n946 ^ n929 ;
  assign n942 = n928 ^ n924 ;
  assign n943 = n925 & ~n942 ;
  assign n944 = n943 ^ n921 ;
  assign n948 = n947 ^ n944 ;
  assign n939 = n917 ^ n913 ;
  assign n940 = n914 & ~n939 ;
  assign n941 = n940 ^ n910 ;
  assign n954 = n944 ^ n941 ;
  assign n955 = ~n948 & n954 ;
  assign n956 = n955 ^ n941 ;
  assign n873 = x257 ^ x129 ;
  assign n839 = x277 ^ x149 ;
  assign n837 = x275 ^ x147 ;
  assign n836 = x276 ^ x148 ;
  assign n838 = n837 ^ n836 ;
  assign n840 = n839 ^ n838 ;
  assign n834 = x274 ^ x146 ;
  assign n832 = x280 ^ x152 ;
  assign n830 = x278 ^ x150 ;
  assign n829 = x279 ^ x151 ;
  assign n831 = n830 ^ n829 ;
  assign n833 = n832 ^ n831 ;
  assign n835 = n834 ^ n833 ;
  assign n841 = n840 ^ n835 ;
  assign n812 = x282 ^ x154 ;
  assign n811 = x283 ^ x155 ;
  assign n813 = n812 ^ n811 ;
  assign n810 = x284 ^ x156 ;
  assign n814 = n813 ^ n810 ;
  assign n808 = x281 ^ x153 ;
  assign n805 = x285 ^ x157 ;
  assign n804 = x286 ^ x158 ;
  assign n806 = n805 ^ n804 ;
  assign n803 = x287 ^ x159 ;
  assign n807 = n806 ^ n803 ;
  assign n809 = n808 ^ n807 ;
  assign n827 = n814 ^ n809 ;
  assign n826 = x273 ^ x145 ;
  assign n828 = n827 ^ n826 ;
  assign n872 = n841 ^ n828 ;
  assign n874 = n873 ^ n872 ;
  assign n903 = n902 ^ n887 ;
  assign n904 = n903 ^ n873 ;
  assign n905 = n874 & ~n904 ;
  assign n906 = n905 ^ n872 ;
  assign n853 = n839 ^ n837 ;
  assign n854 = n838 & ~n853 ;
  assign n855 = n854 ^ n836 ;
  assign n849 = n832 ^ n830 ;
  assign n850 = n831 & ~n849 ;
  assign n851 = n850 ^ n829 ;
  assign n846 = n840 ^ n834 ;
  assign n847 = n835 & ~n846 ;
  assign n848 = n847 ^ n833 ;
  assign n852 = n851 ^ n848 ;
  assign n856 = n855 ^ n852 ;
  assign n842 = n841 ^ n827 ;
  assign n843 = n828 & ~n842 ;
  assign n844 = n843 ^ n826 ;
  assign n822 = n811 ^ n810 ;
  assign n823 = ~n813 & n822 ;
  assign n824 = n823 ^ n810 ;
  assign n818 = n804 ^ n803 ;
  assign n819 = ~n806 & n818 ;
  assign n820 = n819 ^ n803 ;
  assign n815 = n814 ^ n808 ;
  assign n816 = n809 & ~n815 ;
  assign n817 = n816 ^ n807 ;
  assign n821 = n820 ^ n817 ;
  assign n825 = n824 ^ n821 ;
  assign n845 = n844 ^ n825 ;
  assign n871 = n856 ^ n845 ;
  assign n907 = n906 ^ n871 ;
  assign n934 = n933 ^ n918 ;
  assign n935 = n934 ^ n871 ;
  assign n936 = n907 & ~n935 ;
  assign n937 = n936 ^ n906 ;
  assign n864 = n855 ^ n851 ;
  assign n865 = n852 & ~n864 ;
  assign n866 = n865 ^ n848 ;
  assign n860 = n824 ^ n820 ;
  assign n861 = n821 & ~n860 ;
  assign n862 = n861 ^ n817 ;
  assign n857 = n856 ^ n844 ;
  assign n858 = n845 & ~n857 ;
  assign n859 = n858 ^ n825 ;
  assign n863 = n862 ^ n859 ;
  assign n870 = n866 ^ n863 ;
  assign n938 = n937 ^ n870 ;
  assign n949 = n948 ^ n941 ;
  assign n950 = n949 ^ n937 ;
  assign n951 = n938 & ~n950 ;
  assign n952 = n951 ^ n870 ;
  assign n867 = n866 ^ n862 ;
  assign n868 = n863 & ~n867 ;
  assign n869 = n868 ^ n859 ;
  assign n953 = n952 ^ n869 ;
  assign n957 = n956 ^ n953 ;
  assign n958 = n934 ^ n907 ;
  assign n959 = n903 ^ n874 ;
  assign n960 = x256 ^ x128 ;
  assign n961 = n959 & n960 ;
  assign n962 = n958 & n961 ;
  assign n963 = n949 ^ n938 ;
  assign n964 = n962 & n963 ;
  assign n965 = n957 & n964 ;
  assign n966 = n956 ^ n952 ;
  assign n967 = n953 & ~n966 ;
  assign n968 = n967 ^ n869 ;
  assign n969 = n965 & n968 ;
  assign n970 = n802 & ~n969 ;
  assign n971 = n970 ^ n802 ;
  assign n972 = ~n800 & n971 ;
  assign n973 = ~n798 & n972 ;
  assign n974 = n973 ^ n972 ;
  assign n975 = n974 ^ n798 ;
  assign n976 = n975 ^ n972 ;
  assign n977 = n971 ^ n800 ;
  assign n978 = n977 ^ n972 ;
  assign n1077 = x258 ^ x98 ;
  assign n1074 = x266 ^ x106 ;
  assign n1072 = x272 ^ x112 ;
  assign n1070 = x270 ^ x110 ;
  assign n1069 = x271 ^ x111 ;
  assign n1071 = n1070 ^ n1069 ;
  assign n1073 = n1072 ^ n1071 ;
  assign n1075 = n1074 ^ n1073 ;
  assign n1067 = x269 ^ x109 ;
  assign n1065 = x267 ^ x107 ;
  assign n1064 = x268 ^ x108 ;
  assign n1066 = n1065 ^ n1064 ;
  assign n1068 = n1067 ^ n1066 ;
  assign n1076 = n1075 ^ n1068 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1061 = x259 ^ x99 ;
  assign n1059 = x265 ^ x105 ;
  assign n1057 = x263 ^ x103 ;
  assign n1056 = x264 ^ x104 ;
  assign n1058 = n1057 ^ n1056 ;
  assign n1060 = n1059 ^ n1058 ;
  assign n1062 = n1061 ^ n1060 ;
  assign n1054 = x262 ^ x102 ;
  assign n1052 = x260 ^ x100 ;
  assign n1051 = x261 ^ x101 ;
  assign n1053 = n1052 ^ n1051 ;
  assign n1055 = n1054 ^ n1053 ;
  assign n1063 = n1062 ^ n1055 ;
  assign n1106 = n1077 ^ n1063 ;
  assign n1107 = n1078 & ~n1106 ;
  assign n1108 = n1107 ^ n1076 ;
  assign n1102 = n1067 ^ n1065 ;
  assign n1103 = n1066 & ~n1102 ;
  assign n1104 = n1103 ^ n1064 ;
  assign n1098 = n1072 ^ n1070 ;
  assign n1099 = n1071 & ~n1098 ;
  assign n1100 = n1099 ^ n1069 ;
  assign n1095 = n1073 ^ n1068 ;
  assign n1096 = ~n1075 & n1095 ;
  assign n1097 = n1096 ^ n1068 ;
  assign n1101 = n1100 ^ n1097 ;
  assign n1105 = n1104 ^ n1101 ;
  assign n1109 = n1108 ^ n1105 ;
  assign n1091 = n1054 ^ n1052 ;
  assign n1092 = n1053 & ~n1091 ;
  assign n1093 = n1092 ^ n1051 ;
  assign n1087 = n1060 ^ n1055 ;
  assign n1088 = ~n1062 & n1087 ;
  assign n1089 = n1088 ^ n1055 ;
  assign n1084 = n1059 ^ n1057 ;
  assign n1085 = n1058 & ~n1084 ;
  assign n1086 = n1085 ^ n1056 ;
  assign n1090 = n1089 ^ n1086 ;
  assign n1094 = n1093 ^ n1090 ;
  assign n1121 = n1108 ^ n1094 ;
  assign n1122 = n1109 & ~n1121 ;
  assign n1123 = n1122 ^ n1105 ;
  assign n1118 = n1104 ^ n1100 ;
  assign n1119 = n1101 & ~n1118 ;
  assign n1120 = n1119 ^ n1097 ;
  assign n1124 = n1123 ^ n1120 ;
  assign n1115 = n1093 ^ n1089 ;
  assign n1116 = n1090 & ~n1115 ;
  assign n1117 = n1116 ^ n1086 ;
  assign n1130 = n1120 ^ n1117 ;
  assign n1131 = ~n1124 & n1130 ;
  assign n1132 = n1131 ^ n1117 ;
  assign n1049 = x257 ^ x97 ;
  assign n1015 = x277 ^ x117 ;
  assign n1013 = x275 ^ x115 ;
  assign n1012 = x276 ^ x116 ;
  assign n1014 = n1013 ^ n1012 ;
  assign n1016 = n1015 ^ n1014 ;
  assign n1010 = x274 ^ x114 ;
  assign n1008 = x280 ^ x120 ;
  assign n1006 = x278 ^ x118 ;
  assign n1005 = x279 ^ x119 ;
  assign n1007 = n1006 ^ n1005 ;
  assign n1009 = n1008 ^ n1007 ;
  assign n1011 = n1010 ^ n1009 ;
  assign n1017 = n1016 ^ n1011 ;
  assign n988 = x282 ^ x122 ;
  assign n987 = x283 ^ x123 ;
  assign n989 = n988 ^ n987 ;
  assign n986 = x284 ^ x124 ;
  assign n990 = n989 ^ n986 ;
  assign n984 = x281 ^ x121 ;
  assign n981 = x285 ^ x125 ;
  assign n980 = x286 ^ x126 ;
  assign n982 = n981 ^ n980 ;
  assign n979 = x287 ^ x127 ;
  assign n983 = n982 ^ n979 ;
  assign n985 = n984 ^ n983 ;
  assign n1003 = n990 ^ n985 ;
  assign n1002 = x273 ^ x113 ;
  assign n1004 = n1003 ^ n1002 ;
  assign n1048 = n1017 ^ n1004 ;
  assign n1050 = n1049 ^ n1048 ;
  assign n1079 = n1078 ^ n1063 ;
  assign n1080 = n1079 ^ n1049 ;
  assign n1081 = n1050 & ~n1080 ;
  assign n1082 = n1081 ^ n1048 ;
  assign n1029 = n1015 ^ n1013 ;
  assign n1030 = n1014 & ~n1029 ;
  assign n1031 = n1030 ^ n1012 ;
  assign n1025 = n1008 ^ n1006 ;
  assign n1026 = n1007 & ~n1025 ;
  assign n1027 = n1026 ^ n1005 ;
  assign n1022 = n1016 ^ n1010 ;
  assign n1023 = n1011 & ~n1022 ;
  assign n1024 = n1023 ^ n1009 ;
  assign n1028 = n1027 ^ n1024 ;
  assign n1032 = n1031 ^ n1028 ;
  assign n1018 = n1017 ^ n1003 ;
  assign n1019 = n1004 & ~n1018 ;
  assign n1020 = n1019 ^ n1002 ;
  assign n998 = n987 ^ n986 ;
  assign n999 = ~n989 & n998 ;
  assign n1000 = n999 ^ n986 ;
  assign n994 = n980 ^ n979 ;
  assign n995 = ~n982 & n994 ;
  assign n996 = n995 ^ n979 ;
  assign n991 = n990 ^ n984 ;
  assign n992 = n985 & ~n991 ;
  assign n993 = n992 ^ n983 ;
  assign n997 = n996 ^ n993 ;
  assign n1001 = n1000 ^ n997 ;
  assign n1021 = n1020 ^ n1001 ;
  assign n1047 = n1032 ^ n1021 ;
  assign n1083 = n1082 ^ n1047 ;
  assign n1110 = n1109 ^ n1094 ;
  assign n1111 = n1110 ^ n1047 ;
  assign n1112 = n1083 & ~n1111 ;
  assign n1113 = n1112 ^ n1082 ;
  assign n1040 = n1031 ^ n1027 ;
  assign n1041 = n1028 & ~n1040 ;
  assign n1042 = n1041 ^ n1024 ;
  assign n1036 = n1000 ^ n996 ;
  assign n1037 = n997 & ~n1036 ;
  assign n1038 = n1037 ^ n993 ;
  assign n1033 = n1032 ^ n1020 ;
  assign n1034 = n1021 & ~n1033 ;
  assign n1035 = n1034 ^ n1001 ;
  assign n1039 = n1038 ^ n1035 ;
  assign n1046 = n1042 ^ n1039 ;
  assign n1114 = n1113 ^ n1046 ;
  assign n1125 = n1124 ^ n1117 ;
  assign n1126 = n1125 ^ n1113 ;
  assign n1127 = n1114 & ~n1126 ;
  assign n1128 = n1127 ^ n1046 ;
  assign n1043 = n1042 ^ n1038 ;
  assign n1044 = n1039 & ~n1043 ;
  assign n1045 = n1044 ^ n1035 ;
  assign n1129 = n1128 ^ n1045 ;
  assign n1133 = n1132 ^ n1129 ;
  assign n1134 = n1110 ^ n1083 ;
  assign n1135 = n1079 ^ n1050 ;
  assign n1136 = x256 ^ x96 ;
  assign n1137 = n1135 & n1136 ;
  assign n1138 = n1134 & n1137 ;
  assign n1139 = n1125 ^ n1114 ;
  assign n1140 = n1138 & n1139 ;
  assign n1141 = n1133 & n1140 ;
  assign n1142 = n1132 ^ n1128 ;
  assign n1143 = n1129 & ~n1142 ;
  assign n1144 = n1143 ^ n1045 ;
  assign n1145 = n1141 & n1144 ;
  assign n1146 = ~n978 & ~n1145 ;
  assign n1147 = n1146 ^ n978 ;
  assign n1148 = n976 & ~n1147 ;
  assign n1149 = n974 & ~n1148 ;
  assign n1150 = n1149 ^ n1148 ;
  assign n1151 = n1147 ^ n976 ;
  assign n1152 = n1151 ^ n1148 ;
  assign n1251 = x258 ^ x66 ;
  assign n1248 = x266 ^ x74 ;
  assign n1246 = x272 ^ x80 ;
  assign n1244 = x270 ^ x78 ;
  assign n1243 = x271 ^ x79 ;
  assign n1245 = n1244 ^ n1243 ;
  assign n1247 = n1246 ^ n1245 ;
  assign n1249 = n1248 ^ n1247 ;
  assign n1241 = x269 ^ x77 ;
  assign n1239 = x267 ^ x75 ;
  assign n1238 = x268 ^ x76 ;
  assign n1240 = n1239 ^ n1238 ;
  assign n1242 = n1241 ^ n1240 ;
  assign n1250 = n1249 ^ n1242 ;
  assign n1252 = n1251 ^ n1250 ;
  assign n1235 = x259 ^ x67 ;
  assign n1233 = x265 ^ x73 ;
  assign n1231 = x263 ^ x71 ;
  assign n1230 = x264 ^ x72 ;
  assign n1232 = n1231 ^ n1230 ;
  assign n1234 = n1233 ^ n1232 ;
  assign n1236 = n1235 ^ n1234 ;
  assign n1228 = x262 ^ x70 ;
  assign n1226 = x260 ^ x68 ;
  assign n1225 = x261 ^ x69 ;
  assign n1227 = n1226 ^ n1225 ;
  assign n1229 = n1228 ^ n1227 ;
  assign n1237 = n1236 ^ n1229 ;
  assign n1280 = n1251 ^ n1237 ;
  assign n1281 = n1252 & ~n1280 ;
  assign n1282 = n1281 ^ n1250 ;
  assign n1276 = n1241 ^ n1239 ;
  assign n1277 = n1240 & ~n1276 ;
  assign n1278 = n1277 ^ n1238 ;
  assign n1272 = n1246 ^ n1244 ;
  assign n1273 = n1245 & ~n1272 ;
  assign n1274 = n1273 ^ n1243 ;
  assign n1269 = n1247 ^ n1242 ;
  assign n1270 = ~n1249 & n1269 ;
  assign n1271 = n1270 ^ n1242 ;
  assign n1275 = n1274 ^ n1271 ;
  assign n1279 = n1278 ^ n1275 ;
  assign n1283 = n1282 ^ n1279 ;
  assign n1265 = n1228 ^ n1226 ;
  assign n1266 = n1227 & ~n1265 ;
  assign n1267 = n1266 ^ n1225 ;
  assign n1261 = n1234 ^ n1229 ;
  assign n1262 = ~n1236 & n1261 ;
  assign n1263 = n1262 ^ n1229 ;
  assign n1258 = n1233 ^ n1231 ;
  assign n1259 = n1232 & ~n1258 ;
  assign n1260 = n1259 ^ n1230 ;
  assign n1264 = n1263 ^ n1260 ;
  assign n1268 = n1267 ^ n1264 ;
  assign n1295 = n1282 ^ n1268 ;
  assign n1296 = n1283 & ~n1295 ;
  assign n1297 = n1296 ^ n1279 ;
  assign n1292 = n1278 ^ n1274 ;
  assign n1293 = n1275 & ~n1292 ;
  assign n1294 = n1293 ^ n1271 ;
  assign n1298 = n1297 ^ n1294 ;
  assign n1289 = n1267 ^ n1263 ;
  assign n1290 = n1264 & ~n1289 ;
  assign n1291 = n1290 ^ n1260 ;
  assign n1304 = n1294 ^ n1291 ;
  assign n1305 = ~n1298 & n1304 ;
  assign n1306 = n1305 ^ n1291 ;
  assign n1223 = x257 ^ x65 ;
  assign n1189 = x277 ^ x85 ;
  assign n1187 = x275 ^ x83 ;
  assign n1186 = x276 ^ x84 ;
  assign n1188 = n1187 ^ n1186 ;
  assign n1190 = n1189 ^ n1188 ;
  assign n1184 = x274 ^ x82 ;
  assign n1182 = x280 ^ x88 ;
  assign n1180 = x278 ^ x86 ;
  assign n1179 = x279 ^ x87 ;
  assign n1181 = n1180 ^ n1179 ;
  assign n1183 = n1182 ^ n1181 ;
  assign n1185 = n1184 ^ n1183 ;
  assign n1191 = n1190 ^ n1185 ;
  assign n1162 = x282 ^ x90 ;
  assign n1161 = x283 ^ x91 ;
  assign n1163 = n1162 ^ n1161 ;
  assign n1160 = x284 ^ x92 ;
  assign n1164 = n1163 ^ n1160 ;
  assign n1158 = x281 ^ x89 ;
  assign n1155 = x285 ^ x93 ;
  assign n1154 = x286 ^ x94 ;
  assign n1156 = n1155 ^ n1154 ;
  assign n1153 = x287 ^ x95 ;
  assign n1157 = n1156 ^ n1153 ;
  assign n1159 = n1158 ^ n1157 ;
  assign n1177 = n1164 ^ n1159 ;
  assign n1176 = x273 ^ x81 ;
  assign n1178 = n1177 ^ n1176 ;
  assign n1222 = n1191 ^ n1178 ;
  assign n1224 = n1223 ^ n1222 ;
  assign n1253 = n1252 ^ n1237 ;
  assign n1254 = n1253 ^ n1223 ;
  assign n1255 = n1224 & ~n1254 ;
  assign n1256 = n1255 ^ n1222 ;
  assign n1203 = n1189 ^ n1187 ;
  assign n1204 = n1188 & ~n1203 ;
  assign n1205 = n1204 ^ n1186 ;
  assign n1199 = n1182 ^ n1180 ;
  assign n1200 = n1181 & ~n1199 ;
  assign n1201 = n1200 ^ n1179 ;
  assign n1196 = n1190 ^ n1184 ;
  assign n1197 = n1185 & ~n1196 ;
  assign n1198 = n1197 ^ n1183 ;
  assign n1202 = n1201 ^ n1198 ;
  assign n1206 = n1205 ^ n1202 ;
  assign n1192 = n1191 ^ n1177 ;
  assign n1193 = n1178 & ~n1192 ;
  assign n1194 = n1193 ^ n1176 ;
  assign n1172 = n1161 ^ n1160 ;
  assign n1173 = ~n1163 & n1172 ;
  assign n1174 = n1173 ^ n1160 ;
  assign n1168 = n1154 ^ n1153 ;
  assign n1169 = ~n1156 & n1168 ;
  assign n1170 = n1169 ^ n1153 ;
  assign n1165 = n1164 ^ n1158 ;
  assign n1166 = n1159 & ~n1165 ;
  assign n1167 = n1166 ^ n1157 ;
  assign n1171 = n1170 ^ n1167 ;
  assign n1175 = n1174 ^ n1171 ;
  assign n1195 = n1194 ^ n1175 ;
  assign n1221 = n1206 ^ n1195 ;
  assign n1257 = n1256 ^ n1221 ;
  assign n1284 = n1283 ^ n1268 ;
  assign n1285 = n1284 ^ n1221 ;
  assign n1286 = n1257 & ~n1285 ;
  assign n1287 = n1286 ^ n1256 ;
  assign n1214 = n1205 ^ n1201 ;
  assign n1215 = n1202 & ~n1214 ;
  assign n1216 = n1215 ^ n1198 ;
  assign n1210 = n1174 ^ n1170 ;
  assign n1211 = n1171 & ~n1210 ;
  assign n1212 = n1211 ^ n1167 ;
  assign n1207 = n1206 ^ n1194 ;
  assign n1208 = n1195 & ~n1207 ;
  assign n1209 = n1208 ^ n1175 ;
  assign n1213 = n1212 ^ n1209 ;
  assign n1220 = n1216 ^ n1213 ;
  assign n1288 = n1287 ^ n1220 ;
  assign n1299 = n1298 ^ n1291 ;
  assign n1300 = n1299 ^ n1287 ;
  assign n1301 = n1288 & ~n1300 ;
  assign n1302 = n1301 ^ n1220 ;
  assign n1217 = n1216 ^ n1212 ;
  assign n1218 = n1213 & ~n1217 ;
  assign n1219 = n1218 ^ n1209 ;
  assign n1303 = n1302 ^ n1219 ;
  assign n1307 = n1306 ^ n1303 ;
  assign n1308 = n1284 ^ n1257 ;
  assign n1309 = n1253 ^ n1224 ;
  assign n1310 = x256 ^ x64 ;
  assign n1311 = n1309 & n1310 ;
  assign n1312 = n1308 & n1311 ;
  assign n1313 = n1299 ^ n1288 ;
  assign n1314 = n1312 & n1313 ;
  assign n1315 = n1307 & n1314 ;
  assign n1316 = n1306 ^ n1302 ;
  assign n1317 = n1303 & ~n1316 ;
  assign n1318 = n1317 ^ n1219 ;
  assign n1319 = n1315 & n1318 ;
  assign n1320 = ~n1152 & ~n1319 ;
  assign n1321 = n1320 ^ n1152 ;
  assign n1322 = n1150 & ~n1321 ;
  assign n1494 = n1149 ^ n974 ;
  assign n1495 = n1322 & ~n1494 ;
  assign n1496 = n1495 ^ n1322 ;
  assign n1497 = n1496 ^ n1494 ;
  assign n1498 = n1497 ^ n1322 ;
  assign n1323 = n1321 ^ n1150 ;
  assign n1324 = n1323 ^ n1322 ;
  assign n1423 = x258 ^ x34 ;
  assign n1420 = x266 ^ x42 ;
  assign n1418 = x272 ^ x48 ;
  assign n1416 = x270 ^ x46 ;
  assign n1415 = x271 ^ x47 ;
  assign n1417 = n1416 ^ n1415 ;
  assign n1419 = n1418 ^ n1417 ;
  assign n1421 = n1420 ^ n1419 ;
  assign n1413 = x269 ^ x45 ;
  assign n1411 = x267 ^ x43 ;
  assign n1410 = x268 ^ x44 ;
  assign n1412 = n1411 ^ n1410 ;
  assign n1414 = n1413 ^ n1412 ;
  assign n1422 = n1421 ^ n1414 ;
  assign n1424 = n1423 ^ n1422 ;
  assign n1407 = x259 ^ x35 ;
  assign n1405 = x265 ^ x41 ;
  assign n1403 = x263 ^ x39 ;
  assign n1402 = x264 ^ x40 ;
  assign n1404 = n1403 ^ n1402 ;
  assign n1406 = n1405 ^ n1404 ;
  assign n1408 = n1407 ^ n1406 ;
  assign n1400 = x262 ^ x38 ;
  assign n1398 = x260 ^ x36 ;
  assign n1397 = x261 ^ x37 ;
  assign n1399 = n1398 ^ n1397 ;
  assign n1401 = n1400 ^ n1399 ;
  assign n1409 = n1408 ^ n1401 ;
  assign n1452 = n1423 ^ n1409 ;
  assign n1453 = n1424 & ~n1452 ;
  assign n1454 = n1453 ^ n1422 ;
  assign n1448 = n1413 ^ n1411 ;
  assign n1449 = n1412 & ~n1448 ;
  assign n1450 = n1449 ^ n1410 ;
  assign n1444 = n1418 ^ n1416 ;
  assign n1445 = n1417 & ~n1444 ;
  assign n1446 = n1445 ^ n1415 ;
  assign n1441 = n1419 ^ n1414 ;
  assign n1442 = ~n1421 & n1441 ;
  assign n1443 = n1442 ^ n1414 ;
  assign n1447 = n1446 ^ n1443 ;
  assign n1451 = n1450 ^ n1447 ;
  assign n1455 = n1454 ^ n1451 ;
  assign n1437 = n1400 ^ n1398 ;
  assign n1438 = n1399 & ~n1437 ;
  assign n1439 = n1438 ^ n1397 ;
  assign n1433 = n1406 ^ n1401 ;
  assign n1434 = ~n1408 & n1433 ;
  assign n1435 = n1434 ^ n1401 ;
  assign n1430 = n1405 ^ n1403 ;
  assign n1431 = n1404 & ~n1430 ;
  assign n1432 = n1431 ^ n1402 ;
  assign n1436 = n1435 ^ n1432 ;
  assign n1440 = n1439 ^ n1436 ;
  assign n1467 = n1454 ^ n1440 ;
  assign n1468 = n1455 & ~n1467 ;
  assign n1469 = n1468 ^ n1451 ;
  assign n1464 = n1450 ^ n1446 ;
  assign n1465 = n1447 & ~n1464 ;
  assign n1466 = n1465 ^ n1443 ;
  assign n1470 = n1469 ^ n1466 ;
  assign n1461 = n1439 ^ n1435 ;
  assign n1462 = n1436 & ~n1461 ;
  assign n1463 = n1462 ^ n1432 ;
  assign n1476 = n1466 ^ n1463 ;
  assign n1477 = ~n1470 & n1476 ;
  assign n1478 = n1477 ^ n1463 ;
  assign n1395 = x257 ^ x33 ;
  assign n1361 = x277 ^ x53 ;
  assign n1359 = x275 ^ x51 ;
  assign n1358 = x276 ^ x52 ;
  assign n1360 = n1359 ^ n1358 ;
  assign n1362 = n1361 ^ n1360 ;
  assign n1356 = x274 ^ x50 ;
  assign n1354 = x280 ^ x56 ;
  assign n1352 = x278 ^ x54 ;
  assign n1351 = x279 ^ x55 ;
  assign n1353 = n1352 ^ n1351 ;
  assign n1355 = n1354 ^ n1353 ;
  assign n1357 = n1356 ^ n1355 ;
  assign n1363 = n1362 ^ n1357 ;
  assign n1334 = x282 ^ x58 ;
  assign n1333 = x283 ^ x59 ;
  assign n1335 = n1334 ^ n1333 ;
  assign n1332 = x284 ^ x60 ;
  assign n1336 = n1335 ^ n1332 ;
  assign n1330 = x281 ^ x57 ;
  assign n1327 = x285 ^ x61 ;
  assign n1326 = x286 ^ x62 ;
  assign n1328 = n1327 ^ n1326 ;
  assign n1325 = x287 ^ x63 ;
  assign n1329 = n1328 ^ n1325 ;
  assign n1331 = n1330 ^ n1329 ;
  assign n1349 = n1336 ^ n1331 ;
  assign n1348 = x273 ^ x49 ;
  assign n1350 = n1349 ^ n1348 ;
  assign n1394 = n1363 ^ n1350 ;
  assign n1396 = n1395 ^ n1394 ;
  assign n1425 = n1424 ^ n1409 ;
  assign n1426 = n1425 ^ n1395 ;
  assign n1427 = n1396 & ~n1426 ;
  assign n1428 = n1427 ^ n1394 ;
  assign n1375 = n1361 ^ n1359 ;
  assign n1376 = n1360 & ~n1375 ;
  assign n1377 = n1376 ^ n1358 ;
  assign n1371 = n1354 ^ n1352 ;
  assign n1372 = n1353 & ~n1371 ;
  assign n1373 = n1372 ^ n1351 ;
  assign n1368 = n1362 ^ n1356 ;
  assign n1369 = n1357 & ~n1368 ;
  assign n1370 = n1369 ^ n1355 ;
  assign n1374 = n1373 ^ n1370 ;
  assign n1378 = n1377 ^ n1374 ;
  assign n1364 = n1363 ^ n1349 ;
  assign n1365 = n1350 & ~n1364 ;
  assign n1366 = n1365 ^ n1348 ;
  assign n1344 = n1333 ^ n1332 ;
  assign n1345 = ~n1335 & n1344 ;
  assign n1346 = n1345 ^ n1332 ;
  assign n1340 = n1326 ^ n1325 ;
  assign n1341 = ~n1328 & n1340 ;
  assign n1342 = n1341 ^ n1325 ;
  assign n1337 = n1336 ^ n1330 ;
  assign n1338 = n1331 & ~n1337 ;
  assign n1339 = n1338 ^ n1329 ;
  assign n1343 = n1342 ^ n1339 ;
  assign n1347 = n1346 ^ n1343 ;
  assign n1367 = n1366 ^ n1347 ;
  assign n1393 = n1378 ^ n1367 ;
  assign n1429 = n1428 ^ n1393 ;
  assign n1456 = n1455 ^ n1440 ;
  assign n1457 = n1456 ^ n1393 ;
  assign n1458 = n1429 & ~n1457 ;
  assign n1459 = n1458 ^ n1428 ;
  assign n1386 = n1377 ^ n1373 ;
  assign n1387 = n1374 & ~n1386 ;
  assign n1388 = n1387 ^ n1370 ;
  assign n1382 = n1346 ^ n1342 ;
  assign n1383 = n1343 & ~n1382 ;
  assign n1384 = n1383 ^ n1339 ;
  assign n1379 = n1378 ^ n1366 ;
  assign n1380 = n1367 & ~n1379 ;
  assign n1381 = n1380 ^ n1347 ;
  assign n1385 = n1384 ^ n1381 ;
  assign n1392 = n1388 ^ n1385 ;
  assign n1460 = n1459 ^ n1392 ;
  assign n1471 = n1470 ^ n1463 ;
  assign n1472 = n1471 ^ n1459 ;
  assign n1473 = n1460 & ~n1472 ;
  assign n1474 = n1473 ^ n1392 ;
  assign n1389 = n1388 ^ n1384 ;
  assign n1390 = n1385 & ~n1389 ;
  assign n1391 = n1390 ^ n1381 ;
  assign n1475 = n1474 ^ n1391 ;
  assign n1479 = n1478 ^ n1475 ;
  assign n1480 = n1456 ^ n1429 ;
  assign n1481 = n1425 ^ n1396 ;
  assign n1482 = x256 ^ x32 ;
  assign n1483 = n1481 & n1482 ;
  assign n1484 = n1480 & n1483 ;
  assign n1485 = n1471 ^ n1460 ;
  assign n1486 = n1484 & n1485 ;
  assign n1487 = n1479 & n1486 ;
  assign n1488 = n1478 ^ n1474 ;
  assign n1489 = n1475 & ~n1488 ;
  assign n1490 = n1489 ^ n1391 ;
  assign n1491 = n1487 & n1490 ;
  assign n1492 = ~n1324 & ~n1491 ;
  assign n1493 = n1492 ^ n1324 ;
  assign n2014 = n1498 ^ n1493 ;
  assign n1499 = ~n1493 & n1498 ;
  assign n2165 = n2014 ^ n1499 ;
  assign n2264 = x258 ^ x2 ;
  assign n2261 = x266 ^ x10 ;
  assign n2259 = x272 ^ x16 ;
  assign n2257 = x270 ^ x14 ;
  assign n2256 = x271 ^ x15 ;
  assign n2258 = n2257 ^ n2256 ;
  assign n2260 = n2259 ^ n2258 ;
  assign n2262 = n2261 ^ n2260 ;
  assign n2254 = x269 ^ x13 ;
  assign n2252 = x267 ^ x11 ;
  assign n2251 = x268 ^ x12 ;
  assign n2253 = n2252 ^ n2251 ;
  assign n2255 = n2254 ^ n2253 ;
  assign n2263 = n2262 ^ n2255 ;
  assign n2265 = n2264 ^ n2263 ;
  assign n2248 = x259 ^ x3 ;
  assign n2246 = x265 ^ x9 ;
  assign n2244 = x263 ^ x7 ;
  assign n2243 = x264 ^ x8 ;
  assign n2245 = n2244 ^ n2243 ;
  assign n2247 = n2246 ^ n2245 ;
  assign n2249 = n2248 ^ n2247 ;
  assign n2241 = x262 ^ x6 ;
  assign n2239 = x260 ^ x4 ;
  assign n2238 = x261 ^ x5 ;
  assign n2240 = n2239 ^ n2238 ;
  assign n2242 = n2241 ^ n2240 ;
  assign n2250 = n2249 ^ n2242 ;
  assign n2293 = n2264 ^ n2250 ;
  assign n2294 = n2265 & ~n2293 ;
  assign n2295 = n2294 ^ n2263 ;
  assign n2289 = n2254 ^ n2252 ;
  assign n2290 = n2253 & ~n2289 ;
  assign n2291 = n2290 ^ n2251 ;
  assign n2285 = n2259 ^ n2257 ;
  assign n2286 = n2258 & ~n2285 ;
  assign n2287 = n2286 ^ n2256 ;
  assign n2282 = n2260 ^ n2255 ;
  assign n2283 = ~n2262 & n2282 ;
  assign n2284 = n2283 ^ n2255 ;
  assign n2288 = n2287 ^ n2284 ;
  assign n2292 = n2291 ^ n2288 ;
  assign n2296 = n2295 ^ n2292 ;
  assign n2278 = n2241 ^ n2239 ;
  assign n2279 = n2240 & ~n2278 ;
  assign n2280 = n2279 ^ n2238 ;
  assign n2274 = n2247 ^ n2242 ;
  assign n2275 = ~n2249 & n2274 ;
  assign n2276 = n2275 ^ n2242 ;
  assign n2271 = n2246 ^ n2244 ;
  assign n2272 = n2245 & ~n2271 ;
  assign n2273 = n2272 ^ n2243 ;
  assign n2277 = n2276 ^ n2273 ;
  assign n2281 = n2280 ^ n2277 ;
  assign n2308 = n2295 ^ n2281 ;
  assign n2309 = n2296 & ~n2308 ;
  assign n2310 = n2309 ^ n2292 ;
  assign n2305 = n2291 ^ n2287 ;
  assign n2306 = n2288 & ~n2305 ;
  assign n2307 = n2306 ^ n2284 ;
  assign n2311 = n2310 ^ n2307 ;
  assign n2302 = n2280 ^ n2276 ;
  assign n2303 = n2277 & ~n2302 ;
  assign n2304 = n2303 ^ n2273 ;
  assign n2317 = n2307 ^ n2304 ;
  assign n2318 = ~n2311 & n2317 ;
  assign n2319 = n2318 ^ n2304 ;
  assign n2236 = x257 ^ x1 ;
  assign n2202 = x277 ^ x21 ;
  assign n2200 = x275 ^ x19 ;
  assign n2199 = x276 ^ x20 ;
  assign n2201 = n2200 ^ n2199 ;
  assign n2203 = n2202 ^ n2201 ;
  assign n2197 = x274 ^ x18 ;
  assign n2195 = x280 ^ x24 ;
  assign n2193 = x278 ^ x22 ;
  assign n2192 = x279 ^ x23 ;
  assign n2194 = n2193 ^ n2192 ;
  assign n2196 = n2195 ^ n2194 ;
  assign n2198 = n2197 ^ n2196 ;
  assign n2204 = n2203 ^ n2198 ;
  assign n2175 = x282 ^ x26 ;
  assign n2174 = x283 ^ x27 ;
  assign n2176 = n2175 ^ n2174 ;
  assign n2173 = x284 ^ x28 ;
  assign n2177 = n2176 ^ n2173 ;
  assign n2171 = x281 ^ x25 ;
  assign n2168 = x285 ^ x29 ;
  assign n2167 = x286 ^ x30 ;
  assign n2169 = n2168 ^ n2167 ;
  assign n2166 = x287 ^ x31 ;
  assign n2170 = n2169 ^ n2166 ;
  assign n2172 = n2171 ^ n2170 ;
  assign n2190 = n2177 ^ n2172 ;
  assign n2189 = x273 ^ x17 ;
  assign n2191 = n2190 ^ n2189 ;
  assign n2235 = n2204 ^ n2191 ;
  assign n2237 = n2236 ^ n2235 ;
  assign n2266 = n2265 ^ n2250 ;
  assign n2267 = n2266 ^ n2236 ;
  assign n2268 = n2237 & ~n2267 ;
  assign n2269 = n2268 ^ n2235 ;
  assign n2216 = n2202 ^ n2200 ;
  assign n2217 = n2201 & ~n2216 ;
  assign n2218 = n2217 ^ n2199 ;
  assign n2212 = n2195 ^ n2193 ;
  assign n2213 = n2194 & ~n2212 ;
  assign n2214 = n2213 ^ n2192 ;
  assign n2209 = n2203 ^ n2197 ;
  assign n2210 = n2198 & ~n2209 ;
  assign n2211 = n2210 ^ n2196 ;
  assign n2215 = n2214 ^ n2211 ;
  assign n2219 = n2218 ^ n2215 ;
  assign n2205 = n2204 ^ n2190 ;
  assign n2206 = n2191 & ~n2205 ;
  assign n2207 = n2206 ^ n2189 ;
  assign n2185 = n2174 ^ n2173 ;
  assign n2186 = ~n2176 & n2185 ;
  assign n2187 = n2186 ^ n2173 ;
  assign n2181 = n2167 ^ n2166 ;
  assign n2182 = ~n2169 & n2181 ;
  assign n2183 = n2182 ^ n2166 ;
  assign n2178 = n2177 ^ n2171 ;
  assign n2179 = n2172 & ~n2178 ;
  assign n2180 = n2179 ^ n2170 ;
  assign n2184 = n2183 ^ n2180 ;
  assign n2188 = n2187 ^ n2184 ;
  assign n2208 = n2207 ^ n2188 ;
  assign n2234 = n2219 ^ n2208 ;
  assign n2270 = n2269 ^ n2234 ;
  assign n2297 = n2296 ^ n2281 ;
  assign n2298 = n2297 ^ n2234 ;
  assign n2299 = n2270 & ~n2298 ;
  assign n2300 = n2299 ^ n2269 ;
  assign n2227 = n2218 ^ n2214 ;
  assign n2228 = n2215 & ~n2227 ;
  assign n2229 = n2228 ^ n2211 ;
  assign n2223 = n2187 ^ n2183 ;
  assign n2224 = n2184 & ~n2223 ;
  assign n2225 = n2224 ^ n2180 ;
  assign n2220 = n2219 ^ n2207 ;
  assign n2221 = n2208 & ~n2220 ;
  assign n2222 = n2221 ^ n2188 ;
  assign n2226 = n2225 ^ n2222 ;
  assign n2233 = n2229 ^ n2226 ;
  assign n2301 = n2300 ^ n2233 ;
  assign n2312 = n2311 ^ n2304 ;
  assign n2313 = n2312 ^ n2300 ;
  assign n2314 = n2301 & ~n2313 ;
  assign n2315 = n2314 ^ n2233 ;
  assign n2230 = n2229 ^ n2225 ;
  assign n2231 = n2226 & ~n2230 ;
  assign n2232 = n2231 ^ n2222 ;
  assign n2316 = n2315 ^ n2232 ;
  assign n2320 = n2319 ^ n2316 ;
  assign n2321 = n2297 ^ n2270 ;
  assign n2322 = n2266 ^ n2237 ;
  assign n2323 = x256 ^ x0 ;
  assign n2324 = n2322 & n2323 ;
  assign n2325 = n2321 & n2324 ;
  assign n2326 = n2312 ^ n2301 ;
  assign n2327 = n2325 & n2326 ;
  assign n2328 = n2320 & n2327 ;
  assign n2329 = n2319 ^ n2315 ;
  assign n2330 = n2316 & ~n2329 ;
  assign n2331 = n2330 ^ n2232 ;
  assign n2332 = n2328 & n2331 ;
  assign n2333 = ~n2165 & ~n2332 ;
  assign n2334 = n2333 ^ n2165 ;
  assign n2161 = ~n1496 & n1499 ;
  assign n2162 = n2161 ^ n1499 ;
  assign n2163 = n2162 ^ n1496 ;
  assign n2164 = n2163 ^ n1499 ;
  assign n2335 = n2334 ^ n2164 ;
  assign n1537 = n454 ^ n451 ;
  assign n1505 = n621 ^ n618 ;
  assign n1506 = n1505 ^ n789 ;
  assign n1507 = n789 & ~n1505 ;
  assign n1508 = n1507 ^ n792 ;
  assign n1509 = n1507 ^ n1506 ;
  assign n1511 = n787 ^ n786 ;
  assign n1510 = n617 ^ n606 ;
  assign n1512 = n1511 ^ n1510 ;
  assign n1514 = n605 ^ n600 ;
  assign n1513 = n785 ^ n780 ;
  assign n1515 = n1514 ^ n1513 ;
  assign n1517 = n603 ^ n602 ;
  assign n1518 = n783 ^ n782 ;
  assign n1519 = ~n1517 & n1518 ;
  assign n1516 = n604 ^ n601 ;
  assign n1520 = n1519 ^ n1516 ;
  assign n1521 = n784 ^ n781 ;
  assign n1522 = n1521 ^ n1519 ;
  assign n1523 = ~n1520 & ~n1522 ;
  assign n1524 = n1523 ^ n1516 ;
  assign n1525 = n1524 ^ n1513 ;
  assign n1526 = ~n1515 & n1525 ;
  assign n1527 = n1526 ^ n1514 ;
  assign n1528 = n1527 ^ n1510 ;
  assign n1529 = ~n1512 & n1528 ;
  assign n1530 = n1529 ^ n1510 ;
  assign n1531 = ~n1509 & ~n1530 ;
  assign n1532 = ~n1508 & ~n1531 ;
  assign n1533 = n795 & ~n1532 ;
  assign n1534 = n1506 & ~n1533 ;
  assign n1504 = n789 ^ n622 ;
  assign n1535 = n1534 ^ n1504 ;
  assign n1536 = n1535 ^ n622 ;
  assign n1538 = n1537 ^ n1536 ;
  assign n1571 = n1536 ^ n455 ;
  assign n1540 = n1512 & ~n1533 ;
  assign n1541 = n1540 ^ n1511 ;
  assign n1539 = n450 ^ n443 ;
  assign n1542 = n1541 ^ n1539 ;
  assign n1546 = n449 ^ n448 ;
  assign n1543 = n1515 & ~n1533 ;
  assign n1544 = n1543 ^ n1515 ;
  assign n1545 = n1544 ^ n1514 ;
  assign n1547 = n1546 ^ n1545 ;
  assign n1552 = n447 ^ n444 ;
  assign n1548 = n1521 ^ n1516 ;
  assign n1549 = n1533 & n1548 ;
  assign n1550 = n1549 ^ n1548 ;
  assign n1551 = n1550 ^ n1521 ;
  assign n1553 = n1552 ^ n1551 ;
  assign n1554 = n446 ^ n445 ;
  assign n1555 = n1518 ^ n1517 ;
  assign n1556 = ~n1533 & n1555 ;
  assign n1557 = n1556 ^ n1555 ;
  assign n1558 = n1557 ^ n1517 ;
  assign n1559 = n1554 & ~n1558 ;
  assign n1560 = n1559 ^ n1551 ;
  assign n1561 = ~n1553 & ~n1560 ;
  assign n1562 = n1561 ^ n1551 ;
  assign n1563 = n1562 ^ n1545 ;
  assign n1564 = ~n1547 & n1563 ;
  assign n1565 = n1564 ^ n1545 ;
  assign n1566 = n1565 ^ n1539 ;
  assign n1567 = ~n1542 & ~n1566 ;
  assign n1568 = n1567 ^ n1539 ;
  assign n1569 = n1568 ^ n1537 ;
  assign n1570 = ~n1538 & ~n1569 ;
  assign n1572 = n1571 ^ n1570 ;
  assign n1573 = ~n801 & n1572 ;
  assign n1574 = n1573 ^ n793 ;
  assign n1575 = n1538 & n1574 ;
  assign n1615 = n1575 ^ n1536 ;
  assign n1614 = n1534 ^ n1505 ;
  assign n1616 = n1615 ^ n1614 ;
  assign n1617 = ~n1614 & n1615 ;
  assign n1618 = n1617 ^ n797 ;
  assign n1619 = n1617 ^ n1616 ;
  assign n1621 = n1540 ^ n1510 ;
  assign n1582 = n1542 & n1574 ;
  assign n1620 = n1582 ^ n1541 ;
  assign n1622 = n1621 ^ n1620 ;
  assign n1625 = n1543 ^ n1514 ;
  assign n1586 = n1547 & n1574 ;
  assign n1623 = n1586 ^ n1547 ;
  assign n1624 = n1623 ^ n1546 ;
  assign n1626 = n1625 ^ n1624 ;
  assign n1589 = n1553 & n1574 ;
  assign n1628 = n1589 ^ n1553 ;
  assign n1629 = n1628 ^ n1552 ;
  assign n1627 = n1549 ^ n1521 ;
  assign n1630 = n1629 ^ n1627 ;
  assign n1631 = n1556 ^ n1517 ;
  assign n1594 = n1558 ^ n1554 ;
  assign n1595 = n1574 & n1594 ;
  assign n1632 = n1595 ^ n1594 ;
  assign n1633 = n1632 ^ n1554 ;
  assign n1634 = ~n1631 & n1633 ;
  assign n1635 = n1634 ^ n1627 ;
  assign n1636 = ~n1630 & ~n1635 ;
  assign n1637 = n1636 ^ n1627 ;
  assign n1638 = n1637 ^ n1624 ;
  assign n1639 = ~n1626 & ~n1638 ;
  assign n1640 = n1639 ^ n1624 ;
  assign n1641 = n1640 ^ n1620 ;
  assign n1642 = ~n1622 & n1641 ;
  assign n1643 = n1642 ^ n1620 ;
  assign n1644 = ~n1619 & n1643 ;
  assign n1645 = ~n1618 & ~n1644 ;
  assign n1646 = n799 & ~n1645 ;
  assign n1647 = n1616 & ~n1646 ;
  assign n1730 = n1647 ^ n1614 ;
  assign n1648 = n1647 ^ n1615 ;
  assign n1577 = n968 ^ n965 ;
  assign n1576 = n1575 ^ n1537 ;
  assign n1578 = n1577 ^ n1576 ;
  assign n1579 = n1576 & ~n1577 ;
  assign n1580 = ~n970 & ~n1579 ;
  assign n1583 = n1582 ^ n1539 ;
  assign n1581 = n964 ^ n957 ;
  assign n1584 = n1583 ^ n1581 ;
  assign n1587 = n1586 ^ n1546 ;
  assign n1585 = n963 ^ n962 ;
  assign n1588 = n1587 ^ n1585 ;
  assign n1591 = n961 ^ n958 ;
  assign n1590 = n1589 ^ n1552 ;
  assign n1592 = n1591 ^ n1590 ;
  assign n1593 = n960 ^ n959 ;
  assign n1596 = n1595 ^ n1554 ;
  assign n1597 = n1593 & ~n1596 ;
  assign n1598 = n1597 ^ n1590 ;
  assign n1599 = ~n1592 & ~n1598 ;
  assign n1600 = n1599 ^ n1590 ;
  assign n1601 = n1600 ^ n1587 ;
  assign n1602 = ~n1588 & ~n1601 ;
  assign n1603 = n1602 ^ n1585 ;
  assign n1604 = n1603 ^ n1581 ;
  assign n1605 = ~n1584 & n1604 ;
  assign n1606 = n1605 ^ n1581 ;
  assign n1607 = n1580 & n1606 ;
  assign n1608 = n1578 ^ n969 ;
  assign n1609 = n1608 ^ n1579 ;
  assign n1610 = ~n802 & n1609 ;
  assign n1611 = ~n1607 & ~n1610 ;
  assign n1612 = n1578 & ~n1611 ;
  assign n1613 = n1612 ^ n1577 ;
  assign n1649 = n1648 ^ n1613 ;
  assign n1652 = n1584 & n1611 ;
  assign n1653 = n1652 ^ n1583 ;
  assign n1650 = n1622 & ~n1646 ;
  assign n1651 = n1650 ^ n1620 ;
  assign n1654 = n1653 ^ n1651 ;
  assign n1657 = n1626 & ~n1646 ;
  assign n1658 = n1657 ^ n1626 ;
  assign n1659 = n1658 ^ n1625 ;
  assign n1655 = n1588 & ~n1611 ;
  assign n1656 = n1655 ^ n1585 ;
  assign n1660 = n1659 ^ n1656 ;
  assign n1663 = n1630 & n1646 ;
  assign n1664 = n1663 ^ n1630 ;
  assign n1665 = n1664 ^ n1629 ;
  assign n1661 = n1592 & ~n1611 ;
  assign n1662 = n1661 ^ n1591 ;
  assign n1666 = n1665 ^ n1662 ;
  assign n1667 = n1596 ^ n1593 ;
  assign n1668 = ~n1611 & n1667 ;
  assign n1669 = n1668 ^ n1593 ;
  assign n1670 = n1633 ^ n1631 ;
  assign n1671 = ~n1646 & n1670 ;
  assign n1672 = n1671 ^ n1670 ;
  assign n1673 = n1672 ^ n1631 ;
  assign n1674 = n1669 & ~n1673 ;
  assign n1675 = n1674 ^ n1662 ;
  assign n1676 = ~n1666 & n1675 ;
  assign n1677 = n1676 ^ n1662 ;
  assign n1678 = n1677 ^ n1656 ;
  assign n1679 = ~n1660 & n1678 ;
  assign n1680 = n1679 ^ n1656 ;
  assign n1681 = n1680 ^ n1651 ;
  assign n1682 = ~n1654 & n1681 ;
  assign n1683 = n1682 ^ n1653 ;
  assign n1684 = n1683 ^ n1648 ;
  assign n1685 = ~n1649 & n1684 ;
  assign n1686 = n1685 ^ n1613 ;
  assign n1687 = n1686 ^ n971 ;
  assign n1688 = n977 & ~n1687 ;
  assign n1689 = n1688 ^ n800 ;
  assign n1690 = n1649 & ~n1689 ;
  assign n1691 = n1690 ^ n1613 ;
  assign n1728 = n1691 ^ n1648 ;
  assign n1729 = n1728 ^ n1613 ;
  assign n1731 = n1730 ^ n1729 ;
  assign n1732 = n972 ^ n798 ;
  assign n1735 = n1650 ^ n1621 ;
  assign n1695 = n1654 & n1689 ;
  assign n1733 = n1695 ^ n1654 ;
  assign n1734 = n1733 ^ n1651 ;
  assign n1736 = n1735 ^ n1734 ;
  assign n1739 = n1657 ^ n1625 ;
  assign n1700 = n1660 & n1689 ;
  assign n1737 = n1700 ^ n1660 ;
  assign n1738 = n1737 ^ n1659 ;
  assign n1740 = n1739 ^ n1738 ;
  assign n1743 = n1663 ^ n1629 ;
  assign n1703 = n1666 & n1689 ;
  assign n1741 = n1703 ^ n1666 ;
  assign n1742 = n1741 ^ n1665 ;
  assign n1744 = n1743 ^ n1742 ;
  assign n1708 = n1673 ^ n1669 ;
  assign n1709 = ~n1689 & n1708 ;
  assign n1745 = n1709 ^ n1708 ;
  assign n1746 = n1745 ^ n1669 ;
  assign n1747 = n1671 ^ n1631 ;
  assign n1748 = n1746 & ~n1747 ;
  assign n1749 = n1748 ^ n1742 ;
  assign n1750 = ~n1744 & n1749 ;
  assign n1751 = n1750 ^ n1742 ;
  assign n1752 = n1751 ^ n1738 ;
  assign n1753 = ~n1740 & n1752 ;
  assign n1754 = n1753 ^ n1738 ;
  assign n1755 = n1754 ^ n1734 ;
  assign n1756 = ~n1736 & n1755 ;
  assign n1757 = n1756 ^ n1734 ;
  assign n1758 = n1757 ^ n1729 ;
  assign n1759 = ~n1731 & n1758 ;
  assign n1760 = n1759 ^ n1729 ;
  assign n1761 = n1760 ^ n972 ;
  assign n1762 = ~n1732 & ~n1761 ;
  assign n1763 = n1762 ^ n798 ;
  assign n1764 = n1731 & n1763 ;
  assign n1849 = n1764 ^ n1730 ;
  assign n1765 = n1764 ^ n1729 ;
  assign n1503 = n1144 ^ n1141 ;
  assign n1692 = n1691 ^ n1503 ;
  assign n1693 = ~n1503 & n1691 ;
  assign n1694 = ~n1146 & ~n1693 ;
  assign n1697 = n1140 ^ n1133 ;
  assign n1696 = n1695 ^ n1651 ;
  assign n1698 = n1697 ^ n1696 ;
  assign n1701 = n1700 ^ n1659 ;
  assign n1699 = n1139 ^ n1138 ;
  assign n1702 = n1701 ^ n1699 ;
  assign n1705 = n1137 ^ n1134 ;
  assign n1704 = n1703 ^ n1665 ;
  assign n1706 = n1705 ^ n1704 ;
  assign n1707 = n1136 ^ n1135 ;
  assign n1710 = n1709 ^ n1669 ;
  assign n1711 = n1707 & ~n1710 ;
  assign n1712 = n1711 ^ n1704 ;
  assign n1713 = ~n1706 & ~n1712 ;
  assign n1714 = n1713 ^ n1704 ;
  assign n1715 = n1714 ^ n1701 ;
  assign n1716 = ~n1702 & ~n1715 ;
  assign n1717 = n1716 ^ n1699 ;
  assign n1718 = n1717 ^ n1696 ;
  assign n1719 = ~n1698 & ~n1718 ;
  assign n1720 = n1719 ^ n1696 ;
  assign n1721 = n1694 & ~n1720 ;
  assign n1722 = n1692 ^ n1145 ;
  assign n1723 = n1722 ^ n1693 ;
  assign n1724 = n978 & n1723 ;
  assign n1725 = ~n1721 & ~n1724 ;
  assign n1726 = n1692 & n1725 ;
  assign n1727 = n1726 ^ n1691 ;
  assign n1766 = n1765 ^ n1727 ;
  assign n1769 = ~n1734 & n1735 ;
  assign n1772 = n1763 & n1769 ;
  assign n1773 = n1772 ^ n1734 ;
  assign n1770 = n1769 ^ n1736 ;
  assign n1771 = n1763 & n1770 ;
  assign n1774 = n1773 ^ n1771 ;
  assign n1767 = n1698 & ~n1725 ;
  assign n1768 = n1767 ^ n1697 ;
  assign n1775 = n1774 ^ n1768 ;
  assign n1779 = n1702 & ~n1725 ;
  assign n1780 = n1779 ^ n1699 ;
  assign n1776 = n1740 & n1763 ;
  assign n1777 = n1776 ^ n1740 ;
  assign n1778 = n1777 ^ n1739 ;
  assign n1781 = n1780 ^ n1778 ;
  assign n1784 = n1744 & n1763 ;
  assign n1785 = n1784 ^ n1744 ;
  assign n1786 = n1785 ^ n1743 ;
  assign n1782 = n1706 & ~n1725 ;
  assign n1783 = n1782 ^ n1705 ;
  assign n1787 = n1786 ^ n1783 ;
  assign n1788 = n1710 ^ n1707 ;
  assign n1789 = ~n1725 & n1788 ;
  assign n1790 = n1789 ^ n1707 ;
  assign n1791 = n1747 ^ n1746 ;
  assign n1792 = ~n1763 & n1791 ;
  assign n1793 = n1792 ^ n1791 ;
  assign n1794 = n1793 ^ n1746 ;
  assign n1795 = n1790 & ~n1794 ;
  assign n1796 = n1795 ^ n1783 ;
  assign n1797 = ~n1787 & n1796 ;
  assign n1798 = n1797 ^ n1783 ;
  assign n1799 = n1798 ^ n1778 ;
  assign n1800 = ~n1781 & ~n1799 ;
  assign n1801 = n1800 ^ n1778 ;
  assign n1802 = n1801 ^ n1774 ;
  assign n1803 = ~n1775 & ~n1802 ;
  assign n1804 = n1803 ^ n1768 ;
  assign n1805 = n1804 ^ n1765 ;
  assign n1806 = ~n1766 & n1805 ;
  assign n1807 = n1806 ^ n1727 ;
  assign n1808 = n1807 ^ n1147 ;
  assign n1809 = n1151 & n1808 ;
  assign n1810 = n1809 ^ n976 ;
  assign n1811 = n1766 & n1810 ;
  assign n1812 = n1811 ^ n1727 ;
  assign n1850 = n1812 ^ n1765 ;
  assign n1851 = n1850 ^ n1727 ;
  assign n1889 = ~n1849 & n1851 ;
  assign n1890 = n1149 & n1889 ;
  assign n1852 = n1851 ^ n1849 ;
  assign n1853 = n1148 ^ n974 ;
  assign n1856 = n1772 ^ n1771 ;
  assign n1857 = n1856 ^ n1735 ;
  assign n1819 = n1775 & ~n1810 ;
  assign n1854 = n1819 ^ n1775 ;
  assign n1855 = n1854 ^ n1774 ;
  assign n1858 = n1857 ^ n1855 ;
  assign n1823 = n1781 & ~n1810 ;
  assign n1860 = n1823 ^ n1781 ;
  assign n1861 = n1860 ^ n1778 ;
  assign n1859 = n1776 ^ n1739 ;
  assign n1862 = n1861 ^ n1859 ;
  assign n1827 = n1787 & ~n1810 ;
  assign n1864 = n1827 ^ n1787 ;
  assign n1865 = n1864 ^ n1786 ;
  assign n1863 = n1784 ^ n1743 ;
  assign n1866 = n1865 ^ n1863 ;
  assign n1867 = n1792 ^ n1746 ;
  assign n1832 = n1794 ^ n1790 ;
  assign n1833 = n1810 & n1832 ;
  assign n1868 = n1833 ^ n1832 ;
  assign n1869 = n1868 ^ n1790 ;
  assign n1870 = ~n1867 & n1869 ;
  assign n1871 = n1870 ^ n1865 ;
  assign n1872 = ~n1866 & n1871 ;
  assign n1873 = n1872 ^ n1865 ;
  assign n1874 = n1873 ^ n1859 ;
  assign n1875 = ~n1862 & ~n1874 ;
  assign n1876 = n1875 ^ n1859 ;
  assign n1877 = n1876 ^ n1855 ;
  assign n1878 = ~n1858 & ~n1877 ;
  assign n1879 = n1878 ^ n1855 ;
  assign n1880 = n1879 ^ n1851 ;
  assign n1881 = ~n1852 & ~n1880 ;
  assign n1882 = n1881 ^ n1849 ;
  assign n1883 = n1882 ^ n974 ;
  assign n1884 = ~n1853 & ~n1883 ;
  assign n1885 = n1884 ^ n1148 ;
  assign n1886 = n1852 & ~n1885 ;
  assign n1887 = n1849 & ~n1886 ;
  assign n1888 = n1887 ^ n1852 ;
  assign n1891 = n1890 ^ n1888 ;
  assign n1502 = n1318 ^ n1315 ;
  assign n1813 = n1812 ^ n1502 ;
  assign n1815 = ~n1502 & n1812 ;
  assign n1814 = n1813 ^ n1319 ;
  assign n1816 = n1815 ^ n1814 ;
  assign n1817 = n1152 & n1816 ;
  assign n1818 = ~n1320 & ~n1815 ;
  assign n1821 = n1314 ^ n1307 ;
  assign n1820 = n1819 ^ n1774 ;
  assign n1822 = n1821 ^ n1820 ;
  assign n1825 = n1313 ^ n1312 ;
  assign n1824 = n1823 ^ n1778 ;
  assign n1826 = n1825 ^ n1824 ;
  assign n1829 = n1311 ^ n1308 ;
  assign n1828 = n1827 ^ n1786 ;
  assign n1830 = n1829 ^ n1828 ;
  assign n1831 = n1310 ^ n1309 ;
  assign n1834 = n1833 ^ n1790 ;
  assign n1835 = n1831 & ~n1834 ;
  assign n1836 = n1835 ^ n1828 ;
  assign n1837 = ~n1830 & ~n1836 ;
  assign n1838 = n1837 ^ n1828 ;
  assign n1839 = n1838 ^ n1825 ;
  assign n1840 = ~n1826 & ~n1839 ;
  assign n1841 = n1840 ^ n1825 ;
  assign n1842 = n1841 ^ n1820 ;
  assign n1843 = ~n1822 & ~n1842 ;
  assign n1844 = n1843 ^ n1820 ;
  assign n1845 = n1818 & ~n1844 ;
  assign n1846 = ~n1817 & ~n1845 ;
  assign n1847 = n1813 & ~n1846 ;
  assign n1848 = n1847 ^ n1502 ;
  assign n1892 = n1891 ^ n1848 ;
  assign n1895 = n1858 & ~n1885 ;
  assign n1896 = n1895 ^ n1855 ;
  assign n1893 = n1822 & ~n1846 ;
  assign n1894 = n1893 ^ n1821 ;
  assign n1897 = n1896 ^ n1894 ;
  assign n1901 = n1826 & ~n1846 ;
  assign n1902 = n1901 ^ n1825 ;
  assign n1898 = n1862 & ~n1885 ;
  assign n1899 = n1898 ^ n1862 ;
  assign n1900 = n1899 ^ n1859 ;
  assign n1903 = n1902 ^ n1900 ;
  assign n1906 = n1866 & n1885 ;
  assign n1907 = n1906 ^ n1866 ;
  assign n1908 = n1907 ^ n1865 ;
  assign n1904 = n1830 & ~n1846 ;
  assign n1905 = n1904 ^ n1829 ;
  assign n1909 = n1908 ^ n1905 ;
  assign n1910 = n1834 ^ n1831 ;
  assign n1911 = ~n1846 & n1910 ;
  assign n1912 = n1911 ^ n1831 ;
  assign n1913 = n1869 ^ n1867 ;
  assign n1914 = ~n1885 & n1913 ;
  assign n1915 = n1914 ^ n1913 ;
  assign n1916 = n1915 ^ n1867 ;
  assign n1917 = n1912 & ~n1916 ;
  assign n1918 = n1917 ^ n1905 ;
  assign n1919 = ~n1909 & n1918 ;
  assign n1920 = n1919 ^ n1905 ;
  assign n1921 = n1920 ^ n1900 ;
  assign n1922 = ~n1903 & ~n1921 ;
  assign n1923 = n1922 ^ n1900 ;
  assign n1924 = n1923 ^ n1894 ;
  assign n1925 = ~n1897 & n1924 ;
  assign n1926 = n1925 ^ n1896 ;
  assign n1927 = n1926 ^ n1891 ;
  assign n1928 = ~n1892 & ~n1927 ;
  assign n1929 = n1928 ^ n1848 ;
  assign n1930 = n1929 ^ n1150 ;
  assign n1931 = n1323 & n1930 ;
  assign n1932 = n1931 ^ n1321 ;
  assign n1933 = n1892 & n1932 ;
  assign n1934 = n1933 ^ n1848 ;
  assign n1972 = n1934 ^ n1891 ;
  assign n1973 = n1972 ^ n1848 ;
  assign n1974 = n1890 ^ n1887 ;
  assign n2007 = n1973 & ~n1974 ;
  assign n2011 = n1497 & n2007 ;
  assign n2059 = n2011 ^ n1974 ;
  assign n1971 = n1494 ^ n1322 ;
  assign n1975 = n1974 ^ n1973 ;
  assign n1978 = n1895 ^ n1857 ;
  assign n1941 = n1897 & ~n1932 ;
  assign n1976 = n1941 ^ n1897 ;
  assign n1977 = n1976 ^ n1896 ;
  assign n1979 = n1978 ^ n1977 ;
  assign n1982 = n1898 ^ n1859 ;
  assign n1945 = n1903 & ~n1932 ;
  assign n1980 = n1945 ^ n1903 ;
  assign n1981 = n1980 ^ n1900 ;
  assign n1983 = n1982 ^ n1981 ;
  assign n1949 = n1909 & ~n1932 ;
  assign n1985 = n1949 ^ n1909 ;
  assign n1986 = n1985 ^ n1908 ;
  assign n1984 = n1906 ^ n1865 ;
  assign n1987 = n1986 ^ n1984 ;
  assign n1988 = n1914 ^ n1867 ;
  assign n1954 = n1916 ^ n1912 ;
  assign n1955 = n1932 & n1954 ;
  assign n1989 = n1955 ^ n1954 ;
  assign n1990 = n1989 ^ n1912 ;
  assign n1991 = ~n1988 & n1990 ;
  assign n1992 = n1991 ^ n1986 ;
  assign n1993 = ~n1987 & n1992 ;
  assign n1994 = n1993 ^ n1986 ;
  assign n1995 = n1994 ^ n1981 ;
  assign n1996 = ~n1983 & n1995 ;
  assign n1997 = n1996 ^ n1981 ;
  assign n1998 = n1997 ^ n1978 ;
  assign n1999 = ~n1979 & ~n1998 ;
  assign n2000 = n1999 ^ n1978 ;
  assign n2001 = n2000 ^ n1973 ;
  assign n2002 = ~n1975 & ~n2001 ;
  assign n2003 = n2002 ^ n1973 ;
  assign n2004 = n2003 ^ n1494 ;
  assign n2005 = ~n1971 & n2004 ;
  assign n2006 = n2005 ^ n1322 ;
  assign n2008 = n2007 ^ n1975 ;
  assign n2009 = ~n2006 & n2008 ;
  assign n2060 = n2059 ^ n2009 ;
  assign n2010 = n2009 ^ n1973 ;
  assign n2012 = n2011 ^ n2010 ;
  assign n1501 = n1490 ^ n1487 ;
  assign n1935 = n1934 ^ n1501 ;
  assign n1937 = ~n1501 & n1934 ;
  assign n1936 = n1935 ^ n1491 ;
  assign n1938 = n1937 ^ n1936 ;
  assign n1939 = n1324 & n1938 ;
  assign n1940 = ~n1492 & ~n1937 ;
  assign n1943 = n1486 ^ n1479 ;
  assign n1942 = n1941 ^ n1896 ;
  assign n1944 = n1943 ^ n1942 ;
  assign n1947 = n1485 ^ n1484 ;
  assign n1946 = n1945 ^ n1900 ;
  assign n1948 = n1947 ^ n1946 ;
  assign n1951 = n1483 ^ n1480 ;
  assign n1950 = n1949 ^ n1908 ;
  assign n1952 = n1951 ^ n1950 ;
  assign n1953 = n1482 ^ n1481 ;
  assign n1956 = n1955 ^ n1912 ;
  assign n1957 = n1953 & ~n1956 ;
  assign n1958 = n1957 ^ n1950 ;
  assign n1959 = ~n1952 & ~n1958 ;
  assign n1960 = n1959 ^ n1950 ;
  assign n1961 = n1960 ^ n1947 ;
  assign n1962 = ~n1948 & ~n1961 ;
  assign n1963 = n1962 ^ n1947 ;
  assign n1964 = n1963 ^ n1942 ;
  assign n1965 = ~n1944 & ~n1964 ;
  assign n1966 = n1965 ^ n1942 ;
  assign n1967 = n1940 & ~n1966 ;
  assign n1968 = ~n1939 & ~n1967 ;
  assign n1969 = n1935 & ~n1968 ;
  assign n1970 = n1969 ^ n1501 ;
  assign n2013 = n2012 ^ n1970 ;
  assign n2017 = n1944 & ~n1968 ;
  assign n2018 = n2017 ^ n1943 ;
  assign n2015 = n1979 & ~n2006 ;
  assign n2016 = n2015 ^ n1977 ;
  assign n2019 = n2018 ^ n2016 ;
  assign n2023 = n1948 & ~n1968 ;
  assign n2024 = n2023 ^ n1947 ;
  assign n2020 = n1983 & ~n2006 ;
  assign n2021 = n2020 ^ n1983 ;
  assign n2022 = n2021 ^ n1982 ;
  assign n2025 = n2024 ^ n2022 ;
  assign n2028 = n1987 & n2006 ;
  assign n2029 = n2028 ^ n1987 ;
  assign n2030 = n2029 ^ n1986 ;
  assign n2026 = n1952 & ~n1968 ;
  assign n2027 = n2026 ^ n1951 ;
  assign n2031 = n2030 ^ n2027 ;
  assign n2032 = n1956 ^ n1953 ;
  assign n2033 = ~n1968 & n2032 ;
  assign n2034 = n2033 ^ n1953 ;
  assign n2035 = n1990 ^ n1988 ;
  assign n2036 = ~n2006 & n2035 ;
  assign n2037 = n2036 ^ n2035 ;
  assign n2038 = n2037 ^ n1988 ;
  assign n2039 = n2034 & ~n2038 ;
  assign n2040 = n2039 ^ n2027 ;
  assign n2041 = ~n2031 & n2040 ;
  assign n2042 = n2041 ^ n2027 ;
  assign n2043 = n2042 ^ n2022 ;
  assign n2044 = ~n2025 & ~n2043 ;
  assign n2045 = n2044 ^ n2022 ;
  assign n2046 = n2045 ^ n2018 ;
  assign n2047 = ~n2019 & n2046 ;
  assign n2048 = n2047 ^ n2016 ;
  assign n2049 = n2048 ^ n2012 ;
  assign n2050 = ~n2013 & ~n2049 ;
  assign n2051 = n2050 ^ n1970 ;
  assign n2052 = n2051 ^ n1498 ;
  assign n2053 = n2014 & n2052 ;
  assign n2054 = n2053 ^ n1493 ;
  assign n2055 = n2013 & n2054 ;
  assign n2056 = n2055 ^ n1970 ;
  assign n2057 = n2056 ^ n2012 ;
  assign n2058 = n2057 ^ n1970 ;
  assign n2061 = n2060 ^ n2058 ;
  assign n1500 = n1499 ^ n1496 ;
  assign n2063 = n2019 & ~n2054 ;
  assign n2064 = n2063 ^ n2019 ;
  assign n2065 = n2064 ^ n2016 ;
  assign n2062 = n2015 ^ n1978 ;
  assign n2066 = n2065 ^ n2062 ;
  assign n2070 = n2020 ^ n1982 ;
  assign n2067 = n2025 & ~n2054 ;
  assign n2068 = n2067 ^ n2025 ;
  assign n2069 = n2068 ^ n2022 ;
  assign n2071 = n2070 ^ n2069 ;
  assign n2075 = n2028 ^ n1986 ;
  assign n2072 = n2031 & ~n2054 ;
  assign n2073 = n2072 ^ n2031 ;
  assign n2074 = n2073 ^ n2030 ;
  assign n2076 = n2075 ^ n2074 ;
  assign n2077 = n2036 ^ n1988 ;
  assign n2078 = n2038 ^ n2034 ;
  assign n2079 = n2054 & n2078 ;
  assign n2080 = n2079 ^ n2078 ;
  assign n2081 = n2080 ^ n2034 ;
  assign n2082 = ~n2077 & n2081 ;
  assign n2083 = n2082 ^ n2075 ;
  assign n2084 = ~n2076 & ~n2083 ;
  assign n2085 = n2084 ^ n2075 ;
  assign n2086 = n2085 ^ n2069 ;
  assign n2087 = ~n2071 & ~n2086 ;
  assign n2088 = n2087 ^ n2069 ;
  assign n2089 = n2088 ^ n2062 ;
  assign n2090 = ~n2066 & ~n2089 ;
  assign n2091 = n2090 ^ n2062 ;
  assign n2092 = n2091 ^ n2058 ;
  assign n2093 = ~n2061 & ~n2092 ;
  assign n2094 = n2093 ^ n2058 ;
  assign n2095 = n2094 ^ n1499 ;
  assign n2096 = ~n1500 & ~n2095 ;
  assign n2097 = n2096 ^ n1496 ;
  assign n2368 = n2061 & n2097 ;
  assign n2369 = n2368 ^ n2058 ;
  assign n2336 = n2331 ^ n2328 ;
  assign n2337 = n2336 ^ n2056 ;
  assign n2339 = n2056 & ~n2336 ;
  assign n2338 = n2337 ^ n2332 ;
  assign n2340 = n2339 ^ n2338 ;
  assign n2341 = n2165 & n2340 ;
  assign n2342 = ~n2333 & ~n2339 ;
  assign n2344 = n2063 ^ n2016 ;
  assign n2343 = n2327 ^ n2320 ;
  assign n2345 = n2344 ^ n2343 ;
  assign n2347 = n2326 ^ n2325 ;
  assign n2346 = n2067 ^ n2022 ;
  assign n2348 = n2347 ^ n2346 ;
  assign n2350 = n2072 ^ n2030 ;
  assign n2349 = n2324 ^ n2321 ;
  assign n2351 = n2350 ^ n2349 ;
  assign n2352 = n2323 ^ n2322 ;
  assign n2353 = n2079 ^ n2034 ;
  assign n2354 = n2352 & ~n2353 ;
  assign n2355 = n2354 ^ n2349 ;
  assign n2356 = ~n2351 & n2355 ;
  assign n2357 = n2356 ^ n2349 ;
  assign n2358 = n2357 ^ n2347 ;
  assign n2359 = ~n2348 & n2358 ;
  assign n2360 = n2359 ^ n2347 ;
  assign n2361 = n2360 ^ n2343 ;
  assign n2362 = ~n2345 & n2361 ;
  assign n2363 = n2362 ^ n2343 ;
  assign n2364 = n2342 & n2363 ;
  assign n2365 = ~n2341 & ~n2364 ;
  assign n2366 = n2337 & ~n2365 ;
  assign n2367 = n2366 ^ n2336 ;
  assign n2370 = n2369 ^ n2367 ;
  assign n2373 = n2345 & ~n2365 ;
  assign n2374 = n2373 ^ n2343 ;
  assign n2371 = n2066 & n2097 ;
  assign n2372 = n2371 ^ n2065 ;
  assign n2375 = n2374 ^ n2372 ;
  assign n2378 = n2071 & n2097 ;
  assign n2379 = n2378 ^ n2071 ;
  assign n2380 = n2379 ^ n2070 ;
  assign n2376 = n2348 & ~n2365 ;
  assign n2377 = n2376 ^ n2347 ;
  assign n2381 = n2380 ^ n2377 ;
  assign n2385 = n2351 & n2365 ;
  assign n2386 = n2385 ^ n2350 ;
  assign n2382 = n2076 & n2097 ;
  assign n2383 = n2382 ^ n2076 ;
  assign n2384 = n2383 ^ n2075 ;
  assign n2387 = n2386 ^ n2384 ;
  assign n2388 = n2353 ^ n2352 ;
  assign n2389 = ~n2365 & n2388 ;
  assign n2390 = n2389 ^ n2352 ;
  assign n2391 = n2081 ^ n2077 ;
  assign n2392 = n2097 & n2391 ;
  assign n2393 = n2392 ^ n2391 ;
  assign n2394 = n2393 ^ n2077 ;
  assign n2395 = n2390 & ~n2394 ;
  assign n2396 = n2395 ^ n2384 ;
  assign n2397 = ~n2387 & ~n2396 ;
  assign n2398 = n2397 ^ n2384 ;
  assign n2399 = n2398 ^ n2377 ;
  assign n2400 = ~n2381 & ~n2399 ;
  assign n2401 = n2400 ^ n2377 ;
  assign n2402 = n2401 ^ n2372 ;
  assign n2403 = ~n2375 & n2402 ;
  assign n2404 = n2403 ^ n2374 ;
  assign n2405 = n2404 ^ n2367 ;
  assign n2406 = ~n2370 & ~n2405 ;
  assign n2407 = n2406 ^ n2369 ;
  assign n2408 = n2407 ^ n2334 ;
  assign n2409 = n2335 & ~n2408 ;
  assign n2410 = n2409 ^ n2164 ;
  assign n2098 = x224 ^ x192 ;
  assign n2099 = n1533 & n2098 ;
  assign n2100 = n2099 ^ n2098 ;
  assign n2101 = n2100 ^ x192 ;
  assign n2102 = n2101 ^ x160 ;
  assign n2103 = n1574 & n2102 ;
  assign n2109 = n2103 ^ n2102 ;
  assign n2110 = n2109 ^ x160 ;
  assign n2108 = n2099 ^ x192 ;
  assign n2111 = n2110 ^ n2108 ;
  assign n2112 = ~n1646 & n2111 ;
  assign n2122 = n2112 ^ n2111 ;
  assign n2123 = n2122 ^ n2110 ;
  assign n2113 = n2112 ^ n2110 ;
  assign n2104 = n2103 ^ x160 ;
  assign n2105 = n2104 ^ x128 ;
  assign n2106 = ~n1611 & n2105 ;
  assign n2107 = n2106 ^ x128 ;
  assign n2114 = n2113 ^ n2107 ;
  assign n2115 = n1689 & n2114 ;
  assign n2120 = n2115 ^ n2114 ;
  assign n2121 = n2120 ^ n2113 ;
  assign n2124 = n2123 ^ n2121 ;
  assign n2125 = ~n1763 & n2124 ;
  assign n2135 = n2125 ^ n2124 ;
  assign n2136 = n2135 ^ n2123 ;
  assign n2126 = n2125 ^ n2123 ;
  assign n2116 = n2115 ^ n2113 ;
  assign n2117 = n2116 ^ x96 ;
  assign n2118 = ~n1725 & n2117 ;
  assign n2119 = n2118 ^ x96 ;
  assign n2127 = n2126 ^ n2119 ;
  assign n2128 = ~n1810 & n2127 ;
  assign n2133 = n2128 ^ n2127 ;
  assign n2134 = n2133 ^ n2126 ;
  assign n2137 = n2136 ^ n2134 ;
  assign n2138 = n1885 & n2137 ;
  assign n2144 = n2138 ^ n2137 ;
  assign n2145 = n2144 ^ n2136 ;
  assign n2139 = n2138 ^ n2136 ;
  assign n2129 = n2128 ^ n2126 ;
  assign n2130 = n2129 ^ x64 ;
  assign n2131 = ~n1846 & n2130 ;
  assign n2132 = n2131 ^ x64 ;
  assign n2140 = n2139 ^ n2132 ;
  assign n2141 = ~n1932 & n2140 ;
  assign n2142 = n2141 ^ n2140 ;
  assign n2143 = n2142 ^ n2139 ;
  assign n2146 = n2145 ^ n2143 ;
  assign n2147 = ~n2006 & n2146 ;
  assign n2153 = n2147 ^ n2146 ;
  assign n2154 = n2153 ^ n2145 ;
  assign n2149 = n2141 ^ n2139 ;
  assign n2150 = n2149 ^ x32 ;
  assign n2151 = ~n1968 & n2150 ;
  assign n2152 = n2151 ^ x32 ;
  assign n2155 = n2154 ^ n2152 ;
  assign n2156 = n2054 & n2155 ;
  assign n2413 = n2156 ^ n2155 ;
  assign n2414 = n2413 ^ n2154 ;
  assign n2415 = n2414 ^ x0 ;
  assign n2416 = ~n2365 & n2415 ;
  assign n2417 = n2416 ^ x0 ;
  assign n2157 = n2156 ^ n2154 ;
  assign n2148 = n2147 ^ n2145 ;
  assign n2158 = n2157 ^ n2148 ;
  assign n2159 = ~n2097 & n2158 ;
  assign n2411 = n2159 ^ n2158 ;
  assign n2412 = n2411 ^ n2157 ;
  assign n2418 = n2417 ^ n2412 ;
  assign n2419 = n2410 & n2418 ;
  assign n2420 = n2419 ^ n2418 ;
  assign n2421 = n2420 ^ n2417 ;
  assign n2160 = n2159 ^ n2157 ;
  assign n2422 = n2421 ^ n2160 ;
  assign n2423 = n2164 & ~n2334 ;
  assign n2424 = n2423 ^ n2162 ;
  assign n2429 = n2371 ^ n2062 ;
  assign n2427 = n2375 & n2410 ;
  assign n2428 = n2427 ^ n2372 ;
  assign n2430 = n2429 ^ n2428 ;
  assign n2433 = n2378 ^ n2070 ;
  assign n2431 = n2381 & n2410 ;
  assign n2432 = n2431 ^ n2380 ;
  assign n2434 = n2433 ^ n2432 ;
  assign n2437 = n2382 ^ n2075 ;
  assign n2435 = n2387 & ~n2410 ;
  assign n2436 = n2435 ^ n2386 ;
  assign n2438 = n2437 ^ n2436 ;
  assign n2439 = n2392 ^ n2077 ;
  assign n2440 = n2394 ^ n2390 ;
  assign n2441 = n2410 & n2440 ;
  assign n2442 = n2441 ^ n2394 ;
  assign n2443 = ~n2439 & n2442 ;
  assign n2444 = n2443 ^ n2436 ;
  assign n2445 = ~n2438 & n2444 ;
  assign n2446 = n2445 ^ n2436 ;
  assign n2447 = n2446 ^ n2433 ;
  assign n2448 = ~n2434 & n2447 ;
  assign n2449 = n2448 ^ n2432 ;
  assign n2450 = n2449 ^ n2428 ;
  assign n2451 = ~n2430 & ~n2450 ;
  assign n2452 = n2451 ^ n2429 ;
  assign n2425 = n2370 & n2410 ;
  assign n2426 = n2425 ^ n2369 ;
  assign n2453 = n2452 ^ n2426 ;
  assign n2454 = n2368 ^ n2060 ;
  assign n2455 = n2454 ^ n2426 ;
  assign n2456 = ~n2453 & ~n2455 ;
  assign n2457 = n2456 ^ n2426 ;
  assign n2458 = n2457 ^ n2423 ;
  assign n2459 = ~n2424 & ~n2458 ;
  assign n2460 = n2459 ^ n2162 ;
  assign n2461 = n2422 & n2460 ;
  assign n2462 = n2461 ^ n2422 ;
  assign n2463 = n2462 ^ n2421 ;
  assign n2464 = x225 ^ x193 ;
  assign n2465 = n1533 & n2464 ;
  assign n2467 = n2465 ^ n2464 ;
  assign n2468 = n2467 ^ x193 ;
  assign n2469 = n2468 ^ x161 ;
  assign n2470 = n1574 & n2469 ;
  assign n2471 = n2470 ^ n2469 ;
  assign n2472 = n2471 ^ x161 ;
  assign n2466 = n2465 ^ x193 ;
  assign n2473 = n2472 ^ n2466 ;
  assign n2474 = n1646 & n2473 ;
  assign n2480 = n2474 ^ n2473 ;
  assign n2481 = n2480 ^ n2472 ;
  assign n2476 = n2470 ^ x161 ;
  assign n2477 = n2476 ^ x129 ;
  assign n2478 = ~n1611 & n2477 ;
  assign n2479 = n2478 ^ x129 ;
  assign n2482 = n2481 ^ n2479 ;
  assign n2483 = ~n1689 & n2482 ;
  assign n2489 = n2483 ^ n2482 ;
  assign n2490 = n2489 ^ n2481 ;
  assign n2491 = n2490 ^ x97 ;
  assign n2492 = ~n1725 & n2491 ;
  assign n2493 = n2492 ^ x97 ;
  assign n2484 = n2483 ^ n2481 ;
  assign n2475 = n2474 ^ n2472 ;
  assign n2485 = n2484 ^ n2475 ;
  assign n2486 = ~n1763 & n2485 ;
  assign n2487 = n2486 ^ n2485 ;
  assign n2488 = n2487 ^ n2484 ;
  assign n2494 = n2493 ^ n2488 ;
  assign n2495 = ~n1810 & n2494 ;
  assign n2502 = n2495 ^ n2494 ;
  assign n2503 = n2502 ^ n2493 ;
  assign n2504 = n2503 ^ x65 ;
  assign n2505 = ~n1846 & n2504 ;
  assign n2506 = n2505 ^ x65 ;
  assign n2497 = n2486 ^ n2484 ;
  assign n2496 = n2495 ^ n2493 ;
  assign n2498 = n2497 ^ n2496 ;
  assign n2499 = ~n1885 & n2498 ;
  assign n2500 = n2499 ^ n2498 ;
  assign n2501 = n2500 ^ n2497 ;
  assign n2507 = n2506 ^ n2501 ;
  assign n2508 = ~n1932 & n2507 ;
  assign n2515 = n2508 ^ n2507 ;
  assign n2516 = n2515 ^ n2506 ;
  assign n2517 = n2516 ^ x33 ;
  assign n2518 = ~n1968 & n2517 ;
  assign n2519 = n2518 ^ x33 ;
  assign n2510 = n2499 ^ n2497 ;
  assign n2509 = n2508 ^ n2506 ;
  assign n2511 = n2510 ^ n2509 ;
  assign n2512 = ~n2006 & n2511 ;
  assign n2513 = n2512 ^ n2511 ;
  assign n2514 = n2513 ^ n2510 ;
  assign n2520 = n2519 ^ n2514 ;
  assign n2521 = n2054 & n2520 ;
  assign n2527 = n2521 ^ n2520 ;
  assign n2528 = n2527 ^ n2519 ;
  assign n2526 = n2512 ^ n2510 ;
  assign n2529 = n2528 ^ n2526 ;
  assign n2530 = n2097 & n2529 ;
  assign n2536 = n2530 ^ n2529 ;
  assign n2537 = n2536 ^ n2528 ;
  assign n2531 = n2530 ^ n2528 ;
  assign n2522 = n2521 ^ n2519 ;
  assign n2523 = n2522 ^ x1 ;
  assign n2524 = ~n2365 & n2523 ;
  assign n2525 = n2524 ^ x1 ;
  assign n2532 = n2531 ^ n2525 ;
  assign n2533 = ~n2410 & n2532 ;
  assign n2534 = n2533 ^ n2532 ;
  assign n2535 = n2534 ^ n2531 ;
  assign n2538 = n2537 ^ n2535 ;
  assign n2539 = ~n2460 & n2538 ;
  assign n2540 = n2539 ^ n2538 ;
  assign n2541 = n2540 ^ n2537 ;
  assign n2542 = x226 ^ x194 ;
  assign n2543 = n1533 & n2542 ;
  assign n2545 = n2543 ^ n2542 ;
  assign n2546 = n2545 ^ x194 ;
  assign n2547 = n2546 ^ x162 ;
  assign n2548 = n1574 & n2547 ;
  assign n2549 = n2548 ^ n2547 ;
  assign n2550 = n2549 ^ x162 ;
  assign n2544 = n2543 ^ x194 ;
  assign n2551 = n2550 ^ n2544 ;
  assign n2552 = n1646 & n2551 ;
  assign n2558 = n2552 ^ n2551 ;
  assign n2559 = n2558 ^ n2550 ;
  assign n2554 = n2548 ^ x162 ;
  assign n2555 = n2554 ^ x130 ;
  assign n2556 = ~n1611 & n2555 ;
  assign n2557 = n2556 ^ x130 ;
  assign n2560 = n2559 ^ n2557 ;
  assign n2561 = ~n1689 & n2560 ;
  assign n2567 = n2561 ^ n2560 ;
  assign n2568 = n2567 ^ n2559 ;
  assign n2569 = n2568 ^ x98 ;
  assign n2570 = ~n1725 & n2569 ;
  assign n2571 = n2570 ^ x98 ;
  assign n2562 = n2561 ^ n2559 ;
  assign n2553 = n2552 ^ n2550 ;
  assign n2563 = n2562 ^ n2553 ;
  assign n2564 = ~n1763 & n2563 ;
  assign n2565 = n2564 ^ n2563 ;
  assign n2566 = n2565 ^ n2562 ;
  assign n2572 = n2571 ^ n2566 ;
  assign n2573 = ~n1810 & n2572 ;
  assign n2580 = n2573 ^ n2572 ;
  assign n2581 = n2580 ^ n2571 ;
  assign n2582 = n2581 ^ x66 ;
  assign n2583 = ~n1846 & n2582 ;
  assign n2584 = n2583 ^ x66 ;
  assign n2575 = n2564 ^ n2562 ;
  assign n2574 = n2573 ^ n2571 ;
  assign n2576 = n2575 ^ n2574 ;
  assign n2577 = ~n1885 & n2576 ;
  assign n2578 = n2577 ^ n2576 ;
  assign n2579 = n2578 ^ n2575 ;
  assign n2585 = n2584 ^ n2579 ;
  assign n2586 = ~n1932 & n2585 ;
  assign n2593 = n2586 ^ n2585 ;
  assign n2594 = n2593 ^ n2584 ;
  assign n2595 = n2594 ^ x34 ;
  assign n2596 = ~n1968 & n2595 ;
  assign n2597 = n2596 ^ x34 ;
  assign n2588 = n2577 ^ n2575 ;
  assign n2587 = n2586 ^ n2584 ;
  assign n2589 = n2588 ^ n2587 ;
  assign n2590 = ~n2006 & n2589 ;
  assign n2591 = n2590 ^ n2589 ;
  assign n2592 = n2591 ^ n2588 ;
  assign n2598 = n2597 ^ n2592 ;
  assign n2599 = n2054 & n2598 ;
  assign n2605 = n2599 ^ n2598 ;
  assign n2606 = n2605 ^ n2597 ;
  assign n2604 = n2590 ^ n2588 ;
  assign n2607 = n2606 ^ n2604 ;
  assign n2608 = n2097 & n2607 ;
  assign n2614 = n2608 ^ n2607 ;
  assign n2615 = n2614 ^ n2606 ;
  assign n2609 = n2608 ^ n2606 ;
  assign n2600 = n2599 ^ n2597 ;
  assign n2601 = n2600 ^ x2 ;
  assign n2602 = ~n2365 & n2601 ;
  assign n2603 = n2602 ^ x2 ;
  assign n2610 = n2609 ^ n2603 ;
  assign n2611 = ~n2410 & n2610 ;
  assign n2612 = n2611 ^ n2610 ;
  assign n2613 = n2612 ^ n2609 ;
  assign n2616 = n2615 ^ n2613 ;
  assign n2617 = ~n2460 & n2616 ;
  assign n2618 = n2617 ^ n2616 ;
  assign n2619 = n2618 ^ n2615 ;
  assign n2620 = x227 ^ x195 ;
  assign n2621 = n1533 & n2620 ;
  assign n2623 = n2621 ^ n2620 ;
  assign n2624 = n2623 ^ x195 ;
  assign n2625 = n2624 ^ x163 ;
  assign n2626 = n1574 & n2625 ;
  assign n2627 = n2626 ^ n2625 ;
  assign n2628 = n2627 ^ x163 ;
  assign n2622 = n2621 ^ x195 ;
  assign n2629 = n2628 ^ n2622 ;
  assign n2630 = n1646 & n2629 ;
  assign n2636 = n2630 ^ n2629 ;
  assign n2637 = n2636 ^ n2628 ;
  assign n2632 = n2626 ^ x163 ;
  assign n2633 = n2632 ^ x131 ;
  assign n2634 = ~n1611 & n2633 ;
  assign n2635 = n2634 ^ x131 ;
  assign n2638 = n2637 ^ n2635 ;
  assign n2639 = ~n1689 & n2638 ;
  assign n2645 = n2639 ^ n2638 ;
  assign n2646 = n2645 ^ n2637 ;
  assign n2647 = n2646 ^ x99 ;
  assign n2648 = ~n1725 & n2647 ;
  assign n2649 = n2648 ^ x99 ;
  assign n2640 = n2639 ^ n2637 ;
  assign n2631 = n2630 ^ n2628 ;
  assign n2641 = n2640 ^ n2631 ;
  assign n2642 = ~n1763 & n2641 ;
  assign n2643 = n2642 ^ n2641 ;
  assign n2644 = n2643 ^ n2640 ;
  assign n2650 = n2649 ^ n2644 ;
  assign n2651 = ~n1810 & n2650 ;
  assign n2658 = n2651 ^ n2650 ;
  assign n2659 = n2658 ^ n2649 ;
  assign n2660 = n2659 ^ x67 ;
  assign n2661 = ~n1846 & n2660 ;
  assign n2662 = n2661 ^ x67 ;
  assign n2653 = n2642 ^ n2640 ;
  assign n2652 = n2651 ^ n2649 ;
  assign n2654 = n2653 ^ n2652 ;
  assign n2655 = ~n1885 & n2654 ;
  assign n2656 = n2655 ^ n2654 ;
  assign n2657 = n2656 ^ n2653 ;
  assign n2663 = n2662 ^ n2657 ;
  assign n2664 = ~n1932 & n2663 ;
  assign n2671 = n2664 ^ n2663 ;
  assign n2672 = n2671 ^ n2662 ;
  assign n2673 = n2672 ^ x35 ;
  assign n2674 = ~n1968 & n2673 ;
  assign n2675 = n2674 ^ x35 ;
  assign n2666 = n2655 ^ n2653 ;
  assign n2665 = n2664 ^ n2662 ;
  assign n2667 = n2666 ^ n2665 ;
  assign n2668 = ~n2006 & n2667 ;
  assign n2669 = n2668 ^ n2667 ;
  assign n2670 = n2669 ^ n2666 ;
  assign n2676 = n2675 ^ n2670 ;
  assign n2677 = n2054 & n2676 ;
  assign n2683 = n2677 ^ n2676 ;
  assign n2684 = n2683 ^ n2675 ;
  assign n2682 = n2668 ^ n2666 ;
  assign n2685 = n2684 ^ n2682 ;
  assign n2686 = n2097 & n2685 ;
  assign n2692 = n2686 ^ n2685 ;
  assign n2693 = n2692 ^ n2684 ;
  assign n2687 = n2686 ^ n2684 ;
  assign n2678 = n2677 ^ n2675 ;
  assign n2679 = n2678 ^ x3 ;
  assign n2680 = ~n2365 & n2679 ;
  assign n2681 = n2680 ^ x3 ;
  assign n2688 = n2687 ^ n2681 ;
  assign n2689 = ~n2410 & n2688 ;
  assign n2690 = n2689 ^ n2688 ;
  assign n2691 = n2690 ^ n2687 ;
  assign n2694 = n2693 ^ n2691 ;
  assign n2695 = ~n2460 & n2694 ;
  assign n2696 = n2695 ^ n2694 ;
  assign n2697 = n2696 ^ n2693 ;
  assign n2698 = x228 ^ x196 ;
  assign n2699 = n1533 & n2698 ;
  assign n2701 = n2699 ^ n2698 ;
  assign n2702 = n2701 ^ x196 ;
  assign n2703 = n2702 ^ x164 ;
  assign n2704 = n1574 & n2703 ;
  assign n2705 = n2704 ^ n2703 ;
  assign n2706 = n2705 ^ x164 ;
  assign n2700 = n2699 ^ x196 ;
  assign n2707 = n2706 ^ n2700 ;
  assign n2708 = n1646 & n2707 ;
  assign n2714 = n2708 ^ n2707 ;
  assign n2715 = n2714 ^ n2706 ;
  assign n2710 = n2704 ^ x164 ;
  assign n2711 = n2710 ^ x132 ;
  assign n2712 = ~n1611 & n2711 ;
  assign n2713 = n2712 ^ x132 ;
  assign n2716 = n2715 ^ n2713 ;
  assign n2717 = ~n1689 & n2716 ;
  assign n2723 = n2717 ^ n2716 ;
  assign n2724 = n2723 ^ n2715 ;
  assign n2725 = n2724 ^ x100 ;
  assign n2726 = ~n1725 & n2725 ;
  assign n2727 = n2726 ^ x100 ;
  assign n2718 = n2717 ^ n2715 ;
  assign n2709 = n2708 ^ n2706 ;
  assign n2719 = n2718 ^ n2709 ;
  assign n2720 = ~n1763 & n2719 ;
  assign n2721 = n2720 ^ n2719 ;
  assign n2722 = n2721 ^ n2718 ;
  assign n2728 = n2727 ^ n2722 ;
  assign n2729 = ~n1810 & n2728 ;
  assign n2736 = n2729 ^ n2728 ;
  assign n2737 = n2736 ^ n2727 ;
  assign n2738 = n2737 ^ x68 ;
  assign n2739 = ~n1846 & n2738 ;
  assign n2740 = n2739 ^ x68 ;
  assign n2731 = n2720 ^ n2718 ;
  assign n2730 = n2729 ^ n2727 ;
  assign n2732 = n2731 ^ n2730 ;
  assign n2733 = ~n1885 & n2732 ;
  assign n2734 = n2733 ^ n2732 ;
  assign n2735 = n2734 ^ n2731 ;
  assign n2741 = n2740 ^ n2735 ;
  assign n2742 = ~n1932 & n2741 ;
  assign n2749 = n2742 ^ n2741 ;
  assign n2750 = n2749 ^ n2740 ;
  assign n2751 = n2750 ^ x36 ;
  assign n2752 = ~n1968 & n2751 ;
  assign n2753 = n2752 ^ x36 ;
  assign n2744 = n2733 ^ n2731 ;
  assign n2743 = n2742 ^ n2740 ;
  assign n2745 = n2744 ^ n2743 ;
  assign n2746 = ~n2006 & n2745 ;
  assign n2747 = n2746 ^ n2745 ;
  assign n2748 = n2747 ^ n2744 ;
  assign n2754 = n2753 ^ n2748 ;
  assign n2755 = n2054 & n2754 ;
  assign n2761 = n2755 ^ n2754 ;
  assign n2762 = n2761 ^ n2753 ;
  assign n2760 = n2746 ^ n2744 ;
  assign n2763 = n2762 ^ n2760 ;
  assign n2764 = n2097 & n2763 ;
  assign n2770 = n2764 ^ n2763 ;
  assign n2771 = n2770 ^ n2762 ;
  assign n2765 = n2764 ^ n2762 ;
  assign n2756 = n2755 ^ n2753 ;
  assign n2757 = n2756 ^ x4 ;
  assign n2758 = ~n2365 & n2757 ;
  assign n2759 = n2758 ^ x4 ;
  assign n2766 = n2765 ^ n2759 ;
  assign n2767 = ~n2410 & n2766 ;
  assign n2768 = n2767 ^ n2766 ;
  assign n2769 = n2768 ^ n2765 ;
  assign n2772 = n2771 ^ n2769 ;
  assign n2773 = ~n2460 & n2772 ;
  assign n2774 = n2773 ^ n2772 ;
  assign n2775 = n2774 ^ n2771 ;
  assign n2776 = x229 ^ x197 ;
  assign n2777 = n1533 & n2776 ;
  assign n2779 = n2777 ^ n2776 ;
  assign n2780 = n2779 ^ x197 ;
  assign n2781 = n2780 ^ x165 ;
  assign n2782 = n1574 & n2781 ;
  assign n2783 = n2782 ^ n2781 ;
  assign n2784 = n2783 ^ x165 ;
  assign n2778 = n2777 ^ x197 ;
  assign n2785 = n2784 ^ n2778 ;
  assign n2786 = n1646 & n2785 ;
  assign n2792 = n2786 ^ n2785 ;
  assign n2793 = n2792 ^ n2784 ;
  assign n2788 = n2782 ^ x165 ;
  assign n2789 = n2788 ^ x133 ;
  assign n2790 = ~n1611 & n2789 ;
  assign n2791 = n2790 ^ x133 ;
  assign n2794 = n2793 ^ n2791 ;
  assign n2795 = ~n1689 & n2794 ;
  assign n2801 = n2795 ^ n2794 ;
  assign n2802 = n2801 ^ n2793 ;
  assign n2803 = n2802 ^ x101 ;
  assign n2804 = ~n1725 & n2803 ;
  assign n2805 = n2804 ^ x101 ;
  assign n2796 = n2795 ^ n2793 ;
  assign n2787 = n2786 ^ n2784 ;
  assign n2797 = n2796 ^ n2787 ;
  assign n2798 = ~n1763 & n2797 ;
  assign n2799 = n2798 ^ n2797 ;
  assign n2800 = n2799 ^ n2796 ;
  assign n2806 = n2805 ^ n2800 ;
  assign n2807 = ~n1810 & n2806 ;
  assign n2814 = n2807 ^ n2806 ;
  assign n2815 = n2814 ^ n2805 ;
  assign n2816 = n2815 ^ x69 ;
  assign n2817 = ~n1846 & n2816 ;
  assign n2818 = n2817 ^ x69 ;
  assign n2809 = n2798 ^ n2796 ;
  assign n2808 = n2807 ^ n2805 ;
  assign n2810 = n2809 ^ n2808 ;
  assign n2811 = ~n1885 & n2810 ;
  assign n2812 = n2811 ^ n2810 ;
  assign n2813 = n2812 ^ n2809 ;
  assign n2819 = n2818 ^ n2813 ;
  assign n2820 = ~n1932 & n2819 ;
  assign n2827 = n2820 ^ n2819 ;
  assign n2828 = n2827 ^ n2818 ;
  assign n2829 = n2828 ^ x37 ;
  assign n2830 = ~n1968 & n2829 ;
  assign n2831 = n2830 ^ x37 ;
  assign n2822 = n2811 ^ n2809 ;
  assign n2821 = n2820 ^ n2818 ;
  assign n2823 = n2822 ^ n2821 ;
  assign n2824 = ~n2006 & n2823 ;
  assign n2825 = n2824 ^ n2823 ;
  assign n2826 = n2825 ^ n2822 ;
  assign n2832 = n2831 ^ n2826 ;
  assign n2833 = n2054 & n2832 ;
  assign n2839 = n2833 ^ n2832 ;
  assign n2840 = n2839 ^ n2831 ;
  assign n2838 = n2824 ^ n2822 ;
  assign n2841 = n2840 ^ n2838 ;
  assign n2842 = n2097 & n2841 ;
  assign n2848 = n2842 ^ n2841 ;
  assign n2849 = n2848 ^ n2840 ;
  assign n2843 = n2842 ^ n2840 ;
  assign n2834 = n2833 ^ n2831 ;
  assign n2835 = n2834 ^ x5 ;
  assign n2836 = ~n2365 & n2835 ;
  assign n2837 = n2836 ^ x5 ;
  assign n2844 = n2843 ^ n2837 ;
  assign n2845 = ~n2410 & n2844 ;
  assign n2846 = n2845 ^ n2844 ;
  assign n2847 = n2846 ^ n2843 ;
  assign n2850 = n2849 ^ n2847 ;
  assign n2851 = ~n2460 & n2850 ;
  assign n2852 = n2851 ^ n2850 ;
  assign n2853 = n2852 ^ n2849 ;
  assign n2854 = x230 ^ x198 ;
  assign n2855 = n1533 & n2854 ;
  assign n2857 = n2855 ^ n2854 ;
  assign n2858 = n2857 ^ x198 ;
  assign n2859 = n2858 ^ x166 ;
  assign n2860 = n1574 & n2859 ;
  assign n2861 = n2860 ^ n2859 ;
  assign n2862 = n2861 ^ x166 ;
  assign n2856 = n2855 ^ x198 ;
  assign n2863 = n2862 ^ n2856 ;
  assign n2864 = n1646 & n2863 ;
  assign n2870 = n2864 ^ n2863 ;
  assign n2871 = n2870 ^ n2862 ;
  assign n2866 = n2860 ^ x166 ;
  assign n2867 = n2866 ^ x134 ;
  assign n2868 = ~n1611 & n2867 ;
  assign n2869 = n2868 ^ x134 ;
  assign n2872 = n2871 ^ n2869 ;
  assign n2873 = ~n1689 & n2872 ;
  assign n2879 = n2873 ^ n2872 ;
  assign n2880 = n2879 ^ n2871 ;
  assign n2881 = n2880 ^ x102 ;
  assign n2882 = ~n1725 & n2881 ;
  assign n2883 = n2882 ^ x102 ;
  assign n2874 = n2873 ^ n2871 ;
  assign n2865 = n2864 ^ n2862 ;
  assign n2875 = n2874 ^ n2865 ;
  assign n2876 = ~n1763 & n2875 ;
  assign n2877 = n2876 ^ n2875 ;
  assign n2878 = n2877 ^ n2874 ;
  assign n2884 = n2883 ^ n2878 ;
  assign n2885 = ~n1810 & n2884 ;
  assign n2892 = n2885 ^ n2884 ;
  assign n2893 = n2892 ^ n2883 ;
  assign n2894 = n2893 ^ x70 ;
  assign n2895 = ~n1846 & n2894 ;
  assign n2896 = n2895 ^ x70 ;
  assign n2887 = n2876 ^ n2874 ;
  assign n2886 = n2885 ^ n2883 ;
  assign n2888 = n2887 ^ n2886 ;
  assign n2889 = ~n1885 & n2888 ;
  assign n2890 = n2889 ^ n2888 ;
  assign n2891 = n2890 ^ n2887 ;
  assign n2897 = n2896 ^ n2891 ;
  assign n2898 = ~n1932 & n2897 ;
  assign n2905 = n2898 ^ n2897 ;
  assign n2906 = n2905 ^ n2896 ;
  assign n2907 = n2906 ^ x38 ;
  assign n2908 = ~n1968 & n2907 ;
  assign n2909 = n2908 ^ x38 ;
  assign n2900 = n2889 ^ n2887 ;
  assign n2899 = n2898 ^ n2896 ;
  assign n2901 = n2900 ^ n2899 ;
  assign n2902 = ~n2006 & n2901 ;
  assign n2903 = n2902 ^ n2901 ;
  assign n2904 = n2903 ^ n2900 ;
  assign n2910 = n2909 ^ n2904 ;
  assign n2911 = n2054 & n2910 ;
  assign n2917 = n2911 ^ n2910 ;
  assign n2918 = n2917 ^ n2909 ;
  assign n2916 = n2902 ^ n2900 ;
  assign n2919 = n2918 ^ n2916 ;
  assign n2920 = n2097 & n2919 ;
  assign n2926 = n2920 ^ n2919 ;
  assign n2927 = n2926 ^ n2918 ;
  assign n2921 = n2920 ^ n2918 ;
  assign n2912 = n2911 ^ n2909 ;
  assign n2913 = n2912 ^ x6 ;
  assign n2914 = ~n2365 & n2913 ;
  assign n2915 = n2914 ^ x6 ;
  assign n2922 = n2921 ^ n2915 ;
  assign n2923 = ~n2410 & n2922 ;
  assign n2924 = n2923 ^ n2922 ;
  assign n2925 = n2924 ^ n2921 ;
  assign n2928 = n2927 ^ n2925 ;
  assign n2929 = ~n2460 & n2928 ;
  assign n2930 = n2929 ^ n2928 ;
  assign n2931 = n2930 ^ n2927 ;
  assign n2932 = x231 ^ x199 ;
  assign n2933 = n1533 & n2932 ;
  assign n2935 = n2933 ^ n2932 ;
  assign n2936 = n2935 ^ x199 ;
  assign n2937 = n2936 ^ x167 ;
  assign n2938 = n1574 & n2937 ;
  assign n2939 = n2938 ^ n2937 ;
  assign n2940 = n2939 ^ x167 ;
  assign n2934 = n2933 ^ x199 ;
  assign n2941 = n2940 ^ n2934 ;
  assign n2942 = n1646 & n2941 ;
  assign n2948 = n2942 ^ n2941 ;
  assign n2949 = n2948 ^ n2940 ;
  assign n2944 = n2938 ^ x167 ;
  assign n2945 = n2944 ^ x135 ;
  assign n2946 = ~n1611 & n2945 ;
  assign n2947 = n2946 ^ x135 ;
  assign n2950 = n2949 ^ n2947 ;
  assign n2951 = ~n1689 & n2950 ;
  assign n2957 = n2951 ^ n2950 ;
  assign n2958 = n2957 ^ n2949 ;
  assign n2959 = n2958 ^ x103 ;
  assign n2960 = ~n1725 & n2959 ;
  assign n2961 = n2960 ^ x103 ;
  assign n2952 = n2951 ^ n2949 ;
  assign n2943 = n2942 ^ n2940 ;
  assign n2953 = n2952 ^ n2943 ;
  assign n2954 = ~n1763 & n2953 ;
  assign n2955 = n2954 ^ n2953 ;
  assign n2956 = n2955 ^ n2952 ;
  assign n2962 = n2961 ^ n2956 ;
  assign n2963 = ~n1810 & n2962 ;
  assign n2970 = n2963 ^ n2962 ;
  assign n2971 = n2970 ^ n2961 ;
  assign n2972 = n2971 ^ x71 ;
  assign n2973 = ~n1846 & n2972 ;
  assign n2974 = n2973 ^ x71 ;
  assign n2965 = n2954 ^ n2952 ;
  assign n2964 = n2963 ^ n2961 ;
  assign n2966 = n2965 ^ n2964 ;
  assign n2967 = ~n1885 & n2966 ;
  assign n2968 = n2967 ^ n2966 ;
  assign n2969 = n2968 ^ n2965 ;
  assign n2975 = n2974 ^ n2969 ;
  assign n2976 = ~n1932 & n2975 ;
  assign n2983 = n2976 ^ n2975 ;
  assign n2984 = n2983 ^ n2974 ;
  assign n2985 = n2984 ^ x39 ;
  assign n2986 = ~n1968 & n2985 ;
  assign n2987 = n2986 ^ x39 ;
  assign n2978 = n2967 ^ n2965 ;
  assign n2977 = n2976 ^ n2974 ;
  assign n2979 = n2978 ^ n2977 ;
  assign n2980 = ~n2006 & n2979 ;
  assign n2981 = n2980 ^ n2979 ;
  assign n2982 = n2981 ^ n2978 ;
  assign n2988 = n2987 ^ n2982 ;
  assign n2989 = n2054 & n2988 ;
  assign n2995 = n2989 ^ n2988 ;
  assign n2996 = n2995 ^ n2987 ;
  assign n2994 = n2980 ^ n2978 ;
  assign n2997 = n2996 ^ n2994 ;
  assign n2998 = n2097 & n2997 ;
  assign n3004 = n2998 ^ n2997 ;
  assign n3005 = n3004 ^ n2996 ;
  assign n2999 = n2998 ^ n2996 ;
  assign n2990 = n2989 ^ n2987 ;
  assign n2991 = n2990 ^ x7 ;
  assign n2992 = ~n2365 & n2991 ;
  assign n2993 = n2992 ^ x7 ;
  assign n3000 = n2999 ^ n2993 ;
  assign n3001 = ~n2410 & n3000 ;
  assign n3002 = n3001 ^ n3000 ;
  assign n3003 = n3002 ^ n2999 ;
  assign n3006 = n3005 ^ n3003 ;
  assign n3007 = ~n2460 & n3006 ;
  assign n3008 = n3007 ^ n3006 ;
  assign n3009 = n3008 ^ n3005 ;
  assign n3010 = x232 ^ x200 ;
  assign n3011 = n1533 & n3010 ;
  assign n3013 = n3011 ^ n3010 ;
  assign n3014 = n3013 ^ x200 ;
  assign n3015 = n3014 ^ x168 ;
  assign n3016 = n1574 & n3015 ;
  assign n3017 = n3016 ^ n3015 ;
  assign n3018 = n3017 ^ x168 ;
  assign n3012 = n3011 ^ x200 ;
  assign n3019 = n3018 ^ n3012 ;
  assign n3020 = n1646 & n3019 ;
  assign n3026 = n3020 ^ n3019 ;
  assign n3027 = n3026 ^ n3018 ;
  assign n3022 = n3016 ^ x168 ;
  assign n3023 = n3022 ^ x136 ;
  assign n3024 = ~n1611 & n3023 ;
  assign n3025 = n3024 ^ x136 ;
  assign n3028 = n3027 ^ n3025 ;
  assign n3029 = ~n1689 & n3028 ;
  assign n3035 = n3029 ^ n3028 ;
  assign n3036 = n3035 ^ n3027 ;
  assign n3037 = n3036 ^ x104 ;
  assign n3038 = ~n1725 & n3037 ;
  assign n3039 = n3038 ^ x104 ;
  assign n3030 = n3029 ^ n3027 ;
  assign n3021 = n3020 ^ n3018 ;
  assign n3031 = n3030 ^ n3021 ;
  assign n3032 = ~n1763 & n3031 ;
  assign n3033 = n3032 ^ n3031 ;
  assign n3034 = n3033 ^ n3030 ;
  assign n3040 = n3039 ^ n3034 ;
  assign n3041 = ~n1810 & n3040 ;
  assign n3048 = n3041 ^ n3040 ;
  assign n3049 = n3048 ^ n3039 ;
  assign n3050 = n3049 ^ x72 ;
  assign n3051 = ~n1846 & n3050 ;
  assign n3052 = n3051 ^ x72 ;
  assign n3043 = n3032 ^ n3030 ;
  assign n3042 = n3041 ^ n3039 ;
  assign n3044 = n3043 ^ n3042 ;
  assign n3045 = ~n1885 & n3044 ;
  assign n3046 = n3045 ^ n3044 ;
  assign n3047 = n3046 ^ n3043 ;
  assign n3053 = n3052 ^ n3047 ;
  assign n3054 = ~n1932 & n3053 ;
  assign n3061 = n3054 ^ n3053 ;
  assign n3062 = n3061 ^ n3052 ;
  assign n3063 = n3062 ^ x40 ;
  assign n3064 = ~n1968 & n3063 ;
  assign n3065 = n3064 ^ x40 ;
  assign n3056 = n3045 ^ n3043 ;
  assign n3055 = n3054 ^ n3052 ;
  assign n3057 = n3056 ^ n3055 ;
  assign n3058 = ~n2006 & n3057 ;
  assign n3059 = n3058 ^ n3057 ;
  assign n3060 = n3059 ^ n3056 ;
  assign n3066 = n3065 ^ n3060 ;
  assign n3067 = n2054 & n3066 ;
  assign n3073 = n3067 ^ n3066 ;
  assign n3074 = n3073 ^ n3065 ;
  assign n3072 = n3058 ^ n3056 ;
  assign n3075 = n3074 ^ n3072 ;
  assign n3076 = n2097 & n3075 ;
  assign n3082 = n3076 ^ n3075 ;
  assign n3083 = n3082 ^ n3074 ;
  assign n3077 = n3076 ^ n3074 ;
  assign n3068 = n3067 ^ n3065 ;
  assign n3069 = n3068 ^ x8 ;
  assign n3070 = ~n2365 & n3069 ;
  assign n3071 = n3070 ^ x8 ;
  assign n3078 = n3077 ^ n3071 ;
  assign n3079 = ~n2410 & n3078 ;
  assign n3080 = n3079 ^ n3078 ;
  assign n3081 = n3080 ^ n3077 ;
  assign n3084 = n3083 ^ n3081 ;
  assign n3085 = ~n2460 & n3084 ;
  assign n3086 = n3085 ^ n3084 ;
  assign n3087 = n3086 ^ n3083 ;
  assign n3088 = x233 ^ x201 ;
  assign n3089 = n1533 & n3088 ;
  assign n3091 = n3089 ^ n3088 ;
  assign n3092 = n3091 ^ x201 ;
  assign n3093 = n3092 ^ x169 ;
  assign n3094 = n1574 & n3093 ;
  assign n3095 = n3094 ^ n3093 ;
  assign n3096 = n3095 ^ x169 ;
  assign n3090 = n3089 ^ x201 ;
  assign n3097 = n3096 ^ n3090 ;
  assign n3098 = n1646 & n3097 ;
  assign n3104 = n3098 ^ n3097 ;
  assign n3105 = n3104 ^ n3096 ;
  assign n3100 = n3094 ^ x169 ;
  assign n3101 = n3100 ^ x137 ;
  assign n3102 = ~n1611 & n3101 ;
  assign n3103 = n3102 ^ x137 ;
  assign n3106 = n3105 ^ n3103 ;
  assign n3107 = ~n1689 & n3106 ;
  assign n3113 = n3107 ^ n3106 ;
  assign n3114 = n3113 ^ n3105 ;
  assign n3115 = n3114 ^ x105 ;
  assign n3116 = ~n1725 & n3115 ;
  assign n3117 = n3116 ^ x105 ;
  assign n3108 = n3107 ^ n3105 ;
  assign n3099 = n3098 ^ n3096 ;
  assign n3109 = n3108 ^ n3099 ;
  assign n3110 = ~n1763 & n3109 ;
  assign n3111 = n3110 ^ n3109 ;
  assign n3112 = n3111 ^ n3108 ;
  assign n3118 = n3117 ^ n3112 ;
  assign n3119 = ~n1810 & n3118 ;
  assign n3126 = n3119 ^ n3118 ;
  assign n3127 = n3126 ^ n3117 ;
  assign n3128 = n3127 ^ x73 ;
  assign n3129 = ~n1846 & n3128 ;
  assign n3130 = n3129 ^ x73 ;
  assign n3121 = n3110 ^ n3108 ;
  assign n3120 = n3119 ^ n3117 ;
  assign n3122 = n3121 ^ n3120 ;
  assign n3123 = ~n1885 & n3122 ;
  assign n3124 = n3123 ^ n3122 ;
  assign n3125 = n3124 ^ n3121 ;
  assign n3131 = n3130 ^ n3125 ;
  assign n3132 = ~n1932 & n3131 ;
  assign n3139 = n3132 ^ n3131 ;
  assign n3140 = n3139 ^ n3130 ;
  assign n3141 = n3140 ^ x41 ;
  assign n3142 = ~n1968 & n3141 ;
  assign n3143 = n3142 ^ x41 ;
  assign n3134 = n3123 ^ n3121 ;
  assign n3133 = n3132 ^ n3130 ;
  assign n3135 = n3134 ^ n3133 ;
  assign n3136 = ~n2006 & n3135 ;
  assign n3137 = n3136 ^ n3135 ;
  assign n3138 = n3137 ^ n3134 ;
  assign n3144 = n3143 ^ n3138 ;
  assign n3145 = n2054 & n3144 ;
  assign n3151 = n3145 ^ n3144 ;
  assign n3152 = n3151 ^ n3143 ;
  assign n3150 = n3136 ^ n3134 ;
  assign n3153 = n3152 ^ n3150 ;
  assign n3154 = n2097 & n3153 ;
  assign n3160 = n3154 ^ n3153 ;
  assign n3161 = n3160 ^ n3152 ;
  assign n3155 = n3154 ^ n3152 ;
  assign n3146 = n3145 ^ n3143 ;
  assign n3147 = n3146 ^ x9 ;
  assign n3148 = ~n2365 & n3147 ;
  assign n3149 = n3148 ^ x9 ;
  assign n3156 = n3155 ^ n3149 ;
  assign n3157 = ~n2410 & n3156 ;
  assign n3158 = n3157 ^ n3156 ;
  assign n3159 = n3158 ^ n3155 ;
  assign n3162 = n3161 ^ n3159 ;
  assign n3163 = ~n2460 & n3162 ;
  assign n3164 = n3163 ^ n3162 ;
  assign n3165 = n3164 ^ n3161 ;
  assign n3166 = x234 ^ x202 ;
  assign n3167 = n1533 & n3166 ;
  assign n3169 = n3167 ^ n3166 ;
  assign n3170 = n3169 ^ x202 ;
  assign n3171 = n3170 ^ x170 ;
  assign n3172 = n1574 & n3171 ;
  assign n3173 = n3172 ^ n3171 ;
  assign n3174 = n3173 ^ x170 ;
  assign n3168 = n3167 ^ x202 ;
  assign n3175 = n3174 ^ n3168 ;
  assign n3176 = n1646 & n3175 ;
  assign n3182 = n3176 ^ n3175 ;
  assign n3183 = n3182 ^ n3174 ;
  assign n3178 = n3172 ^ x170 ;
  assign n3179 = n3178 ^ x138 ;
  assign n3180 = ~n1611 & n3179 ;
  assign n3181 = n3180 ^ x138 ;
  assign n3184 = n3183 ^ n3181 ;
  assign n3185 = ~n1689 & n3184 ;
  assign n3191 = n3185 ^ n3184 ;
  assign n3192 = n3191 ^ n3183 ;
  assign n3193 = n3192 ^ x106 ;
  assign n3194 = ~n1725 & n3193 ;
  assign n3195 = n3194 ^ x106 ;
  assign n3186 = n3185 ^ n3183 ;
  assign n3177 = n3176 ^ n3174 ;
  assign n3187 = n3186 ^ n3177 ;
  assign n3188 = ~n1763 & n3187 ;
  assign n3189 = n3188 ^ n3187 ;
  assign n3190 = n3189 ^ n3186 ;
  assign n3196 = n3195 ^ n3190 ;
  assign n3197 = ~n1810 & n3196 ;
  assign n3204 = n3197 ^ n3196 ;
  assign n3205 = n3204 ^ n3195 ;
  assign n3206 = n3205 ^ x74 ;
  assign n3207 = ~n1846 & n3206 ;
  assign n3208 = n3207 ^ x74 ;
  assign n3199 = n3188 ^ n3186 ;
  assign n3198 = n3197 ^ n3195 ;
  assign n3200 = n3199 ^ n3198 ;
  assign n3201 = ~n1885 & n3200 ;
  assign n3202 = n3201 ^ n3200 ;
  assign n3203 = n3202 ^ n3199 ;
  assign n3209 = n3208 ^ n3203 ;
  assign n3210 = ~n1932 & n3209 ;
  assign n3217 = n3210 ^ n3209 ;
  assign n3218 = n3217 ^ n3208 ;
  assign n3219 = n3218 ^ x42 ;
  assign n3220 = ~n1968 & n3219 ;
  assign n3221 = n3220 ^ x42 ;
  assign n3212 = n3201 ^ n3199 ;
  assign n3211 = n3210 ^ n3208 ;
  assign n3213 = n3212 ^ n3211 ;
  assign n3214 = ~n2006 & n3213 ;
  assign n3215 = n3214 ^ n3213 ;
  assign n3216 = n3215 ^ n3212 ;
  assign n3222 = n3221 ^ n3216 ;
  assign n3223 = n2054 & n3222 ;
  assign n3229 = n3223 ^ n3222 ;
  assign n3230 = n3229 ^ n3221 ;
  assign n3228 = n3214 ^ n3212 ;
  assign n3231 = n3230 ^ n3228 ;
  assign n3232 = n2097 & n3231 ;
  assign n3238 = n3232 ^ n3231 ;
  assign n3239 = n3238 ^ n3230 ;
  assign n3233 = n3232 ^ n3230 ;
  assign n3224 = n3223 ^ n3221 ;
  assign n3225 = n3224 ^ x10 ;
  assign n3226 = ~n2365 & n3225 ;
  assign n3227 = n3226 ^ x10 ;
  assign n3234 = n3233 ^ n3227 ;
  assign n3235 = ~n2410 & n3234 ;
  assign n3236 = n3235 ^ n3234 ;
  assign n3237 = n3236 ^ n3233 ;
  assign n3240 = n3239 ^ n3237 ;
  assign n3241 = ~n2460 & n3240 ;
  assign n3242 = n3241 ^ n3240 ;
  assign n3243 = n3242 ^ n3239 ;
  assign n3244 = x235 ^ x203 ;
  assign n3245 = n1533 & n3244 ;
  assign n3247 = n3245 ^ n3244 ;
  assign n3248 = n3247 ^ x203 ;
  assign n3249 = n3248 ^ x171 ;
  assign n3250 = n1574 & n3249 ;
  assign n3251 = n3250 ^ n3249 ;
  assign n3252 = n3251 ^ x171 ;
  assign n3246 = n3245 ^ x203 ;
  assign n3253 = n3252 ^ n3246 ;
  assign n3254 = n1646 & n3253 ;
  assign n3260 = n3254 ^ n3253 ;
  assign n3261 = n3260 ^ n3252 ;
  assign n3256 = n3250 ^ x171 ;
  assign n3257 = n3256 ^ x139 ;
  assign n3258 = ~n1611 & n3257 ;
  assign n3259 = n3258 ^ x139 ;
  assign n3262 = n3261 ^ n3259 ;
  assign n3263 = ~n1689 & n3262 ;
  assign n3269 = n3263 ^ n3262 ;
  assign n3270 = n3269 ^ n3261 ;
  assign n3271 = n3270 ^ x107 ;
  assign n3272 = ~n1725 & n3271 ;
  assign n3273 = n3272 ^ x107 ;
  assign n3264 = n3263 ^ n3261 ;
  assign n3255 = n3254 ^ n3252 ;
  assign n3265 = n3264 ^ n3255 ;
  assign n3266 = ~n1763 & n3265 ;
  assign n3267 = n3266 ^ n3265 ;
  assign n3268 = n3267 ^ n3264 ;
  assign n3274 = n3273 ^ n3268 ;
  assign n3275 = ~n1810 & n3274 ;
  assign n3282 = n3275 ^ n3274 ;
  assign n3283 = n3282 ^ n3273 ;
  assign n3284 = n3283 ^ x75 ;
  assign n3285 = ~n1846 & n3284 ;
  assign n3286 = n3285 ^ x75 ;
  assign n3277 = n3266 ^ n3264 ;
  assign n3276 = n3275 ^ n3273 ;
  assign n3278 = n3277 ^ n3276 ;
  assign n3279 = ~n1885 & n3278 ;
  assign n3280 = n3279 ^ n3278 ;
  assign n3281 = n3280 ^ n3277 ;
  assign n3287 = n3286 ^ n3281 ;
  assign n3288 = ~n1932 & n3287 ;
  assign n3295 = n3288 ^ n3287 ;
  assign n3296 = n3295 ^ n3286 ;
  assign n3297 = n3296 ^ x43 ;
  assign n3298 = ~n1968 & n3297 ;
  assign n3299 = n3298 ^ x43 ;
  assign n3290 = n3279 ^ n3277 ;
  assign n3289 = n3288 ^ n3286 ;
  assign n3291 = n3290 ^ n3289 ;
  assign n3292 = ~n2006 & n3291 ;
  assign n3293 = n3292 ^ n3291 ;
  assign n3294 = n3293 ^ n3290 ;
  assign n3300 = n3299 ^ n3294 ;
  assign n3301 = n2054 & n3300 ;
  assign n3307 = n3301 ^ n3300 ;
  assign n3308 = n3307 ^ n3299 ;
  assign n3306 = n3292 ^ n3290 ;
  assign n3309 = n3308 ^ n3306 ;
  assign n3310 = n2097 & n3309 ;
  assign n3316 = n3310 ^ n3309 ;
  assign n3317 = n3316 ^ n3308 ;
  assign n3311 = n3310 ^ n3308 ;
  assign n3302 = n3301 ^ n3299 ;
  assign n3303 = n3302 ^ x11 ;
  assign n3304 = ~n2365 & n3303 ;
  assign n3305 = n3304 ^ x11 ;
  assign n3312 = n3311 ^ n3305 ;
  assign n3313 = ~n2410 & n3312 ;
  assign n3314 = n3313 ^ n3312 ;
  assign n3315 = n3314 ^ n3311 ;
  assign n3318 = n3317 ^ n3315 ;
  assign n3319 = ~n2460 & n3318 ;
  assign n3320 = n3319 ^ n3318 ;
  assign n3321 = n3320 ^ n3317 ;
  assign n3322 = x236 ^ x204 ;
  assign n3323 = n1533 & n3322 ;
  assign n3325 = n3323 ^ n3322 ;
  assign n3326 = n3325 ^ x204 ;
  assign n3327 = n3326 ^ x172 ;
  assign n3328 = n1574 & n3327 ;
  assign n3329 = n3328 ^ n3327 ;
  assign n3330 = n3329 ^ x172 ;
  assign n3324 = n3323 ^ x204 ;
  assign n3331 = n3330 ^ n3324 ;
  assign n3332 = n1646 & n3331 ;
  assign n3338 = n3332 ^ n3331 ;
  assign n3339 = n3338 ^ n3330 ;
  assign n3334 = n3328 ^ x172 ;
  assign n3335 = n3334 ^ x140 ;
  assign n3336 = ~n1611 & n3335 ;
  assign n3337 = n3336 ^ x140 ;
  assign n3340 = n3339 ^ n3337 ;
  assign n3341 = ~n1689 & n3340 ;
  assign n3347 = n3341 ^ n3340 ;
  assign n3348 = n3347 ^ n3339 ;
  assign n3349 = n3348 ^ x108 ;
  assign n3350 = ~n1725 & n3349 ;
  assign n3351 = n3350 ^ x108 ;
  assign n3342 = n3341 ^ n3339 ;
  assign n3333 = n3332 ^ n3330 ;
  assign n3343 = n3342 ^ n3333 ;
  assign n3344 = ~n1763 & n3343 ;
  assign n3345 = n3344 ^ n3343 ;
  assign n3346 = n3345 ^ n3342 ;
  assign n3352 = n3351 ^ n3346 ;
  assign n3353 = ~n1810 & n3352 ;
  assign n3360 = n3353 ^ n3352 ;
  assign n3361 = n3360 ^ n3351 ;
  assign n3362 = n3361 ^ x76 ;
  assign n3363 = ~n1846 & n3362 ;
  assign n3364 = n3363 ^ x76 ;
  assign n3355 = n3344 ^ n3342 ;
  assign n3354 = n3353 ^ n3351 ;
  assign n3356 = n3355 ^ n3354 ;
  assign n3357 = ~n1885 & n3356 ;
  assign n3358 = n3357 ^ n3356 ;
  assign n3359 = n3358 ^ n3355 ;
  assign n3365 = n3364 ^ n3359 ;
  assign n3366 = ~n1932 & n3365 ;
  assign n3373 = n3366 ^ n3365 ;
  assign n3374 = n3373 ^ n3364 ;
  assign n3375 = n3374 ^ x44 ;
  assign n3376 = ~n1968 & n3375 ;
  assign n3377 = n3376 ^ x44 ;
  assign n3368 = n3357 ^ n3355 ;
  assign n3367 = n3366 ^ n3364 ;
  assign n3369 = n3368 ^ n3367 ;
  assign n3370 = ~n2006 & n3369 ;
  assign n3371 = n3370 ^ n3369 ;
  assign n3372 = n3371 ^ n3368 ;
  assign n3378 = n3377 ^ n3372 ;
  assign n3379 = n2054 & n3378 ;
  assign n3385 = n3379 ^ n3378 ;
  assign n3386 = n3385 ^ n3377 ;
  assign n3384 = n3370 ^ n3368 ;
  assign n3387 = n3386 ^ n3384 ;
  assign n3388 = n2097 & n3387 ;
  assign n3394 = n3388 ^ n3387 ;
  assign n3395 = n3394 ^ n3386 ;
  assign n3389 = n3388 ^ n3386 ;
  assign n3380 = n3379 ^ n3377 ;
  assign n3381 = n3380 ^ x12 ;
  assign n3382 = ~n2365 & n3381 ;
  assign n3383 = n3382 ^ x12 ;
  assign n3390 = n3389 ^ n3383 ;
  assign n3391 = ~n2410 & n3390 ;
  assign n3392 = n3391 ^ n3390 ;
  assign n3393 = n3392 ^ n3389 ;
  assign n3396 = n3395 ^ n3393 ;
  assign n3397 = ~n2460 & n3396 ;
  assign n3398 = n3397 ^ n3396 ;
  assign n3399 = n3398 ^ n3395 ;
  assign n3400 = x237 ^ x205 ;
  assign n3401 = n1533 & n3400 ;
  assign n3403 = n3401 ^ n3400 ;
  assign n3404 = n3403 ^ x205 ;
  assign n3405 = n3404 ^ x173 ;
  assign n3406 = n1574 & n3405 ;
  assign n3407 = n3406 ^ n3405 ;
  assign n3408 = n3407 ^ x173 ;
  assign n3402 = n3401 ^ x205 ;
  assign n3409 = n3408 ^ n3402 ;
  assign n3410 = n1646 & n3409 ;
  assign n3416 = n3410 ^ n3409 ;
  assign n3417 = n3416 ^ n3408 ;
  assign n3412 = n3406 ^ x173 ;
  assign n3413 = n3412 ^ x141 ;
  assign n3414 = ~n1611 & n3413 ;
  assign n3415 = n3414 ^ x141 ;
  assign n3418 = n3417 ^ n3415 ;
  assign n3419 = ~n1689 & n3418 ;
  assign n3425 = n3419 ^ n3418 ;
  assign n3426 = n3425 ^ n3417 ;
  assign n3427 = n3426 ^ x109 ;
  assign n3428 = ~n1725 & n3427 ;
  assign n3429 = n3428 ^ x109 ;
  assign n3420 = n3419 ^ n3417 ;
  assign n3411 = n3410 ^ n3408 ;
  assign n3421 = n3420 ^ n3411 ;
  assign n3422 = ~n1763 & n3421 ;
  assign n3423 = n3422 ^ n3421 ;
  assign n3424 = n3423 ^ n3420 ;
  assign n3430 = n3429 ^ n3424 ;
  assign n3431 = ~n1810 & n3430 ;
  assign n3438 = n3431 ^ n3430 ;
  assign n3439 = n3438 ^ n3429 ;
  assign n3440 = n3439 ^ x77 ;
  assign n3441 = ~n1846 & n3440 ;
  assign n3442 = n3441 ^ x77 ;
  assign n3433 = n3422 ^ n3420 ;
  assign n3432 = n3431 ^ n3429 ;
  assign n3434 = n3433 ^ n3432 ;
  assign n3435 = ~n1885 & n3434 ;
  assign n3436 = n3435 ^ n3434 ;
  assign n3437 = n3436 ^ n3433 ;
  assign n3443 = n3442 ^ n3437 ;
  assign n3444 = ~n1932 & n3443 ;
  assign n3451 = n3444 ^ n3443 ;
  assign n3452 = n3451 ^ n3442 ;
  assign n3453 = n3452 ^ x45 ;
  assign n3454 = ~n1968 & n3453 ;
  assign n3455 = n3454 ^ x45 ;
  assign n3446 = n3435 ^ n3433 ;
  assign n3445 = n3444 ^ n3442 ;
  assign n3447 = n3446 ^ n3445 ;
  assign n3448 = ~n2006 & n3447 ;
  assign n3449 = n3448 ^ n3447 ;
  assign n3450 = n3449 ^ n3446 ;
  assign n3456 = n3455 ^ n3450 ;
  assign n3457 = n2054 & n3456 ;
  assign n3463 = n3457 ^ n3456 ;
  assign n3464 = n3463 ^ n3455 ;
  assign n3462 = n3448 ^ n3446 ;
  assign n3465 = n3464 ^ n3462 ;
  assign n3466 = n2097 & n3465 ;
  assign n3472 = n3466 ^ n3465 ;
  assign n3473 = n3472 ^ n3464 ;
  assign n3467 = n3466 ^ n3464 ;
  assign n3458 = n3457 ^ n3455 ;
  assign n3459 = n3458 ^ x13 ;
  assign n3460 = ~n2365 & n3459 ;
  assign n3461 = n3460 ^ x13 ;
  assign n3468 = n3467 ^ n3461 ;
  assign n3469 = ~n2410 & n3468 ;
  assign n3470 = n3469 ^ n3468 ;
  assign n3471 = n3470 ^ n3467 ;
  assign n3474 = n3473 ^ n3471 ;
  assign n3475 = ~n2460 & n3474 ;
  assign n3476 = n3475 ^ n3474 ;
  assign n3477 = n3476 ^ n3473 ;
  assign n3478 = x238 ^ x206 ;
  assign n3479 = n1533 & n3478 ;
  assign n3481 = n3479 ^ n3478 ;
  assign n3482 = n3481 ^ x206 ;
  assign n3483 = n3482 ^ x174 ;
  assign n3484 = n1574 & n3483 ;
  assign n3485 = n3484 ^ n3483 ;
  assign n3486 = n3485 ^ x174 ;
  assign n3480 = n3479 ^ x206 ;
  assign n3487 = n3486 ^ n3480 ;
  assign n3488 = n1646 & n3487 ;
  assign n3494 = n3488 ^ n3487 ;
  assign n3495 = n3494 ^ n3486 ;
  assign n3490 = n3484 ^ x174 ;
  assign n3491 = n3490 ^ x142 ;
  assign n3492 = ~n1611 & n3491 ;
  assign n3493 = n3492 ^ x142 ;
  assign n3496 = n3495 ^ n3493 ;
  assign n3497 = ~n1689 & n3496 ;
  assign n3503 = n3497 ^ n3496 ;
  assign n3504 = n3503 ^ n3495 ;
  assign n3505 = n3504 ^ x110 ;
  assign n3506 = ~n1725 & n3505 ;
  assign n3507 = n3506 ^ x110 ;
  assign n3498 = n3497 ^ n3495 ;
  assign n3489 = n3488 ^ n3486 ;
  assign n3499 = n3498 ^ n3489 ;
  assign n3500 = ~n1763 & n3499 ;
  assign n3501 = n3500 ^ n3499 ;
  assign n3502 = n3501 ^ n3498 ;
  assign n3508 = n3507 ^ n3502 ;
  assign n3509 = ~n1810 & n3508 ;
  assign n3516 = n3509 ^ n3508 ;
  assign n3517 = n3516 ^ n3507 ;
  assign n3518 = n3517 ^ x78 ;
  assign n3519 = ~n1846 & n3518 ;
  assign n3520 = n3519 ^ x78 ;
  assign n3511 = n3500 ^ n3498 ;
  assign n3510 = n3509 ^ n3507 ;
  assign n3512 = n3511 ^ n3510 ;
  assign n3513 = ~n1885 & n3512 ;
  assign n3514 = n3513 ^ n3512 ;
  assign n3515 = n3514 ^ n3511 ;
  assign n3521 = n3520 ^ n3515 ;
  assign n3522 = ~n1932 & n3521 ;
  assign n3529 = n3522 ^ n3521 ;
  assign n3530 = n3529 ^ n3520 ;
  assign n3531 = n3530 ^ x46 ;
  assign n3532 = ~n1968 & n3531 ;
  assign n3533 = n3532 ^ x46 ;
  assign n3524 = n3513 ^ n3511 ;
  assign n3523 = n3522 ^ n3520 ;
  assign n3525 = n3524 ^ n3523 ;
  assign n3526 = ~n2006 & n3525 ;
  assign n3527 = n3526 ^ n3525 ;
  assign n3528 = n3527 ^ n3524 ;
  assign n3534 = n3533 ^ n3528 ;
  assign n3535 = n2054 & n3534 ;
  assign n3541 = n3535 ^ n3534 ;
  assign n3542 = n3541 ^ n3533 ;
  assign n3540 = n3526 ^ n3524 ;
  assign n3543 = n3542 ^ n3540 ;
  assign n3544 = n2097 & n3543 ;
  assign n3550 = n3544 ^ n3543 ;
  assign n3551 = n3550 ^ n3542 ;
  assign n3545 = n3544 ^ n3542 ;
  assign n3536 = n3535 ^ n3533 ;
  assign n3537 = n3536 ^ x14 ;
  assign n3538 = ~n2365 & n3537 ;
  assign n3539 = n3538 ^ x14 ;
  assign n3546 = n3545 ^ n3539 ;
  assign n3547 = ~n2410 & n3546 ;
  assign n3548 = n3547 ^ n3546 ;
  assign n3549 = n3548 ^ n3545 ;
  assign n3552 = n3551 ^ n3549 ;
  assign n3553 = ~n2460 & n3552 ;
  assign n3554 = n3553 ^ n3552 ;
  assign n3555 = n3554 ^ n3551 ;
  assign n3556 = x239 ^ x207 ;
  assign n3557 = n1533 & n3556 ;
  assign n3559 = n3557 ^ n3556 ;
  assign n3560 = n3559 ^ x207 ;
  assign n3561 = n3560 ^ x175 ;
  assign n3562 = n1574 & n3561 ;
  assign n3563 = n3562 ^ n3561 ;
  assign n3564 = n3563 ^ x175 ;
  assign n3558 = n3557 ^ x207 ;
  assign n3565 = n3564 ^ n3558 ;
  assign n3566 = n1646 & n3565 ;
  assign n3572 = n3566 ^ n3565 ;
  assign n3573 = n3572 ^ n3564 ;
  assign n3568 = n3562 ^ x175 ;
  assign n3569 = n3568 ^ x143 ;
  assign n3570 = ~n1611 & n3569 ;
  assign n3571 = n3570 ^ x143 ;
  assign n3574 = n3573 ^ n3571 ;
  assign n3575 = ~n1689 & n3574 ;
  assign n3581 = n3575 ^ n3574 ;
  assign n3582 = n3581 ^ n3573 ;
  assign n3583 = n3582 ^ x111 ;
  assign n3584 = ~n1725 & n3583 ;
  assign n3585 = n3584 ^ x111 ;
  assign n3576 = n3575 ^ n3573 ;
  assign n3567 = n3566 ^ n3564 ;
  assign n3577 = n3576 ^ n3567 ;
  assign n3578 = ~n1763 & n3577 ;
  assign n3579 = n3578 ^ n3577 ;
  assign n3580 = n3579 ^ n3576 ;
  assign n3586 = n3585 ^ n3580 ;
  assign n3587 = ~n1810 & n3586 ;
  assign n3594 = n3587 ^ n3586 ;
  assign n3595 = n3594 ^ n3585 ;
  assign n3596 = n3595 ^ x79 ;
  assign n3597 = ~n1846 & n3596 ;
  assign n3598 = n3597 ^ x79 ;
  assign n3589 = n3578 ^ n3576 ;
  assign n3588 = n3587 ^ n3585 ;
  assign n3590 = n3589 ^ n3588 ;
  assign n3591 = ~n1885 & n3590 ;
  assign n3592 = n3591 ^ n3590 ;
  assign n3593 = n3592 ^ n3589 ;
  assign n3599 = n3598 ^ n3593 ;
  assign n3600 = ~n1932 & n3599 ;
  assign n3607 = n3600 ^ n3599 ;
  assign n3608 = n3607 ^ n3598 ;
  assign n3609 = n3608 ^ x47 ;
  assign n3610 = ~n1968 & n3609 ;
  assign n3611 = n3610 ^ x47 ;
  assign n3602 = n3591 ^ n3589 ;
  assign n3601 = n3600 ^ n3598 ;
  assign n3603 = n3602 ^ n3601 ;
  assign n3604 = ~n2006 & n3603 ;
  assign n3605 = n3604 ^ n3603 ;
  assign n3606 = n3605 ^ n3602 ;
  assign n3612 = n3611 ^ n3606 ;
  assign n3613 = n2054 & n3612 ;
  assign n3619 = n3613 ^ n3612 ;
  assign n3620 = n3619 ^ n3611 ;
  assign n3618 = n3604 ^ n3602 ;
  assign n3621 = n3620 ^ n3618 ;
  assign n3622 = n2097 & n3621 ;
  assign n3628 = n3622 ^ n3621 ;
  assign n3629 = n3628 ^ n3620 ;
  assign n3623 = n3622 ^ n3620 ;
  assign n3614 = n3613 ^ n3611 ;
  assign n3615 = n3614 ^ x15 ;
  assign n3616 = ~n2365 & n3615 ;
  assign n3617 = n3616 ^ x15 ;
  assign n3624 = n3623 ^ n3617 ;
  assign n3625 = ~n2410 & n3624 ;
  assign n3626 = n3625 ^ n3624 ;
  assign n3627 = n3626 ^ n3623 ;
  assign n3630 = n3629 ^ n3627 ;
  assign n3631 = ~n2460 & n3630 ;
  assign n3632 = n3631 ^ n3630 ;
  assign n3633 = n3632 ^ n3629 ;
  assign n3634 = x240 ^ x208 ;
  assign n3635 = n1533 & n3634 ;
  assign n3637 = n3635 ^ n3634 ;
  assign n3638 = n3637 ^ x208 ;
  assign n3639 = n3638 ^ x176 ;
  assign n3640 = n1574 & n3639 ;
  assign n3641 = n3640 ^ n3639 ;
  assign n3642 = n3641 ^ x176 ;
  assign n3636 = n3635 ^ x208 ;
  assign n3643 = n3642 ^ n3636 ;
  assign n3644 = n1646 & n3643 ;
  assign n3650 = n3644 ^ n3643 ;
  assign n3651 = n3650 ^ n3642 ;
  assign n3646 = n3640 ^ x176 ;
  assign n3647 = n3646 ^ x144 ;
  assign n3648 = ~n1611 & n3647 ;
  assign n3649 = n3648 ^ x144 ;
  assign n3652 = n3651 ^ n3649 ;
  assign n3653 = ~n1689 & n3652 ;
  assign n3659 = n3653 ^ n3652 ;
  assign n3660 = n3659 ^ n3651 ;
  assign n3661 = n3660 ^ x112 ;
  assign n3662 = ~n1725 & n3661 ;
  assign n3663 = n3662 ^ x112 ;
  assign n3654 = n3653 ^ n3651 ;
  assign n3645 = n3644 ^ n3642 ;
  assign n3655 = n3654 ^ n3645 ;
  assign n3656 = ~n1763 & n3655 ;
  assign n3657 = n3656 ^ n3655 ;
  assign n3658 = n3657 ^ n3654 ;
  assign n3664 = n3663 ^ n3658 ;
  assign n3665 = ~n1810 & n3664 ;
  assign n3672 = n3665 ^ n3664 ;
  assign n3673 = n3672 ^ n3663 ;
  assign n3674 = n3673 ^ x80 ;
  assign n3675 = ~n1846 & n3674 ;
  assign n3676 = n3675 ^ x80 ;
  assign n3667 = n3656 ^ n3654 ;
  assign n3666 = n3665 ^ n3663 ;
  assign n3668 = n3667 ^ n3666 ;
  assign n3669 = ~n1885 & n3668 ;
  assign n3670 = n3669 ^ n3668 ;
  assign n3671 = n3670 ^ n3667 ;
  assign n3677 = n3676 ^ n3671 ;
  assign n3678 = ~n1932 & n3677 ;
  assign n3685 = n3678 ^ n3677 ;
  assign n3686 = n3685 ^ n3676 ;
  assign n3687 = n3686 ^ x48 ;
  assign n3688 = ~n1968 & n3687 ;
  assign n3689 = n3688 ^ x48 ;
  assign n3680 = n3669 ^ n3667 ;
  assign n3679 = n3678 ^ n3676 ;
  assign n3681 = n3680 ^ n3679 ;
  assign n3682 = ~n2006 & n3681 ;
  assign n3683 = n3682 ^ n3681 ;
  assign n3684 = n3683 ^ n3680 ;
  assign n3690 = n3689 ^ n3684 ;
  assign n3691 = n2054 & n3690 ;
  assign n3697 = n3691 ^ n3690 ;
  assign n3698 = n3697 ^ n3689 ;
  assign n3696 = n3682 ^ n3680 ;
  assign n3699 = n3698 ^ n3696 ;
  assign n3700 = n2097 & n3699 ;
  assign n3706 = n3700 ^ n3699 ;
  assign n3707 = n3706 ^ n3698 ;
  assign n3701 = n3700 ^ n3698 ;
  assign n3692 = n3691 ^ n3689 ;
  assign n3693 = n3692 ^ x16 ;
  assign n3694 = ~n2365 & n3693 ;
  assign n3695 = n3694 ^ x16 ;
  assign n3702 = n3701 ^ n3695 ;
  assign n3703 = ~n2410 & n3702 ;
  assign n3704 = n3703 ^ n3702 ;
  assign n3705 = n3704 ^ n3701 ;
  assign n3708 = n3707 ^ n3705 ;
  assign n3709 = ~n2460 & n3708 ;
  assign n3710 = n3709 ^ n3708 ;
  assign n3711 = n3710 ^ n3707 ;
  assign n3712 = x241 ^ x209 ;
  assign n3713 = n1533 & n3712 ;
  assign n3715 = n3713 ^ n3712 ;
  assign n3716 = n3715 ^ x209 ;
  assign n3717 = n3716 ^ x177 ;
  assign n3718 = n1574 & n3717 ;
  assign n3719 = n3718 ^ n3717 ;
  assign n3720 = n3719 ^ x177 ;
  assign n3714 = n3713 ^ x209 ;
  assign n3721 = n3720 ^ n3714 ;
  assign n3722 = n1646 & n3721 ;
  assign n3728 = n3722 ^ n3721 ;
  assign n3729 = n3728 ^ n3720 ;
  assign n3724 = n3718 ^ x177 ;
  assign n3725 = n3724 ^ x145 ;
  assign n3726 = ~n1611 & n3725 ;
  assign n3727 = n3726 ^ x145 ;
  assign n3730 = n3729 ^ n3727 ;
  assign n3731 = ~n1689 & n3730 ;
  assign n3737 = n3731 ^ n3730 ;
  assign n3738 = n3737 ^ n3729 ;
  assign n3739 = n3738 ^ x113 ;
  assign n3740 = ~n1725 & n3739 ;
  assign n3741 = n3740 ^ x113 ;
  assign n3732 = n3731 ^ n3729 ;
  assign n3723 = n3722 ^ n3720 ;
  assign n3733 = n3732 ^ n3723 ;
  assign n3734 = ~n1763 & n3733 ;
  assign n3735 = n3734 ^ n3733 ;
  assign n3736 = n3735 ^ n3732 ;
  assign n3742 = n3741 ^ n3736 ;
  assign n3743 = ~n1810 & n3742 ;
  assign n3750 = n3743 ^ n3742 ;
  assign n3751 = n3750 ^ n3741 ;
  assign n3752 = n3751 ^ x81 ;
  assign n3753 = ~n1846 & n3752 ;
  assign n3754 = n3753 ^ x81 ;
  assign n3745 = n3734 ^ n3732 ;
  assign n3744 = n3743 ^ n3741 ;
  assign n3746 = n3745 ^ n3744 ;
  assign n3747 = ~n1885 & n3746 ;
  assign n3748 = n3747 ^ n3746 ;
  assign n3749 = n3748 ^ n3745 ;
  assign n3755 = n3754 ^ n3749 ;
  assign n3756 = ~n1932 & n3755 ;
  assign n3763 = n3756 ^ n3755 ;
  assign n3764 = n3763 ^ n3754 ;
  assign n3765 = n3764 ^ x49 ;
  assign n3766 = ~n1968 & n3765 ;
  assign n3767 = n3766 ^ x49 ;
  assign n3758 = n3747 ^ n3745 ;
  assign n3757 = n3756 ^ n3754 ;
  assign n3759 = n3758 ^ n3757 ;
  assign n3760 = ~n2006 & n3759 ;
  assign n3761 = n3760 ^ n3759 ;
  assign n3762 = n3761 ^ n3758 ;
  assign n3768 = n3767 ^ n3762 ;
  assign n3769 = n2054 & n3768 ;
  assign n3775 = n3769 ^ n3768 ;
  assign n3776 = n3775 ^ n3767 ;
  assign n3774 = n3760 ^ n3758 ;
  assign n3777 = n3776 ^ n3774 ;
  assign n3778 = n2097 & n3777 ;
  assign n3784 = n3778 ^ n3777 ;
  assign n3785 = n3784 ^ n3776 ;
  assign n3779 = n3778 ^ n3776 ;
  assign n3770 = n3769 ^ n3767 ;
  assign n3771 = n3770 ^ x17 ;
  assign n3772 = ~n2365 & n3771 ;
  assign n3773 = n3772 ^ x17 ;
  assign n3780 = n3779 ^ n3773 ;
  assign n3781 = ~n2410 & n3780 ;
  assign n3782 = n3781 ^ n3780 ;
  assign n3783 = n3782 ^ n3779 ;
  assign n3786 = n3785 ^ n3783 ;
  assign n3787 = ~n2460 & n3786 ;
  assign n3788 = n3787 ^ n3786 ;
  assign n3789 = n3788 ^ n3785 ;
  assign n3790 = x242 ^ x210 ;
  assign n3791 = n1533 & n3790 ;
  assign n3793 = n3791 ^ n3790 ;
  assign n3794 = n3793 ^ x210 ;
  assign n3795 = n3794 ^ x178 ;
  assign n3796 = n1574 & n3795 ;
  assign n3797 = n3796 ^ n3795 ;
  assign n3798 = n3797 ^ x178 ;
  assign n3792 = n3791 ^ x210 ;
  assign n3799 = n3798 ^ n3792 ;
  assign n3800 = n1646 & n3799 ;
  assign n3806 = n3800 ^ n3799 ;
  assign n3807 = n3806 ^ n3798 ;
  assign n3802 = n3796 ^ x178 ;
  assign n3803 = n3802 ^ x146 ;
  assign n3804 = ~n1611 & n3803 ;
  assign n3805 = n3804 ^ x146 ;
  assign n3808 = n3807 ^ n3805 ;
  assign n3809 = ~n1689 & n3808 ;
  assign n3815 = n3809 ^ n3808 ;
  assign n3816 = n3815 ^ n3807 ;
  assign n3817 = n3816 ^ x114 ;
  assign n3818 = ~n1725 & n3817 ;
  assign n3819 = n3818 ^ x114 ;
  assign n3810 = n3809 ^ n3807 ;
  assign n3801 = n3800 ^ n3798 ;
  assign n3811 = n3810 ^ n3801 ;
  assign n3812 = ~n1763 & n3811 ;
  assign n3813 = n3812 ^ n3811 ;
  assign n3814 = n3813 ^ n3810 ;
  assign n3820 = n3819 ^ n3814 ;
  assign n3821 = ~n1810 & n3820 ;
  assign n3828 = n3821 ^ n3820 ;
  assign n3829 = n3828 ^ n3819 ;
  assign n3830 = n3829 ^ x82 ;
  assign n3831 = ~n1846 & n3830 ;
  assign n3832 = n3831 ^ x82 ;
  assign n3823 = n3812 ^ n3810 ;
  assign n3822 = n3821 ^ n3819 ;
  assign n3824 = n3823 ^ n3822 ;
  assign n3825 = ~n1885 & n3824 ;
  assign n3826 = n3825 ^ n3824 ;
  assign n3827 = n3826 ^ n3823 ;
  assign n3833 = n3832 ^ n3827 ;
  assign n3834 = ~n1932 & n3833 ;
  assign n3841 = n3834 ^ n3833 ;
  assign n3842 = n3841 ^ n3832 ;
  assign n3843 = n3842 ^ x50 ;
  assign n3844 = ~n1968 & n3843 ;
  assign n3845 = n3844 ^ x50 ;
  assign n3836 = n3825 ^ n3823 ;
  assign n3835 = n3834 ^ n3832 ;
  assign n3837 = n3836 ^ n3835 ;
  assign n3838 = ~n2006 & n3837 ;
  assign n3839 = n3838 ^ n3837 ;
  assign n3840 = n3839 ^ n3836 ;
  assign n3846 = n3845 ^ n3840 ;
  assign n3847 = n2054 & n3846 ;
  assign n3853 = n3847 ^ n3846 ;
  assign n3854 = n3853 ^ n3845 ;
  assign n3852 = n3838 ^ n3836 ;
  assign n3855 = n3854 ^ n3852 ;
  assign n3856 = n2097 & n3855 ;
  assign n3862 = n3856 ^ n3855 ;
  assign n3863 = n3862 ^ n3854 ;
  assign n3857 = n3856 ^ n3854 ;
  assign n3848 = n3847 ^ n3845 ;
  assign n3849 = n3848 ^ x18 ;
  assign n3850 = ~n2365 & n3849 ;
  assign n3851 = n3850 ^ x18 ;
  assign n3858 = n3857 ^ n3851 ;
  assign n3859 = ~n2410 & n3858 ;
  assign n3860 = n3859 ^ n3858 ;
  assign n3861 = n3860 ^ n3857 ;
  assign n3864 = n3863 ^ n3861 ;
  assign n3865 = ~n2460 & n3864 ;
  assign n3866 = n3865 ^ n3864 ;
  assign n3867 = n3866 ^ n3863 ;
  assign n3868 = x243 ^ x211 ;
  assign n3869 = n1533 & n3868 ;
  assign n3871 = n3869 ^ n3868 ;
  assign n3872 = n3871 ^ x211 ;
  assign n3873 = n3872 ^ x179 ;
  assign n3874 = n1574 & n3873 ;
  assign n3875 = n3874 ^ n3873 ;
  assign n3876 = n3875 ^ x179 ;
  assign n3870 = n3869 ^ x211 ;
  assign n3877 = n3876 ^ n3870 ;
  assign n3878 = n1646 & n3877 ;
  assign n3884 = n3878 ^ n3877 ;
  assign n3885 = n3884 ^ n3876 ;
  assign n3880 = n3874 ^ x179 ;
  assign n3881 = n3880 ^ x147 ;
  assign n3882 = ~n1611 & n3881 ;
  assign n3883 = n3882 ^ x147 ;
  assign n3886 = n3885 ^ n3883 ;
  assign n3887 = ~n1689 & n3886 ;
  assign n3893 = n3887 ^ n3886 ;
  assign n3894 = n3893 ^ n3885 ;
  assign n3895 = n3894 ^ x115 ;
  assign n3896 = ~n1725 & n3895 ;
  assign n3897 = n3896 ^ x115 ;
  assign n3888 = n3887 ^ n3885 ;
  assign n3879 = n3878 ^ n3876 ;
  assign n3889 = n3888 ^ n3879 ;
  assign n3890 = ~n1763 & n3889 ;
  assign n3891 = n3890 ^ n3889 ;
  assign n3892 = n3891 ^ n3888 ;
  assign n3898 = n3897 ^ n3892 ;
  assign n3899 = ~n1810 & n3898 ;
  assign n3906 = n3899 ^ n3898 ;
  assign n3907 = n3906 ^ n3897 ;
  assign n3908 = n3907 ^ x83 ;
  assign n3909 = ~n1846 & n3908 ;
  assign n3910 = n3909 ^ x83 ;
  assign n3901 = n3890 ^ n3888 ;
  assign n3900 = n3899 ^ n3897 ;
  assign n3902 = n3901 ^ n3900 ;
  assign n3903 = ~n1885 & n3902 ;
  assign n3904 = n3903 ^ n3902 ;
  assign n3905 = n3904 ^ n3901 ;
  assign n3911 = n3910 ^ n3905 ;
  assign n3912 = ~n1932 & n3911 ;
  assign n3919 = n3912 ^ n3911 ;
  assign n3920 = n3919 ^ n3910 ;
  assign n3921 = n3920 ^ x51 ;
  assign n3922 = ~n1968 & n3921 ;
  assign n3923 = n3922 ^ x51 ;
  assign n3914 = n3903 ^ n3901 ;
  assign n3913 = n3912 ^ n3910 ;
  assign n3915 = n3914 ^ n3913 ;
  assign n3916 = ~n2006 & n3915 ;
  assign n3917 = n3916 ^ n3915 ;
  assign n3918 = n3917 ^ n3914 ;
  assign n3924 = n3923 ^ n3918 ;
  assign n3925 = n2054 & n3924 ;
  assign n3931 = n3925 ^ n3924 ;
  assign n3932 = n3931 ^ n3923 ;
  assign n3930 = n3916 ^ n3914 ;
  assign n3933 = n3932 ^ n3930 ;
  assign n3934 = n2097 & n3933 ;
  assign n3940 = n3934 ^ n3933 ;
  assign n3941 = n3940 ^ n3932 ;
  assign n3935 = n3934 ^ n3932 ;
  assign n3926 = n3925 ^ n3923 ;
  assign n3927 = n3926 ^ x19 ;
  assign n3928 = ~n2365 & n3927 ;
  assign n3929 = n3928 ^ x19 ;
  assign n3936 = n3935 ^ n3929 ;
  assign n3937 = ~n2410 & n3936 ;
  assign n3938 = n3937 ^ n3936 ;
  assign n3939 = n3938 ^ n3935 ;
  assign n3942 = n3941 ^ n3939 ;
  assign n3943 = ~n2460 & n3942 ;
  assign n3944 = n3943 ^ n3942 ;
  assign n3945 = n3944 ^ n3941 ;
  assign n3946 = x244 ^ x212 ;
  assign n3947 = n1533 & n3946 ;
  assign n3949 = n3947 ^ n3946 ;
  assign n3950 = n3949 ^ x212 ;
  assign n3951 = n3950 ^ x180 ;
  assign n3952 = n1574 & n3951 ;
  assign n3953 = n3952 ^ n3951 ;
  assign n3954 = n3953 ^ x180 ;
  assign n3948 = n3947 ^ x212 ;
  assign n3955 = n3954 ^ n3948 ;
  assign n3956 = n1646 & n3955 ;
  assign n3962 = n3956 ^ n3955 ;
  assign n3963 = n3962 ^ n3954 ;
  assign n3958 = n3952 ^ x180 ;
  assign n3959 = n3958 ^ x148 ;
  assign n3960 = ~n1611 & n3959 ;
  assign n3961 = n3960 ^ x148 ;
  assign n3964 = n3963 ^ n3961 ;
  assign n3965 = ~n1689 & n3964 ;
  assign n3971 = n3965 ^ n3964 ;
  assign n3972 = n3971 ^ n3963 ;
  assign n3973 = n3972 ^ x116 ;
  assign n3974 = ~n1725 & n3973 ;
  assign n3975 = n3974 ^ x116 ;
  assign n3966 = n3965 ^ n3963 ;
  assign n3957 = n3956 ^ n3954 ;
  assign n3967 = n3966 ^ n3957 ;
  assign n3968 = ~n1763 & n3967 ;
  assign n3969 = n3968 ^ n3967 ;
  assign n3970 = n3969 ^ n3966 ;
  assign n3976 = n3975 ^ n3970 ;
  assign n3977 = ~n1810 & n3976 ;
  assign n3984 = n3977 ^ n3976 ;
  assign n3985 = n3984 ^ n3975 ;
  assign n3986 = n3985 ^ x84 ;
  assign n3987 = ~n1846 & n3986 ;
  assign n3988 = n3987 ^ x84 ;
  assign n3979 = n3968 ^ n3966 ;
  assign n3978 = n3977 ^ n3975 ;
  assign n3980 = n3979 ^ n3978 ;
  assign n3981 = ~n1885 & n3980 ;
  assign n3982 = n3981 ^ n3980 ;
  assign n3983 = n3982 ^ n3979 ;
  assign n3989 = n3988 ^ n3983 ;
  assign n3990 = ~n1932 & n3989 ;
  assign n3997 = n3990 ^ n3989 ;
  assign n3998 = n3997 ^ n3988 ;
  assign n3999 = n3998 ^ x52 ;
  assign n4000 = ~n1968 & n3999 ;
  assign n4001 = n4000 ^ x52 ;
  assign n3992 = n3981 ^ n3979 ;
  assign n3991 = n3990 ^ n3988 ;
  assign n3993 = n3992 ^ n3991 ;
  assign n3994 = ~n2006 & n3993 ;
  assign n3995 = n3994 ^ n3993 ;
  assign n3996 = n3995 ^ n3992 ;
  assign n4002 = n4001 ^ n3996 ;
  assign n4003 = n2054 & n4002 ;
  assign n4009 = n4003 ^ n4002 ;
  assign n4010 = n4009 ^ n4001 ;
  assign n4008 = n3994 ^ n3992 ;
  assign n4011 = n4010 ^ n4008 ;
  assign n4012 = n2097 & n4011 ;
  assign n4018 = n4012 ^ n4011 ;
  assign n4019 = n4018 ^ n4010 ;
  assign n4013 = n4012 ^ n4010 ;
  assign n4004 = n4003 ^ n4001 ;
  assign n4005 = n4004 ^ x20 ;
  assign n4006 = ~n2365 & n4005 ;
  assign n4007 = n4006 ^ x20 ;
  assign n4014 = n4013 ^ n4007 ;
  assign n4015 = ~n2410 & n4014 ;
  assign n4016 = n4015 ^ n4014 ;
  assign n4017 = n4016 ^ n4013 ;
  assign n4020 = n4019 ^ n4017 ;
  assign n4021 = ~n2460 & n4020 ;
  assign n4022 = n4021 ^ n4020 ;
  assign n4023 = n4022 ^ n4019 ;
  assign n4024 = x245 ^ x213 ;
  assign n4025 = n1533 & n4024 ;
  assign n4027 = n4025 ^ n4024 ;
  assign n4028 = n4027 ^ x213 ;
  assign n4029 = n4028 ^ x181 ;
  assign n4030 = n1574 & n4029 ;
  assign n4031 = n4030 ^ n4029 ;
  assign n4032 = n4031 ^ x181 ;
  assign n4026 = n4025 ^ x213 ;
  assign n4033 = n4032 ^ n4026 ;
  assign n4034 = n1646 & n4033 ;
  assign n4040 = n4034 ^ n4033 ;
  assign n4041 = n4040 ^ n4032 ;
  assign n4036 = n4030 ^ x181 ;
  assign n4037 = n4036 ^ x149 ;
  assign n4038 = ~n1611 & n4037 ;
  assign n4039 = n4038 ^ x149 ;
  assign n4042 = n4041 ^ n4039 ;
  assign n4043 = ~n1689 & n4042 ;
  assign n4049 = n4043 ^ n4042 ;
  assign n4050 = n4049 ^ n4041 ;
  assign n4051 = n4050 ^ x117 ;
  assign n4052 = ~n1725 & n4051 ;
  assign n4053 = n4052 ^ x117 ;
  assign n4044 = n4043 ^ n4041 ;
  assign n4035 = n4034 ^ n4032 ;
  assign n4045 = n4044 ^ n4035 ;
  assign n4046 = ~n1763 & n4045 ;
  assign n4047 = n4046 ^ n4045 ;
  assign n4048 = n4047 ^ n4044 ;
  assign n4054 = n4053 ^ n4048 ;
  assign n4055 = ~n1810 & n4054 ;
  assign n4062 = n4055 ^ n4054 ;
  assign n4063 = n4062 ^ n4053 ;
  assign n4064 = n4063 ^ x85 ;
  assign n4065 = ~n1846 & n4064 ;
  assign n4066 = n4065 ^ x85 ;
  assign n4057 = n4046 ^ n4044 ;
  assign n4056 = n4055 ^ n4053 ;
  assign n4058 = n4057 ^ n4056 ;
  assign n4059 = ~n1885 & n4058 ;
  assign n4060 = n4059 ^ n4058 ;
  assign n4061 = n4060 ^ n4057 ;
  assign n4067 = n4066 ^ n4061 ;
  assign n4068 = ~n1932 & n4067 ;
  assign n4075 = n4068 ^ n4067 ;
  assign n4076 = n4075 ^ n4066 ;
  assign n4077 = n4076 ^ x53 ;
  assign n4078 = ~n1968 & n4077 ;
  assign n4079 = n4078 ^ x53 ;
  assign n4070 = n4059 ^ n4057 ;
  assign n4069 = n4068 ^ n4066 ;
  assign n4071 = n4070 ^ n4069 ;
  assign n4072 = ~n2006 & n4071 ;
  assign n4073 = n4072 ^ n4071 ;
  assign n4074 = n4073 ^ n4070 ;
  assign n4080 = n4079 ^ n4074 ;
  assign n4081 = n2054 & n4080 ;
  assign n4087 = n4081 ^ n4080 ;
  assign n4088 = n4087 ^ n4079 ;
  assign n4086 = n4072 ^ n4070 ;
  assign n4089 = n4088 ^ n4086 ;
  assign n4090 = n2097 & n4089 ;
  assign n4096 = n4090 ^ n4089 ;
  assign n4097 = n4096 ^ n4088 ;
  assign n4091 = n4090 ^ n4088 ;
  assign n4082 = n4081 ^ n4079 ;
  assign n4083 = n4082 ^ x21 ;
  assign n4084 = ~n2365 & n4083 ;
  assign n4085 = n4084 ^ x21 ;
  assign n4092 = n4091 ^ n4085 ;
  assign n4093 = ~n2410 & n4092 ;
  assign n4094 = n4093 ^ n4092 ;
  assign n4095 = n4094 ^ n4091 ;
  assign n4098 = n4097 ^ n4095 ;
  assign n4099 = ~n2460 & n4098 ;
  assign n4100 = n4099 ^ n4098 ;
  assign n4101 = n4100 ^ n4097 ;
  assign n4102 = x246 ^ x214 ;
  assign n4103 = n1533 & n4102 ;
  assign n4105 = n4103 ^ n4102 ;
  assign n4106 = n4105 ^ x214 ;
  assign n4107 = n4106 ^ x182 ;
  assign n4108 = n1574 & n4107 ;
  assign n4109 = n4108 ^ n4107 ;
  assign n4110 = n4109 ^ x182 ;
  assign n4104 = n4103 ^ x214 ;
  assign n4111 = n4110 ^ n4104 ;
  assign n4112 = n1646 & n4111 ;
  assign n4118 = n4112 ^ n4111 ;
  assign n4119 = n4118 ^ n4110 ;
  assign n4114 = n4108 ^ x182 ;
  assign n4115 = n4114 ^ x150 ;
  assign n4116 = ~n1611 & n4115 ;
  assign n4117 = n4116 ^ x150 ;
  assign n4120 = n4119 ^ n4117 ;
  assign n4121 = ~n1689 & n4120 ;
  assign n4127 = n4121 ^ n4120 ;
  assign n4128 = n4127 ^ n4119 ;
  assign n4129 = n4128 ^ x118 ;
  assign n4130 = ~n1725 & n4129 ;
  assign n4131 = n4130 ^ x118 ;
  assign n4122 = n4121 ^ n4119 ;
  assign n4113 = n4112 ^ n4110 ;
  assign n4123 = n4122 ^ n4113 ;
  assign n4124 = ~n1763 & n4123 ;
  assign n4125 = n4124 ^ n4123 ;
  assign n4126 = n4125 ^ n4122 ;
  assign n4132 = n4131 ^ n4126 ;
  assign n4133 = ~n1810 & n4132 ;
  assign n4140 = n4133 ^ n4132 ;
  assign n4141 = n4140 ^ n4131 ;
  assign n4142 = n4141 ^ x86 ;
  assign n4143 = ~n1846 & n4142 ;
  assign n4144 = n4143 ^ x86 ;
  assign n4135 = n4124 ^ n4122 ;
  assign n4134 = n4133 ^ n4131 ;
  assign n4136 = n4135 ^ n4134 ;
  assign n4137 = ~n1885 & n4136 ;
  assign n4138 = n4137 ^ n4136 ;
  assign n4139 = n4138 ^ n4135 ;
  assign n4145 = n4144 ^ n4139 ;
  assign n4146 = ~n1932 & n4145 ;
  assign n4153 = n4146 ^ n4145 ;
  assign n4154 = n4153 ^ n4144 ;
  assign n4155 = n4154 ^ x54 ;
  assign n4156 = ~n1968 & n4155 ;
  assign n4157 = n4156 ^ x54 ;
  assign n4148 = n4137 ^ n4135 ;
  assign n4147 = n4146 ^ n4144 ;
  assign n4149 = n4148 ^ n4147 ;
  assign n4150 = ~n2006 & n4149 ;
  assign n4151 = n4150 ^ n4149 ;
  assign n4152 = n4151 ^ n4148 ;
  assign n4158 = n4157 ^ n4152 ;
  assign n4159 = n2054 & n4158 ;
  assign n4165 = n4159 ^ n4158 ;
  assign n4166 = n4165 ^ n4157 ;
  assign n4164 = n4150 ^ n4148 ;
  assign n4167 = n4166 ^ n4164 ;
  assign n4168 = n2097 & n4167 ;
  assign n4174 = n4168 ^ n4167 ;
  assign n4175 = n4174 ^ n4166 ;
  assign n4169 = n4168 ^ n4166 ;
  assign n4160 = n4159 ^ n4157 ;
  assign n4161 = n4160 ^ x22 ;
  assign n4162 = ~n2365 & n4161 ;
  assign n4163 = n4162 ^ x22 ;
  assign n4170 = n4169 ^ n4163 ;
  assign n4171 = ~n2410 & n4170 ;
  assign n4172 = n4171 ^ n4170 ;
  assign n4173 = n4172 ^ n4169 ;
  assign n4176 = n4175 ^ n4173 ;
  assign n4177 = ~n2460 & n4176 ;
  assign n4178 = n4177 ^ n4176 ;
  assign n4179 = n4178 ^ n4175 ;
  assign n4180 = x247 ^ x215 ;
  assign n4181 = n1533 & n4180 ;
  assign n4183 = n4181 ^ n4180 ;
  assign n4184 = n4183 ^ x215 ;
  assign n4185 = n4184 ^ x183 ;
  assign n4186 = n1574 & n4185 ;
  assign n4187 = n4186 ^ n4185 ;
  assign n4188 = n4187 ^ x183 ;
  assign n4182 = n4181 ^ x215 ;
  assign n4189 = n4188 ^ n4182 ;
  assign n4190 = n1646 & n4189 ;
  assign n4196 = n4190 ^ n4189 ;
  assign n4197 = n4196 ^ n4188 ;
  assign n4192 = n4186 ^ x183 ;
  assign n4193 = n4192 ^ x151 ;
  assign n4194 = ~n1611 & n4193 ;
  assign n4195 = n4194 ^ x151 ;
  assign n4198 = n4197 ^ n4195 ;
  assign n4199 = ~n1689 & n4198 ;
  assign n4205 = n4199 ^ n4198 ;
  assign n4206 = n4205 ^ n4197 ;
  assign n4207 = n4206 ^ x119 ;
  assign n4208 = ~n1725 & n4207 ;
  assign n4209 = n4208 ^ x119 ;
  assign n4200 = n4199 ^ n4197 ;
  assign n4191 = n4190 ^ n4188 ;
  assign n4201 = n4200 ^ n4191 ;
  assign n4202 = ~n1763 & n4201 ;
  assign n4203 = n4202 ^ n4201 ;
  assign n4204 = n4203 ^ n4200 ;
  assign n4210 = n4209 ^ n4204 ;
  assign n4211 = ~n1810 & n4210 ;
  assign n4218 = n4211 ^ n4210 ;
  assign n4219 = n4218 ^ n4209 ;
  assign n4220 = n4219 ^ x87 ;
  assign n4221 = ~n1846 & n4220 ;
  assign n4222 = n4221 ^ x87 ;
  assign n4213 = n4202 ^ n4200 ;
  assign n4212 = n4211 ^ n4209 ;
  assign n4214 = n4213 ^ n4212 ;
  assign n4215 = ~n1885 & n4214 ;
  assign n4216 = n4215 ^ n4214 ;
  assign n4217 = n4216 ^ n4213 ;
  assign n4223 = n4222 ^ n4217 ;
  assign n4224 = ~n1932 & n4223 ;
  assign n4231 = n4224 ^ n4223 ;
  assign n4232 = n4231 ^ n4222 ;
  assign n4233 = n4232 ^ x55 ;
  assign n4234 = ~n1968 & n4233 ;
  assign n4235 = n4234 ^ x55 ;
  assign n4226 = n4215 ^ n4213 ;
  assign n4225 = n4224 ^ n4222 ;
  assign n4227 = n4226 ^ n4225 ;
  assign n4228 = ~n2006 & n4227 ;
  assign n4229 = n4228 ^ n4227 ;
  assign n4230 = n4229 ^ n4226 ;
  assign n4236 = n4235 ^ n4230 ;
  assign n4237 = n2054 & n4236 ;
  assign n4243 = n4237 ^ n4236 ;
  assign n4244 = n4243 ^ n4235 ;
  assign n4242 = n4228 ^ n4226 ;
  assign n4245 = n4244 ^ n4242 ;
  assign n4246 = n2097 & n4245 ;
  assign n4252 = n4246 ^ n4245 ;
  assign n4253 = n4252 ^ n4244 ;
  assign n4247 = n4246 ^ n4244 ;
  assign n4238 = n4237 ^ n4235 ;
  assign n4239 = n4238 ^ x23 ;
  assign n4240 = ~n2365 & n4239 ;
  assign n4241 = n4240 ^ x23 ;
  assign n4248 = n4247 ^ n4241 ;
  assign n4249 = ~n2410 & n4248 ;
  assign n4250 = n4249 ^ n4248 ;
  assign n4251 = n4250 ^ n4247 ;
  assign n4254 = n4253 ^ n4251 ;
  assign n4255 = ~n2460 & n4254 ;
  assign n4256 = n4255 ^ n4254 ;
  assign n4257 = n4256 ^ n4253 ;
  assign n4258 = x248 ^ x216 ;
  assign n4259 = n1533 & n4258 ;
  assign n4261 = n4259 ^ n4258 ;
  assign n4262 = n4261 ^ x216 ;
  assign n4263 = n4262 ^ x184 ;
  assign n4264 = n1574 & n4263 ;
  assign n4265 = n4264 ^ n4263 ;
  assign n4266 = n4265 ^ x184 ;
  assign n4260 = n4259 ^ x216 ;
  assign n4267 = n4266 ^ n4260 ;
  assign n4268 = n1646 & n4267 ;
  assign n4274 = n4268 ^ n4267 ;
  assign n4275 = n4274 ^ n4266 ;
  assign n4270 = n4264 ^ x184 ;
  assign n4271 = n4270 ^ x152 ;
  assign n4272 = ~n1611 & n4271 ;
  assign n4273 = n4272 ^ x152 ;
  assign n4276 = n4275 ^ n4273 ;
  assign n4277 = ~n1689 & n4276 ;
  assign n4283 = n4277 ^ n4276 ;
  assign n4284 = n4283 ^ n4275 ;
  assign n4285 = n4284 ^ x120 ;
  assign n4286 = ~n1725 & n4285 ;
  assign n4287 = n4286 ^ x120 ;
  assign n4278 = n4277 ^ n4275 ;
  assign n4269 = n4268 ^ n4266 ;
  assign n4279 = n4278 ^ n4269 ;
  assign n4280 = ~n1763 & n4279 ;
  assign n4281 = n4280 ^ n4279 ;
  assign n4282 = n4281 ^ n4278 ;
  assign n4288 = n4287 ^ n4282 ;
  assign n4289 = ~n1810 & n4288 ;
  assign n4296 = n4289 ^ n4288 ;
  assign n4297 = n4296 ^ n4287 ;
  assign n4298 = n4297 ^ x88 ;
  assign n4299 = ~n1846 & n4298 ;
  assign n4300 = n4299 ^ x88 ;
  assign n4291 = n4280 ^ n4278 ;
  assign n4290 = n4289 ^ n4287 ;
  assign n4292 = n4291 ^ n4290 ;
  assign n4293 = ~n1885 & n4292 ;
  assign n4294 = n4293 ^ n4292 ;
  assign n4295 = n4294 ^ n4291 ;
  assign n4301 = n4300 ^ n4295 ;
  assign n4302 = ~n1932 & n4301 ;
  assign n4309 = n4302 ^ n4301 ;
  assign n4310 = n4309 ^ n4300 ;
  assign n4311 = n4310 ^ x56 ;
  assign n4312 = ~n1968 & n4311 ;
  assign n4313 = n4312 ^ x56 ;
  assign n4304 = n4293 ^ n4291 ;
  assign n4303 = n4302 ^ n4300 ;
  assign n4305 = n4304 ^ n4303 ;
  assign n4306 = ~n2006 & n4305 ;
  assign n4307 = n4306 ^ n4305 ;
  assign n4308 = n4307 ^ n4304 ;
  assign n4314 = n4313 ^ n4308 ;
  assign n4315 = n2054 & n4314 ;
  assign n4321 = n4315 ^ n4314 ;
  assign n4322 = n4321 ^ n4313 ;
  assign n4320 = n4306 ^ n4304 ;
  assign n4323 = n4322 ^ n4320 ;
  assign n4324 = n2097 & n4323 ;
  assign n4330 = n4324 ^ n4323 ;
  assign n4331 = n4330 ^ n4322 ;
  assign n4325 = n4324 ^ n4322 ;
  assign n4316 = n4315 ^ n4313 ;
  assign n4317 = n4316 ^ x24 ;
  assign n4318 = ~n2365 & n4317 ;
  assign n4319 = n4318 ^ x24 ;
  assign n4326 = n4325 ^ n4319 ;
  assign n4327 = ~n2410 & n4326 ;
  assign n4328 = n4327 ^ n4326 ;
  assign n4329 = n4328 ^ n4325 ;
  assign n4332 = n4331 ^ n4329 ;
  assign n4333 = ~n2460 & n4332 ;
  assign n4334 = n4333 ^ n4332 ;
  assign n4335 = n4334 ^ n4331 ;
  assign n4336 = x249 ^ x217 ;
  assign n4337 = n1533 & n4336 ;
  assign n4339 = n4337 ^ n4336 ;
  assign n4340 = n4339 ^ x217 ;
  assign n4341 = n4340 ^ x185 ;
  assign n4342 = n1574 & n4341 ;
  assign n4343 = n4342 ^ n4341 ;
  assign n4344 = n4343 ^ x185 ;
  assign n4338 = n4337 ^ x217 ;
  assign n4345 = n4344 ^ n4338 ;
  assign n4346 = n1646 & n4345 ;
  assign n4352 = n4346 ^ n4345 ;
  assign n4353 = n4352 ^ n4344 ;
  assign n4348 = n4342 ^ x185 ;
  assign n4349 = n4348 ^ x153 ;
  assign n4350 = ~n1611 & n4349 ;
  assign n4351 = n4350 ^ x153 ;
  assign n4354 = n4353 ^ n4351 ;
  assign n4355 = ~n1689 & n4354 ;
  assign n4361 = n4355 ^ n4354 ;
  assign n4362 = n4361 ^ n4353 ;
  assign n4363 = n4362 ^ x121 ;
  assign n4364 = ~n1725 & n4363 ;
  assign n4365 = n4364 ^ x121 ;
  assign n4356 = n4355 ^ n4353 ;
  assign n4347 = n4346 ^ n4344 ;
  assign n4357 = n4356 ^ n4347 ;
  assign n4358 = ~n1763 & n4357 ;
  assign n4359 = n4358 ^ n4357 ;
  assign n4360 = n4359 ^ n4356 ;
  assign n4366 = n4365 ^ n4360 ;
  assign n4367 = ~n1810 & n4366 ;
  assign n4374 = n4367 ^ n4366 ;
  assign n4375 = n4374 ^ n4365 ;
  assign n4376 = n4375 ^ x89 ;
  assign n4377 = ~n1846 & n4376 ;
  assign n4378 = n4377 ^ x89 ;
  assign n4369 = n4358 ^ n4356 ;
  assign n4368 = n4367 ^ n4365 ;
  assign n4370 = n4369 ^ n4368 ;
  assign n4371 = ~n1885 & n4370 ;
  assign n4372 = n4371 ^ n4370 ;
  assign n4373 = n4372 ^ n4369 ;
  assign n4379 = n4378 ^ n4373 ;
  assign n4380 = ~n1932 & n4379 ;
  assign n4387 = n4380 ^ n4379 ;
  assign n4388 = n4387 ^ n4378 ;
  assign n4389 = n4388 ^ x57 ;
  assign n4390 = ~n1968 & n4389 ;
  assign n4391 = n4390 ^ x57 ;
  assign n4382 = n4371 ^ n4369 ;
  assign n4381 = n4380 ^ n4378 ;
  assign n4383 = n4382 ^ n4381 ;
  assign n4384 = ~n2006 & n4383 ;
  assign n4385 = n4384 ^ n4383 ;
  assign n4386 = n4385 ^ n4382 ;
  assign n4392 = n4391 ^ n4386 ;
  assign n4393 = n2054 & n4392 ;
  assign n4399 = n4393 ^ n4392 ;
  assign n4400 = n4399 ^ n4391 ;
  assign n4398 = n4384 ^ n4382 ;
  assign n4401 = n4400 ^ n4398 ;
  assign n4402 = n2097 & n4401 ;
  assign n4408 = n4402 ^ n4401 ;
  assign n4409 = n4408 ^ n4400 ;
  assign n4403 = n4402 ^ n4400 ;
  assign n4394 = n4393 ^ n4391 ;
  assign n4395 = n4394 ^ x25 ;
  assign n4396 = ~n2365 & n4395 ;
  assign n4397 = n4396 ^ x25 ;
  assign n4404 = n4403 ^ n4397 ;
  assign n4405 = ~n2410 & n4404 ;
  assign n4406 = n4405 ^ n4404 ;
  assign n4407 = n4406 ^ n4403 ;
  assign n4410 = n4409 ^ n4407 ;
  assign n4411 = ~n2460 & n4410 ;
  assign n4412 = n4411 ^ n4410 ;
  assign n4413 = n4412 ^ n4409 ;
  assign n4414 = x250 ^ x218 ;
  assign n4415 = n1533 & n4414 ;
  assign n4417 = n4415 ^ n4414 ;
  assign n4418 = n4417 ^ x218 ;
  assign n4419 = n4418 ^ x186 ;
  assign n4420 = n1574 & n4419 ;
  assign n4421 = n4420 ^ n4419 ;
  assign n4422 = n4421 ^ x186 ;
  assign n4416 = n4415 ^ x218 ;
  assign n4423 = n4422 ^ n4416 ;
  assign n4424 = n1646 & n4423 ;
  assign n4430 = n4424 ^ n4423 ;
  assign n4431 = n4430 ^ n4422 ;
  assign n4426 = n4420 ^ x186 ;
  assign n4427 = n4426 ^ x154 ;
  assign n4428 = ~n1611 & n4427 ;
  assign n4429 = n4428 ^ x154 ;
  assign n4432 = n4431 ^ n4429 ;
  assign n4433 = ~n1689 & n4432 ;
  assign n4439 = n4433 ^ n4432 ;
  assign n4440 = n4439 ^ n4431 ;
  assign n4441 = n4440 ^ x122 ;
  assign n4442 = ~n1725 & n4441 ;
  assign n4443 = n4442 ^ x122 ;
  assign n4434 = n4433 ^ n4431 ;
  assign n4425 = n4424 ^ n4422 ;
  assign n4435 = n4434 ^ n4425 ;
  assign n4436 = ~n1763 & n4435 ;
  assign n4437 = n4436 ^ n4435 ;
  assign n4438 = n4437 ^ n4434 ;
  assign n4444 = n4443 ^ n4438 ;
  assign n4445 = ~n1810 & n4444 ;
  assign n4452 = n4445 ^ n4444 ;
  assign n4453 = n4452 ^ n4443 ;
  assign n4454 = n4453 ^ x90 ;
  assign n4455 = ~n1846 & n4454 ;
  assign n4456 = n4455 ^ x90 ;
  assign n4447 = n4436 ^ n4434 ;
  assign n4446 = n4445 ^ n4443 ;
  assign n4448 = n4447 ^ n4446 ;
  assign n4449 = ~n1885 & n4448 ;
  assign n4450 = n4449 ^ n4448 ;
  assign n4451 = n4450 ^ n4447 ;
  assign n4457 = n4456 ^ n4451 ;
  assign n4458 = ~n1932 & n4457 ;
  assign n4465 = n4458 ^ n4457 ;
  assign n4466 = n4465 ^ n4456 ;
  assign n4467 = n4466 ^ x58 ;
  assign n4468 = ~n1968 & n4467 ;
  assign n4469 = n4468 ^ x58 ;
  assign n4460 = n4449 ^ n4447 ;
  assign n4459 = n4458 ^ n4456 ;
  assign n4461 = n4460 ^ n4459 ;
  assign n4462 = ~n2006 & n4461 ;
  assign n4463 = n4462 ^ n4461 ;
  assign n4464 = n4463 ^ n4460 ;
  assign n4470 = n4469 ^ n4464 ;
  assign n4471 = n2054 & n4470 ;
  assign n4477 = n4471 ^ n4470 ;
  assign n4478 = n4477 ^ n4469 ;
  assign n4476 = n4462 ^ n4460 ;
  assign n4479 = n4478 ^ n4476 ;
  assign n4480 = n2097 & n4479 ;
  assign n4486 = n4480 ^ n4479 ;
  assign n4487 = n4486 ^ n4478 ;
  assign n4481 = n4480 ^ n4478 ;
  assign n4472 = n4471 ^ n4469 ;
  assign n4473 = n4472 ^ x26 ;
  assign n4474 = ~n2365 & n4473 ;
  assign n4475 = n4474 ^ x26 ;
  assign n4482 = n4481 ^ n4475 ;
  assign n4483 = ~n2410 & n4482 ;
  assign n4484 = n4483 ^ n4482 ;
  assign n4485 = n4484 ^ n4481 ;
  assign n4488 = n4487 ^ n4485 ;
  assign n4489 = ~n2460 & n4488 ;
  assign n4490 = n4489 ^ n4488 ;
  assign n4491 = n4490 ^ n4487 ;
  assign n4492 = x251 ^ x219 ;
  assign n4493 = n1533 & n4492 ;
  assign n4495 = n4493 ^ n4492 ;
  assign n4496 = n4495 ^ x219 ;
  assign n4497 = n4496 ^ x187 ;
  assign n4498 = n1574 & n4497 ;
  assign n4499 = n4498 ^ n4497 ;
  assign n4500 = n4499 ^ x187 ;
  assign n4494 = n4493 ^ x219 ;
  assign n4501 = n4500 ^ n4494 ;
  assign n4502 = n1646 & n4501 ;
  assign n4508 = n4502 ^ n4501 ;
  assign n4509 = n4508 ^ n4500 ;
  assign n4504 = n4498 ^ x187 ;
  assign n4505 = n4504 ^ x155 ;
  assign n4506 = ~n1611 & n4505 ;
  assign n4507 = n4506 ^ x155 ;
  assign n4510 = n4509 ^ n4507 ;
  assign n4511 = ~n1689 & n4510 ;
  assign n4517 = n4511 ^ n4510 ;
  assign n4518 = n4517 ^ n4509 ;
  assign n4519 = n4518 ^ x123 ;
  assign n4520 = ~n1725 & n4519 ;
  assign n4521 = n4520 ^ x123 ;
  assign n4512 = n4511 ^ n4509 ;
  assign n4503 = n4502 ^ n4500 ;
  assign n4513 = n4512 ^ n4503 ;
  assign n4514 = ~n1763 & n4513 ;
  assign n4515 = n4514 ^ n4513 ;
  assign n4516 = n4515 ^ n4512 ;
  assign n4522 = n4521 ^ n4516 ;
  assign n4523 = ~n1810 & n4522 ;
  assign n4530 = n4523 ^ n4522 ;
  assign n4531 = n4530 ^ n4521 ;
  assign n4532 = n4531 ^ x91 ;
  assign n4533 = ~n1846 & n4532 ;
  assign n4534 = n4533 ^ x91 ;
  assign n4525 = n4514 ^ n4512 ;
  assign n4524 = n4523 ^ n4521 ;
  assign n4526 = n4525 ^ n4524 ;
  assign n4527 = ~n1885 & n4526 ;
  assign n4528 = n4527 ^ n4526 ;
  assign n4529 = n4528 ^ n4525 ;
  assign n4535 = n4534 ^ n4529 ;
  assign n4536 = ~n1932 & n4535 ;
  assign n4543 = n4536 ^ n4535 ;
  assign n4544 = n4543 ^ n4534 ;
  assign n4545 = n4544 ^ x59 ;
  assign n4546 = ~n1968 & n4545 ;
  assign n4547 = n4546 ^ x59 ;
  assign n4538 = n4527 ^ n4525 ;
  assign n4537 = n4536 ^ n4534 ;
  assign n4539 = n4538 ^ n4537 ;
  assign n4540 = ~n2006 & n4539 ;
  assign n4541 = n4540 ^ n4539 ;
  assign n4542 = n4541 ^ n4538 ;
  assign n4548 = n4547 ^ n4542 ;
  assign n4549 = n2054 & n4548 ;
  assign n4555 = n4549 ^ n4548 ;
  assign n4556 = n4555 ^ n4547 ;
  assign n4554 = n4540 ^ n4538 ;
  assign n4557 = n4556 ^ n4554 ;
  assign n4558 = n2097 & n4557 ;
  assign n4564 = n4558 ^ n4557 ;
  assign n4565 = n4564 ^ n4556 ;
  assign n4559 = n4558 ^ n4556 ;
  assign n4550 = n4549 ^ n4547 ;
  assign n4551 = n4550 ^ x27 ;
  assign n4552 = ~n2365 & n4551 ;
  assign n4553 = n4552 ^ x27 ;
  assign n4560 = n4559 ^ n4553 ;
  assign n4561 = ~n2410 & n4560 ;
  assign n4562 = n4561 ^ n4560 ;
  assign n4563 = n4562 ^ n4559 ;
  assign n4566 = n4565 ^ n4563 ;
  assign n4567 = ~n2460 & n4566 ;
  assign n4568 = n4567 ^ n4566 ;
  assign n4569 = n4568 ^ n4565 ;
  assign n4570 = x252 ^ x220 ;
  assign n4571 = n1533 & n4570 ;
  assign n4573 = n4571 ^ n4570 ;
  assign n4574 = n4573 ^ x220 ;
  assign n4575 = n4574 ^ x188 ;
  assign n4576 = n1574 & n4575 ;
  assign n4577 = n4576 ^ n4575 ;
  assign n4578 = n4577 ^ x188 ;
  assign n4572 = n4571 ^ x220 ;
  assign n4579 = n4578 ^ n4572 ;
  assign n4580 = n1646 & n4579 ;
  assign n4586 = n4580 ^ n4579 ;
  assign n4587 = n4586 ^ n4578 ;
  assign n4582 = n4576 ^ x188 ;
  assign n4583 = n4582 ^ x156 ;
  assign n4584 = ~n1611 & n4583 ;
  assign n4585 = n4584 ^ x156 ;
  assign n4588 = n4587 ^ n4585 ;
  assign n4589 = ~n1689 & n4588 ;
  assign n4595 = n4589 ^ n4588 ;
  assign n4596 = n4595 ^ n4587 ;
  assign n4597 = n4596 ^ x124 ;
  assign n4598 = ~n1725 & n4597 ;
  assign n4599 = n4598 ^ x124 ;
  assign n4590 = n4589 ^ n4587 ;
  assign n4581 = n4580 ^ n4578 ;
  assign n4591 = n4590 ^ n4581 ;
  assign n4592 = ~n1763 & n4591 ;
  assign n4593 = n4592 ^ n4591 ;
  assign n4594 = n4593 ^ n4590 ;
  assign n4600 = n4599 ^ n4594 ;
  assign n4601 = ~n1810 & n4600 ;
  assign n4608 = n4601 ^ n4600 ;
  assign n4609 = n4608 ^ n4599 ;
  assign n4610 = n4609 ^ x92 ;
  assign n4611 = ~n1846 & n4610 ;
  assign n4612 = n4611 ^ x92 ;
  assign n4603 = n4592 ^ n4590 ;
  assign n4602 = n4601 ^ n4599 ;
  assign n4604 = n4603 ^ n4602 ;
  assign n4605 = ~n1885 & n4604 ;
  assign n4606 = n4605 ^ n4604 ;
  assign n4607 = n4606 ^ n4603 ;
  assign n4613 = n4612 ^ n4607 ;
  assign n4614 = ~n1932 & n4613 ;
  assign n4621 = n4614 ^ n4613 ;
  assign n4622 = n4621 ^ n4612 ;
  assign n4623 = n4622 ^ x60 ;
  assign n4624 = ~n1968 & n4623 ;
  assign n4625 = n4624 ^ x60 ;
  assign n4616 = n4605 ^ n4603 ;
  assign n4615 = n4614 ^ n4612 ;
  assign n4617 = n4616 ^ n4615 ;
  assign n4618 = ~n2006 & n4617 ;
  assign n4619 = n4618 ^ n4617 ;
  assign n4620 = n4619 ^ n4616 ;
  assign n4626 = n4625 ^ n4620 ;
  assign n4627 = n2054 & n4626 ;
  assign n4633 = n4627 ^ n4626 ;
  assign n4634 = n4633 ^ n4625 ;
  assign n4632 = n4618 ^ n4616 ;
  assign n4635 = n4634 ^ n4632 ;
  assign n4636 = n2097 & n4635 ;
  assign n4642 = n4636 ^ n4635 ;
  assign n4643 = n4642 ^ n4634 ;
  assign n4637 = n4636 ^ n4634 ;
  assign n4628 = n4627 ^ n4625 ;
  assign n4629 = n4628 ^ x28 ;
  assign n4630 = ~n2365 & n4629 ;
  assign n4631 = n4630 ^ x28 ;
  assign n4638 = n4637 ^ n4631 ;
  assign n4639 = ~n2410 & n4638 ;
  assign n4640 = n4639 ^ n4638 ;
  assign n4641 = n4640 ^ n4637 ;
  assign n4644 = n4643 ^ n4641 ;
  assign n4645 = ~n2460 & n4644 ;
  assign n4646 = n4645 ^ n4644 ;
  assign n4647 = n4646 ^ n4643 ;
  assign n4648 = x253 ^ x221 ;
  assign n4649 = n1533 & n4648 ;
  assign n4651 = n4649 ^ n4648 ;
  assign n4652 = n4651 ^ x221 ;
  assign n4653 = n4652 ^ x189 ;
  assign n4654 = n1574 & n4653 ;
  assign n4655 = n4654 ^ n4653 ;
  assign n4656 = n4655 ^ x189 ;
  assign n4650 = n4649 ^ x221 ;
  assign n4657 = n4656 ^ n4650 ;
  assign n4658 = n1646 & n4657 ;
  assign n4664 = n4658 ^ n4657 ;
  assign n4665 = n4664 ^ n4656 ;
  assign n4660 = n4654 ^ x189 ;
  assign n4661 = n4660 ^ x157 ;
  assign n4662 = ~n1611 & n4661 ;
  assign n4663 = n4662 ^ x157 ;
  assign n4666 = n4665 ^ n4663 ;
  assign n4667 = ~n1689 & n4666 ;
  assign n4673 = n4667 ^ n4666 ;
  assign n4674 = n4673 ^ n4665 ;
  assign n4675 = n4674 ^ x125 ;
  assign n4676 = ~n1725 & n4675 ;
  assign n4677 = n4676 ^ x125 ;
  assign n4668 = n4667 ^ n4665 ;
  assign n4659 = n4658 ^ n4656 ;
  assign n4669 = n4668 ^ n4659 ;
  assign n4670 = ~n1763 & n4669 ;
  assign n4671 = n4670 ^ n4669 ;
  assign n4672 = n4671 ^ n4668 ;
  assign n4678 = n4677 ^ n4672 ;
  assign n4679 = ~n1810 & n4678 ;
  assign n4686 = n4679 ^ n4678 ;
  assign n4687 = n4686 ^ n4677 ;
  assign n4688 = n4687 ^ x93 ;
  assign n4689 = ~n1846 & n4688 ;
  assign n4690 = n4689 ^ x93 ;
  assign n4681 = n4670 ^ n4668 ;
  assign n4680 = n4679 ^ n4677 ;
  assign n4682 = n4681 ^ n4680 ;
  assign n4683 = ~n1885 & n4682 ;
  assign n4684 = n4683 ^ n4682 ;
  assign n4685 = n4684 ^ n4681 ;
  assign n4691 = n4690 ^ n4685 ;
  assign n4692 = ~n1932 & n4691 ;
  assign n4699 = n4692 ^ n4691 ;
  assign n4700 = n4699 ^ n4690 ;
  assign n4701 = n4700 ^ x61 ;
  assign n4702 = ~n1968 & n4701 ;
  assign n4703 = n4702 ^ x61 ;
  assign n4694 = n4683 ^ n4681 ;
  assign n4693 = n4692 ^ n4690 ;
  assign n4695 = n4694 ^ n4693 ;
  assign n4696 = ~n2006 & n4695 ;
  assign n4697 = n4696 ^ n4695 ;
  assign n4698 = n4697 ^ n4694 ;
  assign n4704 = n4703 ^ n4698 ;
  assign n4705 = n2054 & n4704 ;
  assign n4711 = n4705 ^ n4704 ;
  assign n4712 = n4711 ^ n4703 ;
  assign n4710 = n4696 ^ n4694 ;
  assign n4713 = n4712 ^ n4710 ;
  assign n4714 = n2097 & n4713 ;
  assign n4720 = n4714 ^ n4713 ;
  assign n4721 = n4720 ^ n4712 ;
  assign n4715 = n4714 ^ n4712 ;
  assign n4706 = n4705 ^ n4703 ;
  assign n4707 = n4706 ^ x29 ;
  assign n4708 = ~n2365 & n4707 ;
  assign n4709 = n4708 ^ x29 ;
  assign n4716 = n4715 ^ n4709 ;
  assign n4717 = ~n2410 & n4716 ;
  assign n4718 = n4717 ^ n4716 ;
  assign n4719 = n4718 ^ n4715 ;
  assign n4722 = n4721 ^ n4719 ;
  assign n4723 = ~n2460 & n4722 ;
  assign n4724 = n4723 ^ n4722 ;
  assign n4725 = n4724 ^ n4721 ;
  assign n4726 = x254 ^ x222 ;
  assign n4727 = n1533 & n4726 ;
  assign n4729 = n4727 ^ n4726 ;
  assign n4730 = n4729 ^ x222 ;
  assign n4731 = n4730 ^ x190 ;
  assign n4732 = n1574 & n4731 ;
  assign n4733 = n4732 ^ n4731 ;
  assign n4734 = n4733 ^ x190 ;
  assign n4728 = n4727 ^ x222 ;
  assign n4735 = n4734 ^ n4728 ;
  assign n4736 = n1646 & n4735 ;
  assign n4742 = n4736 ^ n4735 ;
  assign n4743 = n4742 ^ n4734 ;
  assign n4738 = n4732 ^ x190 ;
  assign n4739 = n4738 ^ x158 ;
  assign n4740 = ~n1611 & n4739 ;
  assign n4741 = n4740 ^ x158 ;
  assign n4744 = n4743 ^ n4741 ;
  assign n4745 = ~n1689 & n4744 ;
  assign n4751 = n4745 ^ n4744 ;
  assign n4752 = n4751 ^ n4743 ;
  assign n4753 = n4752 ^ x126 ;
  assign n4754 = ~n1725 & n4753 ;
  assign n4755 = n4754 ^ x126 ;
  assign n4746 = n4745 ^ n4743 ;
  assign n4737 = n4736 ^ n4734 ;
  assign n4747 = n4746 ^ n4737 ;
  assign n4748 = ~n1763 & n4747 ;
  assign n4749 = n4748 ^ n4747 ;
  assign n4750 = n4749 ^ n4746 ;
  assign n4756 = n4755 ^ n4750 ;
  assign n4757 = ~n1810 & n4756 ;
  assign n4764 = n4757 ^ n4756 ;
  assign n4765 = n4764 ^ n4755 ;
  assign n4766 = n4765 ^ x94 ;
  assign n4767 = ~n1846 & n4766 ;
  assign n4768 = n4767 ^ x94 ;
  assign n4759 = n4748 ^ n4746 ;
  assign n4758 = n4757 ^ n4755 ;
  assign n4760 = n4759 ^ n4758 ;
  assign n4761 = ~n1885 & n4760 ;
  assign n4762 = n4761 ^ n4760 ;
  assign n4763 = n4762 ^ n4759 ;
  assign n4769 = n4768 ^ n4763 ;
  assign n4770 = ~n1932 & n4769 ;
  assign n4777 = n4770 ^ n4769 ;
  assign n4778 = n4777 ^ n4768 ;
  assign n4779 = n4778 ^ x62 ;
  assign n4780 = ~n1968 & n4779 ;
  assign n4781 = n4780 ^ x62 ;
  assign n4772 = n4761 ^ n4759 ;
  assign n4771 = n4770 ^ n4768 ;
  assign n4773 = n4772 ^ n4771 ;
  assign n4774 = ~n2006 & n4773 ;
  assign n4775 = n4774 ^ n4773 ;
  assign n4776 = n4775 ^ n4772 ;
  assign n4782 = n4781 ^ n4776 ;
  assign n4783 = n2054 & n4782 ;
  assign n4789 = n4783 ^ n4782 ;
  assign n4790 = n4789 ^ n4781 ;
  assign n4788 = n4774 ^ n4772 ;
  assign n4791 = n4790 ^ n4788 ;
  assign n4792 = n2097 & n4791 ;
  assign n4798 = n4792 ^ n4791 ;
  assign n4799 = n4798 ^ n4790 ;
  assign n4793 = n4792 ^ n4790 ;
  assign n4784 = n4783 ^ n4781 ;
  assign n4785 = n4784 ^ x30 ;
  assign n4786 = ~n2365 & n4785 ;
  assign n4787 = n4786 ^ x30 ;
  assign n4794 = n4793 ^ n4787 ;
  assign n4795 = ~n2410 & n4794 ;
  assign n4796 = n4795 ^ n4794 ;
  assign n4797 = n4796 ^ n4793 ;
  assign n4800 = n4799 ^ n4797 ;
  assign n4801 = ~n2460 & n4800 ;
  assign n4802 = n4801 ^ n4800 ;
  assign n4803 = n4802 ^ n4799 ;
  assign n4804 = x255 ^ x223 ;
  assign n4805 = n1533 & n4804 ;
  assign n4807 = n4805 ^ n4804 ;
  assign n4808 = n4807 ^ x223 ;
  assign n4809 = n4808 ^ x191 ;
  assign n4810 = n1574 & n4809 ;
  assign n4811 = n4810 ^ n4809 ;
  assign n4812 = n4811 ^ x191 ;
  assign n4806 = n4805 ^ x223 ;
  assign n4813 = n4812 ^ n4806 ;
  assign n4814 = n1646 & n4813 ;
  assign n4820 = n4814 ^ n4813 ;
  assign n4821 = n4820 ^ n4812 ;
  assign n4816 = n4810 ^ x191 ;
  assign n4817 = n4816 ^ x159 ;
  assign n4818 = ~n1611 & n4817 ;
  assign n4819 = n4818 ^ x159 ;
  assign n4822 = n4821 ^ n4819 ;
  assign n4823 = ~n1689 & n4822 ;
  assign n4829 = n4823 ^ n4822 ;
  assign n4830 = n4829 ^ n4821 ;
  assign n4831 = n4830 ^ x127 ;
  assign n4832 = ~n1725 & n4831 ;
  assign n4833 = n4832 ^ x127 ;
  assign n4824 = n4823 ^ n4821 ;
  assign n4815 = n4814 ^ n4812 ;
  assign n4825 = n4824 ^ n4815 ;
  assign n4826 = ~n1763 & n4825 ;
  assign n4827 = n4826 ^ n4825 ;
  assign n4828 = n4827 ^ n4824 ;
  assign n4834 = n4833 ^ n4828 ;
  assign n4835 = ~n1810 & n4834 ;
  assign n4842 = n4835 ^ n4834 ;
  assign n4843 = n4842 ^ n4833 ;
  assign n4844 = n4843 ^ x95 ;
  assign n4845 = ~n1846 & n4844 ;
  assign n4846 = n4845 ^ x95 ;
  assign n4837 = n4826 ^ n4824 ;
  assign n4836 = n4835 ^ n4833 ;
  assign n4838 = n4837 ^ n4836 ;
  assign n4839 = ~n1885 & n4838 ;
  assign n4840 = n4839 ^ n4838 ;
  assign n4841 = n4840 ^ n4837 ;
  assign n4847 = n4846 ^ n4841 ;
  assign n4848 = ~n1932 & n4847 ;
  assign n4855 = n4848 ^ n4847 ;
  assign n4856 = n4855 ^ n4846 ;
  assign n4857 = n4856 ^ x63 ;
  assign n4858 = ~n1968 & n4857 ;
  assign n4859 = n4858 ^ x63 ;
  assign n4850 = n4839 ^ n4837 ;
  assign n4849 = n4848 ^ n4846 ;
  assign n4851 = n4850 ^ n4849 ;
  assign n4852 = ~n2006 & n4851 ;
  assign n4853 = n4852 ^ n4851 ;
  assign n4854 = n4853 ^ n4850 ;
  assign n4860 = n4859 ^ n4854 ;
  assign n4861 = n2054 & n4860 ;
  assign n4867 = n4861 ^ n4860 ;
  assign n4868 = n4867 ^ n4859 ;
  assign n4866 = n4852 ^ n4850 ;
  assign n4869 = n4868 ^ n4866 ;
  assign n4870 = n2097 & n4869 ;
  assign n4876 = n4870 ^ n4869 ;
  assign n4877 = n4876 ^ n4868 ;
  assign n4871 = n4870 ^ n4868 ;
  assign n4862 = n4861 ^ n4859 ;
  assign n4863 = n4862 ^ x31 ;
  assign n4864 = ~n2365 & n4863 ;
  assign n4865 = n4864 ^ x31 ;
  assign n4872 = n4871 ^ n4865 ;
  assign n4873 = ~n2410 & n4872 ;
  assign n4874 = n4873 ^ n4872 ;
  assign n4875 = n4874 ^ n4871 ;
  assign n4878 = n4877 ^ n4875 ;
  assign n4879 = ~n2460 & n4878 ;
  assign n4880 = n4879 ^ n4878 ;
  assign n4881 = n4880 ^ n4877 ;
  assign n4882 = n2461 ^ n2421 ;
  assign n4883 = n2539 ^ n2537 ;
  assign n4884 = n2617 ^ n2615 ;
  assign n4885 = n2695 ^ n2693 ;
  assign n4886 = n2773 ^ n2771 ;
  assign n4887 = n2851 ^ n2849 ;
  assign n4888 = n2929 ^ n2927 ;
  assign n4889 = n3007 ^ n3005 ;
  assign n4890 = n3085 ^ n3083 ;
  assign n4891 = n3163 ^ n3161 ;
  assign n4892 = n3241 ^ n3239 ;
  assign n4893 = n3319 ^ n3317 ;
  assign n4894 = n3397 ^ n3395 ;
  assign n4895 = n3475 ^ n3473 ;
  assign n4896 = n3553 ^ n3551 ;
  assign n4897 = n3631 ^ n3629 ;
  assign n4898 = n3709 ^ n3707 ;
  assign n4899 = n3787 ^ n3785 ;
  assign n4900 = n3865 ^ n3863 ;
  assign n4901 = n3943 ^ n3941 ;
  assign n4902 = n4021 ^ n4019 ;
  assign n4903 = n4099 ^ n4097 ;
  assign n4904 = n4177 ^ n4175 ;
  assign n4905 = n4255 ^ n4253 ;
  assign n4906 = n4333 ^ n4331 ;
  assign n4907 = n4411 ^ n4409 ;
  assign n4908 = n4489 ^ n4487 ;
  assign n4909 = n4567 ^ n4565 ;
  assign n4910 = n4645 ^ n4643 ;
  assign n4911 = n4723 ^ n4721 ;
  assign n4912 = n4801 ^ n4799 ;
  assign n4913 = n4879 ^ n4877 ;
  assign n4914 = n2419 ^ n2417 ;
  assign n4915 = n2533 ^ n2531 ;
  assign n4916 = n2611 ^ n2609 ;
  assign n4917 = n2689 ^ n2687 ;
  assign n4918 = n2767 ^ n2765 ;
  assign n4919 = n2845 ^ n2843 ;
  assign n4920 = n2923 ^ n2921 ;
  assign n4921 = n3001 ^ n2999 ;
  assign n4922 = n3079 ^ n3077 ;
  assign n4923 = n3157 ^ n3155 ;
  assign n4924 = n3235 ^ n3233 ;
  assign n4925 = n3313 ^ n3311 ;
  assign n4926 = n3391 ^ n3389 ;
  assign n4927 = n3469 ^ n3467 ;
  assign n4928 = n3547 ^ n3545 ;
  assign n4929 = n3625 ^ n3623 ;
  assign n4930 = n3703 ^ n3701 ;
  assign n4931 = n3781 ^ n3779 ;
  assign n4932 = n3859 ^ n3857 ;
  assign n4933 = n3937 ^ n3935 ;
  assign n4934 = n4015 ^ n4013 ;
  assign n4935 = n4093 ^ n4091 ;
  assign n4936 = n4171 ^ n4169 ;
  assign n4937 = n4249 ^ n4247 ;
  assign n4938 = n4327 ^ n4325 ;
  assign n4939 = n4405 ^ n4403 ;
  assign n4940 = n4483 ^ n4481 ;
  assign n4941 = n4561 ^ n4559 ;
  assign n4942 = n4639 ^ n4637 ;
  assign n4943 = n4717 ^ n4715 ;
  assign n4944 = n4795 ^ n4793 ;
  assign n4945 = n4873 ^ n4871 ;
  assign y0 = n2463 ;
  assign y1 = n2541 ;
  assign y2 = n2619 ;
  assign y3 = n2697 ;
  assign y4 = n2775 ;
  assign y5 = n2853 ;
  assign y6 = n2931 ;
  assign y7 = n3009 ;
  assign y8 = n3087 ;
  assign y9 = n3165 ;
  assign y10 = n3243 ;
  assign y11 = n3321 ;
  assign y12 = n3399 ;
  assign y13 = n3477 ;
  assign y14 = n3555 ;
  assign y15 = n3633 ;
  assign y16 = n3711 ;
  assign y17 = n3789 ;
  assign y18 = n3867 ;
  assign y19 = n3945 ;
  assign y20 = n4023 ;
  assign y21 = n4101 ;
  assign y22 = n4179 ;
  assign y23 = n4257 ;
  assign y24 = n4335 ;
  assign y25 = n4413 ;
  assign y26 = n4491 ;
  assign y27 = n4569 ;
  assign y28 = n4647 ;
  assign y29 = n4725 ;
  assign y30 = n4803 ;
  assign y31 = n4881 ;
  assign y32 = n4882 ;
  assign y33 = n4883 ;
  assign y34 = n4884 ;
  assign y35 = n4885 ;
  assign y36 = n4886 ;
  assign y37 = n4887 ;
  assign y38 = n4888 ;
  assign y39 = n4889 ;
  assign y40 = n4890 ;
  assign y41 = n4891 ;
  assign y42 = n4892 ;
  assign y43 = n4893 ;
  assign y44 = n4894 ;
  assign y45 = n4895 ;
  assign y46 = n4896 ;
  assign y47 = n4897 ;
  assign y48 = n4898 ;
  assign y49 = n4899 ;
  assign y50 = n4900 ;
  assign y51 = n4901 ;
  assign y52 = n4902 ;
  assign y53 = n4903 ;
  assign y54 = n4904 ;
  assign y55 = n4905 ;
  assign y56 = n4906 ;
  assign y57 = n4907 ;
  assign y58 = n4908 ;
  assign y59 = n4909 ;
  assign y60 = n4910 ;
  assign y61 = n4911 ;
  assign y62 = n4912 ;
  assign y63 = n4913 ;
  assign y64 = n4914 ;
  assign y65 = n4915 ;
  assign y66 = n4916 ;
  assign y67 = n4917 ;
  assign y68 = n4918 ;
  assign y69 = n4919 ;
  assign y70 = n4920 ;
  assign y71 = n4921 ;
  assign y72 = n4922 ;
  assign y73 = n4923 ;
  assign y74 = n4924 ;
  assign y75 = n4925 ;
  assign y76 = n4926 ;
  assign y77 = n4927 ;
  assign y78 = n4928 ;
  assign y79 = n4929 ;
  assign y80 = n4930 ;
  assign y81 = n4931 ;
  assign y82 = n4932 ;
  assign y83 = n4933 ;
  assign y84 = n4934 ;
  assign y85 = n4935 ;
  assign y86 = n4936 ;
  assign y87 = n4937 ;
  assign y88 = n4938 ;
  assign y89 = n4939 ;
  assign y90 = n4940 ;
  assign y91 = n4941 ;
  assign y92 = n4942 ;
  assign y93 = n4943 ;
  assign y94 = n4944 ;
  assign y95 = n4945 ;
endmodule
