// 16 parties, each holding 32-bit data
module auction_N_4_W_32_opt( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 ;
  assign n520 = ~x31 & ~x63 ;
  assign n521 = ~x95 & ~x127 ;
  assign n522 = n520 & n521 ;
  assign n523 = ~x159 & ~x191 ;
  assign n524 = ~x223 & ~x255 ;
  assign n525 = n523 & n524 ;
  assign n526 = n522 & n525 ;
  assign n513 = ~x287 & ~x319 ;
  assign n514 = ~x351 & ~x383 ;
  assign n515 = n513 & n514 ;
  assign n516 = ~x415 & ~x447 ;
  assign n517 = ~x479 & ~x511 ;
  assign n518 = n516 & n517 ;
  assign n519 = n515 & n518 ;
  assign n527 = n526 ^ n519 ;
  assign n2518 = x446 ^ x414 ;
  assign n2519 = x447 ^ x415 ;
  assign n2521 = x444 ^ x412 ;
  assign n2523 = x442 ^ x410 ;
  assign n2525 = x440 ^ x408 ;
  assign n2527 = x438 ^ x406 ;
  assign n2529 = x436 ^ x404 ;
  assign n2531 = x434 ^ x402 ;
  assign n2533 = x432 ^ x400 ;
  assign n2535 = x430 ^ x398 ;
  assign n2537 = x428 ^ x396 ;
  assign n2539 = x426 ^ x394 ;
  assign n2541 = x424 ^ x392 ;
  assign n2543 = x422 ^ x390 ;
  assign n2545 = x420 ^ x388 ;
  assign n2547 = x418 ^ x386 ;
  assign n2549 = x384 & ~x416 ;
  assign n2550 = n2549 ^ x418 ;
  assign n2548 = x418 ^ x385 ;
  assign n2551 = n2550 ^ n2548 ;
  assign n2552 = x417 ^ x385 ;
  assign n2553 = n2551 & ~n2552 ;
  assign n2554 = n2553 ^ n2548 ;
  assign n2555 = ~n2547 & n2554 ;
  assign n2556 = n2555 ^ x386 ;
  assign n2557 = n2556 ^ x420 ;
  assign n2546 = x420 ^ x387 ;
  assign n2558 = n2557 ^ n2546 ;
  assign n2559 = x419 ^ x387 ;
  assign n2560 = n2558 & ~n2559 ;
  assign n2561 = n2560 ^ n2546 ;
  assign n2562 = ~n2545 & n2561 ;
  assign n2563 = n2562 ^ x388 ;
  assign n2564 = n2563 ^ x422 ;
  assign n2544 = x422 ^ x389 ;
  assign n2565 = n2564 ^ n2544 ;
  assign n2566 = x421 ^ x389 ;
  assign n2567 = n2565 & ~n2566 ;
  assign n2568 = n2567 ^ n2544 ;
  assign n2569 = ~n2543 & n2568 ;
  assign n2570 = n2569 ^ x390 ;
  assign n2571 = n2570 ^ x424 ;
  assign n2542 = x424 ^ x391 ;
  assign n2572 = n2571 ^ n2542 ;
  assign n2573 = x423 ^ x391 ;
  assign n2574 = n2572 & ~n2573 ;
  assign n2575 = n2574 ^ n2542 ;
  assign n2576 = ~n2541 & n2575 ;
  assign n2577 = n2576 ^ x392 ;
  assign n2578 = n2577 ^ x426 ;
  assign n2540 = x426 ^ x393 ;
  assign n2579 = n2578 ^ n2540 ;
  assign n2580 = x425 ^ x393 ;
  assign n2581 = n2579 & ~n2580 ;
  assign n2582 = n2581 ^ n2540 ;
  assign n2583 = ~n2539 & n2582 ;
  assign n2584 = n2583 ^ x394 ;
  assign n2585 = n2584 ^ x428 ;
  assign n2538 = x428 ^ x395 ;
  assign n2586 = n2585 ^ n2538 ;
  assign n2587 = x427 ^ x395 ;
  assign n2588 = n2586 & ~n2587 ;
  assign n2589 = n2588 ^ n2538 ;
  assign n2590 = ~n2537 & n2589 ;
  assign n2591 = n2590 ^ x396 ;
  assign n2592 = n2591 ^ x430 ;
  assign n2536 = x430 ^ x397 ;
  assign n2593 = n2592 ^ n2536 ;
  assign n2594 = x429 ^ x397 ;
  assign n2595 = n2593 & ~n2594 ;
  assign n2596 = n2595 ^ n2536 ;
  assign n2597 = ~n2535 & n2596 ;
  assign n2598 = n2597 ^ x398 ;
  assign n2599 = n2598 ^ x432 ;
  assign n2534 = x432 ^ x399 ;
  assign n2600 = n2599 ^ n2534 ;
  assign n2601 = x431 ^ x399 ;
  assign n2602 = n2600 & ~n2601 ;
  assign n2603 = n2602 ^ n2534 ;
  assign n2604 = ~n2533 & n2603 ;
  assign n2605 = n2604 ^ x400 ;
  assign n2606 = n2605 ^ x434 ;
  assign n2532 = x434 ^ x401 ;
  assign n2607 = n2606 ^ n2532 ;
  assign n2608 = x433 ^ x401 ;
  assign n2609 = n2607 & ~n2608 ;
  assign n2610 = n2609 ^ n2532 ;
  assign n2611 = ~n2531 & n2610 ;
  assign n2612 = n2611 ^ x402 ;
  assign n2613 = n2612 ^ x436 ;
  assign n2530 = x436 ^ x403 ;
  assign n2614 = n2613 ^ n2530 ;
  assign n2615 = x435 ^ x403 ;
  assign n2616 = n2614 & ~n2615 ;
  assign n2617 = n2616 ^ n2530 ;
  assign n2618 = ~n2529 & n2617 ;
  assign n2619 = n2618 ^ x404 ;
  assign n2620 = n2619 ^ x438 ;
  assign n2528 = x438 ^ x405 ;
  assign n2621 = n2620 ^ n2528 ;
  assign n2622 = x437 ^ x405 ;
  assign n2623 = n2621 & ~n2622 ;
  assign n2624 = n2623 ^ n2528 ;
  assign n2625 = ~n2527 & n2624 ;
  assign n2626 = n2625 ^ x406 ;
  assign n2627 = n2626 ^ x440 ;
  assign n2526 = x440 ^ x407 ;
  assign n2628 = n2627 ^ n2526 ;
  assign n2629 = x439 ^ x407 ;
  assign n2630 = n2628 & ~n2629 ;
  assign n2631 = n2630 ^ n2526 ;
  assign n2632 = ~n2525 & n2631 ;
  assign n2633 = n2632 ^ x408 ;
  assign n2634 = n2633 ^ x442 ;
  assign n2524 = x442 ^ x409 ;
  assign n2635 = n2634 ^ n2524 ;
  assign n2636 = x441 ^ x409 ;
  assign n2637 = n2635 & ~n2636 ;
  assign n2638 = n2637 ^ n2524 ;
  assign n2639 = ~n2523 & n2638 ;
  assign n2640 = n2639 ^ x410 ;
  assign n2641 = n2640 ^ x444 ;
  assign n2522 = x444 ^ x411 ;
  assign n2642 = n2641 ^ n2522 ;
  assign n2643 = x443 ^ x411 ;
  assign n2644 = n2642 & ~n2643 ;
  assign n2645 = n2644 ^ n2522 ;
  assign n2646 = ~n2521 & n2645 ;
  assign n2647 = n2646 ^ x412 ;
  assign n2648 = n2647 ^ x446 ;
  assign n2520 = x446 ^ x413 ;
  assign n2649 = n2648 ^ n2520 ;
  assign n2650 = x445 ^ x413 ;
  assign n2651 = n2649 & ~n2650 ;
  assign n2652 = n2651 ^ n2520 ;
  assign n2653 = ~n2518 & n2652 ;
  assign n2654 = n2653 ^ x414 ;
  assign n2655 = n2654 ^ x447 ;
  assign n2656 = ~n2519 & n2655 ;
  assign n2657 = n2656 ^ x415 ;
  assign n2658 = n2518 & ~n2657 ;
  assign n2659 = n2658 ^ x414 ;
  assign n2376 = x510 ^ x478 ;
  assign n2377 = x511 ^ x479 ;
  assign n2379 = x508 ^ x476 ;
  assign n2381 = x506 ^ x474 ;
  assign n2383 = x504 ^ x472 ;
  assign n2385 = x502 ^ x470 ;
  assign n2387 = x500 ^ x468 ;
  assign n2389 = x498 ^ x466 ;
  assign n2391 = x496 ^ x464 ;
  assign n2393 = x494 ^ x462 ;
  assign n2395 = x492 ^ x460 ;
  assign n2397 = x490 ^ x458 ;
  assign n2399 = x488 ^ x456 ;
  assign n2401 = x486 ^ x454 ;
  assign n2403 = x484 ^ x452 ;
  assign n2405 = x482 ^ x450 ;
  assign n2407 = x448 & ~x480 ;
  assign n2408 = n2407 ^ x482 ;
  assign n2406 = x482 ^ x449 ;
  assign n2409 = n2408 ^ n2406 ;
  assign n2410 = x481 ^ x449 ;
  assign n2411 = n2409 & ~n2410 ;
  assign n2412 = n2411 ^ n2406 ;
  assign n2413 = ~n2405 & n2412 ;
  assign n2414 = n2413 ^ x450 ;
  assign n2415 = n2414 ^ x484 ;
  assign n2404 = x484 ^ x451 ;
  assign n2416 = n2415 ^ n2404 ;
  assign n2417 = x483 ^ x451 ;
  assign n2418 = n2416 & ~n2417 ;
  assign n2419 = n2418 ^ n2404 ;
  assign n2420 = ~n2403 & n2419 ;
  assign n2421 = n2420 ^ x452 ;
  assign n2422 = n2421 ^ x486 ;
  assign n2402 = x486 ^ x453 ;
  assign n2423 = n2422 ^ n2402 ;
  assign n2424 = x485 ^ x453 ;
  assign n2425 = n2423 & ~n2424 ;
  assign n2426 = n2425 ^ n2402 ;
  assign n2427 = ~n2401 & n2426 ;
  assign n2428 = n2427 ^ x454 ;
  assign n2429 = n2428 ^ x488 ;
  assign n2400 = x488 ^ x455 ;
  assign n2430 = n2429 ^ n2400 ;
  assign n2431 = x487 ^ x455 ;
  assign n2432 = n2430 & ~n2431 ;
  assign n2433 = n2432 ^ n2400 ;
  assign n2434 = ~n2399 & n2433 ;
  assign n2435 = n2434 ^ x456 ;
  assign n2436 = n2435 ^ x490 ;
  assign n2398 = x490 ^ x457 ;
  assign n2437 = n2436 ^ n2398 ;
  assign n2438 = x489 ^ x457 ;
  assign n2439 = n2437 & ~n2438 ;
  assign n2440 = n2439 ^ n2398 ;
  assign n2441 = ~n2397 & n2440 ;
  assign n2442 = n2441 ^ x458 ;
  assign n2443 = n2442 ^ x492 ;
  assign n2396 = x492 ^ x459 ;
  assign n2444 = n2443 ^ n2396 ;
  assign n2445 = x491 ^ x459 ;
  assign n2446 = n2444 & ~n2445 ;
  assign n2447 = n2446 ^ n2396 ;
  assign n2448 = ~n2395 & n2447 ;
  assign n2449 = n2448 ^ x460 ;
  assign n2450 = n2449 ^ x494 ;
  assign n2394 = x494 ^ x461 ;
  assign n2451 = n2450 ^ n2394 ;
  assign n2452 = x493 ^ x461 ;
  assign n2453 = n2451 & ~n2452 ;
  assign n2454 = n2453 ^ n2394 ;
  assign n2455 = ~n2393 & n2454 ;
  assign n2456 = n2455 ^ x462 ;
  assign n2457 = n2456 ^ x496 ;
  assign n2392 = x496 ^ x463 ;
  assign n2458 = n2457 ^ n2392 ;
  assign n2459 = x495 ^ x463 ;
  assign n2460 = n2458 & ~n2459 ;
  assign n2461 = n2460 ^ n2392 ;
  assign n2462 = ~n2391 & n2461 ;
  assign n2463 = n2462 ^ x464 ;
  assign n2464 = n2463 ^ x498 ;
  assign n2390 = x498 ^ x465 ;
  assign n2465 = n2464 ^ n2390 ;
  assign n2466 = x497 ^ x465 ;
  assign n2467 = n2465 & ~n2466 ;
  assign n2468 = n2467 ^ n2390 ;
  assign n2469 = ~n2389 & n2468 ;
  assign n2470 = n2469 ^ x466 ;
  assign n2471 = n2470 ^ x500 ;
  assign n2388 = x500 ^ x467 ;
  assign n2472 = n2471 ^ n2388 ;
  assign n2473 = x499 ^ x467 ;
  assign n2474 = n2472 & ~n2473 ;
  assign n2475 = n2474 ^ n2388 ;
  assign n2476 = ~n2387 & n2475 ;
  assign n2477 = n2476 ^ x468 ;
  assign n2478 = n2477 ^ x502 ;
  assign n2386 = x502 ^ x469 ;
  assign n2479 = n2478 ^ n2386 ;
  assign n2480 = x501 ^ x469 ;
  assign n2481 = n2479 & ~n2480 ;
  assign n2482 = n2481 ^ n2386 ;
  assign n2483 = ~n2385 & n2482 ;
  assign n2484 = n2483 ^ x470 ;
  assign n2485 = n2484 ^ x504 ;
  assign n2384 = x504 ^ x471 ;
  assign n2486 = n2485 ^ n2384 ;
  assign n2487 = x503 ^ x471 ;
  assign n2488 = n2486 & ~n2487 ;
  assign n2489 = n2488 ^ n2384 ;
  assign n2490 = ~n2383 & n2489 ;
  assign n2491 = n2490 ^ x472 ;
  assign n2492 = n2491 ^ x506 ;
  assign n2382 = x506 ^ x473 ;
  assign n2493 = n2492 ^ n2382 ;
  assign n2494 = x505 ^ x473 ;
  assign n2495 = n2493 & ~n2494 ;
  assign n2496 = n2495 ^ n2382 ;
  assign n2497 = ~n2381 & n2496 ;
  assign n2498 = n2497 ^ x474 ;
  assign n2499 = n2498 ^ x508 ;
  assign n2380 = x508 ^ x475 ;
  assign n2500 = n2499 ^ n2380 ;
  assign n2501 = x507 ^ x475 ;
  assign n2502 = n2500 & ~n2501 ;
  assign n2503 = n2502 ^ n2380 ;
  assign n2504 = ~n2379 & n2503 ;
  assign n2505 = n2504 ^ x476 ;
  assign n2506 = n2505 ^ x510 ;
  assign n2378 = x510 ^ x477 ;
  assign n2507 = n2506 ^ n2378 ;
  assign n2508 = x509 ^ x477 ;
  assign n2509 = n2507 & ~n2508 ;
  assign n2510 = n2509 ^ n2378 ;
  assign n2511 = ~n2376 & n2510 ;
  assign n2512 = n2511 ^ x478 ;
  assign n2513 = n2512 ^ x511 ;
  assign n2514 = ~n2377 & n2513 ;
  assign n2515 = n2514 ^ x479 ;
  assign n2516 = n2376 & ~n2515 ;
  assign n2517 = n2516 ^ x478 ;
  assign n2660 = n2659 ^ n2517 ;
  assign n2661 = n517 ^ n516 ;
  assign n2664 = n2508 & ~n2515 ;
  assign n2665 = n2664 ^ x477 ;
  assign n2662 = n2650 & ~n2657 ;
  assign n2663 = n2662 ^ x413 ;
  assign n2666 = n2665 ^ n2663 ;
  assign n2669 = n2379 & ~n2515 ;
  assign n2670 = n2669 ^ x476 ;
  assign n2667 = n2521 & ~n2657 ;
  assign n2668 = n2667 ^ x412 ;
  assign n2671 = n2670 ^ n2668 ;
  assign n2674 = n2643 & ~n2657 ;
  assign n2675 = n2674 ^ x411 ;
  assign n2672 = n2501 & ~n2515 ;
  assign n2673 = n2672 ^ x475 ;
  assign n2676 = n2675 ^ n2673 ;
  assign n2679 = n2381 & ~n2515 ;
  assign n2680 = n2679 ^ x474 ;
  assign n2677 = n2523 & ~n2657 ;
  assign n2678 = n2677 ^ x410 ;
  assign n2681 = n2680 ^ n2678 ;
  assign n2684 = n2494 & ~n2515 ;
  assign n2685 = n2684 ^ x473 ;
  assign n2682 = n2636 & ~n2657 ;
  assign n2683 = n2682 ^ x409 ;
  assign n2686 = n2685 ^ n2683 ;
  assign n2689 = n2383 & ~n2515 ;
  assign n2690 = n2689 ^ x472 ;
  assign n2687 = n2525 & ~n2657 ;
  assign n2688 = n2687 ^ x408 ;
  assign n2691 = n2690 ^ n2688 ;
  assign n2694 = n2629 & ~n2657 ;
  assign n2695 = n2694 ^ x407 ;
  assign n2692 = n2487 & ~n2515 ;
  assign n2693 = n2692 ^ x471 ;
  assign n2696 = n2695 ^ n2693 ;
  assign n2699 = n2385 & ~n2515 ;
  assign n2700 = n2699 ^ x470 ;
  assign n2697 = n2527 & ~n2657 ;
  assign n2698 = n2697 ^ x406 ;
  assign n2701 = n2700 ^ n2698 ;
  assign n2704 = n2622 & ~n2657 ;
  assign n2705 = n2704 ^ x405 ;
  assign n2702 = n2480 & ~n2515 ;
  assign n2703 = n2702 ^ x469 ;
  assign n2706 = n2705 ^ n2703 ;
  assign n2709 = n2387 & ~n2515 ;
  assign n2710 = n2709 ^ x468 ;
  assign n2707 = n2529 & ~n2657 ;
  assign n2708 = n2707 ^ x404 ;
  assign n2711 = n2710 ^ n2708 ;
  assign n2714 = n2615 & ~n2657 ;
  assign n2715 = n2714 ^ x403 ;
  assign n2712 = n2473 & ~n2515 ;
  assign n2713 = n2712 ^ x467 ;
  assign n2716 = n2715 ^ n2713 ;
  assign n2719 = n2389 & ~n2515 ;
  assign n2720 = n2719 ^ x466 ;
  assign n2717 = n2531 & ~n2657 ;
  assign n2718 = n2717 ^ x402 ;
  assign n2721 = n2720 ^ n2718 ;
  assign n2724 = n2608 & ~n2657 ;
  assign n2725 = n2724 ^ x401 ;
  assign n2722 = n2466 & ~n2515 ;
  assign n2723 = n2722 ^ x465 ;
  assign n2726 = n2725 ^ n2723 ;
  assign n2729 = n2391 & ~n2515 ;
  assign n2730 = n2729 ^ x464 ;
  assign n2727 = n2533 & ~n2657 ;
  assign n2728 = n2727 ^ x400 ;
  assign n2731 = n2730 ^ n2728 ;
  assign n2734 = n2601 & ~n2657 ;
  assign n2735 = n2734 ^ x399 ;
  assign n2732 = n2459 & ~n2515 ;
  assign n2733 = n2732 ^ x463 ;
  assign n2736 = n2735 ^ n2733 ;
  assign n2739 = n2393 & ~n2515 ;
  assign n2740 = n2739 ^ x462 ;
  assign n2737 = n2535 & ~n2657 ;
  assign n2738 = n2737 ^ x398 ;
  assign n2741 = n2740 ^ n2738 ;
  assign n2744 = n2594 & ~n2657 ;
  assign n2745 = n2744 ^ x397 ;
  assign n2742 = n2452 & ~n2515 ;
  assign n2743 = n2742 ^ x461 ;
  assign n2746 = n2745 ^ n2743 ;
  assign n2749 = n2395 & ~n2515 ;
  assign n2750 = n2749 ^ x460 ;
  assign n2747 = n2537 & ~n2657 ;
  assign n2748 = n2747 ^ x396 ;
  assign n2751 = n2750 ^ n2748 ;
  assign n2754 = n2587 & ~n2657 ;
  assign n2755 = n2754 ^ x395 ;
  assign n2752 = n2445 & ~n2515 ;
  assign n2753 = n2752 ^ x459 ;
  assign n2756 = n2755 ^ n2753 ;
  assign n2759 = n2397 & ~n2515 ;
  assign n2760 = n2759 ^ x458 ;
  assign n2757 = n2539 & ~n2657 ;
  assign n2758 = n2757 ^ x394 ;
  assign n2761 = n2760 ^ n2758 ;
  assign n2764 = n2580 & ~n2657 ;
  assign n2765 = n2764 ^ x393 ;
  assign n2762 = n2438 & ~n2515 ;
  assign n2763 = n2762 ^ x457 ;
  assign n2766 = n2765 ^ n2763 ;
  assign n2769 = n2399 & ~n2515 ;
  assign n2770 = n2769 ^ x456 ;
  assign n2767 = n2541 & ~n2657 ;
  assign n2768 = n2767 ^ x392 ;
  assign n2771 = n2770 ^ n2768 ;
  assign n2774 = n2573 & ~n2657 ;
  assign n2775 = n2774 ^ x391 ;
  assign n2772 = n2431 & ~n2515 ;
  assign n2773 = n2772 ^ x455 ;
  assign n2776 = n2775 ^ n2773 ;
  assign n2779 = n2401 & ~n2515 ;
  assign n2780 = n2779 ^ x454 ;
  assign n2777 = n2543 & ~n2657 ;
  assign n2778 = n2777 ^ x390 ;
  assign n2781 = n2780 ^ n2778 ;
  assign n2784 = n2566 & ~n2657 ;
  assign n2785 = n2784 ^ x389 ;
  assign n2782 = n2424 & ~n2515 ;
  assign n2783 = n2782 ^ x453 ;
  assign n2786 = n2785 ^ n2783 ;
  assign n2789 = n2403 & ~n2515 ;
  assign n2790 = n2789 ^ x452 ;
  assign n2787 = n2545 & ~n2657 ;
  assign n2788 = n2787 ^ x388 ;
  assign n2791 = n2790 ^ n2788 ;
  assign n2794 = n2559 & ~n2657 ;
  assign n2795 = n2794 ^ x387 ;
  assign n2792 = n2417 & ~n2515 ;
  assign n2793 = n2792 ^ x451 ;
  assign n2796 = n2795 ^ n2793 ;
  assign n2799 = n2547 & ~n2657 ;
  assign n2800 = n2799 ^ x386 ;
  assign n2797 = n2405 & ~n2515 ;
  assign n2798 = n2797 ^ x450 ;
  assign n2801 = n2800 ^ n2798 ;
  assign n2804 = n2410 & ~n2515 ;
  assign n2805 = n2804 ^ x449 ;
  assign n2802 = n2552 & ~n2657 ;
  assign n2803 = n2802 ^ x385 ;
  assign n2806 = n2805 ^ n2803 ;
  assign n2807 = x480 ^ x448 ;
  assign n2808 = ~n2515 & n2807 ;
  assign n2809 = n2808 ^ x448 ;
  assign n2810 = x416 ^ x384 ;
  assign n2811 = ~n2657 & n2810 ;
  assign n2812 = n2811 ^ x384 ;
  assign n2813 = ~n2809 & n2812 ;
  assign n2814 = n2813 ^ n2805 ;
  assign n2815 = ~n2806 & ~n2814 ;
  assign n2816 = n2815 ^ n2805 ;
  assign n2817 = n2816 ^ n2800 ;
  assign n2818 = ~n2801 & ~n2817 ;
  assign n2819 = n2818 ^ n2800 ;
  assign n2820 = n2819 ^ n2795 ;
  assign n2821 = ~n2796 & n2820 ;
  assign n2822 = n2821 ^ n2795 ;
  assign n2823 = n2822 ^ n2788 ;
  assign n2824 = ~n2791 & n2823 ;
  assign n2825 = n2824 ^ n2788 ;
  assign n2826 = n2825 ^ n2785 ;
  assign n2827 = ~n2786 & n2826 ;
  assign n2828 = n2827 ^ n2785 ;
  assign n2829 = n2828 ^ n2778 ;
  assign n2830 = ~n2781 & n2829 ;
  assign n2831 = n2830 ^ n2778 ;
  assign n2832 = n2831 ^ n2775 ;
  assign n2833 = ~n2776 & n2832 ;
  assign n2834 = n2833 ^ n2775 ;
  assign n2835 = n2834 ^ n2768 ;
  assign n2836 = ~n2771 & n2835 ;
  assign n2837 = n2836 ^ n2768 ;
  assign n2838 = n2837 ^ n2765 ;
  assign n2839 = ~n2766 & n2838 ;
  assign n2840 = n2839 ^ n2765 ;
  assign n2841 = n2840 ^ n2758 ;
  assign n2842 = ~n2761 & n2841 ;
  assign n2843 = n2842 ^ n2758 ;
  assign n2844 = n2843 ^ n2755 ;
  assign n2845 = ~n2756 & n2844 ;
  assign n2846 = n2845 ^ n2755 ;
  assign n2847 = n2846 ^ n2748 ;
  assign n2848 = ~n2751 & n2847 ;
  assign n2849 = n2848 ^ n2748 ;
  assign n2850 = n2849 ^ n2745 ;
  assign n2851 = ~n2746 & n2850 ;
  assign n2852 = n2851 ^ n2745 ;
  assign n2853 = n2852 ^ n2738 ;
  assign n2854 = ~n2741 & n2853 ;
  assign n2855 = n2854 ^ n2738 ;
  assign n2856 = n2855 ^ n2735 ;
  assign n2857 = ~n2736 & n2856 ;
  assign n2858 = n2857 ^ n2735 ;
  assign n2859 = n2858 ^ n2728 ;
  assign n2860 = ~n2731 & n2859 ;
  assign n2861 = n2860 ^ n2728 ;
  assign n2862 = n2861 ^ n2725 ;
  assign n2863 = ~n2726 & n2862 ;
  assign n2864 = n2863 ^ n2725 ;
  assign n2865 = n2864 ^ n2718 ;
  assign n2866 = ~n2721 & n2865 ;
  assign n2867 = n2866 ^ n2718 ;
  assign n2868 = n2867 ^ n2715 ;
  assign n2869 = ~n2716 & n2868 ;
  assign n2870 = n2869 ^ n2715 ;
  assign n2871 = n2870 ^ n2708 ;
  assign n2872 = ~n2711 & n2871 ;
  assign n2873 = n2872 ^ n2708 ;
  assign n2874 = n2873 ^ n2705 ;
  assign n2875 = ~n2706 & n2874 ;
  assign n2876 = n2875 ^ n2705 ;
  assign n2877 = n2876 ^ n2698 ;
  assign n2878 = ~n2701 & n2877 ;
  assign n2879 = n2878 ^ n2698 ;
  assign n2880 = n2879 ^ n2695 ;
  assign n2881 = ~n2696 & n2880 ;
  assign n2882 = n2881 ^ n2695 ;
  assign n2883 = n2882 ^ n2688 ;
  assign n2884 = ~n2691 & n2883 ;
  assign n2885 = n2884 ^ n2688 ;
  assign n2886 = n2885 ^ n2685 ;
  assign n2887 = ~n2686 & ~n2886 ;
  assign n2888 = n2887 ^ n2685 ;
  assign n2889 = n2888 ^ n2678 ;
  assign n2890 = ~n2681 & ~n2889 ;
  assign n2891 = n2890 ^ n2678 ;
  assign n2892 = n2891 ^ n2675 ;
  assign n2893 = ~n2676 & n2892 ;
  assign n2894 = n2893 ^ n2675 ;
  assign n2895 = n2894 ^ n2670 ;
  assign n2896 = ~n2671 & ~n2895 ;
  assign n2897 = n2896 ^ n2670 ;
  assign n2898 = n2897 ^ n2665 ;
  assign n2899 = ~n2666 & ~n2898 ;
  assign n2900 = n2899 ^ n2663 ;
  assign n2901 = n2900 ^ n2659 ;
  assign n2902 = ~n2660 & ~n2901 ;
  assign n2903 = n2902 ^ n2517 ;
  assign n2904 = n2903 ^ n517 ;
  assign n2905 = ~n2661 & n2904 ;
  assign n2906 = n2905 ^ n516 ;
  assign n2907 = n2660 & ~n2906 ;
  assign n2908 = n2907 ^ n2517 ;
  assign n1985 = x382 ^ x350 ;
  assign n1986 = x383 ^ x351 ;
  assign n1988 = x380 ^ x348 ;
  assign n1990 = x378 ^ x346 ;
  assign n1992 = x376 ^ x344 ;
  assign n1994 = x374 ^ x342 ;
  assign n1996 = x372 ^ x340 ;
  assign n1998 = x370 ^ x338 ;
  assign n2000 = x368 ^ x336 ;
  assign n2002 = x366 ^ x334 ;
  assign n2004 = x364 ^ x332 ;
  assign n2006 = x362 ^ x330 ;
  assign n2008 = x360 ^ x328 ;
  assign n2010 = x358 ^ x326 ;
  assign n2012 = x356 ^ x324 ;
  assign n2014 = x354 ^ x322 ;
  assign n2016 = x320 & ~x352 ;
  assign n2017 = n2016 ^ x354 ;
  assign n2015 = x354 ^ x321 ;
  assign n2018 = n2017 ^ n2015 ;
  assign n2019 = x353 ^ x321 ;
  assign n2020 = n2018 & ~n2019 ;
  assign n2021 = n2020 ^ n2015 ;
  assign n2022 = ~n2014 & n2021 ;
  assign n2023 = n2022 ^ x322 ;
  assign n2024 = n2023 ^ x356 ;
  assign n2013 = x356 ^ x323 ;
  assign n2025 = n2024 ^ n2013 ;
  assign n2026 = x355 ^ x323 ;
  assign n2027 = n2025 & ~n2026 ;
  assign n2028 = n2027 ^ n2013 ;
  assign n2029 = ~n2012 & n2028 ;
  assign n2030 = n2029 ^ x324 ;
  assign n2031 = n2030 ^ x358 ;
  assign n2011 = x358 ^ x325 ;
  assign n2032 = n2031 ^ n2011 ;
  assign n2033 = x357 ^ x325 ;
  assign n2034 = n2032 & ~n2033 ;
  assign n2035 = n2034 ^ n2011 ;
  assign n2036 = ~n2010 & n2035 ;
  assign n2037 = n2036 ^ x326 ;
  assign n2038 = n2037 ^ x360 ;
  assign n2009 = x360 ^ x327 ;
  assign n2039 = n2038 ^ n2009 ;
  assign n2040 = x359 ^ x327 ;
  assign n2041 = n2039 & ~n2040 ;
  assign n2042 = n2041 ^ n2009 ;
  assign n2043 = ~n2008 & n2042 ;
  assign n2044 = n2043 ^ x328 ;
  assign n2045 = n2044 ^ x362 ;
  assign n2007 = x362 ^ x329 ;
  assign n2046 = n2045 ^ n2007 ;
  assign n2047 = x361 ^ x329 ;
  assign n2048 = n2046 & ~n2047 ;
  assign n2049 = n2048 ^ n2007 ;
  assign n2050 = ~n2006 & n2049 ;
  assign n2051 = n2050 ^ x330 ;
  assign n2052 = n2051 ^ x364 ;
  assign n2005 = x364 ^ x331 ;
  assign n2053 = n2052 ^ n2005 ;
  assign n2054 = x363 ^ x331 ;
  assign n2055 = n2053 & ~n2054 ;
  assign n2056 = n2055 ^ n2005 ;
  assign n2057 = ~n2004 & n2056 ;
  assign n2058 = n2057 ^ x332 ;
  assign n2059 = n2058 ^ x366 ;
  assign n2003 = x366 ^ x333 ;
  assign n2060 = n2059 ^ n2003 ;
  assign n2061 = x365 ^ x333 ;
  assign n2062 = n2060 & ~n2061 ;
  assign n2063 = n2062 ^ n2003 ;
  assign n2064 = ~n2002 & n2063 ;
  assign n2065 = n2064 ^ x334 ;
  assign n2066 = n2065 ^ x368 ;
  assign n2001 = x368 ^ x335 ;
  assign n2067 = n2066 ^ n2001 ;
  assign n2068 = x367 ^ x335 ;
  assign n2069 = n2067 & ~n2068 ;
  assign n2070 = n2069 ^ n2001 ;
  assign n2071 = ~n2000 & n2070 ;
  assign n2072 = n2071 ^ x336 ;
  assign n2073 = n2072 ^ x370 ;
  assign n1999 = x370 ^ x337 ;
  assign n2074 = n2073 ^ n1999 ;
  assign n2075 = x369 ^ x337 ;
  assign n2076 = n2074 & ~n2075 ;
  assign n2077 = n2076 ^ n1999 ;
  assign n2078 = ~n1998 & n2077 ;
  assign n2079 = n2078 ^ x338 ;
  assign n2080 = n2079 ^ x372 ;
  assign n1997 = x372 ^ x339 ;
  assign n2081 = n2080 ^ n1997 ;
  assign n2082 = x371 ^ x339 ;
  assign n2083 = n2081 & ~n2082 ;
  assign n2084 = n2083 ^ n1997 ;
  assign n2085 = ~n1996 & n2084 ;
  assign n2086 = n2085 ^ x340 ;
  assign n2087 = n2086 ^ x374 ;
  assign n1995 = x374 ^ x341 ;
  assign n2088 = n2087 ^ n1995 ;
  assign n2089 = x373 ^ x341 ;
  assign n2090 = n2088 & ~n2089 ;
  assign n2091 = n2090 ^ n1995 ;
  assign n2092 = ~n1994 & n2091 ;
  assign n2093 = n2092 ^ x342 ;
  assign n2094 = n2093 ^ x376 ;
  assign n1993 = x376 ^ x343 ;
  assign n2095 = n2094 ^ n1993 ;
  assign n2096 = x375 ^ x343 ;
  assign n2097 = n2095 & ~n2096 ;
  assign n2098 = n2097 ^ n1993 ;
  assign n2099 = ~n1992 & n2098 ;
  assign n2100 = n2099 ^ x344 ;
  assign n2101 = n2100 ^ x378 ;
  assign n1991 = x378 ^ x345 ;
  assign n2102 = n2101 ^ n1991 ;
  assign n2103 = x377 ^ x345 ;
  assign n2104 = n2102 & ~n2103 ;
  assign n2105 = n2104 ^ n1991 ;
  assign n2106 = ~n1990 & n2105 ;
  assign n2107 = n2106 ^ x346 ;
  assign n2108 = n2107 ^ x380 ;
  assign n1989 = x380 ^ x347 ;
  assign n2109 = n2108 ^ n1989 ;
  assign n2110 = x379 ^ x347 ;
  assign n2111 = n2109 & ~n2110 ;
  assign n2112 = n2111 ^ n1989 ;
  assign n2113 = ~n1988 & n2112 ;
  assign n2114 = n2113 ^ x348 ;
  assign n2115 = n2114 ^ x382 ;
  assign n1987 = x382 ^ x349 ;
  assign n2116 = n2115 ^ n1987 ;
  assign n2117 = x381 ^ x349 ;
  assign n2118 = n2116 & ~n2117 ;
  assign n2119 = n2118 ^ n1987 ;
  assign n2120 = ~n1985 & n2119 ;
  assign n2121 = n2120 ^ x350 ;
  assign n2122 = n2121 ^ x383 ;
  assign n2123 = ~n1986 & n2122 ;
  assign n2124 = n2123 ^ x351 ;
  assign n2125 = n1985 & ~n2124 ;
  assign n2126 = n2125 ^ x350 ;
  assign n1843 = x318 ^ x286 ;
  assign n1844 = x319 ^ x287 ;
  assign n1846 = x316 ^ x284 ;
  assign n1848 = x314 ^ x282 ;
  assign n1850 = x312 ^ x280 ;
  assign n1852 = x310 ^ x278 ;
  assign n1854 = x308 ^ x276 ;
  assign n1856 = x306 ^ x274 ;
  assign n1858 = x304 ^ x272 ;
  assign n1860 = x302 ^ x270 ;
  assign n1862 = x300 ^ x268 ;
  assign n1864 = x298 ^ x266 ;
  assign n1866 = x296 ^ x264 ;
  assign n1868 = x294 ^ x262 ;
  assign n1870 = x292 ^ x260 ;
  assign n1872 = x290 ^ x258 ;
  assign n1874 = x256 & ~x288 ;
  assign n1875 = n1874 ^ x290 ;
  assign n1873 = x290 ^ x257 ;
  assign n1876 = n1875 ^ n1873 ;
  assign n1877 = x289 ^ x257 ;
  assign n1878 = n1876 & ~n1877 ;
  assign n1879 = n1878 ^ n1873 ;
  assign n1880 = ~n1872 & n1879 ;
  assign n1881 = n1880 ^ x258 ;
  assign n1882 = n1881 ^ x292 ;
  assign n1871 = x292 ^ x259 ;
  assign n1883 = n1882 ^ n1871 ;
  assign n1884 = x291 ^ x259 ;
  assign n1885 = n1883 & ~n1884 ;
  assign n1886 = n1885 ^ n1871 ;
  assign n1887 = ~n1870 & n1886 ;
  assign n1888 = n1887 ^ x260 ;
  assign n1889 = n1888 ^ x294 ;
  assign n1869 = x294 ^ x261 ;
  assign n1890 = n1889 ^ n1869 ;
  assign n1891 = x293 ^ x261 ;
  assign n1892 = n1890 & ~n1891 ;
  assign n1893 = n1892 ^ n1869 ;
  assign n1894 = ~n1868 & n1893 ;
  assign n1895 = n1894 ^ x262 ;
  assign n1896 = n1895 ^ x296 ;
  assign n1867 = x296 ^ x263 ;
  assign n1897 = n1896 ^ n1867 ;
  assign n1898 = x295 ^ x263 ;
  assign n1899 = n1897 & ~n1898 ;
  assign n1900 = n1899 ^ n1867 ;
  assign n1901 = ~n1866 & n1900 ;
  assign n1902 = n1901 ^ x264 ;
  assign n1903 = n1902 ^ x298 ;
  assign n1865 = x298 ^ x265 ;
  assign n1904 = n1903 ^ n1865 ;
  assign n1905 = x297 ^ x265 ;
  assign n1906 = n1904 & ~n1905 ;
  assign n1907 = n1906 ^ n1865 ;
  assign n1908 = ~n1864 & n1907 ;
  assign n1909 = n1908 ^ x266 ;
  assign n1910 = n1909 ^ x300 ;
  assign n1863 = x300 ^ x267 ;
  assign n1911 = n1910 ^ n1863 ;
  assign n1912 = x299 ^ x267 ;
  assign n1913 = n1911 & ~n1912 ;
  assign n1914 = n1913 ^ n1863 ;
  assign n1915 = ~n1862 & n1914 ;
  assign n1916 = n1915 ^ x268 ;
  assign n1917 = n1916 ^ x302 ;
  assign n1861 = x302 ^ x269 ;
  assign n1918 = n1917 ^ n1861 ;
  assign n1919 = x301 ^ x269 ;
  assign n1920 = n1918 & ~n1919 ;
  assign n1921 = n1920 ^ n1861 ;
  assign n1922 = ~n1860 & n1921 ;
  assign n1923 = n1922 ^ x270 ;
  assign n1924 = n1923 ^ x304 ;
  assign n1859 = x304 ^ x271 ;
  assign n1925 = n1924 ^ n1859 ;
  assign n1926 = x303 ^ x271 ;
  assign n1927 = n1925 & ~n1926 ;
  assign n1928 = n1927 ^ n1859 ;
  assign n1929 = ~n1858 & n1928 ;
  assign n1930 = n1929 ^ x272 ;
  assign n1931 = n1930 ^ x306 ;
  assign n1857 = x306 ^ x273 ;
  assign n1932 = n1931 ^ n1857 ;
  assign n1933 = x305 ^ x273 ;
  assign n1934 = n1932 & ~n1933 ;
  assign n1935 = n1934 ^ n1857 ;
  assign n1936 = ~n1856 & n1935 ;
  assign n1937 = n1936 ^ x274 ;
  assign n1938 = n1937 ^ x308 ;
  assign n1855 = x308 ^ x275 ;
  assign n1939 = n1938 ^ n1855 ;
  assign n1940 = x307 ^ x275 ;
  assign n1941 = n1939 & ~n1940 ;
  assign n1942 = n1941 ^ n1855 ;
  assign n1943 = ~n1854 & n1942 ;
  assign n1944 = n1943 ^ x276 ;
  assign n1945 = n1944 ^ x310 ;
  assign n1853 = x310 ^ x277 ;
  assign n1946 = n1945 ^ n1853 ;
  assign n1947 = x309 ^ x277 ;
  assign n1948 = n1946 & ~n1947 ;
  assign n1949 = n1948 ^ n1853 ;
  assign n1950 = ~n1852 & n1949 ;
  assign n1951 = n1950 ^ x278 ;
  assign n1952 = n1951 ^ x312 ;
  assign n1851 = x312 ^ x279 ;
  assign n1953 = n1952 ^ n1851 ;
  assign n1954 = x311 ^ x279 ;
  assign n1955 = n1953 & ~n1954 ;
  assign n1956 = n1955 ^ n1851 ;
  assign n1957 = ~n1850 & n1956 ;
  assign n1958 = n1957 ^ x280 ;
  assign n1959 = n1958 ^ x314 ;
  assign n1849 = x314 ^ x281 ;
  assign n1960 = n1959 ^ n1849 ;
  assign n1961 = x313 ^ x281 ;
  assign n1962 = n1960 & ~n1961 ;
  assign n1963 = n1962 ^ n1849 ;
  assign n1964 = ~n1848 & n1963 ;
  assign n1965 = n1964 ^ x282 ;
  assign n1966 = n1965 ^ x316 ;
  assign n1847 = x316 ^ x283 ;
  assign n1967 = n1966 ^ n1847 ;
  assign n1968 = x315 ^ x283 ;
  assign n1969 = n1967 & ~n1968 ;
  assign n1970 = n1969 ^ n1847 ;
  assign n1971 = ~n1846 & n1970 ;
  assign n1972 = n1971 ^ x284 ;
  assign n1973 = n1972 ^ x318 ;
  assign n1845 = x318 ^ x285 ;
  assign n1974 = n1973 ^ n1845 ;
  assign n1975 = x317 ^ x285 ;
  assign n1976 = n1974 & ~n1975 ;
  assign n1977 = n1976 ^ n1845 ;
  assign n1978 = ~n1843 & n1977 ;
  assign n1979 = n1978 ^ x286 ;
  assign n1980 = n1979 ^ x319 ;
  assign n1981 = ~n1844 & n1980 ;
  assign n1982 = n1981 ^ x287 ;
  assign n1983 = n1843 & ~n1982 ;
  assign n1984 = n1983 ^ x286 ;
  assign n2127 = n2126 ^ n1984 ;
  assign n2128 = n514 ^ n513 ;
  assign n2131 = n2117 & ~n2124 ;
  assign n2132 = n2131 ^ x349 ;
  assign n2129 = n1975 & ~n1982 ;
  assign n2130 = n2129 ^ x285 ;
  assign n2133 = n2132 ^ n2130 ;
  assign n2136 = n1988 & ~n2124 ;
  assign n2137 = n2136 ^ x348 ;
  assign n2134 = n1846 & ~n1982 ;
  assign n2135 = n2134 ^ x284 ;
  assign n2138 = n2137 ^ n2135 ;
  assign n2141 = n1968 & ~n1982 ;
  assign n2142 = n2141 ^ x283 ;
  assign n2139 = n2110 & ~n2124 ;
  assign n2140 = n2139 ^ x347 ;
  assign n2143 = n2142 ^ n2140 ;
  assign n2146 = n1990 & ~n2124 ;
  assign n2147 = n2146 ^ x346 ;
  assign n2144 = n1848 & ~n1982 ;
  assign n2145 = n2144 ^ x282 ;
  assign n2148 = n2147 ^ n2145 ;
  assign n2151 = n1961 & ~n1982 ;
  assign n2152 = n2151 ^ x281 ;
  assign n2149 = n2103 & ~n2124 ;
  assign n2150 = n2149 ^ x345 ;
  assign n2153 = n2152 ^ n2150 ;
  assign n2156 = n1992 & ~n2124 ;
  assign n2157 = n2156 ^ x344 ;
  assign n2154 = n1850 & ~n1982 ;
  assign n2155 = n2154 ^ x280 ;
  assign n2158 = n2157 ^ n2155 ;
  assign n2161 = n1954 & ~n1982 ;
  assign n2162 = n2161 ^ x279 ;
  assign n2159 = n2096 & ~n2124 ;
  assign n2160 = n2159 ^ x343 ;
  assign n2163 = n2162 ^ n2160 ;
  assign n2166 = n1994 & ~n2124 ;
  assign n2167 = n2166 ^ x342 ;
  assign n2164 = n1852 & ~n1982 ;
  assign n2165 = n2164 ^ x278 ;
  assign n2168 = n2167 ^ n2165 ;
  assign n2171 = n1947 & ~n1982 ;
  assign n2172 = n2171 ^ x277 ;
  assign n2169 = n2089 & ~n2124 ;
  assign n2170 = n2169 ^ x341 ;
  assign n2173 = n2172 ^ n2170 ;
  assign n2176 = n1996 & ~n2124 ;
  assign n2177 = n2176 ^ x340 ;
  assign n2174 = n1854 & ~n1982 ;
  assign n2175 = n2174 ^ x276 ;
  assign n2178 = n2177 ^ n2175 ;
  assign n2181 = n1940 & ~n1982 ;
  assign n2182 = n2181 ^ x275 ;
  assign n2179 = n2082 & ~n2124 ;
  assign n2180 = n2179 ^ x339 ;
  assign n2183 = n2182 ^ n2180 ;
  assign n2186 = n1998 & ~n2124 ;
  assign n2187 = n2186 ^ x338 ;
  assign n2184 = n1856 & ~n1982 ;
  assign n2185 = n2184 ^ x274 ;
  assign n2188 = n2187 ^ n2185 ;
  assign n2191 = n1933 & ~n1982 ;
  assign n2192 = n2191 ^ x273 ;
  assign n2189 = n2075 & ~n2124 ;
  assign n2190 = n2189 ^ x337 ;
  assign n2193 = n2192 ^ n2190 ;
  assign n2196 = n2000 & ~n2124 ;
  assign n2197 = n2196 ^ x336 ;
  assign n2194 = n1858 & ~n1982 ;
  assign n2195 = n2194 ^ x272 ;
  assign n2198 = n2197 ^ n2195 ;
  assign n2201 = n1926 & ~n1982 ;
  assign n2202 = n2201 ^ x271 ;
  assign n2199 = n2068 & ~n2124 ;
  assign n2200 = n2199 ^ x335 ;
  assign n2203 = n2202 ^ n2200 ;
  assign n2206 = n2002 & ~n2124 ;
  assign n2207 = n2206 ^ x334 ;
  assign n2204 = n1860 & ~n1982 ;
  assign n2205 = n2204 ^ x270 ;
  assign n2208 = n2207 ^ n2205 ;
  assign n2211 = n1919 & ~n1982 ;
  assign n2212 = n2211 ^ x269 ;
  assign n2209 = n2061 & ~n2124 ;
  assign n2210 = n2209 ^ x333 ;
  assign n2213 = n2212 ^ n2210 ;
  assign n2216 = n2004 & ~n2124 ;
  assign n2217 = n2216 ^ x332 ;
  assign n2214 = n1862 & ~n1982 ;
  assign n2215 = n2214 ^ x268 ;
  assign n2218 = n2217 ^ n2215 ;
  assign n2221 = n1912 & ~n1982 ;
  assign n2222 = n2221 ^ x267 ;
  assign n2219 = n2054 & ~n2124 ;
  assign n2220 = n2219 ^ x331 ;
  assign n2223 = n2222 ^ n2220 ;
  assign n2226 = n2006 & ~n2124 ;
  assign n2227 = n2226 ^ x330 ;
  assign n2224 = n1864 & ~n1982 ;
  assign n2225 = n2224 ^ x266 ;
  assign n2228 = n2227 ^ n2225 ;
  assign n2231 = n1905 & ~n1982 ;
  assign n2232 = n2231 ^ x265 ;
  assign n2229 = n2047 & ~n2124 ;
  assign n2230 = n2229 ^ x329 ;
  assign n2233 = n2232 ^ n2230 ;
  assign n2236 = n2008 & ~n2124 ;
  assign n2237 = n2236 ^ x328 ;
  assign n2234 = n1866 & ~n1982 ;
  assign n2235 = n2234 ^ x264 ;
  assign n2238 = n2237 ^ n2235 ;
  assign n2241 = n1898 & ~n1982 ;
  assign n2242 = n2241 ^ x263 ;
  assign n2239 = n2040 & ~n2124 ;
  assign n2240 = n2239 ^ x327 ;
  assign n2243 = n2242 ^ n2240 ;
  assign n2246 = n1868 & ~n1982 ;
  assign n2247 = n2246 ^ x262 ;
  assign n2244 = n2010 & ~n2124 ;
  assign n2245 = n2244 ^ x326 ;
  assign n2248 = n2247 ^ n2245 ;
  assign n2251 = n1891 & ~n1982 ;
  assign n2252 = n2251 ^ x261 ;
  assign n2249 = n2033 & ~n2124 ;
  assign n2250 = n2249 ^ x325 ;
  assign n2253 = n2252 ^ n2250 ;
  assign n2256 = n2012 & ~n2124 ;
  assign n2257 = n2256 ^ x324 ;
  assign n2254 = n1870 & ~n1982 ;
  assign n2255 = n2254 ^ x260 ;
  assign n2258 = n2257 ^ n2255 ;
  assign n2261 = n1884 & ~n1982 ;
  assign n2262 = n2261 ^ x259 ;
  assign n2259 = n2026 & ~n2124 ;
  assign n2260 = n2259 ^ x323 ;
  assign n2263 = n2262 ^ n2260 ;
  assign n2266 = n1872 & ~n1982 ;
  assign n2267 = n2266 ^ x258 ;
  assign n2264 = n2014 & ~n2124 ;
  assign n2265 = n2264 ^ x322 ;
  assign n2268 = n2267 ^ n2265 ;
  assign n2271 = n2019 & ~n2124 ;
  assign n2272 = n2271 ^ x321 ;
  assign n2269 = n1877 & ~n1982 ;
  assign n2270 = n2269 ^ x257 ;
  assign n2273 = n2272 ^ n2270 ;
  assign n2274 = x352 ^ x320 ;
  assign n2275 = ~n2124 & n2274 ;
  assign n2276 = n2275 ^ x320 ;
  assign n2277 = x288 ^ x256 ;
  assign n2278 = ~n1982 & n2277 ;
  assign n2279 = n2278 ^ x256 ;
  assign n2280 = ~n2276 & n2279 ;
  assign n2281 = n2280 ^ n2272 ;
  assign n2282 = ~n2273 & ~n2281 ;
  assign n2283 = n2282 ^ n2272 ;
  assign n2284 = n2283 ^ n2267 ;
  assign n2285 = ~n2268 & ~n2284 ;
  assign n2286 = n2285 ^ n2267 ;
  assign n2287 = n2286 ^ n2262 ;
  assign n2288 = ~n2263 & n2287 ;
  assign n2289 = n2288 ^ n2262 ;
  assign n2290 = n2289 ^ n2255 ;
  assign n2291 = ~n2258 & n2290 ;
  assign n2292 = n2291 ^ n2255 ;
  assign n2293 = n2292 ^ n2252 ;
  assign n2294 = ~n2253 & n2293 ;
  assign n2295 = n2294 ^ n2252 ;
  assign n2296 = n2295 ^ n2245 ;
  assign n2297 = ~n2248 & ~n2296 ;
  assign n2298 = n2297 ^ n2245 ;
  assign n2299 = n2298 ^ n2242 ;
  assign n2300 = ~n2243 & ~n2299 ;
  assign n2301 = n2300 ^ n2242 ;
  assign n2302 = n2301 ^ n2235 ;
  assign n2303 = ~n2238 & n2302 ;
  assign n2304 = n2303 ^ n2235 ;
  assign n2305 = n2304 ^ n2232 ;
  assign n2306 = ~n2233 & n2305 ;
  assign n2307 = n2306 ^ n2232 ;
  assign n2308 = n2307 ^ n2225 ;
  assign n2309 = ~n2228 & n2308 ;
  assign n2310 = n2309 ^ n2225 ;
  assign n2311 = n2310 ^ n2222 ;
  assign n2312 = ~n2223 & n2311 ;
  assign n2313 = n2312 ^ n2222 ;
  assign n2314 = n2313 ^ n2215 ;
  assign n2315 = ~n2218 & n2314 ;
  assign n2316 = n2315 ^ n2215 ;
  assign n2317 = n2316 ^ n2212 ;
  assign n2318 = ~n2213 & n2317 ;
  assign n2319 = n2318 ^ n2212 ;
  assign n2320 = n2319 ^ n2205 ;
  assign n2321 = ~n2208 & n2320 ;
  assign n2322 = n2321 ^ n2205 ;
  assign n2323 = n2322 ^ n2202 ;
  assign n2324 = ~n2203 & n2323 ;
  assign n2325 = n2324 ^ n2202 ;
  assign n2326 = n2325 ^ n2195 ;
  assign n2327 = ~n2198 & n2326 ;
  assign n2328 = n2327 ^ n2195 ;
  assign n2329 = n2328 ^ n2192 ;
  assign n2330 = ~n2193 & n2329 ;
  assign n2331 = n2330 ^ n2192 ;
  assign n2332 = n2331 ^ n2185 ;
  assign n2333 = ~n2188 & n2332 ;
  assign n2334 = n2333 ^ n2185 ;
  assign n2335 = n2334 ^ n2182 ;
  assign n2336 = ~n2183 & n2335 ;
  assign n2337 = n2336 ^ n2182 ;
  assign n2338 = n2337 ^ n2175 ;
  assign n2339 = ~n2178 & n2338 ;
  assign n2340 = n2339 ^ n2175 ;
  assign n2341 = n2340 ^ n2172 ;
  assign n2342 = ~n2173 & n2341 ;
  assign n2343 = n2342 ^ n2172 ;
  assign n2344 = n2343 ^ n2165 ;
  assign n2345 = ~n2168 & n2344 ;
  assign n2346 = n2345 ^ n2165 ;
  assign n2347 = n2346 ^ n2162 ;
  assign n2348 = ~n2163 & n2347 ;
  assign n2349 = n2348 ^ n2162 ;
  assign n2350 = n2349 ^ n2155 ;
  assign n2351 = ~n2158 & n2350 ;
  assign n2352 = n2351 ^ n2155 ;
  assign n2353 = n2352 ^ n2152 ;
  assign n2354 = ~n2153 & n2353 ;
  assign n2355 = n2354 ^ n2152 ;
  assign n2356 = n2355 ^ n2145 ;
  assign n2357 = ~n2148 & n2356 ;
  assign n2358 = n2357 ^ n2145 ;
  assign n2359 = n2358 ^ n2142 ;
  assign n2360 = ~n2143 & n2359 ;
  assign n2361 = n2360 ^ n2142 ;
  assign n2362 = n2361 ^ n2137 ;
  assign n2363 = ~n2138 & ~n2362 ;
  assign n2364 = n2363 ^ n2137 ;
  assign n2365 = n2364 ^ n2132 ;
  assign n2366 = ~n2133 & ~n2365 ;
  assign n2367 = n2366 ^ n2130 ;
  assign n2368 = n2367 ^ n2126 ;
  assign n2369 = ~n2127 & n2368 ;
  assign n2370 = n2369 ^ n1984 ;
  assign n2371 = n2370 ^ n514 ;
  assign n2372 = ~n2128 & ~n2371 ;
  assign n2373 = n2372 ^ n513 ;
  assign n2374 = n2127 & n2373 ;
  assign n2375 = n2374 ^ n1984 ;
  assign n2909 = n2908 ^ n2375 ;
  assign n2910 = n518 ^ n515 ;
  assign n2913 = n2666 & ~n2906 ;
  assign n2914 = n2913 ^ n2665 ;
  assign n2911 = n2133 & ~n2373 ;
  assign n2912 = n2911 ^ n2132 ;
  assign n2915 = n2914 ^ n2912 ;
  assign n2918 = n2138 & ~n2373 ;
  assign n2919 = n2918 ^ n2137 ;
  assign n2916 = n2671 & ~n2906 ;
  assign n2917 = n2916 ^ n2670 ;
  assign n2920 = n2919 ^ n2917 ;
  assign n2923 = n2143 & n2373 ;
  assign n2924 = n2923 ^ n2142 ;
  assign n2921 = n2676 & n2906 ;
  assign n2922 = n2921 ^ n2675 ;
  assign n2925 = n2924 ^ n2922 ;
  assign n2928 = n2148 & n2373 ;
  assign n2929 = n2928 ^ n2145 ;
  assign n2926 = n2681 & n2906 ;
  assign n2927 = n2926 ^ n2678 ;
  assign n2930 = n2929 ^ n2927 ;
  assign n2933 = n2153 & ~n2373 ;
  assign n2934 = n2933 ^ n2150 ;
  assign n2931 = n2686 & n2906 ;
  assign n2932 = n2931 ^ n2683 ;
  assign n2935 = n2934 ^ n2932 ;
  assign n2938 = n2691 & ~n2906 ;
  assign n2939 = n2938 ^ n2690 ;
  assign n2936 = n2158 & ~n2373 ;
  assign n2937 = n2936 ^ n2157 ;
  assign n2940 = n2939 ^ n2937 ;
  assign n2943 = n2163 & n2373 ;
  assign n2944 = n2943 ^ n2162 ;
  assign n2941 = n2696 & n2906 ;
  assign n2942 = n2941 ^ n2695 ;
  assign n2945 = n2944 ^ n2942 ;
  assign n2948 = n2168 & n2373 ;
  assign n2949 = n2948 ^ n2165 ;
  assign n2946 = n2701 & n2906 ;
  assign n2947 = n2946 ^ n2698 ;
  assign n2950 = n2949 ^ n2947 ;
  assign n2953 = n2706 & ~n2906 ;
  assign n2954 = n2953 ^ n2703 ;
  assign n2951 = n2173 & ~n2373 ;
  assign n2952 = n2951 ^ n2170 ;
  assign n2955 = n2954 ^ n2952 ;
  assign n2958 = n2711 & ~n2906 ;
  assign n2959 = n2958 ^ n2710 ;
  assign n2956 = n2178 & ~n2373 ;
  assign n2957 = n2956 ^ n2177 ;
  assign n2960 = n2959 ^ n2957 ;
  assign n2963 = n2183 & n2373 ;
  assign n2964 = n2963 ^ n2182 ;
  assign n2961 = n2716 & n2906 ;
  assign n2962 = n2961 ^ n2715 ;
  assign n2965 = n2964 ^ n2962 ;
  assign n2968 = n2188 & n2373 ;
  assign n2969 = n2968 ^ n2185 ;
  assign n2966 = n2721 & n2906 ;
  assign n2967 = n2966 ^ n2718 ;
  assign n2970 = n2969 ^ n2967 ;
  assign n2973 = n2726 & ~n2906 ;
  assign n2974 = n2973 ^ n2723 ;
  assign n2971 = n2193 & ~n2373 ;
  assign n2972 = n2971 ^ n2190 ;
  assign n2975 = n2974 ^ n2972 ;
  assign n2978 = n2731 & ~n2906 ;
  assign n2979 = n2978 ^ n2730 ;
  assign n2976 = n2198 & ~n2373 ;
  assign n2977 = n2976 ^ n2197 ;
  assign n2980 = n2979 ^ n2977 ;
  assign n2983 = n2203 & n2373 ;
  assign n2984 = n2983 ^ n2202 ;
  assign n2981 = n2736 & n2906 ;
  assign n2982 = n2981 ^ n2735 ;
  assign n2985 = n2984 ^ n2982 ;
  assign n2988 = n2208 & n2373 ;
  assign n2989 = n2988 ^ n2205 ;
  assign n2986 = n2741 & n2906 ;
  assign n2987 = n2986 ^ n2738 ;
  assign n2990 = n2989 ^ n2987 ;
  assign n2993 = n2746 & ~n2906 ;
  assign n2994 = n2993 ^ n2743 ;
  assign n2991 = n2213 & ~n2373 ;
  assign n2992 = n2991 ^ n2210 ;
  assign n2995 = n2994 ^ n2992 ;
  assign n2998 = n2751 & ~n2906 ;
  assign n2999 = n2998 ^ n2750 ;
  assign n2996 = n2218 & ~n2373 ;
  assign n2997 = n2996 ^ n2217 ;
  assign n3000 = n2999 ^ n2997 ;
  assign n3003 = n2223 & n2373 ;
  assign n3004 = n3003 ^ n2222 ;
  assign n3001 = n2756 & n2906 ;
  assign n3002 = n3001 ^ n2755 ;
  assign n3005 = n3004 ^ n3002 ;
  assign n3008 = n2228 & n2373 ;
  assign n3009 = n3008 ^ n2225 ;
  assign n3006 = n2761 & n2906 ;
  assign n3007 = n3006 ^ n2758 ;
  assign n3010 = n3009 ^ n3007 ;
  assign n3013 = n2766 & ~n2906 ;
  assign n3014 = n3013 ^ n2763 ;
  assign n3011 = n2233 & ~n2373 ;
  assign n3012 = n3011 ^ n2230 ;
  assign n3015 = n3014 ^ n3012 ;
  assign n3018 = n2771 & ~n2906 ;
  assign n3019 = n3018 ^ n2770 ;
  assign n3016 = n2238 & ~n2373 ;
  assign n3017 = n3016 ^ n2237 ;
  assign n3020 = n3019 ^ n3017 ;
  assign n3023 = n2243 & n2373 ;
  assign n3024 = n3023 ^ n2242 ;
  assign n3021 = n2776 & n2906 ;
  assign n3022 = n3021 ^ n2775 ;
  assign n3025 = n3024 ^ n3022 ;
  assign n3028 = n2248 & ~n2373 ;
  assign n3029 = n3028 ^ n2245 ;
  assign n3026 = n2781 & n2906 ;
  assign n3027 = n3026 ^ n2778 ;
  assign n3030 = n3029 ^ n3027 ;
  assign n3033 = n2786 & ~n2906 ;
  assign n3034 = n3033 ^ n2783 ;
  assign n3031 = n2253 & ~n2373 ;
  assign n3032 = n3031 ^ n2250 ;
  assign n3035 = n3034 ^ n3032 ;
  assign n3038 = n2791 & ~n2906 ;
  assign n3039 = n3038 ^ n2790 ;
  assign n3036 = n2258 & ~n2373 ;
  assign n3037 = n3036 ^ n2257 ;
  assign n3040 = n3039 ^ n3037 ;
  assign n3043 = n2796 & n2906 ;
  assign n3044 = n3043 ^ n2795 ;
  assign n3041 = n2263 & n2373 ;
  assign n3042 = n3041 ^ n2262 ;
  assign n3045 = n3044 ^ n3042 ;
  assign n3048 = n2268 & ~n2373 ;
  assign n3049 = n3048 ^ n2265 ;
  assign n3046 = n2801 & ~n2906 ;
  assign n3047 = n3046 ^ n2798 ;
  assign n3050 = n3049 ^ n3047 ;
  assign n3053 = n2806 & n2906 ;
  assign n3054 = n3053 ^ n2803 ;
  assign n3051 = n2273 & n2373 ;
  assign n3052 = n3051 ^ n2270 ;
  assign n3055 = n3054 ^ n3052 ;
  assign n3056 = n2812 ^ n2809 ;
  assign n3057 = ~n2906 & n3056 ;
  assign n3058 = n3057 ^ n2809 ;
  assign n3059 = n2279 ^ n2276 ;
  assign n3060 = ~n2373 & n3059 ;
  assign n3061 = n3060 ^ n2276 ;
  assign n3062 = ~n3058 & n3061 ;
  assign n3063 = n3062 ^ n3054 ;
  assign n3064 = ~n3055 & ~n3063 ;
  assign n3065 = n3064 ^ n3054 ;
  assign n3066 = n3065 ^ n3047 ;
  assign n3067 = ~n3050 & n3066 ;
  assign n3068 = n3067 ^ n3047 ;
  assign n3069 = n3068 ^ n3044 ;
  assign n3070 = ~n3045 & n3069 ;
  assign n3071 = n3070 ^ n3044 ;
  assign n3072 = n3071 ^ n3037 ;
  assign n3073 = ~n3040 & ~n3072 ;
  assign n3074 = n3073 ^ n3037 ;
  assign n3075 = n3074 ^ n3034 ;
  assign n3076 = ~n3035 & ~n3075 ;
  assign n3077 = n3076 ^ n3034 ;
  assign n3078 = n3077 ^ n3027 ;
  assign n3079 = ~n3030 & n3078 ;
  assign n3080 = n3079 ^ n3027 ;
  assign n3081 = n3080 ^ n3024 ;
  assign n3082 = ~n3025 & ~n3081 ;
  assign n3083 = n3082 ^ n3024 ;
  assign n3084 = n3083 ^ n3017 ;
  assign n3085 = ~n3020 & n3084 ;
  assign n3086 = n3085 ^ n3017 ;
  assign n3087 = n3086 ^ n3014 ;
  assign n3088 = ~n3015 & ~n3087 ;
  assign n3089 = n3088 ^ n3014 ;
  assign n3090 = n3089 ^ n3007 ;
  assign n3091 = ~n3010 & n3090 ;
  assign n3092 = n3091 ^ n3007 ;
  assign n3093 = n3092 ^ n3004 ;
  assign n3094 = ~n3005 & ~n3093 ;
  assign n3095 = n3094 ^ n3004 ;
  assign n3096 = n3095 ^ n2997 ;
  assign n3097 = ~n3000 & n3096 ;
  assign n3098 = n3097 ^ n2997 ;
  assign n3099 = n3098 ^ n2994 ;
  assign n3100 = ~n2995 & ~n3099 ;
  assign n3101 = n3100 ^ n2994 ;
  assign n3102 = n3101 ^ n2987 ;
  assign n3103 = ~n2990 & n3102 ;
  assign n3104 = n3103 ^ n2987 ;
  assign n3105 = n3104 ^ n2984 ;
  assign n3106 = ~n2985 & ~n3105 ;
  assign n3107 = n3106 ^ n2984 ;
  assign n3108 = n3107 ^ n2977 ;
  assign n3109 = ~n2980 & n3108 ;
  assign n3110 = n3109 ^ n2977 ;
  assign n3111 = n3110 ^ n2974 ;
  assign n3112 = ~n2975 & ~n3111 ;
  assign n3113 = n3112 ^ n2974 ;
  assign n3114 = n3113 ^ n2967 ;
  assign n3115 = ~n2970 & n3114 ;
  assign n3116 = n3115 ^ n2967 ;
  assign n3117 = n3116 ^ n2964 ;
  assign n3118 = ~n2965 & ~n3117 ;
  assign n3119 = n3118 ^ n2964 ;
  assign n3120 = n3119 ^ n2957 ;
  assign n3121 = ~n2960 & n3120 ;
  assign n3122 = n3121 ^ n2957 ;
  assign n3123 = n3122 ^ n2954 ;
  assign n3124 = ~n2955 & ~n3123 ;
  assign n3125 = n3124 ^ n2954 ;
  assign n3126 = n3125 ^ n2947 ;
  assign n3127 = ~n2950 & n3126 ;
  assign n3128 = n3127 ^ n2947 ;
  assign n3129 = n3128 ^ n2944 ;
  assign n3130 = ~n2945 & ~n3129 ;
  assign n3131 = n3130 ^ n2944 ;
  assign n3132 = n3131 ^ n2937 ;
  assign n3133 = ~n2940 & n3132 ;
  assign n3134 = n3133 ^ n2937 ;
  assign n3135 = n3134 ^ n2934 ;
  assign n3136 = ~n2935 & n3135 ;
  assign n3137 = n3136 ^ n2934 ;
  assign n3138 = n3137 ^ n2927 ;
  assign n3139 = ~n2930 & ~n3138 ;
  assign n3140 = n3139 ^ n2927 ;
  assign n3141 = n3140 ^ n2924 ;
  assign n3142 = ~n2925 & ~n3141 ;
  assign n3143 = n3142 ^ n2924 ;
  assign n3144 = n3143 ^ n2917 ;
  assign n3145 = ~n2920 & ~n3144 ;
  assign n3146 = n3145 ^ n2917 ;
  assign n3147 = n3146 ^ n2912 ;
  assign n3148 = ~n2915 & ~n3147 ;
  assign n3149 = n3148 ^ n2912 ;
  assign n3150 = n3149 ^ n2375 ;
  assign n3151 = ~n2909 & ~n3150 ;
  assign n3152 = n3151 ^ n2908 ;
  assign n3153 = n3152 ^ n518 ;
  assign n3154 = ~n2910 & n3153 ;
  assign n3155 = n3154 ^ n515 ;
  assign n3156 = n2909 & n3155 ;
  assign n3157 = n3156 ^ n2375 ;
  assign n1203 = x190 ^ x158 ;
  assign n1204 = x191 ^ x159 ;
  assign n1206 = x188 ^ x156 ;
  assign n1208 = x186 ^ x154 ;
  assign n1210 = x184 ^ x152 ;
  assign n1212 = x182 ^ x150 ;
  assign n1214 = x180 ^ x148 ;
  assign n1216 = x178 ^ x146 ;
  assign n1218 = x176 ^ x144 ;
  assign n1220 = x174 ^ x142 ;
  assign n1222 = x172 ^ x140 ;
  assign n1224 = x170 ^ x138 ;
  assign n1226 = x168 ^ x136 ;
  assign n1228 = x166 ^ x134 ;
  assign n1230 = x164 ^ x132 ;
  assign n1232 = x162 ^ x130 ;
  assign n1234 = x128 & ~x160 ;
  assign n1235 = n1234 ^ x162 ;
  assign n1233 = x162 ^ x129 ;
  assign n1236 = n1235 ^ n1233 ;
  assign n1237 = x161 ^ x129 ;
  assign n1238 = n1236 & ~n1237 ;
  assign n1239 = n1238 ^ n1233 ;
  assign n1240 = ~n1232 & n1239 ;
  assign n1241 = n1240 ^ x130 ;
  assign n1242 = n1241 ^ x164 ;
  assign n1231 = x164 ^ x131 ;
  assign n1243 = n1242 ^ n1231 ;
  assign n1244 = x163 ^ x131 ;
  assign n1245 = n1243 & ~n1244 ;
  assign n1246 = n1245 ^ n1231 ;
  assign n1247 = ~n1230 & n1246 ;
  assign n1248 = n1247 ^ x132 ;
  assign n1249 = n1248 ^ x166 ;
  assign n1229 = x166 ^ x133 ;
  assign n1250 = n1249 ^ n1229 ;
  assign n1251 = x165 ^ x133 ;
  assign n1252 = n1250 & ~n1251 ;
  assign n1253 = n1252 ^ n1229 ;
  assign n1254 = ~n1228 & n1253 ;
  assign n1255 = n1254 ^ x134 ;
  assign n1256 = n1255 ^ x168 ;
  assign n1227 = x168 ^ x135 ;
  assign n1257 = n1256 ^ n1227 ;
  assign n1258 = x167 ^ x135 ;
  assign n1259 = n1257 & ~n1258 ;
  assign n1260 = n1259 ^ n1227 ;
  assign n1261 = ~n1226 & n1260 ;
  assign n1262 = n1261 ^ x136 ;
  assign n1263 = n1262 ^ x170 ;
  assign n1225 = x170 ^ x137 ;
  assign n1264 = n1263 ^ n1225 ;
  assign n1265 = x169 ^ x137 ;
  assign n1266 = n1264 & ~n1265 ;
  assign n1267 = n1266 ^ n1225 ;
  assign n1268 = ~n1224 & n1267 ;
  assign n1269 = n1268 ^ x138 ;
  assign n1270 = n1269 ^ x172 ;
  assign n1223 = x172 ^ x139 ;
  assign n1271 = n1270 ^ n1223 ;
  assign n1272 = x171 ^ x139 ;
  assign n1273 = n1271 & ~n1272 ;
  assign n1274 = n1273 ^ n1223 ;
  assign n1275 = ~n1222 & n1274 ;
  assign n1276 = n1275 ^ x140 ;
  assign n1277 = n1276 ^ x174 ;
  assign n1221 = x174 ^ x141 ;
  assign n1278 = n1277 ^ n1221 ;
  assign n1279 = x173 ^ x141 ;
  assign n1280 = n1278 & ~n1279 ;
  assign n1281 = n1280 ^ n1221 ;
  assign n1282 = ~n1220 & n1281 ;
  assign n1283 = n1282 ^ x142 ;
  assign n1284 = n1283 ^ x176 ;
  assign n1219 = x176 ^ x143 ;
  assign n1285 = n1284 ^ n1219 ;
  assign n1286 = x175 ^ x143 ;
  assign n1287 = n1285 & ~n1286 ;
  assign n1288 = n1287 ^ n1219 ;
  assign n1289 = ~n1218 & n1288 ;
  assign n1290 = n1289 ^ x144 ;
  assign n1291 = n1290 ^ x178 ;
  assign n1217 = x178 ^ x145 ;
  assign n1292 = n1291 ^ n1217 ;
  assign n1293 = x177 ^ x145 ;
  assign n1294 = n1292 & ~n1293 ;
  assign n1295 = n1294 ^ n1217 ;
  assign n1296 = ~n1216 & n1295 ;
  assign n1297 = n1296 ^ x146 ;
  assign n1298 = n1297 ^ x180 ;
  assign n1215 = x180 ^ x147 ;
  assign n1299 = n1298 ^ n1215 ;
  assign n1300 = x179 ^ x147 ;
  assign n1301 = n1299 & ~n1300 ;
  assign n1302 = n1301 ^ n1215 ;
  assign n1303 = ~n1214 & n1302 ;
  assign n1304 = n1303 ^ x148 ;
  assign n1305 = n1304 ^ x182 ;
  assign n1213 = x182 ^ x149 ;
  assign n1306 = n1305 ^ n1213 ;
  assign n1307 = x181 ^ x149 ;
  assign n1308 = n1306 & ~n1307 ;
  assign n1309 = n1308 ^ n1213 ;
  assign n1310 = ~n1212 & n1309 ;
  assign n1311 = n1310 ^ x150 ;
  assign n1312 = n1311 ^ x184 ;
  assign n1211 = x184 ^ x151 ;
  assign n1313 = n1312 ^ n1211 ;
  assign n1314 = x183 ^ x151 ;
  assign n1315 = n1313 & ~n1314 ;
  assign n1316 = n1315 ^ n1211 ;
  assign n1317 = ~n1210 & n1316 ;
  assign n1318 = n1317 ^ x152 ;
  assign n1319 = n1318 ^ x186 ;
  assign n1209 = x186 ^ x153 ;
  assign n1320 = n1319 ^ n1209 ;
  assign n1321 = x185 ^ x153 ;
  assign n1322 = n1320 & ~n1321 ;
  assign n1323 = n1322 ^ n1209 ;
  assign n1324 = ~n1208 & n1323 ;
  assign n1325 = n1324 ^ x154 ;
  assign n1326 = n1325 ^ x188 ;
  assign n1207 = x188 ^ x155 ;
  assign n1327 = n1326 ^ n1207 ;
  assign n1328 = x187 ^ x155 ;
  assign n1329 = n1327 & ~n1328 ;
  assign n1330 = n1329 ^ n1207 ;
  assign n1331 = ~n1206 & n1330 ;
  assign n1332 = n1331 ^ x156 ;
  assign n1333 = n1332 ^ x190 ;
  assign n1205 = x190 ^ x157 ;
  assign n1334 = n1333 ^ n1205 ;
  assign n1335 = x189 ^ x157 ;
  assign n1336 = n1334 & ~n1335 ;
  assign n1337 = n1336 ^ n1205 ;
  assign n1338 = ~n1203 & n1337 ;
  assign n1339 = n1338 ^ x158 ;
  assign n1340 = n1339 ^ x191 ;
  assign n1341 = ~n1204 & n1340 ;
  assign n1342 = n1341 ^ x159 ;
  assign n1343 = n1203 & ~n1342 ;
  assign n1344 = n1343 ^ x158 ;
  assign n1061 = x254 ^ x222 ;
  assign n1062 = x255 ^ x223 ;
  assign n1064 = x252 ^ x220 ;
  assign n1066 = x250 ^ x218 ;
  assign n1068 = x248 ^ x216 ;
  assign n1070 = x246 ^ x214 ;
  assign n1072 = x244 ^ x212 ;
  assign n1074 = x242 ^ x210 ;
  assign n1076 = x240 ^ x208 ;
  assign n1078 = x238 ^ x206 ;
  assign n1080 = x236 ^ x204 ;
  assign n1082 = x234 ^ x202 ;
  assign n1084 = x232 ^ x200 ;
  assign n1086 = x230 ^ x198 ;
  assign n1088 = x228 ^ x196 ;
  assign n1090 = x226 ^ x194 ;
  assign n1092 = x192 & ~x224 ;
  assign n1093 = n1092 ^ x226 ;
  assign n1091 = x226 ^ x193 ;
  assign n1094 = n1093 ^ n1091 ;
  assign n1095 = x225 ^ x193 ;
  assign n1096 = n1094 & ~n1095 ;
  assign n1097 = n1096 ^ n1091 ;
  assign n1098 = ~n1090 & n1097 ;
  assign n1099 = n1098 ^ x194 ;
  assign n1100 = n1099 ^ x228 ;
  assign n1089 = x228 ^ x195 ;
  assign n1101 = n1100 ^ n1089 ;
  assign n1102 = x227 ^ x195 ;
  assign n1103 = n1101 & ~n1102 ;
  assign n1104 = n1103 ^ n1089 ;
  assign n1105 = ~n1088 & n1104 ;
  assign n1106 = n1105 ^ x196 ;
  assign n1107 = n1106 ^ x230 ;
  assign n1087 = x230 ^ x197 ;
  assign n1108 = n1107 ^ n1087 ;
  assign n1109 = x229 ^ x197 ;
  assign n1110 = n1108 & ~n1109 ;
  assign n1111 = n1110 ^ n1087 ;
  assign n1112 = ~n1086 & n1111 ;
  assign n1113 = n1112 ^ x198 ;
  assign n1114 = n1113 ^ x232 ;
  assign n1085 = x232 ^ x199 ;
  assign n1115 = n1114 ^ n1085 ;
  assign n1116 = x231 ^ x199 ;
  assign n1117 = n1115 & ~n1116 ;
  assign n1118 = n1117 ^ n1085 ;
  assign n1119 = ~n1084 & n1118 ;
  assign n1120 = n1119 ^ x200 ;
  assign n1121 = n1120 ^ x234 ;
  assign n1083 = x234 ^ x201 ;
  assign n1122 = n1121 ^ n1083 ;
  assign n1123 = x233 ^ x201 ;
  assign n1124 = n1122 & ~n1123 ;
  assign n1125 = n1124 ^ n1083 ;
  assign n1126 = ~n1082 & n1125 ;
  assign n1127 = n1126 ^ x202 ;
  assign n1128 = n1127 ^ x236 ;
  assign n1081 = x236 ^ x203 ;
  assign n1129 = n1128 ^ n1081 ;
  assign n1130 = x235 ^ x203 ;
  assign n1131 = n1129 & ~n1130 ;
  assign n1132 = n1131 ^ n1081 ;
  assign n1133 = ~n1080 & n1132 ;
  assign n1134 = n1133 ^ x204 ;
  assign n1135 = n1134 ^ x238 ;
  assign n1079 = x238 ^ x205 ;
  assign n1136 = n1135 ^ n1079 ;
  assign n1137 = x237 ^ x205 ;
  assign n1138 = n1136 & ~n1137 ;
  assign n1139 = n1138 ^ n1079 ;
  assign n1140 = ~n1078 & n1139 ;
  assign n1141 = n1140 ^ x206 ;
  assign n1142 = n1141 ^ x240 ;
  assign n1077 = x240 ^ x207 ;
  assign n1143 = n1142 ^ n1077 ;
  assign n1144 = x239 ^ x207 ;
  assign n1145 = n1143 & ~n1144 ;
  assign n1146 = n1145 ^ n1077 ;
  assign n1147 = ~n1076 & n1146 ;
  assign n1148 = n1147 ^ x208 ;
  assign n1149 = n1148 ^ x242 ;
  assign n1075 = x242 ^ x209 ;
  assign n1150 = n1149 ^ n1075 ;
  assign n1151 = x241 ^ x209 ;
  assign n1152 = n1150 & ~n1151 ;
  assign n1153 = n1152 ^ n1075 ;
  assign n1154 = ~n1074 & n1153 ;
  assign n1155 = n1154 ^ x210 ;
  assign n1156 = n1155 ^ x244 ;
  assign n1073 = x244 ^ x211 ;
  assign n1157 = n1156 ^ n1073 ;
  assign n1158 = x243 ^ x211 ;
  assign n1159 = n1157 & ~n1158 ;
  assign n1160 = n1159 ^ n1073 ;
  assign n1161 = ~n1072 & n1160 ;
  assign n1162 = n1161 ^ x212 ;
  assign n1163 = n1162 ^ x246 ;
  assign n1071 = x246 ^ x213 ;
  assign n1164 = n1163 ^ n1071 ;
  assign n1165 = x245 ^ x213 ;
  assign n1166 = n1164 & ~n1165 ;
  assign n1167 = n1166 ^ n1071 ;
  assign n1168 = ~n1070 & n1167 ;
  assign n1169 = n1168 ^ x214 ;
  assign n1170 = n1169 ^ x248 ;
  assign n1069 = x248 ^ x215 ;
  assign n1171 = n1170 ^ n1069 ;
  assign n1172 = x247 ^ x215 ;
  assign n1173 = n1171 & ~n1172 ;
  assign n1174 = n1173 ^ n1069 ;
  assign n1175 = ~n1068 & n1174 ;
  assign n1176 = n1175 ^ x216 ;
  assign n1177 = n1176 ^ x250 ;
  assign n1067 = x250 ^ x217 ;
  assign n1178 = n1177 ^ n1067 ;
  assign n1179 = x249 ^ x217 ;
  assign n1180 = n1178 & ~n1179 ;
  assign n1181 = n1180 ^ n1067 ;
  assign n1182 = ~n1066 & n1181 ;
  assign n1183 = n1182 ^ x218 ;
  assign n1184 = n1183 ^ x252 ;
  assign n1065 = x252 ^ x219 ;
  assign n1185 = n1184 ^ n1065 ;
  assign n1186 = x251 ^ x219 ;
  assign n1187 = n1185 & ~n1186 ;
  assign n1188 = n1187 ^ n1065 ;
  assign n1189 = ~n1064 & n1188 ;
  assign n1190 = n1189 ^ x220 ;
  assign n1191 = n1190 ^ x254 ;
  assign n1063 = x254 ^ x221 ;
  assign n1192 = n1191 ^ n1063 ;
  assign n1193 = x253 ^ x221 ;
  assign n1194 = n1192 & ~n1193 ;
  assign n1195 = n1194 ^ n1063 ;
  assign n1196 = ~n1061 & n1195 ;
  assign n1197 = n1196 ^ x222 ;
  assign n1198 = n1197 ^ x255 ;
  assign n1199 = ~n1062 & n1198 ;
  assign n1200 = n1199 ^ x223 ;
  assign n1201 = n1061 & ~n1200 ;
  assign n1202 = n1201 ^ x222 ;
  assign n1345 = n1344 ^ n1202 ;
  assign n1346 = n524 ^ n523 ;
  assign n1349 = n1193 & ~n1200 ;
  assign n1350 = n1349 ^ x221 ;
  assign n1347 = n1335 & ~n1342 ;
  assign n1348 = n1347 ^ x157 ;
  assign n1351 = n1350 ^ n1348 ;
  assign n1354 = n1064 & ~n1200 ;
  assign n1355 = n1354 ^ x220 ;
  assign n1352 = n1206 & ~n1342 ;
  assign n1353 = n1352 ^ x156 ;
  assign n1356 = n1355 ^ n1353 ;
  assign n1359 = n1328 & ~n1342 ;
  assign n1360 = n1359 ^ x155 ;
  assign n1357 = n1186 & ~n1200 ;
  assign n1358 = n1357 ^ x219 ;
  assign n1361 = n1360 ^ n1358 ;
  assign n1364 = n1066 & ~n1200 ;
  assign n1365 = n1364 ^ x218 ;
  assign n1362 = n1208 & ~n1342 ;
  assign n1363 = n1362 ^ x154 ;
  assign n1366 = n1365 ^ n1363 ;
  assign n1369 = n1321 & ~n1342 ;
  assign n1370 = n1369 ^ x153 ;
  assign n1367 = n1179 & ~n1200 ;
  assign n1368 = n1367 ^ x217 ;
  assign n1371 = n1370 ^ n1368 ;
  assign n1374 = n1068 & ~n1200 ;
  assign n1375 = n1374 ^ x216 ;
  assign n1372 = n1210 & ~n1342 ;
  assign n1373 = n1372 ^ x152 ;
  assign n1376 = n1375 ^ n1373 ;
  assign n1379 = n1314 & ~n1342 ;
  assign n1380 = n1379 ^ x151 ;
  assign n1377 = n1172 & ~n1200 ;
  assign n1378 = n1377 ^ x215 ;
  assign n1381 = n1380 ^ n1378 ;
  assign n1384 = n1070 & ~n1200 ;
  assign n1385 = n1384 ^ x214 ;
  assign n1382 = n1212 & ~n1342 ;
  assign n1383 = n1382 ^ x150 ;
  assign n1386 = n1385 ^ n1383 ;
  assign n1389 = n1307 & ~n1342 ;
  assign n1390 = n1389 ^ x149 ;
  assign n1387 = n1165 & ~n1200 ;
  assign n1388 = n1387 ^ x213 ;
  assign n1391 = n1390 ^ n1388 ;
  assign n1394 = n1072 & ~n1200 ;
  assign n1395 = n1394 ^ x212 ;
  assign n1392 = n1214 & ~n1342 ;
  assign n1393 = n1392 ^ x148 ;
  assign n1396 = n1395 ^ n1393 ;
  assign n1399 = n1300 & ~n1342 ;
  assign n1400 = n1399 ^ x147 ;
  assign n1397 = n1158 & ~n1200 ;
  assign n1398 = n1397 ^ x211 ;
  assign n1401 = n1400 ^ n1398 ;
  assign n1404 = n1074 & ~n1200 ;
  assign n1405 = n1404 ^ x210 ;
  assign n1402 = n1216 & ~n1342 ;
  assign n1403 = n1402 ^ x146 ;
  assign n1406 = n1405 ^ n1403 ;
  assign n1409 = n1293 & ~n1342 ;
  assign n1410 = n1409 ^ x145 ;
  assign n1407 = n1151 & ~n1200 ;
  assign n1408 = n1407 ^ x209 ;
  assign n1411 = n1410 ^ n1408 ;
  assign n1414 = n1076 & ~n1200 ;
  assign n1415 = n1414 ^ x208 ;
  assign n1412 = n1218 & ~n1342 ;
  assign n1413 = n1412 ^ x144 ;
  assign n1416 = n1415 ^ n1413 ;
  assign n1419 = n1286 & ~n1342 ;
  assign n1420 = n1419 ^ x143 ;
  assign n1417 = n1144 & ~n1200 ;
  assign n1418 = n1417 ^ x207 ;
  assign n1421 = n1420 ^ n1418 ;
  assign n1424 = n1078 & ~n1200 ;
  assign n1425 = n1424 ^ x206 ;
  assign n1422 = n1220 & ~n1342 ;
  assign n1423 = n1422 ^ x142 ;
  assign n1426 = n1425 ^ n1423 ;
  assign n1429 = n1279 & ~n1342 ;
  assign n1430 = n1429 ^ x141 ;
  assign n1427 = n1137 & ~n1200 ;
  assign n1428 = n1427 ^ x205 ;
  assign n1431 = n1430 ^ n1428 ;
  assign n1434 = n1080 & ~n1200 ;
  assign n1435 = n1434 ^ x204 ;
  assign n1432 = n1222 & ~n1342 ;
  assign n1433 = n1432 ^ x140 ;
  assign n1436 = n1435 ^ n1433 ;
  assign n1439 = n1272 & ~n1342 ;
  assign n1440 = n1439 ^ x139 ;
  assign n1437 = n1130 & ~n1200 ;
  assign n1438 = n1437 ^ x203 ;
  assign n1441 = n1440 ^ n1438 ;
  assign n1444 = n1082 & ~n1200 ;
  assign n1445 = n1444 ^ x202 ;
  assign n1442 = n1224 & ~n1342 ;
  assign n1443 = n1442 ^ x138 ;
  assign n1446 = n1445 ^ n1443 ;
  assign n1449 = n1265 & ~n1342 ;
  assign n1450 = n1449 ^ x137 ;
  assign n1447 = n1123 & ~n1200 ;
  assign n1448 = n1447 ^ x201 ;
  assign n1451 = n1450 ^ n1448 ;
  assign n1454 = n1084 & ~n1200 ;
  assign n1455 = n1454 ^ x200 ;
  assign n1452 = n1226 & ~n1342 ;
  assign n1453 = n1452 ^ x136 ;
  assign n1456 = n1455 ^ n1453 ;
  assign n1459 = n1258 & ~n1342 ;
  assign n1460 = n1459 ^ x135 ;
  assign n1457 = n1116 & ~n1200 ;
  assign n1458 = n1457 ^ x199 ;
  assign n1461 = n1460 ^ n1458 ;
  assign n1464 = n1086 & ~n1200 ;
  assign n1465 = n1464 ^ x198 ;
  assign n1462 = n1228 & ~n1342 ;
  assign n1463 = n1462 ^ x134 ;
  assign n1466 = n1465 ^ n1463 ;
  assign n1469 = n1251 & ~n1342 ;
  assign n1470 = n1469 ^ x133 ;
  assign n1467 = n1109 & ~n1200 ;
  assign n1468 = n1467 ^ x197 ;
  assign n1471 = n1470 ^ n1468 ;
  assign n1474 = n1088 & ~n1200 ;
  assign n1475 = n1474 ^ x196 ;
  assign n1472 = n1230 & ~n1342 ;
  assign n1473 = n1472 ^ x132 ;
  assign n1476 = n1475 ^ n1473 ;
  assign n1479 = n1102 & ~n1200 ;
  assign n1480 = n1479 ^ x195 ;
  assign n1477 = n1244 & ~n1342 ;
  assign n1478 = n1477 ^ x131 ;
  assign n1481 = n1480 ^ n1478 ;
  assign n1484 = n1232 & ~n1342 ;
  assign n1485 = n1484 ^ x130 ;
  assign n1482 = n1090 & ~n1200 ;
  assign n1483 = n1482 ^ x194 ;
  assign n1486 = n1485 ^ n1483 ;
  assign n1489 = n1095 & ~n1200 ;
  assign n1490 = n1489 ^ x193 ;
  assign n1487 = n1237 & ~n1342 ;
  assign n1488 = n1487 ^ x129 ;
  assign n1491 = n1490 ^ n1488 ;
  assign n1492 = x224 ^ x192 ;
  assign n1493 = ~n1200 & n1492 ;
  assign n1494 = n1493 ^ x192 ;
  assign n1495 = x160 ^ x128 ;
  assign n1496 = ~n1342 & n1495 ;
  assign n1497 = n1496 ^ x128 ;
  assign n1498 = ~n1494 & n1497 ;
  assign n1499 = n1498 ^ n1490 ;
  assign n1500 = ~n1491 & ~n1499 ;
  assign n1501 = n1500 ^ n1490 ;
  assign n1502 = n1501 ^ n1485 ;
  assign n1503 = ~n1486 & ~n1502 ;
  assign n1504 = n1503 ^ n1485 ;
  assign n1505 = n1504 ^ n1480 ;
  assign n1506 = ~n1481 & ~n1505 ;
  assign n1507 = n1506 ^ n1480 ;
  assign n1508 = n1507 ^ n1473 ;
  assign n1509 = ~n1476 & ~n1508 ;
  assign n1510 = n1509 ^ n1473 ;
  assign n1511 = n1510 ^ n1470 ;
  assign n1512 = ~n1471 & n1511 ;
  assign n1513 = n1512 ^ n1470 ;
  assign n1514 = n1513 ^ n1463 ;
  assign n1515 = ~n1466 & n1514 ;
  assign n1516 = n1515 ^ n1463 ;
  assign n1517 = n1516 ^ n1460 ;
  assign n1518 = ~n1461 & n1517 ;
  assign n1519 = n1518 ^ n1460 ;
  assign n1520 = n1519 ^ n1453 ;
  assign n1521 = ~n1456 & n1520 ;
  assign n1522 = n1521 ^ n1453 ;
  assign n1523 = n1522 ^ n1450 ;
  assign n1524 = ~n1451 & n1523 ;
  assign n1525 = n1524 ^ n1450 ;
  assign n1526 = n1525 ^ n1443 ;
  assign n1527 = ~n1446 & n1526 ;
  assign n1528 = n1527 ^ n1443 ;
  assign n1529 = n1528 ^ n1440 ;
  assign n1530 = ~n1441 & n1529 ;
  assign n1531 = n1530 ^ n1440 ;
  assign n1532 = n1531 ^ n1433 ;
  assign n1533 = ~n1436 & n1532 ;
  assign n1534 = n1533 ^ n1433 ;
  assign n1535 = n1534 ^ n1430 ;
  assign n1536 = ~n1431 & n1535 ;
  assign n1537 = n1536 ^ n1430 ;
  assign n1538 = n1537 ^ n1423 ;
  assign n1539 = ~n1426 & n1538 ;
  assign n1540 = n1539 ^ n1423 ;
  assign n1541 = n1540 ^ n1420 ;
  assign n1542 = ~n1421 & n1541 ;
  assign n1543 = n1542 ^ n1420 ;
  assign n1544 = n1543 ^ n1413 ;
  assign n1545 = ~n1416 & n1544 ;
  assign n1546 = n1545 ^ n1413 ;
  assign n1547 = n1546 ^ n1410 ;
  assign n1548 = ~n1411 & n1547 ;
  assign n1549 = n1548 ^ n1410 ;
  assign n1550 = n1549 ^ n1403 ;
  assign n1551 = ~n1406 & n1550 ;
  assign n1552 = n1551 ^ n1403 ;
  assign n1553 = n1552 ^ n1400 ;
  assign n1554 = ~n1401 & n1553 ;
  assign n1555 = n1554 ^ n1400 ;
  assign n1556 = n1555 ^ n1393 ;
  assign n1557 = ~n1396 & n1556 ;
  assign n1558 = n1557 ^ n1393 ;
  assign n1559 = n1558 ^ n1390 ;
  assign n1560 = ~n1391 & n1559 ;
  assign n1561 = n1560 ^ n1390 ;
  assign n1562 = n1561 ^ n1383 ;
  assign n1563 = ~n1386 & n1562 ;
  assign n1564 = n1563 ^ n1383 ;
  assign n1565 = n1564 ^ n1380 ;
  assign n1566 = ~n1381 & n1565 ;
  assign n1567 = n1566 ^ n1380 ;
  assign n1568 = n1567 ^ n1373 ;
  assign n1569 = ~n1376 & n1568 ;
  assign n1570 = n1569 ^ n1373 ;
  assign n1571 = n1570 ^ n1370 ;
  assign n1572 = ~n1371 & n1571 ;
  assign n1573 = n1572 ^ n1370 ;
  assign n1574 = n1573 ^ n1363 ;
  assign n1575 = ~n1366 & n1574 ;
  assign n1576 = n1575 ^ n1363 ;
  assign n1577 = n1576 ^ n1360 ;
  assign n1578 = ~n1361 & n1577 ;
  assign n1579 = n1578 ^ n1360 ;
  assign n1580 = n1579 ^ n1355 ;
  assign n1581 = ~n1356 & ~n1580 ;
  assign n1582 = n1581 ^ n1355 ;
  assign n1583 = n1582 ^ n1350 ;
  assign n1584 = ~n1351 & ~n1583 ;
  assign n1585 = n1584 ^ n1348 ;
  assign n1586 = n1585 ^ n1344 ;
  assign n1587 = ~n1345 & ~n1586 ;
  assign n1588 = n1587 ^ n1202 ;
  assign n1589 = n1588 ^ n524 ;
  assign n1590 = ~n1346 & n1589 ;
  assign n1591 = n1590 ^ n523 ;
  assign n1592 = n1345 & ~n1591 ;
  assign n1593 = n1592 ^ n1202 ;
  assign n670 = x126 ^ x94 ;
  assign n671 = x127 ^ x95 ;
  assign n673 = x124 ^ x92 ;
  assign n675 = x122 ^ x90 ;
  assign n677 = x120 ^ x88 ;
  assign n679 = x118 ^ x86 ;
  assign n681 = x116 ^ x84 ;
  assign n683 = x114 ^ x82 ;
  assign n685 = x112 ^ x80 ;
  assign n687 = x110 ^ x78 ;
  assign n689 = x108 ^ x76 ;
  assign n691 = x106 ^ x74 ;
  assign n693 = x104 ^ x72 ;
  assign n695 = x102 ^ x70 ;
  assign n697 = x100 ^ x68 ;
  assign n699 = x98 ^ x66 ;
  assign n701 = x64 & ~x96 ;
  assign n702 = n701 ^ x98 ;
  assign n700 = x98 ^ x65 ;
  assign n703 = n702 ^ n700 ;
  assign n704 = x97 ^ x65 ;
  assign n705 = n703 & ~n704 ;
  assign n706 = n705 ^ n700 ;
  assign n707 = ~n699 & n706 ;
  assign n708 = n707 ^ x66 ;
  assign n709 = n708 ^ x100 ;
  assign n698 = x100 ^ x67 ;
  assign n710 = n709 ^ n698 ;
  assign n711 = x99 ^ x67 ;
  assign n712 = n710 & ~n711 ;
  assign n713 = n712 ^ n698 ;
  assign n714 = ~n697 & n713 ;
  assign n715 = n714 ^ x68 ;
  assign n716 = n715 ^ x102 ;
  assign n696 = x102 ^ x69 ;
  assign n717 = n716 ^ n696 ;
  assign n718 = x101 ^ x69 ;
  assign n719 = n717 & ~n718 ;
  assign n720 = n719 ^ n696 ;
  assign n721 = ~n695 & n720 ;
  assign n722 = n721 ^ x70 ;
  assign n723 = n722 ^ x104 ;
  assign n694 = x104 ^ x71 ;
  assign n724 = n723 ^ n694 ;
  assign n725 = x103 ^ x71 ;
  assign n726 = n724 & ~n725 ;
  assign n727 = n726 ^ n694 ;
  assign n728 = ~n693 & n727 ;
  assign n729 = n728 ^ x72 ;
  assign n730 = n729 ^ x106 ;
  assign n692 = x106 ^ x73 ;
  assign n731 = n730 ^ n692 ;
  assign n732 = x105 ^ x73 ;
  assign n733 = n731 & ~n732 ;
  assign n734 = n733 ^ n692 ;
  assign n735 = ~n691 & n734 ;
  assign n736 = n735 ^ x74 ;
  assign n737 = n736 ^ x108 ;
  assign n690 = x108 ^ x75 ;
  assign n738 = n737 ^ n690 ;
  assign n739 = x107 ^ x75 ;
  assign n740 = n738 & ~n739 ;
  assign n741 = n740 ^ n690 ;
  assign n742 = ~n689 & n741 ;
  assign n743 = n742 ^ x76 ;
  assign n744 = n743 ^ x110 ;
  assign n688 = x110 ^ x77 ;
  assign n745 = n744 ^ n688 ;
  assign n746 = x109 ^ x77 ;
  assign n747 = n745 & ~n746 ;
  assign n748 = n747 ^ n688 ;
  assign n749 = ~n687 & n748 ;
  assign n750 = n749 ^ x78 ;
  assign n751 = n750 ^ x112 ;
  assign n686 = x112 ^ x79 ;
  assign n752 = n751 ^ n686 ;
  assign n753 = x111 ^ x79 ;
  assign n754 = n752 & ~n753 ;
  assign n755 = n754 ^ n686 ;
  assign n756 = ~n685 & n755 ;
  assign n757 = n756 ^ x80 ;
  assign n758 = n757 ^ x114 ;
  assign n684 = x114 ^ x81 ;
  assign n759 = n758 ^ n684 ;
  assign n760 = x113 ^ x81 ;
  assign n761 = n759 & ~n760 ;
  assign n762 = n761 ^ n684 ;
  assign n763 = ~n683 & n762 ;
  assign n764 = n763 ^ x82 ;
  assign n765 = n764 ^ x116 ;
  assign n682 = x116 ^ x83 ;
  assign n766 = n765 ^ n682 ;
  assign n767 = x115 ^ x83 ;
  assign n768 = n766 & ~n767 ;
  assign n769 = n768 ^ n682 ;
  assign n770 = ~n681 & n769 ;
  assign n771 = n770 ^ x84 ;
  assign n772 = n771 ^ x118 ;
  assign n680 = x118 ^ x85 ;
  assign n773 = n772 ^ n680 ;
  assign n774 = x117 ^ x85 ;
  assign n775 = n773 & ~n774 ;
  assign n776 = n775 ^ n680 ;
  assign n777 = ~n679 & n776 ;
  assign n778 = n777 ^ x86 ;
  assign n779 = n778 ^ x120 ;
  assign n678 = x120 ^ x87 ;
  assign n780 = n779 ^ n678 ;
  assign n781 = x119 ^ x87 ;
  assign n782 = n780 & ~n781 ;
  assign n783 = n782 ^ n678 ;
  assign n784 = ~n677 & n783 ;
  assign n785 = n784 ^ x88 ;
  assign n786 = n785 ^ x122 ;
  assign n676 = x122 ^ x89 ;
  assign n787 = n786 ^ n676 ;
  assign n788 = x121 ^ x89 ;
  assign n789 = n787 & ~n788 ;
  assign n790 = n789 ^ n676 ;
  assign n791 = ~n675 & n790 ;
  assign n792 = n791 ^ x90 ;
  assign n793 = n792 ^ x124 ;
  assign n674 = x124 ^ x91 ;
  assign n794 = n793 ^ n674 ;
  assign n795 = x123 ^ x91 ;
  assign n796 = n794 & ~n795 ;
  assign n797 = n796 ^ n674 ;
  assign n798 = ~n673 & n797 ;
  assign n799 = n798 ^ x92 ;
  assign n800 = n799 ^ x126 ;
  assign n672 = x126 ^ x93 ;
  assign n801 = n800 ^ n672 ;
  assign n802 = x125 ^ x93 ;
  assign n803 = n801 & ~n802 ;
  assign n804 = n803 ^ n672 ;
  assign n805 = ~n670 & n804 ;
  assign n806 = n805 ^ x94 ;
  assign n807 = n806 ^ x127 ;
  assign n808 = ~n671 & n807 ;
  assign n809 = n808 ^ x95 ;
  assign n810 = n670 & ~n809 ;
  assign n811 = n810 ^ x94 ;
  assign n528 = x62 ^ x30 ;
  assign n529 = x63 ^ x31 ;
  assign n531 = x60 ^ x28 ;
  assign n533 = x58 ^ x26 ;
  assign n535 = x56 ^ x24 ;
  assign n537 = x54 ^ x22 ;
  assign n539 = x52 ^ x20 ;
  assign n541 = x50 ^ x18 ;
  assign n543 = x48 ^ x16 ;
  assign n545 = x46 ^ x14 ;
  assign n547 = x44 ^ x12 ;
  assign n549 = x42 ^ x10 ;
  assign n551 = x40 ^ x8 ;
  assign n553 = x38 ^ x6 ;
  assign n555 = x36 ^ x4 ;
  assign n557 = x34 ^ x2 ;
  assign n559 = x0 & ~x32 ;
  assign n560 = n559 ^ x34 ;
  assign n558 = x34 ^ x1 ;
  assign n561 = n560 ^ n558 ;
  assign n562 = x33 ^ x1 ;
  assign n563 = n561 & ~n562 ;
  assign n564 = n563 ^ n558 ;
  assign n565 = ~n557 & n564 ;
  assign n566 = n565 ^ x2 ;
  assign n567 = n566 ^ x36 ;
  assign n556 = x36 ^ x3 ;
  assign n568 = n567 ^ n556 ;
  assign n569 = x35 ^ x3 ;
  assign n570 = n568 & ~n569 ;
  assign n571 = n570 ^ n556 ;
  assign n572 = ~n555 & n571 ;
  assign n573 = n572 ^ x4 ;
  assign n574 = n573 ^ x38 ;
  assign n554 = x38 ^ x5 ;
  assign n575 = n574 ^ n554 ;
  assign n576 = x37 ^ x5 ;
  assign n577 = n575 & ~n576 ;
  assign n578 = n577 ^ n554 ;
  assign n579 = ~n553 & n578 ;
  assign n580 = n579 ^ x6 ;
  assign n581 = n580 ^ x40 ;
  assign n552 = x40 ^ x7 ;
  assign n582 = n581 ^ n552 ;
  assign n583 = x39 ^ x7 ;
  assign n584 = n582 & ~n583 ;
  assign n585 = n584 ^ n552 ;
  assign n586 = ~n551 & n585 ;
  assign n587 = n586 ^ x8 ;
  assign n588 = n587 ^ x42 ;
  assign n550 = x42 ^ x9 ;
  assign n589 = n588 ^ n550 ;
  assign n590 = x41 ^ x9 ;
  assign n591 = n589 & ~n590 ;
  assign n592 = n591 ^ n550 ;
  assign n593 = ~n549 & n592 ;
  assign n594 = n593 ^ x10 ;
  assign n595 = n594 ^ x44 ;
  assign n548 = x44 ^ x11 ;
  assign n596 = n595 ^ n548 ;
  assign n597 = x43 ^ x11 ;
  assign n598 = n596 & ~n597 ;
  assign n599 = n598 ^ n548 ;
  assign n600 = ~n547 & n599 ;
  assign n601 = n600 ^ x12 ;
  assign n602 = n601 ^ x46 ;
  assign n546 = x46 ^ x13 ;
  assign n603 = n602 ^ n546 ;
  assign n604 = x45 ^ x13 ;
  assign n605 = n603 & ~n604 ;
  assign n606 = n605 ^ n546 ;
  assign n607 = ~n545 & n606 ;
  assign n608 = n607 ^ x14 ;
  assign n609 = n608 ^ x48 ;
  assign n544 = x48 ^ x15 ;
  assign n610 = n609 ^ n544 ;
  assign n611 = x47 ^ x15 ;
  assign n612 = n610 & ~n611 ;
  assign n613 = n612 ^ n544 ;
  assign n614 = ~n543 & n613 ;
  assign n615 = n614 ^ x16 ;
  assign n616 = n615 ^ x50 ;
  assign n542 = x50 ^ x17 ;
  assign n617 = n616 ^ n542 ;
  assign n618 = x49 ^ x17 ;
  assign n619 = n617 & ~n618 ;
  assign n620 = n619 ^ n542 ;
  assign n621 = ~n541 & n620 ;
  assign n622 = n621 ^ x18 ;
  assign n623 = n622 ^ x52 ;
  assign n540 = x52 ^ x19 ;
  assign n624 = n623 ^ n540 ;
  assign n625 = x51 ^ x19 ;
  assign n626 = n624 & ~n625 ;
  assign n627 = n626 ^ n540 ;
  assign n628 = ~n539 & n627 ;
  assign n629 = n628 ^ x20 ;
  assign n630 = n629 ^ x54 ;
  assign n538 = x54 ^ x21 ;
  assign n631 = n630 ^ n538 ;
  assign n632 = x53 ^ x21 ;
  assign n633 = n631 & ~n632 ;
  assign n634 = n633 ^ n538 ;
  assign n635 = ~n537 & n634 ;
  assign n636 = n635 ^ x22 ;
  assign n637 = n636 ^ x56 ;
  assign n536 = x56 ^ x23 ;
  assign n638 = n637 ^ n536 ;
  assign n639 = x55 ^ x23 ;
  assign n640 = n638 & ~n639 ;
  assign n641 = n640 ^ n536 ;
  assign n642 = ~n535 & n641 ;
  assign n643 = n642 ^ x24 ;
  assign n644 = n643 ^ x58 ;
  assign n534 = x58 ^ x25 ;
  assign n645 = n644 ^ n534 ;
  assign n646 = x57 ^ x25 ;
  assign n647 = n645 & ~n646 ;
  assign n648 = n647 ^ n534 ;
  assign n649 = ~n533 & n648 ;
  assign n650 = n649 ^ x26 ;
  assign n651 = n650 ^ x60 ;
  assign n532 = x60 ^ x27 ;
  assign n652 = n651 ^ n532 ;
  assign n653 = x59 ^ x27 ;
  assign n654 = n652 & ~n653 ;
  assign n655 = n654 ^ n532 ;
  assign n656 = ~n531 & n655 ;
  assign n657 = n656 ^ x28 ;
  assign n658 = n657 ^ x62 ;
  assign n530 = x62 ^ x29 ;
  assign n659 = n658 ^ n530 ;
  assign n660 = x61 ^ x29 ;
  assign n661 = n659 & ~n660 ;
  assign n662 = n661 ^ n530 ;
  assign n663 = ~n528 & n662 ;
  assign n664 = n663 ^ x30 ;
  assign n665 = n664 ^ x63 ;
  assign n666 = ~n529 & n665 ;
  assign n667 = n666 ^ x31 ;
  assign n668 = n528 & ~n667 ;
  assign n669 = n668 ^ x30 ;
  assign n812 = n811 ^ n669 ;
  assign n813 = n521 ^ n520 ;
  assign n816 = n802 & ~n809 ;
  assign n817 = n816 ^ x93 ;
  assign n814 = n660 & ~n667 ;
  assign n815 = n814 ^ x29 ;
  assign n818 = n817 ^ n815 ;
  assign n821 = n673 & ~n809 ;
  assign n822 = n821 ^ x92 ;
  assign n819 = n531 & ~n667 ;
  assign n820 = n819 ^ x28 ;
  assign n823 = n822 ^ n820 ;
  assign n826 = n653 & ~n667 ;
  assign n827 = n826 ^ x27 ;
  assign n824 = n795 & ~n809 ;
  assign n825 = n824 ^ x91 ;
  assign n828 = n827 ^ n825 ;
  assign n831 = n675 & ~n809 ;
  assign n832 = n831 ^ x90 ;
  assign n829 = n533 & ~n667 ;
  assign n830 = n829 ^ x26 ;
  assign n833 = n832 ^ n830 ;
  assign n836 = n646 & ~n667 ;
  assign n837 = n836 ^ x25 ;
  assign n834 = n788 & ~n809 ;
  assign n835 = n834 ^ x89 ;
  assign n838 = n837 ^ n835 ;
  assign n841 = n677 & ~n809 ;
  assign n842 = n841 ^ x88 ;
  assign n839 = n535 & ~n667 ;
  assign n840 = n839 ^ x24 ;
  assign n843 = n842 ^ n840 ;
  assign n846 = n639 & ~n667 ;
  assign n847 = n846 ^ x23 ;
  assign n844 = n781 & ~n809 ;
  assign n845 = n844 ^ x87 ;
  assign n848 = n847 ^ n845 ;
  assign n851 = n679 & ~n809 ;
  assign n852 = n851 ^ x86 ;
  assign n849 = n537 & ~n667 ;
  assign n850 = n849 ^ x22 ;
  assign n853 = n852 ^ n850 ;
  assign n856 = n632 & ~n667 ;
  assign n857 = n856 ^ x21 ;
  assign n854 = n774 & ~n809 ;
  assign n855 = n854 ^ x85 ;
  assign n858 = n857 ^ n855 ;
  assign n861 = n681 & ~n809 ;
  assign n862 = n861 ^ x84 ;
  assign n859 = n539 & ~n667 ;
  assign n860 = n859 ^ x20 ;
  assign n863 = n862 ^ n860 ;
  assign n866 = n625 & ~n667 ;
  assign n867 = n866 ^ x19 ;
  assign n864 = n767 & ~n809 ;
  assign n865 = n864 ^ x83 ;
  assign n868 = n867 ^ n865 ;
  assign n871 = n683 & ~n809 ;
  assign n872 = n871 ^ x82 ;
  assign n869 = n541 & ~n667 ;
  assign n870 = n869 ^ x18 ;
  assign n873 = n872 ^ n870 ;
  assign n876 = n618 & ~n667 ;
  assign n877 = n876 ^ x17 ;
  assign n874 = n760 & ~n809 ;
  assign n875 = n874 ^ x81 ;
  assign n878 = n877 ^ n875 ;
  assign n881 = n685 & ~n809 ;
  assign n882 = n881 ^ x80 ;
  assign n879 = n543 & ~n667 ;
  assign n880 = n879 ^ x16 ;
  assign n883 = n882 ^ n880 ;
  assign n886 = n611 & ~n667 ;
  assign n887 = n886 ^ x15 ;
  assign n884 = n753 & ~n809 ;
  assign n885 = n884 ^ x79 ;
  assign n888 = n887 ^ n885 ;
  assign n891 = n687 & ~n809 ;
  assign n892 = n891 ^ x78 ;
  assign n889 = n545 & ~n667 ;
  assign n890 = n889 ^ x14 ;
  assign n893 = n892 ^ n890 ;
  assign n896 = n604 & ~n667 ;
  assign n897 = n896 ^ x13 ;
  assign n894 = n746 & ~n809 ;
  assign n895 = n894 ^ x77 ;
  assign n898 = n897 ^ n895 ;
  assign n901 = n689 & ~n809 ;
  assign n902 = n901 ^ x76 ;
  assign n899 = n547 & ~n667 ;
  assign n900 = n899 ^ x12 ;
  assign n903 = n902 ^ n900 ;
  assign n906 = n597 & ~n667 ;
  assign n907 = n906 ^ x11 ;
  assign n904 = n739 & ~n809 ;
  assign n905 = n904 ^ x75 ;
  assign n908 = n907 ^ n905 ;
  assign n911 = n691 & ~n809 ;
  assign n912 = n911 ^ x74 ;
  assign n909 = n549 & ~n667 ;
  assign n910 = n909 ^ x10 ;
  assign n913 = n912 ^ n910 ;
  assign n916 = n590 & ~n667 ;
  assign n917 = n916 ^ x9 ;
  assign n914 = n732 & ~n809 ;
  assign n915 = n914 ^ x73 ;
  assign n918 = n917 ^ n915 ;
  assign n921 = n693 & ~n809 ;
  assign n922 = n921 ^ x72 ;
  assign n919 = n551 & ~n667 ;
  assign n920 = n919 ^ x8 ;
  assign n923 = n922 ^ n920 ;
  assign n926 = n583 & ~n667 ;
  assign n927 = n926 ^ x7 ;
  assign n924 = n725 & ~n809 ;
  assign n925 = n924 ^ x71 ;
  assign n928 = n927 ^ n925 ;
  assign n931 = n553 & ~n667 ;
  assign n932 = n931 ^ x6 ;
  assign n929 = n695 & ~n809 ;
  assign n930 = n929 ^ x70 ;
  assign n933 = n932 ^ n930 ;
  assign n936 = n576 & ~n667 ;
  assign n937 = n936 ^ x5 ;
  assign n934 = n718 & ~n809 ;
  assign n935 = n934 ^ x69 ;
  assign n938 = n937 ^ n935 ;
  assign n941 = n555 & ~n667 ;
  assign n942 = n941 ^ x4 ;
  assign n939 = n697 & ~n809 ;
  assign n940 = n939 ^ x68 ;
  assign n943 = n942 ^ n940 ;
  assign n946 = n569 & ~n667 ;
  assign n947 = n946 ^ x3 ;
  assign n944 = n711 & ~n809 ;
  assign n945 = n944 ^ x67 ;
  assign n948 = n947 ^ n945 ;
  assign n951 = n557 & ~n667 ;
  assign n952 = n951 ^ x2 ;
  assign n949 = n699 & ~n809 ;
  assign n950 = n949 ^ x66 ;
  assign n953 = n952 ^ n950 ;
  assign n956 = n704 & ~n809 ;
  assign n957 = n956 ^ x65 ;
  assign n954 = n562 & ~n667 ;
  assign n955 = n954 ^ x1 ;
  assign n958 = n957 ^ n955 ;
  assign n959 = x32 ^ x0 ;
  assign n960 = ~n667 & n959 ;
  assign n961 = n960 ^ x0 ;
  assign n962 = x96 ^ x64 ;
  assign n963 = ~n809 & n962 ;
  assign n964 = n963 ^ x64 ;
  assign n965 = n961 & ~n964 ;
  assign n966 = n965 ^ n957 ;
  assign n967 = ~n958 & ~n966 ;
  assign n968 = n967 ^ n957 ;
  assign n969 = n968 ^ n952 ;
  assign n970 = ~n953 & ~n969 ;
  assign n971 = n970 ^ n952 ;
  assign n972 = n971 ^ n947 ;
  assign n973 = ~n948 & n972 ;
  assign n974 = n973 ^ n947 ;
  assign n975 = n974 ^ n940 ;
  assign n976 = ~n943 & ~n975 ;
  assign n977 = n976 ^ n940 ;
  assign n978 = n977 ^ n937 ;
  assign n979 = ~n938 & ~n978 ;
  assign n980 = n979 ^ n937 ;
  assign n981 = n980 ^ n930 ;
  assign n982 = ~n933 & ~n981 ;
  assign n983 = n982 ^ n930 ;
  assign n984 = n983 ^ n927 ;
  assign n985 = ~n928 & ~n984 ;
  assign n986 = n985 ^ n927 ;
  assign n987 = n986 ^ n920 ;
  assign n988 = ~n923 & n987 ;
  assign n989 = n988 ^ n920 ;
  assign n990 = n989 ^ n917 ;
  assign n991 = ~n918 & n990 ;
  assign n992 = n991 ^ n917 ;
  assign n993 = n992 ^ n910 ;
  assign n994 = ~n913 & n993 ;
  assign n995 = n994 ^ n910 ;
  assign n996 = n995 ^ n907 ;
  assign n997 = ~n908 & n996 ;
  assign n998 = n997 ^ n907 ;
  assign n999 = n998 ^ n900 ;
  assign n1000 = ~n903 & n999 ;
  assign n1001 = n1000 ^ n900 ;
  assign n1002 = n1001 ^ n897 ;
  assign n1003 = ~n898 & n1002 ;
  assign n1004 = n1003 ^ n897 ;
  assign n1005 = n1004 ^ n890 ;
  assign n1006 = ~n893 & n1005 ;
  assign n1007 = n1006 ^ n890 ;
  assign n1008 = n1007 ^ n887 ;
  assign n1009 = ~n888 & n1008 ;
  assign n1010 = n1009 ^ n887 ;
  assign n1011 = n1010 ^ n880 ;
  assign n1012 = ~n883 & n1011 ;
  assign n1013 = n1012 ^ n880 ;
  assign n1014 = n1013 ^ n877 ;
  assign n1015 = ~n878 & n1014 ;
  assign n1016 = n1015 ^ n877 ;
  assign n1017 = n1016 ^ n870 ;
  assign n1018 = ~n873 & n1017 ;
  assign n1019 = n1018 ^ n870 ;
  assign n1020 = n1019 ^ n867 ;
  assign n1021 = ~n868 & n1020 ;
  assign n1022 = n1021 ^ n867 ;
  assign n1023 = n1022 ^ n860 ;
  assign n1024 = ~n863 & n1023 ;
  assign n1025 = n1024 ^ n860 ;
  assign n1026 = n1025 ^ n857 ;
  assign n1027 = ~n858 & n1026 ;
  assign n1028 = n1027 ^ n857 ;
  assign n1029 = n1028 ^ n850 ;
  assign n1030 = ~n853 & n1029 ;
  assign n1031 = n1030 ^ n850 ;
  assign n1032 = n1031 ^ n847 ;
  assign n1033 = ~n848 & n1032 ;
  assign n1034 = n1033 ^ n847 ;
  assign n1035 = n1034 ^ n840 ;
  assign n1036 = ~n843 & n1035 ;
  assign n1037 = n1036 ^ n840 ;
  assign n1038 = n1037 ^ n837 ;
  assign n1039 = ~n838 & n1038 ;
  assign n1040 = n1039 ^ n837 ;
  assign n1041 = n1040 ^ n830 ;
  assign n1042 = ~n833 & n1041 ;
  assign n1043 = n1042 ^ n830 ;
  assign n1044 = n1043 ^ n827 ;
  assign n1045 = ~n828 & n1044 ;
  assign n1046 = n1045 ^ n827 ;
  assign n1047 = n1046 ^ n822 ;
  assign n1048 = ~n823 & ~n1047 ;
  assign n1049 = n1048 ^ n822 ;
  assign n1050 = n1049 ^ n817 ;
  assign n1051 = ~n818 & ~n1050 ;
  assign n1052 = n1051 ^ n815 ;
  assign n1053 = n1052 ^ n811 ;
  assign n1054 = ~n812 & n1053 ;
  assign n1055 = n1054 ^ n669 ;
  assign n1056 = n1055 ^ n521 ;
  assign n1057 = ~n813 & ~n1056 ;
  assign n1058 = n1057 ^ n520 ;
  assign n1059 = n812 & n1058 ;
  assign n1060 = n1059 ^ n669 ;
  assign n1594 = n1593 ^ n1060 ;
  assign n1595 = n525 ^ n522 ;
  assign n1598 = n1351 & ~n1591 ;
  assign n1599 = n1598 ^ n1350 ;
  assign n1596 = n818 & ~n1058 ;
  assign n1597 = n1596 ^ n817 ;
  assign n1600 = n1599 ^ n1597 ;
  assign n1603 = n823 & ~n1058 ;
  assign n1604 = n1603 ^ n822 ;
  assign n1601 = n1356 & ~n1591 ;
  assign n1602 = n1601 ^ n1355 ;
  assign n1605 = n1604 ^ n1602 ;
  assign n1608 = n828 & n1058 ;
  assign n1609 = n1608 ^ n827 ;
  assign n1606 = n1361 & n1591 ;
  assign n1607 = n1606 ^ n1360 ;
  assign n1610 = n1609 ^ n1607 ;
  assign n1613 = n833 & n1058 ;
  assign n1614 = n1613 ^ n830 ;
  assign n1611 = n1366 & n1591 ;
  assign n1612 = n1611 ^ n1363 ;
  assign n1615 = n1614 ^ n1612 ;
  assign n1618 = n838 & ~n1058 ;
  assign n1619 = n1618 ^ n835 ;
  assign n1616 = n1371 & ~n1591 ;
  assign n1617 = n1616 ^ n1368 ;
  assign n1620 = n1619 ^ n1617 ;
  assign n1623 = n1376 & ~n1591 ;
  assign n1624 = n1623 ^ n1375 ;
  assign n1621 = n843 & ~n1058 ;
  assign n1622 = n1621 ^ n842 ;
  assign n1625 = n1624 ^ n1622 ;
  assign n1628 = n848 & n1058 ;
  assign n1629 = n1628 ^ n847 ;
  assign n1626 = n1381 & n1591 ;
  assign n1627 = n1626 ^ n1380 ;
  assign n1630 = n1629 ^ n1627 ;
  assign n1633 = n853 & n1058 ;
  assign n1634 = n1633 ^ n850 ;
  assign n1631 = n1386 & n1591 ;
  assign n1632 = n1631 ^ n1383 ;
  assign n1635 = n1634 ^ n1632 ;
  assign n1638 = n1391 & ~n1591 ;
  assign n1639 = n1638 ^ n1388 ;
  assign n1636 = n858 & ~n1058 ;
  assign n1637 = n1636 ^ n855 ;
  assign n1640 = n1639 ^ n1637 ;
  assign n1643 = n1396 & ~n1591 ;
  assign n1644 = n1643 ^ n1395 ;
  assign n1641 = n863 & ~n1058 ;
  assign n1642 = n1641 ^ n862 ;
  assign n1645 = n1644 ^ n1642 ;
  assign n1648 = n868 & n1058 ;
  assign n1649 = n1648 ^ n867 ;
  assign n1646 = n1401 & n1591 ;
  assign n1647 = n1646 ^ n1400 ;
  assign n1650 = n1649 ^ n1647 ;
  assign n1653 = n873 & n1058 ;
  assign n1654 = n1653 ^ n870 ;
  assign n1651 = n1406 & n1591 ;
  assign n1652 = n1651 ^ n1403 ;
  assign n1655 = n1654 ^ n1652 ;
  assign n1658 = n1411 & ~n1591 ;
  assign n1659 = n1658 ^ n1408 ;
  assign n1656 = n878 & ~n1058 ;
  assign n1657 = n1656 ^ n875 ;
  assign n1660 = n1659 ^ n1657 ;
  assign n1663 = n1416 & ~n1591 ;
  assign n1664 = n1663 ^ n1415 ;
  assign n1661 = n883 & ~n1058 ;
  assign n1662 = n1661 ^ n882 ;
  assign n1665 = n1664 ^ n1662 ;
  assign n1668 = n888 & n1058 ;
  assign n1669 = n1668 ^ n887 ;
  assign n1666 = n1421 & n1591 ;
  assign n1667 = n1666 ^ n1420 ;
  assign n1670 = n1669 ^ n1667 ;
  assign n1673 = n893 & n1058 ;
  assign n1674 = n1673 ^ n890 ;
  assign n1671 = n1426 & n1591 ;
  assign n1672 = n1671 ^ n1423 ;
  assign n1675 = n1674 ^ n1672 ;
  assign n1678 = n1431 & ~n1591 ;
  assign n1679 = n1678 ^ n1428 ;
  assign n1676 = n898 & ~n1058 ;
  assign n1677 = n1676 ^ n895 ;
  assign n1680 = n1679 ^ n1677 ;
  assign n1683 = n1436 & ~n1591 ;
  assign n1684 = n1683 ^ n1435 ;
  assign n1681 = n903 & ~n1058 ;
  assign n1682 = n1681 ^ n902 ;
  assign n1685 = n1684 ^ n1682 ;
  assign n1688 = n908 & n1058 ;
  assign n1689 = n1688 ^ n907 ;
  assign n1686 = n1441 & n1591 ;
  assign n1687 = n1686 ^ n1440 ;
  assign n1690 = n1689 ^ n1687 ;
  assign n1693 = n913 & n1058 ;
  assign n1694 = n1693 ^ n910 ;
  assign n1691 = n1446 & n1591 ;
  assign n1692 = n1691 ^ n1443 ;
  assign n1695 = n1694 ^ n1692 ;
  assign n1698 = n1451 & ~n1591 ;
  assign n1699 = n1698 ^ n1448 ;
  assign n1696 = n918 & ~n1058 ;
  assign n1697 = n1696 ^ n915 ;
  assign n1700 = n1699 ^ n1697 ;
  assign n1703 = n1456 & ~n1591 ;
  assign n1704 = n1703 ^ n1455 ;
  assign n1701 = n923 & ~n1058 ;
  assign n1702 = n1701 ^ n922 ;
  assign n1705 = n1704 ^ n1702 ;
  assign n1708 = n928 & n1058 ;
  assign n1709 = n1708 ^ n927 ;
  assign n1706 = n1461 & n1591 ;
  assign n1707 = n1706 ^ n1460 ;
  assign n1710 = n1709 ^ n1707 ;
  assign n1713 = n933 & ~n1058 ;
  assign n1714 = n1713 ^ n930 ;
  assign n1711 = n1466 & n1591 ;
  assign n1712 = n1711 ^ n1463 ;
  assign n1715 = n1714 ^ n1712 ;
  assign n1718 = n1471 & ~n1591 ;
  assign n1719 = n1718 ^ n1468 ;
  assign n1716 = n938 & ~n1058 ;
  assign n1717 = n1716 ^ n935 ;
  assign n1720 = n1719 ^ n1717 ;
  assign n1723 = n943 & n1058 ;
  assign n1724 = n1723 ^ n942 ;
  assign n1721 = n1476 & ~n1591 ;
  assign n1722 = n1721 ^ n1475 ;
  assign n1725 = n1724 ^ n1722 ;
  assign n1728 = n948 & n1058 ;
  assign n1729 = n1728 ^ n947 ;
  assign n1726 = n1481 & ~n1591 ;
  assign n1727 = n1726 ^ n1480 ;
  assign n1730 = n1729 ^ n1727 ;
  assign n1733 = n953 & ~n1058 ;
  assign n1734 = n1733 ^ n950 ;
  assign n1731 = n1486 & ~n1591 ;
  assign n1732 = n1731 ^ n1483 ;
  assign n1735 = n1734 ^ n1732 ;
  assign n1738 = n1491 & n1591 ;
  assign n1739 = n1738 ^ n1488 ;
  assign n1736 = n958 & n1058 ;
  assign n1737 = n1736 ^ n955 ;
  assign n1740 = n1739 ^ n1737 ;
  assign n1741 = n1497 ^ n1494 ;
  assign n1742 = ~n1591 & n1741 ;
  assign n1743 = n1742 ^ n1494 ;
  assign n1744 = n964 ^ n961 ;
  assign n1745 = n1058 & n1744 ;
  assign n1746 = n1745 ^ n961 ;
  assign n1747 = ~n1743 & n1746 ;
  assign n1748 = n1747 ^ n1739 ;
  assign n1749 = ~n1740 & ~n1748 ;
  assign n1750 = n1749 ^ n1739 ;
  assign n1751 = n1750 ^ n1732 ;
  assign n1752 = ~n1735 & n1751 ;
  assign n1753 = n1752 ^ n1732 ;
  assign n1754 = n1753 ^ n1729 ;
  assign n1755 = ~n1730 & ~n1754 ;
  assign n1756 = n1755 ^ n1729 ;
  assign n1757 = n1756 ^ n1722 ;
  assign n1758 = ~n1725 & ~n1757 ;
  assign n1759 = n1758 ^ n1722 ;
  assign n1760 = n1759 ^ n1719 ;
  assign n1761 = ~n1720 & n1760 ;
  assign n1762 = n1761 ^ n1719 ;
  assign n1763 = n1762 ^ n1712 ;
  assign n1764 = ~n1715 & n1763 ;
  assign n1765 = n1764 ^ n1712 ;
  assign n1766 = n1765 ^ n1709 ;
  assign n1767 = ~n1710 & ~n1766 ;
  assign n1768 = n1767 ^ n1709 ;
  assign n1769 = n1768 ^ n1702 ;
  assign n1770 = ~n1705 & n1769 ;
  assign n1771 = n1770 ^ n1702 ;
  assign n1772 = n1771 ^ n1699 ;
  assign n1773 = ~n1700 & ~n1772 ;
  assign n1774 = n1773 ^ n1699 ;
  assign n1775 = n1774 ^ n1692 ;
  assign n1776 = ~n1695 & n1775 ;
  assign n1777 = n1776 ^ n1692 ;
  assign n1778 = n1777 ^ n1689 ;
  assign n1779 = ~n1690 & ~n1778 ;
  assign n1780 = n1779 ^ n1689 ;
  assign n1781 = n1780 ^ n1682 ;
  assign n1782 = ~n1685 & n1781 ;
  assign n1783 = n1782 ^ n1682 ;
  assign n1784 = n1783 ^ n1679 ;
  assign n1785 = ~n1680 & ~n1784 ;
  assign n1786 = n1785 ^ n1679 ;
  assign n1787 = n1786 ^ n1672 ;
  assign n1788 = ~n1675 & n1787 ;
  assign n1789 = n1788 ^ n1672 ;
  assign n1790 = n1789 ^ n1669 ;
  assign n1791 = ~n1670 & ~n1790 ;
  assign n1792 = n1791 ^ n1669 ;
  assign n1793 = n1792 ^ n1662 ;
  assign n1794 = ~n1665 & n1793 ;
  assign n1795 = n1794 ^ n1662 ;
  assign n1796 = n1795 ^ n1659 ;
  assign n1797 = ~n1660 & ~n1796 ;
  assign n1798 = n1797 ^ n1659 ;
  assign n1799 = n1798 ^ n1652 ;
  assign n1800 = ~n1655 & n1799 ;
  assign n1801 = n1800 ^ n1652 ;
  assign n1802 = n1801 ^ n1649 ;
  assign n1803 = ~n1650 & ~n1802 ;
  assign n1804 = n1803 ^ n1649 ;
  assign n1805 = n1804 ^ n1642 ;
  assign n1806 = ~n1645 & n1805 ;
  assign n1807 = n1806 ^ n1642 ;
  assign n1808 = n1807 ^ n1639 ;
  assign n1809 = ~n1640 & ~n1808 ;
  assign n1810 = n1809 ^ n1639 ;
  assign n1811 = n1810 ^ n1632 ;
  assign n1812 = ~n1635 & n1811 ;
  assign n1813 = n1812 ^ n1632 ;
  assign n1814 = n1813 ^ n1629 ;
  assign n1815 = ~n1630 & ~n1814 ;
  assign n1816 = n1815 ^ n1629 ;
  assign n1817 = n1816 ^ n1622 ;
  assign n1818 = ~n1625 & n1817 ;
  assign n1819 = n1818 ^ n1622 ;
  assign n1820 = n1819 ^ n1619 ;
  assign n1821 = ~n1620 & n1820 ;
  assign n1822 = n1821 ^ n1619 ;
  assign n1823 = n1822 ^ n1612 ;
  assign n1824 = ~n1615 & ~n1823 ;
  assign n1825 = n1824 ^ n1612 ;
  assign n1826 = n1825 ^ n1609 ;
  assign n1827 = ~n1610 & ~n1826 ;
  assign n1828 = n1827 ^ n1609 ;
  assign n1829 = n1828 ^ n1602 ;
  assign n1830 = ~n1605 & ~n1829 ;
  assign n1831 = n1830 ^ n1602 ;
  assign n1832 = n1831 ^ n1597 ;
  assign n1833 = ~n1600 & ~n1832 ;
  assign n1834 = n1833 ^ n1597 ;
  assign n1835 = n1834 ^ n1060 ;
  assign n1836 = ~n1594 & ~n1835 ;
  assign n1837 = n1836 ^ n1593 ;
  assign n1838 = n1837 ^ n525 ;
  assign n1839 = ~n1595 & n1838 ;
  assign n1840 = n1839 ^ n522 ;
  assign n1841 = n1594 & n1840 ;
  assign n1842 = n1841 ^ n1060 ;
  assign n3158 = n3157 ^ n1842 ;
  assign n3161 = n1600 & n1840 ;
  assign n3162 = n3161 ^ n1597 ;
  assign n3159 = n2915 & n3155 ;
  assign n3160 = n3159 ^ n2912 ;
  assign n3163 = n3162 ^ n3160 ;
  assign n3166 = n1605 & n1840 ;
  assign n3167 = n3166 ^ n1604 ;
  assign n3164 = n2920 & n3155 ;
  assign n3165 = n3164 ^ n2919 ;
  assign n3168 = n3167 ^ n3165 ;
  assign n3171 = n2925 & n3155 ;
  assign n3172 = n3171 ^ n2924 ;
  assign n3169 = n1610 & n1840 ;
  assign n3170 = n3169 ^ n1609 ;
  assign n3173 = n3172 ^ n3170 ;
  assign n3176 = n1615 & ~n1840 ;
  assign n3177 = n3176 ^ n1612 ;
  assign n3174 = n2930 & ~n3155 ;
  assign n3175 = n3174 ^ n2927 ;
  assign n3178 = n3177 ^ n3175 ;
  assign n3181 = n2935 & ~n3155 ;
  assign n3182 = n3181 ^ n2932 ;
  assign n3179 = n1620 & ~n1840 ;
  assign n3180 = n3179 ^ n1617 ;
  assign n3183 = n3182 ^ n3180 ;
  assign n3186 = n1625 & ~n1840 ;
  assign n3187 = n3186 ^ n1624 ;
  assign n3184 = n2940 & ~n3155 ;
  assign n3185 = n3184 ^ n2939 ;
  assign n3188 = n3187 ^ n3185 ;
  assign n3372 = n1630 & n1840 ;
  assign n3373 = n3372 ^ n1629 ;
  assign n3191 = n1635 & ~n1840 ;
  assign n3192 = n3191 ^ n1632 ;
  assign n3189 = n2950 & ~n3155 ;
  assign n3190 = n3189 ^ n2947 ;
  assign n3193 = n3192 ^ n3190 ;
  assign n3196 = n2955 & n3155 ;
  assign n3197 = n3196 ^ n2952 ;
  assign n3194 = n1640 & n1840 ;
  assign n3195 = n3194 ^ n1637 ;
  assign n3198 = n3197 ^ n3195 ;
  assign n3201 = n2960 & ~n3155 ;
  assign n3202 = n3201 ^ n2959 ;
  assign n3199 = n1645 & ~n1840 ;
  assign n3200 = n3199 ^ n1644 ;
  assign n3203 = n3202 ^ n3200 ;
  assign n3355 = n1650 & n1840 ;
  assign n3356 = n3355 ^ n1649 ;
  assign n3206 = n1655 & ~n1840 ;
  assign n3207 = n3206 ^ n1652 ;
  assign n3204 = n2970 & ~n3155 ;
  assign n3205 = n3204 ^ n2967 ;
  assign n3208 = n3207 ^ n3205 ;
  assign n3211 = n1660 & n1840 ;
  assign n3212 = n3211 ^ n1657 ;
  assign n3209 = n2975 & n3155 ;
  assign n3210 = n3209 ^ n2972 ;
  assign n3213 = n3212 ^ n3210 ;
  assign n3216 = n2980 & ~n3155 ;
  assign n3217 = n3216 ^ n2979 ;
  assign n3214 = n1665 & ~n1840 ;
  assign n3215 = n3214 ^ n1664 ;
  assign n3218 = n3217 ^ n3215 ;
  assign n3338 = n1670 & n1840 ;
  assign n3339 = n3338 ^ n1669 ;
  assign n3221 = n1675 & ~n1840 ;
  assign n3222 = n3221 ^ n1672 ;
  assign n3219 = n2990 & ~n3155 ;
  assign n3220 = n3219 ^ n2987 ;
  assign n3223 = n3222 ^ n3220 ;
  assign n3226 = n1680 & n1840 ;
  assign n3227 = n3226 ^ n1677 ;
  assign n3224 = n2995 & n3155 ;
  assign n3225 = n3224 ^ n2992 ;
  assign n3228 = n3227 ^ n3225 ;
  assign n3231 = n3000 & ~n3155 ;
  assign n3232 = n3231 ^ n2999 ;
  assign n3229 = n1685 & ~n1840 ;
  assign n3230 = n3229 ^ n1684 ;
  assign n3233 = n3232 ^ n3230 ;
  assign n3321 = n1690 & n1840 ;
  assign n3322 = n3321 ^ n1689 ;
  assign n3236 = n1695 & ~n1840 ;
  assign n3237 = n3236 ^ n1692 ;
  assign n3234 = n3010 & ~n3155 ;
  assign n3235 = n3234 ^ n3007 ;
  assign n3238 = n3237 ^ n3235 ;
  assign n3241 = n3015 & n3155 ;
  assign n3242 = n3241 ^ n3012 ;
  assign n3239 = n1700 & n1840 ;
  assign n3240 = n3239 ^ n1697 ;
  assign n3243 = n3242 ^ n3240 ;
  assign n3246 = n3020 & ~n3155 ;
  assign n3247 = n3246 ^ n3019 ;
  assign n3244 = n1705 & ~n1840 ;
  assign n3245 = n3244 ^ n1704 ;
  assign n3248 = n3247 ^ n3245 ;
  assign n3251 = n3025 & n3155 ;
  assign n3252 = n3251 ^ n3024 ;
  assign n3249 = n1710 & n1840 ;
  assign n3250 = n3249 ^ n1709 ;
  assign n3253 = n3252 ^ n3250 ;
  assign n3256 = n1715 & ~n1840 ;
  assign n3257 = n3256 ^ n1712 ;
  assign n3254 = n3030 & ~n3155 ;
  assign n3255 = n3254 ^ n3027 ;
  assign n3258 = n3257 ^ n3255 ;
  assign n3261 = n3035 & n3155 ;
  assign n3262 = n3261 ^ n3032 ;
  assign n3259 = n1720 & n1840 ;
  assign n3260 = n3259 ^ n1717 ;
  assign n3263 = n3262 ^ n3260 ;
  assign n3266 = n1725 & n1840 ;
  assign n3267 = n3266 ^ n1724 ;
  assign n3264 = n3040 & ~n3155 ;
  assign n3265 = n3264 ^ n3039 ;
  assign n3268 = n3267 ^ n3265 ;
  assign n3271 = n1730 & n1840 ;
  assign n3272 = n3271 ^ n1729 ;
  assign n3299 = n3272 ^ n3267 ;
  assign n3269 = n3045 & ~n3155 ;
  assign n3270 = n3269 ^ n3044 ;
  assign n3273 = n3272 ^ n3270 ;
  assign n3276 = n1735 & ~n1840 ;
  assign n3277 = n3276 ^ n1732 ;
  assign n3274 = n3050 & ~n3155 ;
  assign n3275 = n3274 ^ n3047 ;
  assign n3278 = n3277 ^ n3275 ;
  assign n3281 = n3055 & n3155 ;
  assign n3282 = n3281 ^ n3052 ;
  assign n3279 = n1740 & n1840 ;
  assign n3280 = n3279 ^ n1737 ;
  assign n3283 = n3282 ^ n3280 ;
  assign n3284 = n3061 ^ n3058 ;
  assign n3285 = ~n3155 & n3284 ;
  assign n3286 = n3285 ^ n3058 ;
  assign n3287 = n1746 ^ n1743 ;
  assign n3288 = ~n1840 & n3287 ;
  assign n3289 = n3288 ^ n1743 ;
  assign n3290 = ~n3286 & n3289 ;
  assign n3291 = n3290 ^ n3282 ;
  assign n3292 = ~n3283 & ~n3291 ;
  assign n3293 = n3292 ^ n3282 ;
  assign n3294 = n3293 ^ n3277 ;
  assign n3295 = ~n3278 & ~n3294 ;
  assign n3296 = n3295 ^ n3277 ;
  assign n3297 = n3296 ^ n3270 ;
  assign n3298 = ~n3273 & n3297 ;
  assign n3300 = n3299 ^ n3298 ;
  assign n3301 = ~n3268 & ~n3300 ;
  assign n3302 = n3301 ^ n3265 ;
  assign n3303 = n3302 ^ n3262 ;
  assign n3304 = ~n3263 & ~n3303 ;
  assign n3305 = n3304 ^ n3260 ;
  assign n3306 = n3305 ^ n3257 ;
  assign n3307 = ~n3258 & n3306 ;
  assign n3308 = n3307 ^ n3257 ;
  assign n3309 = n3308 ^ n3250 ;
  assign n3310 = ~n3253 & n3309 ;
  assign n3311 = n3310 ^ n3250 ;
  assign n3312 = n3311 ^ n3245 ;
  assign n3313 = ~n3248 & n3312 ;
  assign n3314 = n3313 ^ n3245 ;
  assign n3315 = n3314 ^ n3242 ;
  assign n3316 = ~n3243 & n3315 ;
  assign n3317 = n3316 ^ n3240 ;
  assign n3318 = n3317 ^ n3237 ;
  assign n3319 = ~n3238 & ~n3318 ;
  assign n3320 = n3319 ^ n3235 ;
  assign n3323 = n3322 ^ n3320 ;
  assign n3324 = n3005 & n3155 ;
  assign n3325 = n3324 ^ n3004 ;
  assign n3326 = n3325 ^ n3320 ;
  assign n3327 = ~n3323 & n3326 ;
  assign n3328 = n3327 ^ n3320 ;
  assign n3329 = n3328 ^ n3232 ;
  assign n3330 = ~n3233 & n3329 ;
  assign n3331 = n3330 ^ n3232 ;
  assign n3332 = n3331 ^ n3225 ;
  assign n3333 = ~n3228 & ~n3332 ;
  assign n3334 = n3333 ^ n3227 ;
  assign n3335 = n3334 ^ n3222 ;
  assign n3336 = ~n3223 & ~n3335 ;
  assign n3337 = n3336 ^ n3220 ;
  assign n3340 = n3339 ^ n3337 ;
  assign n3341 = n2985 & n3155 ;
  assign n3342 = n3341 ^ n2984 ;
  assign n3343 = n3342 ^ n3337 ;
  assign n3344 = ~n3340 & n3343 ;
  assign n3345 = n3344 ^ n3337 ;
  assign n3346 = n3345 ^ n3217 ;
  assign n3347 = ~n3218 & n3346 ;
  assign n3348 = n3347 ^ n3217 ;
  assign n3349 = n3348 ^ n3212 ;
  assign n3350 = ~n3213 & n3349 ;
  assign n3351 = n3350 ^ n3210 ;
  assign n3352 = n3351 ^ n3207 ;
  assign n3353 = ~n3208 & n3352 ;
  assign n3354 = n3353 ^ n3205 ;
  assign n3357 = n3356 ^ n3354 ;
  assign n3358 = n2965 & n3155 ;
  assign n3359 = n3358 ^ n2964 ;
  assign n3360 = n3359 ^ n3354 ;
  assign n3361 = ~n3357 & n3360 ;
  assign n3362 = n3361 ^ n3354 ;
  assign n3363 = n3362 ^ n3202 ;
  assign n3364 = ~n3203 & n3363 ;
  assign n3365 = n3364 ^ n3202 ;
  assign n3366 = n3365 ^ n3195 ;
  assign n3367 = ~n3198 & n3366 ;
  assign n3368 = n3367 ^ n3197 ;
  assign n3369 = n3368 ^ n3192 ;
  assign n3370 = ~n3193 & n3369 ;
  assign n3371 = n3370 ^ n3190 ;
  assign n3374 = n3373 ^ n3371 ;
  assign n3375 = n2945 & n3155 ;
  assign n3376 = n3375 ^ n2944 ;
  assign n3377 = n3376 ^ n3371 ;
  assign n3378 = ~n3374 & n3377 ;
  assign n3379 = n3378 ^ n3371 ;
  assign n3380 = n3379 ^ n3185 ;
  assign n3381 = ~n3188 & ~n3380 ;
  assign n3382 = n3381 ^ n3187 ;
  assign n3383 = n3382 ^ n3182 ;
  assign n3384 = ~n3183 & n3383 ;
  assign n3385 = n3384 ^ n3180 ;
  assign n3386 = n3385 ^ n3177 ;
  assign n3387 = ~n3178 & ~n3386 ;
  assign n3388 = n3387 ^ n3175 ;
  assign n3389 = n3388 ^ n3172 ;
  assign n3390 = ~n3173 & n3389 ;
  assign n3391 = n3390 ^ n3172 ;
  assign n3392 = n3391 ^ n3165 ;
  assign n3393 = ~n3168 & n3392 ;
  assign n3394 = n3393 ^ n3165 ;
  assign n3395 = n3394 ^ n3160 ;
  assign n3396 = ~n3163 & n3395 ;
  assign n3397 = n3396 ^ n3160 ;
  assign n3398 = n3397 ^ n1842 ;
  assign n3399 = ~n3158 & n3398 ;
  assign n3400 = n3399 ^ n3157 ;
  assign n3401 = n3400 ^ n526 ;
  assign n3402 = ~n527 & ~n3401 ;
  assign n3403 = n3402 ^ n519 ;
  assign n3404 = n3155 ^ n1840 ;
  assign n3405 = ~n3403 & n3404 ;
  assign n3406 = n3405 ^ n1840 ;
  assign n3410 = n1058 & ~n3406 ;
  assign n3411 = n1591 & n1840 ;
  assign n3412 = ~n3410 & ~n3411 ;
  assign n3407 = n2373 & ~n3406 ;
  assign n3408 = n2906 & n3155 ;
  assign n3409 = ~n3407 & ~n3408 ;
  assign n3413 = n3412 ^ n3409 ;
  assign n3414 = n3403 & n3413 ;
  assign n3415 = n3414 ^ n3409 ;
  assign n3428 = n809 ^ n667 ;
  assign n3429 = n3415 & n3428 ;
  assign n3430 = n3429 ^ n809 ;
  assign n3425 = n1342 ^ n1200 ;
  assign n3426 = n3415 & n3425 ;
  assign n3427 = n3426 ^ n1200 ;
  assign n3431 = n3430 ^ n3427 ;
  assign n3432 = n3406 & n3431 ;
  assign n3433 = n3432 ^ n3430 ;
  assign n3419 = n2124 ^ n1982 ;
  assign n3420 = n3415 & n3419 ;
  assign n3421 = n3420 ^ n2124 ;
  assign n3416 = n2657 ^ n2515 ;
  assign n3417 = n3415 & n3416 ;
  assign n3418 = n3417 ^ n2515 ;
  assign n3422 = n3421 ^ n3418 ;
  assign n3423 = n3406 & n3422 ;
  assign n3424 = n3423 ^ n3421 ;
  assign n3434 = n3433 ^ n3424 ;
  assign n3435 = n3403 & n3434 ;
  assign n3436 = n3435 ^ n3424 ;
  assign n3437 = n3289 ^ n3286 ;
  assign n3438 = n3403 & n3437 ;
  assign n3439 = n3438 ^ n3286 ;
  assign n3440 = n3283 & ~n3403 ;
  assign n3441 = n3440 ^ n3280 ;
  assign n3442 = n3278 & n3403 ;
  assign n3443 = n3442 ^ n3275 ;
  assign n3444 = n3273 & n3403 ;
  assign n3445 = n3444 ^ n3270 ;
  assign n3446 = n3268 & n3403 ;
  assign n3447 = n3446 ^ n3265 ;
  assign n3448 = n3263 & ~n3403 ;
  assign n3449 = n3448 ^ n3260 ;
  assign n3450 = n3258 & n3403 ;
  assign n3451 = n3450 ^ n3255 ;
  assign n3452 = n3253 & ~n3403 ;
  assign n3453 = n3452 ^ n3250 ;
  assign n3454 = n3248 & n3403 ;
  assign n3455 = n3454 ^ n3247 ;
  assign n3456 = n3243 & ~n3403 ;
  assign n3457 = n3456 ^ n3240 ;
  assign n3458 = n3238 & n3403 ;
  assign n3459 = n3458 ^ n3235 ;
  assign n3460 = n3325 ^ n3322 ;
  assign n3461 = n3403 & n3460 ;
  assign n3462 = n3461 ^ n3325 ;
  assign n3463 = n3233 & ~n3403 ;
  assign n3464 = n3463 ^ n3230 ;
  assign n3465 = n3228 & ~n3403 ;
  assign n3466 = n3465 ^ n3227 ;
  assign n3467 = n3223 & n3403 ;
  assign n3468 = n3467 ^ n3220 ;
  assign n3469 = n3342 ^ n3339 ;
  assign n3470 = n3403 & n3469 ;
  assign n3471 = n3470 ^ n3342 ;
  assign n3472 = n3218 & ~n3403 ;
  assign n3473 = n3472 ^ n3215 ;
  assign n3474 = n3213 & ~n3403 ;
  assign n3475 = n3474 ^ n3212 ;
  assign n3476 = n3208 & n3403 ;
  assign n3477 = n3476 ^ n3205 ;
  assign n3478 = n3359 ^ n3356 ;
  assign n3479 = n3403 & n3478 ;
  assign n3480 = n3479 ^ n3359 ;
  assign n3481 = n3203 & ~n3403 ;
  assign n3482 = n3481 ^ n3200 ;
  assign n3483 = n3198 & ~n3403 ;
  assign n3484 = n3483 ^ n3195 ;
  assign n3485 = n3193 & n3403 ;
  assign n3486 = n3485 ^ n3190 ;
  assign n3487 = n3376 ^ n3373 ;
  assign n3488 = n3403 & n3487 ;
  assign n3489 = n3488 ^ n3376 ;
  assign n3490 = n3188 & ~n3403 ;
  assign n3491 = n3490 ^ n3187 ;
  assign n3492 = n3183 & ~n3403 ;
  assign n3493 = n3492 ^ n3180 ;
  assign n3494 = n3178 & n3403 ;
  assign n3495 = n3494 ^ n3175 ;
  assign n3496 = n3173 & ~n3403 ;
  assign n3497 = n3496 ^ n3170 ;
  assign n3498 = n3168 & n3403 ;
  assign n3499 = n3498 ^ n3165 ;
  assign n3500 = n3163 & ~n3403 ;
  assign n3501 = n3500 ^ n3162 ;
  assign n3502 = n3158 & n3403 ;
  assign n3503 = n3502 ^ n3157 ;
  assign n3504 = n519 & n526 ;
  assign y0 = ~n3436 ;
  assign y1 = ~n3415 ;
  assign y2 = n3406 ;
  assign y3 = ~n3403 ;
  assign y4 = n3439 ;
  assign y5 = n3441 ;
  assign y6 = n3443 ;
  assign y7 = n3445 ;
  assign y8 = n3447 ;
  assign y9 = n3449 ;
  assign y10 = n3451 ;
  assign y11 = n3453 ;
  assign y12 = n3455 ;
  assign y13 = n3457 ;
  assign y14 = n3459 ;
  assign y15 = n3462 ;
  assign y16 = n3464 ;
  assign y17 = n3466 ;
  assign y18 = n3468 ;
  assign y19 = n3471 ;
  assign y20 = n3473 ;
  assign y21 = n3475 ;
  assign y22 = n3477 ;
  assign y23 = n3480 ;
  assign y24 = n3482 ;
  assign y25 = n3484 ;
  assign y26 = n3486 ;
  assign y27 = n3489 ;
  assign y28 = n3491 ;
  assign y29 = n3493 ;
  assign y30 = n3495 ;
  assign y31 = n3497 ;
  assign y32 = n3499 ;
  assign y33 = n3501 ;
  assign y34 = n3503 ;
  assign y35 = ~n3504 ;
endmodule
