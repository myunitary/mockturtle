// eight voters and four candidate
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 ;
  assign n25 = ~x14 & x15 ;
  assign n57 = n25 ^ x15 ;
  assign n127 = n57 ^ x14 ;
  assign n24 = ~x12 & x13 ;
  assign n56 = n24 ^ x13 ;
  assign n126 = n56 ^ x12 ;
  assign n128 = n127 ^ n126 ;
  assign n27 = ~x10 & x11 ;
  assign n59 = n27 ^ x11 ;
  assign n125 = n59 ^ x10 ;
  assign n135 = n126 ^ n125 ;
  assign n136 = ~n128 & n135 ;
  assign n137 = n136 ^ n125 ;
  assign n129 = n128 ^ n125 ;
  assign n29 = ~x2 & x3 ;
  assign n61 = n29 ^ x3 ;
  assign n124 = n61 ^ x2 ;
  assign n130 = n129 ^ n124 ;
  assign n20 = ~x4 & x5 ;
  assign n54 = n20 ^ x5 ;
  assign n120 = n54 ^ x4 ;
  assign n18 = ~x8 & x9 ;
  assign n52 = n18 ^ x9 ;
  assign n118 = n52 ^ x8 ;
  assign n17 = ~x6 & x7 ;
  assign n51 = n17 ^ x7 ;
  assign n117 = n51 ^ x6 ;
  assign n119 = n118 ^ n117 ;
  assign n131 = n120 ^ n119 ;
  assign n132 = n131 ^ n129 ;
  assign n133 = n130 & ~n132 ;
  assign n134 = n133 ^ n124 ;
  assign n138 = n137 ^ n134 ;
  assign n121 = n120 ^ n117 ;
  assign n122 = ~n119 & n121 ;
  assign n123 = n122 ^ n120 ;
  assign n139 = n138 ^ n123 ;
  assign n140 = n131 ^ n130 ;
  assign n40 = ~x0 & x1 ;
  assign n50 = n40 ^ x1 ;
  assign n141 = n50 ^ x0 ;
  assign n142 = n140 & n141 ;
  assign n143 = n139 & n142 ;
  assign n144 = n137 ^ n123 ;
  assign n145 = n138 & ~n144 ;
  assign n146 = n145 ^ n134 ;
  assign n148 = ~n143 & ~n146 ;
  assign n147 = n146 ^ n143 ;
  assign n149 = n148 ^ n147 ;
  assign n94 = n27 ^ x10 ;
  assign n93 = n24 ^ x12 ;
  assign n95 = n94 ^ n93 ;
  assign n92 = n25 ^ x14 ;
  assign n102 = n93 ^ n92 ;
  assign n103 = ~n95 & n102 ;
  assign n104 = n103 ^ n92 ;
  assign n96 = n95 ^ n92 ;
  assign n91 = n29 ^ x2 ;
  assign n97 = n96 ^ n91 ;
  assign n87 = n18 ^ x8 ;
  assign n85 = n17 ^ x6 ;
  assign n84 = n20 ^ x4 ;
  assign n86 = n85 ^ n84 ;
  assign n98 = n87 ^ n86 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = n97 & ~n99 ;
  assign n101 = n100 ^ n91 ;
  assign n105 = n104 ^ n101 ;
  assign n88 = n87 ^ n84 ;
  assign n89 = ~n86 & n88 ;
  assign n90 = n89 ^ n87 ;
  assign n106 = n105 ^ n90 ;
  assign n107 = n98 ^ n97 ;
  assign n108 = n40 ^ x0 ;
  assign n109 = ~n107 & ~n108 ;
  assign n110 = ~n106 & n109 ;
  assign n111 = n104 ^ n90 ;
  assign n112 = n105 & ~n111 ;
  assign n113 = n112 ^ n101 ;
  assign n115 = ~n110 & n113 ;
  assign n114 = n113 ^ n110 ;
  assign n116 = n115 ^ n114 ;
  assign n150 = n149 ^ n116 ;
  assign n58 = n57 ^ n56 ;
  assign n60 = n59 ^ n58 ;
  assign n62 = n61 ^ n60 ;
  assign n53 = n52 ^ n51 ;
  assign n55 = n54 ^ n53 ;
  assign n63 = n62 ^ n55 ;
  assign n64 = n50 & n63 ;
  assign n71 = n61 ^ n55 ;
  assign n72 = n62 & ~n71 ;
  assign n73 = n72 ^ n60 ;
  assign n68 = n59 ^ n56 ;
  assign n69 = ~n58 & n68 ;
  assign n70 = n69 ^ n59 ;
  assign n74 = n73 ^ n70 ;
  assign n65 = n54 ^ n51 ;
  assign n66 = ~n53 & n65 ;
  assign n67 = n66 ^ n54 ;
  assign n75 = n74 ^ n67 ;
  assign n76 = n64 & n75 ;
  assign n77 = n73 ^ n67 ;
  assign n78 = n74 & ~n77 ;
  assign n79 = n78 ^ n70 ;
  assign n81 = ~n76 & ~n79 ;
  assign n80 = n79 ^ n76 ;
  assign n82 = n81 ^ n80 ;
  assign n26 = n25 ^ n24 ;
  assign n35 = n27 ^ n25 ;
  assign n36 = n26 & ~n35 ;
  assign n37 = n36 ^ n24 ;
  assign n28 = n27 ^ n26 ;
  assign n30 = n29 ^ n28 ;
  assign n19 = n18 ^ n17 ;
  assign n31 = n20 ^ n19 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n30 & ~n32 ;
  assign n34 = n33 ^ n28 ;
  assign n38 = n37 ^ n34 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n19 & ~n21 ;
  assign n23 = n22 ^ n17 ;
  assign n39 = n38 ^ n23 ;
  assign n41 = n31 ^ n30 ;
  assign n42 = n40 & n41 ;
  assign n43 = n39 & n42 ;
  assign n44 = n37 ^ n23 ;
  assign n45 = n38 & ~n44 ;
  assign n46 = n45 ^ n34 ;
  assign n48 = ~n43 & ~n46 ;
  assign n47 = n46 ^ n43 ;
  assign n49 = n48 ^ n47 ;
  assign n83 = n82 ^ n49 ;
  assign n151 = n150 ^ n83 ;
  assign n154 = n115 & n148 ;
  assign n155 = n154 ^ n150 ;
  assign n152 = n48 & n81 ;
  assign n153 = n152 ^ n83 ;
  assign n156 = n155 ^ n153 ;
  assign n157 = n80 ^ n47 ;
  assign n161 = n75 ^ n64 ;
  assign n158 = n63 ^ n50 ;
  assign n159 = n41 ^ n40 ;
  assign n160 = ~n158 & n159 ;
  assign n162 = n161 ^ n160 ;
  assign n163 = n160 ^ n42 ;
  assign n164 = n163 ^ n39 ;
  assign n165 = ~n162 & ~n164 ;
  assign n166 = n165 ^ n161 ;
  assign n167 = n166 ^ n47 ;
  assign n168 = ~n157 & n167 ;
  assign n169 = n168 ^ n80 ;
  assign n170 = n169 ^ n82 ;
  assign n171 = ~n83 & n170 ;
  assign n172 = n171 ^ n49 ;
  assign n196 = n42 ^ n39 ;
  assign n197 = n196 ^ n161 ;
  assign n198 = ~n172 & n197 ;
  assign n199 = n198 ^ n161 ;
  assign n173 = n159 ^ n158 ;
  assign n174 = ~n172 & n173 ;
  assign n175 = n174 ^ n158 ;
  assign n177 = n141 ^ n140 ;
  assign n176 = n108 ^ n107 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = n147 ^ n114 ;
  assign n181 = n142 ^ n139 ;
  assign n180 = n109 ^ n106 ;
  assign n182 = n181 ^ n180 ;
  assign n183 = n176 & ~n177 ;
  assign n184 = n183 ^ n180 ;
  assign n185 = ~n182 & ~n184 ;
  assign n186 = n185 ^ n183 ;
  assign n187 = n186 ^ n114 ;
  assign n188 = n179 & ~n187 ;
  assign n189 = n188 ^ n114 ;
  assign n190 = n189 ^ n149 ;
  assign n191 = n150 & n190 ;
  assign n192 = n191 ^ n116 ;
  assign n193 = n178 & ~n192 ;
  assign n194 = n193 ^ n176 ;
  assign n195 = ~n175 & n194 ;
  assign n200 = n199 ^ n195 ;
  assign n201 = ~n182 & ~n192 ;
  assign n202 = n201 ^ n180 ;
  assign n203 = n202 ^ n199 ;
  assign n204 = ~n200 & ~n203 ;
  assign n205 = n204 ^ n195 ;
  assign n206 = n205 ^ n153 ;
  assign n207 = n156 & ~n206 ;
  assign n208 = n207 ^ n155 ;
  assign n209 = n208 ^ n83 ;
  assign n210 = n151 & n209 ;
  assign n211 = n210 ^ n150 ;
  assign n212 = n192 ^ n172 ;
  assign n213 = ~n211 & ~n212 ;
  assign n214 = n213 ^ n172 ;
  assign y0 = n214 ;
  assign y1 = n211 ;
endmodule
