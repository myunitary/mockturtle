module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 ;
  assign n730 = x0 & ~x8 ;
  assign n695 = x8 ^ x0 ;
  assign n728 = x1 & ~x9 ;
  assign n729 = ~n695 & n728 ;
  assign n731 = n730 ^ n729 ;
  assign n696 = x9 ^ x1 ;
  assign n697 = ~n695 & ~n696 ;
  assign n725 = x2 & ~x10 ;
  assign n698 = x10 ^ x2 ;
  assign n723 = x3 & ~x11 ;
  assign n724 = ~n698 & n723 ;
  assign n726 = n725 ^ n724 ;
  assign n727 = n697 & n726 ;
  assign n732 = n731 ^ n727 ;
  assign n699 = x11 ^ x3 ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = n697 & n700 ;
  assign n719 = x4 & ~x12 ;
  assign n702 = x12 ^ x4 ;
  assign n717 = x5 & ~x13 ;
  assign n718 = ~n702 & n717 ;
  assign n720 = n719 ^ n718 ;
  assign n703 = x13 ^ x5 ;
  assign n704 = ~n702 & ~n703 ;
  assign n714 = x6 & ~x14 ;
  assign n705 = x14 ^ x6 ;
  assign n710 = x7 & x15 ;
  assign n711 = n710 ^ x7 ;
  assign n712 = n705 & n711 ;
  assign n713 = n712 ^ n711 ;
  assign n715 = n714 ^ n713 ;
  assign n716 = n704 & n715 ;
  assign n721 = n720 ^ n716 ;
  assign n722 = n701 & n721 ;
  assign n733 = n732 ^ n722 ;
  assign n706 = x15 ^ x7 ;
  assign n707 = ~n705 & ~n706 ;
  assign n708 = n704 & n707 ;
  assign n709 = n701 & n708 ;
  assign n734 = n733 ^ n709 ;
  assign n631 = x0 & ~x16 ;
  assign n596 = x16 ^ x0 ;
  assign n629 = x1 & ~x17 ;
  assign n630 = ~n596 & n629 ;
  assign n632 = n631 ^ n630 ;
  assign n597 = x17 ^ x1 ;
  assign n598 = ~n596 & ~n597 ;
  assign n626 = x2 & ~x18 ;
  assign n599 = x18 ^ x2 ;
  assign n624 = x3 & ~x19 ;
  assign n625 = ~n599 & n624 ;
  assign n627 = n626 ^ n625 ;
  assign n628 = n598 & n627 ;
  assign n633 = n632 ^ n628 ;
  assign n600 = x19 ^ x3 ;
  assign n601 = ~n599 & ~n600 ;
  assign n602 = n598 & n601 ;
  assign n620 = x4 & ~x20 ;
  assign n603 = x20 ^ x4 ;
  assign n618 = x5 & ~x21 ;
  assign n619 = ~n603 & n618 ;
  assign n621 = n620 ^ n619 ;
  assign n604 = x21 ^ x5 ;
  assign n605 = ~n603 & ~n604 ;
  assign n615 = x6 & ~x22 ;
  assign n606 = x22 ^ x6 ;
  assign n611 = x7 & x23 ;
  assign n612 = n611 ^ x7 ;
  assign n613 = n606 & n612 ;
  assign n614 = n613 ^ n612 ;
  assign n616 = n615 ^ n614 ;
  assign n617 = n605 & n616 ;
  assign n622 = n621 ^ n617 ;
  assign n623 = n602 & n622 ;
  assign n634 = n633 ^ n623 ;
  assign n607 = x23 ^ x7 ;
  assign n608 = ~n606 & ~n607 ;
  assign n609 = n605 & n608 ;
  assign n610 = n602 & n609 ;
  assign n635 = n634 ^ n610 ;
  assign n755 = n734 ^ n635 ;
  assign n388 = x0 & ~x32 ;
  assign n353 = x32 ^ x0 ;
  assign n386 = x1 & ~x33 ;
  assign n387 = ~n353 & n386 ;
  assign n389 = n388 ^ n387 ;
  assign n354 = x33 ^ x1 ;
  assign n355 = ~n353 & ~n354 ;
  assign n383 = x2 & ~x34 ;
  assign n356 = x34 ^ x2 ;
  assign n381 = x3 & ~x35 ;
  assign n382 = ~n356 & n381 ;
  assign n384 = n383 ^ n382 ;
  assign n385 = n355 & n384 ;
  assign n390 = n389 ^ n385 ;
  assign n357 = x35 ^ x3 ;
  assign n358 = ~n356 & ~n357 ;
  assign n359 = n355 & n358 ;
  assign n377 = x4 & ~x36 ;
  assign n360 = x36 ^ x4 ;
  assign n375 = x5 & ~x37 ;
  assign n376 = ~n360 & n375 ;
  assign n378 = n377 ^ n376 ;
  assign n361 = x37 ^ x5 ;
  assign n362 = ~n360 & ~n361 ;
  assign n372 = x6 & ~x38 ;
  assign n363 = x38 ^ x6 ;
  assign n368 = x7 & x39 ;
  assign n369 = n368 ^ x7 ;
  assign n370 = n363 & n369 ;
  assign n371 = n370 ^ n369 ;
  assign n373 = n372 ^ n371 ;
  assign n374 = n362 & n373 ;
  assign n379 = n378 ^ n374 ;
  assign n380 = n359 & n379 ;
  assign n391 = n390 ^ n380 ;
  assign n364 = x39 ^ x7 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = n362 & n365 ;
  assign n367 = n359 & n366 ;
  assign n392 = n391 ^ n367 ;
  assign n165 = x0 & ~x40 ;
  assign n130 = x40 ^ x0 ;
  assign n163 = x1 & ~x41 ;
  assign n164 = ~n130 & n163 ;
  assign n166 = n165 ^ n164 ;
  assign n131 = x41 ^ x1 ;
  assign n132 = ~n130 & ~n131 ;
  assign n160 = x2 & ~x42 ;
  assign n133 = x42 ^ x2 ;
  assign n158 = x3 & ~x43 ;
  assign n159 = ~n133 & n158 ;
  assign n161 = n160 ^ n159 ;
  assign n162 = n132 & n161 ;
  assign n167 = n166 ^ n162 ;
  assign n134 = x43 ^ x3 ;
  assign n135 = ~n133 & ~n134 ;
  assign n136 = n132 & n135 ;
  assign n154 = x4 & ~x44 ;
  assign n137 = x44 ^ x4 ;
  assign n152 = x5 & ~x45 ;
  assign n153 = ~n137 & n152 ;
  assign n155 = n154 ^ n153 ;
  assign n138 = x45 ^ x5 ;
  assign n139 = ~n137 & ~n138 ;
  assign n149 = x6 & ~x46 ;
  assign n140 = x46 ^ x6 ;
  assign n145 = x7 & x47 ;
  assign n146 = n145 ^ x7 ;
  assign n147 = n140 & n146 ;
  assign n148 = n147 ^ n146 ;
  assign n150 = n149 ^ n148 ;
  assign n151 = n139 & n150 ;
  assign n156 = n155 ^ n151 ;
  assign n157 = n136 & n156 ;
  assign n168 = n167 ^ n157 ;
  assign n141 = x47 ^ x7 ;
  assign n142 = ~n140 & ~n141 ;
  assign n143 = n139 & n142 ;
  assign n144 = n136 & n143 ;
  assign n169 = n168 ^ n144 ;
  assign n756 = n392 ^ n169 ;
  assign n572 = x0 & ~x24 ;
  assign n537 = x24 ^ x0 ;
  assign n570 = x1 & ~x25 ;
  assign n571 = ~n537 & n570 ;
  assign n573 = n572 ^ n571 ;
  assign n538 = x25 ^ x1 ;
  assign n539 = ~n537 & ~n538 ;
  assign n567 = x2 & ~x26 ;
  assign n540 = x26 ^ x2 ;
  assign n565 = x3 & ~x27 ;
  assign n566 = ~n540 & n565 ;
  assign n568 = n567 ^ n566 ;
  assign n569 = n539 & n568 ;
  assign n574 = n573 ^ n569 ;
  assign n541 = x27 ^ x3 ;
  assign n542 = ~n540 & ~n541 ;
  assign n543 = n539 & n542 ;
  assign n561 = x4 & ~x28 ;
  assign n544 = x28 ^ x4 ;
  assign n559 = x5 & ~x29 ;
  assign n560 = ~n544 & n559 ;
  assign n562 = n561 ^ n560 ;
  assign n545 = x29 ^ x5 ;
  assign n546 = ~n544 & ~n545 ;
  assign n556 = x6 & ~x30 ;
  assign n547 = x30 ^ x6 ;
  assign n552 = x7 & x31 ;
  assign n553 = n552 ^ x7 ;
  assign n554 = n547 & n553 ;
  assign n555 = n554 ^ n553 ;
  assign n557 = n556 ^ n555 ;
  assign n558 = n546 & n557 ;
  assign n563 = n562 ^ n558 ;
  assign n564 = n543 & n563 ;
  assign n575 = n574 ^ n564 ;
  assign n548 = x31 ^ x7 ;
  assign n549 = ~n547 & ~n548 ;
  assign n550 = n546 & n549 ;
  assign n551 = n543 & n550 ;
  assign n576 = n575 ^ n551 ;
  assign n757 = n756 ^ n576 ;
  assign n758 = n755 & n757 ;
  assign n754 = n635 & n734 ;
  assign n759 = n758 ^ n754 ;
  assign n761 = n576 & n756 ;
  assign n760 = n169 & n392 ;
  assign n762 = n761 ^ n760 ;
  assign n763 = n762 ^ n758 ;
  assign n764 = n759 & n763 ;
  assign n765 = n764 ^ n758 ;
  assign n766 = n757 ^ n755 ;
  assign n767 = n762 ^ n759 ;
  assign n768 = ~n766 & ~n767 ;
  assign n769 = ~n765 & n768 ;
  assign n770 = x0 & n769 ;
  assign n671 = x8 & ~x16 ;
  assign n636 = x16 ^ x8 ;
  assign n669 = x9 & ~x17 ;
  assign n670 = ~n636 & n669 ;
  assign n672 = n671 ^ n670 ;
  assign n637 = x17 ^ x9 ;
  assign n638 = ~n636 & ~n637 ;
  assign n666 = x10 & ~x18 ;
  assign n639 = x18 ^ x10 ;
  assign n664 = x11 & ~x19 ;
  assign n665 = ~n639 & n664 ;
  assign n667 = n666 ^ n665 ;
  assign n668 = n638 & n667 ;
  assign n673 = n672 ^ n668 ;
  assign n640 = x19 ^ x11 ;
  assign n641 = ~n639 & ~n640 ;
  assign n642 = n638 & n641 ;
  assign n660 = x12 & ~x20 ;
  assign n643 = x20 ^ x12 ;
  assign n658 = x13 & ~x21 ;
  assign n659 = ~n643 & n658 ;
  assign n661 = n660 ^ n659 ;
  assign n644 = x21 ^ x13 ;
  assign n645 = ~n643 & ~n644 ;
  assign n655 = x14 & ~x22 ;
  assign n646 = x22 ^ x14 ;
  assign n651 = x15 & x23 ;
  assign n652 = n651 ^ x15 ;
  assign n653 = n646 & n652 ;
  assign n654 = n653 ^ n652 ;
  assign n656 = n655 ^ n654 ;
  assign n657 = n645 & n656 ;
  assign n662 = n661 ^ n657 ;
  assign n663 = n642 & n662 ;
  assign n674 = n673 ^ n663 ;
  assign n647 = x23 ^ x15 ;
  assign n648 = ~n646 & ~n647 ;
  assign n649 = n645 & n648 ;
  assign n650 = n642 & n649 ;
  assign n675 = n674 ^ n650 ;
  assign n737 = n734 ^ n675 ;
  assign n347 = x8 & ~x32 ;
  assign n312 = x32 ^ x8 ;
  assign n345 = x9 & ~x33 ;
  assign n346 = ~n312 & n345 ;
  assign n348 = n347 ^ n346 ;
  assign n313 = x33 ^ x9 ;
  assign n314 = ~n312 & ~n313 ;
  assign n342 = x10 & ~x34 ;
  assign n315 = x34 ^ x10 ;
  assign n340 = x11 & ~x35 ;
  assign n341 = ~n315 & n340 ;
  assign n343 = n342 ^ n341 ;
  assign n344 = n314 & n343 ;
  assign n349 = n348 ^ n344 ;
  assign n316 = x35 ^ x11 ;
  assign n317 = ~n315 & ~n316 ;
  assign n318 = n314 & n317 ;
  assign n336 = x12 & ~x36 ;
  assign n319 = x36 ^ x12 ;
  assign n334 = x13 & ~x37 ;
  assign n335 = ~n319 & n334 ;
  assign n337 = n336 ^ n335 ;
  assign n320 = x37 ^ x13 ;
  assign n321 = ~n319 & ~n320 ;
  assign n331 = x14 & ~x38 ;
  assign n322 = x38 ^ x14 ;
  assign n327 = x15 & x39 ;
  assign n328 = n327 ^ x15 ;
  assign n329 = n322 & n328 ;
  assign n330 = n329 ^ n328 ;
  assign n332 = n331 ^ n330 ;
  assign n333 = n321 & n332 ;
  assign n338 = n337 ^ n333 ;
  assign n339 = n318 & n338 ;
  assign n350 = n349 ^ n339 ;
  assign n323 = x39 ^ x15 ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = n321 & n324 ;
  assign n326 = n318 & n325 ;
  assign n351 = n350 ^ n326 ;
  assign n124 = x8 & ~x40 ;
  assign n89 = x40 ^ x8 ;
  assign n122 = x9 & ~x41 ;
  assign n123 = ~n89 & n122 ;
  assign n125 = n124 ^ n123 ;
  assign n90 = x41 ^ x9 ;
  assign n91 = ~n89 & ~n90 ;
  assign n119 = x10 & ~x42 ;
  assign n92 = x42 ^ x10 ;
  assign n117 = x11 & ~x43 ;
  assign n118 = ~n92 & n117 ;
  assign n120 = n119 ^ n118 ;
  assign n121 = n91 & n120 ;
  assign n126 = n125 ^ n121 ;
  assign n93 = x43 ^ x11 ;
  assign n94 = ~n92 & ~n93 ;
  assign n95 = n91 & n94 ;
  assign n113 = x12 & ~x44 ;
  assign n96 = x44 ^ x12 ;
  assign n111 = x13 & ~x45 ;
  assign n112 = ~n96 & n111 ;
  assign n114 = n113 ^ n112 ;
  assign n97 = x45 ^ x13 ;
  assign n98 = ~n96 & ~n97 ;
  assign n108 = x14 & ~x46 ;
  assign n99 = x46 ^ x14 ;
  assign n104 = x15 & x47 ;
  assign n105 = n104 ^ x15 ;
  assign n106 = n99 & n105 ;
  assign n107 = n106 ^ n105 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = n98 & n109 ;
  assign n115 = n114 ^ n110 ;
  assign n116 = n95 & n115 ;
  assign n127 = n126 ^ n116 ;
  assign n100 = x47 ^ x15 ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = n98 & n101 ;
  assign n103 = n95 & n102 ;
  assign n128 = n127 ^ n103 ;
  assign n738 = n351 ^ n128 ;
  assign n531 = x8 & ~x24 ;
  assign n496 = x24 ^ x8 ;
  assign n529 = x9 & ~x25 ;
  assign n530 = ~n496 & n529 ;
  assign n532 = n531 ^ n530 ;
  assign n497 = x25 ^ x9 ;
  assign n498 = ~n496 & ~n497 ;
  assign n526 = x10 & ~x26 ;
  assign n499 = x26 ^ x10 ;
  assign n524 = x11 & ~x27 ;
  assign n525 = ~n499 & n524 ;
  assign n527 = n526 ^ n525 ;
  assign n528 = n498 & n527 ;
  assign n533 = n532 ^ n528 ;
  assign n500 = x27 ^ x11 ;
  assign n501 = ~n499 & ~n500 ;
  assign n502 = n498 & n501 ;
  assign n520 = x12 & ~x28 ;
  assign n503 = x28 ^ x12 ;
  assign n518 = x13 & ~x29 ;
  assign n519 = ~n503 & n518 ;
  assign n521 = n520 ^ n519 ;
  assign n504 = x29 ^ x13 ;
  assign n505 = ~n503 & ~n504 ;
  assign n515 = x14 & ~x30 ;
  assign n506 = x30 ^ x14 ;
  assign n511 = x15 & x31 ;
  assign n512 = n511 ^ x15 ;
  assign n513 = n506 & n512 ;
  assign n514 = n513 ^ n512 ;
  assign n516 = n515 ^ n514 ;
  assign n517 = n505 & n516 ;
  assign n522 = n521 ^ n517 ;
  assign n523 = n502 & n522 ;
  assign n534 = n533 ^ n523 ;
  assign n507 = x31 ^ x15 ;
  assign n508 = ~n506 & ~n507 ;
  assign n509 = n505 & n508 ;
  assign n510 = n502 & n509 ;
  assign n535 = n534 ^ n510 ;
  assign n739 = n738 ^ n535 ;
  assign n740 = n737 & n739 ;
  assign n741 = n740 ^ n739 ;
  assign n735 = n675 & n734 ;
  assign n736 = n735 ^ n675 ;
  assign n742 = n741 ^ n736 ;
  assign n744 = n535 & n738 ;
  assign n743 = n128 & n351 ;
  assign n745 = n744 ^ n743 ;
  assign n746 = n745 ^ n741 ;
  assign n747 = n742 & n746 ;
  assign n748 = n747 ^ n741 ;
  assign n749 = n739 ^ n737 ;
  assign n750 = n745 ^ n742 ;
  assign n751 = n749 & ~n750 ;
  assign n752 = ~n748 & n751 ;
  assign n753 = x8 & n752 ;
  assign n771 = n770 ^ n753 ;
  assign n679 = n675 ^ n635 ;
  assign n307 = x16 & ~x32 ;
  assign n272 = x32 ^ x16 ;
  assign n305 = x17 & ~x33 ;
  assign n306 = ~n272 & n305 ;
  assign n308 = n307 ^ n306 ;
  assign n273 = x33 ^ x17 ;
  assign n274 = ~n272 & ~n273 ;
  assign n302 = x18 & ~x34 ;
  assign n275 = x34 ^ x18 ;
  assign n300 = x19 & ~x35 ;
  assign n301 = ~n275 & n300 ;
  assign n303 = n302 ^ n301 ;
  assign n304 = n274 & n303 ;
  assign n309 = n308 ^ n304 ;
  assign n276 = x35 ^ x19 ;
  assign n277 = ~n275 & ~n276 ;
  assign n278 = n274 & n277 ;
  assign n296 = x20 & ~x36 ;
  assign n279 = x36 ^ x20 ;
  assign n294 = x21 & ~x37 ;
  assign n295 = ~n279 & n294 ;
  assign n297 = n296 ^ n295 ;
  assign n280 = x37 ^ x21 ;
  assign n281 = ~n279 & ~n280 ;
  assign n291 = x22 & ~x38 ;
  assign n282 = x38 ^ x22 ;
  assign n287 = x23 & x39 ;
  assign n288 = n287 ^ x23 ;
  assign n289 = n282 & n288 ;
  assign n290 = n289 ^ n288 ;
  assign n292 = n291 ^ n290 ;
  assign n293 = n281 & n292 ;
  assign n298 = n297 ^ n293 ;
  assign n299 = n278 & n298 ;
  assign n310 = n309 ^ n299 ;
  assign n283 = x39 ^ x23 ;
  assign n284 = ~n282 & ~n283 ;
  assign n285 = n281 & n284 ;
  assign n286 = n278 & n285 ;
  assign n311 = n310 ^ n286 ;
  assign n84 = x16 & ~x40 ;
  assign n49 = x40 ^ x16 ;
  assign n82 = x17 & ~x41 ;
  assign n83 = ~n49 & n82 ;
  assign n85 = n84 ^ n83 ;
  assign n50 = x41 ^ x17 ;
  assign n51 = ~n49 & ~n50 ;
  assign n79 = x18 & ~x42 ;
  assign n52 = x42 ^ x18 ;
  assign n77 = x19 & ~x43 ;
  assign n78 = ~n52 & n77 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n51 & n80 ;
  assign n86 = n85 ^ n81 ;
  assign n53 = x43 ^ x19 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n51 & n54 ;
  assign n73 = x20 & ~x44 ;
  assign n56 = x44 ^ x20 ;
  assign n71 = x21 & ~x45 ;
  assign n72 = ~n56 & n71 ;
  assign n74 = n73 ^ n72 ;
  assign n57 = x45 ^ x21 ;
  assign n58 = ~n56 & ~n57 ;
  assign n68 = x22 & ~x46 ;
  assign n59 = x46 ^ x22 ;
  assign n64 = x23 & x47 ;
  assign n65 = n64 ^ x23 ;
  assign n66 = n59 & n65 ;
  assign n67 = n66 ^ n65 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n58 & n69 ;
  assign n75 = n74 ^ n70 ;
  assign n76 = n55 & n75 ;
  assign n87 = n86 ^ n76 ;
  assign n60 = x47 ^ x23 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = n58 & n61 ;
  assign n63 = n55 & n62 ;
  assign n88 = n87 ^ n63 ;
  assign n680 = n311 ^ n88 ;
  assign n491 = x16 & ~x24 ;
  assign n456 = x24 ^ x16 ;
  assign n489 = x17 & ~x25 ;
  assign n490 = ~n456 & n489 ;
  assign n492 = n491 ^ n490 ;
  assign n457 = x25 ^ x17 ;
  assign n458 = ~n456 & ~n457 ;
  assign n486 = x18 & ~x26 ;
  assign n459 = x26 ^ x18 ;
  assign n484 = x19 & ~x27 ;
  assign n485 = ~n459 & n484 ;
  assign n487 = n486 ^ n485 ;
  assign n488 = n458 & n487 ;
  assign n493 = n492 ^ n488 ;
  assign n460 = x27 ^ x19 ;
  assign n461 = ~n459 & ~n460 ;
  assign n462 = n458 & n461 ;
  assign n480 = x20 & ~x28 ;
  assign n463 = x28 ^ x20 ;
  assign n478 = x21 & ~x29 ;
  assign n479 = ~n463 & n478 ;
  assign n481 = n480 ^ n479 ;
  assign n464 = x29 ^ x21 ;
  assign n465 = ~n463 & ~n464 ;
  assign n475 = x22 & ~x30 ;
  assign n466 = x30 ^ x22 ;
  assign n471 = x23 & x31 ;
  assign n472 = n471 ^ x23 ;
  assign n473 = n466 & n472 ;
  assign n474 = n473 ^ n472 ;
  assign n476 = n475 ^ n474 ;
  assign n477 = n465 & n476 ;
  assign n482 = n481 ^ n477 ;
  assign n483 = n462 & n482 ;
  assign n494 = n493 ^ n483 ;
  assign n467 = x31 ^ x23 ;
  assign n468 = ~n466 & ~n467 ;
  assign n469 = n465 & n468 ;
  assign n470 = n462 & n469 ;
  assign n495 = n494 ^ n470 ;
  assign n681 = n680 ^ n495 ;
  assign n682 = n679 & n681 ;
  assign n676 = n635 & n675 ;
  assign n677 = n676 ^ n675 ;
  assign n678 = n677 ^ n635 ;
  assign n683 = n682 ^ n678 ;
  assign n685 = n495 & n680 ;
  assign n684 = n88 & n311 ;
  assign n686 = n685 ^ n684 ;
  assign n687 = n686 ^ n682 ;
  assign n688 = ~n683 & n687 ;
  assign n689 = n688 ^ n682 ;
  assign n690 = n681 ^ n679 ;
  assign n691 = n686 ^ n683 ;
  assign n692 = ~n690 & n691 ;
  assign n693 = ~n689 & n692 ;
  assign n694 = x16 & n693 ;
  assign n772 = n771 ^ n694 ;
  assign n536 = n535 ^ n495 ;
  assign n583 = n536 & n576 ;
  assign n584 = n583 ^ n536 ;
  assign n580 = n495 & n535 ;
  assign n581 = n580 ^ n495 ;
  assign n582 = n581 ^ n535 ;
  assign n585 = n584 ^ n582 ;
  assign n429 = x24 & ~x32 ;
  assign n394 = x32 ^ x24 ;
  assign n427 = x25 & ~x33 ;
  assign n428 = ~n394 & n427 ;
  assign n430 = n429 ^ n428 ;
  assign n395 = x33 ^ x25 ;
  assign n396 = ~n394 & ~n395 ;
  assign n424 = x26 & ~x34 ;
  assign n397 = x34 ^ x26 ;
  assign n422 = x27 & ~x35 ;
  assign n423 = ~n397 & n422 ;
  assign n425 = n424 ^ n423 ;
  assign n426 = n396 & n425 ;
  assign n431 = n430 ^ n426 ;
  assign n398 = x35 ^ x27 ;
  assign n399 = ~n397 & ~n398 ;
  assign n400 = n396 & n399 ;
  assign n418 = x28 & ~x36 ;
  assign n401 = x36 ^ x28 ;
  assign n416 = x29 & ~x37 ;
  assign n417 = ~n401 & n416 ;
  assign n419 = n418 ^ n417 ;
  assign n402 = x37 ^ x29 ;
  assign n403 = ~n401 & ~n402 ;
  assign n413 = x30 & ~x38 ;
  assign n404 = x38 ^ x30 ;
  assign n409 = x31 & x39 ;
  assign n410 = n409 ^ x31 ;
  assign n411 = n404 & n410 ;
  assign n412 = n411 ^ n410 ;
  assign n414 = n413 ^ n412 ;
  assign n415 = n403 & n414 ;
  assign n420 = n419 ^ n415 ;
  assign n421 = n400 & n420 ;
  assign n432 = n431 ^ n421 ;
  assign n405 = x39 ^ x31 ;
  assign n406 = ~n404 & ~n405 ;
  assign n407 = n403 & n406 ;
  assign n408 = n400 & n407 ;
  assign n433 = n432 ^ n408 ;
  assign n246 = x24 & ~x40 ;
  assign n211 = x40 ^ x24 ;
  assign n244 = x25 & ~x41 ;
  assign n245 = ~n211 & n244 ;
  assign n247 = n246 ^ n245 ;
  assign n212 = x41 ^ x25 ;
  assign n213 = ~n211 & ~n212 ;
  assign n241 = x26 & ~x42 ;
  assign n214 = x42 ^ x26 ;
  assign n239 = x27 & ~x43 ;
  assign n240 = ~n214 & n239 ;
  assign n242 = n241 ^ n240 ;
  assign n243 = n213 & n242 ;
  assign n248 = n247 ^ n243 ;
  assign n215 = x43 ^ x27 ;
  assign n216 = ~n214 & ~n215 ;
  assign n217 = n213 & n216 ;
  assign n235 = x28 & ~x44 ;
  assign n218 = x44 ^ x28 ;
  assign n233 = x29 & ~x45 ;
  assign n234 = ~n218 & n233 ;
  assign n236 = n235 ^ n234 ;
  assign n219 = x45 ^ x29 ;
  assign n220 = ~n218 & ~n219 ;
  assign n230 = x30 & ~x46 ;
  assign n221 = x46 ^ x30 ;
  assign n226 = x31 & x47 ;
  assign n227 = n226 ^ x31 ;
  assign n228 = n221 & n227 ;
  assign n229 = n228 ^ n227 ;
  assign n231 = n230 ^ n229 ;
  assign n232 = n220 & n231 ;
  assign n237 = n236 ^ n232 ;
  assign n238 = n217 & n237 ;
  assign n249 = n248 ^ n238 ;
  assign n222 = x47 ^ x31 ;
  assign n223 = ~n221 & ~n222 ;
  assign n224 = n220 & n223 ;
  assign n225 = n217 & n224 ;
  assign n250 = n249 ^ n225 ;
  assign n455 = n433 ^ n250 ;
  assign n577 = n576 ^ n536 ;
  assign n578 = n455 & n577 ;
  assign n579 = n578 ^ n455 ;
  assign n586 = n585 ^ n579 ;
  assign n587 = n250 & n433 ;
  assign n588 = n587 ^ n579 ;
  assign n589 = ~n586 & n588 ;
  assign n590 = n589 ^ n579 ;
  assign n591 = n577 ^ n455 ;
  assign n592 = n587 ^ n586 ;
  assign n593 = n591 & n592 ;
  assign n594 = ~n590 & n593 ;
  assign n595 = x24 & n594 ;
  assign n773 = n772 ^ n595 ;
  assign n352 = n351 ^ n311 ;
  assign n441 = n352 & n392 ;
  assign n442 = n441 ^ n352 ;
  assign n438 = n311 & n351 ;
  assign n439 = n438 ^ n311 ;
  assign n440 = n439 ^ n351 ;
  assign n443 = n442 ^ n440 ;
  assign n393 = n392 ^ n352 ;
  assign n206 = x32 & ~x40 ;
  assign n171 = x40 ^ x32 ;
  assign n204 = x33 & ~x41 ;
  assign n205 = ~n171 & n204 ;
  assign n207 = n206 ^ n205 ;
  assign n172 = x41 ^ x33 ;
  assign n173 = ~n171 & ~n172 ;
  assign n201 = x34 & ~x42 ;
  assign n174 = x42 ^ x34 ;
  assign n199 = x35 & ~x43 ;
  assign n200 = ~n174 & n199 ;
  assign n202 = n201 ^ n200 ;
  assign n203 = n173 & n202 ;
  assign n208 = n207 ^ n203 ;
  assign n175 = x43 ^ x35 ;
  assign n176 = ~n174 & ~n175 ;
  assign n177 = n173 & n176 ;
  assign n195 = x36 & ~x44 ;
  assign n178 = x44 ^ x36 ;
  assign n193 = x37 & ~x45 ;
  assign n194 = ~n178 & n193 ;
  assign n196 = n195 ^ n194 ;
  assign n179 = x45 ^ x37 ;
  assign n180 = ~n178 & ~n179 ;
  assign n190 = x38 & ~x46 ;
  assign n181 = x46 ^ x38 ;
  assign n186 = x39 & x47 ;
  assign n187 = n186 ^ x39 ;
  assign n188 = n181 & n187 ;
  assign n189 = n188 ^ n187 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = n180 & n191 ;
  assign n197 = n196 ^ n192 ;
  assign n198 = n177 & n197 ;
  assign n209 = n208 ^ n198 ;
  assign n182 = x47 ^ x39 ;
  assign n183 = ~n181 & ~n182 ;
  assign n184 = n180 & n183 ;
  assign n185 = n177 & n184 ;
  assign n210 = n209 ^ n185 ;
  assign n434 = n433 ^ n210 ;
  assign n435 = n393 & n434 ;
  assign n436 = n435 ^ n434 ;
  assign n437 = n436 ^ n393 ;
  assign n444 = n443 ^ n437 ;
  assign n445 = n210 & n433 ;
  assign n446 = n445 ^ n210 ;
  assign n447 = n446 ^ n437 ;
  assign n448 = n444 & ~n447 ;
  assign n449 = n448 ^ n437 ;
  assign n450 = n434 ^ n393 ;
  assign n451 = n446 ^ n444 ;
  assign n452 = ~n450 & ~n451 ;
  assign n453 = n449 & n452 ;
  assign n454 = x32 & n453 ;
  assign n774 = n773 ^ n454 ;
  assign n129 = n128 ^ n88 ;
  assign n257 = n129 & n169 ;
  assign n258 = n257 ^ n129 ;
  assign n254 = n88 & n128 ;
  assign n255 = n254 ^ n88 ;
  assign n256 = n255 ^ n128 ;
  assign n259 = n258 ^ n256 ;
  assign n170 = n169 ^ n129 ;
  assign n251 = n250 ^ n210 ;
  assign n252 = n170 & n251 ;
  assign n253 = n252 ^ n251 ;
  assign n260 = n259 ^ n253 ;
  assign n261 = n210 & n250 ;
  assign n262 = n261 ^ n210 ;
  assign n263 = n262 ^ n250 ;
  assign n264 = n263 ^ n253 ;
  assign n265 = ~n260 & ~n264 ;
  assign n266 = n265 ^ n253 ;
  assign n267 = n251 ^ n170 ;
  assign n268 = n263 ^ n260 ;
  assign n269 = n267 & ~n268 ;
  assign n270 = ~n266 & n269 ;
  assign n271 = x40 & n270 ;
  assign n775 = n774 ^ n271 ;
  assign n781 = x1 & n769 ;
  assign n780 = x9 & n752 ;
  assign n782 = n781 ^ n780 ;
  assign n779 = x17 & n693 ;
  assign n783 = n782 ^ n779 ;
  assign n778 = x25 & n594 ;
  assign n784 = n783 ^ n778 ;
  assign n777 = x33 & n453 ;
  assign n785 = n784 ^ n777 ;
  assign n776 = x41 & n270 ;
  assign n786 = n785 ^ n776 ;
  assign n792 = x2 & n769 ;
  assign n791 = x10 & n752 ;
  assign n793 = n792 ^ n791 ;
  assign n790 = x18 & n693 ;
  assign n794 = n793 ^ n790 ;
  assign n789 = x26 & n594 ;
  assign n795 = n794 ^ n789 ;
  assign n788 = x34 & n453 ;
  assign n796 = n795 ^ n788 ;
  assign n787 = x42 & n270 ;
  assign n797 = n796 ^ n787 ;
  assign n803 = x3 & n769 ;
  assign n802 = x11 & n752 ;
  assign n804 = n803 ^ n802 ;
  assign n801 = x19 & n693 ;
  assign n805 = n804 ^ n801 ;
  assign n800 = x27 & n594 ;
  assign n806 = n805 ^ n800 ;
  assign n799 = x35 & n453 ;
  assign n807 = n806 ^ n799 ;
  assign n798 = x43 & n270 ;
  assign n808 = n807 ^ n798 ;
  assign n814 = x4 & n769 ;
  assign n813 = x12 & n752 ;
  assign n815 = n814 ^ n813 ;
  assign n812 = x20 & n693 ;
  assign n816 = n815 ^ n812 ;
  assign n811 = x28 & n594 ;
  assign n817 = n816 ^ n811 ;
  assign n810 = x36 & n453 ;
  assign n818 = n817 ^ n810 ;
  assign n809 = x44 & n270 ;
  assign n819 = n818 ^ n809 ;
  assign n825 = x5 & n769 ;
  assign n824 = x13 & n752 ;
  assign n826 = n825 ^ n824 ;
  assign n823 = x21 & n693 ;
  assign n827 = n826 ^ n823 ;
  assign n822 = x29 & n594 ;
  assign n828 = n827 ^ n822 ;
  assign n821 = x37 & n453 ;
  assign n829 = n828 ^ n821 ;
  assign n820 = x45 & n270 ;
  assign n830 = n829 ^ n820 ;
  assign n836 = x6 & n769 ;
  assign n835 = x14 & n752 ;
  assign n837 = n836 ^ n835 ;
  assign n834 = x22 & n693 ;
  assign n838 = n837 ^ n834 ;
  assign n833 = x30 & n594 ;
  assign n839 = n838 ^ n833 ;
  assign n832 = x38 & n453 ;
  assign n840 = n839 ^ n832 ;
  assign n831 = x46 & n270 ;
  assign n841 = n840 ^ n831 ;
  assign n847 = x7 & n769 ;
  assign n846 = x15 & n752 ;
  assign n848 = n847 ^ n846 ;
  assign n845 = x23 & n693 ;
  assign n849 = n848 ^ n845 ;
  assign n844 = x31 & n594 ;
  assign n850 = n849 ^ n844 ;
  assign n843 = x39 & n453 ;
  assign n851 = n850 ^ n843 ;
  assign n842 = x47 & n270 ;
  assign n852 = n851 ^ n842 ;
  assign n868 = n766 & ~n767 ;
  assign n869 = ~n765 & n868 ;
  assign n870 = x0 & n869 ;
  assign n865 = ~n749 & ~n750 ;
  assign n866 = ~n748 & n865 ;
  assign n867 = x8 & n866 ;
  assign n871 = n870 ^ n867 ;
  assign n862 = n690 & n691 ;
  assign n863 = ~n689 & n862 ;
  assign n864 = x16 & n863 ;
  assign n872 = n871 ^ n864 ;
  assign n859 = ~n591 & n592 ;
  assign n860 = ~n590 & n859 ;
  assign n861 = x24 & n860 ;
  assign n873 = n872 ^ n861 ;
  assign n856 = n450 & ~n451 ;
  assign n857 = n449 & n856 ;
  assign n858 = x32 & n857 ;
  assign n874 = n873 ^ n858 ;
  assign n853 = ~n267 & ~n268 ;
  assign n854 = ~n266 & n853 ;
  assign n855 = x40 & n854 ;
  assign n875 = n874 ^ n855 ;
  assign n881 = x1 & n869 ;
  assign n880 = x9 & n866 ;
  assign n882 = n881 ^ n880 ;
  assign n879 = x17 & n863 ;
  assign n883 = n882 ^ n879 ;
  assign n878 = x25 & n860 ;
  assign n884 = n883 ^ n878 ;
  assign n877 = x33 & n857 ;
  assign n885 = n884 ^ n877 ;
  assign n876 = x41 & n854 ;
  assign n886 = n885 ^ n876 ;
  assign n892 = x2 & n869 ;
  assign n891 = x10 & n866 ;
  assign n893 = n892 ^ n891 ;
  assign n890 = x18 & n863 ;
  assign n894 = n893 ^ n890 ;
  assign n889 = x26 & n860 ;
  assign n895 = n894 ^ n889 ;
  assign n888 = x34 & n857 ;
  assign n896 = n895 ^ n888 ;
  assign n887 = x42 & n854 ;
  assign n897 = n896 ^ n887 ;
  assign n903 = x3 & n869 ;
  assign n902 = x11 & n866 ;
  assign n904 = n903 ^ n902 ;
  assign n901 = x19 & n863 ;
  assign n905 = n904 ^ n901 ;
  assign n900 = x27 & n860 ;
  assign n906 = n905 ^ n900 ;
  assign n899 = x35 & n857 ;
  assign n907 = n906 ^ n899 ;
  assign n898 = x43 & n854 ;
  assign n908 = n907 ^ n898 ;
  assign n914 = x4 & n869 ;
  assign n913 = x12 & n866 ;
  assign n915 = n914 ^ n913 ;
  assign n912 = x20 & n863 ;
  assign n916 = n915 ^ n912 ;
  assign n911 = x28 & n860 ;
  assign n917 = n916 ^ n911 ;
  assign n910 = x36 & n857 ;
  assign n918 = n917 ^ n910 ;
  assign n909 = x44 & n854 ;
  assign n919 = n918 ^ n909 ;
  assign n925 = x5 & n869 ;
  assign n924 = x13 & n866 ;
  assign n926 = n925 ^ n924 ;
  assign n923 = x21 & n863 ;
  assign n927 = n926 ^ n923 ;
  assign n922 = x29 & n860 ;
  assign n928 = n927 ^ n922 ;
  assign n921 = x37 & n857 ;
  assign n929 = n928 ^ n921 ;
  assign n920 = x45 & n854 ;
  assign n930 = n929 ^ n920 ;
  assign n936 = x6 & n869 ;
  assign n935 = x14 & n866 ;
  assign n937 = n936 ^ n935 ;
  assign n934 = x22 & n863 ;
  assign n938 = n937 ^ n934 ;
  assign n933 = x30 & n860 ;
  assign n939 = n938 ^ n933 ;
  assign n932 = x38 & n857 ;
  assign n940 = n939 ^ n932 ;
  assign n931 = x46 & n854 ;
  assign n941 = n940 ^ n931 ;
  assign n947 = x7 & n869 ;
  assign n946 = x15 & n866 ;
  assign n948 = n947 ^ n946 ;
  assign n945 = x23 & n863 ;
  assign n949 = n948 ^ n945 ;
  assign n944 = x31 & n860 ;
  assign n950 = n949 ^ n944 ;
  assign n943 = x39 & n857 ;
  assign n951 = n950 ^ n943 ;
  assign n942 = x47 & n854 ;
  assign n952 = n951 ^ n942 ;
  assign n968 = ~n766 & n767 ;
  assign n969 = ~n765 & n968 ;
  assign n970 = x0 & n969 ;
  assign n965 = n749 & n750 ;
  assign n966 = ~n748 & n965 ;
  assign n967 = x8 & n966 ;
  assign n971 = n970 ^ n967 ;
  assign n962 = ~n690 & ~n691 ;
  assign n963 = ~n689 & n962 ;
  assign n964 = x16 & n963 ;
  assign n972 = n971 ^ n964 ;
  assign n959 = n591 & ~n592 ;
  assign n960 = ~n590 & n959 ;
  assign n961 = x24 & n960 ;
  assign n973 = n972 ^ n961 ;
  assign n956 = ~n450 & n451 ;
  assign n957 = n449 & n956 ;
  assign n958 = x32 & n957 ;
  assign n974 = n973 ^ n958 ;
  assign n953 = n267 & n268 ;
  assign n954 = ~n266 & n953 ;
  assign n955 = x40 & n954 ;
  assign n975 = n974 ^ n955 ;
  assign n981 = x1 & n969 ;
  assign n980 = x9 & n966 ;
  assign n982 = n981 ^ n980 ;
  assign n979 = x17 & n963 ;
  assign n983 = n982 ^ n979 ;
  assign n978 = x25 & n960 ;
  assign n984 = n983 ^ n978 ;
  assign n977 = x33 & n957 ;
  assign n985 = n984 ^ n977 ;
  assign n976 = x41 & n954 ;
  assign n986 = n985 ^ n976 ;
  assign n992 = x2 & n969 ;
  assign n991 = x10 & n966 ;
  assign n993 = n992 ^ n991 ;
  assign n990 = x18 & n963 ;
  assign n994 = n993 ^ n990 ;
  assign n989 = x26 & n960 ;
  assign n995 = n994 ^ n989 ;
  assign n988 = x34 & n957 ;
  assign n996 = n995 ^ n988 ;
  assign n987 = x42 & n954 ;
  assign n997 = n996 ^ n987 ;
  assign n1003 = x3 & n969 ;
  assign n1002 = x11 & n966 ;
  assign n1004 = n1003 ^ n1002 ;
  assign n1001 = x19 & n963 ;
  assign n1005 = n1004 ^ n1001 ;
  assign n1000 = x27 & n960 ;
  assign n1006 = n1005 ^ n1000 ;
  assign n999 = x35 & n957 ;
  assign n1007 = n1006 ^ n999 ;
  assign n998 = x43 & n954 ;
  assign n1008 = n1007 ^ n998 ;
  assign n1014 = x4 & n969 ;
  assign n1013 = x12 & n966 ;
  assign n1015 = n1014 ^ n1013 ;
  assign n1012 = x20 & n963 ;
  assign n1016 = n1015 ^ n1012 ;
  assign n1011 = x28 & n960 ;
  assign n1017 = n1016 ^ n1011 ;
  assign n1010 = x36 & n957 ;
  assign n1018 = n1017 ^ n1010 ;
  assign n1009 = x44 & n954 ;
  assign n1019 = n1018 ^ n1009 ;
  assign n1025 = x5 & n969 ;
  assign n1024 = x13 & n966 ;
  assign n1026 = n1025 ^ n1024 ;
  assign n1023 = x21 & n963 ;
  assign n1027 = n1026 ^ n1023 ;
  assign n1022 = x29 & n960 ;
  assign n1028 = n1027 ^ n1022 ;
  assign n1021 = x37 & n957 ;
  assign n1029 = n1028 ^ n1021 ;
  assign n1020 = x45 & n954 ;
  assign n1030 = n1029 ^ n1020 ;
  assign n1036 = x6 & n969 ;
  assign n1035 = x14 & n966 ;
  assign n1037 = n1036 ^ n1035 ;
  assign n1034 = x22 & n963 ;
  assign n1038 = n1037 ^ n1034 ;
  assign n1033 = x30 & n960 ;
  assign n1039 = n1038 ^ n1033 ;
  assign n1032 = x38 & n957 ;
  assign n1040 = n1039 ^ n1032 ;
  assign n1031 = x46 & n954 ;
  assign n1041 = n1040 ^ n1031 ;
  assign n1047 = x7 & n969 ;
  assign n1046 = x15 & n966 ;
  assign n1048 = n1047 ^ n1046 ;
  assign n1045 = x23 & n963 ;
  assign n1049 = n1048 ^ n1045 ;
  assign n1044 = x31 & n960 ;
  assign n1050 = n1049 ^ n1044 ;
  assign n1043 = x39 & n957 ;
  assign n1051 = n1050 ^ n1043 ;
  assign n1042 = x47 & n954 ;
  assign n1052 = n1051 ^ n1042 ;
  assign n1068 = n766 & n767 ;
  assign n1069 = ~n765 & n1068 ;
  assign n1070 = x0 & n1069 ;
  assign n1065 = ~n749 & n750 ;
  assign n1066 = ~n748 & n1065 ;
  assign n1067 = x8 & n1066 ;
  assign n1071 = n1070 ^ n1067 ;
  assign n1062 = n690 & ~n691 ;
  assign n1063 = ~n689 & n1062 ;
  assign n1064 = x16 & n1063 ;
  assign n1072 = n1071 ^ n1064 ;
  assign n1059 = ~n591 & ~n592 ;
  assign n1060 = ~n590 & n1059 ;
  assign n1061 = x24 & n1060 ;
  assign n1073 = n1072 ^ n1061 ;
  assign n1056 = n450 & n451 ;
  assign n1057 = n449 & n1056 ;
  assign n1058 = x32 & n1057 ;
  assign n1074 = n1073 ^ n1058 ;
  assign n1053 = ~n267 & n268 ;
  assign n1054 = ~n266 & n1053 ;
  assign n1055 = x40 & n1054 ;
  assign n1075 = n1074 ^ n1055 ;
  assign n1081 = x1 & n1069 ;
  assign n1080 = x9 & n1066 ;
  assign n1082 = n1081 ^ n1080 ;
  assign n1079 = x17 & n1063 ;
  assign n1083 = n1082 ^ n1079 ;
  assign n1078 = x25 & n1060 ;
  assign n1084 = n1083 ^ n1078 ;
  assign n1077 = x33 & n1057 ;
  assign n1085 = n1084 ^ n1077 ;
  assign n1076 = x41 & n1054 ;
  assign n1086 = n1085 ^ n1076 ;
  assign n1092 = x2 & n1069 ;
  assign n1091 = x10 & n1066 ;
  assign n1093 = n1092 ^ n1091 ;
  assign n1090 = x18 & n1063 ;
  assign n1094 = n1093 ^ n1090 ;
  assign n1089 = x26 & n1060 ;
  assign n1095 = n1094 ^ n1089 ;
  assign n1088 = x34 & n1057 ;
  assign n1096 = n1095 ^ n1088 ;
  assign n1087 = x42 & n1054 ;
  assign n1097 = n1096 ^ n1087 ;
  assign n1103 = x3 & n1069 ;
  assign n1102 = x11 & n1066 ;
  assign n1104 = n1103 ^ n1102 ;
  assign n1101 = x19 & n1063 ;
  assign n1105 = n1104 ^ n1101 ;
  assign n1100 = x27 & n1060 ;
  assign n1106 = n1105 ^ n1100 ;
  assign n1099 = x35 & n1057 ;
  assign n1107 = n1106 ^ n1099 ;
  assign n1098 = x43 & n1054 ;
  assign n1108 = n1107 ^ n1098 ;
  assign n1114 = x4 & n1069 ;
  assign n1113 = x12 & n1066 ;
  assign n1115 = n1114 ^ n1113 ;
  assign n1112 = x20 & n1063 ;
  assign n1116 = n1115 ^ n1112 ;
  assign n1111 = x28 & n1060 ;
  assign n1117 = n1116 ^ n1111 ;
  assign n1110 = x36 & n1057 ;
  assign n1118 = n1117 ^ n1110 ;
  assign n1109 = x44 & n1054 ;
  assign n1119 = n1118 ^ n1109 ;
  assign n1125 = x5 & n1069 ;
  assign n1124 = x13 & n1066 ;
  assign n1126 = n1125 ^ n1124 ;
  assign n1123 = x21 & n1063 ;
  assign n1127 = n1126 ^ n1123 ;
  assign n1122 = x29 & n1060 ;
  assign n1128 = n1127 ^ n1122 ;
  assign n1121 = x37 & n1057 ;
  assign n1129 = n1128 ^ n1121 ;
  assign n1120 = x45 & n1054 ;
  assign n1130 = n1129 ^ n1120 ;
  assign n1136 = x6 & n1069 ;
  assign n1135 = x14 & n1066 ;
  assign n1137 = n1136 ^ n1135 ;
  assign n1134 = x22 & n1063 ;
  assign n1138 = n1137 ^ n1134 ;
  assign n1133 = x30 & n1060 ;
  assign n1139 = n1138 ^ n1133 ;
  assign n1132 = x38 & n1057 ;
  assign n1140 = n1139 ^ n1132 ;
  assign n1131 = x46 & n1054 ;
  assign n1141 = n1140 ^ n1131 ;
  assign n1147 = x7 & n1069 ;
  assign n1146 = x15 & n1066 ;
  assign n1148 = n1147 ^ n1146 ;
  assign n1145 = x23 & n1063 ;
  assign n1149 = n1148 ^ n1145 ;
  assign n1144 = x31 & n1060 ;
  assign n1150 = n1149 ^ n1144 ;
  assign n1143 = x39 & n1057 ;
  assign n1151 = n1150 ^ n1143 ;
  assign n1142 = x47 & n1054 ;
  assign n1152 = n1151 ^ n1142 ;
  assign n1163 = n765 & n768 ;
  assign n1164 = x0 & n1163 ;
  assign n1161 = n748 & n751 ;
  assign n1162 = x8 & n1161 ;
  assign n1165 = n1164 ^ n1162 ;
  assign n1159 = n689 & n692 ;
  assign n1160 = x16 & n1159 ;
  assign n1166 = n1165 ^ n1160 ;
  assign n1157 = n590 & n593 ;
  assign n1158 = x24 & n1157 ;
  assign n1167 = n1166 ^ n1158 ;
  assign n1155 = ~n449 & n452 ;
  assign n1156 = x32 & n1155 ;
  assign n1168 = n1167 ^ n1156 ;
  assign n1153 = n266 & n269 ;
  assign n1154 = x40 & n1153 ;
  assign n1169 = n1168 ^ n1154 ;
  assign n1175 = x1 & n1163 ;
  assign n1174 = x9 & n1161 ;
  assign n1176 = n1175 ^ n1174 ;
  assign n1173 = x17 & n1159 ;
  assign n1177 = n1176 ^ n1173 ;
  assign n1172 = x25 & n1157 ;
  assign n1178 = n1177 ^ n1172 ;
  assign n1171 = x33 & n1155 ;
  assign n1179 = n1178 ^ n1171 ;
  assign n1170 = x41 & n1153 ;
  assign n1180 = n1179 ^ n1170 ;
  assign n1186 = x2 & n1163 ;
  assign n1185 = x10 & n1161 ;
  assign n1187 = n1186 ^ n1185 ;
  assign n1184 = x18 & n1159 ;
  assign n1188 = n1187 ^ n1184 ;
  assign n1183 = x26 & n1157 ;
  assign n1189 = n1188 ^ n1183 ;
  assign n1182 = x34 & n1155 ;
  assign n1190 = n1189 ^ n1182 ;
  assign n1181 = x42 & n1153 ;
  assign n1191 = n1190 ^ n1181 ;
  assign n1197 = x3 & n1163 ;
  assign n1196 = x11 & n1161 ;
  assign n1198 = n1197 ^ n1196 ;
  assign n1195 = x19 & n1159 ;
  assign n1199 = n1198 ^ n1195 ;
  assign n1194 = x27 & n1157 ;
  assign n1200 = n1199 ^ n1194 ;
  assign n1193 = x35 & n1155 ;
  assign n1201 = n1200 ^ n1193 ;
  assign n1192 = x43 & n1153 ;
  assign n1202 = n1201 ^ n1192 ;
  assign n1208 = x4 & n1163 ;
  assign n1207 = x12 & n1161 ;
  assign n1209 = n1208 ^ n1207 ;
  assign n1206 = x20 & n1159 ;
  assign n1210 = n1209 ^ n1206 ;
  assign n1205 = x28 & n1157 ;
  assign n1211 = n1210 ^ n1205 ;
  assign n1204 = x36 & n1155 ;
  assign n1212 = n1211 ^ n1204 ;
  assign n1203 = x44 & n1153 ;
  assign n1213 = n1212 ^ n1203 ;
  assign n1219 = x5 & n1163 ;
  assign n1218 = x13 & n1161 ;
  assign n1220 = n1219 ^ n1218 ;
  assign n1217 = x21 & n1159 ;
  assign n1221 = n1220 ^ n1217 ;
  assign n1216 = x29 & n1157 ;
  assign n1222 = n1221 ^ n1216 ;
  assign n1215 = x37 & n1155 ;
  assign n1223 = n1222 ^ n1215 ;
  assign n1214 = x45 & n1153 ;
  assign n1224 = n1223 ^ n1214 ;
  assign n1230 = x6 & n1163 ;
  assign n1229 = x14 & n1161 ;
  assign n1231 = n1230 ^ n1229 ;
  assign n1228 = x22 & n1159 ;
  assign n1232 = n1231 ^ n1228 ;
  assign n1227 = x30 & n1157 ;
  assign n1233 = n1232 ^ n1227 ;
  assign n1226 = x38 & n1155 ;
  assign n1234 = n1233 ^ n1226 ;
  assign n1225 = x46 & n1153 ;
  assign n1235 = n1234 ^ n1225 ;
  assign n1241 = x7 & n1163 ;
  assign n1240 = x15 & n1161 ;
  assign n1242 = n1241 ^ n1240 ;
  assign n1239 = x23 & n1159 ;
  assign n1243 = n1242 ^ n1239 ;
  assign n1238 = x31 & n1157 ;
  assign n1244 = n1243 ^ n1238 ;
  assign n1237 = x39 & n1155 ;
  assign n1245 = n1244 ^ n1237 ;
  assign n1236 = x47 & n1153 ;
  assign n1246 = n1245 ^ n1236 ;
  assign n1257 = n765 & n868 ;
  assign n1258 = x0 & n1257 ;
  assign n1255 = n748 & n865 ;
  assign n1256 = x8 & n1255 ;
  assign n1259 = n1258 ^ n1256 ;
  assign n1253 = n689 & n862 ;
  assign n1254 = x16 & n1253 ;
  assign n1260 = n1259 ^ n1254 ;
  assign n1251 = n590 & n859 ;
  assign n1252 = x24 & n1251 ;
  assign n1261 = n1260 ^ n1252 ;
  assign n1249 = ~n449 & n856 ;
  assign n1250 = x32 & n1249 ;
  assign n1262 = n1261 ^ n1250 ;
  assign n1247 = n266 & n853 ;
  assign n1248 = x40 & n1247 ;
  assign n1263 = n1262 ^ n1248 ;
  assign n1269 = x1 & n1257 ;
  assign n1268 = x9 & n1255 ;
  assign n1270 = n1269 ^ n1268 ;
  assign n1267 = x17 & n1253 ;
  assign n1271 = n1270 ^ n1267 ;
  assign n1266 = x25 & n1251 ;
  assign n1272 = n1271 ^ n1266 ;
  assign n1265 = x33 & n1249 ;
  assign n1273 = n1272 ^ n1265 ;
  assign n1264 = x41 & n1247 ;
  assign n1274 = n1273 ^ n1264 ;
  assign n1280 = x2 & n1257 ;
  assign n1279 = x10 & n1255 ;
  assign n1281 = n1280 ^ n1279 ;
  assign n1278 = x18 & n1253 ;
  assign n1282 = n1281 ^ n1278 ;
  assign n1277 = x26 & n1251 ;
  assign n1283 = n1282 ^ n1277 ;
  assign n1276 = x34 & n1249 ;
  assign n1284 = n1283 ^ n1276 ;
  assign n1275 = x42 & n1247 ;
  assign n1285 = n1284 ^ n1275 ;
  assign n1291 = x3 & n1257 ;
  assign n1290 = x11 & n1255 ;
  assign n1292 = n1291 ^ n1290 ;
  assign n1289 = x19 & n1253 ;
  assign n1293 = n1292 ^ n1289 ;
  assign n1288 = x27 & n1251 ;
  assign n1294 = n1293 ^ n1288 ;
  assign n1287 = x35 & n1249 ;
  assign n1295 = n1294 ^ n1287 ;
  assign n1286 = x43 & n1247 ;
  assign n1296 = n1295 ^ n1286 ;
  assign n1302 = x4 & n1257 ;
  assign n1301 = x12 & n1255 ;
  assign n1303 = n1302 ^ n1301 ;
  assign n1300 = x20 & n1253 ;
  assign n1304 = n1303 ^ n1300 ;
  assign n1299 = x28 & n1251 ;
  assign n1305 = n1304 ^ n1299 ;
  assign n1298 = x36 & n1249 ;
  assign n1306 = n1305 ^ n1298 ;
  assign n1297 = x44 & n1247 ;
  assign n1307 = n1306 ^ n1297 ;
  assign n1313 = x5 & n1257 ;
  assign n1312 = x13 & n1255 ;
  assign n1314 = n1313 ^ n1312 ;
  assign n1311 = x21 & n1253 ;
  assign n1315 = n1314 ^ n1311 ;
  assign n1310 = x29 & n1251 ;
  assign n1316 = n1315 ^ n1310 ;
  assign n1309 = x37 & n1249 ;
  assign n1317 = n1316 ^ n1309 ;
  assign n1308 = x45 & n1247 ;
  assign n1318 = n1317 ^ n1308 ;
  assign n1324 = x6 & n1257 ;
  assign n1323 = x14 & n1255 ;
  assign n1325 = n1324 ^ n1323 ;
  assign n1322 = x22 & n1253 ;
  assign n1326 = n1325 ^ n1322 ;
  assign n1321 = x30 & n1251 ;
  assign n1327 = n1326 ^ n1321 ;
  assign n1320 = x38 & n1249 ;
  assign n1328 = n1327 ^ n1320 ;
  assign n1319 = x46 & n1247 ;
  assign n1329 = n1328 ^ n1319 ;
  assign n1335 = x7 & n1257 ;
  assign n1334 = x15 & n1255 ;
  assign n1336 = n1335 ^ n1334 ;
  assign n1333 = x23 & n1253 ;
  assign n1337 = n1336 ^ n1333 ;
  assign n1332 = x31 & n1251 ;
  assign n1338 = n1337 ^ n1332 ;
  assign n1331 = x39 & n1249 ;
  assign n1339 = n1338 ^ n1331 ;
  assign n1330 = x47 & n1247 ;
  assign n1340 = n1339 ^ n1330 ;
  assign y0 = n775 ;
  assign y1 = n786 ;
  assign y2 = n797 ;
  assign y3 = n808 ;
  assign y4 = n819 ;
  assign y5 = n830 ;
  assign y6 = n841 ;
  assign y7 = n852 ;
  assign y8 = n875 ;
  assign y9 = n886 ;
  assign y10 = n897 ;
  assign y11 = n908 ;
  assign y12 = n919 ;
  assign y13 = n930 ;
  assign y14 = n941 ;
  assign y15 = n952 ;
  assign y16 = n975 ;
  assign y17 = n986 ;
  assign y18 = n997 ;
  assign y19 = n1008 ;
  assign y20 = n1019 ;
  assign y21 = n1030 ;
  assign y22 = n1041 ;
  assign y23 = n1052 ;
  assign y24 = n1075 ;
  assign y25 = n1086 ;
  assign y26 = n1097 ;
  assign y27 = n1108 ;
  assign y28 = n1119 ;
  assign y29 = n1130 ;
  assign y30 = n1141 ;
  assign y31 = n1152 ;
  assign y32 = n1169 ;
  assign y33 = n1180 ;
  assign y34 = n1191 ;
  assign y35 = n1202 ;
  assign y36 = n1213 ;
  assign y37 = n1224 ;
  assign y38 = n1235 ;
  assign y39 = n1246 ;
  assign y40 = n1263 ;
  assign y41 = n1274 ;
  assign y42 = n1285 ;
  assign y43 = n1296 ;
  assign y44 = n1307 ;
  assign y45 = n1318 ;
  assign y46 = n1329 ;
  assign y47 = n1340 ;
endmodule
