module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 ;
  assign n18 = x9 ^ x1 ;
  assign n17 = x0 & x8 ;
  assign n19 = n18 ^ n17 ;
  assign n22 = x10 ^ x2 ;
  assign n21 = x1 & x9 ;
  assign n23 = n22 ^ n21 ;
  assign n20 = n17 & n18 ;
  assign n24 = n23 ^ n20 ;
  assign n33 = x11 ^ x3 ;
  assign n32 = x2 & x10 ;
  assign n34 = n33 ^ n32 ;
  assign n30 = n21 & n22 ;
  assign n27 = ~x1 & n22 ;
  assign n28 = n17 & n27 ;
  assign n25 = ~x9 & n22 ;
  assign n26 = n17 & n25 ;
  assign n29 = n28 ^ n26 ;
  assign n31 = n30 ^ n29 ;
  assign n35 = n34 ^ n31 ;
  assign n40 = x12 ^ x4 ;
  assign n39 = x3 & x11 ;
  assign n41 = n40 ^ n39 ;
  assign n37 = n31 & n34 ;
  assign n36 = n32 & n33 ;
  assign n38 = n37 ^ n36 ;
  assign n42 = n41 ^ n38 ;
  assign n50 = x13 ^ x5 ;
  assign n49 = x4 & x12 ;
  assign n51 = n50 ^ n49 ;
  assign n46 = n36 & n41 ;
  assign n45 = n39 & n40 ;
  assign n47 = n46 ^ n45 ;
  assign n43 = n34 & n41 ;
  assign n44 = n31 & n43 ;
  assign n48 = n47 ^ n44 ;
  assign n52 = n51 ^ n48 ;
  assign n57 = x14 ^ x6 ;
  assign n56 = x5 & x13 ;
  assign n58 = n57 ^ n56 ;
  assign n54 = n48 & n51 ;
  assign n53 = n49 & n50 ;
  assign n55 = n54 ^ n53 ;
  assign n59 = n58 ^ n55 ;
  assign n67 = x15 ^ x7 ;
  assign n66 = x6 & x14 ;
  assign n68 = n67 ^ n66 ;
  assign n63 = n53 & n58 ;
  assign n62 = n56 & n57 ;
  assign n64 = n63 ^ n62 ;
  assign n60 = n51 & n58 ;
  assign n61 = n48 & n60 ;
  assign n65 = n64 ^ n61 ;
  assign n69 = n68 ^ n65 ;
  assign n76 = x7 & x15 ;
  assign n77 = n76 ^ n67 ;
  assign n73 = n64 & n68 ;
  assign n72 = n66 & n67 ;
  assign n74 = n73 ^ n72 ;
  assign n70 = n60 & n68 ;
  assign n71 = n48 & n70 ;
  assign n75 = n74 ^ n71 ;
  assign n78 = n77 ^ n75 ;
  assign y0 = n19 ;
  assign y1 = n24 ;
  assign y2 = n35 ;
  assign y3 = n42 ;
  assign y4 = n52 ;
  assign y5 = n59 ;
  assign y6 = n69 ;
  assign y7 = n78 ;
endmodule
