module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 ;
  assign n68 = x8 ^ x0 ;
  assign n69 = x9 ^ x1 ;
  assign n70 = n68 & n69 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = x10 ^ x2 ;
  assign n103 = x3 & x11 ;
  assign n104 = n103 ^ x3 ;
  assign n105 = n73 & n104 ;
  assign n106 = n105 ^ n104 ;
  assign n102 = x2 & ~x10 ;
  assign n107 = n106 ^ n102 ;
  assign n388 = ~n72 & n107 ;
  assign n98 = x1 & ~x9 ;
  assign n99 = ~n68 & n98 ;
  assign n97 = x0 & ~x8 ;
  assign n100 = n99 ^ n97 ;
  assign n389 = n388 ^ n100 ;
  assign n50 = x12 ^ x4 ;
  assign n54 = x13 ^ x5 ;
  assign n55 = n50 & n54 ;
  assign n56 = n55 ^ n50 ;
  assign n57 = n56 ^ n54 ;
  assign n59 = x14 ^ x6 ;
  assign n60 = x7 & x15 ;
  assign n61 = n60 ^ x7 ;
  assign n62 = n59 & n61 ;
  assign n63 = n62 ^ n61 ;
  assign n58 = x6 & ~x14 ;
  assign n64 = n63 ^ n58 ;
  assign n65 = n57 & n64 ;
  assign n66 = n65 ^ n64 ;
  assign n51 = x5 & ~x13 ;
  assign n52 = ~n50 & n51 ;
  assign n49 = x4 & ~x12 ;
  assign n53 = n52 ^ n49 ;
  assign n67 = n66 ^ n53 ;
  assign n74 = x11 ^ x3 ;
  assign n75 = n73 & n74 ;
  assign n76 = n75 ^ n73 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = n72 & n77 ;
  assign n79 = n78 ^ n72 ;
  assign n80 = n79 ^ n77 ;
  assign n387 = n67 & ~n80 ;
  assign n390 = n389 ^ n387 ;
  assign n84 = x15 ^ x7 ;
  assign n85 = n59 & n84 ;
  assign n86 = n85 ^ n59 ;
  assign n87 = n86 ^ n84 ;
  assign n88 = n57 & n87 ;
  assign n89 = n88 ^ n57 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = n80 & n90 ;
  assign n92 = n91 ^ n80 ;
  assign n93 = n92 ^ n90 ;
  assign n391 = n390 ^ n93 ;
  assign n460 = x10 & ~n391 ;
  assign n459 = x2 & n391 ;
  assign n461 = n460 ^ n459 ;
  assign n120 = x4 & ~n72 ;
  assign n121 = n107 & n120 ;
  assign n119 = x4 & n100 ;
  assign n122 = n121 ^ n119 ;
  assign n123 = n122 ^ x4 ;
  assign n116 = x4 & n93 ;
  assign n117 = n116 ^ x4 ;
  assign n118 = n117 ^ x4 ;
  assign n124 = n123 ^ n118 ;
  assign n113 = x4 & n80 ;
  assign n114 = n113 ^ x4 ;
  assign n115 = n67 & n114 ;
  assign n125 = n124 ^ n115 ;
  assign n108 = x12 & ~n72 ;
  assign n109 = n107 & n108 ;
  assign n101 = x12 & n100 ;
  assign n110 = n109 ^ n101 ;
  assign n94 = x12 & n93 ;
  assign n95 = n94 ^ x12 ;
  assign n96 = n95 ^ x12 ;
  assign n111 = n110 ^ n96 ;
  assign n81 = x12 & n80 ;
  assign n82 = n81 ^ x12 ;
  assign n83 = n67 & n82 ;
  assign n112 = n111 ^ n83 ;
  assign n126 = n125 ^ n112 ;
  assign n244 = n126 ^ x20 ;
  assign n264 = x5 & ~n72 ;
  assign n265 = n107 & n264 ;
  assign n263 = x5 & n100 ;
  assign n266 = n265 ^ n263 ;
  assign n267 = n266 ^ x5 ;
  assign n260 = x5 & n93 ;
  assign n261 = n260 ^ x5 ;
  assign n262 = n261 ^ x5 ;
  assign n268 = n267 ^ n262 ;
  assign n257 = x5 & n80 ;
  assign n258 = n257 ^ x5 ;
  assign n259 = n67 & n258 ;
  assign n269 = n268 ^ n259 ;
  assign n252 = x13 & ~n72 ;
  assign n253 = n107 & n252 ;
  assign n251 = x13 & n100 ;
  assign n254 = n253 ^ n251 ;
  assign n248 = x13 & n93 ;
  assign n249 = n248 ^ x13 ;
  assign n250 = n249 ^ x13 ;
  assign n255 = n254 ^ n250 ;
  assign n245 = x13 & n80 ;
  assign n246 = n245 ^ x13 ;
  assign n247 = n67 & n246 ;
  assign n256 = n255 ^ n247 ;
  assign n270 = n269 ^ n256 ;
  assign n271 = n270 ^ x21 ;
  assign n272 = n244 & n271 ;
  assign n273 = n272 ^ n244 ;
  assign n274 = n273 ^ n271 ;
  assign n294 = x6 & ~n72 ;
  assign n295 = n107 & n294 ;
  assign n293 = x6 & n100 ;
  assign n296 = n295 ^ n293 ;
  assign n297 = n296 ^ x6 ;
  assign n290 = x6 & n93 ;
  assign n291 = n290 ^ x6 ;
  assign n292 = n291 ^ x6 ;
  assign n298 = n297 ^ n292 ;
  assign n287 = x6 & n80 ;
  assign n288 = n287 ^ x6 ;
  assign n289 = n67 & n288 ;
  assign n299 = n298 ^ n289 ;
  assign n282 = x14 & ~n72 ;
  assign n283 = n107 & n282 ;
  assign n281 = x14 & n100 ;
  assign n284 = n283 ^ n281 ;
  assign n278 = x14 & n93 ;
  assign n279 = n278 ^ x14 ;
  assign n280 = n279 ^ x14 ;
  assign n285 = n284 ^ n280 ;
  assign n275 = x14 & n80 ;
  assign n276 = n275 ^ x14 ;
  assign n277 = n67 & n276 ;
  assign n286 = n285 ^ n277 ;
  assign n300 = n299 ^ n286 ;
  assign n301 = n300 ^ x22 ;
  assign n322 = x7 & ~n72 ;
  assign n323 = n107 & n322 ;
  assign n321 = x7 & ~n100 ;
  assign n324 = n323 ^ n321 ;
  assign n318 = x7 & n93 ;
  assign n319 = n318 ^ x7 ;
  assign n320 = n319 ^ x7 ;
  assign n325 = n324 ^ n320 ;
  assign n315 = x7 & n80 ;
  assign n316 = n315 ^ x7 ;
  assign n317 = n67 & n316 ;
  assign n326 = n325 ^ n317 ;
  assign n309 = x15 & ~n72 ;
  assign n310 = n107 & n309 ;
  assign n308 = x15 & ~n100 ;
  assign n311 = n310 ^ n308 ;
  assign n305 = x15 & n93 ;
  assign n306 = n305 ^ x15 ;
  assign n307 = n306 ^ x15 ;
  assign n312 = n311 ^ n307 ;
  assign n302 = x15 & n80 ;
  assign n303 = n302 ^ x15 ;
  assign n304 = n67 & n303 ;
  assign n313 = n312 ^ n304 ;
  assign n314 = n313 ^ x15 ;
  assign n327 = n326 ^ n314 ;
  assign n361 = x23 & n327 ;
  assign n362 = n361 ^ n327 ;
  assign n363 = n301 & n362 ;
  assign n364 = n363 ^ n362 ;
  assign n360 = ~x22 & n300 ;
  assign n365 = n364 ^ n360 ;
  assign n366 = n274 & n365 ;
  assign n367 = n366 ^ n365 ;
  assign n357 = ~x21 & n270 ;
  assign n358 = ~n244 & n357 ;
  assign n356 = ~x20 & n126 ;
  assign n359 = n358 ^ n356 ;
  assign n368 = n367 ^ n359 ;
  assign n146 = x0 & ~n72 ;
  assign n147 = n107 & n146 ;
  assign n145 = x0 & n100 ;
  assign n148 = n147 ^ n145 ;
  assign n149 = n148 ^ x0 ;
  assign n142 = x0 & n93 ;
  assign n143 = n142 ^ x0 ;
  assign n144 = n143 ^ x0 ;
  assign n150 = n149 ^ n144 ;
  assign n139 = x0 & n80 ;
  assign n140 = n139 ^ x0 ;
  assign n141 = n67 & n140 ;
  assign n151 = n150 ^ n141 ;
  assign n134 = x8 & ~n72 ;
  assign n135 = n107 & n134 ;
  assign n133 = x8 & n100 ;
  assign n136 = n135 ^ n133 ;
  assign n130 = x8 & n93 ;
  assign n131 = n130 ^ x8 ;
  assign n132 = n131 ^ x8 ;
  assign n137 = n136 ^ n132 ;
  assign n127 = x8 & n80 ;
  assign n128 = n127 ^ x8 ;
  assign n129 = n67 & n128 ;
  assign n138 = n137 ^ n129 ;
  assign n152 = n151 ^ n138 ;
  assign n153 = n152 ^ x16 ;
  assign n173 = x1 & ~n72 ;
  assign n174 = n107 & n173 ;
  assign n172 = x1 & n100 ;
  assign n175 = n174 ^ n172 ;
  assign n176 = n175 ^ x1 ;
  assign n169 = x1 & n93 ;
  assign n170 = n169 ^ x1 ;
  assign n171 = n170 ^ x1 ;
  assign n177 = n176 ^ n171 ;
  assign n166 = x1 & n80 ;
  assign n167 = n166 ^ x1 ;
  assign n168 = n67 & n167 ;
  assign n178 = n177 ^ n168 ;
  assign n161 = x9 & ~n72 ;
  assign n162 = n107 & n161 ;
  assign n160 = x9 & n100 ;
  assign n163 = n162 ^ n160 ;
  assign n157 = x9 & n93 ;
  assign n158 = n157 ^ x9 ;
  assign n159 = n158 ^ x9 ;
  assign n164 = n163 ^ n159 ;
  assign n154 = x9 & n80 ;
  assign n155 = n154 ^ x9 ;
  assign n156 = n67 & n155 ;
  assign n165 = n164 ^ n156 ;
  assign n179 = n178 ^ n165 ;
  assign n180 = n179 ^ x17 ;
  assign n181 = n153 & n180 ;
  assign n182 = n181 ^ n153 ;
  assign n183 = n182 ^ n180 ;
  assign n203 = x2 & ~n72 ;
  assign n204 = n107 & n203 ;
  assign n202 = x2 & n100 ;
  assign n205 = n204 ^ n202 ;
  assign n206 = n205 ^ x2 ;
  assign n199 = x2 & n93 ;
  assign n200 = n199 ^ x2 ;
  assign n201 = n200 ^ x2 ;
  assign n207 = n206 ^ n201 ;
  assign n196 = x2 & n80 ;
  assign n197 = n196 ^ x2 ;
  assign n198 = n67 & n197 ;
  assign n208 = n207 ^ n198 ;
  assign n191 = x10 & ~n72 ;
  assign n192 = n107 & n191 ;
  assign n190 = x10 & n100 ;
  assign n193 = n192 ^ n190 ;
  assign n187 = x10 & n93 ;
  assign n188 = n187 ^ x10 ;
  assign n189 = n188 ^ x10 ;
  assign n194 = n193 ^ n189 ;
  assign n184 = x10 & n80 ;
  assign n185 = n184 ^ x10 ;
  assign n186 = n67 & n185 ;
  assign n195 = n194 ^ n186 ;
  assign n209 = n208 ^ n195 ;
  assign n210 = n209 ^ x18 ;
  assign n230 = x3 & ~n72 ;
  assign n231 = n107 & n230 ;
  assign n229 = x3 & n100 ;
  assign n232 = n231 ^ n229 ;
  assign n233 = n232 ^ x3 ;
  assign n226 = x3 & n93 ;
  assign n227 = n226 ^ x3 ;
  assign n228 = n227 ^ x3 ;
  assign n234 = n233 ^ n228 ;
  assign n223 = x3 & n80 ;
  assign n224 = n223 ^ x3 ;
  assign n225 = n67 & n224 ;
  assign n235 = n234 ^ n225 ;
  assign n218 = x11 & ~n72 ;
  assign n219 = n107 & n218 ;
  assign n217 = x11 & n100 ;
  assign n220 = n219 ^ n217 ;
  assign n214 = x11 & n93 ;
  assign n215 = n214 ^ x11 ;
  assign n216 = n215 ^ x11 ;
  assign n221 = n220 ^ n216 ;
  assign n211 = x11 & n80 ;
  assign n212 = n211 ^ x11 ;
  assign n213 = n67 & n212 ;
  assign n222 = n221 ^ n213 ;
  assign n236 = n235 ^ n222 ;
  assign n237 = n236 ^ x19 ;
  assign n238 = n210 & n237 ;
  assign n239 = n238 ^ n210 ;
  assign n240 = n239 ^ n237 ;
  assign n241 = n183 & n240 ;
  assign n242 = n241 ^ n183 ;
  assign n243 = n242 ^ n240 ;
  assign n416 = x16 & n243 ;
  assign n417 = n416 ^ x16 ;
  assign n418 = n368 & n417 ;
  assign n328 = n327 ^ x23 ;
  assign n329 = n301 & n328 ;
  assign n330 = n329 ^ n301 ;
  assign n331 = n330 ^ n328 ;
  assign n332 = n274 & n331 ;
  assign n333 = n332 ^ n274 ;
  assign n334 = n333 ^ n331 ;
  assign n335 = n243 & n334 ;
  assign n336 = n335 ^ n243 ;
  assign n337 = n336 ^ n334 ;
  assign n412 = x16 & n337 ;
  assign n413 = n412 ^ x16 ;
  assign n414 = n413 ^ x16 ;
  assign n347 = x19 & n236 ;
  assign n348 = n347 ^ n236 ;
  assign n349 = n210 & n348 ;
  assign n350 = n349 ^ n348 ;
  assign n346 = ~x18 & n209 ;
  assign n351 = n350 ^ n346 ;
  assign n408 = x16 & ~n183 ;
  assign n409 = n351 & n408 ;
  assign n342 = ~x17 & n179 ;
  assign n343 = ~n153 & n342 ;
  assign n341 = ~x16 & n152 ;
  assign n344 = n343 ^ n341 ;
  assign n407 = x16 & n344 ;
  assign n410 = n409 ^ n407 ;
  assign n411 = n410 ^ x16 ;
  assign n415 = n414 ^ n411 ;
  assign n419 = n418 ^ n415 ;
  assign n403 = n152 & n243 ;
  assign n404 = n403 ^ n152 ;
  assign n405 = n368 & n404 ;
  assign n399 = n152 & ~n183 ;
  assign n400 = n351 & n399 ;
  assign n398 = n152 & n344 ;
  assign n401 = n400 ^ n398 ;
  assign n395 = n152 & n337 ;
  assign n396 = n395 ^ n152 ;
  assign n397 = n396 ^ n152 ;
  assign n402 = n401 ^ n397 ;
  assign n406 = n405 ^ n402 ;
  assign n420 = n419 ^ n406 ;
  assign n393 = x8 & ~n391 ;
  assign n392 = x0 & n391 ;
  assign n394 = n393 ^ n392 ;
  assign n422 = n420 ^ n394 ;
  assign n450 = x9 & ~n391 ;
  assign n449 = x1 & n391 ;
  assign n451 = n450 ^ n449 ;
  assign n444 = x17 & n243 ;
  assign n445 = n444 ^ x17 ;
  assign n446 = n368 & n445 ;
  assign n440 = x17 & n337 ;
  assign n441 = n440 ^ x17 ;
  assign n442 = n441 ^ x17 ;
  assign n436 = x17 & ~n183 ;
  assign n437 = n351 & n436 ;
  assign n435 = x17 & n344 ;
  assign n438 = n437 ^ n435 ;
  assign n439 = n438 ^ x17 ;
  assign n443 = n442 ^ n439 ;
  assign n447 = n446 ^ n443 ;
  assign n431 = n179 & n243 ;
  assign n432 = n431 ^ n179 ;
  assign n433 = n368 & n432 ;
  assign n427 = n179 & ~n183 ;
  assign n428 = n351 & n427 ;
  assign n426 = n179 & n344 ;
  assign n429 = n428 ^ n426 ;
  assign n423 = n179 & n337 ;
  assign n424 = n423 ^ n179 ;
  assign n425 = n424 ^ n179 ;
  assign n430 = n429 ^ n425 ;
  assign n434 = n433 ^ n430 ;
  assign n448 = n447 ^ n434 ;
  assign n455 = n451 ^ n448 ;
  assign n456 = n422 & n455 ;
  assign n457 = n456 ^ n422 ;
  assign n458 = n457 ^ n455 ;
  assign n483 = x18 & n243 ;
  assign n484 = n483 ^ x18 ;
  assign n485 = n368 & n484 ;
  assign n479 = x18 & n337 ;
  assign n480 = n479 ^ x18 ;
  assign n481 = n480 ^ x18 ;
  assign n475 = x18 & ~n183 ;
  assign n476 = n351 & n475 ;
  assign n474 = x18 & n344 ;
  assign n477 = n476 ^ n474 ;
  assign n478 = n477 ^ x18 ;
  assign n482 = n481 ^ n478 ;
  assign n486 = n485 ^ n482 ;
  assign n470 = n209 & n243 ;
  assign n471 = n470 ^ n209 ;
  assign n472 = n368 & n471 ;
  assign n466 = ~n183 & n209 ;
  assign n467 = n351 & n466 ;
  assign n465 = n209 & n344 ;
  assign n468 = n467 ^ n465 ;
  assign n462 = n209 & n337 ;
  assign n463 = n462 ^ n209 ;
  assign n464 = n463 ^ n209 ;
  assign n469 = n468 ^ n464 ;
  assign n473 = n472 ^ n469 ;
  assign n487 = n486 ^ n473 ;
  assign n489 = n487 ^ n461 ;
  assign n514 = x19 & n243 ;
  assign n515 = n514 ^ x19 ;
  assign n516 = n368 & n515 ;
  assign n510 = x19 & n337 ;
  assign n511 = n510 ^ x19 ;
  assign n512 = n511 ^ x19 ;
  assign n506 = x19 & ~n183 ;
  assign n507 = n351 & n506 ;
  assign n505 = x19 & n344 ;
  assign n508 = n507 ^ n505 ;
  assign n509 = n508 ^ x19 ;
  assign n513 = n512 ^ n509 ;
  assign n517 = n516 ^ n513 ;
  assign n501 = n236 & n243 ;
  assign n502 = n501 ^ n236 ;
  assign n503 = n368 & n502 ;
  assign n497 = ~n183 & n236 ;
  assign n498 = n351 & n497 ;
  assign n496 = n236 & n344 ;
  assign n499 = n498 ^ n496 ;
  assign n493 = n236 & n337 ;
  assign n494 = n493 ^ n236 ;
  assign n495 = n494 ^ n236 ;
  assign n500 = n499 ^ n495 ;
  assign n504 = n503 ^ n500 ;
  assign n518 = n517 ^ n504 ;
  assign n491 = x11 & ~n391 ;
  assign n490 = x3 & n391 ;
  assign n492 = n491 ^ n490 ;
  assign n527 = n518 ^ n492 ;
  assign n528 = n489 & n527 ;
  assign n529 = n528 ^ n489 ;
  assign n530 = n529 ^ n527 ;
  assign n531 = n458 & n530 ;
  assign n532 = n531 ^ n458 ;
  assign n533 = n532 ^ n530 ;
  assign n535 = x12 & ~n391 ;
  assign n534 = x4 & n391 ;
  assign n536 = n535 ^ n534 ;
  assign n382 = x20 & n243 ;
  assign n383 = n382 ^ x20 ;
  assign n384 = n368 & n383 ;
  assign n378 = x20 & n337 ;
  assign n379 = n378 ^ x20 ;
  assign n380 = n379 ^ x20 ;
  assign n374 = x20 & ~n183 ;
  assign n375 = n351 & n374 ;
  assign n373 = x20 & n344 ;
  assign n376 = n375 ^ n373 ;
  assign n377 = n376 ^ x20 ;
  assign n381 = n380 ^ n377 ;
  assign n385 = n384 ^ n381 ;
  assign n369 = n126 & n243 ;
  assign n370 = n369 ^ n126 ;
  assign n371 = n368 & n370 ;
  assign n352 = n126 & ~n183 ;
  assign n353 = n351 & n352 ;
  assign n345 = n126 & n344 ;
  assign n354 = n353 ^ n345 ;
  assign n338 = n126 & n337 ;
  assign n339 = n338 ^ n126 ;
  assign n340 = n339 ^ n126 ;
  assign n355 = n354 ^ n340 ;
  assign n372 = n371 ^ n355 ;
  assign n386 = n385 ^ n372 ;
  assign n538 = n536 ^ n386 ;
  assign n563 = x21 & n243 ;
  assign n564 = n563 ^ x21 ;
  assign n565 = n368 & n564 ;
  assign n559 = x21 & n337 ;
  assign n560 = n559 ^ x21 ;
  assign n561 = n560 ^ x21 ;
  assign n555 = x21 & ~n183 ;
  assign n556 = n351 & n555 ;
  assign n554 = x21 & n344 ;
  assign n557 = n556 ^ n554 ;
  assign n558 = n557 ^ x21 ;
  assign n562 = n561 ^ n558 ;
  assign n566 = n565 ^ n562 ;
  assign n550 = n243 & n270 ;
  assign n551 = n550 ^ n270 ;
  assign n552 = n368 & n551 ;
  assign n546 = ~n183 & n270 ;
  assign n547 = n351 & n546 ;
  assign n545 = n270 & n344 ;
  assign n548 = n547 ^ n545 ;
  assign n542 = n270 & n337 ;
  assign n543 = n542 ^ n270 ;
  assign n544 = n543 ^ n270 ;
  assign n549 = n548 ^ n544 ;
  assign n553 = n552 ^ n549 ;
  assign n567 = n566 ^ n553 ;
  assign n540 = x13 & ~n391 ;
  assign n539 = x5 & n391 ;
  assign n541 = n540 ^ n539 ;
  assign n573 = n567 ^ n541 ;
  assign n574 = n538 & n573 ;
  assign n575 = n574 ^ n538 ;
  assign n576 = n575 ^ n573 ;
  assign n601 = x22 & n243 ;
  assign n602 = n601 ^ x22 ;
  assign n603 = n368 & n602 ;
  assign n597 = x22 & n337 ;
  assign n598 = n597 ^ x22 ;
  assign n599 = n598 ^ x22 ;
  assign n593 = x22 & ~n183 ;
  assign n594 = n351 & n593 ;
  assign n592 = x22 & n344 ;
  assign n595 = n594 ^ n592 ;
  assign n596 = n595 ^ x22 ;
  assign n600 = n599 ^ n596 ;
  assign n604 = n603 ^ n600 ;
  assign n588 = n243 & n300 ;
  assign n589 = n588 ^ n300 ;
  assign n590 = n368 & n589 ;
  assign n584 = ~n183 & n300 ;
  assign n585 = n351 & n584 ;
  assign n583 = n300 & n344 ;
  assign n586 = n585 ^ n583 ;
  assign n580 = n300 & n337 ;
  assign n581 = n580 ^ n300 ;
  assign n582 = n581 ^ n300 ;
  assign n587 = n586 ^ n582 ;
  assign n591 = n590 ^ n587 ;
  assign n605 = n604 ^ n591 ;
  assign n578 = x14 & ~n391 ;
  assign n577 = x6 & n391 ;
  assign n579 = n578 ^ n577 ;
  assign n608 = n605 ^ n579 ;
  assign n673 = x23 & ~n183 ;
  assign n674 = n351 & n673 ;
  assign n672 = x23 & n344 ;
  assign n675 = n674 ^ n672 ;
  assign n676 = n675 ^ x23 ;
  assign n669 = x23 & n337 ;
  assign n670 = n669 ^ x23 ;
  assign n671 = n670 ^ x23 ;
  assign n677 = n676 ^ n671 ;
  assign n666 = x23 & n243 ;
  assign n667 = n666 ^ x23 ;
  assign n668 = n368 & n667 ;
  assign n678 = n677 ^ n668 ;
  assign n659 = ~n183 & n327 ;
  assign n660 = n351 & n659 ;
  assign n658 = n327 & n344 ;
  assign n661 = n660 ^ n658 ;
  assign n662 = n661 ^ n327 ;
  assign n655 = n327 & n337 ;
  assign n656 = n655 ^ n327 ;
  assign n657 = n656 ^ n327 ;
  assign n663 = n662 ^ n657 ;
  assign n652 = n243 & n327 ;
  assign n653 = n652 ^ n327 ;
  assign n654 = n368 & n653 ;
  assign n664 = n663 ^ n654 ;
  assign n665 = n664 ^ n327 ;
  assign n679 = n678 ^ n665 ;
  assign n609 = x7 & ~n389 ;
  assign n610 = n609 ^ n318 ;
  assign n611 = n610 ^ n317 ;
  assign n612 = n611 ^ x7 ;
  assign n613 = n612 ^ n313 ;
  assign n680 = n679 ^ n613 ;
  assign n681 = n608 & n680 ;
  assign n682 = n681 ^ n608 ;
  assign n683 = n682 ^ n680 ;
  assign n684 = n576 & n683 ;
  assign n685 = n684 ^ n576 ;
  assign n686 = n685 ^ n683 ;
  assign n687 = n533 & n686 ;
  assign n688 = n687 ^ n533 ;
  assign n689 = n688 ^ n686 ;
  assign n627 = x23 & n613 ;
  assign n635 = ~n183 & n627 ;
  assign n636 = n351 & n635 ;
  assign n634 = n344 & n627 ;
  assign n637 = n636 ^ n634 ;
  assign n638 = n637 ^ n627 ;
  assign n631 = n337 & n627 ;
  assign n632 = n631 ^ n627 ;
  assign n633 = n632 ^ n627 ;
  assign n639 = n638 ^ n633 ;
  assign n628 = n243 & n627 ;
  assign n629 = n628 ^ n627 ;
  assign n630 = n368 & n629 ;
  assign n640 = n639 ^ n630 ;
  assign n614 = n327 & n613 ;
  assign n622 = ~n183 & n614 ;
  assign n623 = n351 & n622 ;
  assign n621 = n344 & n614 ;
  assign n624 = n623 ^ n621 ;
  assign n618 = n337 & n614 ;
  assign n619 = n618 ^ n614 ;
  assign n620 = n619 ^ n614 ;
  assign n625 = n624 ^ n620 ;
  assign n615 = n243 & n614 ;
  assign n616 = n615 ^ n614 ;
  assign n617 = n368 & n616 ;
  assign n626 = n625 ^ n617 ;
  assign n641 = n640 ^ n626 ;
  assign n642 = n641 ^ n613 ;
  assign n643 = n608 & n642 ;
  assign n644 = n643 ^ n642 ;
  assign n606 = n579 & n605 ;
  assign n607 = n606 ^ n579 ;
  assign n645 = n644 ^ n607 ;
  assign n646 = n576 & n645 ;
  assign n647 = n646 ^ n645 ;
  assign n568 = n541 & n567 ;
  assign n569 = n568 ^ n541 ;
  assign n570 = n538 & n569 ;
  assign n571 = n570 ^ n569 ;
  assign n537 = ~n386 & n536 ;
  assign n572 = n571 ^ n537 ;
  assign n648 = n647 ^ n572 ;
  assign n649 = n533 & n648 ;
  assign n650 = n649 ^ n648 ;
  assign n519 = n492 & n518 ;
  assign n520 = n519 ^ n492 ;
  assign n521 = n489 & n520 ;
  assign n522 = n521 ^ n520 ;
  assign n488 = n461 & ~n487 ;
  assign n523 = n522 ^ n488 ;
  assign n524 = n458 & n523 ;
  assign n525 = n524 ^ n523 ;
  assign n452 = ~n448 & n451 ;
  assign n453 = ~n422 & n452 ;
  assign n421 = n394 & ~n420 ;
  assign n454 = n453 ^ n421 ;
  assign n526 = n525 ^ n454 ;
  assign n651 = n650 ^ n526 ;
  assign n690 = n689 ^ n651 ;
  assign n949 = n461 & n690 ;
  assign n950 = n949 ^ n461 ;
  assign n946 = n487 & n690 ;
  assign n947 = n946 ^ n487 ;
  assign n948 = n947 ^ n487 ;
  assign n951 = n950 ^ n948 ;
  assign n705 = n401 ^ n152 ;
  assign n706 = n705 ^ n397 ;
  assign n707 = n706 ^ n405 ;
  assign n703 = n414 ^ n410 ;
  assign n704 = n703 ^ n418 ;
  assign n708 = n707 ^ n704 ;
  assign n710 = n708 ^ x24 ;
  assign n713 = n429 ^ n179 ;
  assign n714 = n713 ^ n425 ;
  assign n715 = n714 ^ n433 ;
  assign n711 = n442 ^ n438 ;
  assign n712 = n711 ^ n446 ;
  assign n716 = n715 ^ n712 ;
  assign n720 = n716 ^ x25 ;
  assign n721 = n710 & n720 ;
  assign n722 = n721 ^ n710 ;
  assign n723 = n722 ^ n720 ;
  assign n726 = n468 ^ n209 ;
  assign n727 = n726 ^ n464 ;
  assign n728 = n727 ^ n472 ;
  assign n724 = n481 ^ n477 ;
  assign n725 = n724 ^ n485 ;
  assign n729 = n728 ^ n725 ;
  assign n731 = n729 ^ x26 ;
  assign n734 = n499 ^ n236 ;
  assign n735 = n734 ^ n495 ;
  assign n736 = n735 ^ n503 ;
  assign n732 = n512 ^ n508 ;
  assign n733 = n732 ^ n516 ;
  assign n737 = n736 ^ n733 ;
  assign n746 = n737 ^ x27 ;
  assign n747 = n731 & n746 ;
  assign n748 = n747 ^ n731 ;
  assign n749 = n748 ^ n746 ;
  assign n750 = n723 & n749 ;
  assign n751 = n750 ^ n723 ;
  assign n752 = n751 ^ n749 ;
  assign n699 = n354 ^ n126 ;
  assign n700 = n699 ^ n340 ;
  assign n701 = n700 ^ n371 ;
  assign n697 = n380 ^ n376 ;
  assign n698 = n697 ^ n384 ;
  assign n702 = n701 ^ n698 ;
  assign n754 = n702 ^ x28 ;
  assign n757 = n548 ^ n270 ;
  assign n758 = n757 ^ n544 ;
  assign n759 = n758 ^ n552 ;
  assign n755 = n561 ^ n557 ;
  assign n756 = n755 ^ n565 ;
  assign n760 = n759 ^ n756 ;
  assign n766 = n760 ^ x29 ;
  assign n767 = n754 & n766 ;
  assign n768 = n767 ^ n754 ;
  assign n769 = n768 ^ n766 ;
  assign n815 = n599 ^ n595 ;
  assign n816 = n815 ^ n603 ;
  assign n811 = n586 ^ n300 ;
  assign n812 = n811 ^ n582 ;
  assign n813 = n812 ^ n590 ;
  assign n837 = n816 ^ n813 ;
  assign n838 = n837 ^ x30 ;
  assign n807 = n678 ^ x23 ;
  assign n808 = n807 ^ n664 ;
  assign n839 = n808 ^ x31 ;
  assign n840 = n838 & n839 ;
  assign n841 = n840 ^ n838 ;
  assign n842 = n841 ^ n839 ;
  assign n843 = n769 & n842 ;
  assign n844 = n843 ^ n769 ;
  assign n845 = n844 ^ n842 ;
  assign n846 = n752 & n845 ;
  assign n847 = n846 ^ n752 ;
  assign n848 = n847 ^ n845 ;
  assign n774 = ~n183 & n351 ;
  assign n775 = n774 ^ n344 ;
  assign n821 = x22 & ~x30 ;
  assign n825 = ~n775 & n821 ;
  assign n824 = n337 & n821 ;
  assign n826 = n825 ^ n824 ;
  assign n822 = ~n243 & n821 ;
  assign n823 = n368 & n822 ;
  assign n827 = n826 ^ n823 ;
  assign n828 = n827 ^ n821 ;
  assign n793 = x23 & x31 ;
  assign n801 = ~n183 & n793 ;
  assign n802 = n351 & n801 ;
  assign n800 = n344 & n793 ;
  assign n803 = n802 ^ n800 ;
  assign n797 = n337 & n793 ;
  assign n798 = n797 ^ n793 ;
  assign n799 = n798 ^ n793 ;
  assign n804 = n803 ^ n799 ;
  assign n794 = n243 & n793 ;
  assign n795 = n794 ^ n793 ;
  assign n796 = n368 & n795 ;
  assign n805 = n804 ^ n796 ;
  assign n779 = x31 & n327 ;
  assign n787 = ~n183 & n779 ;
  assign n788 = n351 & n787 ;
  assign n786 = n344 & n779 ;
  assign n789 = n788 ^ n786 ;
  assign n790 = n789 ^ n779 ;
  assign n783 = n337 & n779 ;
  assign n784 = n783 ^ n779 ;
  assign n785 = n784 ^ n779 ;
  assign n791 = n790 ^ n785 ;
  assign n780 = n243 & n779 ;
  assign n781 = n780 ^ n779 ;
  assign n782 = n368 & n781 ;
  assign n792 = n791 ^ n782 ;
  assign n806 = n805 ^ n792 ;
  assign n809 = n808 ^ n806 ;
  assign n817 = n809 & n816 ;
  assign n814 = n809 & n813 ;
  assign n818 = n817 ^ n814 ;
  assign n810 = x30 & n809 ;
  assign n819 = n818 ^ n810 ;
  assign n820 = n819 ^ n809 ;
  assign n829 = n828 ^ n820 ;
  assign n770 = ~x30 & n300 ;
  assign n776 = n770 & ~n775 ;
  assign n773 = n337 & n770 ;
  assign n777 = n776 ^ n773 ;
  assign n771 = ~n243 & n770 ;
  assign n772 = n368 & n771 ;
  assign n778 = n777 ^ n772 ;
  assign n830 = n829 ^ n778 ;
  assign n831 = n769 & n830 ;
  assign n832 = n831 ^ n830 ;
  assign n761 = x29 & n760 ;
  assign n762 = n761 ^ n760 ;
  assign n763 = n754 & n762 ;
  assign n764 = n763 ^ n762 ;
  assign n753 = ~x28 & n702 ;
  assign n765 = n764 ^ n753 ;
  assign n833 = n832 ^ n765 ;
  assign n834 = n752 & n833 ;
  assign n835 = n834 ^ n833 ;
  assign n738 = x27 & n737 ;
  assign n739 = n738 ^ n737 ;
  assign n740 = n731 & n739 ;
  assign n741 = n740 ^ n739 ;
  assign n730 = ~x26 & n729 ;
  assign n742 = n741 ^ n730 ;
  assign n743 = n723 & n742 ;
  assign n744 = n743 ^ n742 ;
  assign n717 = ~x25 & n716 ;
  assign n718 = ~n710 & n717 ;
  assign n709 = ~x24 & n708 ;
  assign n719 = n718 ^ n709 ;
  assign n745 = n744 ^ n719 ;
  assign n836 = n835 ^ n745 ;
  assign n849 = n848 ^ n836 ;
  assign n943 = x26 & n849 ;
  assign n944 = n943 ^ x26 ;
  assign n940 = n729 & n849 ;
  assign n941 = n940 ^ n729 ;
  assign n942 = n941 ^ n729 ;
  assign n945 = n944 ^ n942 ;
  assign n952 = n951 ^ n945 ;
  assign n956 = n492 & n690 ;
  assign n957 = n956 ^ n492 ;
  assign n953 = n518 & n690 ;
  assign n954 = n953 ^ n518 ;
  assign n955 = n954 ^ n518 ;
  assign n958 = n957 ^ n955 ;
  assign n962 = x27 & n849 ;
  assign n963 = n962 ^ x27 ;
  assign n959 = n737 & n849 ;
  assign n960 = n959 ^ n737 ;
  assign n961 = n960 ^ n737 ;
  assign n964 = n963 ^ n961 ;
  assign n994 = n958 & n964 ;
  assign n995 = n994 ^ n958 ;
  assign n996 = n952 & n995 ;
  assign n997 = n996 ^ n995 ;
  assign n993 = ~n945 & n951 ;
  assign n998 = n997 ^ n993 ;
  assign n920 = x24 & n849 ;
  assign n921 = n920 ^ x24 ;
  assign n917 = n708 & n849 ;
  assign n918 = n917 ^ n708 ;
  assign n919 = n918 ^ n708 ;
  assign n922 = n921 ^ n919 ;
  assign n914 = n394 & n690 ;
  assign n915 = n914 ^ n394 ;
  assign n911 = n420 & n690 ;
  assign n912 = n911 ^ n420 ;
  assign n913 = n912 ^ n420 ;
  assign n916 = n915 ^ n913 ;
  assign n923 = n922 ^ n916 ;
  assign n933 = x25 & n849 ;
  assign n934 = n933 ^ x25 ;
  assign n930 = n716 & n849 ;
  assign n931 = n930 ^ n716 ;
  assign n932 = n931 ^ n716 ;
  assign n935 = n934 ^ n932 ;
  assign n927 = n451 & n690 ;
  assign n928 = n927 ^ n451 ;
  assign n924 = n448 & n690 ;
  assign n925 = n924 ^ n448 ;
  assign n926 = n925 ^ n448 ;
  assign n929 = n928 ^ n926 ;
  assign n936 = n935 ^ n929 ;
  assign n937 = n923 & n936 ;
  assign n938 = n937 ^ n923 ;
  assign n939 = n938 ^ n936 ;
  assign n1081 = ~n939 & n945 ;
  assign n1082 = n998 & n1081 ;
  assign n989 = n929 & ~n935 ;
  assign n990 = ~n923 & n989 ;
  assign n988 = n916 & ~n922 ;
  assign n991 = n990 ^ n988 ;
  assign n1080 = n945 & n991 ;
  assign n1083 = n1082 ^ n1080 ;
  assign n1084 = n1083 ^ n945 ;
  assign n965 = n964 ^ n958 ;
  assign n966 = n952 & n965 ;
  assign n967 = n966 ^ n952 ;
  assign n968 = n967 ^ n965 ;
  assign n969 = n939 & n968 ;
  assign n970 = n969 ^ n939 ;
  assign n971 = n970 ^ n968 ;
  assign n853 = x28 & n849 ;
  assign n854 = n853 ^ x28 ;
  assign n850 = n702 & n849 ;
  assign n851 = n850 ^ n702 ;
  assign n852 = n851 ^ n702 ;
  assign n855 = n854 ^ n852 ;
  assign n694 = n536 & n690 ;
  assign n695 = n694 ^ n536 ;
  assign n691 = n386 & n690 ;
  assign n692 = n691 ^ n386 ;
  assign n693 = n692 ^ n386 ;
  assign n696 = n695 ^ n693 ;
  assign n857 = n855 ^ n696 ;
  assign n867 = x29 & n849 ;
  assign n868 = n867 ^ x29 ;
  assign n864 = n760 & n849 ;
  assign n865 = n864 ^ n760 ;
  assign n866 = n865 ^ n760 ;
  assign n869 = n868 ^ n866 ;
  assign n861 = n541 & n690 ;
  assign n862 = n861 ^ n541 ;
  assign n858 = n567 & n690 ;
  assign n859 = n858 ^ n567 ;
  assign n860 = n859 ^ n567 ;
  assign n863 = n862 ^ n860 ;
  assign n873 = n869 ^ n863 ;
  assign n874 = n857 & n873 ;
  assign n875 = n874 ^ n857 ;
  assign n876 = n875 ^ n873 ;
  assign n886 = x30 & n849 ;
  assign n887 = n886 ^ x30 ;
  assign n883 = n837 & n849 ;
  assign n884 = n883 ^ n837 ;
  assign n885 = n884 ^ n837 ;
  assign n888 = n887 ^ n885 ;
  assign n880 = n579 & n690 ;
  assign n881 = n880 ^ n579 ;
  assign n877 = n605 & n690 ;
  assign n878 = n877 ^ n605 ;
  assign n879 = n878 ^ n605 ;
  assign n882 = n881 ^ n879 ;
  assign n890 = n888 ^ n882 ;
  assign n900 = n613 & n690 ;
  assign n901 = n900 ^ n613 ;
  assign n897 = n679 & n690 ;
  assign n898 = n897 ^ n679 ;
  assign n899 = n898 ^ n679 ;
  assign n902 = n901 ^ n899 ;
  assign n894 = x31 & n849 ;
  assign n895 = n894 ^ x31 ;
  assign n891 = n808 & n849 ;
  assign n892 = n891 ^ n808 ;
  assign n893 = n892 ^ n808 ;
  assign n896 = n895 ^ n893 ;
  assign n975 = n902 ^ n896 ;
  assign n976 = n890 & n975 ;
  assign n977 = n976 ^ n890 ;
  assign n978 = n977 ^ n975 ;
  assign n979 = n876 & n978 ;
  assign n980 = n979 ^ n876 ;
  assign n981 = n980 ^ n978 ;
  assign n982 = n971 & n981 ;
  assign n983 = n982 ^ n971 ;
  assign n984 = n983 ^ n981 ;
  assign n1077 = n945 & n984 ;
  assign n1078 = n1077 ^ n945 ;
  assign n1079 = n1078 ^ n945 ;
  assign n1085 = n1084 ^ n1079 ;
  assign n903 = n896 & n902 ;
  assign n904 = n903 ^ n902 ;
  assign n905 = n890 & n904 ;
  assign n906 = n905 ^ n904 ;
  assign n889 = n882 & ~n888 ;
  assign n907 = n906 ^ n889 ;
  assign n908 = n876 & n907 ;
  assign n909 = n908 ^ n907 ;
  assign n870 = n863 & ~n869 ;
  assign n871 = ~n857 & n870 ;
  assign n856 = n696 & ~n855 ;
  assign n872 = n871 ^ n856 ;
  assign n910 = n909 ^ n872 ;
  assign n1074 = n945 & n971 ;
  assign n1075 = n1074 ^ n945 ;
  assign n1076 = n910 & n1075 ;
  assign n1086 = n1085 ^ n1076 ;
  assign n1511 = n1086 ^ n945 ;
  assign n1067 = ~n939 & n951 ;
  assign n1068 = n998 & n1067 ;
  assign n1066 = n951 & n991 ;
  assign n1069 = n1068 ^ n1066 ;
  assign n1070 = n1069 ^ n951 ;
  assign n1063 = n951 & n984 ;
  assign n1064 = n1063 ^ n951 ;
  assign n1065 = n1064 ^ n951 ;
  assign n1071 = n1070 ^ n1065 ;
  assign n1060 = n951 & n971 ;
  assign n1061 = n1060 ^ n951 ;
  assign n1062 = n910 & n1061 ;
  assign n1072 = n1071 ^ n1062 ;
  assign n1512 = n1511 ^ n1072 ;
  assign n1329 = n921 ^ x24 ;
  assign n1330 = n1329 ^ n918 ;
  assign n1332 = n1330 ^ x32 ;
  assign n1333 = n934 ^ x25 ;
  assign n1334 = n1333 ^ n931 ;
  assign n1338 = n1334 ^ x33 ;
  assign n1339 = n1332 & n1338 ;
  assign n1340 = n1339 ^ n1332 ;
  assign n1341 = n1340 ^ n1338 ;
  assign n1342 = n944 ^ x26 ;
  assign n1343 = n1342 ^ n941 ;
  assign n1345 = n1343 ^ x34 ;
  assign n1351 = n963 ^ x27 ;
  assign n1352 = n1351 ^ n960 ;
  assign n1359 = n1352 ^ x35 ;
  assign n1360 = n1345 & n1359 ;
  assign n1361 = n1360 ^ n1345 ;
  assign n1362 = n1361 ^ n1359 ;
  assign n1363 = n1341 & n1362 ;
  assign n1364 = n1363 ^ n1341 ;
  assign n1365 = n1364 ^ n1362 ;
  assign n1327 = n854 ^ x28 ;
  assign n1328 = n1327 ^ n851 ;
  assign n1367 = n1328 ^ x36 ;
  assign n1373 = n868 ^ x29 ;
  assign n1374 = n1373 ^ n865 ;
  assign n1379 = n1374 ^ x37 ;
  assign n1380 = n1367 & n1379 ;
  assign n1381 = n1380 ^ n1367 ;
  assign n1382 = n1381 ^ n1379 ;
  assign n1404 = n887 ^ x30 ;
  assign n1419 = n1404 ^ n884 ;
  assign n1420 = n1419 ^ x38 ;
  assign n1400 = n895 ^ x31 ;
  assign n1401 = n1400 ^ n892 ;
  assign n1421 = n1401 ^ x39 ;
  assign n1422 = n1420 & n1421 ;
  assign n1423 = n1422 ^ n1420 ;
  assign n1424 = n1423 ^ n1421 ;
  assign n1425 = n1382 & n1424 ;
  assign n1426 = n1425 ^ n1382 ;
  assign n1427 = n1426 ^ n1424 ;
  assign n1428 = n1365 & n1427 ;
  assign n1429 = n1428 ^ n1365 ;
  assign n1430 = n1429 ^ n1427 ;
  assign n1409 = x30 & ~x38 ;
  assign n1410 = n849 & n1409 ;
  assign n1395 = x31 & x39 ;
  assign n1396 = n849 & n1395 ;
  assign n1397 = n1396 ^ n1395 ;
  assign n1398 = n1397 ^ n1395 ;
  assign n1392 = x39 & n808 ;
  assign n1393 = n849 & n1392 ;
  assign n1394 = n1393 ^ n1392 ;
  assign n1399 = n1398 ^ n1394 ;
  assign n1402 = n1401 ^ n1399 ;
  assign n1405 = n1402 & n1404 ;
  assign n1403 = n884 & n1402 ;
  assign n1406 = n1405 ^ n1403 ;
  assign n1388 = x31 & x38 ;
  assign n1389 = ~x39 & n1388 ;
  assign n1390 = n849 & n1389 ;
  assign n1385 = x38 & ~x39 ;
  assign n1386 = n808 & n1385 ;
  assign n1387 = ~n849 & n1386 ;
  assign n1391 = n1390 ^ n1387 ;
  assign n1407 = n1406 ^ n1391 ;
  assign n1408 = n1407 ^ n1402 ;
  assign n1411 = n1410 ^ n1408 ;
  assign n1383 = ~x38 & n837 ;
  assign n1384 = ~n849 & n1383 ;
  assign n1412 = n1411 ^ n1384 ;
  assign n1413 = n1382 & n1412 ;
  assign n1414 = n1413 ^ n1412 ;
  assign n1370 = x29 & x37 ;
  assign n1371 = n849 & n1370 ;
  assign n1368 = x37 & n760 ;
  assign n1369 = ~n849 & n1368 ;
  assign n1372 = n1371 ^ n1369 ;
  assign n1375 = n1374 ^ n1372 ;
  assign n1376 = n1367 & n1375 ;
  assign n1377 = n1376 ^ n1375 ;
  assign n1366 = ~x36 & n1328 ;
  assign n1378 = n1377 ^ n1366 ;
  assign n1415 = n1414 ^ n1378 ;
  assign n1416 = n1365 & n1415 ;
  assign n1417 = n1416 ^ n1415 ;
  assign n1348 = x27 & x35 ;
  assign n1349 = n849 & n1348 ;
  assign n1346 = x35 & n737 ;
  assign n1347 = ~n849 & n1346 ;
  assign n1350 = n1349 ^ n1347 ;
  assign n1353 = n1352 ^ n1350 ;
  assign n1354 = n1345 & n1353 ;
  assign n1355 = n1354 ^ n1353 ;
  assign n1344 = ~x34 & n1343 ;
  assign n1356 = n1355 ^ n1344 ;
  assign n1357 = ~n1341 & n1356 ;
  assign n1335 = ~x33 & n1334 ;
  assign n1336 = ~n1332 & n1335 ;
  assign n1331 = ~x32 & n1330 ;
  assign n1337 = n1336 ^ n1331 ;
  assign n1358 = n1357 ^ n1337 ;
  assign n1418 = n1417 ^ n1358 ;
  assign n1431 = n1430 ^ n1418 ;
  assign n1508 = x34 & n1431 ;
  assign n1509 = n1508 ^ x34 ;
  assign n1505 = n1343 & n1431 ;
  assign n1506 = n1505 ^ n1343 ;
  assign n1507 = n1506 ^ n1343 ;
  assign n1510 = n1509 ^ n1507 ;
  assign n1513 = n1512 ^ n1510 ;
  assign n1112 = ~n939 & n964 ;
  assign n1113 = n998 & n1112 ;
  assign n1111 = n964 & n991 ;
  assign n1114 = n1113 ^ n1111 ;
  assign n1115 = n1114 ^ n964 ;
  assign n1108 = n964 & n984 ;
  assign n1109 = n1108 ^ n964 ;
  assign n1110 = n1109 ^ n964 ;
  assign n1116 = n1115 ^ n1110 ;
  assign n1105 = n964 & n971 ;
  assign n1106 = n1105 ^ n964 ;
  assign n1107 = n910 & n1106 ;
  assign n1117 = n1116 ^ n1107 ;
  assign n1514 = n1117 ^ n964 ;
  assign n1098 = ~n939 & n958 ;
  assign n1099 = n998 & n1098 ;
  assign n1097 = n958 & n991 ;
  assign n1100 = n1099 ^ n1097 ;
  assign n1101 = n1100 ^ n958 ;
  assign n1094 = n958 & n984 ;
  assign n1095 = n1094 ^ n958 ;
  assign n1096 = n1095 ^ n958 ;
  assign n1102 = n1101 ^ n1096 ;
  assign n1091 = n958 & n971 ;
  assign n1092 = n1091 ^ n958 ;
  assign n1093 = n910 & n1092 ;
  assign n1103 = n1102 ^ n1093 ;
  assign n1515 = n1514 ^ n1103 ;
  assign n1519 = x35 & n1431 ;
  assign n1520 = n1519 ^ x35 ;
  assign n1516 = n1352 & n1431 ;
  assign n1517 = n1516 ^ n1352 ;
  assign n1518 = n1517 ^ n1352 ;
  assign n1521 = n1520 ^ n1518 ;
  assign n1551 = n1515 & n1521 ;
  assign n1552 = n1551 ^ n1515 ;
  assign n1553 = n1513 & n1552 ;
  assign n1554 = n1553 ^ n1552 ;
  assign n1550 = ~n1510 & n1512 ;
  assign n1555 = n1554 ^ n1550 ;
  assign n1489 = x32 & n1431 ;
  assign n1490 = n1489 ^ x32 ;
  assign n1486 = n1330 & n1431 ;
  assign n1487 = n1486 ^ n1330 ;
  assign n1488 = n1487 ^ n1330 ;
  assign n1491 = n1490 ^ n1488 ;
  assign n1013 = n922 & ~n939 ;
  assign n1014 = n998 & n1013 ;
  assign n1012 = n922 & n991 ;
  assign n1015 = n1014 ^ n1012 ;
  assign n1016 = n1015 ^ n922 ;
  assign n1009 = n922 & n984 ;
  assign n1010 = n1009 ^ n922 ;
  assign n1011 = n1010 ^ n922 ;
  assign n1017 = n1016 ^ n1011 ;
  assign n1006 = n922 & n971 ;
  assign n1007 = n1006 ^ n922 ;
  assign n1008 = n910 & n1007 ;
  assign n1018 = n1017 ^ n1008 ;
  assign n1484 = n1018 ^ n922 ;
  assign n999 = n916 & ~n939 ;
  assign n1000 = n998 & n999 ;
  assign n992 = n916 & n991 ;
  assign n1001 = n1000 ^ n992 ;
  assign n1002 = n1001 ^ n916 ;
  assign n985 = n916 & n984 ;
  assign n986 = n985 ^ n916 ;
  assign n987 = n986 ^ n916 ;
  assign n1003 = n1002 ^ n987 ;
  assign n972 = n916 & n971 ;
  assign n973 = n972 ^ n916 ;
  assign n974 = n910 & n973 ;
  assign n1004 = n1003 ^ n974 ;
  assign n1485 = n1484 ^ n1004 ;
  assign n1492 = n1491 ^ n1485 ;
  assign n1498 = x33 & n1431 ;
  assign n1499 = n1498 ^ x33 ;
  assign n1495 = n1334 & n1431 ;
  assign n1496 = n1495 ^ n1334 ;
  assign n1497 = n1496 ^ n1334 ;
  assign n1500 = n1499 ^ n1497 ;
  assign n1044 = n935 & ~n939 ;
  assign n1045 = n998 & n1044 ;
  assign n1043 = n935 & n991 ;
  assign n1046 = n1045 ^ n1043 ;
  assign n1047 = n1046 ^ n935 ;
  assign n1040 = n935 & n984 ;
  assign n1041 = n1040 ^ n935 ;
  assign n1042 = n1041 ^ n935 ;
  assign n1048 = n1047 ^ n1042 ;
  assign n1037 = n935 & n971 ;
  assign n1038 = n1037 ^ n935 ;
  assign n1039 = n910 & n1038 ;
  assign n1049 = n1048 ^ n1039 ;
  assign n1493 = n1049 ^ n935 ;
  assign n1030 = n929 & ~n939 ;
  assign n1031 = n998 & n1030 ;
  assign n1029 = n929 & n991 ;
  assign n1032 = n1031 ^ n1029 ;
  assign n1033 = n1032 ^ n929 ;
  assign n1026 = n929 & n984 ;
  assign n1027 = n1026 ^ n929 ;
  assign n1028 = n1027 ^ n929 ;
  assign n1034 = n1033 ^ n1028 ;
  assign n1023 = n929 & n971 ;
  assign n1024 = n1023 ^ n929 ;
  assign n1025 = n910 & n1024 ;
  assign n1035 = n1034 ^ n1025 ;
  assign n1494 = n1493 ^ n1035 ;
  assign n1501 = n1500 ^ n1494 ;
  assign n1502 = n1492 & n1501 ;
  assign n1503 = n1502 ^ n1492 ;
  assign n1504 = n1503 ^ n1501 ;
  assign n1792 = ~n1504 & n1510 ;
  assign n1793 = n1555 & n1792 ;
  assign n1546 = n1494 & ~n1500 ;
  assign n1547 = ~n1492 & n1546 ;
  assign n1545 = n1485 & ~n1491 ;
  assign n1548 = n1547 ^ n1545 ;
  assign n1791 = n1510 & n1548 ;
  assign n1794 = n1793 ^ n1791 ;
  assign n1795 = n1794 ^ n1510 ;
  assign n1522 = n1521 ^ n1515 ;
  assign n1523 = n1513 & n1522 ;
  assign n1524 = n1523 ^ n1513 ;
  assign n1525 = n1524 ^ n1522 ;
  assign n1526 = n1504 & n1525 ;
  assign n1527 = n1526 ^ n1504 ;
  assign n1528 = n1527 ^ n1525 ;
  assign n1435 = x36 & n1431 ;
  assign n1436 = n1435 ^ x36 ;
  assign n1432 = n1328 & n1431 ;
  assign n1433 = n1432 ^ n1328 ;
  assign n1434 = n1433 ^ n1328 ;
  assign n1437 = n1436 ^ n1434 ;
  assign n1156 = n855 & ~n939 ;
  assign n1157 = n998 & n1156 ;
  assign n1155 = n855 & n991 ;
  assign n1158 = n1157 ^ n1155 ;
  assign n1159 = n1158 ^ n855 ;
  assign n1152 = n855 & n984 ;
  assign n1153 = n1152 ^ n855 ;
  assign n1154 = n1153 ^ n855 ;
  assign n1160 = n1159 ^ n1154 ;
  assign n1149 = n855 & n971 ;
  assign n1150 = n1149 ^ n855 ;
  assign n1151 = n910 & n1150 ;
  assign n1161 = n1160 ^ n1151 ;
  assign n1325 = n1161 ^ n855 ;
  assign n1142 = n696 & ~n939 ;
  assign n1143 = n998 & n1142 ;
  assign n1141 = n696 & n991 ;
  assign n1144 = n1143 ^ n1141 ;
  assign n1145 = n1144 ^ n696 ;
  assign n1138 = n696 & n984 ;
  assign n1139 = n1138 ^ n696 ;
  assign n1140 = n1139 ^ n696 ;
  assign n1146 = n1145 ^ n1140 ;
  assign n1135 = n696 & n971 ;
  assign n1136 = n1135 ^ n696 ;
  assign n1137 = n910 & n1136 ;
  assign n1147 = n1146 ^ n1137 ;
  assign n1326 = n1325 ^ n1147 ;
  assign n1439 = n1437 ^ n1326 ;
  assign n1445 = x37 & n1431 ;
  assign n1446 = n1445 ^ x37 ;
  assign n1442 = n1374 & n1431 ;
  assign n1443 = n1442 ^ n1374 ;
  assign n1444 = n1443 ^ n1374 ;
  assign n1447 = n1446 ^ n1444 ;
  assign n1187 = n869 & ~n939 ;
  assign n1188 = n998 & n1187 ;
  assign n1186 = n869 & n991 ;
  assign n1189 = n1188 ^ n1186 ;
  assign n1190 = n1189 ^ n869 ;
  assign n1183 = n869 & n984 ;
  assign n1184 = n1183 ^ n869 ;
  assign n1185 = n1184 ^ n869 ;
  assign n1191 = n1190 ^ n1185 ;
  assign n1180 = n869 & n971 ;
  assign n1181 = n1180 ^ n869 ;
  assign n1182 = n910 & n1181 ;
  assign n1192 = n1191 ^ n1182 ;
  assign n1440 = n1192 ^ n869 ;
  assign n1173 = n863 & ~n939 ;
  assign n1174 = n998 & n1173 ;
  assign n1172 = n863 & n991 ;
  assign n1175 = n1174 ^ n1172 ;
  assign n1176 = n1175 ^ n863 ;
  assign n1169 = n863 & n984 ;
  assign n1170 = n1169 ^ n863 ;
  assign n1171 = n1170 ^ n863 ;
  assign n1177 = n1176 ^ n1171 ;
  assign n1166 = n863 & n971 ;
  assign n1167 = n1166 ^ n863 ;
  assign n1168 = n910 & n1167 ;
  assign n1178 = n1177 ^ n1168 ;
  assign n1441 = n1440 ^ n1178 ;
  assign n1453 = n1447 ^ n1441 ;
  assign n1454 = n1439 & n1453 ;
  assign n1455 = n1454 ^ n1439 ;
  assign n1456 = n1455 ^ n1453 ;
  assign n1462 = x38 & n1431 ;
  assign n1463 = n1462 ^ x38 ;
  assign n1459 = n1419 & n1431 ;
  assign n1460 = n1459 ^ n1419 ;
  assign n1461 = n1460 ^ n1419 ;
  assign n1464 = n1463 ^ n1461 ;
  assign n1225 = n888 & ~n939 ;
  assign n1226 = n998 & n1225 ;
  assign n1224 = n888 & n991 ;
  assign n1227 = n1226 ^ n1224 ;
  assign n1228 = n1227 ^ n888 ;
  assign n1221 = n888 & n984 ;
  assign n1222 = n1221 ^ n888 ;
  assign n1223 = n1222 ^ n888 ;
  assign n1229 = n1228 ^ n1223 ;
  assign n1218 = n888 & n971 ;
  assign n1219 = n1218 ^ n888 ;
  assign n1220 = n910 & n1219 ;
  assign n1230 = n1229 ^ n1220 ;
  assign n1457 = n1230 ^ n888 ;
  assign n1211 = n882 & ~n939 ;
  assign n1212 = n998 & n1211 ;
  assign n1210 = n882 & n991 ;
  assign n1213 = n1212 ^ n1210 ;
  assign n1214 = n1213 ^ n882 ;
  assign n1207 = n882 & n984 ;
  assign n1208 = n1207 ^ n882 ;
  assign n1209 = n1208 ^ n882 ;
  assign n1215 = n1214 ^ n1209 ;
  assign n1204 = n882 & n971 ;
  assign n1205 = n1204 ^ n882 ;
  assign n1206 = n910 & n1205 ;
  assign n1216 = n1215 ^ n1206 ;
  assign n1458 = n1457 ^ n1216 ;
  assign n1467 = n1464 ^ n1458 ;
  assign n1297 = n896 & ~n939 ;
  assign n1298 = n998 & n1297 ;
  assign n1296 = n896 & n991 ;
  assign n1299 = n1298 ^ n1296 ;
  assign n1300 = n1299 ^ n896 ;
  assign n1293 = n896 & n984 ;
  assign n1294 = n1293 ^ n896 ;
  assign n1295 = n1294 ^ n896 ;
  assign n1301 = n1300 ^ n1295 ;
  assign n1290 = n896 & n971 ;
  assign n1291 = n1290 ^ n896 ;
  assign n1292 = n910 & n1291 ;
  assign n1302 = n1301 ^ n1292 ;
  assign n1474 = n1302 ^ n896 ;
  assign n1283 = n902 & ~n939 ;
  assign n1284 = n998 & n1283 ;
  assign n1282 = n902 & n991 ;
  assign n1285 = n1284 ^ n1282 ;
  assign n1286 = n1285 ^ n902 ;
  assign n1279 = n902 & n984 ;
  assign n1280 = n1279 ^ n902 ;
  assign n1281 = n1280 ^ n902 ;
  assign n1287 = n1286 ^ n1281 ;
  assign n1276 = n902 & n971 ;
  assign n1277 = n1276 ^ n902 ;
  assign n1278 = n910 & n1277 ;
  assign n1288 = n1287 ^ n1278 ;
  assign n1475 = n1474 ^ n1288 ;
  assign n1471 = x39 & n1431 ;
  assign n1472 = n1471 ^ x39 ;
  assign n1468 = n1401 & n1431 ;
  assign n1469 = n1468 ^ n1401 ;
  assign n1470 = n1469 ^ n1401 ;
  assign n1473 = n1472 ^ n1470 ;
  assign n1532 = n1475 ^ n1473 ;
  assign n1533 = n1467 & n1532 ;
  assign n1534 = n1533 ^ n1467 ;
  assign n1535 = n1534 ^ n1532 ;
  assign n1536 = n1456 & n1535 ;
  assign n1537 = n1536 ^ n1456 ;
  assign n1538 = n1537 ^ n1535 ;
  assign n1539 = n1528 & n1538 ;
  assign n1540 = n1539 ^ n1528 ;
  assign n1541 = n1540 ^ n1538 ;
  assign n1788 = n1510 & n1541 ;
  assign n1789 = n1788 ^ n1510 ;
  assign n1790 = n1789 ^ n1510 ;
  assign n1796 = n1795 ^ n1790 ;
  assign n1476 = n1473 & n1475 ;
  assign n1477 = n1476 ^ n1475 ;
  assign n1478 = n1467 & n1477 ;
  assign n1479 = n1478 ^ n1477 ;
  assign n1465 = n1458 & n1464 ;
  assign n1466 = n1465 ^ n1458 ;
  assign n1480 = n1479 ^ n1466 ;
  assign n1481 = n1456 & n1480 ;
  assign n1482 = n1481 ^ n1480 ;
  assign n1448 = n1441 & n1447 ;
  assign n1449 = n1448 ^ n1441 ;
  assign n1450 = n1439 & n1449 ;
  assign n1451 = n1450 ^ n1449 ;
  assign n1438 = n1326 & ~n1437 ;
  assign n1452 = n1451 ^ n1438 ;
  assign n1483 = n1482 ^ n1452 ;
  assign n1785 = n1510 & n1528 ;
  assign n1786 = n1785 ^ n1510 ;
  assign n1787 = n1483 & n1786 ;
  assign n1797 = n1796 ^ n1787 ;
  assign n2333 = n1797 ^ n1510 ;
  assign n1778 = ~n1504 & n1512 ;
  assign n1779 = n1555 & n1778 ;
  assign n1777 = n1512 & n1548 ;
  assign n1780 = n1779 ^ n1777 ;
  assign n1781 = n1780 ^ n1512 ;
  assign n1774 = n1512 & n1541 ;
  assign n1775 = n1774 ^ n1512 ;
  assign n1776 = n1775 ^ n1512 ;
  assign n1782 = n1781 ^ n1776 ;
  assign n1771 = n1512 & n1528 ;
  assign n1772 = n1771 ^ n1512 ;
  assign n1773 = n1483 & n1772 ;
  assign n1783 = n1782 ^ n1773 ;
  assign n2334 = n2333 ^ n1783 ;
  assign n2165 = n1490 ^ x32 ;
  assign n2166 = n2165 ^ n1487 ;
  assign n2168 = n2166 ^ x40 ;
  assign n2169 = n1499 ^ x33 ;
  assign n2170 = n2169 ^ n1496 ;
  assign n2174 = n2170 ^ x41 ;
  assign n2175 = n2168 & n2174 ;
  assign n2176 = n2175 ^ n2168 ;
  assign n2177 = n2176 ^ n2174 ;
  assign n2178 = n1509 ^ x34 ;
  assign n2179 = n2178 ^ n1506 ;
  assign n2181 = n2179 ^ x42 ;
  assign n2187 = n1520 ^ x35 ;
  assign n2188 = n2187 ^ n1517 ;
  assign n2195 = n2188 ^ x43 ;
  assign n2196 = n2181 & n2195 ;
  assign n2197 = n2196 ^ n2181 ;
  assign n2198 = n2197 ^ n2195 ;
  assign n2199 = n2177 & n2198 ;
  assign n2200 = n2199 ^ n2177 ;
  assign n2201 = n2200 ^ n2198 ;
  assign n2163 = n1436 ^ x36 ;
  assign n2164 = n2163 ^ n1433 ;
  assign n2203 = n2164 ^ x44 ;
  assign n2209 = n1446 ^ x37 ;
  assign n2210 = n2209 ^ n1443 ;
  assign n2215 = n2210 ^ x45 ;
  assign n2216 = n2203 & n2215 ;
  assign n2217 = n2216 ^ n2203 ;
  assign n2218 = n2217 ^ n2215 ;
  assign n2240 = n1463 ^ x38 ;
  assign n2255 = n2240 ^ n1460 ;
  assign n2256 = n2255 ^ x46 ;
  assign n2236 = n1472 ^ x39 ;
  assign n2237 = n2236 ^ n1469 ;
  assign n2257 = n2237 ^ x47 ;
  assign n2258 = n2256 & n2257 ;
  assign n2259 = n2258 ^ n2256 ;
  assign n2260 = n2259 ^ n2257 ;
  assign n2261 = n2218 & n2260 ;
  assign n2262 = n2261 ^ n2218 ;
  assign n2263 = n2262 ^ n2260 ;
  assign n2264 = n2201 & n2263 ;
  assign n2265 = n2264 ^ n2201 ;
  assign n2266 = n2265 ^ n2263 ;
  assign n2245 = x38 & ~x46 ;
  assign n2246 = n1431 & n2245 ;
  assign n2231 = x39 & x47 ;
  assign n2232 = n1431 & n2231 ;
  assign n2233 = n2232 ^ n2231 ;
  assign n2234 = n2233 ^ n2231 ;
  assign n2228 = x47 & n1401 ;
  assign n2229 = n1431 & n2228 ;
  assign n2230 = n2229 ^ n2228 ;
  assign n2235 = n2234 ^ n2230 ;
  assign n2238 = n2237 ^ n2235 ;
  assign n2241 = n2238 & n2240 ;
  assign n2239 = n1460 & n2238 ;
  assign n2242 = n2241 ^ n2239 ;
  assign n2224 = x39 & x46 ;
  assign n2225 = ~x47 & n2224 ;
  assign n2226 = n1431 & n2225 ;
  assign n2221 = x46 & ~x47 ;
  assign n2222 = n1401 & n2221 ;
  assign n2223 = ~n1431 & n2222 ;
  assign n2227 = n2226 ^ n2223 ;
  assign n2243 = n2242 ^ n2227 ;
  assign n2244 = n2243 ^ n2238 ;
  assign n2247 = n2246 ^ n2244 ;
  assign n2219 = ~x46 & n1419 ;
  assign n2220 = ~n1431 & n2219 ;
  assign n2248 = n2247 ^ n2220 ;
  assign n2249 = n2218 & n2248 ;
  assign n2250 = n2249 ^ n2248 ;
  assign n2206 = x37 & x45 ;
  assign n2207 = n1431 & n2206 ;
  assign n2204 = x45 & n1374 ;
  assign n2205 = ~n1431 & n2204 ;
  assign n2208 = n2207 ^ n2205 ;
  assign n2211 = n2210 ^ n2208 ;
  assign n2212 = n2203 & n2211 ;
  assign n2213 = n2212 ^ n2211 ;
  assign n2202 = ~x44 & n2164 ;
  assign n2214 = n2213 ^ n2202 ;
  assign n2251 = n2250 ^ n2214 ;
  assign n2252 = n2201 & n2251 ;
  assign n2253 = n2252 ^ n2251 ;
  assign n2184 = x35 & x43 ;
  assign n2185 = n1431 & n2184 ;
  assign n2182 = x43 & n1352 ;
  assign n2183 = ~n1431 & n2182 ;
  assign n2186 = n2185 ^ n2183 ;
  assign n2189 = n2188 ^ n2186 ;
  assign n2190 = n2181 & n2189 ;
  assign n2191 = n2190 ^ n2189 ;
  assign n2180 = ~x42 & n2179 ;
  assign n2192 = n2191 ^ n2180 ;
  assign n2193 = ~n2177 & n2192 ;
  assign n2171 = ~x41 & n2170 ;
  assign n2172 = ~n2168 & n2171 ;
  assign n2167 = ~x40 & n2166 ;
  assign n2173 = n2172 ^ n2167 ;
  assign n2194 = n2193 ^ n2173 ;
  assign n2254 = n2253 ^ n2194 ;
  assign n2267 = n2266 ^ n2254 ;
  assign n2331 = x42 & ~n2267 ;
  assign n2329 = n2179 & ~n2267 ;
  assign n2330 = n2329 ^ n2179 ;
  assign n2332 = n2331 ^ n2330 ;
  assign n2335 = n2334 ^ n2332 ;
  assign n1833 = ~n1504 & n1521 ;
  assign n1834 = n1555 & n1833 ;
  assign n1832 = n1521 & n1548 ;
  assign n1835 = n1834 ^ n1832 ;
  assign n1836 = n1835 ^ n1521 ;
  assign n1829 = n1521 & n1541 ;
  assign n1830 = n1829 ^ n1521 ;
  assign n1831 = n1830 ^ n1521 ;
  assign n1837 = n1836 ^ n1831 ;
  assign n1826 = n1521 & n1528 ;
  assign n1827 = n1826 ^ n1521 ;
  assign n1828 = n1483 & n1827 ;
  assign n1838 = n1837 ^ n1828 ;
  assign n2336 = n1838 ^ n1521 ;
  assign n1819 = ~n1504 & n1515 ;
  assign n1820 = n1555 & n1819 ;
  assign n1818 = n1515 & n1548 ;
  assign n1821 = n1820 ^ n1818 ;
  assign n1822 = n1821 ^ n1515 ;
  assign n1815 = n1515 & n1541 ;
  assign n1816 = n1815 ^ n1515 ;
  assign n1817 = n1816 ^ n1515 ;
  assign n1823 = n1822 ^ n1817 ;
  assign n1812 = n1515 & n1528 ;
  assign n1813 = n1812 ^ n1515 ;
  assign n1814 = n1483 & n1813 ;
  assign n1824 = n1823 ^ n1814 ;
  assign n2337 = n2336 ^ n1824 ;
  assign n2340 = x43 & ~n2267 ;
  assign n2338 = n2188 & ~n2267 ;
  assign n2339 = n2338 ^ n2188 ;
  assign n2341 = n2340 ^ n2339 ;
  assign n2370 = n2337 & n2341 ;
  assign n2371 = n2370 ^ n2337 ;
  assign n2372 = n2335 & n2371 ;
  assign n2373 = n2372 ^ n2371 ;
  assign n2369 = ~n2332 & n2334 ;
  assign n2374 = n2373 ^ n2369 ;
  assign n2316 = x40 & ~n2267 ;
  assign n2314 = n2166 & ~n2267 ;
  assign n2315 = n2314 ^ n2166 ;
  assign n2317 = n2316 ^ n2315 ;
  assign n1725 = n1491 & ~n1504 ;
  assign n1726 = n1555 & n1725 ;
  assign n1724 = n1491 & n1548 ;
  assign n1727 = n1726 ^ n1724 ;
  assign n1728 = n1727 ^ n1491 ;
  assign n1721 = n1491 & n1541 ;
  assign n1722 = n1721 ^ n1491 ;
  assign n1723 = n1722 ^ n1491 ;
  assign n1729 = n1728 ^ n1723 ;
  assign n1718 = n1491 & n1528 ;
  assign n1719 = n1718 ^ n1491 ;
  assign n1720 = n1483 & n1719 ;
  assign n1730 = n1729 ^ n1720 ;
  assign n2312 = n1730 ^ n1491 ;
  assign n1711 = n1485 & ~n1504 ;
  assign n1712 = n1555 & n1711 ;
  assign n1710 = n1485 & n1548 ;
  assign n1713 = n1712 ^ n1710 ;
  assign n1714 = n1713 ^ n1485 ;
  assign n1707 = n1485 & n1541 ;
  assign n1708 = n1707 ^ n1485 ;
  assign n1709 = n1708 ^ n1485 ;
  assign n1715 = n1714 ^ n1709 ;
  assign n1704 = n1485 & n1528 ;
  assign n1705 = n1704 ^ n1485 ;
  assign n1706 = n1483 & n1705 ;
  assign n1716 = n1715 ^ n1706 ;
  assign n2313 = n2312 ^ n1716 ;
  assign n2318 = n2317 ^ n2313 ;
  assign n1760 = n1500 & ~n1504 ;
  assign n1761 = n1555 & n1760 ;
  assign n1759 = n1500 & n1548 ;
  assign n1762 = n1761 ^ n1759 ;
  assign n1763 = n1762 ^ n1500 ;
  assign n1756 = n1500 & n1541 ;
  assign n1757 = n1756 ^ n1500 ;
  assign n1758 = n1757 ^ n1500 ;
  assign n1764 = n1763 ^ n1758 ;
  assign n1753 = n1500 & n1528 ;
  assign n1754 = n1753 ^ n1500 ;
  assign n1755 = n1483 & n1754 ;
  assign n1765 = n1764 ^ n1755 ;
  assign n2323 = n1765 ^ n1500 ;
  assign n1746 = n1494 & ~n1504 ;
  assign n1747 = n1555 & n1746 ;
  assign n1745 = n1494 & n1548 ;
  assign n1748 = n1747 ^ n1745 ;
  assign n1749 = n1748 ^ n1494 ;
  assign n1742 = n1494 & n1541 ;
  assign n1743 = n1742 ^ n1494 ;
  assign n1744 = n1743 ^ n1494 ;
  assign n1750 = n1749 ^ n1744 ;
  assign n1739 = n1494 & n1528 ;
  assign n1740 = n1739 ^ n1494 ;
  assign n1741 = n1483 & n1740 ;
  assign n1751 = n1750 ^ n1741 ;
  assign n2324 = n2323 ^ n1751 ;
  assign n2321 = x41 & ~n2267 ;
  assign n2319 = n2170 & ~n2267 ;
  assign n2320 = n2319 ^ n2170 ;
  assign n2322 = n2321 ^ n2320 ;
  assign n2325 = n2324 ^ n2322 ;
  assign n2326 = n2318 & n2325 ;
  assign n2327 = n2326 ^ n2318 ;
  assign n2328 = n2327 ^ n2325 ;
  assign n2515 = n2317 & ~n2328 ;
  assign n2516 = n2374 & n2515 ;
  assign n2365 = ~n2322 & n2324 ;
  assign n2366 = ~n2318 & n2365 ;
  assign n2364 = n2313 & ~n2317 ;
  assign n2367 = n2366 ^ n2364 ;
  assign n2514 = n2317 & ~n2367 ;
  assign n2517 = n2516 ^ n2514 ;
  assign n2342 = n2341 ^ n2337 ;
  assign n2343 = n2335 & n2342 ;
  assign n2344 = n2343 ^ n2335 ;
  assign n2345 = n2344 ^ n2342 ;
  assign n2346 = n2328 & n2345 ;
  assign n2347 = n2346 ^ n2328 ;
  assign n2348 = n2347 ^ n2345 ;
  assign n2270 = x44 & ~n2267 ;
  assign n2268 = n2164 & ~n2267 ;
  assign n2269 = n2268 ^ n2164 ;
  assign n2271 = n2270 ^ n2269 ;
  assign n1570 = n1437 & ~n1504 ;
  assign n1571 = n1555 & n1570 ;
  assign n1569 = n1437 & n1548 ;
  assign n1572 = n1571 ^ n1569 ;
  assign n1573 = n1572 ^ n1437 ;
  assign n1566 = n1437 & n1541 ;
  assign n1567 = n1566 ^ n1437 ;
  assign n1568 = n1567 ^ n1437 ;
  assign n1574 = n1573 ^ n1568 ;
  assign n1563 = n1437 & n1528 ;
  assign n1564 = n1563 ^ n1437 ;
  assign n1565 = n1483 & n1564 ;
  assign n1575 = n1574 ^ n1565 ;
  assign n2161 = n1575 ^ n1437 ;
  assign n1556 = n1326 & ~n1504 ;
  assign n1557 = n1555 & n1556 ;
  assign n1549 = n1326 & n1548 ;
  assign n1558 = n1557 ^ n1549 ;
  assign n1559 = n1558 ^ n1326 ;
  assign n1542 = n1326 & n1541 ;
  assign n1543 = n1542 ^ n1326 ;
  assign n1544 = n1543 ^ n1326 ;
  assign n1560 = n1559 ^ n1544 ;
  assign n1529 = n1326 & n1528 ;
  assign n1530 = n1529 ^ n1326 ;
  assign n1531 = n1483 & n1530 ;
  assign n1561 = n1560 ^ n1531 ;
  assign n2162 = n2161 ^ n1561 ;
  assign n2273 = n2271 ^ n2162 ;
  assign n2278 = x45 & ~n2267 ;
  assign n2276 = n2210 & ~n2267 ;
  assign n2277 = n2276 ^ n2210 ;
  assign n2279 = n2278 ^ n2277 ;
  assign n1606 = n1447 & ~n1504 ;
  assign n1607 = n1555 & n1606 ;
  assign n1605 = n1447 & n1548 ;
  assign n1608 = n1607 ^ n1605 ;
  assign n1609 = n1608 ^ n1447 ;
  assign n1602 = n1447 & n1541 ;
  assign n1603 = n1602 ^ n1447 ;
  assign n1604 = n1603 ^ n1447 ;
  assign n1610 = n1609 ^ n1604 ;
  assign n1599 = n1447 & n1528 ;
  assign n1600 = n1599 ^ n1447 ;
  assign n1601 = n1483 & n1600 ;
  assign n1611 = n1610 ^ n1601 ;
  assign n2274 = n1611 ^ n1447 ;
  assign n1592 = n1441 & ~n1504 ;
  assign n1593 = n1555 & n1592 ;
  assign n1591 = n1441 & n1548 ;
  assign n1594 = n1593 ^ n1591 ;
  assign n1595 = n1594 ^ n1441 ;
  assign n1588 = n1441 & n1541 ;
  assign n1589 = n1588 ^ n1441 ;
  assign n1590 = n1589 ^ n1441 ;
  assign n1596 = n1595 ^ n1590 ;
  assign n1585 = n1441 & n1528 ;
  assign n1586 = n1585 ^ n1441 ;
  assign n1587 = n1483 & n1586 ;
  assign n1597 = n1596 ^ n1587 ;
  assign n2275 = n2274 ^ n1597 ;
  assign n2285 = n2279 ^ n2275 ;
  assign n2286 = n2273 & n2285 ;
  assign n2287 = n2286 ^ n2273 ;
  assign n2288 = n2287 ^ n2285 ;
  assign n2293 = x46 & ~n2267 ;
  assign n2291 = n2255 & ~n2267 ;
  assign n2292 = n2291 ^ n2255 ;
  assign n2294 = n2293 ^ n2292 ;
  assign n1649 = n1464 & ~n1504 ;
  assign n1650 = n1555 & n1649 ;
  assign n1648 = n1464 & n1548 ;
  assign n1651 = n1650 ^ n1648 ;
  assign n1652 = n1651 ^ n1464 ;
  assign n1645 = n1464 & n1541 ;
  assign n1646 = n1645 ^ n1464 ;
  assign n1647 = n1646 ^ n1464 ;
  assign n1653 = n1652 ^ n1647 ;
  assign n1642 = n1464 & n1528 ;
  assign n1643 = n1642 ^ n1464 ;
  assign n1644 = n1483 & n1643 ;
  assign n1654 = n1653 ^ n1644 ;
  assign n2289 = n1654 ^ n1464 ;
  assign n1635 = n1458 & ~n1504 ;
  assign n1636 = n1555 & n1635 ;
  assign n1634 = n1458 & n1548 ;
  assign n1637 = n1636 ^ n1634 ;
  assign n1638 = n1637 ^ n1458 ;
  assign n1631 = n1458 & n1541 ;
  assign n1632 = n1631 ^ n1458 ;
  assign n1633 = n1632 ^ n1458 ;
  assign n1639 = n1638 ^ n1633 ;
  assign n1628 = n1458 & n1528 ;
  assign n1629 = n1628 ^ n1458 ;
  assign n1630 = n1483 & n1629 ;
  assign n1640 = n1639 ^ n1630 ;
  assign n2290 = n2289 ^ n1640 ;
  assign n2297 = n2294 ^ n2290 ;
  assign n2302 = x47 & ~n2267 ;
  assign n2300 = n2237 & ~n2267 ;
  assign n2301 = n2300 ^ n2237 ;
  assign n2303 = n2302 ^ n2301 ;
  assign n1680 = n1473 & ~n1504 ;
  assign n1681 = n1555 & n1680 ;
  assign n1679 = n1473 & n1548 ;
  assign n1682 = n1681 ^ n1679 ;
  assign n1683 = n1682 ^ n1473 ;
  assign n1676 = n1473 & n1541 ;
  assign n1677 = n1676 ^ n1473 ;
  assign n1678 = n1677 ^ n1473 ;
  assign n1684 = n1683 ^ n1678 ;
  assign n1673 = n1473 & n1528 ;
  assign n1674 = n1673 ^ n1473 ;
  assign n1675 = n1483 & n1674 ;
  assign n1685 = n1684 ^ n1675 ;
  assign n2298 = n1685 ^ n1473 ;
  assign n1666 = n1475 & ~n1504 ;
  assign n1667 = n1555 & n1666 ;
  assign n1665 = n1475 & n1548 ;
  assign n1668 = n1667 ^ n1665 ;
  assign n1669 = n1668 ^ n1475 ;
  assign n1662 = n1475 & n1541 ;
  assign n1663 = n1662 ^ n1475 ;
  assign n1664 = n1663 ^ n1475 ;
  assign n1670 = n1669 ^ n1664 ;
  assign n1659 = n1475 & n1528 ;
  assign n1660 = n1659 ^ n1475 ;
  assign n1661 = n1483 & n1660 ;
  assign n1671 = n1670 ^ n1661 ;
  assign n2299 = n2298 ^ n1671 ;
  assign n2352 = n2303 ^ n2299 ;
  assign n2353 = n2297 & n2352 ;
  assign n2354 = n2353 ^ n2297 ;
  assign n2355 = n2354 ^ n2352 ;
  assign n2356 = n2288 & n2355 ;
  assign n2357 = n2356 ^ n2288 ;
  assign n2358 = n2357 ^ n2355 ;
  assign n2359 = n2348 & n2358 ;
  assign n2360 = n2359 ^ n2348 ;
  assign n2361 = n2360 ^ n2358 ;
  assign n2512 = n2317 & ~n2361 ;
  assign n2513 = n2512 ^ n2317 ;
  assign n2518 = n2517 ^ n2513 ;
  assign n2304 = n2299 & n2303 ;
  assign n2305 = n2304 ^ n2299 ;
  assign n2306 = n2297 & n2305 ;
  assign n2307 = n2306 ^ n2305 ;
  assign n2295 = n2290 & n2294 ;
  assign n2296 = n2295 ^ n2290 ;
  assign n2308 = n2307 ^ n2296 ;
  assign n2309 = n2288 & n2308 ;
  assign n2310 = n2309 ^ n2308 ;
  assign n2280 = n2275 & n2279 ;
  assign n2281 = n2280 ^ n2275 ;
  assign n2282 = n2273 & n2281 ;
  assign n2283 = n2282 ^ n2281 ;
  assign n2272 = n2162 & ~n2271 ;
  assign n2284 = n2283 ^ n2272 ;
  assign n2311 = n2310 ^ n2284 ;
  assign n2509 = n2317 & n2348 ;
  assign n2510 = n2509 ^ n2317 ;
  assign n2511 = n2311 & n2510 ;
  assign n2519 = n2518 ^ n2511 ;
  assign n2503 = n2313 & ~n2328 ;
  assign n2504 = n2374 & n2503 ;
  assign n2502 = n2313 & ~n2367 ;
  assign n2505 = n2504 ^ n2502 ;
  assign n2500 = n2313 & ~n2361 ;
  assign n2501 = n2500 ^ n2313 ;
  assign n2506 = n2505 ^ n2501 ;
  assign n2497 = n2313 & n2348 ;
  assign n2498 = n2497 ^ n2313 ;
  assign n2499 = n2311 & n2498 ;
  assign n2507 = n2506 ^ n2499 ;
  assign n2508 = n2507 ^ n2313 ;
  assign n2520 = n2519 ^ n2508 ;
  assign n1059 = n949 ^ n947 ;
  assign n1020 = n914 ^ n912 ;
  assign n1005 = n1004 ^ n916 ;
  assign n1019 = n1018 ^ n1005 ;
  assign n1022 = n1020 ^ n1019 ;
  assign n1051 = n927 ^ n925 ;
  assign n1036 = n1035 ^ n929 ;
  assign n1050 = n1049 ^ n1036 ;
  assign n1055 = n1051 ^ n1050 ;
  assign n1056 = n1022 & n1055 ;
  assign n1057 = n1056 ^ n1022 ;
  assign n1058 = n1057 ^ n1055 ;
  assign n1073 = n1072 ^ n951 ;
  assign n1087 = n1086 ^ n1073 ;
  assign n1089 = n1087 ^ n1059 ;
  assign n1104 = n1103 ^ n958 ;
  assign n1118 = n1117 ^ n1104 ;
  assign n1090 = n956 ^ n954 ;
  assign n1127 = n1118 ^ n1090 ;
  assign n1128 = n1089 & n1127 ;
  assign n1129 = n1128 ^ n1089 ;
  assign n1130 = n1129 ^ n1127 ;
  assign n1131 = n1058 & n1130 ;
  assign n1132 = n1131 ^ n1058 ;
  assign n1133 = n1132 ^ n1130 ;
  assign n1148 = n1147 ^ n696 ;
  assign n1162 = n1161 ^ n1148 ;
  assign n1134 = n694 ^ n692 ;
  assign n1164 = n1162 ^ n1134 ;
  assign n1179 = n1178 ^ n863 ;
  assign n1193 = n1192 ^ n1179 ;
  assign n1165 = n861 ^ n859 ;
  assign n1199 = n1193 ^ n1165 ;
  assign n1200 = n1164 & n1199 ;
  assign n1201 = n1200 ^ n1164 ;
  assign n1202 = n1201 ^ n1199 ;
  assign n1217 = n1216 ^ n882 ;
  assign n1231 = n1230 ^ n1217 ;
  assign n1203 = n880 ^ n878 ;
  assign n1234 = n1231 ^ n1203 ;
  assign n1289 = n1288 ^ n902 ;
  assign n1303 = n1302 ^ n1289 ;
  assign n1235 = n900 ^ n898 ;
  assign n1304 = n1303 ^ n1235 ;
  assign n1305 = n1234 & n1304 ;
  assign n1306 = n1305 ^ n1234 ;
  assign n1307 = n1306 ^ n1304 ;
  assign n1308 = n1202 & n1307 ;
  assign n1309 = n1308 ^ n1202 ;
  assign n1310 = n1309 ^ n1307 ;
  assign n1311 = n1133 & n1310 ;
  assign n1312 = n1311 ^ n1133 ;
  assign n1313 = n1312 ^ n1310 ;
  assign n1251 = n896 & n1235 ;
  assign n1259 = ~n939 & n1251 ;
  assign n1260 = n998 & n1259 ;
  assign n1258 = n991 & n1251 ;
  assign n1261 = n1260 ^ n1258 ;
  assign n1262 = n1261 ^ n1251 ;
  assign n1255 = n984 & n1251 ;
  assign n1256 = n1255 ^ n1251 ;
  assign n1257 = n1256 ^ n1251 ;
  assign n1263 = n1262 ^ n1257 ;
  assign n1252 = n971 & n1251 ;
  assign n1253 = n1252 ^ n1251 ;
  assign n1254 = n910 & n1253 ;
  assign n1264 = n1263 ^ n1254 ;
  assign n1236 = n902 & n1235 ;
  assign n1244 = ~n939 & n1236 ;
  assign n1245 = n998 & n1244 ;
  assign n1243 = n991 & n1236 ;
  assign n1246 = n1245 ^ n1243 ;
  assign n1247 = n1246 ^ n1236 ;
  assign n1240 = n984 & n1236 ;
  assign n1241 = n1240 ^ n1236 ;
  assign n1242 = n1241 ^ n1236 ;
  assign n1248 = n1247 ^ n1242 ;
  assign n1237 = n971 & n1236 ;
  assign n1238 = n1237 ^ n1236 ;
  assign n1239 = n910 & n1238 ;
  assign n1249 = n1248 ^ n1239 ;
  assign n1250 = n1249 ^ n1236 ;
  assign n1265 = n1264 ^ n1250 ;
  assign n1266 = n1265 ^ n1235 ;
  assign n1267 = n1234 & n1266 ;
  assign n1268 = n1267 ^ n1266 ;
  assign n1232 = n1203 & n1231 ;
  assign n1233 = n1232 ^ n1203 ;
  assign n1269 = n1268 ^ n1233 ;
  assign n1270 = n1202 & n1269 ;
  assign n1271 = n1270 ^ n1269 ;
  assign n1194 = n1165 & n1193 ;
  assign n1195 = n1194 ^ n1165 ;
  assign n1196 = n1164 & n1195 ;
  assign n1197 = n1196 ^ n1195 ;
  assign n1163 = n1134 & ~n1162 ;
  assign n1198 = n1197 ^ n1163 ;
  assign n1272 = n1271 ^ n1198 ;
  assign n1273 = n1133 & n1272 ;
  assign n1274 = n1273 ^ n1272 ;
  assign n1119 = n1090 & n1118 ;
  assign n1120 = n1119 ^ n1090 ;
  assign n1121 = n1089 & n1120 ;
  assign n1122 = n1121 ^ n1120 ;
  assign n1088 = n1059 & ~n1087 ;
  assign n1123 = n1122 ^ n1088 ;
  assign n1124 = n1058 & n1123 ;
  assign n1125 = n1124 ^ n1123 ;
  assign n1052 = ~n1050 & n1051 ;
  assign n1053 = ~n1022 & n1052 ;
  assign n1021 = ~n1019 & n1020 ;
  assign n1054 = n1053 ^ n1021 ;
  assign n1126 = n1125 ^ n1054 ;
  assign n1275 = n1274 ^ n1126 ;
  assign n1314 = n1313 ^ n1275 ;
  assign n1802 = n1059 & n1314 ;
  assign n1803 = n1802 ^ n1059 ;
  assign n1799 = n1087 & n1314 ;
  assign n1800 = n1799 ^ n1087 ;
  assign n1801 = n1800 ^ n1087 ;
  assign n1804 = n1803 ^ n1801 ;
  assign n1784 = n1783 ^ n1512 ;
  assign n1798 = n1797 ^ n1784 ;
  assign n1805 = n1804 ^ n1798 ;
  assign n1809 = n1090 & n1314 ;
  assign n1810 = n1809 ^ n1090 ;
  assign n1806 = n1118 & n1314 ;
  assign n1807 = n1806 ^ n1118 ;
  assign n1808 = n1807 ^ n1118 ;
  assign n1811 = n1810 ^ n1808 ;
  assign n1825 = n1824 ^ n1515 ;
  assign n1839 = n1838 ^ n1825 ;
  assign n1868 = n1811 & n1839 ;
  assign n1869 = n1868 ^ n1811 ;
  assign n1870 = n1805 & n1869 ;
  assign n1871 = n1870 ^ n1869 ;
  assign n1867 = ~n1798 & n1804 ;
  assign n1872 = n1871 ^ n1867 ;
  assign n1717 = n1716 ^ n1485 ;
  assign n1731 = n1730 ^ n1717 ;
  assign n1317 = n1020 & n1314 ;
  assign n1702 = n1317 ^ n1020 ;
  assign n1315 = n1019 & n1314 ;
  assign n1316 = n1315 ^ n1019 ;
  assign n1701 = n1316 ^ n1019 ;
  assign n1703 = n1702 ^ n1701 ;
  assign n1732 = n1731 ^ n1703 ;
  assign n1752 = n1751 ^ n1494 ;
  assign n1766 = n1765 ^ n1752 ;
  assign n1736 = n1051 & n1314 ;
  assign n1737 = n1736 ^ n1051 ;
  assign n1733 = n1050 & n1314 ;
  assign n1734 = n1733 ^ n1050 ;
  assign n1735 = n1734 ^ n1050 ;
  assign n1738 = n1737 ^ n1735 ;
  assign n1767 = n1766 ^ n1738 ;
  assign n1768 = n1732 & n1767 ;
  assign n1769 = n1768 ^ n1732 ;
  assign n1770 = n1769 ^ n1767 ;
  assign n1885 = n1731 & ~n1770 ;
  assign n1886 = n1872 & n1885 ;
  assign n1863 = n1738 & ~n1766 ;
  assign n1864 = ~n1732 & n1863 ;
  assign n1862 = n1703 & ~n1731 ;
  assign n1865 = n1864 ^ n1862 ;
  assign n1884 = n1731 & ~n1865 ;
  assign n1887 = n1886 ^ n1884 ;
  assign n1840 = n1839 ^ n1811 ;
  assign n1841 = n1805 & n1840 ;
  assign n1842 = n1841 ^ n1805 ;
  assign n1843 = n1842 ^ n1840 ;
  assign n1844 = n1770 & n1843 ;
  assign n1845 = n1844 ^ n1770 ;
  assign n1846 = n1845 ^ n1843 ;
  assign n1562 = n1561 ^ n1326 ;
  assign n1576 = n1575 ^ n1562 ;
  assign n1322 = n1134 & n1314 ;
  assign n1323 = n1322 ^ n1134 ;
  assign n1319 = n1162 & n1314 ;
  assign n1320 = n1319 ^ n1162 ;
  assign n1321 = n1320 ^ n1162 ;
  assign n1324 = n1323 ^ n1321 ;
  assign n1578 = n1576 ^ n1324 ;
  assign n1598 = n1597 ^ n1441 ;
  assign n1612 = n1611 ^ n1598 ;
  assign n1582 = n1165 & n1314 ;
  assign n1583 = n1582 ^ n1165 ;
  assign n1579 = n1193 & n1314 ;
  assign n1580 = n1579 ^ n1193 ;
  assign n1581 = n1580 ^ n1193 ;
  assign n1584 = n1583 ^ n1581 ;
  assign n1618 = n1612 ^ n1584 ;
  assign n1619 = n1578 & n1618 ;
  assign n1620 = n1619 ^ n1578 ;
  assign n1621 = n1620 ^ n1618 ;
  assign n1641 = n1640 ^ n1458 ;
  assign n1655 = n1654 ^ n1641 ;
  assign n1625 = n1203 & n1314 ;
  assign n1626 = n1625 ^ n1203 ;
  assign n1622 = n1231 & n1314 ;
  assign n1623 = n1622 ^ n1231 ;
  assign n1624 = n1623 ^ n1231 ;
  assign n1627 = n1626 ^ n1624 ;
  assign n1658 = n1655 ^ n1627 ;
  assign n1690 = n1235 & n1314 ;
  assign n1691 = n1690 ^ n1235 ;
  assign n1687 = n1303 & n1314 ;
  assign n1688 = n1687 ^ n1303 ;
  assign n1689 = n1688 ^ n1303 ;
  assign n1692 = n1691 ^ n1689 ;
  assign n1672 = n1671 ^ n1475 ;
  assign n1686 = n1685 ^ n1672 ;
  assign n1850 = n1692 ^ n1686 ;
  assign n1851 = n1658 & n1850 ;
  assign n1852 = n1851 ^ n1658 ;
  assign n1853 = n1852 ^ n1850 ;
  assign n1854 = n1621 & n1853 ;
  assign n1855 = n1854 ^ n1621 ;
  assign n1856 = n1855 ^ n1853 ;
  assign n1857 = n1846 & n1856 ;
  assign n1858 = n1857 ^ n1846 ;
  assign n1859 = n1858 ^ n1856 ;
  assign n1882 = n1731 & ~n1859 ;
  assign n1883 = n1882 ^ n1731 ;
  assign n1888 = n1887 ^ n1883 ;
  assign n1693 = n1686 & n1692 ;
  assign n1694 = n1693 ^ n1692 ;
  assign n1695 = n1658 & n1694 ;
  assign n1696 = n1695 ^ n1694 ;
  assign n1656 = n1627 & n1655 ;
  assign n1657 = n1656 ^ n1627 ;
  assign n1697 = n1696 ^ n1657 ;
  assign n1698 = n1621 & n1697 ;
  assign n1699 = n1698 ^ n1697 ;
  assign n1613 = n1584 & n1612 ;
  assign n1614 = n1613 ^ n1584 ;
  assign n1615 = n1578 & n1614 ;
  assign n1616 = n1615 ^ n1614 ;
  assign n1577 = n1324 & ~n1576 ;
  assign n1617 = n1616 ^ n1577 ;
  assign n1700 = n1699 ^ n1617 ;
  assign n1879 = n1731 & n1846 ;
  assign n1880 = n1879 ^ n1731 ;
  assign n1881 = n1700 & n1880 ;
  assign n1889 = n1888 ^ n1881 ;
  assign n2495 = n1889 ^ n1731 ;
  assign n1873 = n1703 & ~n1770 ;
  assign n1874 = n1872 & n1873 ;
  assign n1866 = n1703 & ~n1865 ;
  assign n1875 = n1874 ^ n1866 ;
  assign n1860 = n1703 & ~n1859 ;
  assign n1861 = n1860 ^ n1703 ;
  assign n1876 = n1875 ^ n1861 ;
  assign n1847 = n1703 & n1846 ;
  assign n1848 = n1847 ^ n1703 ;
  assign n1849 = n1700 & n1848 ;
  assign n1877 = n1876 ^ n1849 ;
  assign n2496 = n2495 ^ n1877 ;
  assign n2521 = n2520 ^ n2496 ;
  assign n2542 = n2322 & ~n2328 ;
  assign n2543 = n2374 & n2542 ;
  assign n2541 = n2322 & ~n2367 ;
  assign n2544 = n2543 ^ n2541 ;
  assign n2539 = n2322 & ~n2361 ;
  assign n2540 = n2539 ^ n2322 ;
  assign n2545 = n2544 ^ n2540 ;
  assign n2536 = n2322 & n2348 ;
  assign n2537 = n2536 ^ n2322 ;
  assign n2538 = n2311 & n2537 ;
  assign n2546 = n2545 ^ n2538 ;
  assign n2530 = n2324 & ~n2328 ;
  assign n2531 = n2374 & n2530 ;
  assign n2529 = n2324 & ~n2367 ;
  assign n2532 = n2531 ^ n2529 ;
  assign n2527 = n2324 & ~n2361 ;
  assign n2528 = n2527 ^ n2324 ;
  assign n2533 = n2532 ^ n2528 ;
  assign n2524 = n2324 & n2348 ;
  assign n2525 = n2524 ^ n2324 ;
  assign n2526 = n2311 & n2525 ;
  assign n2534 = n2533 ^ n2526 ;
  assign n2535 = n2534 ^ n2324 ;
  assign n2547 = n2546 ^ n2535 ;
  assign n1911 = n1766 & ~n1770 ;
  assign n1912 = n1872 & n1911 ;
  assign n1910 = n1766 & ~n1865 ;
  assign n1913 = n1912 ^ n1910 ;
  assign n1908 = n1766 & ~n1859 ;
  assign n1909 = n1908 ^ n1766 ;
  assign n1914 = n1913 ^ n1909 ;
  assign n1905 = n1766 & n1846 ;
  assign n1906 = n1905 ^ n1766 ;
  assign n1907 = n1700 & n1906 ;
  assign n1915 = n1914 ^ n1907 ;
  assign n2522 = n1915 ^ n1766 ;
  assign n1899 = n1738 & ~n1770 ;
  assign n1900 = n1872 & n1899 ;
  assign n1898 = n1738 & ~n1865 ;
  assign n1901 = n1900 ^ n1898 ;
  assign n1896 = n1738 & ~n1859 ;
  assign n1897 = n1896 ^ n1738 ;
  assign n1902 = n1901 ^ n1897 ;
  assign n1893 = n1738 & n1846 ;
  assign n1894 = n1893 ^ n1738 ;
  assign n1895 = n1700 & n1894 ;
  assign n1903 = n1902 ^ n1895 ;
  assign n2523 = n2522 ^ n1903 ;
  assign n2548 = n2547 ^ n2523 ;
  assign n2549 = n2521 & n2548 ;
  assign n2550 = n2549 ^ n2521 ;
  assign n2551 = n2550 ^ n2548 ;
  assign n2572 = ~n2328 & n2332 ;
  assign n2573 = n2374 & n2572 ;
  assign n2571 = n2332 & ~n2367 ;
  assign n2574 = n2573 ^ n2571 ;
  assign n2569 = n2332 & ~n2361 ;
  assign n2570 = n2569 ^ n2332 ;
  assign n2575 = n2574 ^ n2570 ;
  assign n2566 = n2332 & n2348 ;
  assign n2567 = n2566 ^ n2332 ;
  assign n2568 = n2311 & n2567 ;
  assign n2576 = n2575 ^ n2568 ;
  assign n2560 = ~n2328 & n2334 ;
  assign n2561 = n2374 & n2560 ;
  assign n2559 = n2334 & ~n2367 ;
  assign n2562 = n2561 ^ n2559 ;
  assign n2557 = n2334 & ~n2361 ;
  assign n2558 = n2557 ^ n2334 ;
  assign n2563 = n2562 ^ n2558 ;
  assign n2554 = n2334 & n2348 ;
  assign n2555 = n2554 ^ n2334 ;
  assign n2556 = n2311 & n2555 ;
  assign n2564 = n2563 ^ n2556 ;
  assign n2565 = n2564 ^ n2334 ;
  assign n2577 = n2576 ^ n2565 ;
  assign n1944 = ~n1770 & n1798 ;
  assign n1945 = n1872 & n1944 ;
  assign n1943 = n1798 & ~n1865 ;
  assign n1946 = n1945 ^ n1943 ;
  assign n1941 = n1798 & ~n1859 ;
  assign n1942 = n1941 ^ n1798 ;
  assign n1947 = n1946 ^ n1942 ;
  assign n1938 = n1798 & n1846 ;
  assign n1939 = n1938 ^ n1798 ;
  assign n1940 = n1700 & n1939 ;
  assign n1948 = n1947 ^ n1940 ;
  assign n2552 = n1948 ^ n1798 ;
  assign n1932 = ~n1770 & n1804 ;
  assign n1933 = n1872 & n1932 ;
  assign n1931 = n1804 & ~n1865 ;
  assign n1934 = n1933 ^ n1931 ;
  assign n1929 = n1804 & ~n1859 ;
  assign n1930 = n1929 ^ n1804 ;
  assign n1935 = n1934 ^ n1930 ;
  assign n1926 = n1804 & n1846 ;
  assign n1927 = n1926 ^ n1804 ;
  assign n1928 = n1700 & n1927 ;
  assign n1936 = n1935 ^ n1928 ;
  assign n2553 = n2552 ^ n1936 ;
  assign n2578 = n2577 ^ n2553 ;
  assign n1971 = ~n1770 & n1839 ;
  assign n1972 = n1872 & n1971 ;
  assign n1970 = n1839 & ~n1865 ;
  assign n1973 = n1972 ^ n1970 ;
  assign n1968 = n1839 & ~n1859 ;
  assign n1969 = n1968 ^ n1839 ;
  assign n1974 = n1973 ^ n1969 ;
  assign n1965 = n1839 & n1846 ;
  assign n1966 = n1965 ^ n1839 ;
  assign n1967 = n1700 & n1966 ;
  assign n1975 = n1974 ^ n1967 ;
  assign n2579 = n1975 ^ n1839 ;
  assign n1959 = ~n1770 & n1811 ;
  assign n1960 = n1872 & n1959 ;
  assign n1958 = n1811 & ~n1865 ;
  assign n1961 = n1960 ^ n1958 ;
  assign n1956 = n1811 & ~n1859 ;
  assign n1957 = n1956 ^ n1811 ;
  assign n1962 = n1961 ^ n1957 ;
  assign n1953 = n1811 & n1846 ;
  assign n1954 = n1953 ^ n1811 ;
  assign n1955 = n1700 & n1954 ;
  assign n1963 = n1962 ^ n1955 ;
  assign n2580 = n2579 ^ n1963 ;
  assign n2599 = ~n2328 & n2341 ;
  assign n2600 = n2374 & n2599 ;
  assign n2598 = n2341 & ~n2367 ;
  assign n2601 = n2600 ^ n2598 ;
  assign n2596 = n2341 & ~n2361 ;
  assign n2597 = n2596 ^ n2341 ;
  assign n2602 = n2601 ^ n2597 ;
  assign n2593 = n2341 & n2348 ;
  assign n2594 = n2593 ^ n2341 ;
  assign n2595 = n2311 & n2594 ;
  assign n2603 = n2602 ^ n2595 ;
  assign n2587 = ~n2328 & n2337 ;
  assign n2588 = n2374 & n2587 ;
  assign n2586 = n2337 & ~n2367 ;
  assign n2589 = n2588 ^ n2586 ;
  assign n2584 = n2337 & ~n2361 ;
  assign n2585 = n2584 ^ n2337 ;
  assign n2590 = n2589 ^ n2585 ;
  assign n2581 = n2337 & n2348 ;
  assign n2582 = n2581 ^ n2337 ;
  assign n2583 = n2311 & n2582 ;
  assign n2591 = n2590 ^ n2583 ;
  assign n2592 = n2591 ^ n2337 ;
  assign n2604 = n2603 ^ n2592 ;
  assign n2629 = n2580 & n2604 ;
  assign n2630 = n2629 ^ n2580 ;
  assign n2631 = n2578 & n2630 ;
  assign n2632 = n2631 ^ n2630 ;
  assign n2628 = n2553 & ~n2577 ;
  assign n2633 = n2632 ^ n2628 ;
  assign n2634 = n2551 & n2633 ;
  assign n2635 = n2634 ^ n2633 ;
  assign n2625 = n2523 & ~n2547 ;
  assign n2626 = ~n2521 & n2625 ;
  assign n2624 = n2496 & ~n2520 ;
  assign n2627 = n2626 ^ n2624 ;
  assign n2636 = n2635 ^ n2627 ;
  assign n2747 = n2520 & n2636 ;
  assign n2748 = n2747 ^ n2520 ;
  assign n2605 = n2604 ^ n2580 ;
  assign n2606 = n2578 & n2605 ;
  assign n2607 = n2606 ^ n2578 ;
  assign n2608 = n2607 ^ n2605 ;
  assign n2609 = n2551 & n2608 ;
  assign n2610 = n2609 ^ n2551 ;
  assign n2611 = n2610 ^ n2608 ;
  assign n2387 = n2271 & ~n2328 ;
  assign n2388 = n2374 & n2387 ;
  assign n2386 = n2271 & ~n2367 ;
  assign n2389 = n2388 ^ n2386 ;
  assign n2384 = n2271 & ~n2361 ;
  assign n2385 = n2384 ^ n2271 ;
  assign n2390 = n2389 ^ n2385 ;
  assign n2381 = n2271 & n2348 ;
  assign n2382 = n2381 ^ n2271 ;
  assign n2383 = n2311 & n2382 ;
  assign n2391 = n2390 ^ n2383 ;
  assign n2375 = n2162 & ~n2328 ;
  assign n2376 = n2374 & n2375 ;
  assign n2368 = n2162 & ~n2367 ;
  assign n2377 = n2376 ^ n2368 ;
  assign n2362 = n2162 & ~n2361 ;
  assign n2363 = n2362 ^ n2162 ;
  assign n2378 = n2377 ^ n2363 ;
  assign n2349 = n2162 & n2348 ;
  assign n2350 = n2349 ^ n2162 ;
  assign n2351 = n2311 & n2350 ;
  assign n2379 = n2378 ^ n2351 ;
  assign n2380 = n2379 ^ n2162 ;
  assign n2392 = n2391 ^ n2380 ;
  assign n2011 = n1576 & ~n1770 ;
  assign n2012 = n1872 & n2011 ;
  assign n2010 = n1576 & ~n1865 ;
  assign n2013 = n2012 ^ n2010 ;
  assign n2008 = n1576 & ~n1859 ;
  assign n2009 = n2008 ^ n1576 ;
  assign n2014 = n2013 ^ n2009 ;
  assign n2005 = n1576 & n1846 ;
  assign n2006 = n2005 ^ n1576 ;
  assign n2007 = n1700 & n2006 ;
  assign n2015 = n2014 ^ n2007 ;
  assign n2159 = n2015 ^ n1576 ;
  assign n1999 = n1324 & ~n1770 ;
  assign n2000 = n1872 & n1999 ;
  assign n1998 = n1324 & ~n1865 ;
  assign n2001 = n2000 ^ n1998 ;
  assign n1996 = n1324 & ~n1859 ;
  assign n1997 = n1996 ^ n1324 ;
  assign n2002 = n2001 ^ n1997 ;
  assign n1993 = n1324 & n1846 ;
  assign n1994 = n1993 ^ n1324 ;
  assign n1995 = n1700 & n1994 ;
  assign n2003 = n2002 ^ n1995 ;
  assign n2160 = n2159 ^ n2003 ;
  assign n2394 = n2392 ^ n2160 ;
  assign n2415 = n2279 & ~n2328 ;
  assign n2416 = n2374 & n2415 ;
  assign n2414 = n2279 & ~n2367 ;
  assign n2417 = n2416 ^ n2414 ;
  assign n2412 = n2279 & ~n2361 ;
  assign n2413 = n2412 ^ n2279 ;
  assign n2418 = n2417 ^ n2413 ;
  assign n2409 = n2279 & n2348 ;
  assign n2410 = n2409 ^ n2279 ;
  assign n2411 = n2311 & n2410 ;
  assign n2419 = n2418 ^ n2411 ;
  assign n2403 = n2275 & ~n2328 ;
  assign n2404 = n2374 & n2403 ;
  assign n2402 = n2275 & ~n2367 ;
  assign n2405 = n2404 ^ n2402 ;
  assign n2400 = n2275 & ~n2361 ;
  assign n2401 = n2400 ^ n2275 ;
  assign n2406 = n2405 ^ n2401 ;
  assign n2397 = n2275 & n2348 ;
  assign n2398 = n2397 ^ n2275 ;
  assign n2399 = n2311 & n2398 ;
  assign n2407 = n2406 ^ n2399 ;
  assign n2408 = n2407 ^ n2275 ;
  assign n2420 = n2419 ^ n2408 ;
  assign n2038 = n1612 & ~n1770 ;
  assign n2039 = n1872 & n2038 ;
  assign n2037 = n1612 & ~n1865 ;
  assign n2040 = n2039 ^ n2037 ;
  assign n2035 = n1612 & ~n1859 ;
  assign n2036 = n2035 ^ n1612 ;
  assign n2041 = n2040 ^ n2036 ;
  assign n2032 = n1612 & n1846 ;
  assign n2033 = n2032 ^ n1612 ;
  assign n2034 = n1700 & n2033 ;
  assign n2042 = n2041 ^ n2034 ;
  assign n2395 = n2042 ^ n1612 ;
  assign n2026 = n1584 & ~n1770 ;
  assign n2027 = n1872 & n2026 ;
  assign n2025 = n1584 & ~n1865 ;
  assign n2028 = n2027 ^ n2025 ;
  assign n2023 = n1584 & ~n1859 ;
  assign n2024 = n2023 ^ n1584 ;
  assign n2029 = n2028 ^ n2024 ;
  assign n2020 = n1584 & n1846 ;
  assign n2021 = n2020 ^ n1584 ;
  assign n2022 = n1700 & n2021 ;
  assign n2030 = n2029 ^ n2022 ;
  assign n2396 = n2395 ^ n2030 ;
  assign n2426 = n2420 ^ n2396 ;
  assign n2427 = n2394 & n2426 ;
  assign n2428 = n2427 ^ n2394 ;
  assign n2429 = n2428 ^ n2426 ;
  assign n2450 = n2294 & ~n2328 ;
  assign n2451 = n2374 & n2450 ;
  assign n2449 = n2294 & ~n2367 ;
  assign n2452 = n2451 ^ n2449 ;
  assign n2447 = n2294 & ~n2361 ;
  assign n2448 = n2447 ^ n2294 ;
  assign n2453 = n2452 ^ n2448 ;
  assign n2444 = n2294 & n2348 ;
  assign n2445 = n2444 ^ n2294 ;
  assign n2446 = n2311 & n2445 ;
  assign n2454 = n2453 ^ n2446 ;
  assign n2438 = n2290 & ~n2328 ;
  assign n2439 = n2374 & n2438 ;
  assign n2437 = n2290 & ~n2367 ;
  assign n2440 = n2439 ^ n2437 ;
  assign n2435 = n2290 & ~n2361 ;
  assign n2436 = n2435 ^ n2290 ;
  assign n2441 = n2440 ^ n2436 ;
  assign n2432 = n2290 & n2348 ;
  assign n2433 = n2432 ^ n2290 ;
  assign n2434 = n2311 & n2433 ;
  assign n2442 = n2441 ^ n2434 ;
  assign n2443 = n2442 ^ n2290 ;
  assign n2455 = n2454 ^ n2443 ;
  assign n2072 = n1655 & ~n1770 ;
  assign n2073 = n1872 & n2072 ;
  assign n2071 = n1655 & ~n1865 ;
  assign n2074 = n2073 ^ n2071 ;
  assign n2069 = n1655 & ~n1859 ;
  assign n2070 = n2069 ^ n1655 ;
  assign n2075 = n2074 ^ n2070 ;
  assign n2066 = n1655 & n1846 ;
  assign n2067 = n2066 ^ n1655 ;
  assign n2068 = n1700 & n2067 ;
  assign n2076 = n2075 ^ n2068 ;
  assign n2430 = n2076 ^ n1655 ;
  assign n2060 = n1627 & ~n1770 ;
  assign n2061 = n1872 & n2060 ;
  assign n2059 = n1627 & ~n1865 ;
  assign n2062 = n2061 ^ n2059 ;
  assign n2057 = n1627 & ~n1859 ;
  assign n2058 = n2057 ^ n1627 ;
  assign n2063 = n2062 ^ n2058 ;
  assign n2054 = n1627 & n1846 ;
  assign n2055 = n2054 ^ n1627 ;
  assign n2056 = n1700 & n2055 ;
  assign n2064 = n2063 ^ n2056 ;
  assign n2431 = n2430 ^ n2064 ;
  assign n2458 = n2455 ^ n2431 ;
  assign n2480 = n2303 & ~n2328 ;
  assign n2481 = n2374 & n2480 ;
  assign n2479 = n2303 & n2367 ;
  assign n2482 = n2481 ^ n2479 ;
  assign n2483 = n2482 ^ n2303 ;
  assign n2477 = n2303 & ~n2361 ;
  assign n2478 = n2477 ^ n2303 ;
  assign n2484 = n2483 ^ n2478 ;
  assign n2474 = n2303 & n2348 ;
  assign n2475 = n2474 ^ n2303 ;
  assign n2476 = n2311 & n2475 ;
  assign n2485 = n2484 ^ n2476 ;
  assign n2467 = n2299 & ~n2328 ;
  assign n2468 = n2374 & n2467 ;
  assign n2466 = n2299 & n2367 ;
  assign n2469 = n2468 ^ n2466 ;
  assign n2470 = n2469 ^ n2299 ;
  assign n2464 = n2299 & ~n2361 ;
  assign n2465 = n2464 ^ n2299 ;
  assign n2471 = n2470 ^ n2465 ;
  assign n2461 = n2299 & n2348 ;
  assign n2462 = n2461 ^ n2299 ;
  assign n2463 = n2311 & n2462 ;
  assign n2472 = n2471 ^ n2463 ;
  assign n2473 = n2472 ^ n2299 ;
  assign n2486 = n2485 ^ n2473 ;
  assign n2136 = n1686 & ~n1770 ;
  assign n2137 = n1872 & n2136 ;
  assign n2135 = n1686 & n1865 ;
  assign n2138 = n2137 ^ n2135 ;
  assign n2139 = n2138 ^ n1686 ;
  assign n2133 = n1686 & ~n1859 ;
  assign n2134 = n2133 ^ n1686 ;
  assign n2140 = n2139 ^ n2134 ;
  assign n2130 = n1686 & n1846 ;
  assign n2131 = n2130 ^ n1686 ;
  assign n2132 = n1700 & n2131 ;
  assign n2141 = n2140 ^ n2132 ;
  assign n2459 = n2141 ^ n1686 ;
  assign n2123 = n1692 & ~n1770 ;
  assign n2124 = n1872 & n2123 ;
  assign n2122 = n1692 & n1865 ;
  assign n2125 = n2124 ^ n2122 ;
  assign n2126 = n2125 ^ n1692 ;
  assign n2120 = n1692 & ~n1859 ;
  assign n2121 = n2120 ^ n1692 ;
  assign n2127 = n2126 ^ n2121 ;
  assign n2117 = n1692 & n1846 ;
  assign n2118 = n2117 ^ n1692 ;
  assign n2119 = n1700 & n2118 ;
  assign n2128 = n2127 ^ n2119 ;
  assign n2460 = n2459 ^ n2128 ;
  assign n2614 = n2486 ^ n2460 ;
  assign n2615 = n2458 & n2614 ;
  assign n2616 = n2615 ^ n2458 ;
  assign n2617 = n2616 ^ n2614 ;
  assign n2618 = n2429 & n2617 ;
  assign n2619 = n2618 ^ n2429 ;
  assign n2620 = n2619 ^ n2617 ;
  assign n2621 = ~n2611 & ~n2620 ;
  assign n2745 = n2520 & n2621 ;
  assign n2746 = n2745 ^ n2520 ;
  assign n2749 = n2748 ^ n2746 ;
  assign n2487 = n2460 & n2486 ;
  assign n2488 = n2487 ^ n2460 ;
  assign n2489 = n2458 & n2488 ;
  assign n2490 = n2489 ^ n2488 ;
  assign n2456 = n2431 & n2455 ;
  assign n2457 = n2456 ^ n2431 ;
  assign n2491 = n2490 ^ n2457 ;
  assign n2492 = n2429 & n2491 ;
  assign n2493 = n2492 ^ n2491 ;
  assign n2421 = n2396 & n2420 ;
  assign n2422 = n2421 ^ n2396 ;
  assign n2423 = n2394 & n2422 ;
  assign n2424 = n2423 ^ n2422 ;
  assign n2393 = n2160 & ~n2392 ;
  assign n2425 = n2424 ^ n2393 ;
  assign n2494 = n2493 ^ n2425 ;
  assign n2743 = n2520 & ~n2611 ;
  assign n2744 = n2494 & n2743 ;
  assign n2750 = n2749 ^ n2744 ;
  assign n2740 = n2496 & n2636 ;
  assign n2738 = n2496 & n2621 ;
  assign n2739 = n2738 ^ n2496 ;
  assign n2741 = n2740 ^ n2739 ;
  assign n2736 = n2496 & ~n2611 ;
  assign n2737 = n2494 & n2736 ;
  assign n2742 = n2741 ^ n2737 ;
  assign n2751 = n2750 ^ n2742 ;
  assign n1318 = n1317 ^ n1316 ;
  assign n1878 = n1877 ^ n1703 ;
  assign n1890 = n1889 ^ n1878 ;
  assign n1892 = n1890 ^ n1318 ;
  assign n1917 = n1736 ^ n1734 ;
  assign n1904 = n1903 ^ n1738 ;
  assign n1916 = n1915 ^ n1904 ;
  assign n1921 = n1917 ^ n1916 ;
  assign n1922 = n1892 & n1921 ;
  assign n1923 = n1922 ^ n1892 ;
  assign n1924 = n1923 ^ n1921 ;
  assign n1937 = n1936 ^ n1804 ;
  assign n1949 = n1948 ^ n1937 ;
  assign n1925 = n1802 ^ n1800 ;
  assign n1951 = n1949 ^ n1925 ;
  assign n1964 = n1963 ^ n1811 ;
  assign n1976 = n1975 ^ n1964 ;
  assign n1952 = n1809 ^ n1807 ;
  assign n1985 = n1976 ^ n1952 ;
  assign n1986 = n1951 & n1985 ;
  assign n1987 = n1986 ^ n1951 ;
  assign n1988 = n1987 ^ n1985 ;
  assign n1989 = n1924 & n1988 ;
  assign n1990 = n1989 ^ n1924 ;
  assign n1991 = n1990 ^ n1988 ;
  assign n2004 = n2003 ^ n1324 ;
  assign n2016 = n2015 ^ n2004 ;
  assign n1992 = n1322 ^ n1320 ;
  assign n2018 = n2016 ^ n1992 ;
  assign n2031 = n2030 ^ n1584 ;
  assign n2043 = n2042 ^ n2031 ;
  assign n2019 = n1582 ^ n1580 ;
  assign n2049 = n2043 ^ n2019 ;
  assign n2050 = n2018 & n2049 ;
  assign n2051 = n2050 ^ n2018 ;
  assign n2052 = n2051 ^ n2049 ;
  assign n2065 = n2064 ^ n1627 ;
  assign n2077 = n2076 ^ n2065 ;
  assign n2053 = n1625 ^ n1623 ;
  assign n2080 = n2077 ^ n2053 ;
  assign n2129 = n2128 ^ n1692 ;
  assign n2142 = n2141 ^ n2129 ;
  assign n2081 = n1690 ^ n1688 ;
  assign n2143 = n2142 ^ n2081 ;
  assign n2144 = n2080 & n2143 ;
  assign n2145 = n2144 ^ n2080 ;
  assign n2146 = n2145 ^ n2143 ;
  assign n2147 = n2052 & n2146 ;
  assign n2148 = n2147 ^ n2052 ;
  assign n2149 = n2148 ^ n2146 ;
  assign n2150 = ~n1991 & ~n2149 ;
  assign n2095 = n1686 & n2081 ;
  assign n2102 = ~n1770 & n2095 ;
  assign n2103 = n1872 & n2102 ;
  assign n2101 = ~n1865 & n2095 ;
  assign n2104 = n2103 ^ n2101 ;
  assign n2099 = ~n1859 & n2095 ;
  assign n2100 = n2099 ^ n2095 ;
  assign n2105 = n2104 ^ n2100 ;
  assign n2096 = n1846 & n2095 ;
  assign n2097 = n2096 ^ n2095 ;
  assign n2098 = n1700 & n2097 ;
  assign n2106 = n2105 ^ n2098 ;
  assign n2082 = n1692 & n2081 ;
  assign n2089 = ~n1770 & n2082 ;
  assign n2090 = n1872 & n2089 ;
  assign n2088 = ~n1865 & n2082 ;
  assign n2091 = n2090 ^ n2088 ;
  assign n2086 = ~n1859 & n2082 ;
  assign n2087 = n2086 ^ n2082 ;
  assign n2092 = n2091 ^ n2087 ;
  assign n2083 = n1846 & n2082 ;
  assign n2084 = n2083 ^ n2082 ;
  assign n2085 = n1700 & n2084 ;
  assign n2093 = n2092 ^ n2085 ;
  assign n2094 = n2093 ^ n2082 ;
  assign n2107 = n2106 ^ n2094 ;
  assign n2108 = n2107 ^ n2081 ;
  assign n2109 = n2080 & n2108 ;
  assign n2110 = n2109 ^ n2108 ;
  assign n2078 = n2053 & n2077 ;
  assign n2079 = n2078 ^ n2053 ;
  assign n2111 = n2110 ^ n2079 ;
  assign n2112 = n2052 & n2111 ;
  assign n2113 = n2112 ^ n2111 ;
  assign n2044 = n2019 & n2043 ;
  assign n2045 = n2044 ^ n2019 ;
  assign n2046 = n2018 & n2045 ;
  assign n2047 = n2046 ^ n2045 ;
  assign n2017 = n1992 & ~n2016 ;
  assign n2048 = n2047 ^ n2017 ;
  assign n2114 = n2113 ^ n2048 ;
  assign n2115 = ~n1991 & n2114 ;
  assign n1977 = n1952 & n1976 ;
  assign n1978 = n1977 ^ n1952 ;
  assign n1979 = n1951 & n1978 ;
  assign n1980 = n1979 ^ n1978 ;
  assign n1950 = n1925 & ~n1949 ;
  assign n1981 = n1980 ^ n1950 ;
  assign n1982 = n1924 & n1981 ;
  assign n1983 = n1982 ^ n1981 ;
  assign n1918 = ~n1916 & n1917 ;
  assign n1919 = ~n1892 & n1918 ;
  assign n1891 = n1318 & ~n1890 ;
  assign n1920 = n1919 ^ n1891 ;
  assign n1984 = n1983 ^ n1920 ;
  assign n2116 = n2115 ^ n1984 ;
  assign n2151 = n2150 ^ n2116 ;
  assign n2734 = n1318 & n2151 ;
  assign n2153 = n1890 & n2151 ;
  assign n2733 = n2153 ^ n1890 ;
  assign n2735 = n2734 ^ n2733 ;
  assign n2752 = n2751 ^ n2735 ;
  assign n2768 = n2547 & n2636 ;
  assign n2769 = n2768 ^ n2547 ;
  assign n2766 = n2547 & n2621 ;
  assign n2767 = n2766 ^ n2547 ;
  assign n2770 = n2769 ^ n2767 ;
  assign n2764 = n2547 & ~n2611 ;
  assign n2765 = n2494 & n2764 ;
  assign n2771 = n2770 ^ n2765 ;
  assign n2761 = n2523 & n2636 ;
  assign n2759 = n2523 & n2621 ;
  assign n2760 = n2759 ^ n2523 ;
  assign n2762 = n2761 ^ n2760 ;
  assign n2757 = n2523 & ~n2611 ;
  assign n2758 = n2494 & n2757 ;
  assign n2763 = n2762 ^ n2758 ;
  assign n2772 = n2771 ^ n2763 ;
  assign n2755 = n1917 & n2151 ;
  assign n2753 = n1916 & n2151 ;
  assign n2754 = n2753 ^ n1916 ;
  assign n2756 = n2755 ^ n2754 ;
  assign n2773 = n2772 ^ n2756 ;
  assign n2774 = n2752 & n2773 ;
  assign n2775 = n2774 ^ n2752 ;
  assign n2776 = n2775 ^ n2773 ;
  assign n2792 = n2577 & n2636 ;
  assign n2793 = n2792 ^ n2577 ;
  assign n2790 = n2577 & n2621 ;
  assign n2791 = n2790 ^ n2577 ;
  assign n2794 = n2793 ^ n2791 ;
  assign n2788 = n2577 & ~n2611 ;
  assign n2789 = n2494 & n2788 ;
  assign n2795 = n2794 ^ n2789 ;
  assign n2785 = n2553 & n2636 ;
  assign n2783 = n2553 & n2621 ;
  assign n2784 = n2783 ^ n2553 ;
  assign n2786 = n2785 ^ n2784 ;
  assign n2781 = n2553 & ~n2611 ;
  assign n2782 = n2494 & n2781 ;
  assign n2787 = n2786 ^ n2782 ;
  assign n2796 = n2795 ^ n2787 ;
  assign n2779 = n1925 & n2151 ;
  assign n2777 = n1949 & n2151 ;
  assign n2778 = n2777 ^ n1949 ;
  assign n2780 = n2779 ^ n2778 ;
  assign n2797 = n2796 ^ n2780 ;
  assign n2800 = n1952 & n2151 ;
  assign n2798 = n1976 & n2151 ;
  assign n2799 = n2798 ^ n1976 ;
  assign n2801 = n2800 ^ n2799 ;
  assign n2813 = n2604 & n2636 ;
  assign n2814 = n2813 ^ n2604 ;
  assign n2811 = n2604 & n2621 ;
  assign n2812 = n2811 ^ n2604 ;
  assign n2815 = n2814 ^ n2812 ;
  assign n2809 = n2604 & ~n2611 ;
  assign n2810 = n2494 & n2809 ;
  assign n2816 = n2815 ^ n2810 ;
  assign n2806 = n2580 & n2636 ;
  assign n2804 = n2580 & n2621 ;
  assign n2805 = n2804 ^ n2580 ;
  assign n2807 = n2806 ^ n2805 ;
  assign n2802 = n2580 & ~n2611 ;
  assign n2803 = n2494 & n2802 ;
  assign n2808 = n2807 ^ n2803 ;
  assign n2817 = n2816 ^ n2808 ;
  assign n2838 = n2801 & n2817 ;
  assign n2839 = n2838 ^ n2801 ;
  assign n2840 = n2797 & n2839 ;
  assign n2841 = n2840 ^ n2839 ;
  assign n2837 = n2780 & ~n2796 ;
  assign n2842 = n2841 ^ n2837 ;
  assign n2843 = ~n2776 & n2842 ;
  assign n2834 = n2756 & ~n2772 ;
  assign n2835 = ~n2752 & n2834 ;
  assign n2833 = n2735 & ~n2751 ;
  assign n2836 = n2835 ^ n2833 ;
  assign n2844 = n2843 ^ n2836 ;
  assign n2854 = n2751 & n2844 ;
  assign n2855 = n2854 ^ n2751 ;
  assign n2818 = n2817 ^ n2801 ;
  assign n2819 = n2797 & n2818 ;
  assign n2820 = n2819 ^ n2797 ;
  assign n2821 = n2820 ^ n2818 ;
  assign n2822 = ~n2776 & ~n2821 ;
  assign n2644 = n2392 & n2636 ;
  assign n2645 = n2644 ^ n2392 ;
  assign n2642 = n2392 & n2621 ;
  assign n2643 = n2642 ^ n2392 ;
  assign n2646 = n2645 ^ n2643 ;
  assign n2640 = n2392 & ~n2611 ;
  assign n2641 = n2494 & n2640 ;
  assign n2647 = n2646 ^ n2641 ;
  assign n2637 = n2160 & n2636 ;
  assign n2622 = n2160 & n2621 ;
  assign n2623 = n2622 ^ n2160 ;
  assign n2638 = n2637 ^ n2623 ;
  assign n2612 = n2160 & ~n2611 ;
  assign n2613 = n2494 & n2612 ;
  assign n2639 = n2638 ^ n2613 ;
  assign n2648 = n2647 ^ n2639 ;
  assign n2157 = n1992 & n2151 ;
  assign n2155 = n2016 & n2151 ;
  assign n2156 = n2155 ^ n2016 ;
  assign n2158 = n2157 ^ n2156 ;
  assign n2650 = n2648 ^ n2158 ;
  assign n2666 = n2420 & n2636 ;
  assign n2667 = n2666 ^ n2420 ;
  assign n2664 = n2420 & n2621 ;
  assign n2665 = n2664 ^ n2420 ;
  assign n2668 = n2667 ^ n2665 ;
  assign n2662 = n2420 & ~n2611 ;
  assign n2663 = n2494 & n2662 ;
  assign n2669 = n2668 ^ n2663 ;
  assign n2659 = n2396 & n2636 ;
  assign n2657 = n2396 & n2621 ;
  assign n2658 = n2657 ^ n2396 ;
  assign n2660 = n2659 ^ n2658 ;
  assign n2655 = n2396 & ~n2611 ;
  assign n2656 = n2494 & n2655 ;
  assign n2661 = n2660 ^ n2656 ;
  assign n2670 = n2669 ^ n2661 ;
  assign n2653 = n2019 & n2151 ;
  assign n2651 = n2043 & n2151 ;
  assign n2652 = n2651 ^ n2043 ;
  assign n2654 = n2653 ^ n2652 ;
  assign n2674 = n2670 ^ n2654 ;
  assign n2675 = n2650 & n2674 ;
  assign n2676 = n2675 ^ n2650 ;
  assign n2677 = n2676 ^ n2674 ;
  assign n2693 = n2455 & n2636 ;
  assign n2694 = n2693 ^ n2455 ;
  assign n2691 = n2455 & n2621 ;
  assign n2692 = n2691 ^ n2455 ;
  assign n2695 = n2694 ^ n2692 ;
  assign n2689 = n2455 & ~n2611 ;
  assign n2690 = n2494 & n2689 ;
  assign n2696 = n2695 ^ n2690 ;
  assign n2686 = n2431 & n2636 ;
  assign n2684 = n2431 & n2621 ;
  assign n2685 = n2684 ^ n2431 ;
  assign n2687 = n2686 ^ n2685 ;
  assign n2682 = n2431 & ~n2611 ;
  assign n2683 = n2494 & n2682 ;
  assign n2688 = n2687 ^ n2683 ;
  assign n2697 = n2696 ^ n2688 ;
  assign n2680 = n2053 & n2151 ;
  assign n2678 = n2077 & n2151 ;
  assign n2679 = n2678 ^ n2077 ;
  assign n2681 = n2680 ^ n2679 ;
  assign n2699 = n2697 ^ n2681 ;
  assign n2720 = n2486 & ~n2551 ;
  assign n2721 = n2633 & n2720 ;
  assign n2719 = n2486 & ~n2627 ;
  assign n2722 = n2721 ^ n2719 ;
  assign n2717 = n2486 & n2621 ;
  assign n2718 = n2717 ^ n2486 ;
  assign n2723 = n2722 ^ n2718 ;
  assign n2715 = n2486 & ~n2611 ;
  assign n2716 = n2494 & n2715 ;
  assign n2724 = n2723 ^ n2716 ;
  assign n2709 = n2460 & ~n2551 ;
  assign n2710 = n2633 & n2709 ;
  assign n2708 = n2460 & ~n2627 ;
  assign n2711 = n2710 ^ n2708 ;
  assign n2706 = n2460 & n2621 ;
  assign n2707 = n2706 ^ n2460 ;
  assign n2712 = n2711 ^ n2707 ;
  assign n2704 = n2460 & ~n2611 ;
  assign n2705 = n2494 & n2704 ;
  assign n2713 = n2712 ^ n2705 ;
  assign n2714 = n2713 ^ n2460 ;
  assign n2725 = n2724 ^ n2714 ;
  assign n2702 = n2081 & n2151 ;
  assign n2700 = n2142 & n2151 ;
  assign n2701 = n2700 ^ n2142 ;
  assign n2703 = n2702 ^ n2701 ;
  assign n2825 = n2725 ^ n2703 ;
  assign n2826 = n2699 & n2825 ;
  assign n2827 = n2826 ^ n2699 ;
  assign n2828 = n2827 ^ n2825 ;
  assign n2829 = ~n2677 & ~n2828 ;
  assign n2830 = n2822 & n2829 ;
  assign n2852 = n2751 & n2830 ;
  assign n2853 = n2852 ^ n2751 ;
  assign n2856 = n2855 ^ n2853 ;
  assign n2726 = n2703 & n2725 ;
  assign n2727 = n2726 ^ n2703 ;
  assign n2728 = n2699 & n2727 ;
  assign n2729 = n2728 ^ n2727 ;
  assign n2698 = n2681 & ~n2697 ;
  assign n2730 = n2729 ^ n2698 ;
  assign n2731 = ~n2677 & n2730 ;
  assign n2671 = n2654 & ~n2670 ;
  assign n2672 = ~n2650 & n2671 ;
  assign n2649 = n2158 & ~n2648 ;
  assign n2673 = n2672 ^ n2649 ;
  assign n2732 = n2731 ^ n2673 ;
  assign n2850 = n2751 & n2822 ;
  assign n2851 = n2732 & n2850 ;
  assign n2857 = n2856 ^ n2851 ;
  assign n2845 = n2735 & n2844 ;
  assign n2846 = n2845 ^ n2735 ;
  assign n2831 = n2735 & n2830 ;
  assign n2832 = n2831 ^ n2735 ;
  assign n2847 = n2846 ^ n2832 ;
  assign n2823 = n2735 & n2822 ;
  assign n2824 = n2732 & n2823 ;
  assign n2848 = n2847 ^ n2824 ;
  assign n2849 = n2848 ^ n2735 ;
  assign n2858 = n2857 ^ n2849 ;
  assign n2152 = n1318 & ~n2151 ;
  assign n2154 = n2153 ^ n2152 ;
  assign n2860 = n2858 ^ n2154 ;
  assign n2876 = n2772 & n2844 ;
  assign n2877 = n2876 ^ n2772 ;
  assign n2874 = n2772 & n2830 ;
  assign n2875 = n2874 ^ n2772 ;
  assign n2878 = n2877 ^ n2875 ;
  assign n2872 = n2772 & n2822 ;
  assign n2873 = n2732 & n2872 ;
  assign n2879 = n2878 ^ n2873 ;
  assign n2867 = n2756 & n2844 ;
  assign n2868 = n2867 ^ n2756 ;
  assign n2865 = n2756 & n2830 ;
  assign n2866 = n2865 ^ n2756 ;
  assign n2869 = n2868 ^ n2866 ;
  assign n2863 = n2756 & n2822 ;
  assign n2864 = n2732 & n2863 ;
  assign n2870 = n2869 ^ n2864 ;
  assign n2871 = n2870 ^ n2756 ;
  assign n2880 = n2879 ^ n2871 ;
  assign n2861 = n1917 & ~n2151 ;
  assign n2862 = n2861 ^ n2753 ;
  assign n2884 = n2880 ^ n2862 ;
  assign n2885 = n2860 & n2884 ;
  assign n2886 = n2885 ^ n2860 ;
  assign n2887 = n2886 ^ n2884 ;
  assign n2903 = n2796 & n2844 ;
  assign n2904 = n2903 ^ n2796 ;
  assign n2901 = n2796 & n2830 ;
  assign n2902 = n2901 ^ n2796 ;
  assign n2905 = n2904 ^ n2902 ;
  assign n2899 = n2796 & n2822 ;
  assign n2900 = n2732 & n2899 ;
  assign n2906 = n2905 ^ n2900 ;
  assign n2894 = n2780 & n2844 ;
  assign n2895 = n2894 ^ n2780 ;
  assign n2892 = n2780 & n2830 ;
  assign n2893 = n2892 ^ n2780 ;
  assign n2896 = n2895 ^ n2893 ;
  assign n2890 = n2780 & n2822 ;
  assign n2891 = n2732 & n2890 ;
  assign n2897 = n2896 ^ n2891 ;
  assign n2898 = n2897 ^ n2780 ;
  assign n2907 = n2906 ^ n2898 ;
  assign n2888 = n1925 & ~n2151 ;
  assign n2889 = n2888 ^ n2777 ;
  assign n2909 = n2907 ^ n2889 ;
  assign n2940 = n2817 & n2844 ;
  assign n2941 = n2940 ^ n2817 ;
  assign n2938 = n2817 & n2830 ;
  assign n2939 = n2938 ^ n2817 ;
  assign n2942 = n2941 ^ n2939 ;
  assign n2936 = n2817 & n2822 ;
  assign n2937 = n2732 & n2936 ;
  assign n2943 = n2942 ^ n2937 ;
  assign n2931 = n2801 & n2844 ;
  assign n2932 = n2931 ^ n2801 ;
  assign n2929 = n2801 & n2830 ;
  assign n2930 = n2929 ^ n2801 ;
  assign n2933 = n2932 ^ n2930 ;
  assign n2927 = n2801 & n2822 ;
  assign n2928 = n2732 & n2927 ;
  assign n2934 = n2933 ^ n2928 ;
  assign n2935 = n2934 ^ n2801 ;
  assign n2944 = n2943 ^ n2935 ;
  assign n2913 = n1952 & ~n2151 ;
  assign n2914 = n2913 ^ n2798 ;
  assign n2945 = n2944 ^ n2914 ;
  assign n2946 = n2909 & n2945 ;
  assign n2947 = n2946 ^ n2909 ;
  assign n2948 = n2947 ^ n2945 ;
  assign n2949 = n2887 & n2948 ;
  assign n2950 = n2949 ^ n2887 ;
  assign n2951 = n2950 ^ n2948 ;
  assign n2967 = n2648 & n2844 ;
  assign n2968 = n2967 ^ n2648 ;
  assign n2965 = n2648 & n2830 ;
  assign n2966 = n2965 ^ n2648 ;
  assign n2969 = n2968 ^ n2966 ;
  assign n2963 = n2648 & n2822 ;
  assign n2964 = n2732 & n2963 ;
  assign n2970 = n2969 ^ n2964 ;
  assign n2958 = n2158 & n2844 ;
  assign n2959 = n2958 ^ n2158 ;
  assign n2956 = n2158 & n2830 ;
  assign n2957 = n2956 ^ n2158 ;
  assign n2960 = n2959 ^ n2957 ;
  assign n2954 = n2158 & n2822 ;
  assign n2955 = n2732 & n2954 ;
  assign n2961 = n2960 ^ n2955 ;
  assign n2962 = n2961 ^ n2158 ;
  assign n2971 = n2970 ^ n2962 ;
  assign n2952 = n1992 & ~n2151 ;
  assign n2953 = n2952 ^ n2155 ;
  assign n2973 = n2971 ^ n2953 ;
  assign n2998 = n2670 & n2844 ;
  assign n2999 = n2998 ^ n2670 ;
  assign n2996 = n2670 & n2830 ;
  assign n2997 = n2996 ^ n2670 ;
  assign n3000 = n2999 ^ n2997 ;
  assign n2994 = n2670 & n2822 ;
  assign n2995 = n2732 & n2994 ;
  assign n3001 = n3000 ^ n2995 ;
  assign n2989 = n2654 & n2844 ;
  assign n2990 = n2989 ^ n2654 ;
  assign n2987 = n2654 & n2830 ;
  assign n2988 = n2987 ^ n2654 ;
  assign n2991 = n2990 ^ n2988 ;
  assign n2985 = n2654 & n2822 ;
  assign n2986 = n2732 & n2985 ;
  assign n2992 = n2991 ^ n2986 ;
  assign n2993 = n2992 ^ n2654 ;
  assign n3002 = n3001 ^ n2993 ;
  assign n2974 = n2019 & ~n2151 ;
  assign n2975 = n2974 ^ n2651 ;
  assign n3003 = n3002 ^ n2975 ;
  assign n3004 = n2973 & n3003 ;
  assign n3005 = n3004 ^ n2973 ;
  assign n3006 = n3005 ^ n3003 ;
  assign n3028 = n2697 & n2844 ;
  assign n3029 = n3028 ^ n2697 ;
  assign n3026 = n2697 & n2830 ;
  assign n3027 = n3026 ^ n2697 ;
  assign n3030 = n3029 ^ n3027 ;
  assign n3024 = n2697 & n2822 ;
  assign n3025 = n2732 & n3024 ;
  assign n3031 = n3030 ^ n3025 ;
  assign n3019 = n2681 & n2844 ;
  assign n3020 = n3019 ^ n2681 ;
  assign n3017 = n2681 & n2830 ;
  assign n3018 = n3017 ^ n2681 ;
  assign n3021 = n3020 ^ n3018 ;
  assign n3015 = n2681 & n2822 ;
  assign n3016 = n2732 & n3015 ;
  assign n3022 = n3021 ^ n3016 ;
  assign n3023 = n3022 ^ n2681 ;
  assign n3032 = n3031 ^ n3023 ;
  assign n3007 = n2053 & ~n2151 ;
  assign n3008 = n3007 ^ n2678 ;
  assign n3033 = n3032 ^ n3008 ;
  assign n3078 = n2703 & n2844 ;
  assign n3079 = n3078 ^ n2703 ;
  assign n3076 = n2703 & n2830 ;
  assign n3077 = n3076 ^ n2703 ;
  assign n3080 = n3079 ^ n3077 ;
  assign n3074 = n2703 & n2822 ;
  assign n3075 = n2732 & n3074 ;
  assign n3081 = n3080 ^ n3075 ;
  assign n3082 = n3081 ^ n2703 ;
  assign n3070 = n2725 & n2844 ;
  assign n3071 = n3070 ^ n2725 ;
  assign n3068 = n2725 & n2830 ;
  assign n3069 = n3068 ^ n2725 ;
  assign n3072 = n3071 ^ n3069 ;
  assign n3066 = n2725 & n2822 ;
  assign n3067 = n2732 & n3066 ;
  assign n3073 = n3072 ^ n3067 ;
  assign n3083 = n3082 ^ n3073 ;
  assign n3034 = n2081 & ~n2151 ;
  assign n3035 = n3034 ^ n2700 ;
  assign n3084 = n3083 ^ n3035 ;
  assign n3085 = n3033 & n3084 ;
  assign n3086 = n3085 ^ n3033 ;
  assign n3087 = n3086 ^ n3084 ;
  assign n3088 = n3006 & n3087 ;
  assign n3089 = n3088 ^ n3006 ;
  assign n3090 = n3089 ^ n3087 ;
  assign n3091 = n2951 & n3090 ;
  assign n3092 = n3091 ^ n2951 ;
  assign n3093 = n3092 ^ n3090 ;
  assign n3045 = n2703 & n3035 ;
  assign n3050 = n2844 & n3045 ;
  assign n3051 = n3050 ^ n3045 ;
  assign n3048 = n2830 & n3045 ;
  assign n3049 = n3048 ^ n3045 ;
  assign n3052 = n3051 ^ n3049 ;
  assign n3046 = n2822 & n3045 ;
  assign n3047 = n2732 & n3046 ;
  assign n3053 = n3052 ^ n3047 ;
  assign n3054 = n3053 ^ n3045 ;
  assign n3036 = n2725 & n3035 ;
  assign n3041 = n2844 & n3036 ;
  assign n3042 = n3041 ^ n3036 ;
  assign n3039 = n2830 & n3036 ;
  assign n3040 = n3039 ^ n3036 ;
  assign n3043 = n3042 ^ n3040 ;
  assign n3037 = n2822 & n3036 ;
  assign n3038 = n2732 & n3037 ;
  assign n3044 = n3043 ^ n3038 ;
  assign n3055 = n3054 ^ n3044 ;
  assign n3056 = n3055 ^ n3035 ;
  assign n3057 = n3033 & n3056 ;
  assign n3058 = n3057 ^ n3056 ;
  assign n2910 = n2732 & n2822 ;
  assign n2911 = n2910 ^ n2844 ;
  assign n2912 = n2911 ^ n2830 ;
  assign n3012 = ~n2697 & n3008 ;
  assign n3013 = n2912 & n3012 ;
  assign n3009 = ~n2681 & n3008 ;
  assign n3010 = n2912 & n3009 ;
  assign n3011 = n3010 ^ n3009 ;
  assign n3014 = n3013 ^ n3011 ;
  assign n3059 = n3058 ^ n3014 ;
  assign n3060 = n3006 & n3059 ;
  assign n3061 = n3060 ^ n3059 ;
  assign n2979 = ~n2670 & n2975 ;
  assign n2980 = n2912 & n2979 ;
  assign n2976 = ~n2654 & n2975 ;
  assign n2977 = n2912 & n2976 ;
  assign n2978 = n2977 ^ n2976 ;
  assign n2981 = n2980 ^ n2978 ;
  assign n2982 = n2973 & n2981 ;
  assign n2983 = n2982 ^ n2981 ;
  assign n2972 = n2953 & ~n2971 ;
  assign n2984 = n2983 ^ n2972 ;
  assign n3062 = n3061 ^ n2984 ;
  assign n3063 = n2951 & n3062 ;
  assign n3064 = n3063 ^ n3062 ;
  assign n2918 = ~n2817 & n2914 ;
  assign n2919 = n2912 & n2918 ;
  assign n2915 = ~n2801 & n2914 ;
  assign n2916 = n2912 & n2915 ;
  assign n2917 = n2916 ^ n2915 ;
  assign n2920 = n2919 ^ n2917 ;
  assign n2921 = n2909 & n2920 ;
  assign n2922 = n2921 ^ n2920 ;
  assign n2908 = n2889 & ~n2907 ;
  assign n2923 = n2922 ^ n2908 ;
  assign n2924 = n2887 & n2923 ;
  assign n2925 = n2924 ^ n2923 ;
  assign n2881 = n2862 & ~n2880 ;
  assign n2882 = ~n2860 & n2881 ;
  assign n2859 = n2154 & ~n2858 ;
  assign n2883 = n2882 ^ n2859 ;
  assign n2926 = n2925 ^ n2883 ;
  assign n3065 = n3064 ^ n2926 ;
  assign n3094 = n3093 ^ n3065 ;
  assign n3098 = n2858 & n3094 ;
  assign n3099 = n3098 ^ n2858 ;
  assign n3095 = n2154 & n3094 ;
  assign n3096 = n3095 ^ n2154 ;
  assign n3097 = n3096 ^ n2154 ;
  assign n3100 = n3099 ^ n3097 ;
  assign n3104 = n2880 & n3094 ;
  assign n3105 = n3104 ^ n2880 ;
  assign n3101 = n2862 & n3094 ;
  assign n3102 = n3101 ^ n2862 ;
  assign n3103 = n3102 ^ n2862 ;
  assign n3106 = n3105 ^ n3103 ;
  assign n3110 = n2907 & n3094 ;
  assign n3111 = n3110 ^ n2907 ;
  assign n3107 = n2889 & n3094 ;
  assign n3108 = n3107 ^ n2889 ;
  assign n3109 = n3108 ^ n2889 ;
  assign n3112 = n3111 ^ n3109 ;
  assign n3116 = n2944 & n3094 ;
  assign n3117 = n3116 ^ n2944 ;
  assign n3113 = n2914 & n3094 ;
  assign n3114 = n3113 ^ n2914 ;
  assign n3115 = n3114 ^ n2914 ;
  assign n3118 = n3117 ^ n3115 ;
  assign n3122 = n2971 & n3094 ;
  assign n3123 = n3122 ^ n2971 ;
  assign n3119 = n2953 & n3094 ;
  assign n3120 = n3119 ^ n2953 ;
  assign n3121 = n3120 ^ n2953 ;
  assign n3124 = n3123 ^ n3121 ;
  assign n3128 = n3002 & n3094 ;
  assign n3129 = n3128 ^ n3002 ;
  assign n3125 = n2975 & n3094 ;
  assign n3126 = n3125 ^ n2975 ;
  assign n3127 = n3126 ^ n2975 ;
  assign n3130 = n3129 ^ n3127 ;
  assign n3134 = n3032 & n3094 ;
  assign n3135 = n3134 ^ n3032 ;
  assign n3131 = n3008 & n3094 ;
  assign n3132 = n3131 ^ n3008 ;
  assign n3133 = n3132 ^ n3008 ;
  assign n3136 = n3135 ^ n3133 ;
  assign n3140 = n3083 & n3094 ;
  assign n3141 = n3140 ^ n3083 ;
  assign n3137 = n3035 & n3094 ;
  assign n3138 = n3137 ^ n3035 ;
  assign n3139 = n3138 ^ n3035 ;
  assign n3142 = n3141 ^ n3139 ;
  assign n3143 = n3099 ^ n2858 ;
  assign n3144 = n3143 ^ n3096 ;
  assign n3145 = n3105 ^ n2880 ;
  assign n3146 = n3145 ^ n3102 ;
  assign n3147 = n3111 ^ n2907 ;
  assign n3148 = n3147 ^ n3108 ;
  assign n3149 = n3117 ^ n2944 ;
  assign n3150 = n3149 ^ n3114 ;
  assign n3151 = n3123 ^ n2971 ;
  assign n3152 = n3151 ^ n3120 ;
  assign n3153 = n3129 ^ n3002 ;
  assign n3154 = n3153 ^ n3126 ;
  assign n3155 = n3135 ^ n3032 ;
  assign n3156 = n3155 ^ n3132 ;
  assign n3157 = n3141 ^ n3083 ;
  assign n3158 = n3157 ^ n3138 ;
  assign n3159 = n2751 & ~n2912 ;
  assign n3160 = n3159 ^ n2848 ;
  assign n3161 = n2772 & ~n2912 ;
  assign n3162 = n3161 ^ n2870 ;
  assign n3163 = n2796 & ~n2912 ;
  assign n3164 = n3163 ^ n2897 ;
  assign n3165 = n2817 & ~n2912 ;
  assign n3166 = n3165 ^ n2934 ;
  assign n3167 = n2648 & ~n2912 ;
  assign n3168 = n3167 ^ n2961 ;
  assign n3169 = n2670 & ~n2912 ;
  assign n3170 = n3169 ^ n2992 ;
  assign n3171 = n2697 & ~n2912 ;
  assign n3172 = n3171 ^ n3022 ;
  assign n3173 = n2725 & ~n2912 ;
  assign n3174 = n3173 ^ n3081 ;
  assign n3175 = n2494 & ~n2611 ;
  assign n3176 = n3175 ^ n2636 ;
  assign n3177 = n3176 ^ n2621 ;
  assign n3179 = n2496 & n3177 ;
  assign n3178 = n2520 & ~n3177 ;
  assign n3180 = n3179 ^ n3178 ;
  assign n3182 = n2523 & n3177 ;
  assign n3181 = n2547 & ~n3177 ;
  assign n3183 = n3182 ^ n3181 ;
  assign n3185 = n2553 & n3177 ;
  assign n3184 = n2577 & ~n3177 ;
  assign n3186 = n3185 ^ n3184 ;
  assign n3188 = n2580 & n3177 ;
  assign n3187 = n2604 & ~n3177 ;
  assign n3189 = n3188 ^ n3187 ;
  assign n3191 = n2160 & n3177 ;
  assign n3190 = n2392 & ~n3177 ;
  assign n3192 = n3191 ^ n3190 ;
  assign n3194 = n2396 & n3177 ;
  assign n3193 = n2420 & ~n3177 ;
  assign n3195 = n3194 ^ n3193 ;
  assign n3197 = n2431 & n3177 ;
  assign n3196 = n2455 & ~n3177 ;
  assign n3198 = n3197 ^ n3196 ;
  assign n3199 = n2486 & ~n3177 ;
  assign n3200 = n3199 ^ n2713 ;
  assign n3202 = n2328 & n2374 ;
  assign n3203 = n3202 ^ n2374 ;
  assign n3204 = n3203 ^ n2367 ;
  assign n3201 = n2311 & ~n2348 ;
  assign n3205 = n3204 ^ n3201 ;
  assign n3206 = n3205 ^ n2361 ;
  assign n3207 = n2317 & n3206 ;
  assign n3208 = n3207 ^ n2507 ;
  assign n3209 = n2322 & n3206 ;
  assign n3210 = n3209 ^ n2534 ;
  assign n3211 = n2332 & n3206 ;
  assign n3212 = n3211 ^ n2564 ;
  assign n3213 = n2341 & n3206 ;
  assign n3214 = n3213 ^ n2591 ;
  assign n3215 = n2271 & n3206 ;
  assign n3216 = n3215 ^ n2379 ;
  assign n3217 = n2279 & n3206 ;
  assign n3218 = n3217 ^ n2407 ;
  assign n3219 = n2294 & n3206 ;
  assign n3220 = n3219 ^ n2442 ;
  assign n3221 = n2303 & n3206 ;
  assign n3222 = n3221 ^ n2472 ;
  assign n3223 = x40 & n2267 ;
  assign n3224 = n3223 ^ n2314 ;
  assign n3225 = x41 & n2267 ;
  assign n3226 = n3225 ^ n2319 ;
  assign n3227 = x42 & n2267 ;
  assign n3228 = n3227 ^ n2329 ;
  assign n3229 = x43 & n2267 ;
  assign n3230 = n3229 ^ n2338 ;
  assign n3231 = x44 & n2267 ;
  assign n3232 = n3231 ^ n2268 ;
  assign n3233 = x45 & n2267 ;
  assign n3234 = n3233 ^ n2276 ;
  assign n3235 = x46 & n2267 ;
  assign n3236 = n3235 ^ n2291 ;
  assign n3237 = x47 & n2267 ;
  assign n3238 = n3237 ^ n2300 ;
  assign y0 = n3100 ;
  assign y1 = n3106 ;
  assign y2 = n3112 ;
  assign y3 = n3118 ;
  assign y4 = n3124 ;
  assign y5 = n3130 ;
  assign y6 = n3136 ;
  assign y7 = n3142 ;
  assign y8 = n3144 ;
  assign y9 = n3146 ;
  assign y10 = n3148 ;
  assign y11 = n3150 ;
  assign y12 = n3152 ;
  assign y13 = n3154 ;
  assign y14 = n3156 ;
  assign y15 = n3158 ;
  assign y16 = n3160 ;
  assign y17 = n3162 ;
  assign y18 = n3164 ;
  assign y19 = n3166 ;
  assign y20 = n3168 ;
  assign y21 = n3170 ;
  assign y22 = n3172 ;
  assign y23 = n3174 ;
  assign y24 = n3180 ;
  assign y25 = n3183 ;
  assign y26 = n3186 ;
  assign y27 = n3189 ;
  assign y28 = n3192 ;
  assign y29 = n3195 ;
  assign y30 = n3198 ;
  assign y31 = n3200 ;
  assign y32 = n3208 ;
  assign y33 = n3210 ;
  assign y34 = n3212 ;
  assign y35 = n3214 ;
  assign y36 = n3216 ;
  assign y37 = n3218 ;
  assign y38 = n3220 ;
  assign y39 = n3222 ;
  assign y40 = n3224 ;
  assign y41 = n3226 ;
  assign y42 = n3228 ;
  assign y43 = n3230 ;
  assign y44 = n3232 ;
  assign y45 = n3234 ;
  assign y46 = n3236 ;
  assign y47 = n3238 ;
endmodule
