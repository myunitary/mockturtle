module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 ;
  assign n129 = ~x79 & ~x95 ;
  assign n130 = ~x111 & ~x127 ;
  assign n131 = n129 & n130 ;
  assign n132 = ~x15 & ~x31 ;
  assign n133 = ~x47 & ~x63 ;
  assign n134 = n132 & n133 ;
  assign n135 = n131 & ~n134 ;
  assign n136 = ~x15 & x31 ;
  assign n137 = x15 & ~x31 ;
  assign n138 = ~x14 & x30 ;
  assign n139 = x14 & ~x30 ;
  assign n140 = ~x13 & x29 ;
  assign n141 = x13 & ~x29 ;
  assign n142 = ~x12 & x28 ;
  assign n143 = x12 & ~x28 ;
  assign n144 = ~x11 & x27 ;
  assign n145 = x11 & ~x27 ;
  assign n146 = ~x10 & x26 ;
  assign n147 = x10 & ~x26 ;
  assign n148 = ~x9 & x25 ;
  assign n149 = x9 & ~x25 ;
  assign n150 = ~x8 & x24 ;
  assign n151 = x8 & ~x24 ;
  assign n152 = ~x7 & x23 ;
  assign n153 = x7 & ~x23 ;
  assign n154 = ~x6 & x22 ;
  assign n155 = x6 & ~x22 ;
  assign n156 = ~x5 & x21 ;
  assign n157 = x5 & ~x21 ;
  assign n158 = ~x4 & x20 ;
  assign n159 = x4 & ~x20 ;
  assign n160 = ~x3 & x19 ;
  assign n161 = x3 & ~x19 ;
  assign n162 = ~x2 & x18 ;
  assign n163 = x2 & ~x18 ;
  assign n164 = ~x1 & x17 ;
  assign n165 = x1 & ~x17 ;
  assign n166 = x0 & ~x16 ;
  assign n167 = ~n165 & ~n166 ;
  assign n168 = ~n164 & ~n167 ;
  assign n169 = ~n163 & ~n168 ;
  assign n170 = ~n162 & ~n169 ;
  assign n171 = ~n161 & ~n170 ;
  assign n172 = ~n160 & ~n171 ;
  assign n173 = ~n159 & ~n172 ;
  assign n174 = ~n158 & ~n173 ;
  assign n175 = ~n157 & ~n174 ;
  assign n176 = ~n156 & ~n175 ;
  assign n177 = ~n155 & ~n176 ;
  assign n178 = ~n154 & ~n177 ;
  assign n179 = ~n153 & ~n178 ;
  assign n180 = ~n152 & ~n179 ;
  assign n181 = ~n151 & ~n180 ;
  assign n182 = ~n150 & ~n181 ;
  assign n183 = ~n149 & ~n182 ;
  assign n184 = ~n148 & ~n183 ;
  assign n185 = ~n147 & ~n184 ;
  assign n186 = ~n146 & ~n185 ;
  assign n187 = ~n145 & ~n186 ;
  assign n188 = ~n144 & ~n187 ;
  assign n189 = ~n143 & ~n188 ;
  assign n190 = ~n142 & ~n189 ;
  assign n191 = ~n141 & ~n190 ;
  assign n192 = ~n140 & ~n191 ;
  assign n193 = ~n139 & ~n192 ;
  assign n194 = ~n138 & ~n193 ;
  assign n195 = ~n137 & ~n194 ;
  assign n196 = ~n136 & ~n195 ;
  assign n197 = x17 & ~n196 ;
  assign n198 = x1 & n196 ;
  assign n199 = ~n197 & ~n198 ;
  assign n200 = n132 & ~n133 ;
  assign n201 = ~n132 & n133 ;
  assign n202 = ~x47 & x63 ;
  assign n203 = x47 & ~x63 ;
  assign n204 = ~x46 & x62 ;
  assign n205 = x46 & ~x62 ;
  assign n206 = ~x45 & x61 ;
  assign n207 = x45 & ~x61 ;
  assign n208 = ~x44 & x60 ;
  assign n209 = x44 & ~x60 ;
  assign n210 = ~x43 & x59 ;
  assign n211 = x43 & ~x59 ;
  assign n212 = ~x42 & x58 ;
  assign n213 = x42 & ~x58 ;
  assign n214 = ~x41 & x57 ;
  assign n215 = x41 & ~x57 ;
  assign n216 = ~x40 & x56 ;
  assign n217 = x40 & ~x56 ;
  assign n218 = ~x39 & x55 ;
  assign n219 = x39 & ~x55 ;
  assign n220 = ~x38 & x54 ;
  assign n221 = x38 & ~x54 ;
  assign n222 = ~x37 & x53 ;
  assign n223 = x37 & ~x53 ;
  assign n224 = ~x36 & x52 ;
  assign n225 = x36 & ~x52 ;
  assign n226 = ~x35 & x51 ;
  assign n227 = x35 & ~x51 ;
  assign n228 = ~x34 & x50 ;
  assign n229 = x34 & ~x50 ;
  assign n230 = ~x33 & x49 ;
  assign n231 = x33 & ~x49 ;
  assign n232 = x32 & ~x48 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = ~n230 & ~n233 ;
  assign n235 = ~n229 & ~n234 ;
  assign n236 = ~n228 & ~n235 ;
  assign n237 = ~n227 & ~n236 ;
  assign n238 = ~n226 & ~n237 ;
  assign n239 = ~n225 & ~n238 ;
  assign n240 = ~n224 & ~n239 ;
  assign n241 = ~n223 & ~n240 ;
  assign n242 = ~n222 & ~n241 ;
  assign n243 = ~n221 & ~n242 ;
  assign n244 = ~n220 & ~n243 ;
  assign n245 = ~n219 & ~n244 ;
  assign n246 = ~n218 & ~n245 ;
  assign n247 = ~n217 & ~n246 ;
  assign n248 = ~n216 & ~n247 ;
  assign n249 = ~n215 & ~n248 ;
  assign n250 = ~n214 & ~n249 ;
  assign n251 = ~n213 & ~n250 ;
  assign n252 = ~n212 & ~n251 ;
  assign n253 = ~n211 & ~n252 ;
  assign n254 = ~n210 & ~n253 ;
  assign n255 = ~n209 & ~n254 ;
  assign n256 = ~n208 & ~n255 ;
  assign n257 = ~n207 & ~n256 ;
  assign n258 = ~n206 & ~n257 ;
  assign n259 = ~n205 & ~n258 ;
  assign n260 = ~n204 & ~n259 ;
  assign n261 = ~n203 & ~n260 ;
  assign n262 = ~n202 & ~n261 ;
  assign n263 = x62 & ~n262 ;
  assign n264 = x46 & n262 ;
  assign n265 = ~n263 & ~n264 ;
  assign n266 = x30 & ~n196 ;
  assign n267 = x14 & n196 ;
  assign n268 = ~n266 & ~n267 ;
  assign n269 = ~n265 & n268 ;
  assign n270 = x49 & ~n262 ;
  assign n271 = x33 & n262 ;
  assign n272 = ~n270 & ~n271 ;
  assign n273 = n199 & ~n272 ;
  assign n274 = x48 & ~n262 ;
  assign n275 = x32 & n262 ;
  assign n276 = ~n274 & ~n275 ;
  assign n277 = x16 & ~n196 ;
  assign n278 = x0 & n196 ;
  assign n279 = ~n277 & ~n278 ;
  assign n280 = n276 & ~n279 ;
  assign n281 = ~n273 & n280 ;
  assign n282 = x50 & ~n262 ;
  assign n283 = x34 & n262 ;
  assign n284 = ~n282 & ~n283 ;
  assign n285 = x18 & ~n196 ;
  assign n286 = x2 & n196 ;
  assign n287 = ~n285 & ~n286 ;
  assign n288 = n284 & ~n287 ;
  assign n289 = ~n199 & n272 ;
  assign n290 = ~n288 & ~n289 ;
  assign n291 = ~n281 & n290 ;
  assign n292 = x19 & ~n196 ;
  assign n293 = x3 & n196 ;
  assign n294 = ~n292 & ~n293 ;
  assign n295 = x51 & ~n262 ;
  assign n296 = x35 & n262 ;
  assign n297 = ~n295 & ~n296 ;
  assign n298 = n294 & ~n297 ;
  assign n299 = ~n284 & n287 ;
  assign n300 = ~n298 & ~n299 ;
  assign n301 = ~n291 & n300 ;
  assign n302 = x52 & ~n262 ;
  assign n303 = x36 & n262 ;
  assign n304 = ~n302 & ~n303 ;
  assign n305 = x20 & ~n196 ;
  assign n306 = x4 & n196 ;
  assign n307 = ~n305 & ~n306 ;
  assign n308 = n304 & ~n307 ;
  assign n309 = ~n294 & n297 ;
  assign n310 = ~n308 & ~n309 ;
  assign n311 = ~n301 & n310 ;
  assign n312 = x53 & ~n262 ;
  assign n313 = x37 & n262 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = x21 & ~n196 ;
  assign n316 = x5 & n196 ;
  assign n317 = ~n315 & ~n316 ;
  assign n318 = ~n314 & n317 ;
  assign n319 = ~n304 & n307 ;
  assign n320 = ~n318 & ~n319 ;
  assign n321 = ~n311 & n320 ;
  assign n322 = x22 & ~n196 ;
  assign n323 = x6 & n196 ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = x54 & ~n262 ;
  assign n326 = x38 & n262 ;
  assign n327 = ~n325 & ~n326 ;
  assign n328 = ~n324 & n327 ;
  assign n329 = n314 & ~n317 ;
  assign n330 = ~n328 & ~n329 ;
  assign n331 = ~n321 & n330 ;
  assign n332 = x23 & ~n196 ;
  assign n333 = x7 & n196 ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = x55 & ~n262 ;
  assign n336 = x39 & n262 ;
  assign n337 = ~n335 & ~n336 ;
  assign n338 = n334 & ~n337 ;
  assign n339 = n324 & ~n327 ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = ~n331 & n340 ;
  assign n342 = ~n334 & n337 ;
  assign n343 = x24 & ~n196 ;
  assign n344 = x8 & n196 ;
  assign n345 = ~n343 & ~n344 ;
  assign n346 = x56 & ~n262 ;
  assign n347 = x40 & n262 ;
  assign n348 = ~n346 & ~n347 ;
  assign n349 = ~n345 & n348 ;
  assign n350 = ~n342 & ~n349 ;
  assign n351 = ~n341 & n350 ;
  assign n352 = n345 & ~n348 ;
  assign n353 = x57 & ~n262 ;
  assign n354 = x41 & n262 ;
  assign n355 = ~n353 & ~n354 ;
  assign n356 = x25 & ~n196 ;
  assign n357 = x9 & n196 ;
  assign n358 = ~n356 & ~n357 ;
  assign n359 = ~n355 & n358 ;
  assign n360 = ~n352 & ~n359 ;
  assign n361 = ~n351 & n360 ;
  assign n362 = n355 & ~n358 ;
  assign n363 = x26 & ~n196 ;
  assign n364 = x10 & n196 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = x58 & ~n262 ;
  assign n367 = x42 & n262 ;
  assign n368 = ~n366 & ~n367 ;
  assign n369 = ~n365 & n368 ;
  assign n370 = ~n362 & ~n369 ;
  assign n371 = ~n361 & n370 ;
  assign n372 = x27 & ~n196 ;
  assign n373 = x11 & n196 ;
  assign n374 = ~n372 & ~n373 ;
  assign n375 = x59 & ~n262 ;
  assign n376 = x43 & n262 ;
  assign n377 = ~n375 & ~n376 ;
  assign n378 = n374 & ~n377 ;
  assign n379 = n365 & ~n368 ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = ~n371 & n380 ;
  assign n382 = x60 & ~n262 ;
  assign n383 = x44 & n262 ;
  assign n384 = ~n382 & ~n383 ;
  assign n385 = x28 & ~n196 ;
  assign n386 = x12 & n196 ;
  assign n387 = ~n385 & ~n386 ;
  assign n388 = n384 & ~n387 ;
  assign n389 = ~n374 & n377 ;
  assign n390 = ~n388 & ~n389 ;
  assign n391 = ~n381 & n390 ;
  assign n392 = ~n384 & n387 ;
  assign n393 = x29 & ~n196 ;
  assign n394 = x13 & n196 ;
  assign n395 = ~n393 & ~n394 ;
  assign n396 = x61 & ~n262 ;
  assign n397 = x45 & n262 ;
  assign n398 = ~n396 & ~n397 ;
  assign n399 = n395 & ~n398 ;
  assign n400 = ~n392 & ~n399 ;
  assign n401 = ~n391 & n400 ;
  assign n402 = n265 & ~n268 ;
  assign n403 = ~n395 & n398 ;
  assign n404 = ~n402 & ~n403 ;
  assign n405 = ~n401 & n404 ;
  assign n406 = ~n269 & ~n405 ;
  assign n407 = ~n201 & ~n406 ;
  assign n408 = ~n200 & ~n407 ;
  assign n409 = ~n199 & n408 ;
  assign n410 = ~n272 & ~n408 ;
  assign n411 = ~n409 & ~n410 ;
  assign n412 = ~x79 & x95 ;
  assign n413 = x79 & ~x95 ;
  assign n414 = ~x78 & x94 ;
  assign n415 = x78 & ~x94 ;
  assign n416 = ~x77 & x93 ;
  assign n417 = x77 & ~x93 ;
  assign n418 = ~x76 & x92 ;
  assign n419 = x76 & ~x92 ;
  assign n420 = ~x75 & x91 ;
  assign n421 = x75 & ~x91 ;
  assign n422 = ~x74 & x90 ;
  assign n423 = x74 & ~x90 ;
  assign n424 = ~x73 & x89 ;
  assign n425 = x73 & ~x89 ;
  assign n426 = ~x72 & x88 ;
  assign n427 = x72 & ~x88 ;
  assign n428 = ~x71 & x87 ;
  assign n429 = x71 & ~x87 ;
  assign n430 = ~x70 & x86 ;
  assign n431 = x70 & ~x86 ;
  assign n432 = ~x69 & x85 ;
  assign n433 = x69 & ~x85 ;
  assign n434 = ~x68 & x84 ;
  assign n435 = x68 & ~x84 ;
  assign n436 = ~x67 & x83 ;
  assign n437 = x67 & ~x83 ;
  assign n438 = ~x66 & x82 ;
  assign n439 = x66 & ~x82 ;
  assign n440 = ~x65 & x81 ;
  assign n441 = x65 & ~x81 ;
  assign n442 = x64 & ~x80 ;
  assign n443 = ~n441 & ~n442 ;
  assign n444 = ~n440 & ~n443 ;
  assign n445 = ~n439 & ~n444 ;
  assign n446 = ~n438 & ~n445 ;
  assign n447 = ~n437 & ~n446 ;
  assign n448 = ~n436 & ~n447 ;
  assign n449 = ~n435 & ~n448 ;
  assign n450 = ~n434 & ~n449 ;
  assign n451 = ~n433 & ~n450 ;
  assign n452 = ~n432 & ~n451 ;
  assign n453 = ~n431 & ~n452 ;
  assign n454 = ~n430 & ~n453 ;
  assign n455 = ~n429 & ~n454 ;
  assign n456 = ~n428 & ~n455 ;
  assign n457 = ~n427 & ~n456 ;
  assign n458 = ~n426 & ~n457 ;
  assign n459 = ~n425 & ~n458 ;
  assign n460 = ~n424 & ~n459 ;
  assign n461 = ~n423 & ~n460 ;
  assign n462 = ~n422 & ~n461 ;
  assign n463 = ~n421 & ~n462 ;
  assign n464 = ~n420 & ~n463 ;
  assign n465 = ~n419 & ~n464 ;
  assign n466 = ~n418 & ~n465 ;
  assign n467 = ~n417 & ~n466 ;
  assign n468 = ~n416 & ~n467 ;
  assign n469 = ~n415 & ~n468 ;
  assign n470 = ~n414 & ~n469 ;
  assign n471 = ~n413 & ~n470 ;
  assign n472 = ~n412 & ~n471 ;
  assign n473 = x81 & ~n472 ;
  assign n474 = x65 & n472 ;
  assign n475 = ~n473 & ~n474 ;
  assign n476 = n129 & ~n130 ;
  assign n477 = ~n129 & n130 ;
  assign n478 = ~x111 & x127 ;
  assign n479 = x111 & ~x127 ;
  assign n480 = ~x110 & x126 ;
  assign n481 = x110 & ~x126 ;
  assign n482 = ~x109 & x125 ;
  assign n483 = x109 & ~x125 ;
  assign n484 = ~x108 & x124 ;
  assign n485 = x108 & ~x124 ;
  assign n486 = ~x107 & x123 ;
  assign n487 = x107 & ~x123 ;
  assign n488 = ~x106 & x122 ;
  assign n489 = x106 & ~x122 ;
  assign n490 = ~x105 & x121 ;
  assign n491 = x105 & ~x121 ;
  assign n492 = ~x104 & x120 ;
  assign n493 = x104 & ~x120 ;
  assign n494 = ~x103 & x119 ;
  assign n495 = x103 & ~x119 ;
  assign n496 = ~x102 & x118 ;
  assign n497 = x102 & ~x118 ;
  assign n498 = ~x101 & x117 ;
  assign n499 = x101 & ~x117 ;
  assign n500 = ~x100 & x116 ;
  assign n501 = x100 & ~x116 ;
  assign n502 = ~x99 & x115 ;
  assign n503 = x99 & ~x115 ;
  assign n504 = ~x98 & x114 ;
  assign n505 = x98 & ~x114 ;
  assign n506 = ~x97 & x113 ;
  assign n507 = x97 & ~x113 ;
  assign n508 = x96 & ~x112 ;
  assign n509 = ~n507 & ~n508 ;
  assign n510 = ~n506 & ~n509 ;
  assign n511 = ~n505 & ~n510 ;
  assign n512 = ~n504 & ~n511 ;
  assign n513 = ~n503 & ~n512 ;
  assign n514 = ~n502 & ~n513 ;
  assign n515 = ~n501 & ~n514 ;
  assign n516 = ~n500 & ~n515 ;
  assign n517 = ~n499 & ~n516 ;
  assign n518 = ~n498 & ~n517 ;
  assign n519 = ~n497 & ~n518 ;
  assign n520 = ~n496 & ~n519 ;
  assign n521 = ~n495 & ~n520 ;
  assign n522 = ~n494 & ~n521 ;
  assign n523 = ~n493 & ~n522 ;
  assign n524 = ~n492 & ~n523 ;
  assign n525 = ~n491 & ~n524 ;
  assign n526 = ~n490 & ~n525 ;
  assign n527 = ~n489 & ~n526 ;
  assign n528 = ~n488 & ~n527 ;
  assign n529 = ~n487 & ~n528 ;
  assign n530 = ~n486 & ~n529 ;
  assign n531 = ~n485 & ~n530 ;
  assign n532 = ~n484 & ~n531 ;
  assign n533 = ~n483 & ~n532 ;
  assign n534 = ~n482 & ~n533 ;
  assign n535 = ~n481 & ~n534 ;
  assign n536 = ~n480 & ~n535 ;
  assign n537 = ~n479 & ~n536 ;
  assign n538 = ~n478 & ~n537 ;
  assign n539 = x113 & ~n538 ;
  assign n540 = x97 & n538 ;
  assign n541 = ~n539 & ~n540 ;
  assign n542 = n475 & ~n541 ;
  assign n543 = x112 & ~n538 ;
  assign n544 = x96 & n538 ;
  assign n545 = ~n543 & ~n544 ;
  assign n546 = x80 & ~n472 ;
  assign n547 = x64 & n472 ;
  assign n548 = ~n546 & ~n547 ;
  assign n549 = n545 & ~n548 ;
  assign n550 = ~n542 & n549 ;
  assign n551 = x114 & ~n538 ;
  assign n552 = x98 & n538 ;
  assign n553 = ~n551 & ~n552 ;
  assign n554 = x82 & ~n472 ;
  assign n555 = x66 & n472 ;
  assign n556 = ~n554 & ~n555 ;
  assign n557 = n553 & ~n556 ;
  assign n558 = ~n475 & n541 ;
  assign n559 = ~n557 & ~n558 ;
  assign n560 = ~n550 & n559 ;
  assign n561 = ~n553 & n556 ;
  assign n562 = x115 & ~n538 ;
  assign n563 = x99 & n538 ;
  assign n564 = ~n562 & ~n563 ;
  assign n565 = x83 & ~n472 ;
  assign n566 = x67 & n472 ;
  assign n567 = ~n565 & ~n566 ;
  assign n568 = ~n564 & n567 ;
  assign n569 = ~n561 & ~n568 ;
  assign n570 = ~n560 & n569 ;
  assign n571 = x84 & ~n472 ;
  assign n572 = x68 & n472 ;
  assign n573 = ~n571 & ~n572 ;
  assign n574 = x116 & ~n538 ;
  assign n575 = x100 & n538 ;
  assign n576 = ~n574 & ~n575 ;
  assign n577 = ~n573 & n576 ;
  assign n578 = n564 & ~n567 ;
  assign n579 = ~n577 & ~n578 ;
  assign n580 = ~n570 & n579 ;
  assign n581 = x117 & ~n538 ;
  assign n582 = x101 & n538 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = x85 & ~n472 ;
  assign n585 = x69 & n472 ;
  assign n586 = ~n584 & ~n585 ;
  assign n587 = ~n583 & n586 ;
  assign n588 = n573 & ~n576 ;
  assign n589 = ~n587 & ~n588 ;
  assign n590 = ~n580 & n589 ;
  assign n591 = x118 & ~n538 ;
  assign n592 = x102 & n538 ;
  assign n593 = ~n591 & ~n592 ;
  assign n594 = x86 & ~n472 ;
  assign n595 = x70 & n472 ;
  assign n596 = ~n594 & ~n595 ;
  assign n597 = n593 & ~n596 ;
  assign n598 = n583 & ~n586 ;
  assign n599 = ~n597 & ~n598 ;
  assign n600 = ~n590 & n599 ;
  assign n601 = ~n593 & n596 ;
  assign n602 = x87 & ~n472 ;
  assign n603 = x71 & n472 ;
  assign n604 = ~n602 & ~n603 ;
  assign n605 = x119 & ~n538 ;
  assign n606 = x103 & n538 ;
  assign n607 = ~n605 & ~n606 ;
  assign n608 = n604 & ~n607 ;
  assign n609 = ~n601 & ~n608 ;
  assign n610 = ~n600 & n609 ;
  assign n611 = ~n604 & n607 ;
  assign n612 = x120 & ~n538 ;
  assign n613 = x104 & n538 ;
  assign n614 = ~n612 & ~n613 ;
  assign n615 = x88 & ~n472 ;
  assign n616 = x72 & n472 ;
  assign n617 = ~n615 & ~n616 ;
  assign n618 = n614 & ~n617 ;
  assign n619 = ~n611 & ~n618 ;
  assign n620 = ~n610 & n619 ;
  assign n621 = ~n614 & n617 ;
  assign n622 = x121 & ~n538 ;
  assign n623 = x105 & n538 ;
  assign n624 = ~n622 & ~n623 ;
  assign n625 = x89 & ~n472 ;
  assign n626 = x73 & n472 ;
  assign n627 = ~n625 & ~n626 ;
  assign n628 = ~n624 & n627 ;
  assign n629 = ~n621 & ~n628 ;
  assign n630 = ~n620 & n629 ;
  assign n631 = n624 & ~n627 ;
  assign n632 = x90 & ~n472 ;
  assign n633 = x74 & n472 ;
  assign n634 = ~n632 & ~n633 ;
  assign n635 = x122 & ~n538 ;
  assign n636 = x106 & n538 ;
  assign n637 = ~n635 & ~n636 ;
  assign n638 = ~n634 & n637 ;
  assign n639 = ~n631 & ~n638 ;
  assign n640 = ~n630 & n639 ;
  assign n641 = x123 & ~n538 ;
  assign n642 = x107 & n538 ;
  assign n643 = ~n641 & ~n642 ;
  assign n644 = x91 & ~n472 ;
  assign n645 = x75 & n472 ;
  assign n646 = ~n644 & ~n645 ;
  assign n647 = ~n643 & n646 ;
  assign n648 = n634 & ~n637 ;
  assign n649 = ~n647 & ~n648 ;
  assign n650 = ~n640 & n649 ;
  assign n651 = x92 & ~n472 ;
  assign n652 = x76 & n472 ;
  assign n653 = ~n651 & ~n652 ;
  assign n654 = x124 & ~n538 ;
  assign n655 = x108 & n538 ;
  assign n656 = ~n654 & ~n655 ;
  assign n657 = ~n653 & n656 ;
  assign n658 = n643 & ~n646 ;
  assign n659 = ~n657 & ~n658 ;
  assign n660 = ~n650 & n659 ;
  assign n661 = n653 & ~n656 ;
  assign n662 = x93 & ~n472 ;
  assign n663 = x77 & n472 ;
  assign n664 = ~n662 & ~n663 ;
  assign n665 = x125 & ~n538 ;
  assign n666 = x109 & n538 ;
  assign n667 = ~n665 & ~n666 ;
  assign n668 = n664 & ~n667 ;
  assign n669 = ~n661 & ~n668 ;
  assign n670 = ~n660 & n669 ;
  assign n671 = ~n664 & n667 ;
  assign n672 = x94 & ~n472 ;
  assign n673 = x78 & n472 ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = x126 & ~n538 ;
  assign n676 = x110 & n538 ;
  assign n677 = ~n675 & ~n676 ;
  assign n678 = ~n674 & n677 ;
  assign n679 = ~n671 & ~n678 ;
  assign n680 = ~n670 & n679 ;
  assign n681 = n674 & ~n677 ;
  assign n682 = ~n680 & ~n681 ;
  assign n683 = ~n477 & ~n682 ;
  assign n684 = ~n476 & ~n683 ;
  assign n685 = ~n475 & n684 ;
  assign n686 = ~n541 & ~n684 ;
  assign n687 = ~n685 & ~n686 ;
  assign n688 = n411 & ~n687 ;
  assign n689 = ~n548 & n684 ;
  assign n690 = ~n545 & ~n684 ;
  assign n691 = ~n689 & ~n690 ;
  assign n692 = ~n279 & n408 ;
  assign n693 = ~n276 & ~n408 ;
  assign n694 = ~n692 & ~n693 ;
  assign n695 = n691 & ~n694 ;
  assign n696 = ~n688 & n695 ;
  assign n697 = ~n556 & n684 ;
  assign n698 = ~n553 & ~n684 ;
  assign n699 = ~n697 & ~n698 ;
  assign n700 = ~n287 & n408 ;
  assign n701 = ~n284 & ~n408 ;
  assign n702 = ~n700 & ~n701 ;
  assign n703 = n699 & ~n702 ;
  assign n704 = ~n411 & n687 ;
  assign n705 = ~n703 & ~n704 ;
  assign n706 = ~n696 & n705 ;
  assign n707 = ~n699 & n702 ;
  assign n708 = ~n294 & n408 ;
  assign n709 = ~n297 & ~n408 ;
  assign n710 = ~n708 & ~n709 ;
  assign n711 = ~n567 & n684 ;
  assign n712 = ~n564 & ~n684 ;
  assign n713 = ~n711 & ~n712 ;
  assign n714 = n710 & ~n713 ;
  assign n715 = ~n707 & ~n714 ;
  assign n716 = ~n706 & n715 ;
  assign n717 = ~n573 & n684 ;
  assign n718 = ~n576 & ~n684 ;
  assign n719 = ~n717 & ~n718 ;
  assign n720 = ~n307 & n408 ;
  assign n721 = ~n304 & ~n408 ;
  assign n722 = ~n720 & ~n721 ;
  assign n723 = n719 & ~n722 ;
  assign n724 = ~n710 & n713 ;
  assign n725 = ~n723 & ~n724 ;
  assign n726 = ~n716 & n725 ;
  assign n727 = ~n317 & n408 ;
  assign n728 = ~n314 & ~n408 ;
  assign n729 = ~n727 & ~n728 ;
  assign n730 = ~n586 & n684 ;
  assign n731 = ~n583 & ~n684 ;
  assign n732 = ~n730 & ~n731 ;
  assign n733 = n729 & ~n732 ;
  assign n734 = ~n719 & n722 ;
  assign n735 = ~n733 & ~n734 ;
  assign n736 = ~n726 & n735 ;
  assign n737 = ~n324 & n408 ;
  assign n738 = ~n327 & ~n408 ;
  assign n739 = ~n737 & ~n738 ;
  assign n740 = ~n596 & n684 ;
  assign n741 = ~n593 & ~n684 ;
  assign n742 = ~n740 & ~n741 ;
  assign n743 = ~n739 & n742 ;
  assign n744 = ~n729 & n732 ;
  assign n745 = ~n743 & ~n744 ;
  assign n746 = ~n736 & n745 ;
  assign n747 = ~n334 & n408 ;
  assign n748 = ~n337 & ~n408 ;
  assign n749 = ~n747 & ~n748 ;
  assign n750 = ~n604 & n684 ;
  assign n751 = ~n607 & ~n684 ;
  assign n752 = ~n750 & ~n751 ;
  assign n753 = n749 & ~n752 ;
  assign n754 = n739 & ~n742 ;
  assign n755 = ~n753 & ~n754 ;
  assign n756 = ~n746 & n755 ;
  assign n757 = ~n345 & n408 ;
  assign n758 = ~n348 & ~n408 ;
  assign n759 = ~n757 & ~n758 ;
  assign n760 = ~n617 & n684 ;
  assign n761 = ~n614 & ~n684 ;
  assign n762 = ~n760 & ~n761 ;
  assign n763 = ~n759 & n762 ;
  assign n764 = ~n749 & n752 ;
  assign n765 = ~n763 & ~n764 ;
  assign n766 = ~n756 & n765 ;
  assign n767 = ~n358 & n408 ;
  assign n768 = ~n355 & ~n408 ;
  assign n769 = ~n767 & ~n768 ;
  assign n770 = ~n627 & n684 ;
  assign n771 = ~n624 & ~n684 ;
  assign n772 = ~n770 & ~n771 ;
  assign n773 = n769 & ~n772 ;
  assign n774 = n759 & ~n762 ;
  assign n775 = ~n773 & ~n774 ;
  assign n776 = ~n766 & n775 ;
  assign n777 = ~n634 & n684 ;
  assign n778 = ~n637 & ~n684 ;
  assign n779 = ~n777 & ~n778 ;
  assign n780 = ~n365 & n408 ;
  assign n781 = ~n368 & ~n408 ;
  assign n782 = ~n780 & ~n781 ;
  assign n783 = n779 & ~n782 ;
  assign n784 = ~n769 & n772 ;
  assign n785 = ~n783 & ~n784 ;
  assign n786 = ~n776 & n785 ;
  assign n787 = ~n779 & n782 ;
  assign n788 = ~n374 & n408 ;
  assign n789 = ~n377 & ~n408 ;
  assign n790 = ~n788 & ~n789 ;
  assign n791 = ~n646 & n684 ;
  assign n792 = ~n643 & ~n684 ;
  assign n793 = ~n791 & ~n792 ;
  assign n794 = n790 & ~n793 ;
  assign n795 = ~n787 & ~n794 ;
  assign n796 = ~n786 & n795 ;
  assign n797 = ~n790 & n793 ;
  assign n798 = ~n653 & n684 ;
  assign n799 = ~n656 & ~n684 ;
  assign n800 = ~n798 & ~n799 ;
  assign n801 = ~n387 & n408 ;
  assign n802 = ~n384 & ~n408 ;
  assign n803 = ~n801 & ~n802 ;
  assign n804 = n800 & ~n803 ;
  assign n805 = ~n797 & ~n804 ;
  assign n806 = ~n796 & n805 ;
  assign n807 = ~n800 & n803 ;
  assign n808 = ~n664 & n684 ;
  assign n809 = ~n667 & ~n684 ;
  assign n810 = ~n808 & ~n809 ;
  assign n811 = ~n395 & n408 ;
  assign n812 = ~n398 & ~n408 ;
  assign n813 = ~n811 & ~n812 ;
  assign n814 = ~n810 & n813 ;
  assign n815 = ~n807 & ~n814 ;
  assign n816 = ~n806 & n815 ;
  assign n817 = n810 & ~n813 ;
  assign n818 = ~n674 & n684 ;
  assign n819 = ~n677 & ~n684 ;
  assign n820 = ~n818 & ~n819 ;
  assign n821 = ~n268 & n408 ;
  assign n822 = ~n265 & ~n408 ;
  assign n823 = ~n821 & ~n822 ;
  assign n824 = n820 & ~n823 ;
  assign n825 = ~n817 & ~n824 ;
  assign n826 = ~n816 & n825 ;
  assign n827 = ~n131 & n134 ;
  assign n828 = ~n820 & n823 ;
  assign n829 = ~n827 & ~n828 ;
  assign n830 = ~n826 & n829 ;
  assign n831 = ~n135 & ~n830 ;
  assign n832 = ~n684 & n831 ;
  assign n833 = ~n408 & ~n831 ;
  assign n834 = ~n832 & ~n833 ;
  assign n835 = n472 & n834 ;
  assign n836 = n538 & ~n684 ;
  assign n837 = ~n835 & ~n836 ;
  assign n838 = n831 & ~n837 ;
  assign n839 = n196 & n834 ;
  assign n840 = n262 & ~n408 ;
  assign n841 = ~n839 & ~n840 ;
  assign n842 = ~n831 & ~n841 ;
  assign n843 = ~n838 & ~n842 ;
  assign n844 = ~n694 & ~n831 ;
  assign n845 = ~n691 & n831 ;
  assign n846 = ~n844 & ~n845 ;
  assign n847 = ~n411 & ~n831 ;
  assign n848 = ~n687 & n831 ;
  assign n849 = ~n847 & ~n848 ;
  assign n850 = ~n702 & ~n831 ;
  assign n851 = ~n699 & n831 ;
  assign n852 = ~n850 & ~n851 ;
  assign n853 = ~n713 & n831 ;
  assign n854 = ~n710 & ~n831 ;
  assign n855 = ~n853 & ~n854 ;
  assign n856 = ~n722 & ~n831 ;
  assign n857 = ~n719 & n831 ;
  assign n858 = ~n856 & ~n857 ;
  assign n859 = ~n729 & ~n831 ;
  assign n860 = ~n732 & n831 ;
  assign n861 = ~n859 & ~n860 ;
  assign n862 = ~n742 & n831 ;
  assign n863 = ~n739 & ~n831 ;
  assign n864 = ~n862 & ~n863 ;
  assign n865 = ~n749 & ~n831 ;
  assign n866 = ~n752 & n831 ;
  assign n867 = ~n865 & ~n866 ;
  assign n868 = ~n762 & n831 ;
  assign n869 = ~n759 & ~n831 ;
  assign n870 = ~n868 & ~n869 ;
  assign n871 = ~n769 & ~n831 ;
  assign n872 = ~n772 & n831 ;
  assign n873 = ~n871 & ~n872 ;
  assign n874 = n782 & ~n831 ;
  assign n875 = n779 & n831 ;
  assign n876 = ~n874 & ~n875 ;
  assign n877 = ~n793 & n831 ;
  assign n878 = ~n790 & ~n831 ;
  assign n879 = ~n877 & ~n878 ;
  assign n880 = ~n803 & ~n831 ;
  assign n881 = ~n800 & n831 ;
  assign n882 = ~n880 & ~n881 ;
  assign n883 = n813 & ~n831 ;
  assign n884 = n810 & n831 ;
  assign n885 = ~n883 & ~n884 ;
  assign n886 = ~n823 & ~n831 ;
  assign n887 = ~n820 & n831 ;
  assign n888 = ~n886 & ~n887 ;
  assign n889 = n131 & n134 ;
  assign y0 = n843 ;
  assign y1 = ~n834 ;
  assign y2 = n831 ;
  assign y3 = ~n846 ;
  assign y4 = ~n849 ;
  assign y5 = ~n852 ;
  assign y6 = ~n855 ;
  assign y7 = ~n858 ;
  assign y8 = ~n861 ;
  assign y9 = ~n864 ;
  assign y10 = ~n867 ;
  assign y11 = ~n870 ;
  assign y12 = ~n873 ;
  assign y13 = n876 ;
  assign y14 = ~n879 ;
  assign y15 = ~n882 ;
  assign y16 = n885 ;
  assign y17 = ~n888 ;
  assign y18 = ~n889 ;
endmodule
