module bitonic_sort_inc_4_8 (in_array_0, in_array_1, in_array_2, in_array_3, in_array_4, in_array_5, in_array_6, in_array_7, in_array_8, in_array_9, in_array_10, in_array_11, in_array_12, in_array_13, in_array_14, in_array_15, in_array_16, in_array_17, in_array_18, in_array_19, in_array_20, in_array_21, in_array_22, in_array_23, in_array_24, in_array_25, in_array_26, in_array_27, in_array_28, in_array_29, in_array_30, in_array_31, out_array_0, out_array_1, out_array_2, out_array_3, out_array_4, out_array_5, out_array_6, out_array_7, out_array_8, out_array_9, out_array_10, out_array_11, out_array_12, out_array_13, out_array_14, out_array_15, out_array_16, out_array_17, out_array_18, out_array_19, out_array_20, out_array_21, out_array_22, out_array_23, out_array_24, out_array_25, out_array_26, out_array_27, out_array_28, out_array_29, out_array_30, out_array_31);
input in_array_0, in_array_1, in_array_2, in_array_3, in_array_4, in_array_5, in_array_6, in_array_7, in_array_8, in_array_9, in_array_10, in_array_11, in_array_12, in_array_13, in_array_14, in_array_15, in_array_16, in_array_17, in_array_18, in_array_19, in_array_20, in_array_21, in_array_22, in_array_23, in_array_24, in_array_25, in_array_26, in_array_27, in_array_28, in_array_29, in_array_30, in_array_31;
output out_array_0, out_array_1, out_array_2, out_array_3, out_array_4, out_array_5, out_array_6, out_array_7, out_array_8, out_array_9, out_array_10, out_array_11, out_array_12, out_array_13, out_array_14, out_array_15, out_array_16, out_array_17, out_array_18, out_array_19, out_array_20, out_array_21, out_array_22, out_array_23, out_array_24, out_array_25, out_array_26, out_array_27, out_array_28, out_array_29, out_array_30, out_array_31;
wire _0000_, _0001_, _0002_, _0003_, _0004_, _0005_, _0006_, _0007_, _0007__neg, _0008_, _0009_, _0010_, _0011_, _0012_, _0013_, _0014_, _0015_, _0016_, _0017_, _0018_, _0019_, _0020_, _0021_, _0022_, _0023_, _0024_, _0025_, _0026_, _0027_, _0028_, _0029_, _0030_, _0031_, _0032_, _0033_, _0034_, _0035_, _0036_, _0037_, _0038_, _0039_, _0040_, _0041_, _0042_, _0043_, _0044_, _0045_, _0046_, _0047_, _0048_, _0048__neg, _0049_, _0050_, _0051_, _0052_, _0053_, _0054_, _0055_, _0056_, _0057_, _0058_, _0059_, _0060_, _0061_, _0062_, _0063_, _0064_, _0065_, _0066_, _0067_, _0068_, _0069_, _0070_, _0071_, _0071__neg, _0072_, _0072__neg, _0073_, _0074_, _0075_, _0076_, _0076__neg, _0077_, _0078_, _0079_, _0080_, _0080__neg, _0081_, _0082_, _0083_, _0084_, _0085_, _0085__neg, _0086_, _0087_, _0088_, _0089_, _0090_, _0091_, _0092_, _0093_, _0094_, _0095_, _0096_, _0097_, _0097__neg, _0098_, _0099_, _0100_, _0101_, _0102_, _0102__neg, _0103_, _0104_, _0105_, _0106_, _0107_, _0108_, _0109_, _0110_, _0111_, _0112_, _0113_, _0114_, _0115_, _0116_, _0117_, _0118_, _0119_, _0120_, _0121_, _0122_, _0123_, _0124_, _0125_, _0126_, _0127_, _0128_, _0129_, _0130_, _0131_, _0132_, _0133_, _0134_, _0135_, _0136_, _0137_, _0138_, _0139_, _0140_, _0141_, _0142_, _0143_, _0144_, _0145_, _0146_, _0147_, _0148_, _0149_, _0150_, _0151_, _0152_, _0153_, _0153__neg, _0154_, _0155_, _0156_, _0157_, _0158_, _0159_, _0160_, _0161_, _0162_, _0163_, _0164_, _0165_, _0166_, _0167_, _0168_, _0169_, _0170_, _0171_, _0172_, _0173_, _0174_, _0175_, _0176_, _0177_, _0178_, _0179_, _0180_, _0181_, _0182_, _0183_, _0184_, _0185_, _0186_, _0187_, _0188_, _0189_, _0190_, _0191_, _0192_, _0192__neg, _0193_, _0194_, _0195_, _0196_, _0197_, _0198_, _0199_, _0200_, _0201_, _0202_, _0203_, _0204_, _0205_, _0206_, _0207_, _0208_, _0209_, _0210_, _0211_, _0212_, _0213_, _0214_, _0215_, _0216_, _0216__neg, _0217_, _0217__neg, _0218_, _0219_, _0220_, _0221_, _0221__neg, _0222_, _0223_, _0224_, _0225_, _0225__neg, _0226_, _0227_, _0228_, _0229_, _0230_, _0230__neg, _0231_, _0232_, _0233_, _0234_, _0235_, _0236_, _0237_, _0238_, _0239_, _0240_, _0240__neg, _0241_, _0242_, _0243_, _0244_, _0245_, _0246_, _0246__neg, _0247_, _0248_, _0249_, _0250_, _0251_, _0252_, _0253_, _0254_, _0254__neg, _0255_, _0255__neg, _0256_, _0257_, _0258_, _0259_, _0259__neg, _0260_, _0261_, _0262_, _0263_, _0263__neg, _0264_, _0265_, _0266_, _0267_, _0268_, _0268__neg, _0269_, _0270_, _0271_, _0272_, _0273_, _0274_, _0275_, _0276_, _0277_, _0278_, _0279_, _0280_, _0281_, _0282_, _0283_, _0284_, _0285_, _0286_, _0287_, _0288_, _0289_, _0290_, _0291_, _0292_, _0293_, _0294_, _0295_, _0295__neg, _0296_, _0297_, _0298_, _0299_, _0300_, _0301_, _0302_, _0303_, _0304_, _0305_, _0306_, _0307_, _0308_, _0309_, _0310_, _0311_, _0312_, _0313_, _0314_, _0315_, _0316_, _0317_, _0318_, _0319_, _0320_, _0321_, _0322_, _0323_, _0324_, _0325_, _0325__neg, _0326_, _0327_, _0328_, _0329_, _0330_, _0331_, _0332_, _0333_, _0334_, _0335_, _0336_, _0337_, _0338_, _0339_, _0340_, _0341_, _0342_, _0343_, _0344_, _0345_, _0346_, _0347_, _0348_, _0349_, _0350_, _0351_, _0352_, _0352__neg, _0353_, _0353__neg, _0354_, _0355_, _0356_, _0357_, _0357__neg, _0358_, _0359_, _0360_, _0361_, _0361__neg, _0362_, _0363_, _0364_, _0365_, _0366_, _0366__neg, _0367_, _0368_, _0369_, _0370_, _0371_, _0372_, _0373_, _0374_, _0375_, _0376_, _0377_, _0378_, _0379_, _0380_, _0381_, _0382_, _0383_, _0384_, _0385_, _0386_, _0387_, _0388_, _0389_, _0390_, _0390__neg, _0391_, _0391__neg, _0392_, _0393_, _0394_, _0395_, _0395__neg, _0396_, _0397_, _0398_, _0399_, _0399__neg, _0400_, _0401_, _0402_, _0403_, _0404_, _0404__neg, _0405_, _0406_, _0407_, _0408_, _0409_, _0410_, _0411_, _0412_, _0413_, _0414_, _0415_, _0416_, _0417_, _0418_, _0419_, _0420_, _0421_, _0422_, _0423_, _0424_, _0425_, _0426_, _0427_, _0428_, _0429_, _0430_, _0431_, _0432_, _0432__neg, _0433_, _0434_, _0435_, _0436_, _0437_, _0438_, _0439_, _0440_, _0441_, _0442_, _0443_, _0444_, _0445_, _0446_, _0447_, _0448_, _0449_, _0450_, _0451_, _0452_, _0453_, _0454_, _0455_, _0456_, _0457_, _0458_, _0459_, _0460_, _0461_, _0462_, _0462__neg, _0463_, _0464_, _0465_, _0466_, _0467_, _0468_, _0469_, _0470_, _0471_, _0472_, _0473_, _0474_, _0475_, _0476_, _0477_, _0478_, _0479_, _0480_, _0481_, _0482_, _0483_, _0484_, _0485_, _0486_, _0487_, _0488_, _0488__neg, _0489_, _0489__neg, _0490_, _0491_, _0492_, _0493_, _0493__neg, _0494_, _0495_, _0496_, _0497_, _0497__neg, _0498_, _0499_, _0500_, _0501_, _0502_, _0502__neg, _0503_, _0504_, _0505_, _0506_, _0507_, _0508_, _0509_, _0510_, _0511_, _0512_, _0513_, _0514_, _0515_, _0516_, _0517_, _0518_, _0519_, _0520_, _0521_, _0522_, _0523_, _0524_, _0525_, _0526_, _0526__neg, _0527_, _0528_, _0528__neg, _0529_, _0530_, _0531_, _0531__neg, _0532_, _0533_, _0534_, _0535_, _0536_, _0536__neg, _0537_, _0538_, _0539_, _0540_, _0540__neg, _0541_, _0542_, _0543_, _0544_, _0545_, _0546_, _0547_, _0548_, _0549_, _0550_, _0551_, _0552_, _0553_, _0554_, _0555_, _0556_, _0557_, _0558_, _0559_, _0560_, _0561_, _0562_, _0563_, _0564_, _0565_, _0565__neg, _0566_, _0567_, _0567__neg, _0568_, _0569_, _0570_, _0571_, _0572_, _0573_, _0574_, _0575_, _0576_, _0577_, _0578_, _0579_, _0580_, _0580__neg, _0581_, _0582_, _0583_, _0584_, _0585_, _0586_, _0587_, _0588_, _0589_, _0590_, _0591_, _0592_, _0593_, _0594_, _0595_, _0596_, _0597_, _0598_, _0599_, _0600_, _0601_, _0602_, _0603_, _0604_, _0605_, _0606_, _0607_, _0607__neg, _0608_, _0609_, _0610_, _0610__neg, _0611_, _0612_, _0613_, _0614_, _0615_, _0616_, _0617_, _0618_, _0619_, _0620_, _0621_, _0622_, _0623_, _0624_, _0625_, _0625__neg, _0626_, _0627_, _0628_, _0629_, _0630_, _0631_, _0632_, _0633_, _0634_, _0635_, _0636_, _0637_, _0638_, _0639_, _0640_, _0641_, _0642_, _0643_, _0644_, _0645_, _0646_, _0647_, _0648_, _0649_, _0650_, _0651_, _0652_, _0653_, _0654_, _0655_, _0656_, _0657_, _0658_, _0658__neg, _0659_, _0660_, _0661_, _0662_, _0663_, _0664_, _0665_, _0666_, _0667_, _0668_, _0669_, _0670_, _0671_, _0672_, _0673_, _0674_, _0675_, _0676_, _0677_, _0678_, _0679_, _0680_, _0681_, _0682_, _0683_, _0684_, _0685_, _0686_, _0686__neg, _0687_, _0688_, _0689_, _0689__neg, _0690_, _0691_, _0692_, _0692__neg, _0693_, _0694_, _0695_, _0696_, _0697_, _0697__neg, _0698_, _0699_, _0700_, _0701_, _0702_, _0702__neg, _0703_, _0704_, _0705_, _0706_, _0707_, _0708_, _0709_, _0710_, _0711_, _0712_, _0713_, _0714_, _0715_, _0716_, _0717_, _0718_, _0719_, _0720_, _0721_, _0722_, _0723_, _0724_, _0725_, _0726_, _0727_, _0727__neg, _0728_, _0729_, _0729__neg, _0730_, _0731_, _0732_, _0733_, _0734_, _0735_, _0736_, _0737_, _0738_, _0739_, _0740_, _0741_, _0742_, _0742__neg, _0743_, _0744_, _0745_, _0746_, _0747_, _0748_, _0749_, _0750_, _0751_, _0752_, _0753_, _0754_, _0755_, _0756_, _0757_, _0758_, _0759_, _0760_, _0761_, _0762_, _0763_, _0764_, _0765_, _0766_, _0767_, _0768_, _0769_, _0770_, _0770__neg, _0771_, _0772_, _0772__neg, _0773_, _0774_, _0775_, _0776_, _0777_, _0778_, _0779_, _0780_, _0781_, _0782_, _0783_, _0784_, _0785_, _0786_, _0787_, _0788_, _0789_, _0790_, _0791_, _0792_, _0793_;
assign _0550_ = ~in_array_6;
assign _0561_ = in_array_2 ^ in_array_6;
assign _0569_ = ~in_array_0;
assign _0576_ = in_array_4 & _0569_;
assign _0587_ = ~in_array_1;
assign _0598_ = _0576_ ^ _0587_;
assign _0608_ = _0576_ ^ in_array_5;
assign _0615_ = _0608_ & _0598_;
assign _0622_ = _0615_ ^ _0576_;
assign _0633_ = ~in_array_2;
assign _0644_ = _0622_ ^ _0633_;
assign _0655_ = _0622_ ^ in_array_6;
assign _0666_ = _0655_ & _0644_;
assign _0677_ = _0666_ ^ _0622_;
assign _0688_ = ~_0677_;
assign _0699_ = ~in_array_3;
assign _0710_ = _0677_ ^ _0699_;
assign _0721_ = _0677_ ^ in_array_7;
assign _0730_ = _0721_ & _0710_;
assign _0737_ = _0730_ ^ _0688_;
assign _0747_ = _0737_ & _0561_;
assign _0758_ = _0747_ ^ _0550_;
assign _0769_ = in_array_10 ^ in_array_14;
assign _0776_ = ~in_array_8;
assign _0783_ = in_array_12 & _0776_;
assign _0784_ = ~in_array_9;
assign _0785_ = _0783_ ^ _0784_;
assign _0786_ = _0783_ ^ in_array_13;
assign _0787_ = _0786_ & _0785_;
assign _0788_ = _0787_ ^ _0783_;
assign _0789_ = ~in_array_10;
assign _0790_ = _0788_ ^ _0789_;
assign _0791_ = _0788_ ^ in_array_14;
assign _0792_ = _0791_ & _0790_;
assign _0793_ = _0792_ ^ _0788_;
assign _0000_ = ~in_array_11;
assign _0001_ = _0793_ ^ _0000_;
assign _0002_ = _0793_ ^ in_array_15;
assign _0003_ = _0002_ & _0001_;
assign _0004_ = _0003_ ^ _0793_;
assign _0005_ = _0004_ & _0769_;
assign _0006_ = _0005_ ^ in_array_14;
assign _0007__neg = _0006_ ^ _0758_;
assign _0007_ = ~_0007__neg;
assign _0008_ = ~in_array_4;
assign _0009_ = in_array_4 ^ in_array_0;
assign _0010_ = _0009_ & _0737_;
assign _0011_ = _0010_ ^ _0008_;
assign _0012_ = in_array_12 ^ in_array_8;
assign _0013_ = _0012_ & _0004_;
assign _0014_ = _0013_ ^ in_array_12;
assign _0015_ = _0014_ & _0011_;
assign _0016_ = ~in_array_5;
assign _0017_ = in_array_1 ^ in_array_5;
assign _0018_ = _0017_ & _0737_;
assign _0019_ = _0018_ ^ _0016_;
assign _0020_ = _0019_ ^ _0015_;
assign _0021_ = in_array_9 ^ in_array_13;
assign _0022_ = _0021_ & _0004_;
assign _0023_ = _0022_ ^ in_array_13;
assign _0024_ = _0023_ ^ _0015_;
assign _0025_ = _0024_ & _0020_;
assign _0026_ = _0025_ ^ _0015_;
assign _0027_ = ~_0026_;
assign _0028_ = _0026_ ^ _0758_;
assign _0029_ = _0026_ ^ _0006_;
assign _0030_ = _0029_ & _0028_;
assign _0031_ = _0030_ ^ _0027_;
assign _0032_ = ~in_array_7;
assign _0033_ = in_array_3 & _0032_;
assign _0034_ = _0033_ ^ _0032_;
assign _0035_ = ~_0034_;
assign _0036_ = _0035_ ^ _0031_;
assign _0037_ = _0000_ & in_array_15;
assign _0038_ = _0037_ ^ in_array_15;
assign _0039_ = ~_0038_;
assign _0040_ = _0039_ ^ _0031_;
assign _0041_ = _0040_ & _0036_;
assign _0042_ = _0041_ ^ _0031_;
assign _0043_ = _0042_ & _0007_;
assign _0044_ = _0043_ ^ _0758_;
assign _0045_ = _0747_ ^ _0633_;
assign _0046_ = ~_0045_;
assign _0047_ = _0005_ ^ in_array_10;
assign _0048__neg = _0047_ ^ _0045_;
assign _0048_ = ~_0048__neg;
assign _0049_ = _0010_ ^ _0569_;
assign _0050_ = _0013_ ^ in_array_8;
assign _0051_ = _0050_ & _0049_;
assign _0052_ = _0018_ ^ _0587_;
assign _0053_ = _0052_ ^ _0051_;
assign _0054_ = _0022_ ^ in_array_9;
assign _0055_ = _0054_ ^ _0051_;
assign _0056_ = _0055_ & _0053_;
assign _0057_ = _0056_ ^ _0051_;
assign _0058_ = ~_0057_;
assign _0059_ = _0057_ ^ _0045_;
assign _0060_ = _0057_ ^ _0047_;
assign _0061_ = _0060_ & _0059_;
assign _0062_ = _0061_ ^ _0058_;
assign _0063_ = _0033_ ^ in_array_3;
assign _0064_ = _0063_ ^ _0062_;
assign _0065_ = _0037_ ^ _0000_;
assign _0066_ = _0065_ ^ _0062_;
assign _0067_ = _0066_ & _0064_;
assign _0068_ = _0067_ ^ _0062_;
assign _0069_ = _0068_ & _0048_;
assign _0070_ = _0069_ ^ _0046_;
assign _0071__neg = _0070_ ^ _0044_;
assign _0071_ = ~_0071__neg;
assign _0072__neg = _0014_ ^ _0011_;
assign _0072_ = ~_0072__neg;
assign _0073_ = _0072_ & _0042_;
assign _0074_ = _0073_ ^ _0011_;
assign _0075_ = ~_0049_;
assign _0076__neg = _0050_ ^ _0049_;
assign _0076_ = ~_0076__neg;
assign _0077_ = _0076_ & _0068_;
assign _0078_ = _0077_ ^ _0075_;
assign _0079_ = _0078_ & _0074_;
assign _0080__neg = _0023_ ^ _0019_;
assign _0080_ = ~_0080__neg;
assign _0081_ = _0080_ & _0042_;
assign _0082_ = _0081_ ^ _0019_;
assign _0083_ = _0082_ ^ _0079_;
assign _0084_ = ~_0052_;
assign _0085__neg = _0054_ ^ _0052_;
assign _0085_ = ~_0085__neg;
assign _0086_ = _0085_ & _0068_;
assign _0087_ = _0086_ ^ _0084_;
assign _0088_ = _0087_ ^ _0079_;
assign _0089_ = _0088_ & _0083_;
assign _0090_ = _0089_ ^ _0079_;
assign _0091_ = ~_0090_;
assign _0092_ = _0090_ ^ _0044_;
assign _0093_ = _0090_ ^ _0070_;
assign _0094_ = _0093_ & _0092_;
assign _0095_ = _0094_ ^ _0091_;
assign _0096_ = _0094_ ^ _0090_;
assign _0097__neg = _0038_ ^ _0034_;
assign _0097_ = ~_0097__neg;
assign _0098_ = _0097_ & _0042_;
assign _0099_ = _0098_ ^ _0034_;
assign _0100_ = _0099_ ^ _0096_;
assign _0101_ = ~_0063_;
assign _0102__neg = _0065_ ^ _0063_;
assign _0102_ = ~_0102__neg;
assign _0103_ = _0102_ & _0068_;
assign _0104_ = _0103_ ^ _0101_;
assign _0105_ = _0104_ ^ _0095_;
assign _0106_ = _0105_ & _0100_;
assign _0107_ = _0106_ ^ _0095_;
assign _0108_ = _0107_ & _0071_;
assign _0109_ = _0108_ ^ _0044_;
assign _0110_ = ~_0109_;
assign _0111_ = ~in_array_22;
assign _0112_ = in_array_18 ^ in_array_22;
assign _0113_ = ~in_array_16;
assign _0114_ = in_array_20 & _0113_;
assign _0115_ = ~in_array_17;
assign _0116_ = _0114_ ^ _0115_;
assign _0117_ = _0114_ ^ in_array_21;
assign _0118_ = _0117_ & _0116_;
assign _0119_ = _0118_ ^ _0114_;
assign _0120_ = ~in_array_18;
assign _0121_ = _0119_ ^ _0120_;
assign _0122_ = _0119_ ^ in_array_22;
assign _0123_ = _0122_ & _0121_;
assign _0124_ = _0123_ ^ _0119_;
assign _0125_ = ~_0124_;
assign _0126_ = ~in_array_19;
assign _0127_ = _0124_ ^ _0126_;
assign _0128_ = _0124_ ^ in_array_23;
assign _0129_ = _0128_ & _0127_;
assign _0130_ = _0129_ ^ _0125_;
assign _0131_ = _0130_ & _0112_;
assign _0132_ = _0131_ ^ _0111_;
assign _0133_ = in_array_26 ^ in_array_30;
assign _0134_ = ~in_array_24;
assign _0135_ = in_array_28 & _0134_;
assign _0136_ = ~in_array_25;
assign _0137_ = _0135_ ^ _0136_;
assign _0138_ = _0135_ ^ in_array_29;
assign _0139_ = _0138_ & _0137_;
assign _0140_ = _0139_ ^ _0135_;
assign _0141_ = ~in_array_26;
assign _0142_ = _0140_ ^ _0141_;
assign _0143_ = _0140_ ^ in_array_30;
assign _0144_ = _0143_ & _0142_;
assign _0145_ = _0144_ ^ _0140_;
assign _0146_ = ~in_array_27;
assign _0147_ = _0145_ ^ _0146_;
assign _0148_ = _0145_ ^ in_array_31;
assign _0149_ = _0148_ & _0147_;
assign _0150_ = _0149_ ^ _0145_;
assign _0151_ = _0150_ & _0133_;
assign _0152_ = _0151_ ^ in_array_30;
assign _0153__neg = _0152_ ^ _0132_;
assign _0153_ = ~_0153__neg;
assign _0154_ = ~in_array_20;
assign _0155_ = in_array_20 ^ in_array_16;
assign _0156_ = _0155_ & _0130_;
assign _0157_ = _0156_ ^ _0154_;
assign _0158_ = in_array_28 ^ in_array_24;
assign _0159_ = _0158_ & _0150_;
assign _0160_ = _0159_ ^ in_array_28;
assign _0161_ = _0160_ & _0157_;
assign _0162_ = ~in_array_21;
assign _0163_ = in_array_17 ^ in_array_21;
assign _0164_ = _0163_ & _0130_;
assign _0165_ = _0164_ ^ _0162_;
assign _0166_ = _0165_ ^ _0161_;
assign _0167_ = in_array_25 ^ in_array_29;
assign _0168_ = _0167_ & _0150_;
assign _0169_ = _0168_ ^ in_array_29;
assign _0170_ = _0169_ ^ _0161_;
assign _0171_ = _0170_ & _0166_;
assign _0172_ = _0171_ ^ _0161_;
assign _0173_ = _0172_ ^ _0132_;
assign _0174_ = _0172_ ^ _0152_;
assign _0175_ = _0174_ & _0173_;
assign _0176_ = _0175_ ^ _0172_;
assign _0177_ = ~in_array_23;
assign _0178_ = in_array_19 & _0177_;
assign _0179_ = _0178_ ^ _0177_;
assign _0180_ = _0179_ ^ _0176_;
assign _0181_ = _0146_ & in_array_31;
assign _0182_ = _0181_ ^ in_array_31;
assign _0183_ = _0182_ ^ _0176_;
assign _0184_ = _0183_ & _0180_;
assign _0185_ = _0184_ ^ _0176_;
assign _0186_ = _0185_ & _0153_;
assign _0187_ = _0186_ ^ _0132_;
assign _0188_ = ~_0187_;
assign _0189_ = _0131_ ^ _0120_;
assign _0190_ = ~_0189_;
assign _0191_ = _0151_ ^ in_array_26;
assign _0192__neg = _0191_ ^ _0189_;
assign _0192_ = ~_0192__neg;
assign _0193_ = _0156_ ^ _0113_;
assign _0194_ = _0159_ ^ in_array_24;
assign _0195_ = _0194_ & _0193_;
assign _0196_ = _0164_ ^ _0115_;
assign _0197_ = _0196_ ^ _0195_;
assign _0198_ = _0168_ ^ in_array_25;
assign _0199_ = _0198_ ^ _0195_;
assign _0200_ = _0199_ & _0197_;
assign _0201_ = _0200_ ^ _0195_;
assign _0202_ = _0201_ ^ _0189_;
assign _0203_ = _0201_ ^ _0191_;
assign _0204_ = _0203_ & _0202_;
assign _0205_ = _0204_ ^ _0201_;
assign _0206_ = _0178_ ^ in_array_19;
assign _0207_ = ~_0206_;
assign _0208_ = _0207_ ^ _0205_;
assign _0209_ = _0181_ ^ _0146_;
assign _0210_ = ~_0209_;
assign _0211_ = _0210_ ^ _0205_;
assign _0212_ = _0211_ & _0208_;
assign _0213_ = _0212_ ^ _0205_;
assign _0214_ = _0213_ & _0192_;
assign _0215_ = _0214_ ^ _0190_;
assign _0216__neg = _0215_ ^ _0187_;
assign _0216_ = ~_0216__neg;
assign _0217__neg = _0160_ ^ _0157_;
assign _0217_ = ~_0217__neg;
assign _0218_ = _0217_ & _0185_;
assign _0219_ = _0218_ ^ _0157_;
assign _0220_ = ~_0193_;
assign _0221__neg = _0194_ ^ _0193_;
assign _0221_ = ~_0221__neg;
assign _0222_ = _0221_ & _0213_;
assign _0223_ = _0222_ ^ _0220_;
assign _0224_ = _0223_ & _0219_;
assign _0225__neg = _0169_ ^ _0165_;
assign _0225_ = ~_0225__neg;
assign _0226_ = _0225_ & _0185_;
assign _0227_ = _0226_ ^ _0165_;
assign _0228_ = _0227_ ^ _0224_;
assign _0229_ = ~_0196_;
assign _0230__neg = _0198_ ^ _0196_;
assign _0230_ = ~_0230__neg;
assign _0231_ = _0230_ & _0213_;
assign _0232_ = _0231_ ^ _0229_;
assign _0233_ = _0232_ ^ _0224_;
assign _0234_ = _0233_ & _0228_;
assign _0235_ = _0234_ ^ _0224_;
assign _0236_ = _0235_ ^ _0187_;
assign _0237_ = _0235_ ^ _0215_;
assign _0238_ = _0237_ & _0236_;
assign _0239_ = _0238_ ^ _0235_;
assign _0240__neg = _0182_ ^ _0179_;
assign _0240_ = ~_0240__neg;
assign _0241_ = _0240_ & _0185_;
assign _0242_ = _0241_ ^ _0179_;
assign _0243_ = _0242_ ^ _0239_;
assign _0244_ = ~_0235_;
assign _0245_ = _0238_ ^ _0244_;
assign _0246__neg = _0209_ ^ _0206_;
assign _0246_ = ~_0246__neg;
assign _0247_ = _0246_ & _0213_;
assign _0248_ = _0247_ ^ _0207_;
assign _0249_ = _0248_ ^ _0245_;
assign _0250_ = _0249_ & _0243_;
assign _0251_ = _0250_ ^ _0239_;
assign _0252_ = _0251_ & _0216_;
assign _0253_ = _0252_ ^ _0188_;
assign _0254__neg = _0253_ ^ _0109_;
assign _0254_ = ~_0254__neg;
assign _0255__neg = _0078_ ^ _0074_;
assign _0255_ = ~_0255__neg;
assign _0256_ = _0255_ & _0107_;
assign _0257_ = _0256_ ^ _0074_;
assign _0258_ = ~_0219_;
assign _0259__neg = _0223_ ^ _0219_;
assign _0259_ = ~_0259__neg;
assign _0260_ = _0259_ & _0251_;
assign _0261_ = _0260_ ^ _0258_;
assign _0262_ = _0261_ & _0257_;
assign _0263__neg = _0087_ ^ _0082_;
assign _0263_ = ~_0263__neg;
assign _0264_ = _0263_ & _0107_;
assign _0265_ = _0264_ ^ _0082_;
assign _0266_ = _0265_ ^ _0262_;
assign _0267_ = ~_0227_;
assign _0268__neg = _0232_ ^ _0227_;
assign _0268_ = ~_0268__neg;
assign _0269_ = _0268_ & _0251_;
assign _0270_ = _0269_ ^ _0267_;
assign _0271_ = _0270_ ^ _0262_;
assign _0272_ = _0271_ & _0266_;
assign _0273_ = _0272_ ^ _0262_;
assign _0274_ = ~_0273_;
assign _0275_ = _0273_ ^ _0109_;
assign _0276_ = _0273_ ^ _0253_;
assign _0277_ = _0276_ & _0275_;
assign _0278_ = _0277_ ^ _0274_;
assign _0279_ = _0277_ ^ _0273_;
assign _0280_ = _0104_ ^ _0099_;
assign _0281_ = _0280_ & _0107_;
assign _0282_ = _0281_ ^ _0099_;
assign _0283_ = _0282_ ^ _0279_;
assign _0284_ = _0248_ ^ _0242_;
assign _0285_ = _0284_ & _0251_;
assign _0286_ = _0285_ ^ _0242_;
assign _0287_ = _0286_ ^ _0278_;
assign _0288_ = _0287_ & _0283_;
assign _0289_ = _0288_ ^ _0278_;
assign _0290_ = _0289_ & _0254_;
assign _0291_ = _0290_ ^ _0110_;
assign _0292_ = ~_0006_;
assign _0293_ = _0043_ ^ _0292_;
assign _0294_ = _0069_ ^ _0047_;
assign _0295__neg = _0294_ ^ _0293_;
assign _0295_ = ~_0295__neg;
assign _0296_ = ~_0014_;
assign _0297_ = _0073_ ^ _0296_;
assign _0298_ = _0077_ ^ _0050_;
assign _0299_ = _0298_ & _0297_;
assign _0300_ = ~_0023_;
assign _0301_ = _0081_ ^ _0300_;
assign _0302_ = _0301_ ^ _0299_;
assign _0303_ = _0086_ ^ _0054_;
assign _0304_ = _0303_ ^ _0299_;
assign _0305_ = _0304_ & _0302_;
assign _0306_ = _0305_ ^ _0299_;
assign _0307_ = ~_0306_;
assign _0308_ = _0306_ ^ _0293_;
assign _0309_ = _0306_ ^ _0294_;
assign _0310_ = _0309_ & _0308_;
assign _0311_ = _0310_ ^ _0307_;
assign _0312_ = _0310_ ^ _0306_;
assign _0313_ = _0098_ ^ _0039_;
assign _0314_ = _0313_ ^ _0312_;
assign _0315_ = _0103_ ^ _0065_;
assign _0316_ = _0315_ ^ _0311_;
assign _0317_ = _0316_ & _0314_;
assign _0318_ = _0317_ ^ _0311_;
assign _0319_ = _0318_ & _0295_;
assign _0320_ = _0319_ ^ _0293_;
assign _0321_ = ~_0152_;
assign _0322_ = _0186_ ^ _0321_;
assign _0323_ = ~_0322_;
assign _0324_ = _0214_ ^ _0191_;
assign _0325__neg = _0324_ ^ _0322_;
assign _0325_ = ~_0325__neg;
assign _0326_ = ~_0160_;
assign _0327_ = _0218_ ^ _0326_;
assign _0328_ = _0222_ ^ _0194_;
assign _0329_ = _0328_ & _0327_;
assign _0330_ = ~_0169_;
assign _0331_ = _0226_ ^ _0330_;
assign _0332_ = _0331_ ^ _0329_;
assign _0333_ = _0231_ ^ _0198_;
assign _0334_ = _0333_ ^ _0329_;
assign _0335_ = _0334_ & _0332_;
assign _0336_ = _0335_ ^ _0329_;
assign _0337_ = _0336_ ^ _0322_;
assign _0338_ = _0336_ ^ _0324_;
assign _0339_ = _0338_ & _0337_;
assign _0340_ = _0339_ ^ _0336_;
assign _0341_ = ~_0182_;
assign _0342_ = _0241_ ^ _0341_;
assign _0343_ = _0342_ ^ _0340_;
assign _0344_ = ~_0336_;
assign _0345_ = _0339_ ^ _0344_;
assign _0346_ = _0247_ ^ _0209_;
assign _0347_ = _0346_ ^ _0345_;
assign _0348_ = _0347_ & _0343_;
assign _0349_ = _0348_ ^ _0340_;
assign _0350_ = _0349_ & _0325_;
assign _0351_ = _0350_ ^ _0323_;
assign _0352__neg = _0351_ ^ _0320_;
assign _0352_ = ~_0352__neg;
assign _0353__neg = _0298_ ^ _0297_;
assign _0353_ = ~_0353__neg;
assign _0354_ = _0353_ & _0318_;
assign _0355_ = _0354_ ^ _0297_;
assign _0356_ = ~_0327_;
assign _0357__neg = _0328_ ^ _0327_;
assign _0357_ = ~_0357__neg;
assign _0358_ = _0357_ & _0349_;
assign _0359_ = _0358_ ^ _0356_;
assign _0360_ = _0359_ & _0355_;
assign _0361__neg = _0303_ ^ _0301_;
assign _0361_ = ~_0361__neg;
assign _0362_ = _0361_ & _0318_;
assign _0363_ = _0362_ ^ _0301_;
assign _0364_ = _0363_ ^ _0360_;
assign _0365_ = ~_0331_;
assign _0366__neg = _0333_ ^ _0331_;
assign _0366_ = ~_0366__neg;
assign _0367_ = _0366_ & _0349_;
assign _0368_ = _0367_ ^ _0365_;
assign _0369_ = _0368_ ^ _0360_;
assign _0370_ = _0369_ & _0364_;
assign _0371_ = _0370_ ^ _0360_;
assign _0372_ = ~_0371_;
assign _0373_ = _0371_ ^ _0320_;
assign _0374_ = _0371_ ^ _0351_;
assign _0375_ = _0374_ & _0373_;
assign _0376_ = _0375_ ^ _0372_;
assign _0377_ = _0375_ ^ _0371_;
assign _0378_ = _0315_ ^ _0313_;
assign _0379_ = _0378_ & _0318_;
assign _0380_ = _0379_ ^ _0313_;
assign _0381_ = _0380_ ^ _0377_;
assign _0382_ = _0346_ ^ _0342_;
assign _0383_ = _0382_ & _0349_;
assign _0384_ = _0383_ ^ _0342_;
assign _0385_ = _0384_ ^ _0376_;
assign _0386_ = _0385_ & _0381_;
assign _0387_ = _0386_ ^ _0376_;
assign _0388_ = _0387_ & _0352_;
assign _0389_ = _0388_ ^ _0320_;
assign _0390__neg = _0389_ ^ _0291_;
assign _0390_ = ~_0390__neg;
assign _0391__neg = _0359_ ^ _0355_;
assign _0391_ = ~_0391__neg;
assign _0392_ = _0391_ & _0387_;
assign _0393_ = _0392_ ^ _0355_;
assign _0394_ = ~_0257_;
assign _0395__neg = _0261_ ^ _0257_;
assign _0395_ = ~_0395__neg;
assign _0396_ = _0395_ & _0289_;
assign _0397_ = _0396_ ^ _0394_;
assign _0398_ = _0397_ & _0393_;
assign _0399__neg = _0368_ ^ _0363_;
assign _0399_ = ~_0399__neg;
assign _0400_ = _0399_ & _0387_;
assign _0401_ = _0400_ ^ _0363_;
assign _0402_ = _0401_ ^ _0398_;
assign _0403_ = ~_0265_;
assign _0404__neg = _0270_ ^ _0265_;
assign _0404_ = ~_0404__neg;
assign _0405_ = _0404_ & _0289_;
assign _0406_ = _0405_ ^ _0403_;
assign _0407_ = _0406_ ^ _0398_;
assign _0408_ = _0407_ & _0402_;
assign _0409_ = _0408_ ^ _0398_;
assign _0410_ = ~_0409_;
assign _0411_ = _0409_ ^ _0389_;
assign _0412_ = _0409_ ^ _0291_;
assign _0413_ = _0412_ & _0411_;
assign _0414_ = _0413_ ^ _0410_;
assign _0415_ = _0413_ ^ _0409_;
assign _0416_ = _0384_ ^ _0380_;
assign _0417_ = _0416_ & _0387_;
assign _0418_ = _0417_ ^ _0380_;
assign _0419_ = _0418_ ^ _0415_;
assign _0420_ = _0286_ ^ _0282_;
assign _0421_ = _0420_ & _0289_;
assign _0422_ = _0421_ ^ _0282_;
assign _0423_ = _0422_ ^ _0414_;
assign _0424_ = _0423_ & _0419_;
assign _0425_ = _0424_ ^ _0414_;
assign _0426_ = _0425_ & _0390_;
assign _0427_ = _0426_ ^ _0291_;
assign _0428_ = ~_0070_;
assign _0429_ = _0108_ ^ _0428_;
assign _0430_ = ~_0429_;
assign _0431_ = _0252_ ^ _0215_;
assign _0432__neg = _0431_ ^ _0429_;
assign _0432_ = ~_0432__neg;
assign _0433_ = ~_0078_;
assign _0434_ = _0256_ ^ _0433_;
assign _0435_ = _0260_ ^ _0223_;
assign _0436_ = _0435_ & _0434_;
assign _0437_ = ~_0087_;
assign _0438_ = _0264_ ^ _0437_;
assign _0439_ = _0438_ ^ _0436_;
assign _0440_ = _0269_ ^ _0232_;
assign _0441_ = _0440_ ^ _0436_;
assign _0442_ = _0441_ & _0439_;
assign _0443_ = _0442_ ^ _0436_;
assign _0444_ = ~_0443_;
assign _0445_ = _0443_ ^ _0429_;
assign _0446_ = _0443_ ^ _0431_;
assign _0447_ = _0446_ & _0445_;
assign _0448_ = _0447_ ^ _0444_;
assign _0449_ = _0447_ ^ _0443_;
assign _0450_ = _0281_ ^ _0104_;
assign _0451_ = _0450_ ^ _0449_;
assign _0452_ = _0285_ ^ _0248_;
assign _0453_ = _0452_ ^ _0448_;
assign _0454_ = _0453_ & _0451_;
assign _0455_ = _0454_ ^ _0448_;
assign _0456_ = _0455_ & _0432_;
assign _0457_ = _0456_ ^ _0430_;
assign _0458_ = ~_0457_;
assign _0459_ = ~_0294_;
assign _0460_ = _0319_ ^ _0459_;
assign _0461_ = _0350_ ^ _0324_;
assign _0462__neg = _0461_ ^ _0460_;
assign _0462_ = ~_0462__neg;
assign _0463_ = ~_0298_;
assign _0464_ = _0354_ ^ _0463_;
assign _0465_ = _0358_ ^ _0328_;
assign _0466_ = _0465_ & _0464_;
assign _0467_ = ~_0303_;
assign _0468_ = _0362_ ^ _0467_;
assign _0469_ = _0468_ ^ _0466_;
assign _0470_ = _0367_ ^ _0333_;
assign _0471_ = _0470_ ^ _0466_;
assign _0472_ = _0471_ & _0469_;
assign _0473_ = _0472_ ^ _0466_;
assign _0474_ = ~_0473_;
assign _0475_ = _0473_ ^ _0460_;
assign _0476_ = _0473_ ^ _0461_;
assign _0477_ = _0476_ & _0475_;
assign _0478_ = _0477_ ^ _0474_;
assign _0479_ = _0477_ ^ _0473_;
assign _0480_ = _0379_ ^ _0315_;
assign _0481_ = _0480_ ^ _0479_;
assign _0482_ = _0383_ ^ _0346_;
assign _0483_ = _0482_ ^ _0478_;
assign _0484_ = _0483_ & _0481_;
assign _0485_ = _0484_ ^ _0478_;
assign _0486_ = _0485_ & _0462_;
assign _0487_ = _0486_ ^ _0460_;
assign _0488__neg = _0487_ ^ _0457_;
assign _0488_ = ~_0488__neg;
assign _0489__neg = _0465_ ^ _0464_;
assign _0489_ = ~_0489__neg;
assign _0490_ = _0489_ & _0485_;
assign _0491_ = _0490_ ^ _0464_;
assign _0492_ = ~_0434_;
assign _0493__neg = _0435_ ^ _0434_;
assign _0493_ = ~_0493__neg;
assign _0494_ = _0493_ & _0455_;
assign _0495_ = _0494_ ^ _0492_;
assign _0496_ = _0495_ & _0491_;
assign _0497__neg = _0470_ ^ _0468_;
assign _0497_ = ~_0497__neg;
assign _0498_ = _0497_ & _0485_;
assign _0499_ = _0498_ ^ _0468_;
assign _0500_ = _0499_ ^ _0496_;
assign _0501_ = ~_0438_;
assign _0502__neg = _0440_ ^ _0438_;
assign _0502_ = ~_0502__neg;
assign _0503_ = _0502_ & _0455_;
assign _0504_ = _0503_ ^ _0501_;
assign _0505_ = _0504_ ^ _0496_;
assign _0506_ = _0505_ & _0500_;
assign _0507_ = _0506_ ^ _0496_;
assign _0508_ = ~_0507_;
assign _0509_ = _0507_ ^ _0487_;
assign _0510_ = _0507_ ^ _0457_;
assign _0511_ = _0510_ & _0509_;
assign _0512_ = _0511_ ^ _0508_;
assign _0513_ = _0511_ ^ _0507_;
assign _0514_ = _0482_ ^ _0480_;
assign _0515_ = _0514_ & _0485_;
assign _0516_ = _0515_ ^ _0480_;
assign _0517_ = _0516_ ^ _0513_;
assign _0518_ = _0452_ ^ _0450_;
assign _0519_ = _0518_ & _0455_;
assign _0520_ = _0519_ ^ _0450_;
assign _0521_ = _0520_ ^ _0512_;
assign _0522_ = _0521_ & _0517_;
assign _0523_ = _0522_ ^ _0512_;
assign _0524_ = _0523_ & _0488_;
assign _0525_ = _0524_ ^ _0458_;
assign _0526__neg = _0525_ ^ _0427_;
assign _0526_ = ~_0526__neg;
assign _0527_ = ~_0495_;
assign _0528__neg = _0495_ ^ _0491_;
assign _0528_ = ~_0528__neg;
assign _0529_ = _0528_ & _0523_;
assign _0530_ = _0529_ ^ _0527_;
assign _0531__neg = _0397_ ^ _0393_;
assign _0531_ = ~_0531__neg;
assign _0532_ = _0531_ & _0425_;
assign _0533_ = _0532_ ^ _0397_;
assign _0534_ = _0533_ & _0530_;
assign _0535_ = ~_0504_;
assign _0536__neg = _0504_ ^ _0499_;
assign _0536_ = ~_0536__neg;
assign _0537_ = _0536_ & _0523_;
assign _0538_ = _0537_ ^ _0535_;
assign _0539_ = _0538_ ^ _0534_;
assign _0540__neg = _0406_ ^ _0401_;
assign _0540_ = ~_0540__neg;
assign _0541_ = _0540_ & _0425_;
assign _0542_ = _0541_ ^ _0406_;
assign _0543_ = _0542_ ^ _0534_;
assign _0544_ = _0543_ & _0539_;
assign _0545_ = _0544_ ^ _0534_;
assign _0546_ = ~_0545_;
assign _0547_ = _0545_ ^ _0525_;
assign _0548_ = _0545_ ^ _0427_;
assign _0549_ = _0548_ & _0547_;
assign _0551_ = _0549_ ^ _0546_;
assign _0552_ = _0549_ ^ _0545_;
assign _0553_ = _0520_ ^ _0516_;
assign _0554_ = _0553_ & _0523_;
assign _0555_ = _0554_ ^ _0520_;
assign _0556_ = _0555_ ^ _0552_;
assign _0557_ = _0422_ ^ _0418_;
assign _0558_ = _0557_ & _0425_;
assign _0559_ = _0558_ ^ _0422_;
assign _0560_ = _0559_ ^ _0551_;
assign _0562_ = _0560_ & _0556_;
assign _0563_ = _0562_ ^ _0551_;
assign _0564_ = _0563_ & _0526_;
assign out_array_18 = _0564_ ^ _0427_;
assign _0565__neg = _0542_ ^ _0538_;
assign _0565_ = ~_0565__neg;
assign _0566_ = _0565_ & _0563_;
assign out_array_17 = _0566_ ^ _0542_;
assign _0567__neg = _0533_ ^ _0530_;
assign _0567_ = ~_0567__neg;
assign _0568_ = _0567_ & _0563_;
assign out_array_16 = _0568_ ^ _0533_;
assign _0570_ = ~_0525_;
assign out_array_22 = _0564_ ^ _0570_;
assign _0571_ = ~_0538_;
assign out_array_21 = _0566_ ^ _0571_;
assign _0572_ = ~_0530_;
assign out_array_20 = _0568_ ^ _0572_;
assign _0573_ = ~_0559_;
assign _0574_ = _0559_ ^ _0555_;
assign _0575_ = _0574_ & _0563_;
assign out_array_19 = _0575_ ^ _0573_;
assign _0577_ = ~_0389_;
assign _0578_ = _0426_ ^ _0577_;
assign _0579_ = _0524_ ^ _0487_;
assign _0580__neg = _0579_ ^ _0578_;
assign _0580_ = ~_0580__neg;
assign _0581_ = _0529_ ^ _0491_;
assign _0582_ = ~_0393_;
assign _0583_ = _0532_ ^ _0582_;
assign _0584_ = _0583_ & _0581_;
assign _0585_ = _0537_ ^ _0499_;
assign _0586_ = _0585_ ^ _0584_;
assign _0588_ = ~_0401_;
assign _0589_ = _0541_ ^ _0588_;
assign _0590_ = _0589_ ^ _0584_;
assign _0591_ = _0590_ & _0586_;
assign _0592_ = _0591_ ^ _0584_;
assign _0593_ = ~_0592_;
assign _0594_ = _0592_ ^ _0579_;
assign _0595_ = _0592_ ^ _0578_;
assign _0596_ = _0595_ & _0594_;
assign _0597_ = _0596_ ^ _0593_;
assign _0599_ = _0596_ ^ _0592_;
assign _0600_ = _0554_ ^ _0516_;
assign _0601_ = _0600_ ^ _0599_;
assign _0602_ = _0558_ ^ _0418_;
assign _0603_ = _0602_ ^ _0597_;
assign _0604_ = _0603_ & _0601_;
assign _0605_ = _0604_ ^ _0597_;
assign _0606_ = _0605_ & _0580_;
assign out_array_26 = _0606_ ^ _0578_;
assign _0607__neg = _0589_ ^ _0585_;
assign _0607_ = ~_0607__neg;
assign _0609_ = _0607_ & _0605_;
assign out_array_25 = _0609_ ^ _0589_;
assign _0610__neg = _0583_ ^ _0581_;
assign _0610_ = ~_0610__neg;
assign _0611_ = _0610_ & _0605_;
assign out_array_24 = _0611_ ^ _0583_;
assign _0612_ = ~_0579_;
assign out_array_30 = _0606_ ^ _0612_;
assign _0613_ = ~_0585_;
assign out_array_29 = _0609_ ^ _0613_;
assign _0614_ = ~_0581_;
assign out_array_28 = _0611_ ^ _0614_;
assign _0616_ = ~_0602_;
assign _0617_ = _0602_ ^ _0600_;
assign _0618_ = _0617_ & _0605_;
assign out_array_27 = _0618_ ^ _0616_;
assign _0619_ = ~_0555_;
assign out_array_23 = _0575_ ^ _0619_;
assign _0620_ = ~_0600_;
assign out_array_31 = _0618_ ^ _0620_;
assign _0621_ = _0290_ ^ _0253_;
assign _0623_ = ~_0351_;
assign _0624_ = _0388_ ^ _0623_;
assign _0625__neg = _0624_ ^ _0621_;
assign _0625_ = ~_0625__neg;
assign _0626_ = ~_0359_;
assign _0627_ = _0392_ ^ _0626_;
assign _0628_ = _0396_ ^ _0261_;
assign _0629_ = _0628_ & _0627_;
assign _0630_ = ~_0368_;
assign _0631_ = _0400_ ^ _0630_;
assign _0632_ = _0631_ ^ _0629_;
assign _0634_ = _0405_ ^ _0270_;
assign _0635_ = _0634_ ^ _0629_;
assign _0636_ = _0635_ & _0632_;
assign _0637_ = _0636_ ^ _0629_;
assign _0638_ = ~_0637_;
assign _0639_ = _0637_ ^ _0624_;
assign _0640_ = _0637_ ^ _0621_;
assign _0641_ = _0640_ & _0639_;
assign _0642_ = _0641_ ^ _0638_;
assign _0643_ = _0641_ ^ _0637_;
assign _0645_ = _0417_ ^ _0384_;
assign _0646_ = _0645_ ^ _0643_;
assign _0647_ = _0421_ ^ _0286_;
assign _0648_ = _0647_ ^ _0642_;
assign _0649_ = _0648_ & _0646_;
assign _0650_ = _0649_ ^ _0642_;
assign _0651_ = _0650_ & _0625_;
assign _0652_ = _0651_ ^ _0621_;
assign _0653_ = _0456_ ^ _0431_;
assign _0654_ = ~_0653_;
assign _0656_ = ~_0461_;
assign _0657_ = _0486_ ^ _0656_;
assign _0658__neg = _0657_ ^ _0653_;
assign _0658_ = ~_0658__neg;
assign _0659_ = ~_0465_;
assign _0660_ = _0490_ ^ _0659_;
assign _0661_ = _0494_ ^ _0435_;
assign _0662_ = _0661_ & _0660_;
assign _0663_ = ~_0470_;
assign _0664_ = _0498_ ^ _0663_;
assign _0665_ = _0664_ ^ _0662_;
assign _0667_ = _0503_ ^ _0440_;
assign _0668_ = _0667_ ^ _0662_;
assign _0669_ = _0668_ & _0665_;
assign _0670_ = _0669_ ^ _0662_;
assign _0671_ = ~_0670_;
assign _0672_ = _0670_ ^ _0657_;
assign _0673_ = _0670_ ^ _0653_;
assign _0674_ = _0673_ & _0672_;
assign _0675_ = _0674_ ^ _0671_;
assign _0676_ = _0674_ ^ _0670_;
assign _0678_ = _0515_ ^ _0482_;
assign _0679_ = _0678_ ^ _0676_;
assign _0680_ = _0519_ ^ _0452_;
assign _0681_ = _0680_ ^ _0675_;
assign _0682_ = _0681_ & _0679_;
assign _0683_ = _0682_ ^ _0675_;
assign _0684_ = _0683_ & _0658_;
assign _0685_ = _0684_ ^ _0654_;
assign _0686__neg = _0685_ ^ _0652_;
assign _0686_ = ~_0686__neg;
assign _0687_ = ~_0661_;
assign _0689__neg = _0661_ ^ _0660_;
assign _0689_ = ~_0689__neg;
assign _0690_ = _0689_ & _0683_;
assign _0691_ = _0690_ ^ _0687_;
assign _0692__neg = _0628_ ^ _0627_;
assign _0692_ = ~_0692__neg;
assign _0693_ = _0692_ & _0650_;
assign _0694_ = _0693_ ^ _0628_;
assign _0695_ = _0694_ & _0691_;
assign _0696_ = ~_0667_;
assign _0697__neg = _0667_ ^ _0664_;
assign _0697_ = ~_0697__neg;
assign _0698_ = _0697_ & _0683_;
assign _0700_ = _0698_ ^ _0696_;
assign _0701_ = _0700_ ^ _0695_;
assign _0702__neg = _0634_ ^ _0631_;
assign _0702_ = ~_0702__neg;
assign _0703_ = _0702_ & _0650_;
assign _0704_ = _0703_ ^ _0634_;
assign _0705_ = _0704_ ^ _0695_;
assign _0706_ = _0705_ & _0701_;
assign _0707_ = _0706_ ^ _0695_;
assign _0708_ = ~_0707_;
assign _0709_ = _0707_ ^ _0685_;
assign _0711_ = _0707_ ^ _0652_;
assign _0712_ = _0711_ & _0709_;
assign _0713_ = _0712_ ^ _0708_;
assign _0714_ = _0712_ ^ _0707_;
assign _0715_ = _0680_ ^ _0678_;
assign _0716_ = _0715_ & _0683_;
assign _0717_ = _0716_ ^ _0680_;
assign _0718_ = _0717_ ^ _0714_;
assign _0719_ = _0647_ ^ _0645_;
assign _0720_ = _0719_ & _0650_;
assign _0722_ = _0720_ ^ _0647_;
assign _0723_ = _0722_ ^ _0713_;
assign _0724_ = _0723_ & _0718_;
assign _0725_ = _0724_ ^ _0713_;
assign _0726_ = _0725_ & _0686_;
assign out_array_2 = _0726_ ^ _0652_;
assign _0727__neg = _0704_ ^ _0700_;
assign _0727_ = ~_0727__neg;
assign _0728_ = _0727_ & _0725_;
assign out_array_1 = _0728_ ^ _0704_;
assign _0729__neg = _0694_ ^ _0691_;
assign _0729_ = ~_0729__neg;
assign _0731_ = _0729_ & _0725_;
assign out_array_0 = _0731_ ^ _0694_;
assign _0732_ = ~_0685_;
assign out_array_6 = _0726_ ^ _0732_;
assign _0733_ = ~_0700_;
assign out_array_5 = _0728_ ^ _0733_;
assign _0734_ = ~_0691_;
assign out_array_4 = _0731_ ^ _0734_;
assign _0735_ = ~_0722_;
assign _0736_ = _0722_ ^ _0717_;
assign _0738_ = _0736_ & _0725_;
assign out_array_3 = _0738_ ^ _0735_;
assign _0739_ = ~_0624_;
assign _0740_ = _0651_ ^ _0739_;
assign _0741_ = _0684_ ^ _0657_;
assign _0742__neg = _0741_ ^ _0740_;
assign _0742_ = ~_0742__neg;
assign _0743_ = _0690_ ^ _0660_;
assign _0744_ = ~_0627_;
assign _0745_ = _0693_ ^ _0744_;
assign _0746_ = _0745_ & _0743_;
assign _0748_ = _0698_ ^ _0664_;
assign _0749_ = _0748_ ^ _0746_;
assign _0750_ = ~_0631_;
assign _0751_ = _0703_ ^ _0750_;
assign _0752_ = _0751_ ^ _0746_;
assign _0753_ = _0752_ & _0749_;
assign _0754_ = _0753_ ^ _0746_;
assign _0755_ = ~_0754_;
assign _0756_ = _0754_ ^ _0741_;
assign _0757_ = _0754_ ^ _0740_;
assign _0759_ = _0757_ & _0756_;
assign _0760_ = _0759_ ^ _0755_;
assign _0761_ = _0759_ ^ _0754_;
assign _0762_ = _0716_ ^ _0678_;
assign _0763_ = _0762_ ^ _0761_;
assign _0764_ = _0720_ ^ _0645_;
assign _0765_ = _0764_ ^ _0760_;
assign _0766_ = _0765_ & _0763_;
assign _0767_ = _0766_ ^ _0760_;
assign _0768_ = _0767_ & _0742_;
assign out_array_10 = _0768_ ^ _0740_;
assign _0770__neg = _0751_ ^ _0748_;
assign _0770_ = ~_0770__neg;
assign _0771_ = _0770_ & _0767_;
assign out_array_9 = _0771_ ^ _0751_;
assign _0772__neg = _0745_ ^ _0743_;
assign _0772_ = ~_0772__neg;
assign _0773_ = _0772_ & _0767_;
assign out_array_8 = _0773_ ^ _0745_;
assign _0774_ = ~_0741_;
assign out_array_14 = _0768_ ^ _0774_;
assign _0775_ = ~_0748_;
assign out_array_13 = _0771_ ^ _0775_;
assign _0777_ = ~_0743_;
assign out_array_12 = _0773_ ^ _0777_;
assign _0778_ = ~_0764_;
assign _0779_ = _0764_ ^ _0762_;
assign _0780_ = _0779_ & _0767_;
assign out_array_11 = _0780_ ^ _0778_;
assign _0781_ = ~_0717_;
assign out_array_7 = _0738_ ^ _0781_;
assign _0782_ = ~_0762_;
assign out_array_15 = _0780_ ^ _0782_;
endmodule
