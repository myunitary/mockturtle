module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 ;
  assign n188 = x132 & x133 ;
  assign n148 = ~x130 & ~x131 ;
  assign n407 = x78 ^ x77 ;
  assign n408 = x128 & n407 ;
  assign n409 = n408 ^ x78 ;
  assign n404 = x80 ^ x79 ;
  assign n405 = x128 & n404 ;
  assign n406 = n405 ^ x80 ;
  assign n410 = n409 ^ n406 ;
  assign n411 = x129 & n410 ;
  assign n412 = n411 ^ n406 ;
  assign n413 = n148 & n412 ;
  assign n137 = x130 & ~x131 ;
  assign n397 = x74 ^ x73 ;
  assign n398 = x128 & n397 ;
  assign n399 = n398 ^ x74 ;
  assign n394 = x76 ^ x75 ;
  assign n395 = x128 & n394 ;
  assign n396 = n395 ^ x76 ;
  assign n400 = n399 ^ n396 ;
  assign n401 = x129 & n400 ;
  assign n402 = n401 ^ n396 ;
  assign n403 = n137 & n402 ;
  assign n414 = n413 ^ n403 ;
  assign n171 = x130 & x131 ;
  assign n428 = x66 ^ x65 ;
  assign n429 = x128 & n428 ;
  assign n430 = n429 ^ x66 ;
  assign n425 = x68 ^ x67 ;
  assign n426 = x128 & n425 ;
  assign n427 = n426 ^ x68 ;
  assign n431 = n430 ^ n427 ;
  assign n432 = x129 & n431 ;
  assign n433 = n432 ^ n427 ;
  assign n434 = n171 & n433 ;
  assign n160 = ~x130 & x131 ;
  assign n418 = x70 ^ x69 ;
  assign n419 = x128 & n418 ;
  assign n420 = n419 ^ x70 ;
  assign n415 = x72 ^ x71 ;
  assign n416 = x128 & n415 ;
  assign n417 = n416 ^ x72 ;
  assign n421 = n420 ^ n417 ;
  assign n422 = x129 & n421 ;
  assign n423 = n422 ^ n417 ;
  assign n424 = n160 & n423 ;
  assign n435 = n434 ^ n424 ;
  assign n436 = n414 & n435 ;
  assign n437 = n436 ^ n414 ;
  assign n438 = n437 ^ n435 ;
  assign n439 = n188 & n438 ;
  assign n136 = ~x132 & x133 ;
  assign n360 = x94 ^ x93 ;
  assign n361 = x128 & n360 ;
  assign n362 = n361 ^ x94 ;
  assign n357 = x96 ^ x95 ;
  assign n358 = x128 & n357 ;
  assign n359 = n358 ^ x96 ;
  assign n363 = n362 ^ n359 ;
  assign n364 = x129 & n363 ;
  assign n365 = n364 ^ n359 ;
  assign n366 = n148 & n365 ;
  assign n350 = x90 ^ x89 ;
  assign n351 = x128 & n350 ;
  assign n352 = n351 ^ x90 ;
  assign n347 = x92 ^ x91 ;
  assign n348 = x128 & n347 ;
  assign n349 = n348 ^ x92 ;
  assign n353 = n352 ^ n349 ;
  assign n354 = x129 & n353 ;
  assign n355 = n354 ^ n349 ;
  assign n356 = n137 & n355 ;
  assign n367 = n366 ^ n356 ;
  assign n381 = x82 ^ x81 ;
  assign n382 = x128 & n381 ;
  assign n383 = n382 ^ x82 ;
  assign n378 = x84 ^ x83 ;
  assign n379 = x128 & n378 ;
  assign n380 = n379 ^ x84 ;
  assign n384 = n383 ^ n380 ;
  assign n385 = x129 & n384 ;
  assign n386 = n385 ^ n380 ;
  assign n387 = n171 & n386 ;
  assign n371 = x86 ^ x85 ;
  assign n372 = x128 & n371 ;
  assign n373 = n372 ^ x86 ;
  assign n368 = x88 ^ x87 ;
  assign n369 = x128 & n368 ;
  assign n370 = n369 ^ x88 ;
  assign n374 = n373 ^ n370 ;
  assign n375 = x129 & n374 ;
  assign n376 = n375 ^ n370 ;
  assign n377 = n160 & n376 ;
  assign n388 = n387 ^ n377 ;
  assign n389 = n367 & n388 ;
  assign n390 = n389 ^ n367 ;
  assign n391 = n390 ^ n388 ;
  assign n392 = n136 & ~n391 ;
  assign n393 = n392 ^ n136 ;
  assign n440 = n439 ^ n393 ;
  assign n236 = ~x132 & ~x133 ;
  assign n502 = x126 ^ x125 ;
  assign n503 = x128 & n502 ;
  assign n504 = n503 ^ x126 ;
  assign n498 = x127 ^ x0 ;
  assign n499 = x128 & n498 ;
  assign n500 = n499 ^ n498 ;
  assign n501 = n500 ^ x127 ;
  assign n505 = n504 ^ n501 ;
  assign n506 = x129 & n505 ;
  assign n507 = n506 ^ n501 ;
  assign n508 = n148 & n507 ;
  assign n491 = x122 ^ x121 ;
  assign n492 = x128 & n491 ;
  assign n493 = n492 ^ x122 ;
  assign n488 = x124 ^ x123 ;
  assign n489 = x128 & n488 ;
  assign n490 = n489 ^ x124 ;
  assign n494 = n493 ^ n490 ;
  assign n495 = x129 & n494 ;
  assign n496 = n495 ^ n490 ;
  assign n497 = n137 & n496 ;
  assign n509 = n508 ^ n497 ;
  assign n523 = x114 ^ x113 ;
  assign n524 = x128 & n523 ;
  assign n525 = n524 ^ x114 ;
  assign n520 = x116 ^ x115 ;
  assign n521 = x128 & n520 ;
  assign n522 = n521 ^ x116 ;
  assign n526 = n525 ^ n522 ;
  assign n527 = x129 & n526 ;
  assign n528 = n527 ^ n522 ;
  assign n529 = n171 & n528 ;
  assign n513 = x118 ^ x117 ;
  assign n514 = x128 & n513 ;
  assign n515 = n514 ^ x118 ;
  assign n510 = x120 ^ x119 ;
  assign n511 = x128 & n510 ;
  assign n512 = n511 ^ x120 ;
  assign n516 = n515 ^ n512 ;
  assign n517 = x129 & n516 ;
  assign n518 = n517 ^ n512 ;
  assign n519 = n160 & n518 ;
  assign n530 = n529 ^ n519 ;
  assign n531 = n509 & n530 ;
  assign n532 = n531 ^ n509 ;
  assign n533 = n532 ^ n530 ;
  assign n534 = n236 & n533 ;
  assign n314 = x132 & ~x133 ;
  assign n454 = x110 ^ x109 ;
  assign n455 = x128 & n454 ;
  assign n456 = n455 ^ x110 ;
  assign n451 = x112 ^ x111 ;
  assign n452 = x128 & n451 ;
  assign n453 = n452 ^ x112 ;
  assign n457 = n456 ^ n453 ;
  assign n458 = x129 & n457 ;
  assign n459 = n458 ^ n453 ;
  assign n460 = n148 & n459 ;
  assign n444 = x106 ^ x105 ;
  assign n445 = x128 & n444 ;
  assign n446 = n445 ^ x106 ;
  assign n441 = x108 ^ x107 ;
  assign n442 = x128 & n441 ;
  assign n443 = n442 ^ x108 ;
  assign n447 = n446 ^ n443 ;
  assign n448 = x129 & n447 ;
  assign n449 = n448 ^ n443 ;
  assign n450 = n137 & n449 ;
  assign n461 = n460 ^ n450 ;
  assign n475 = x98 ^ x97 ;
  assign n476 = x128 & n475 ;
  assign n477 = n476 ^ x98 ;
  assign n472 = x100 ^ x99 ;
  assign n473 = x128 & n472 ;
  assign n474 = n473 ^ x100 ;
  assign n478 = n477 ^ n474 ;
  assign n479 = x129 & n478 ;
  assign n480 = n479 ^ n474 ;
  assign n481 = n171 & n480 ;
  assign n465 = x102 ^ x101 ;
  assign n466 = x128 & n465 ;
  assign n467 = n466 ^ x102 ;
  assign n462 = x104 ^ x103 ;
  assign n463 = x128 & n462 ;
  assign n464 = n463 ^ x104 ;
  assign n468 = n467 ^ n464 ;
  assign n469 = x129 & n468 ;
  assign n470 = n469 ^ n464 ;
  assign n471 = n160 & n470 ;
  assign n482 = n481 ^ n471 ;
  assign n483 = n461 & n482 ;
  assign n484 = n483 ^ n461 ;
  assign n485 = n484 ^ n482 ;
  assign n486 = n314 & ~n485 ;
  assign n487 = n486 ^ n314 ;
  assign n535 = n534 ^ n487 ;
  assign n536 = n440 & n535 ;
  assign n537 = n536 ^ n440 ;
  assign n538 = n537 ^ n535 ;
  assign n202 = x14 ^ x13 ;
  assign n203 = x128 & n202 ;
  assign n204 = n203 ^ x14 ;
  assign n199 = x16 ^ x15 ;
  assign n200 = x128 & n199 ;
  assign n201 = n200 ^ x16 ;
  assign n205 = n204 ^ n201 ;
  assign n206 = x129 & n205 ;
  assign n207 = n206 ^ n201 ;
  assign n208 = n148 & n207 ;
  assign n192 = x10 ^ x9 ;
  assign n193 = x128 & n192 ;
  assign n194 = n193 ^ x10 ;
  assign n189 = x12 ^ x11 ;
  assign n190 = x128 & n189 ;
  assign n191 = n190 ^ x12 ;
  assign n195 = n194 ^ n191 ;
  assign n196 = x129 & n195 ;
  assign n197 = n196 ^ n191 ;
  assign n198 = n137 & n197 ;
  assign n209 = n208 ^ n198 ;
  assign n223 = x2 ^ x1 ;
  assign n224 = x128 & n223 ;
  assign n225 = n224 ^ x2 ;
  assign n220 = x4 ^ x3 ;
  assign n221 = x128 & n220 ;
  assign n222 = n221 ^ x4 ;
  assign n226 = n225 ^ n222 ;
  assign n227 = x129 & n226 ;
  assign n228 = n227 ^ n222 ;
  assign n229 = n171 & n228 ;
  assign n213 = x6 ^ x5 ;
  assign n214 = x128 & n213 ;
  assign n215 = n214 ^ x6 ;
  assign n210 = x8 ^ x7 ;
  assign n211 = x128 & n210 ;
  assign n212 = n211 ^ x8 ;
  assign n216 = n215 ^ n212 ;
  assign n217 = x129 & n216 ;
  assign n218 = n217 ^ n212 ;
  assign n219 = n160 & n218 ;
  assign n230 = n229 ^ n219 ;
  assign n231 = n209 & n230 ;
  assign n232 = n231 ^ n209 ;
  assign n233 = n232 ^ n230 ;
  assign n234 = n188 & n233 ;
  assign n152 = x30 ^ x29 ;
  assign n153 = x128 & n152 ;
  assign n154 = n153 ^ x30 ;
  assign n149 = x32 ^ x31 ;
  assign n150 = x128 & n149 ;
  assign n151 = n150 ^ x32 ;
  assign n155 = n154 ^ n151 ;
  assign n156 = x129 & n155 ;
  assign n157 = n156 ^ n151 ;
  assign n158 = n148 & n157 ;
  assign n141 = x26 ^ x25 ;
  assign n142 = x128 & n141 ;
  assign n143 = n142 ^ x26 ;
  assign n138 = x28 ^ x27 ;
  assign n139 = x128 & n138 ;
  assign n140 = n139 ^ x28 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = x129 & n144 ;
  assign n146 = n145 ^ n140 ;
  assign n147 = n137 & n146 ;
  assign n159 = n158 ^ n147 ;
  assign n175 = x18 ^ x17 ;
  assign n176 = x128 & n175 ;
  assign n177 = n176 ^ x18 ;
  assign n172 = x20 ^ x19 ;
  assign n173 = x128 & n172 ;
  assign n174 = n173 ^ x20 ;
  assign n178 = n177 ^ n174 ;
  assign n179 = x129 & n178 ;
  assign n180 = n179 ^ n174 ;
  assign n181 = n171 & n180 ;
  assign n164 = x22 ^ x21 ;
  assign n165 = x128 & n164 ;
  assign n166 = n165 ^ x22 ;
  assign n161 = x24 ^ x23 ;
  assign n162 = x128 & n161 ;
  assign n163 = n162 ^ x24 ;
  assign n167 = n166 ^ n163 ;
  assign n168 = x129 & n167 ;
  assign n169 = n168 ^ n163 ;
  assign n170 = n160 & n169 ;
  assign n182 = n181 ^ n170 ;
  assign n183 = n159 & n182 ;
  assign n184 = n183 ^ n159 ;
  assign n185 = n184 ^ n182 ;
  assign n186 = n136 & ~n185 ;
  assign n187 = n186 ^ n136 ;
  assign n235 = n234 ^ n187 ;
  assign n250 = x62 ^ x61 ;
  assign n251 = x128 & n250 ;
  assign n252 = n251 ^ x62 ;
  assign n247 = x64 ^ x63 ;
  assign n248 = x128 & n247 ;
  assign n249 = n248 ^ x64 ;
  assign n253 = n252 ^ n249 ;
  assign n254 = x129 & n253 ;
  assign n255 = n254 ^ n249 ;
  assign n256 = n148 & n255 ;
  assign n240 = x58 ^ x57 ;
  assign n241 = x128 & n240 ;
  assign n242 = n241 ^ x58 ;
  assign n237 = x60 ^ x59 ;
  assign n238 = x128 & n237 ;
  assign n239 = n238 ^ x60 ;
  assign n243 = n242 ^ n239 ;
  assign n244 = x129 & n243 ;
  assign n245 = n244 ^ n239 ;
  assign n246 = n137 & n245 ;
  assign n257 = n256 ^ n246 ;
  assign n271 = x50 ^ x49 ;
  assign n272 = x128 & n271 ;
  assign n273 = n272 ^ x50 ;
  assign n268 = x52 ^ x51 ;
  assign n269 = x128 & n268 ;
  assign n270 = n269 ^ x52 ;
  assign n274 = n273 ^ n270 ;
  assign n275 = x129 & n274 ;
  assign n276 = n275 ^ n270 ;
  assign n277 = n171 & n276 ;
  assign n261 = x54 ^ x53 ;
  assign n262 = x128 & n261 ;
  assign n263 = n262 ^ x54 ;
  assign n258 = x56 ^ x55 ;
  assign n259 = x128 & n258 ;
  assign n260 = n259 ^ x56 ;
  assign n264 = n263 ^ n260 ;
  assign n265 = x129 & n264 ;
  assign n266 = n265 ^ n260 ;
  assign n267 = n160 & n266 ;
  assign n278 = n277 ^ n267 ;
  assign n279 = n257 & n278 ;
  assign n280 = n279 ^ n257 ;
  assign n281 = n280 ^ n278 ;
  assign n282 = n236 & ~n281 ;
  assign n283 = n282 ^ n236 ;
  assign n306 = x34 ^ x33 ;
  assign n307 = x128 & n306 ;
  assign n308 = n307 ^ x34 ;
  assign n303 = x36 ^ x35 ;
  assign n304 = x128 & n303 ;
  assign n305 = n304 ^ x36 ;
  assign n309 = n308 ^ n305 ;
  assign n310 = x129 & n309 ;
  assign n311 = n310 ^ n305 ;
  assign n312 = n171 & n311 ;
  assign n286 = x39 & x128 ;
  assign n284 = x38 & x128 ;
  assign n285 = n284 ^ x38 ;
  assign n287 = n286 ^ n285 ;
  assign n288 = x129 & n287 ;
  assign n289 = n288 ^ n287 ;
  assign n290 = n289 ^ n285 ;
  assign n293 = x37 & x128 ;
  assign n291 = x40 & x128 ;
  assign n292 = n291 ^ x40 ;
  assign n294 = n293 ^ n292 ;
  assign n295 = x129 & n294 ;
  assign n296 = n295 ^ n292 ;
  assign n297 = n290 & n296 ;
  assign n298 = n297 ^ n290 ;
  assign n299 = n298 ^ n296 ;
  assign n300 = n160 & n299 ;
  assign n301 = n300 ^ n160 ;
  assign n302 = n301 ^ n160 ;
  assign n313 = n312 ^ n302 ;
  assign n328 = x46 ^ x45 ;
  assign n329 = x128 & n328 ;
  assign n330 = n329 ^ x46 ;
  assign n325 = x48 ^ x47 ;
  assign n326 = x128 & n325 ;
  assign n327 = n326 ^ x48 ;
  assign n331 = n330 ^ n327 ;
  assign n332 = x129 & n331 ;
  assign n333 = n332 ^ n327 ;
  assign n334 = n148 & n333 ;
  assign n318 = x42 ^ x41 ;
  assign n319 = x128 & n318 ;
  assign n320 = n319 ^ x42 ;
  assign n315 = x44 ^ x43 ;
  assign n316 = x128 & n315 ;
  assign n317 = n316 ^ x44 ;
  assign n321 = n320 ^ n317 ;
  assign n322 = x129 & n321 ;
  assign n323 = n322 ^ n317 ;
  assign n324 = n137 & n323 ;
  assign n335 = n334 ^ n324 ;
  assign n336 = n314 & n335 ;
  assign n337 = n336 ^ n314 ;
  assign n338 = n313 & n337 ;
  assign n339 = n338 ^ n337 ;
  assign n340 = n339 ^ n314 ;
  assign n341 = n283 & n340 ;
  assign n342 = n341 ^ n283 ;
  assign n343 = n342 ^ n340 ;
  assign n344 = n235 & n343 ;
  assign n345 = n344 ^ n235 ;
  assign n346 = n345 ^ n343 ;
  assign n539 = n538 ^ n346 ;
  assign n540 = x134 & n539 ;
  assign n541 = n540 ^ n539 ;
  assign n542 = n541 ^ n346 ;
  assign n948 = x80 & x128 ;
  assign n946 = x79 & x128 ;
  assign n947 = n946 ^ x79 ;
  assign n949 = n948 ^ n947 ;
  assign n950 = x129 & n949 ;
  assign n951 = n950 ^ n949 ;
  assign n952 = n951 ^ n947 ;
  assign n955 = x78 & x128 ;
  assign n953 = x81 & x128 ;
  assign n954 = n953 ^ x81 ;
  assign n956 = n955 ^ n954 ;
  assign n957 = x129 & n956 ;
  assign n958 = n957 ^ n954 ;
  assign n959 = n952 & n958 ;
  assign n960 = n959 ^ n952 ;
  assign n961 = n960 ^ n958 ;
  assign n962 = n148 & n961 ;
  assign n929 = x76 & x128 ;
  assign n927 = x75 & x128 ;
  assign n928 = n927 ^ x75 ;
  assign n930 = n929 ^ n928 ;
  assign n931 = x129 & n930 ;
  assign n932 = n931 ^ n930 ;
  assign n933 = n932 ^ n928 ;
  assign n936 = x74 & x128 ;
  assign n934 = x77 & x128 ;
  assign n935 = n934 ^ x77 ;
  assign n937 = n936 ^ n935 ;
  assign n938 = x129 & n937 ;
  assign n939 = n938 ^ n935 ;
  assign n940 = n933 & n939 ;
  assign n941 = n940 ^ n933 ;
  assign n942 = n941 ^ n939 ;
  assign n943 = n137 & n942 ;
  assign n944 = n943 ^ n137 ;
  assign n945 = n944 ^ n137 ;
  assign n963 = n962 ^ n945 ;
  assign n985 = x68 & x128 ;
  assign n983 = x67 & x128 ;
  assign n984 = n983 ^ x67 ;
  assign n986 = n985 ^ n984 ;
  assign n987 = x129 & n986 ;
  assign n988 = n987 ^ n986 ;
  assign n989 = n988 ^ n984 ;
  assign n992 = x66 & x128 ;
  assign n990 = x69 & x128 ;
  assign n991 = n990 ^ x69 ;
  assign n993 = n992 ^ n991 ;
  assign n994 = x129 & n993 ;
  assign n995 = n994 ^ n991 ;
  assign n996 = n989 & n995 ;
  assign n997 = n996 ^ n989 ;
  assign n998 = n997 ^ n995 ;
  assign n999 = n171 & n998 ;
  assign n966 = x72 & x128 ;
  assign n964 = x71 & x128 ;
  assign n965 = n964 ^ x71 ;
  assign n967 = n966 ^ n965 ;
  assign n968 = x129 & n967 ;
  assign n969 = n968 ^ n967 ;
  assign n970 = n969 ^ n965 ;
  assign n973 = x70 & x128 ;
  assign n971 = x73 & x128 ;
  assign n972 = n971 ^ x73 ;
  assign n974 = n973 ^ n972 ;
  assign n975 = x129 & n974 ;
  assign n976 = n975 ^ n972 ;
  assign n977 = n970 & n976 ;
  assign n978 = n977 ^ n970 ;
  assign n979 = n978 ^ n976 ;
  assign n980 = n160 & n979 ;
  assign n981 = n980 ^ n160 ;
  assign n982 = n981 ^ n160 ;
  assign n1000 = n999 ^ n982 ;
  assign n1001 = n963 & n1000 ;
  assign n1002 = n1001 ^ n963 ;
  assign n1003 = n1002 ^ n1000 ;
  assign n1004 = n188 & n1003 ;
  assign n869 = x96 & x128 ;
  assign n867 = x95 & x128 ;
  assign n868 = n867 ^ x95 ;
  assign n870 = n869 ^ n868 ;
  assign n871 = x129 & n870 ;
  assign n872 = n871 ^ n870 ;
  assign n873 = n872 ^ n868 ;
  assign n876 = x94 & x128 ;
  assign n874 = x97 & x128 ;
  assign n875 = n874 ^ x97 ;
  assign n877 = n876 ^ n875 ;
  assign n878 = x129 & n877 ;
  assign n879 = n878 ^ n875 ;
  assign n880 = n873 & n879 ;
  assign n881 = n880 ^ n873 ;
  assign n882 = n881 ^ n879 ;
  assign n883 = n148 & n882 ;
  assign n850 = x92 & x128 ;
  assign n848 = x91 & x128 ;
  assign n849 = n848 ^ x91 ;
  assign n851 = n850 ^ n849 ;
  assign n852 = x129 & n851 ;
  assign n853 = n852 ^ n851 ;
  assign n854 = n853 ^ n849 ;
  assign n857 = x90 & x128 ;
  assign n855 = x93 & x128 ;
  assign n856 = n855 ^ x93 ;
  assign n858 = n857 ^ n856 ;
  assign n859 = x129 & n858 ;
  assign n860 = n859 ^ n856 ;
  assign n861 = n854 & n860 ;
  assign n862 = n861 ^ n854 ;
  assign n863 = n862 ^ n860 ;
  assign n864 = n137 & n863 ;
  assign n865 = n864 ^ n137 ;
  assign n866 = n865 ^ n137 ;
  assign n884 = n883 ^ n866 ;
  assign n906 = x84 & x128 ;
  assign n904 = x83 & x128 ;
  assign n905 = n904 ^ x83 ;
  assign n907 = n906 ^ n905 ;
  assign n908 = x129 & n907 ;
  assign n909 = n908 ^ n907 ;
  assign n910 = n909 ^ n905 ;
  assign n913 = x82 & x128 ;
  assign n911 = x85 & x128 ;
  assign n912 = n911 ^ x85 ;
  assign n914 = n913 ^ n912 ;
  assign n915 = x129 & n914 ;
  assign n916 = n915 ^ n912 ;
  assign n917 = n910 & n916 ;
  assign n918 = n917 ^ n910 ;
  assign n919 = n918 ^ n916 ;
  assign n920 = n171 & n919 ;
  assign n887 = x88 & x128 ;
  assign n885 = x87 & x128 ;
  assign n886 = n885 ^ x87 ;
  assign n888 = n887 ^ n886 ;
  assign n889 = x129 & n888 ;
  assign n890 = n889 ^ n888 ;
  assign n891 = n890 ^ n886 ;
  assign n894 = x86 & x128 ;
  assign n892 = x89 & x128 ;
  assign n893 = n892 ^ x89 ;
  assign n895 = n894 ^ n893 ;
  assign n896 = x129 & n895 ;
  assign n897 = n896 ^ n893 ;
  assign n898 = n891 & n897 ;
  assign n899 = n898 ^ n891 ;
  assign n900 = n899 ^ n897 ;
  assign n901 = n160 & n900 ;
  assign n902 = n901 ^ n160 ;
  assign n903 = n902 ^ n160 ;
  assign n921 = n920 ^ n903 ;
  assign n922 = n884 & n921 ;
  assign n923 = n922 ^ n884 ;
  assign n924 = n923 ^ n921 ;
  assign n925 = n136 & ~n924 ;
  assign n926 = n925 ^ n136 ;
  assign n1005 = n1004 ^ n926 ;
  assign n1106 = x0 & x128 ;
  assign n1104 = x127 & x128 ;
  assign n1105 = n1104 ^ x127 ;
  assign n1107 = n1106 ^ n1105 ;
  assign n1108 = x129 & n1107 ;
  assign n1109 = n1108 ^ n1107 ;
  assign n1110 = n1109 ^ n1105 ;
  assign n1113 = x126 & x128 ;
  assign n1111 = x1 & x128 ;
  assign n1112 = n1111 ^ x1 ;
  assign n1114 = n1113 ^ n1112 ;
  assign n1115 = x129 & n1114 ;
  assign n1116 = n1115 ^ n1112 ;
  assign n1117 = n1110 & n1116 ;
  assign n1118 = n1117 ^ n1110 ;
  assign n1119 = n1118 ^ n1116 ;
  assign n1120 = n148 & n1119 ;
  assign n1087 = x124 & x128 ;
  assign n1085 = x123 & x128 ;
  assign n1086 = n1085 ^ x123 ;
  assign n1088 = n1087 ^ n1086 ;
  assign n1089 = x129 & n1088 ;
  assign n1090 = n1089 ^ n1088 ;
  assign n1091 = n1090 ^ n1086 ;
  assign n1094 = x122 & x128 ;
  assign n1092 = x125 & x128 ;
  assign n1093 = n1092 ^ x125 ;
  assign n1095 = n1094 ^ n1093 ;
  assign n1096 = x129 & n1095 ;
  assign n1097 = n1096 ^ n1093 ;
  assign n1098 = n1091 & n1097 ;
  assign n1099 = n1098 ^ n1091 ;
  assign n1100 = n1099 ^ n1097 ;
  assign n1101 = n137 & n1100 ;
  assign n1102 = n1101 ^ n137 ;
  assign n1103 = n1102 ^ n137 ;
  assign n1121 = n1120 ^ n1103 ;
  assign n1143 = x116 & x128 ;
  assign n1141 = x115 & x128 ;
  assign n1142 = n1141 ^ x115 ;
  assign n1144 = n1143 ^ n1142 ;
  assign n1145 = x129 & n1144 ;
  assign n1146 = n1145 ^ n1144 ;
  assign n1147 = n1146 ^ n1142 ;
  assign n1150 = x114 & x128 ;
  assign n1148 = x117 & x128 ;
  assign n1149 = n1148 ^ x117 ;
  assign n1151 = n1150 ^ n1149 ;
  assign n1152 = x129 & n1151 ;
  assign n1153 = n1152 ^ n1149 ;
  assign n1154 = n1147 & n1153 ;
  assign n1155 = n1154 ^ n1147 ;
  assign n1156 = n1155 ^ n1153 ;
  assign n1157 = n171 & n1156 ;
  assign n1124 = x120 & x128 ;
  assign n1122 = x119 & x128 ;
  assign n1123 = n1122 ^ x119 ;
  assign n1125 = n1124 ^ n1123 ;
  assign n1126 = x129 & n1125 ;
  assign n1127 = n1126 ^ n1125 ;
  assign n1128 = n1127 ^ n1123 ;
  assign n1131 = x118 & x128 ;
  assign n1129 = x121 & x128 ;
  assign n1130 = n1129 ^ x121 ;
  assign n1132 = n1131 ^ n1130 ;
  assign n1133 = x129 & n1132 ;
  assign n1134 = n1133 ^ n1130 ;
  assign n1135 = n1128 & n1134 ;
  assign n1136 = n1135 ^ n1128 ;
  assign n1137 = n1136 ^ n1134 ;
  assign n1138 = n160 & n1137 ;
  assign n1139 = n1138 ^ n160 ;
  assign n1140 = n1139 ^ n160 ;
  assign n1158 = n1157 ^ n1140 ;
  assign n1159 = n1121 & n1158 ;
  assign n1160 = n1159 ^ n1121 ;
  assign n1161 = n1160 ^ n1158 ;
  assign n1162 = n236 & n1161 ;
  assign n1027 = x112 & x128 ;
  assign n1025 = x111 & x128 ;
  assign n1026 = n1025 ^ x111 ;
  assign n1028 = n1027 ^ n1026 ;
  assign n1029 = x129 & n1028 ;
  assign n1030 = n1029 ^ n1028 ;
  assign n1031 = n1030 ^ n1026 ;
  assign n1034 = x110 & x128 ;
  assign n1032 = x113 & x128 ;
  assign n1033 = n1032 ^ x113 ;
  assign n1035 = n1034 ^ n1033 ;
  assign n1036 = x129 & n1035 ;
  assign n1037 = n1036 ^ n1033 ;
  assign n1038 = n1031 & n1037 ;
  assign n1039 = n1038 ^ n1031 ;
  assign n1040 = n1039 ^ n1037 ;
  assign n1041 = n148 & n1040 ;
  assign n1008 = x108 & x128 ;
  assign n1006 = x107 & x128 ;
  assign n1007 = n1006 ^ x107 ;
  assign n1009 = n1008 ^ n1007 ;
  assign n1010 = x129 & n1009 ;
  assign n1011 = n1010 ^ n1009 ;
  assign n1012 = n1011 ^ n1007 ;
  assign n1015 = x106 & x128 ;
  assign n1013 = x109 & x128 ;
  assign n1014 = n1013 ^ x109 ;
  assign n1016 = n1015 ^ n1014 ;
  assign n1017 = x129 & n1016 ;
  assign n1018 = n1017 ^ n1014 ;
  assign n1019 = n1012 & n1018 ;
  assign n1020 = n1019 ^ n1012 ;
  assign n1021 = n1020 ^ n1018 ;
  assign n1022 = n137 & n1021 ;
  assign n1023 = n1022 ^ n137 ;
  assign n1024 = n1023 ^ n137 ;
  assign n1042 = n1041 ^ n1024 ;
  assign n1064 = x100 & x128 ;
  assign n1062 = x99 & x128 ;
  assign n1063 = n1062 ^ x99 ;
  assign n1065 = n1064 ^ n1063 ;
  assign n1066 = x129 & n1065 ;
  assign n1067 = n1066 ^ n1065 ;
  assign n1068 = n1067 ^ n1063 ;
  assign n1071 = x98 & x128 ;
  assign n1069 = x101 & x128 ;
  assign n1070 = n1069 ^ x101 ;
  assign n1072 = n1071 ^ n1070 ;
  assign n1073 = x129 & n1072 ;
  assign n1074 = n1073 ^ n1070 ;
  assign n1075 = n1068 & n1074 ;
  assign n1076 = n1075 ^ n1068 ;
  assign n1077 = n1076 ^ n1074 ;
  assign n1078 = n171 & n1077 ;
  assign n1045 = x104 & x128 ;
  assign n1043 = x103 & x128 ;
  assign n1044 = n1043 ^ x103 ;
  assign n1046 = n1045 ^ n1044 ;
  assign n1047 = x129 & n1046 ;
  assign n1048 = n1047 ^ n1046 ;
  assign n1049 = n1048 ^ n1044 ;
  assign n1052 = x102 & x128 ;
  assign n1050 = x105 & x128 ;
  assign n1051 = n1050 ^ x105 ;
  assign n1053 = n1052 ^ n1051 ;
  assign n1054 = x129 & n1053 ;
  assign n1055 = n1054 ^ n1051 ;
  assign n1056 = n1049 & n1055 ;
  assign n1057 = n1056 ^ n1049 ;
  assign n1058 = n1057 ^ n1055 ;
  assign n1059 = n160 & n1058 ;
  assign n1060 = n1059 ^ n160 ;
  assign n1061 = n1060 ^ n160 ;
  assign n1079 = n1078 ^ n1061 ;
  assign n1080 = n1042 & n1079 ;
  assign n1081 = n1080 ^ n1042 ;
  assign n1082 = n1081 ^ n1079 ;
  assign n1083 = n314 & ~n1082 ;
  assign n1084 = n1083 ^ n314 ;
  assign n1163 = n1162 ^ n1084 ;
  assign n1164 = n1005 & n1163 ;
  assign n1165 = n1164 ^ n1005 ;
  assign n1166 = n1165 ^ n1163 ;
  assign n643 = x64 & x128 ;
  assign n641 = x63 & x128 ;
  assign n642 = n641 ^ x63 ;
  assign n644 = n643 ^ n642 ;
  assign n645 = x129 & n644 ;
  assign n646 = n645 ^ n644 ;
  assign n647 = n646 ^ n642 ;
  assign n650 = x62 & x128 ;
  assign n648 = x65 & x128 ;
  assign n649 = n648 ^ x65 ;
  assign n651 = n650 ^ n649 ;
  assign n652 = x129 & n651 ;
  assign n653 = n652 ^ n649 ;
  assign n654 = n647 & n653 ;
  assign n655 = n654 ^ n647 ;
  assign n656 = n655 ^ n653 ;
  assign n657 = n148 & n656 ;
  assign n624 = x60 & x128 ;
  assign n622 = x59 & x128 ;
  assign n623 = n622 ^ x59 ;
  assign n625 = n624 ^ n623 ;
  assign n626 = x129 & n625 ;
  assign n627 = n626 ^ n625 ;
  assign n628 = n627 ^ n623 ;
  assign n631 = x58 & x128 ;
  assign n629 = x61 & x128 ;
  assign n630 = n629 ^ x61 ;
  assign n632 = n631 ^ n630 ;
  assign n633 = x129 & n632 ;
  assign n634 = n633 ^ n630 ;
  assign n635 = n628 & n634 ;
  assign n636 = n635 ^ n628 ;
  assign n637 = n636 ^ n634 ;
  assign n638 = n137 & n637 ;
  assign n639 = n638 ^ n137 ;
  assign n640 = n639 ^ n137 ;
  assign n658 = n657 ^ n640 ;
  assign n680 = x52 & x128 ;
  assign n678 = x51 & x128 ;
  assign n679 = n678 ^ x51 ;
  assign n681 = n680 ^ n679 ;
  assign n682 = x129 & n681 ;
  assign n683 = n682 ^ n681 ;
  assign n684 = n683 ^ n679 ;
  assign n687 = x50 & x128 ;
  assign n685 = x53 & x128 ;
  assign n686 = n685 ^ x53 ;
  assign n688 = n687 ^ n686 ;
  assign n689 = x129 & n688 ;
  assign n690 = n689 ^ n686 ;
  assign n691 = n684 & n690 ;
  assign n692 = n691 ^ n684 ;
  assign n693 = n692 ^ n690 ;
  assign n694 = n171 & n693 ;
  assign n661 = x56 & x128 ;
  assign n659 = x55 & x128 ;
  assign n660 = n659 ^ x55 ;
  assign n662 = n661 ^ n660 ;
  assign n663 = x129 & n662 ;
  assign n664 = n663 ^ n662 ;
  assign n665 = n664 ^ n660 ;
  assign n668 = x54 & x128 ;
  assign n666 = x57 & x128 ;
  assign n667 = n666 ^ x57 ;
  assign n669 = n668 ^ n667 ;
  assign n670 = x129 & n669 ;
  assign n671 = n670 ^ n667 ;
  assign n672 = n665 & n671 ;
  assign n673 = n672 ^ n665 ;
  assign n674 = n673 ^ n671 ;
  assign n675 = n160 & n674 ;
  assign n676 = n675 ^ n160 ;
  assign n677 = n676 ^ n160 ;
  assign n695 = n694 ^ n677 ;
  assign n696 = n658 & n695 ;
  assign n697 = n696 ^ n658 ;
  assign n698 = n697 ^ n695 ;
  assign n699 = n236 & n698 ;
  assign n564 = x16 & x128 ;
  assign n562 = x15 & x128 ;
  assign n563 = n562 ^ x15 ;
  assign n565 = n564 ^ n563 ;
  assign n566 = x129 & n565 ;
  assign n567 = n566 ^ n565 ;
  assign n568 = n567 ^ n563 ;
  assign n571 = x14 & x128 ;
  assign n569 = x17 & x128 ;
  assign n570 = n569 ^ x17 ;
  assign n572 = n571 ^ n570 ;
  assign n573 = x129 & n572 ;
  assign n574 = n573 ^ n570 ;
  assign n575 = n568 & n574 ;
  assign n576 = n575 ^ n568 ;
  assign n577 = n576 ^ n574 ;
  assign n578 = n148 & n577 ;
  assign n545 = x12 & x128 ;
  assign n543 = x11 & x128 ;
  assign n544 = n543 ^ x11 ;
  assign n546 = n545 ^ n544 ;
  assign n547 = x129 & n546 ;
  assign n548 = n547 ^ n546 ;
  assign n549 = n548 ^ n544 ;
  assign n552 = x10 & x128 ;
  assign n550 = x13 & x128 ;
  assign n551 = n550 ^ x13 ;
  assign n553 = n552 ^ n551 ;
  assign n554 = x129 & n553 ;
  assign n555 = n554 ^ n551 ;
  assign n556 = n549 & n555 ;
  assign n557 = n556 ^ n549 ;
  assign n558 = n557 ^ n555 ;
  assign n559 = n137 & n558 ;
  assign n560 = n559 ^ n137 ;
  assign n561 = n560 ^ n137 ;
  assign n579 = n578 ^ n561 ;
  assign n601 = x4 & x128 ;
  assign n599 = x3 & x128 ;
  assign n600 = n599 ^ x3 ;
  assign n602 = n601 ^ n600 ;
  assign n603 = x129 & n602 ;
  assign n604 = n603 ^ n602 ;
  assign n605 = n604 ^ n600 ;
  assign n608 = x2 & x128 ;
  assign n606 = x5 & x128 ;
  assign n607 = n606 ^ x5 ;
  assign n609 = n608 ^ n607 ;
  assign n610 = x129 & n609 ;
  assign n611 = n610 ^ n607 ;
  assign n612 = n605 & n611 ;
  assign n613 = n612 ^ n605 ;
  assign n614 = n613 ^ n611 ;
  assign n615 = n171 & n614 ;
  assign n582 = x8 & x128 ;
  assign n580 = x7 & x128 ;
  assign n581 = n580 ^ x7 ;
  assign n583 = n582 ^ n581 ;
  assign n584 = x129 & n583 ;
  assign n585 = n584 ^ n583 ;
  assign n586 = n585 ^ n581 ;
  assign n589 = x6 & x128 ;
  assign n587 = x9 & x128 ;
  assign n588 = n587 ^ x9 ;
  assign n590 = n589 ^ n588 ;
  assign n591 = x129 & n590 ;
  assign n592 = n591 ^ n588 ;
  assign n593 = n586 & n592 ;
  assign n594 = n593 ^ n586 ;
  assign n595 = n594 ^ n592 ;
  assign n596 = n160 & n595 ;
  assign n597 = n596 ^ n160 ;
  assign n598 = n597 ^ n160 ;
  assign n616 = n615 ^ n598 ;
  assign n617 = n579 & n616 ;
  assign n618 = n617 ^ n579 ;
  assign n619 = n618 ^ n616 ;
  assign n620 = n188 & ~n619 ;
  assign n621 = n620 ^ n188 ;
  assign n700 = n699 ^ n621 ;
  assign n795 = x48 & x128 ;
  assign n793 = x47 & x128 ;
  assign n794 = n793 ^ x47 ;
  assign n796 = n795 ^ n794 ;
  assign n797 = x129 & n796 ;
  assign n798 = n797 ^ n796 ;
  assign n799 = n798 ^ n794 ;
  assign n802 = x46 & x128 ;
  assign n800 = x49 & x128 ;
  assign n801 = n800 ^ x49 ;
  assign n803 = n802 ^ n801 ;
  assign n804 = x129 & n803 ;
  assign n805 = n804 ^ n801 ;
  assign n806 = n799 & n805 ;
  assign n807 = n806 ^ n799 ;
  assign n808 = n807 ^ n805 ;
  assign n809 = n148 & n808 ;
  assign n783 = x43 ^ x42 ;
  assign n784 = x128 & n783 ;
  assign n785 = n784 ^ x43 ;
  assign n780 = x45 ^ x44 ;
  assign n781 = x128 & n780 ;
  assign n782 = n781 ^ x45 ;
  assign n786 = n785 ^ n782 ;
  assign n787 = x129 & n786 ;
  assign n788 = n787 ^ x129 ;
  assign n789 = n788 ^ x129 ;
  assign n790 = n789 ^ n782 ;
  assign n791 = n137 & ~n790 ;
  assign n792 = n791 ^ n137 ;
  assign n810 = n809 ^ n792 ;
  assign n825 = x36 & x128 ;
  assign n823 = x35 & x128 ;
  assign n824 = n823 ^ x35 ;
  assign n826 = n825 ^ n824 ;
  assign n827 = x129 & n826 ;
  assign n828 = n827 ^ n826 ;
  assign n829 = n828 ^ n824 ;
  assign n831 = x34 & x128 ;
  assign n830 = n293 ^ x37 ;
  assign n832 = n831 ^ n830 ;
  assign n833 = x129 & n832 ;
  assign n834 = n833 ^ n830 ;
  assign n835 = n829 & n834 ;
  assign n836 = n835 ^ n829 ;
  assign n837 = n836 ^ n834 ;
  assign n838 = n171 & n837 ;
  assign n814 = x41 ^ x40 ;
  assign n815 = x128 & n814 ;
  assign n816 = n815 ^ x41 ;
  assign n811 = x39 ^ x38 ;
  assign n812 = x128 & n811 ;
  assign n813 = n812 ^ x39 ;
  assign n817 = n816 ^ n813 ;
  assign n818 = x129 & n817 ;
  assign n819 = n818 ^ n817 ;
  assign n820 = n819 ^ n813 ;
  assign n821 = n160 & ~n820 ;
  assign n822 = n821 ^ n160 ;
  assign n839 = n838 ^ n822 ;
  assign n840 = n810 & n839 ;
  assign n841 = n840 ^ n810 ;
  assign n842 = n841 ^ n839 ;
  assign n843 = n314 & n842 ;
  assign n722 = x32 & x128 ;
  assign n720 = x31 & x128 ;
  assign n721 = n720 ^ x31 ;
  assign n723 = n722 ^ n721 ;
  assign n724 = x129 & n723 ;
  assign n725 = n724 ^ n723 ;
  assign n726 = n725 ^ n721 ;
  assign n729 = x30 & x128 ;
  assign n727 = x33 & x128 ;
  assign n728 = n727 ^ x33 ;
  assign n730 = n729 ^ n728 ;
  assign n731 = x129 & n730 ;
  assign n732 = n731 ^ n728 ;
  assign n733 = n726 & n732 ;
  assign n734 = n733 ^ n726 ;
  assign n735 = n734 ^ n732 ;
  assign n736 = n148 & n735 ;
  assign n703 = x28 & x128 ;
  assign n701 = x27 & x128 ;
  assign n702 = n701 ^ x27 ;
  assign n704 = n703 ^ n702 ;
  assign n705 = x129 & n704 ;
  assign n706 = n705 ^ n704 ;
  assign n707 = n706 ^ n702 ;
  assign n710 = x26 & x128 ;
  assign n708 = x29 & x128 ;
  assign n709 = n708 ^ x29 ;
  assign n711 = n710 ^ n709 ;
  assign n712 = x129 & n711 ;
  assign n713 = n712 ^ n709 ;
  assign n714 = n707 & n713 ;
  assign n715 = n714 ^ n707 ;
  assign n716 = n715 ^ n713 ;
  assign n717 = n137 & n716 ;
  assign n718 = n717 ^ n137 ;
  assign n719 = n718 ^ n137 ;
  assign n737 = n736 ^ n719 ;
  assign n759 = x20 & x128 ;
  assign n757 = x19 & x128 ;
  assign n758 = n757 ^ x19 ;
  assign n760 = n759 ^ n758 ;
  assign n761 = x129 & n760 ;
  assign n762 = n761 ^ n760 ;
  assign n763 = n762 ^ n758 ;
  assign n766 = x18 & x128 ;
  assign n764 = x21 & x128 ;
  assign n765 = n764 ^ x21 ;
  assign n767 = n766 ^ n765 ;
  assign n768 = x129 & n767 ;
  assign n769 = n768 ^ n765 ;
  assign n770 = n763 & n769 ;
  assign n771 = n770 ^ n763 ;
  assign n772 = n771 ^ n769 ;
  assign n773 = n171 & n772 ;
  assign n740 = x24 & x128 ;
  assign n738 = x23 & x128 ;
  assign n739 = n738 ^ x23 ;
  assign n741 = n740 ^ n739 ;
  assign n742 = x129 & n741 ;
  assign n743 = n742 ^ n741 ;
  assign n744 = n743 ^ n739 ;
  assign n747 = x22 & x128 ;
  assign n745 = x25 & x128 ;
  assign n746 = n745 ^ x25 ;
  assign n748 = n747 ^ n746 ;
  assign n749 = x129 & n748 ;
  assign n750 = n749 ^ n746 ;
  assign n751 = n744 & n750 ;
  assign n752 = n751 ^ n744 ;
  assign n753 = n752 ^ n750 ;
  assign n754 = n160 & n753 ;
  assign n755 = n754 ^ n160 ;
  assign n756 = n755 ^ n160 ;
  assign n774 = n773 ^ n756 ;
  assign n775 = n737 & n774 ;
  assign n776 = n775 ^ n737 ;
  assign n777 = n776 ^ n774 ;
  assign n778 = n136 & ~n777 ;
  assign n779 = n778 ^ n136 ;
  assign n844 = n843 ^ n779 ;
  assign n845 = n700 & n844 ;
  assign n846 = n845 ^ n700 ;
  assign n847 = n846 ^ n844 ;
  assign n1167 = n1166 ^ n847 ;
  assign n1168 = x134 & n1167 ;
  assign n1169 = n1168 ^ n1167 ;
  assign n1170 = n1169 ^ n847 ;
  assign n1318 = n406 ^ n383 ;
  assign n1319 = x129 & n1318 ;
  assign n1320 = n1319 ^ n383 ;
  assign n1321 = n148 & n1320 ;
  assign n1313 = n409 ^ n396 ;
  assign n1314 = x129 & n1313 ;
  assign n1315 = n1314 ^ n1313 ;
  assign n1316 = n1315 ^ n396 ;
  assign n1317 = n137 & n1316 ;
  assign n1322 = n1321 ^ n1317 ;
  assign n1328 = n427 ^ n420 ;
  assign n1329 = x129 & n1328 ;
  assign n1330 = n1329 ^ n420 ;
  assign n1331 = n171 & n1330 ;
  assign n1323 = n417 ^ n399 ;
  assign n1324 = x129 & n1323 ;
  assign n1325 = n1324 ^ n1323 ;
  assign n1326 = n1325 ^ n417 ;
  assign n1327 = n160 & n1326 ;
  assign n1332 = n1331 ^ n1327 ;
  assign n1333 = n1322 & n1332 ;
  assign n1334 = n1333 ^ n1322 ;
  assign n1335 = n1334 ^ n1332 ;
  assign n1336 = n188 & n1335 ;
  assign n1293 = n477 ^ n359 ;
  assign n1294 = x129 & n1293 ;
  assign n1295 = n1294 ^ n477 ;
  assign n1296 = n148 & n1295 ;
  assign n1288 = n362 ^ n349 ;
  assign n1289 = x129 & n1288 ;
  assign n1290 = n1289 ^ n1288 ;
  assign n1291 = n1290 ^ n349 ;
  assign n1292 = n137 & n1291 ;
  assign n1297 = n1296 ^ n1292 ;
  assign n1303 = n380 ^ n373 ;
  assign n1304 = x129 & n1303 ;
  assign n1305 = n1304 ^ n373 ;
  assign n1306 = n171 & n1305 ;
  assign n1298 = n370 ^ n352 ;
  assign n1299 = x129 & n1298 ;
  assign n1300 = n1299 ^ n1298 ;
  assign n1301 = n1300 ^ n370 ;
  assign n1302 = n160 & n1301 ;
  assign n1307 = n1306 ^ n1302 ;
  assign n1308 = n1297 & n1307 ;
  assign n1309 = n1308 ^ n1297 ;
  assign n1310 = n1309 ^ n1307 ;
  assign n1311 = n136 & ~n1310 ;
  assign n1312 = n1311 ^ n136 ;
  assign n1337 = n1336 ^ n1312 ;
  assign n1369 = n501 ^ n225 ;
  assign n1370 = x129 & n1369 ;
  assign n1371 = n1370 ^ n225 ;
  assign n1372 = n148 & n1371 ;
  assign n1364 = n504 ^ n490 ;
  assign n1365 = x129 & n1364 ;
  assign n1366 = n1365 ^ n1364 ;
  assign n1367 = n1366 ^ n490 ;
  assign n1368 = n137 & n1367 ;
  assign n1373 = n1372 ^ n1368 ;
  assign n1379 = n522 ^ n515 ;
  assign n1380 = x129 & n1379 ;
  assign n1381 = n1380 ^ n515 ;
  assign n1382 = n171 & n1381 ;
  assign n1374 = n512 ^ n493 ;
  assign n1375 = x129 & n1374 ;
  assign n1376 = n1375 ^ n1374 ;
  assign n1377 = n1376 ^ n512 ;
  assign n1378 = n160 & n1377 ;
  assign n1383 = n1382 ^ n1378 ;
  assign n1384 = n1373 & n1383 ;
  assign n1385 = n1384 ^ n1373 ;
  assign n1386 = n1385 ^ n1383 ;
  assign n1387 = n236 & n1386 ;
  assign n1343 = n525 ^ n453 ;
  assign n1344 = x129 & n1343 ;
  assign n1345 = n1344 ^ n1343 ;
  assign n1346 = n1345 ^ n453 ;
  assign n1347 = n148 & n1346 ;
  assign n1338 = n456 ^ n443 ;
  assign n1339 = x129 & n1338 ;
  assign n1340 = n1339 ^ n1338 ;
  assign n1341 = n1340 ^ n443 ;
  assign n1342 = n137 & n1341 ;
  assign n1348 = n1347 ^ n1342 ;
  assign n1354 = n474 ^ n467 ;
  assign n1355 = x129 & n1354 ;
  assign n1356 = n1355 ^ n467 ;
  assign n1357 = n171 & n1356 ;
  assign n1349 = n464 ^ n446 ;
  assign n1350 = x129 & n1349 ;
  assign n1351 = n1350 ^ n1349 ;
  assign n1352 = n1351 ^ n464 ;
  assign n1353 = n160 & n1352 ;
  assign n1358 = n1357 ^ n1353 ;
  assign n1359 = n1348 & n1358 ;
  assign n1360 = n1359 ^ n1348 ;
  assign n1361 = n1360 ^ n1358 ;
  assign n1362 = n314 & ~n1361 ;
  assign n1363 = n1362 ^ n314 ;
  assign n1388 = n1387 ^ n1363 ;
  assign n1389 = n1337 & n1388 ;
  assign n1390 = n1389 ^ n1337 ;
  assign n1391 = n1390 ^ n1388 ;
  assign n1201 = n430 ^ n249 ;
  assign n1202 = x129 & n1201 ;
  assign n1203 = n1202 ^ n1201 ;
  assign n1204 = n1203 ^ n249 ;
  assign n1205 = n148 & n1204 ;
  assign n1196 = n252 ^ n239 ;
  assign n1197 = x129 & n1196 ;
  assign n1198 = n1197 ^ n1196 ;
  assign n1199 = n1198 ^ n239 ;
  assign n1200 = n137 & n1199 ;
  assign n1206 = n1205 ^ n1200 ;
  assign n1212 = n270 ^ n263 ;
  assign n1213 = x129 & n1212 ;
  assign n1214 = n1213 ^ n263 ;
  assign n1215 = n171 & n1214 ;
  assign n1207 = n260 ^ n242 ;
  assign n1208 = x129 & n1207 ;
  assign n1209 = n1208 ^ n1207 ;
  assign n1210 = n1209 ^ n260 ;
  assign n1211 = n160 & n1210 ;
  assign n1216 = n1215 ^ n1211 ;
  assign n1217 = n1206 & n1216 ;
  assign n1218 = n1217 ^ n1206 ;
  assign n1219 = n1218 ^ n1216 ;
  assign n1220 = n236 & n1219 ;
  assign n1176 = n201 ^ n177 ;
  assign n1177 = x129 & n1176 ;
  assign n1178 = n1177 ^ n177 ;
  assign n1179 = n148 & n1178 ;
  assign n1171 = n204 ^ n191 ;
  assign n1172 = x129 & n1171 ;
  assign n1173 = n1172 ^ n1171 ;
  assign n1174 = n1173 ^ n191 ;
  assign n1175 = n137 & n1174 ;
  assign n1180 = n1179 ^ n1175 ;
  assign n1186 = n222 ^ n215 ;
  assign n1187 = x129 & n1186 ;
  assign n1188 = n1187 ^ n215 ;
  assign n1189 = n171 & n1188 ;
  assign n1181 = n212 ^ n194 ;
  assign n1182 = x129 & n1181 ;
  assign n1183 = n1182 ^ n1181 ;
  assign n1184 = n1183 ^ n212 ;
  assign n1185 = n160 & n1184 ;
  assign n1190 = n1189 ^ n1185 ;
  assign n1191 = n1180 & n1190 ;
  assign n1192 = n1191 ^ n1180 ;
  assign n1193 = n1192 ^ n1190 ;
  assign n1194 = n188 & ~n1193 ;
  assign n1195 = n1194 ^ n188 ;
  assign n1221 = n1220 ^ n1195 ;
  assign n1252 = n327 ^ n273 ;
  assign n1253 = x129 & n1252 ;
  assign n1254 = n1253 ^ n1252 ;
  assign n1255 = n1254 ^ n327 ;
  assign n1256 = n148 & n1255 ;
  assign n1247 = n330 ^ n317 ;
  assign n1248 = x129 & n1247 ;
  assign n1249 = n1248 ^ n1247 ;
  assign n1250 = n1249 ^ n317 ;
  assign n1251 = n137 & n1250 ;
  assign n1257 = n1256 ^ n1251 ;
  assign n1270 = x38 ^ x37 ;
  assign n1271 = x128 & n1270 ;
  assign n1272 = n1271 ^ x38 ;
  assign n1273 = n1272 ^ n305 ;
  assign n1274 = x129 & n1273 ;
  assign n1275 = n1274 ^ x129 ;
  assign n1276 = n1275 ^ x129 ;
  assign n1277 = n1276 ^ n1272 ;
  assign n1278 = n171 & n1277 ;
  assign n1258 = x40 ^ x39 ;
  assign n1259 = x128 & n1258 ;
  assign n1260 = n1259 ^ x40 ;
  assign n1261 = n1260 ^ n320 ;
  assign n1262 = x129 & n1261 ;
  assign n1263 = n1262 ^ x129 ;
  assign n1264 = n1263 ^ x129 ;
  assign n1265 = n1264 ^ n1261 ;
  assign n1266 = n1265 ^ n1260 ;
  assign n1267 = n160 & n1266 ;
  assign n1268 = n1267 ^ n160 ;
  assign n1269 = n1268 ^ n160 ;
  assign n1279 = n1278 ^ n1269 ;
  assign n1280 = n1257 & n1279 ;
  assign n1281 = n1280 ^ n1257 ;
  assign n1282 = n1281 ^ n1279 ;
  assign n1283 = n314 & n1282 ;
  assign n1227 = n308 ^ n151 ;
  assign n1228 = x129 & n1227 ;
  assign n1229 = n1228 ^ n308 ;
  assign n1230 = n148 & n1229 ;
  assign n1222 = n154 ^ n140 ;
  assign n1223 = x129 & n1222 ;
  assign n1224 = n1223 ^ n1222 ;
  assign n1225 = n1224 ^ n140 ;
  assign n1226 = n137 & n1225 ;
  assign n1231 = n1230 ^ n1226 ;
  assign n1237 = n174 ^ n166 ;
  assign n1238 = x129 & n1237 ;
  assign n1239 = n1238 ^ n166 ;
  assign n1240 = n171 & n1239 ;
  assign n1232 = n163 ^ n143 ;
  assign n1233 = x129 & n1232 ;
  assign n1234 = n1233 ^ n1232 ;
  assign n1235 = n1234 ^ n163 ;
  assign n1236 = n160 & n1235 ;
  assign n1241 = n1240 ^ n1236 ;
  assign n1242 = n1231 & n1241 ;
  assign n1243 = n1242 ^ n1231 ;
  assign n1244 = n1243 ^ n1241 ;
  assign n1245 = n136 & ~n1244 ;
  assign n1246 = n1245 ^ n136 ;
  assign n1284 = n1283 ^ n1246 ;
  assign n1285 = n1221 & n1284 ;
  assign n1286 = n1285 ^ n1221 ;
  assign n1287 = n1286 ^ n1284 ;
  assign n1392 = n1391 ^ n1287 ;
  assign n1393 = x134 & n1392 ;
  assign n1394 = n1393 ^ n1392 ;
  assign n1395 = n1394 ^ n1287 ;
  assign n1695 = n1142 ^ n1027 ;
  assign n1696 = x129 & n1695 ;
  assign n1697 = n1696 ^ n1695 ;
  assign n1698 = n1697 ^ n1027 ;
  assign n1699 = n1150 ^ n1033 ;
  assign n1700 = x129 & n1699 ;
  assign n1701 = n1700 ^ n1699 ;
  assign n1702 = n1701 ^ n1033 ;
  assign n1703 = n1698 & n1702 ;
  assign n1704 = n1703 ^ n1698 ;
  assign n1705 = n1704 ^ n1702 ;
  assign n1706 = n148 & n1705 ;
  assign n1681 = n1026 ^ n1008 ;
  assign n1682 = x129 & n1681 ;
  assign n1683 = n1682 ^ n1681 ;
  assign n1684 = n1683 ^ n1008 ;
  assign n1685 = n1034 ^ n1014 ;
  assign n1686 = x129 & n1685 ;
  assign n1687 = n1686 ^ n1685 ;
  assign n1688 = n1687 ^ n1014 ;
  assign n1689 = n1684 & n1688 ;
  assign n1690 = n1689 ^ n1684 ;
  assign n1691 = n1690 ^ n1688 ;
  assign n1692 = n137 & n1691 ;
  assign n1693 = n1692 ^ n137 ;
  assign n1694 = n1693 ^ n137 ;
  assign n1707 = n1706 ^ n1694 ;
  assign n1722 = n1064 ^ n1044 ;
  assign n1723 = x129 & n1722 ;
  assign n1724 = n1723 ^ n1044 ;
  assign n1725 = n1070 ^ n1052 ;
  assign n1726 = x129 & n1725 ;
  assign n1727 = n1726 ^ n1052 ;
  assign n1728 = n1724 & n1727 ;
  assign n1729 = n1728 ^ n1724 ;
  assign n1730 = n1729 ^ n1727 ;
  assign n1731 = n171 & n1730 ;
  assign n1708 = n1045 ^ n1007 ;
  assign n1709 = x129 & n1708 ;
  assign n1710 = n1709 ^ n1708 ;
  assign n1711 = n1710 ^ n1045 ;
  assign n1712 = n1051 ^ n1015 ;
  assign n1713 = x129 & n1712 ;
  assign n1714 = n1713 ^ n1712 ;
  assign n1715 = n1714 ^ n1051 ;
  assign n1716 = n1711 & n1715 ;
  assign n1717 = n1716 ^ n1711 ;
  assign n1718 = n1717 ^ n1715 ;
  assign n1719 = n160 & n1718 ;
  assign n1720 = n1719 ^ n160 ;
  assign n1721 = n1720 ^ n160 ;
  assign n1732 = n1731 ^ n1721 ;
  assign n1733 = n1707 & n1732 ;
  assign n1734 = n1733 ^ n1707 ;
  assign n1735 = n1734 ^ n1732 ;
  assign n1736 = n314 & n1735 ;
  assign n1640 = n1063 ^ n869 ;
  assign n1641 = x129 & n1640 ;
  assign n1642 = n1641 ^ n1063 ;
  assign n1643 = n1071 ^ n875 ;
  assign n1644 = x129 & n1643 ;
  assign n1645 = n1644 ^ n1071 ;
  assign n1646 = n1642 & n1645 ;
  assign n1647 = n1646 ^ n1642 ;
  assign n1648 = n1647 ^ n1645 ;
  assign n1649 = n148 & n1648 ;
  assign n1626 = n868 ^ n850 ;
  assign n1627 = x129 & n1626 ;
  assign n1628 = n1627 ^ n1626 ;
  assign n1629 = n1628 ^ n850 ;
  assign n1630 = n876 ^ n856 ;
  assign n1631 = x129 & n1630 ;
  assign n1632 = n1631 ^ n1630 ;
  assign n1633 = n1632 ^ n856 ;
  assign n1634 = n1629 & n1633 ;
  assign n1635 = n1634 ^ n1629 ;
  assign n1636 = n1635 ^ n1633 ;
  assign n1637 = n137 & n1636 ;
  assign n1638 = n1637 ^ n137 ;
  assign n1639 = n1638 ^ n137 ;
  assign n1650 = n1649 ^ n1639 ;
  assign n1665 = n906 ^ n886 ;
  assign n1666 = x129 & n1665 ;
  assign n1667 = n1666 ^ n886 ;
  assign n1668 = n912 ^ n894 ;
  assign n1669 = x129 & n1668 ;
  assign n1670 = n1669 ^ n894 ;
  assign n1671 = n1667 & n1670 ;
  assign n1672 = n1671 ^ n1667 ;
  assign n1673 = n1672 ^ n1670 ;
  assign n1674 = n171 & n1673 ;
  assign n1651 = n887 ^ n849 ;
  assign n1652 = x129 & n1651 ;
  assign n1653 = n1652 ^ n1651 ;
  assign n1654 = n1653 ^ n887 ;
  assign n1655 = n893 ^ n857 ;
  assign n1656 = x129 & n1655 ;
  assign n1657 = n1656 ^ n1655 ;
  assign n1658 = n1657 ^ n893 ;
  assign n1659 = n1654 & n1658 ;
  assign n1660 = n1659 ^ n1654 ;
  assign n1661 = n1660 ^ n1658 ;
  assign n1662 = n160 & n1661 ;
  assign n1663 = n1662 ^ n160 ;
  assign n1664 = n1663 ^ n160 ;
  assign n1675 = n1674 ^ n1664 ;
  assign n1676 = n1650 & n1675 ;
  assign n1677 = n1676 ^ n1650 ;
  assign n1678 = n1677 ^ n1675 ;
  assign n1679 = n136 & ~n1678 ;
  assign n1680 = n1679 ^ n136 ;
  assign n1737 = n1736 ^ n1680 ;
  assign n1807 = n1106 ^ n600 ;
  assign n1808 = x129 & n1807 ;
  assign n1809 = n1808 ^ n600 ;
  assign n1810 = n1112 ^ n608 ;
  assign n1811 = x129 & n1810 ;
  assign n1812 = n1811 ^ n608 ;
  assign n1813 = n1809 & n1812 ;
  assign n1814 = n1813 ^ n1809 ;
  assign n1815 = n1814 ^ n1812 ;
  assign n1816 = n148 & n1815 ;
  assign n1793 = n1105 ^ n1087 ;
  assign n1794 = x129 & n1793 ;
  assign n1795 = n1794 ^ n1793 ;
  assign n1796 = n1795 ^ n1087 ;
  assign n1797 = n1113 ^ n1093 ;
  assign n1798 = x129 & n1797 ;
  assign n1799 = n1798 ^ n1797 ;
  assign n1800 = n1799 ^ n1093 ;
  assign n1801 = n1796 & n1800 ;
  assign n1802 = n1801 ^ n1796 ;
  assign n1803 = n1802 ^ n1800 ;
  assign n1804 = n137 & n1803 ;
  assign n1805 = n1804 ^ n137 ;
  assign n1806 = n1805 ^ n137 ;
  assign n1817 = n1816 ^ n1806 ;
  assign n1832 = n1143 ^ n1123 ;
  assign n1833 = x129 & n1832 ;
  assign n1834 = n1833 ^ n1123 ;
  assign n1835 = n1149 ^ n1131 ;
  assign n1836 = x129 & n1835 ;
  assign n1837 = n1836 ^ n1131 ;
  assign n1838 = n1834 & n1837 ;
  assign n1839 = n1838 ^ n1834 ;
  assign n1840 = n1839 ^ n1837 ;
  assign n1841 = n171 & n1840 ;
  assign n1818 = n1124 ^ n1086 ;
  assign n1819 = x129 & n1818 ;
  assign n1820 = n1819 ^ n1818 ;
  assign n1821 = n1820 ^ n1124 ;
  assign n1822 = n1130 ^ n1094 ;
  assign n1823 = x129 & n1822 ;
  assign n1824 = n1823 ^ n1822 ;
  assign n1825 = n1824 ^ n1130 ;
  assign n1826 = n1821 & n1825 ;
  assign n1827 = n1826 ^ n1821 ;
  assign n1828 = n1827 ^ n1825 ;
  assign n1829 = n160 & n1828 ;
  assign n1830 = n1829 ^ n160 ;
  assign n1831 = n1830 ^ n160 ;
  assign n1842 = n1841 ^ n1831 ;
  assign n1843 = n1817 & n1842 ;
  assign n1844 = n1843 ^ n1817 ;
  assign n1845 = n1844 ^ n1842 ;
  assign n1846 = n236 & n1845 ;
  assign n1752 = n948 ^ n905 ;
  assign n1753 = x129 & n1752 ;
  assign n1754 = n1753 ^ n905 ;
  assign n1755 = n954 ^ n913 ;
  assign n1756 = x129 & n1755 ;
  assign n1757 = n1756 ^ n913 ;
  assign n1758 = n1754 & n1757 ;
  assign n1759 = n1758 ^ n1754 ;
  assign n1760 = n1759 ^ n1757 ;
  assign n1761 = n148 & n1760 ;
  assign n1738 = n947 ^ n929 ;
  assign n1739 = x129 & n1738 ;
  assign n1740 = n1739 ^ n1738 ;
  assign n1741 = n1740 ^ n929 ;
  assign n1742 = n955 ^ n935 ;
  assign n1743 = x129 & n1742 ;
  assign n1744 = n1743 ^ n1742 ;
  assign n1745 = n1744 ^ n935 ;
  assign n1746 = n1741 & n1745 ;
  assign n1747 = n1746 ^ n1741 ;
  assign n1748 = n1747 ^ n1745 ;
  assign n1749 = n137 & n1748 ;
  assign n1750 = n1749 ^ n137 ;
  assign n1751 = n1750 ^ n137 ;
  assign n1762 = n1761 ^ n1751 ;
  assign n1777 = n985 ^ n965 ;
  assign n1778 = x129 & n1777 ;
  assign n1779 = n1778 ^ n965 ;
  assign n1780 = n991 ^ n973 ;
  assign n1781 = x129 & n1780 ;
  assign n1782 = n1781 ^ n973 ;
  assign n1783 = n1779 & n1782 ;
  assign n1784 = n1783 ^ n1779 ;
  assign n1785 = n1784 ^ n1782 ;
  assign n1786 = n171 & n1785 ;
  assign n1763 = n966 ^ n928 ;
  assign n1764 = x129 & n1763 ;
  assign n1765 = n1764 ^ n1763 ;
  assign n1766 = n1765 ^ n966 ;
  assign n1767 = n972 ^ n936 ;
  assign n1768 = x129 & n1767 ;
  assign n1769 = n1768 ^ n1767 ;
  assign n1770 = n1769 ^ n972 ;
  assign n1771 = n1766 & n1770 ;
  assign n1772 = n1771 ^ n1766 ;
  assign n1773 = n1772 ^ n1770 ;
  assign n1774 = n160 & n1773 ;
  assign n1775 = n1774 ^ n160 ;
  assign n1776 = n1775 ^ n160 ;
  assign n1787 = n1786 ^ n1776 ;
  assign n1788 = n1762 & n1787 ;
  assign n1789 = n1788 ^ n1762 ;
  assign n1790 = n1789 ^ n1787 ;
  assign n1791 = n188 & ~n1790 ;
  assign n1792 = n1791 ^ n188 ;
  assign n1847 = n1846 ^ n1792 ;
  assign n1848 = n1737 & n1847 ;
  assign n1849 = n1848 ^ n1737 ;
  assign n1850 = n1849 ^ n1847 ;
  assign n1468 = n984 ^ n643 ;
  assign n1469 = x129 & n1468 ;
  assign n1470 = n1469 ^ n1468 ;
  assign n1471 = n1470 ^ n643 ;
  assign n1472 = n992 ^ n649 ;
  assign n1473 = x129 & n1472 ;
  assign n1474 = n1473 ^ n1472 ;
  assign n1475 = n1474 ^ n649 ;
  assign n1476 = n1471 & n1475 ;
  assign n1477 = n1476 ^ n1471 ;
  assign n1478 = n1477 ^ n1475 ;
  assign n1479 = n148 & n1478 ;
  assign n1454 = n642 ^ n624 ;
  assign n1455 = x129 & n1454 ;
  assign n1456 = n1455 ^ n1454 ;
  assign n1457 = n1456 ^ n624 ;
  assign n1458 = n650 ^ n630 ;
  assign n1459 = x129 & n1458 ;
  assign n1460 = n1459 ^ n1458 ;
  assign n1461 = n1460 ^ n630 ;
  assign n1462 = n1457 & n1461 ;
  assign n1463 = n1462 ^ n1457 ;
  assign n1464 = n1463 ^ n1461 ;
  assign n1465 = n137 & n1464 ;
  assign n1466 = n1465 ^ n137 ;
  assign n1467 = n1466 ^ n137 ;
  assign n1480 = n1479 ^ n1467 ;
  assign n1495 = n680 ^ n660 ;
  assign n1496 = x129 & n1495 ;
  assign n1497 = n1496 ^ n660 ;
  assign n1498 = n686 ^ n668 ;
  assign n1499 = x129 & n1498 ;
  assign n1500 = n1499 ^ n668 ;
  assign n1501 = n1497 & n1500 ;
  assign n1502 = n1501 ^ n1497 ;
  assign n1503 = n1502 ^ n1500 ;
  assign n1504 = n171 & n1503 ;
  assign n1481 = n661 ^ n623 ;
  assign n1482 = x129 & n1481 ;
  assign n1483 = n1482 ^ n1481 ;
  assign n1484 = n1483 ^ n661 ;
  assign n1485 = n667 ^ n631 ;
  assign n1486 = x129 & n1485 ;
  assign n1487 = n1486 ^ n1485 ;
  assign n1488 = n1487 ^ n667 ;
  assign n1489 = n1484 & n1488 ;
  assign n1490 = n1489 ^ n1484 ;
  assign n1491 = n1490 ^ n1488 ;
  assign n1492 = n160 & n1491 ;
  assign n1493 = n1492 ^ n160 ;
  assign n1494 = n1493 ^ n160 ;
  assign n1505 = n1504 ^ n1494 ;
  assign n1506 = n1480 & n1505 ;
  assign n1507 = n1506 ^ n1480 ;
  assign n1508 = n1507 ^ n1505 ;
  assign n1509 = n236 & n1508 ;
  assign n1405 = n795 ^ n679 ;
  assign n1406 = x129 & n1405 ;
  assign n1407 = n1406 ^ n1405 ;
  assign n1408 = n1407 ^ n795 ;
  assign n1409 = n801 ^ n687 ;
  assign n1410 = x129 & n1409 ;
  assign n1411 = n1410 ^ n1409 ;
  assign n1412 = n1411 ^ n801 ;
  assign n1413 = n1408 & n1412 ;
  assign n1414 = n1413 ^ n1408 ;
  assign n1415 = n1414 ^ n1412 ;
  assign n1416 = n148 & n1415 ;
  assign n1396 = x47 ^ x46 ;
  assign n1397 = x128 & n1396 ;
  assign n1398 = n1397 ^ x47 ;
  assign n1399 = n1398 ^ n782 ;
  assign n1400 = x129 & ~n1399 ;
  assign n1401 = n1400 ^ x129 ;
  assign n1402 = n1401 ^ n1398 ;
  assign n1403 = n137 & ~n1402 ;
  assign n1404 = n1403 ^ n137 ;
  assign n1417 = n1416 ^ n1404 ;
  assign n1437 = n286 ^ x39 ;
  assign n1438 = n1437 ^ n825 ;
  assign n1439 = x129 & n1438 ;
  assign n1440 = n1439 ^ n1437 ;
  assign n1441 = n830 ^ n284 ;
  assign n1442 = x129 & n1441 ;
  assign n1443 = n1442 ^ n284 ;
  assign n1444 = n1440 & n1443 ;
  assign n1445 = n1444 ^ n1440 ;
  assign n1446 = n1445 ^ n1443 ;
  assign n1447 = n171 & n1446 ;
  assign n1418 = x43 & x128 ;
  assign n1419 = n1418 ^ x43 ;
  assign n1420 = n1419 ^ n291 ;
  assign n1421 = x129 & n1420 ;
  assign n1422 = n1421 ^ n1420 ;
  assign n1423 = n1422 ^ n291 ;
  assign n1426 = x42 & x128 ;
  assign n1424 = x41 & x128 ;
  assign n1425 = n1424 ^ x41 ;
  assign n1427 = n1426 ^ n1425 ;
  assign n1428 = x129 & n1427 ;
  assign n1429 = n1428 ^ n1427 ;
  assign n1430 = n1429 ^ n1425 ;
  assign n1431 = n1423 & n1430 ;
  assign n1432 = n1431 ^ n1423 ;
  assign n1433 = n1432 ^ n1430 ;
  assign n1434 = n160 & n1433 ;
  assign n1435 = n1434 ^ n160 ;
  assign n1436 = n1435 ^ n160 ;
  assign n1448 = n1447 ^ n1436 ;
  assign n1449 = n1417 & n1448 ;
  assign n1450 = n1449 ^ n1417 ;
  assign n1451 = n1450 ^ n1448 ;
  assign n1452 = n314 & ~n1451 ;
  assign n1453 = n1452 ^ n314 ;
  assign n1510 = n1509 ^ n1453 ;
  assign n1582 = n758 ^ n564 ;
  assign n1583 = x129 & n1582 ;
  assign n1584 = n1583 ^ n758 ;
  assign n1585 = n766 ^ n570 ;
  assign n1586 = x129 & n1585 ;
  assign n1587 = n1586 ^ n766 ;
  assign n1588 = n1584 & n1587 ;
  assign n1589 = n1588 ^ n1584 ;
  assign n1590 = n1589 ^ n1587 ;
  assign n1591 = n148 & n1590 ;
  assign n1568 = n563 ^ n545 ;
  assign n1569 = x129 & n1568 ;
  assign n1570 = n1569 ^ n1568 ;
  assign n1571 = n1570 ^ n545 ;
  assign n1572 = n571 ^ n551 ;
  assign n1573 = x129 & n1572 ;
  assign n1574 = n1573 ^ n1572 ;
  assign n1575 = n1574 ^ n551 ;
  assign n1576 = n1571 & n1575 ;
  assign n1577 = n1576 ^ n1571 ;
  assign n1578 = n1577 ^ n1575 ;
  assign n1579 = n137 & n1578 ;
  assign n1580 = n1579 ^ n137 ;
  assign n1581 = n1580 ^ n137 ;
  assign n1592 = n1591 ^ n1581 ;
  assign n1607 = n601 ^ n581 ;
  assign n1608 = x129 & n1607 ;
  assign n1609 = n1608 ^ n581 ;
  assign n1610 = n607 ^ n589 ;
  assign n1611 = x129 & n1610 ;
  assign n1612 = n1611 ^ n589 ;
  assign n1613 = n1609 & n1612 ;
  assign n1614 = n1613 ^ n1609 ;
  assign n1615 = n1614 ^ n1612 ;
  assign n1616 = n171 & n1615 ;
  assign n1593 = n582 ^ n544 ;
  assign n1594 = x129 & n1593 ;
  assign n1595 = n1594 ^ n1593 ;
  assign n1596 = n1595 ^ n582 ;
  assign n1597 = n588 ^ n552 ;
  assign n1598 = x129 & n1597 ;
  assign n1599 = n1598 ^ n1597 ;
  assign n1600 = n1599 ^ n588 ;
  assign n1601 = n1596 & n1600 ;
  assign n1602 = n1601 ^ n1596 ;
  assign n1603 = n1602 ^ n1600 ;
  assign n1604 = n160 & n1603 ;
  assign n1605 = n1604 ^ n160 ;
  assign n1606 = n1605 ^ n160 ;
  assign n1617 = n1616 ^ n1606 ;
  assign n1618 = n1592 & n1617 ;
  assign n1619 = n1618 ^ n1592 ;
  assign n1620 = n1619 ^ n1617 ;
  assign n1621 = n188 & n1620 ;
  assign n1525 = n824 ^ n722 ;
  assign n1526 = x129 & n1525 ;
  assign n1527 = n1526 ^ n1525 ;
  assign n1528 = n1527 ^ n722 ;
  assign n1529 = n831 ^ n728 ;
  assign n1530 = x129 & n1529 ;
  assign n1531 = n1530 ^ n1529 ;
  assign n1532 = n1531 ^ n728 ;
  assign n1533 = n1528 & n1532 ;
  assign n1534 = n1533 ^ n1528 ;
  assign n1535 = n1534 ^ n1532 ;
  assign n1536 = n148 & n1535 ;
  assign n1511 = n721 ^ n703 ;
  assign n1512 = x129 & n1511 ;
  assign n1513 = n1512 ^ n1511 ;
  assign n1514 = n1513 ^ n703 ;
  assign n1515 = n729 ^ n709 ;
  assign n1516 = x129 & n1515 ;
  assign n1517 = n1516 ^ n1515 ;
  assign n1518 = n1517 ^ n709 ;
  assign n1519 = n1514 & n1518 ;
  assign n1520 = n1519 ^ n1514 ;
  assign n1521 = n1520 ^ n1518 ;
  assign n1522 = n137 & n1521 ;
  assign n1523 = n1522 ^ n137 ;
  assign n1524 = n1523 ^ n137 ;
  assign n1537 = n1536 ^ n1524 ;
  assign n1552 = n759 ^ n739 ;
  assign n1553 = x129 & n1552 ;
  assign n1554 = n1553 ^ n739 ;
  assign n1555 = n765 ^ n747 ;
  assign n1556 = x129 & n1555 ;
  assign n1557 = n1556 ^ n747 ;
  assign n1558 = n1554 & n1557 ;
  assign n1559 = n1558 ^ n1554 ;
  assign n1560 = n1559 ^ n1557 ;
  assign n1561 = n171 & n1560 ;
  assign n1538 = n740 ^ n702 ;
  assign n1539 = x129 & n1538 ;
  assign n1540 = n1539 ^ n1538 ;
  assign n1541 = n1540 ^ n740 ;
  assign n1542 = n746 ^ n710 ;
  assign n1543 = x129 & n1542 ;
  assign n1544 = n1543 ^ n1542 ;
  assign n1545 = n1544 ^ n746 ;
  assign n1546 = n1541 & n1545 ;
  assign n1547 = n1546 ^ n1541 ;
  assign n1548 = n1547 ^ n1545 ;
  assign n1549 = n160 & n1548 ;
  assign n1550 = n1549 ^ n160 ;
  assign n1551 = n1550 ^ n160 ;
  assign n1562 = n1561 ^ n1551 ;
  assign n1563 = n1537 & n1562 ;
  assign n1564 = n1563 ^ n1537 ;
  assign n1565 = n1564 ^ n1562 ;
  assign n1566 = n136 & ~n1565 ;
  assign n1567 = n1566 ^ n136 ;
  assign n1622 = n1621 ^ n1567 ;
  assign n1623 = n1510 & n1622 ;
  assign n1624 = n1623 ^ n1510 ;
  assign n1625 = n1624 ^ n1622 ;
  assign n1851 = n1850 ^ n1625 ;
  assign n1852 = x134 & n1851 ;
  assign n1853 = n1852 ^ n1851 ;
  assign n1854 = n1853 ^ n1625 ;
  assign n1917 = n148 & n386 ;
  assign n1916 = n137 & n412 ;
  assign n1918 = n1917 ^ n1916 ;
  assign n1920 = n171 & n423 ;
  assign n1919 = n160 & n402 ;
  assign n1921 = n1920 ^ n1919 ;
  assign n1922 = n1918 & n1921 ;
  assign n1923 = n1922 ^ n1918 ;
  assign n1924 = n1923 ^ n1921 ;
  assign n1925 = n188 & n1924 ;
  assign n1906 = n148 & n480 ;
  assign n1905 = n137 & n365 ;
  assign n1907 = n1906 ^ n1905 ;
  assign n1909 = n171 & n376 ;
  assign n1908 = n160 & n355 ;
  assign n1910 = n1909 ^ n1908 ;
  assign n1911 = n1907 & n1910 ;
  assign n1912 = n1911 ^ n1907 ;
  assign n1913 = n1912 ^ n1910 ;
  assign n1914 = n136 & ~n1913 ;
  assign n1915 = n1914 ^ n136 ;
  assign n1926 = n1925 ^ n1915 ;
  assign n1939 = n148 & n228 ;
  assign n1938 = n137 & n507 ;
  assign n1940 = n1939 ^ n1938 ;
  assign n1942 = n171 & n518 ;
  assign n1941 = n160 & n496 ;
  assign n1943 = n1942 ^ n1941 ;
  assign n1944 = n1940 & n1943 ;
  assign n1945 = n1944 ^ n1940 ;
  assign n1946 = n1945 ^ n1943 ;
  assign n1947 = n236 & n1946 ;
  assign n1928 = n148 & n528 ;
  assign n1927 = n137 & n459 ;
  assign n1929 = n1928 ^ n1927 ;
  assign n1931 = n171 & n470 ;
  assign n1930 = n160 & n449 ;
  assign n1932 = n1931 ^ n1930 ;
  assign n1933 = n1929 & n1932 ;
  assign n1934 = n1933 ^ n1929 ;
  assign n1935 = n1934 ^ n1932 ;
  assign n1936 = n314 & ~n1935 ;
  assign n1937 = n1936 ^ n314 ;
  assign n1948 = n1947 ^ n1937 ;
  assign n1949 = n1926 & n1948 ;
  assign n1950 = n1949 ^ n1926 ;
  assign n1951 = n1950 ^ n1948 ;
  assign n1856 = n171 & n299 ;
  assign n1855 = n160 & n323 ;
  assign n1857 = n1856 ^ n1855 ;
  assign n1859 = n148 & n276 ;
  assign n1858 = n137 & n333 ;
  assign n1860 = n1859 ^ n1858 ;
  assign n1861 = n314 & n1860 ;
  assign n1862 = n1861 ^ n314 ;
  assign n1863 = n1857 & n1862 ;
  assign n1864 = n1863 ^ n1862 ;
  assign n1865 = n1864 ^ n314 ;
  assign n1867 = n148 & n433 ;
  assign n1866 = n137 & n255 ;
  assign n1868 = n1867 ^ n1866 ;
  assign n1870 = n171 & n266 ;
  assign n1869 = n160 & n245 ;
  assign n1871 = n1870 ^ n1869 ;
  assign n1872 = n1868 & n1871 ;
  assign n1873 = n1872 ^ n1868 ;
  assign n1874 = n1873 ^ n1871 ;
  assign n1875 = n236 & ~n1874 ;
  assign n1876 = n1875 ^ n236 ;
  assign n1877 = n1865 & n1876 ;
  assign n1878 = n1877 ^ n1865 ;
  assign n1879 = n1878 ^ n1876 ;
  assign n1892 = n148 & n311 ;
  assign n1891 = n137 & n157 ;
  assign n1893 = n1892 ^ n1891 ;
  assign n1895 = n169 & n171 ;
  assign n1894 = n146 & n160 ;
  assign n1896 = n1895 ^ n1894 ;
  assign n1897 = n1893 & n1896 ;
  assign n1898 = n1897 ^ n1893 ;
  assign n1899 = n1898 ^ n1896 ;
  assign n1900 = n136 & n1899 ;
  assign n1881 = n148 & n180 ;
  assign n1880 = n137 & n207 ;
  assign n1882 = n1881 ^ n1880 ;
  assign n1884 = n171 & n218 ;
  assign n1883 = n160 & n197 ;
  assign n1885 = n1884 ^ n1883 ;
  assign n1886 = n1882 & n1885 ;
  assign n1887 = n1886 ^ n1882 ;
  assign n1888 = n1887 ^ n1885 ;
  assign n1889 = n188 & ~n1888 ;
  assign n1890 = n1889 ^ n188 ;
  assign n1901 = n1900 ^ n1890 ;
  assign n1902 = n1879 & n1901 ;
  assign n1903 = n1902 ^ n1879 ;
  assign n1904 = n1903 ^ n1901 ;
  assign n1952 = n1951 ^ n1904 ;
  assign n1953 = x134 & n1952 ;
  assign n1954 = n1953 ^ n1952 ;
  assign n1955 = n1954 ^ n1904 ;
  assign n2045 = n148 & n919 ;
  assign n2042 = n137 & n961 ;
  assign n2043 = n2042 ^ n137 ;
  assign n2044 = n2043 ^ n137 ;
  assign n2046 = n2045 ^ n2044 ;
  assign n2050 = n171 & n979 ;
  assign n2047 = n160 & n942 ;
  assign n2048 = n2047 ^ n160 ;
  assign n2049 = n2048 ^ n160 ;
  assign n2051 = n2050 ^ n2049 ;
  assign n2052 = n2046 & n2051 ;
  assign n2053 = n2052 ^ n2046 ;
  assign n2054 = n2053 ^ n2051 ;
  assign n2055 = n188 & n2054 ;
  assign n2030 = n148 & n1077 ;
  assign n2027 = n137 & n882 ;
  assign n2028 = n2027 ^ n137 ;
  assign n2029 = n2028 ^ n137 ;
  assign n2031 = n2030 ^ n2029 ;
  assign n2035 = n171 & n900 ;
  assign n2032 = n160 & n863 ;
  assign n2033 = n2032 ^ n160 ;
  assign n2034 = n2033 ^ n160 ;
  assign n2036 = n2035 ^ n2034 ;
  assign n2037 = n2031 & n2036 ;
  assign n2038 = n2037 ^ n2031 ;
  assign n2039 = n2038 ^ n2036 ;
  assign n2040 = n136 & ~n2039 ;
  assign n2041 = n2040 ^ n136 ;
  assign n2056 = n2055 ^ n2041 ;
  assign n2075 = n148 & n614 ;
  assign n2072 = n137 & n1119 ;
  assign n2073 = n2072 ^ n137 ;
  assign n2074 = n2073 ^ n137 ;
  assign n2076 = n2075 ^ n2074 ;
  assign n2080 = n171 & n1137 ;
  assign n2077 = n160 & n1100 ;
  assign n2078 = n2077 ^ n160 ;
  assign n2079 = n2078 ^ n160 ;
  assign n2081 = n2080 ^ n2079 ;
  assign n2082 = n2076 & n2081 ;
  assign n2083 = n2082 ^ n2076 ;
  assign n2084 = n2083 ^ n2081 ;
  assign n2085 = n236 & n2084 ;
  assign n2060 = n148 & n1156 ;
  assign n2057 = n137 & n1040 ;
  assign n2058 = n2057 ^ n137 ;
  assign n2059 = n2058 ^ n137 ;
  assign n2061 = n2060 ^ n2059 ;
  assign n2065 = n171 & n1058 ;
  assign n2062 = n160 & n1021 ;
  assign n2063 = n2062 ^ n160 ;
  assign n2064 = n2063 ^ n160 ;
  assign n2066 = n2065 ^ n2064 ;
  assign n2067 = n2061 & n2066 ;
  assign n2068 = n2067 ^ n2061 ;
  assign n2069 = n2068 ^ n2066 ;
  assign n2070 = n314 & ~n2069 ;
  assign n2071 = n2070 ^ n314 ;
  assign n2086 = n2085 ^ n2071 ;
  assign n2087 = n2056 & n2086 ;
  assign n2088 = n2087 ^ n2056 ;
  assign n2089 = n2088 ^ n2086 ;
  assign n1964 = n148 & n693 ;
  assign n1961 = n137 & n808 ;
  assign n1962 = n1961 ^ n137 ;
  assign n1963 = n1962 ^ n137 ;
  assign n1965 = n1964 ^ n1963 ;
  assign n1959 = n171 & n820 ;
  assign n1956 = n160 & n790 ;
  assign n1957 = n1956 ^ n160 ;
  assign n1958 = n1957 ^ n160 ;
  assign n1960 = n1959 ^ n1958 ;
  assign n1966 = n1965 ^ n1960 ;
  assign n1967 = n1960 ^ n314 ;
  assign n1968 = n314 & n1967 ;
  assign n1969 = n1968 ^ n1967 ;
  assign n1970 = n1969 ^ n314 ;
  assign n1971 = n1970 ^ n1965 ;
  assign n1972 = n1966 & n1971 ;
  assign n1973 = n1972 ^ n1969 ;
  assign n1974 = n1973 ^ n1965 ;
  assign n1978 = n148 & n998 ;
  assign n1975 = n137 & n656 ;
  assign n1976 = n1975 ^ n137 ;
  assign n1977 = n1976 ^ n137 ;
  assign n1979 = n1978 ^ n1977 ;
  assign n1983 = n171 & n674 ;
  assign n1980 = n160 & n637 ;
  assign n1981 = n1980 ^ n160 ;
  assign n1982 = n1981 ^ n160 ;
  assign n1984 = n1983 ^ n1982 ;
  assign n1985 = n1979 & n1984 ;
  assign n1986 = n1985 ^ n1979 ;
  assign n1987 = n1986 ^ n1984 ;
  assign n1988 = n236 & n1987 ;
  assign n1989 = n1988 ^ n236 ;
  assign n1990 = n1989 ^ n236 ;
  assign n1991 = n1974 & n1990 ;
  assign n1992 = n1991 ^ n1974 ;
  assign n1993 = n1992 ^ n1990 ;
  assign n2012 = n148 & n837 ;
  assign n2009 = n137 & n735 ;
  assign n2010 = n2009 ^ n137 ;
  assign n2011 = n2010 ^ n137 ;
  assign n2013 = n2012 ^ n2011 ;
  assign n2017 = n171 & n753 ;
  assign n2014 = n160 & n716 ;
  assign n2015 = n2014 ^ n160 ;
  assign n2016 = n2015 ^ n160 ;
  assign n2018 = n2017 ^ n2016 ;
  assign n2019 = n2013 & n2018 ;
  assign n2020 = n2019 ^ n2013 ;
  assign n2021 = n2020 ^ n2018 ;
  assign n2022 = n136 & n2021 ;
  assign n1997 = n148 & n772 ;
  assign n1994 = n137 & n577 ;
  assign n1995 = n1994 ^ n137 ;
  assign n1996 = n1995 ^ n137 ;
  assign n1998 = n1997 ^ n1996 ;
  assign n2002 = n171 & n595 ;
  assign n1999 = n160 & n558 ;
  assign n2000 = n1999 ^ n160 ;
  assign n2001 = n2000 ^ n160 ;
  assign n2003 = n2002 ^ n2001 ;
  assign n2004 = n1998 & n2003 ;
  assign n2005 = n2004 ^ n1998 ;
  assign n2006 = n2005 ^ n2003 ;
  assign n2007 = n188 & ~n2006 ;
  assign n2008 = n2007 ^ n188 ;
  assign n2023 = n2022 ^ n2008 ;
  assign n2024 = n1993 & n2023 ;
  assign n2025 = n2024 ^ n1993 ;
  assign n2026 = n2025 ^ n2023 ;
  assign n2090 = n2089 ^ n2026 ;
  assign n2091 = x134 & n2090 ;
  assign n2092 = n2091 ^ n2090 ;
  assign n2093 = n2092 ^ n2026 ;
  assign n2153 = n148 & n1305 ;
  assign n2152 = n137 & n1320 ;
  assign n2154 = n2153 ^ n2152 ;
  assign n2156 = n171 & n1326 ;
  assign n2155 = n160 & n1316 ;
  assign n2157 = n2156 ^ n2155 ;
  assign n2158 = n2154 & n2157 ;
  assign n2159 = n2158 ^ n2154 ;
  assign n2160 = n2159 ^ n2157 ;
  assign n2161 = n188 & n2160 ;
  assign n2142 = n148 & n1356 ;
  assign n2141 = n137 & n1295 ;
  assign n2143 = n2142 ^ n2141 ;
  assign n2145 = n171 & n1301 ;
  assign n2144 = n160 & n1291 ;
  assign n2146 = n2145 ^ n2144 ;
  assign n2147 = n2143 & n2146 ;
  assign n2148 = n2147 ^ n2143 ;
  assign n2149 = n2148 ^ n2146 ;
  assign n2150 = n136 & ~n2149 ;
  assign n2151 = n2150 ^ n136 ;
  assign n2162 = n2161 ^ n2151 ;
  assign n2175 = n148 & n1188 ;
  assign n2174 = n137 & n1371 ;
  assign n2176 = n2175 ^ n2174 ;
  assign n2178 = n171 & n1377 ;
  assign n2177 = n160 & n1367 ;
  assign n2179 = n2178 ^ n2177 ;
  assign n2180 = n2176 & n2179 ;
  assign n2181 = n2180 ^ n2176 ;
  assign n2182 = n2181 ^ n2179 ;
  assign n2183 = n236 & n2182 ;
  assign n2164 = n148 & n1381 ;
  assign n2163 = n137 & n1346 ;
  assign n2165 = n2164 ^ n2163 ;
  assign n2167 = n171 & n1352 ;
  assign n2166 = n160 & n1341 ;
  assign n2168 = n2167 ^ n2166 ;
  assign n2169 = n2165 & n2168 ;
  assign n2170 = n2169 ^ n2165 ;
  assign n2171 = n2170 ^ n2168 ;
  assign n2172 = n314 & ~n2171 ;
  assign n2173 = n2172 ^ n314 ;
  assign n2184 = n2183 ^ n2173 ;
  assign n2185 = n2162 & n2184 ;
  assign n2186 = n2185 ^ n2162 ;
  assign n2187 = n2186 ^ n2184 ;
  assign n2106 = n148 & n1214 ;
  assign n2105 = n137 & n1255 ;
  assign n2107 = n2106 ^ n2105 ;
  assign n2109 = n171 & n1266 ;
  assign n2108 = n160 & n1250 ;
  assign n2110 = n2109 ^ n2108 ;
  assign n2111 = n2107 & n2110 ;
  assign n2112 = n2111 ^ n2107 ;
  assign n2113 = n2112 ^ n2110 ;
  assign n2114 = n314 & n2113 ;
  assign n2095 = n148 & n1330 ;
  assign n2094 = n137 & n1204 ;
  assign n2096 = n2095 ^ n2094 ;
  assign n2098 = n171 & n1210 ;
  assign n2097 = n160 & n1199 ;
  assign n2099 = n2098 ^ n2097 ;
  assign n2100 = n2096 & n2099 ;
  assign n2101 = n2100 ^ n2096 ;
  assign n2102 = n2101 ^ n2099 ;
  assign n2103 = n236 & ~n2102 ;
  assign n2104 = n2103 ^ n236 ;
  assign n2115 = n2114 ^ n2104 ;
  assign n2128 = n148 & n1277 ;
  assign n2127 = n137 & n1229 ;
  assign n2129 = n2128 ^ n2127 ;
  assign n2131 = n171 & n1235 ;
  assign n2130 = n160 & n1225 ;
  assign n2132 = n2131 ^ n2130 ;
  assign n2133 = n2129 & n2132 ;
  assign n2134 = n2133 ^ n2129 ;
  assign n2135 = n2134 ^ n2132 ;
  assign n2136 = n136 & n2135 ;
  assign n2117 = n148 & n1239 ;
  assign n2116 = n137 & n1178 ;
  assign n2118 = n2117 ^ n2116 ;
  assign n2120 = n171 & n1184 ;
  assign n2119 = n160 & n1174 ;
  assign n2121 = n2120 ^ n2119 ;
  assign n2122 = n2118 & n2121 ;
  assign n2123 = n2122 ^ n2118 ;
  assign n2124 = n2123 ^ n2121 ;
  assign n2125 = n188 & ~n2124 ;
  assign n2126 = n2125 ^ n188 ;
  assign n2137 = n2136 ^ n2126 ;
  assign n2138 = n2115 & n2137 ;
  assign n2139 = n2138 ^ n2115 ;
  assign n2140 = n2139 ^ n2137 ;
  assign n2188 = n2187 ^ n2140 ;
  assign n2189 = x134 & n2188 ;
  assign n2190 = n2189 ^ n2188 ;
  assign n2191 = n2190 ^ n2140 ;
  assign n2272 = n148 & n1673 ;
  assign n2269 = n137 & n1760 ;
  assign n2270 = n2269 ^ n137 ;
  assign n2271 = n2270 ^ n137 ;
  assign n2273 = n2272 ^ n2271 ;
  assign n2277 = n171 & n1773 ;
  assign n2274 = n160 & n1748 ;
  assign n2275 = n2274 ^ n160 ;
  assign n2276 = n2275 ^ n160 ;
  assign n2278 = n2277 ^ n2276 ;
  assign n2279 = n2273 & n2278 ;
  assign n2280 = n2279 ^ n2273 ;
  assign n2281 = n2280 ^ n2278 ;
  assign n2282 = n188 & n2281 ;
  assign n2257 = n148 & n1730 ;
  assign n2254 = n137 & n1648 ;
  assign n2255 = n2254 ^ n137 ;
  assign n2256 = n2255 ^ n137 ;
  assign n2258 = n2257 ^ n2256 ;
  assign n2262 = n171 & n1661 ;
  assign n2259 = n160 & n1636 ;
  assign n2260 = n2259 ^ n160 ;
  assign n2261 = n2260 ^ n160 ;
  assign n2263 = n2262 ^ n2261 ;
  assign n2264 = n2258 & n2263 ;
  assign n2265 = n2264 ^ n2258 ;
  assign n2266 = n2265 ^ n2263 ;
  assign n2267 = n136 & ~n2266 ;
  assign n2268 = n2267 ^ n136 ;
  assign n2283 = n2282 ^ n2268 ;
  assign n2302 = n148 & n1615 ;
  assign n2299 = n137 & n1815 ;
  assign n2300 = n2299 ^ n137 ;
  assign n2301 = n2300 ^ n137 ;
  assign n2303 = n2302 ^ n2301 ;
  assign n2307 = n171 & n1828 ;
  assign n2304 = n160 & n1803 ;
  assign n2305 = n2304 ^ n160 ;
  assign n2306 = n2305 ^ n160 ;
  assign n2308 = n2307 ^ n2306 ;
  assign n2309 = n2303 & n2308 ;
  assign n2310 = n2309 ^ n2303 ;
  assign n2311 = n2310 ^ n2308 ;
  assign n2312 = n236 & n2311 ;
  assign n2287 = n148 & n1840 ;
  assign n2284 = n137 & n1705 ;
  assign n2285 = n2284 ^ n137 ;
  assign n2286 = n2285 ^ n137 ;
  assign n2288 = n2287 ^ n2286 ;
  assign n2292 = n171 & n1718 ;
  assign n2289 = n160 & n1691 ;
  assign n2290 = n2289 ^ n160 ;
  assign n2291 = n2290 ^ n160 ;
  assign n2293 = n2292 ^ n2291 ;
  assign n2294 = n2288 & n2293 ;
  assign n2295 = n2294 ^ n2288 ;
  assign n2296 = n2295 ^ n2293 ;
  assign n2297 = n314 & ~n2296 ;
  assign n2298 = n2297 ^ n314 ;
  assign n2313 = n2312 ^ n2298 ;
  assign n2314 = n2283 & n2313 ;
  assign n2315 = n2314 ^ n2283 ;
  assign n2316 = n2315 ^ n2313 ;
  assign n2209 = n137 & n1415 ;
  assign n2207 = n160 & ~n1402 ;
  assign n2208 = n2207 ^ n160 ;
  assign n2210 = n2209 ^ n2208 ;
  assign n2214 = n171 & n1433 ;
  assign n2211 = n148 & n1503 ;
  assign n2212 = n2211 ^ n148 ;
  assign n2213 = n2212 ^ n148 ;
  assign n2215 = n2214 ^ n2213 ;
  assign n2216 = n2210 & n2215 ;
  assign n2217 = n2216 ^ n2210 ;
  assign n2218 = n2217 ^ n2215 ;
  assign n2219 = n314 & n2218 ;
  assign n2195 = n148 & n1785 ;
  assign n2192 = n137 & n1478 ;
  assign n2193 = n2192 ^ n137 ;
  assign n2194 = n2193 ^ n137 ;
  assign n2196 = n2195 ^ n2194 ;
  assign n2200 = n171 & n1491 ;
  assign n2197 = n160 & n1464 ;
  assign n2198 = n2197 ^ n160 ;
  assign n2199 = n2198 ^ n160 ;
  assign n2201 = n2200 ^ n2199 ;
  assign n2202 = n2196 & n2201 ;
  assign n2203 = n2202 ^ n2196 ;
  assign n2204 = n2203 ^ n2201 ;
  assign n2205 = n236 & ~n2204 ;
  assign n2206 = n2205 ^ n236 ;
  assign n2220 = n2219 ^ n2206 ;
  assign n2239 = n148 & n1446 ;
  assign n2236 = n137 & n1535 ;
  assign n2237 = n2236 ^ n137 ;
  assign n2238 = n2237 ^ n137 ;
  assign n2240 = n2239 ^ n2238 ;
  assign n2244 = n171 & n1548 ;
  assign n2241 = n160 & n1521 ;
  assign n2242 = n2241 ^ n160 ;
  assign n2243 = n2242 ^ n160 ;
  assign n2245 = n2244 ^ n2243 ;
  assign n2246 = n2240 & n2245 ;
  assign n2247 = n2246 ^ n2240 ;
  assign n2248 = n2247 ^ n2245 ;
  assign n2249 = n136 & n2248 ;
  assign n2224 = n148 & n1560 ;
  assign n2221 = n137 & n1590 ;
  assign n2222 = n2221 ^ n137 ;
  assign n2223 = n2222 ^ n137 ;
  assign n2225 = n2224 ^ n2223 ;
  assign n2229 = n171 & n1603 ;
  assign n2226 = n160 & n1578 ;
  assign n2227 = n2226 ^ n160 ;
  assign n2228 = n2227 ^ n160 ;
  assign n2230 = n2229 ^ n2228 ;
  assign n2231 = n2225 & n2230 ;
  assign n2232 = n2231 ^ n2225 ;
  assign n2233 = n2232 ^ n2230 ;
  assign n2234 = n188 & ~n2233 ;
  assign n2235 = n2234 ^ n188 ;
  assign n2250 = n2249 ^ n2235 ;
  assign n2251 = n2220 & n2250 ;
  assign n2252 = n2251 ^ n2220 ;
  assign n2253 = n2252 ^ n2250 ;
  assign n2317 = n2316 ^ n2253 ;
  assign n2318 = x134 & n2317 ;
  assign n2319 = n2318 ^ n2317 ;
  assign n2320 = n2319 ^ n2253 ;
  assign n2387 = n148 & n376 ;
  assign n2386 = n137 & n386 ;
  assign n2388 = n2387 ^ n2386 ;
  assign n2390 = n171 & n402 ;
  assign n2389 = n160 & n412 ;
  assign n2391 = n2390 ^ n2389 ;
  assign n2392 = n2388 & n2391 ;
  assign n2393 = n2392 ^ n2388 ;
  assign n2394 = n2393 ^ n2391 ;
  assign n2395 = n188 & n2394 ;
  assign n2376 = n148 & n470 ;
  assign n2375 = n137 & n480 ;
  assign n2377 = n2376 ^ n2375 ;
  assign n2379 = n171 & n355 ;
  assign n2378 = n160 & n365 ;
  assign n2380 = n2379 ^ n2378 ;
  assign n2381 = n2377 & n2380 ;
  assign n2382 = n2381 ^ n2377 ;
  assign n2383 = n2382 ^ n2380 ;
  assign n2384 = n136 & ~n2383 ;
  assign n2385 = n2384 ^ n136 ;
  assign n2396 = n2395 ^ n2385 ;
  assign n2409 = n148 & n218 ;
  assign n2408 = n137 & n228 ;
  assign n2410 = n2409 ^ n2408 ;
  assign n2412 = n171 & n496 ;
  assign n2411 = n160 & n507 ;
  assign n2413 = n2412 ^ n2411 ;
  assign n2414 = n2410 & n2413 ;
  assign n2415 = n2414 ^ n2410 ;
  assign n2416 = n2415 ^ n2413 ;
  assign n2417 = n236 & n2416 ;
  assign n2398 = n148 & n518 ;
  assign n2397 = n137 & n528 ;
  assign n2399 = n2398 ^ n2397 ;
  assign n2401 = n171 & n449 ;
  assign n2400 = n160 & n459 ;
  assign n2402 = n2401 ^ n2400 ;
  assign n2403 = n2399 & n2402 ;
  assign n2404 = n2403 ^ n2399 ;
  assign n2405 = n2404 ^ n2402 ;
  assign n2406 = n314 & ~n2405 ;
  assign n2407 = n2406 ^ n314 ;
  assign n2418 = n2417 ^ n2407 ;
  assign n2419 = n2396 & n2418 ;
  assign n2420 = n2419 ^ n2396 ;
  assign n2421 = n2420 ^ n2418 ;
  assign n2333 = n148 & n266 ;
  assign n2332 = n137 & n276 ;
  assign n2334 = n2333 ^ n2332 ;
  assign n2336 = n171 & n323 ;
  assign n2335 = n160 & n333 ;
  assign n2337 = n2336 ^ n2335 ;
  assign n2338 = n2334 & n2337 ;
  assign n2339 = n2338 ^ n2334 ;
  assign n2340 = n2339 ^ n2337 ;
  assign n2341 = n314 & n2340 ;
  assign n2322 = n148 & n423 ;
  assign n2321 = n137 & n433 ;
  assign n2323 = n2322 ^ n2321 ;
  assign n2325 = n171 & n245 ;
  assign n2324 = n160 & n255 ;
  assign n2326 = n2325 ^ n2324 ;
  assign n2327 = n2323 & n2326 ;
  assign n2328 = n2327 ^ n2323 ;
  assign n2329 = n2328 ^ n2326 ;
  assign n2330 = n236 & ~n2329 ;
  assign n2331 = n2330 ^ n236 ;
  assign n2342 = n2341 ^ n2331 ;
  assign n2347 = n148 & n299 ;
  assign n2346 = n137 & n311 ;
  assign n2348 = n2347 ^ n2346 ;
  assign n2344 = n146 & n171 ;
  assign n2343 = n157 & n160 ;
  assign n2345 = n2344 ^ n2343 ;
  assign n2349 = n2348 ^ n2345 ;
  assign n2350 = n2345 ^ n136 ;
  assign n2351 = n136 & n2350 ;
  assign n2352 = n2351 ^ n2350 ;
  assign n2353 = n2352 ^ n136 ;
  assign n2354 = n2353 ^ n2348 ;
  assign n2355 = n2349 & n2354 ;
  assign n2356 = n2355 ^ n2352 ;
  assign n2357 = n2356 ^ n2348 ;
  assign n2359 = n137 & n180 ;
  assign n2358 = n148 & n169 ;
  assign n2360 = n2359 ^ n2358 ;
  assign n2362 = n171 & n197 ;
  assign n2361 = n160 & n207 ;
  assign n2363 = n2362 ^ n2361 ;
  assign n2364 = n2360 & n2363 ;
  assign n2365 = n2364 ^ n2360 ;
  assign n2366 = n2365 ^ n2363 ;
  assign n2367 = n188 & ~n2366 ;
  assign n2368 = n2367 ^ n188 ;
  assign n2369 = n2357 & n2368 ;
  assign n2370 = n2369 ^ n2357 ;
  assign n2371 = n2370 ^ n2368 ;
  assign n2372 = n2342 & n2371 ;
  assign n2373 = n2372 ^ n2342 ;
  assign n2374 = n2373 ^ n2371 ;
  assign n2422 = n2421 ^ n2374 ;
  assign n2423 = x134 & n2422 ;
  assign n2424 = n2423 ^ n2422 ;
  assign n2425 = n2424 ^ n2374 ;
  assign n2507 = n148 & n900 ;
  assign n2504 = n137 & n919 ;
  assign n2505 = n2504 ^ n137 ;
  assign n2506 = n2505 ^ n137 ;
  assign n2508 = n2507 ^ n2506 ;
  assign n2512 = n171 & n942 ;
  assign n2509 = n160 & n961 ;
  assign n2510 = n2509 ^ n160 ;
  assign n2511 = n2510 ^ n160 ;
  assign n2513 = n2512 ^ n2511 ;
  assign n2514 = n2508 & n2513 ;
  assign n2515 = n2514 ^ n2508 ;
  assign n2516 = n2515 ^ n2513 ;
  assign n2517 = n188 & n2516 ;
  assign n2492 = n148 & n1058 ;
  assign n2489 = n137 & n1077 ;
  assign n2490 = n2489 ^ n137 ;
  assign n2491 = n2490 ^ n137 ;
  assign n2493 = n2492 ^ n2491 ;
  assign n2497 = n171 & n863 ;
  assign n2494 = n160 & n882 ;
  assign n2495 = n2494 ^ n160 ;
  assign n2496 = n2495 ^ n160 ;
  assign n2498 = n2497 ^ n2496 ;
  assign n2499 = n2493 & n2498 ;
  assign n2500 = n2499 ^ n2493 ;
  assign n2501 = n2500 ^ n2498 ;
  assign n2502 = n136 & ~n2501 ;
  assign n2503 = n2502 ^ n136 ;
  assign n2518 = n2517 ^ n2503 ;
  assign n2537 = n148 & n595 ;
  assign n2534 = n137 & n614 ;
  assign n2535 = n2534 ^ n137 ;
  assign n2536 = n2535 ^ n137 ;
  assign n2538 = n2537 ^ n2536 ;
  assign n2542 = n171 & n1100 ;
  assign n2539 = n160 & n1119 ;
  assign n2540 = n2539 ^ n160 ;
  assign n2541 = n2540 ^ n160 ;
  assign n2543 = n2542 ^ n2541 ;
  assign n2544 = n2538 & n2543 ;
  assign n2545 = n2544 ^ n2538 ;
  assign n2546 = n2545 ^ n2543 ;
  assign n2547 = n236 & n2546 ;
  assign n2522 = n148 & n1137 ;
  assign n2519 = n137 & n1156 ;
  assign n2520 = n2519 ^ n137 ;
  assign n2521 = n2520 ^ n137 ;
  assign n2523 = n2522 ^ n2521 ;
  assign n2527 = n171 & n1021 ;
  assign n2524 = n160 & n1040 ;
  assign n2525 = n2524 ^ n160 ;
  assign n2526 = n2525 ^ n160 ;
  assign n2528 = n2527 ^ n2526 ;
  assign n2529 = n2523 & n2528 ;
  assign n2530 = n2529 ^ n2523 ;
  assign n2531 = n2530 ^ n2528 ;
  assign n2532 = n314 & ~n2531 ;
  assign n2533 = n2532 ^ n314 ;
  assign n2548 = n2547 ^ n2533 ;
  assign n2549 = n2518 & n2548 ;
  assign n2550 = n2549 ^ n2518 ;
  assign n2551 = n2550 ^ n2548 ;
  assign n2444 = n148 & n674 ;
  assign n2441 = n137 & n693 ;
  assign n2442 = n2441 ^ n137 ;
  assign n2443 = n2442 ^ n137 ;
  assign n2445 = n2444 ^ n2443 ;
  assign n2447 = n160 & n808 ;
  assign n2448 = n2447 ^ n160 ;
  assign n2449 = n2448 ^ n160 ;
  assign n2446 = n171 & n790 ;
  assign n2450 = n2449 ^ n2446 ;
  assign n2451 = n2445 & n2450 ;
  assign n2452 = n2451 ^ n2445 ;
  assign n2453 = n2452 ^ n2450 ;
  assign n2454 = n314 & n2453 ;
  assign n2429 = n148 & n979 ;
  assign n2426 = n137 & n998 ;
  assign n2427 = n2426 ^ n137 ;
  assign n2428 = n2427 ^ n137 ;
  assign n2430 = n2429 ^ n2428 ;
  assign n2434 = n171 & n637 ;
  assign n2431 = n160 & n656 ;
  assign n2432 = n2431 ^ n160 ;
  assign n2433 = n2432 ^ n160 ;
  assign n2435 = n2434 ^ n2433 ;
  assign n2436 = n2430 & n2435 ;
  assign n2437 = n2436 ^ n2430 ;
  assign n2438 = n2437 ^ n2435 ;
  assign n2439 = n236 & ~n2438 ;
  assign n2440 = n2439 ^ n236 ;
  assign n2455 = n2454 ^ n2440 ;
  assign n2472 = n137 & n837 ;
  assign n2473 = n2472 ^ n137 ;
  assign n2474 = n2473 ^ n137 ;
  assign n2471 = n148 & n820 ;
  assign n2475 = n2474 ^ n2471 ;
  assign n2479 = n171 & n716 ;
  assign n2476 = n160 & n735 ;
  assign n2477 = n2476 ^ n160 ;
  assign n2478 = n2477 ^ n160 ;
  assign n2480 = n2479 ^ n2478 ;
  assign n2481 = n2475 & n2480 ;
  assign n2482 = n2481 ^ n2475 ;
  assign n2483 = n2482 ^ n2480 ;
  assign n2484 = n136 & n2483 ;
  assign n2459 = n148 & n753 ;
  assign n2456 = n137 & n772 ;
  assign n2457 = n2456 ^ n137 ;
  assign n2458 = n2457 ^ n137 ;
  assign n2460 = n2459 ^ n2458 ;
  assign n2464 = n171 & n558 ;
  assign n2461 = n160 & n577 ;
  assign n2462 = n2461 ^ n160 ;
  assign n2463 = n2462 ^ n160 ;
  assign n2465 = n2464 ^ n2463 ;
  assign n2466 = n2460 & n2465 ;
  assign n2467 = n2466 ^ n2460 ;
  assign n2468 = n2467 ^ n2465 ;
  assign n2469 = n188 & ~n2468 ;
  assign n2470 = n2469 ^ n188 ;
  assign n2485 = n2484 ^ n2470 ;
  assign n2486 = n2455 & n2485 ;
  assign n2487 = n2486 ^ n2455 ;
  assign n2488 = n2487 ^ n2485 ;
  assign n2552 = n2551 ^ n2488 ;
  assign n2553 = x134 & n2552 ;
  assign n2554 = n2553 ^ n2552 ;
  assign n2555 = n2554 ^ n2488 ;
  assign n2617 = n148 & n1301 ;
  assign n2616 = n137 & n1305 ;
  assign n2618 = n2617 ^ n2616 ;
  assign n2620 = n171 & n1316 ;
  assign n2619 = n160 & n1320 ;
  assign n2621 = n2620 ^ n2619 ;
  assign n2622 = n2618 & n2621 ;
  assign n2623 = n2622 ^ n2618 ;
  assign n2624 = n2623 ^ n2621 ;
  assign n2625 = n188 & n2624 ;
  assign n2606 = n148 & n1352 ;
  assign n2605 = n137 & n1356 ;
  assign n2607 = n2606 ^ n2605 ;
  assign n2609 = n171 & n1291 ;
  assign n2608 = n160 & n1295 ;
  assign n2610 = n2609 ^ n2608 ;
  assign n2611 = n2607 & n2610 ;
  assign n2612 = n2611 ^ n2607 ;
  assign n2613 = n2612 ^ n2610 ;
  assign n2614 = n136 & ~n2613 ;
  assign n2615 = n2614 ^ n136 ;
  assign n2626 = n2625 ^ n2615 ;
  assign n2639 = n148 & n1184 ;
  assign n2638 = n137 & n1188 ;
  assign n2640 = n2639 ^ n2638 ;
  assign n2642 = n171 & n1367 ;
  assign n2641 = n160 & n1371 ;
  assign n2643 = n2642 ^ n2641 ;
  assign n2644 = n2640 & n2643 ;
  assign n2645 = n2644 ^ n2640 ;
  assign n2646 = n2645 ^ n2643 ;
  assign n2647 = n236 & n2646 ;
  assign n2628 = n148 & n1377 ;
  assign n2627 = n137 & n1381 ;
  assign n2629 = n2628 ^ n2627 ;
  assign n2631 = n171 & n1341 ;
  assign n2630 = n160 & n1346 ;
  assign n2632 = n2631 ^ n2630 ;
  assign n2633 = n2629 & n2632 ;
  assign n2634 = n2633 ^ n2629 ;
  assign n2635 = n2634 ^ n2632 ;
  assign n2636 = n314 & ~n2635 ;
  assign n2637 = n2636 ^ n314 ;
  assign n2648 = n2647 ^ n2637 ;
  assign n2649 = n2626 & n2648 ;
  assign n2650 = n2649 ^ n2626 ;
  assign n2651 = n2650 ^ n2648 ;
  assign n2568 = n148 & n1210 ;
  assign n2567 = n137 & n1214 ;
  assign n2569 = n2568 ^ n2567 ;
  assign n2571 = n171 & n1250 ;
  assign n2570 = n160 & n1255 ;
  assign n2572 = n2571 ^ n2570 ;
  assign n2573 = n2569 & n2572 ;
  assign n2574 = n2573 ^ n2569 ;
  assign n2575 = n2574 ^ n2572 ;
  assign n2576 = n314 & n2575 ;
  assign n2557 = n148 & n1326 ;
  assign n2556 = n137 & n1330 ;
  assign n2558 = n2557 ^ n2556 ;
  assign n2560 = n171 & n1199 ;
  assign n2559 = n160 & n1204 ;
  assign n2561 = n2560 ^ n2559 ;
  assign n2562 = n2558 & n2561 ;
  assign n2563 = n2562 ^ n2558 ;
  assign n2564 = n2563 ^ n2561 ;
  assign n2565 = n236 & ~n2564 ;
  assign n2566 = n2565 ^ n236 ;
  assign n2577 = n2576 ^ n2566 ;
  assign n2592 = n148 & n1266 ;
  assign n2589 = n137 & n1277 ;
  assign n2590 = n2589 ^ n137 ;
  assign n2591 = n2590 ^ n137 ;
  assign n2593 = n2592 ^ n2591 ;
  assign n2595 = n171 & n1225 ;
  assign n2594 = n160 & n1229 ;
  assign n2596 = n2595 ^ n2594 ;
  assign n2597 = n2593 & n2596 ;
  assign n2598 = n2597 ^ n2593 ;
  assign n2599 = n2598 ^ n2596 ;
  assign n2600 = n136 & n2599 ;
  assign n2579 = n148 & n1235 ;
  assign n2578 = n137 & n1239 ;
  assign n2580 = n2579 ^ n2578 ;
  assign n2582 = n171 & n1174 ;
  assign n2581 = n160 & n1178 ;
  assign n2583 = n2582 ^ n2581 ;
  assign n2584 = n2580 & n2583 ;
  assign n2585 = n2584 ^ n2580 ;
  assign n2586 = n2585 ^ n2583 ;
  assign n2587 = n188 & ~n2586 ;
  assign n2588 = n2587 ^ n188 ;
  assign n2601 = n2600 ^ n2588 ;
  assign n2602 = n2577 & n2601 ;
  assign n2603 = n2602 ^ n2577 ;
  assign n2604 = n2603 ^ n2601 ;
  assign n2652 = n2651 ^ n2604 ;
  assign n2653 = x134 & n2652 ;
  assign n2654 = n2653 ^ n2652 ;
  assign n2655 = n2654 ^ n2604 ;
  assign n2737 = n148 & n1661 ;
  assign n2734 = n137 & n1673 ;
  assign n2735 = n2734 ^ n137 ;
  assign n2736 = n2735 ^ n137 ;
  assign n2738 = n2737 ^ n2736 ;
  assign n2742 = n171 & n1748 ;
  assign n2739 = n160 & n1760 ;
  assign n2740 = n2739 ^ n160 ;
  assign n2741 = n2740 ^ n160 ;
  assign n2743 = n2742 ^ n2741 ;
  assign n2744 = n2738 & n2743 ;
  assign n2745 = n2744 ^ n2738 ;
  assign n2746 = n2745 ^ n2743 ;
  assign n2747 = n188 & n2746 ;
  assign n2722 = n148 & n1718 ;
  assign n2719 = n137 & n1730 ;
  assign n2720 = n2719 ^ n137 ;
  assign n2721 = n2720 ^ n137 ;
  assign n2723 = n2722 ^ n2721 ;
  assign n2727 = n171 & n1636 ;
  assign n2724 = n160 & n1648 ;
  assign n2725 = n2724 ^ n160 ;
  assign n2726 = n2725 ^ n160 ;
  assign n2728 = n2727 ^ n2726 ;
  assign n2729 = n2723 & n2728 ;
  assign n2730 = n2729 ^ n2723 ;
  assign n2731 = n2730 ^ n2728 ;
  assign n2732 = n136 & ~n2731 ;
  assign n2733 = n2732 ^ n136 ;
  assign n2748 = n2747 ^ n2733 ;
  assign n2767 = n148 & n1603 ;
  assign n2764 = n137 & n1615 ;
  assign n2765 = n2764 ^ n137 ;
  assign n2766 = n2765 ^ n137 ;
  assign n2768 = n2767 ^ n2766 ;
  assign n2772 = n171 & n1803 ;
  assign n2769 = n160 & n1815 ;
  assign n2770 = n2769 ^ n160 ;
  assign n2771 = n2770 ^ n160 ;
  assign n2773 = n2772 ^ n2771 ;
  assign n2774 = n2768 & n2773 ;
  assign n2775 = n2774 ^ n2768 ;
  assign n2776 = n2775 ^ n2773 ;
  assign n2777 = n236 & n2776 ;
  assign n2752 = n148 & n1828 ;
  assign n2749 = n137 & n1840 ;
  assign n2750 = n2749 ^ n137 ;
  assign n2751 = n2750 ^ n137 ;
  assign n2753 = n2752 ^ n2751 ;
  assign n2757 = n171 & n1691 ;
  assign n2754 = n160 & n1705 ;
  assign n2755 = n2754 ^ n160 ;
  assign n2756 = n2755 ^ n160 ;
  assign n2758 = n2757 ^ n2756 ;
  assign n2759 = n2753 & n2758 ;
  assign n2760 = n2759 ^ n2753 ;
  assign n2761 = n2760 ^ n2758 ;
  assign n2762 = n314 & ~n2761 ;
  assign n2763 = n2762 ^ n314 ;
  assign n2778 = n2777 ^ n2763 ;
  assign n2779 = n2748 & n2778 ;
  assign n2780 = n2779 ^ n2748 ;
  assign n2781 = n2780 ^ n2778 ;
  assign n2674 = n148 & n1491 ;
  assign n2671 = n160 & n1415 ;
  assign n2672 = n2671 ^ n160 ;
  assign n2673 = n2672 ^ n160 ;
  assign n2675 = n2674 ^ n2673 ;
  assign n2677 = n137 & n1503 ;
  assign n2678 = n2677 ^ n137 ;
  assign n2679 = n2678 ^ n137 ;
  assign n2676 = n171 & n1402 ;
  assign n2680 = n2679 ^ n2676 ;
  assign n2681 = n2675 & n2680 ;
  assign n2682 = n2681 ^ n2675 ;
  assign n2683 = n2682 ^ n2680 ;
  assign n2684 = n314 & n2683 ;
  assign n2659 = n148 & n1773 ;
  assign n2656 = n137 & n1785 ;
  assign n2657 = n2656 ^ n137 ;
  assign n2658 = n2657 ^ n137 ;
  assign n2660 = n2659 ^ n2658 ;
  assign n2664 = n171 & n1464 ;
  assign n2661 = n160 & n1478 ;
  assign n2662 = n2661 ^ n160 ;
  assign n2663 = n2662 ^ n160 ;
  assign n2665 = n2664 ^ n2663 ;
  assign n2666 = n2660 & n2665 ;
  assign n2667 = n2666 ^ n2660 ;
  assign n2668 = n2667 ^ n2665 ;
  assign n2669 = n236 & ~n2668 ;
  assign n2670 = n2669 ^ n236 ;
  assign n2685 = n2684 ^ n2670 ;
  assign n2704 = n148 & n1433 ;
  assign n2701 = n137 & n1446 ;
  assign n2702 = n2701 ^ n137 ;
  assign n2703 = n2702 ^ n137 ;
  assign n2705 = n2704 ^ n2703 ;
  assign n2709 = n171 & n1521 ;
  assign n2706 = n160 & n1535 ;
  assign n2707 = n2706 ^ n160 ;
  assign n2708 = n2707 ^ n160 ;
  assign n2710 = n2709 ^ n2708 ;
  assign n2711 = n2705 & n2710 ;
  assign n2712 = n2711 ^ n2705 ;
  assign n2713 = n2712 ^ n2710 ;
  assign n2714 = n136 & n2713 ;
  assign n2689 = n148 & n1548 ;
  assign n2686 = n137 & n1560 ;
  assign n2687 = n2686 ^ n137 ;
  assign n2688 = n2687 ^ n137 ;
  assign n2690 = n2689 ^ n2688 ;
  assign n2694 = n171 & n1578 ;
  assign n2691 = n160 & n1590 ;
  assign n2692 = n2691 ^ n160 ;
  assign n2693 = n2692 ^ n160 ;
  assign n2695 = n2694 ^ n2693 ;
  assign n2696 = n2690 & n2695 ;
  assign n2697 = n2696 ^ n2690 ;
  assign n2698 = n2697 ^ n2695 ;
  assign n2699 = n188 & ~n2698 ;
  assign n2700 = n2699 ^ n188 ;
  assign n2715 = n2714 ^ n2700 ;
  assign n2716 = n2685 & n2715 ;
  assign n2717 = n2716 ^ n2685 ;
  assign n2718 = n2717 ^ n2715 ;
  assign n2782 = n2781 ^ n2718 ;
  assign n2783 = x134 & n2782 ;
  assign n2784 = n2783 ^ n2782 ;
  assign n2785 = n2784 ^ n2718 ;
  assign n2854 = n148 & n355 ;
  assign n2853 = n137 & n376 ;
  assign n2855 = n2854 ^ n2853 ;
  assign n2857 = n171 & n412 ;
  assign n2856 = n160 & n386 ;
  assign n2858 = n2857 ^ n2856 ;
  assign n2859 = n2855 & n2858 ;
  assign n2860 = n2859 ^ n2855 ;
  assign n2861 = n2860 ^ n2858 ;
  assign n2862 = n188 & n2861 ;
  assign n2843 = n148 & n449 ;
  assign n2842 = n137 & n470 ;
  assign n2844 = n2843 ^ n2842 ;
  assign n2846 = n171 & n365 ;
  assign n2845 = n160 & n480 ;
  assign n2847 = n2846 ^ n2845 ;
  assign n2848 = n2844 & n2847 ;
  assign n2849 = n2848 ^ n2844 ;
  assign n2850 = n2849 ^ n2847 ;
  assign n2851 = n136 & ~n2850 ;
  assign n2852 = n2851 ^ n136 ;
  assign n2863 = n2862 ^ n2852 ;
  assign n2876 = n148 & n197 ;
  assign n2875 = n137 & n218 ;
  assign n2877 = n2876 ^ n2875 ;
  assign n2879 = n171 & n507 ;
  assign n2878 = n160 & n228 ;
  assign n2880 = n2879 ^ n2878 ;
  assign n2881 = n2877 & n2880 ;
  assign n2882 = n2881 ^ n2877 ;
  assign n2883 = n2882 ^ n2880 ;
  assign n2884 = n236 & n2883 ;
  assign n2865 = n148 & n496 ;
  assign n2864 = n137 & n518 ;
  assign n2866 = n2865 ^ n2864 ;
  assign n2868 = n171 & n459 ;
  assign n2867 = n160 & n528 ;
  assign n2869 = n2868 ^ n2867 ;
  assign n2870 = n2866 & n2869 ;
  assign n2871 = n2870 ^ n2866 ;
  assign n2872 = n2871 ^ n2869 ;
  assign n2873 = n314 & ~n2872 ;
  assign n2874 = n2873 ^ n314 ;
  assign n2885 = n2884 ^ n2874 ;
  assign n2886 = n2863 & n2885 ;
  assign n2887 = n2886 ^ n2863 ;
  assign n2888 = n2887 ^ n2885 ;
  assign n2798 = n148 & n245 ;
  assign n2797 = n137 & n266 ;
  assign n2799 = n2798 ^ n2797 ;
  assign n2801 = n171 & n333 ;
  assign n2800 = n160 & n276 ;
  assign n2802 = n2801 ^ n2800 ;
  assign n2803 = n2799 & n2802 ;
  assign n2804 = n2803 ^ n2799 ;
  assign n2805 = n2804 ^ n2802 ;
  assign n2806 = n314 & n2805 ;
  assign n2787 = n148 & n402 ;
  assign n2786 = n137 & n423 ;
  assign n2788 = n2787 ^ n2786 ;
  assign n2790 = n171 & n255 ;
  assign n2789 = n160 & n433 ;
  assign n2791 = n2790 ^ n2789 ;
  assign n2792 = n2788 & n2791 ;
  assign n2793 = n2792 ^ n2788 ;
  assign n2794 = n2793 ^ n2791 ;
  assign n2795 = n236 & ~n2794 ;
  assign n2796 = n2795 ^ n236 ;
  assign n2807 = n2806 ^ n2796 ;
  assign n2814 = n148 & n323 ;
  assign n2811 = n137 & n299 ;
  assign n2812 = n2811 ^ n137 ;
  assign n2813 = n2812 ^ n137 ;
  assign n2815 = n2814 ^ n2813 ;
  assign n2809 = n157 & n171 ;
  assign n2808 = n160 & n311 ;
  assign n2810 = n2809 ^ n2808 ;
  assign n2816 = n2815 ^ n2810 ;
  assign n2817 = n2810 ^ n136 ;
  assign n2818 = n136 & n2817 ;
  assign n2819 = n2818 ^ n2817 ;
  assign n2820 = n2819 ^ n136 ;
  assign n2821 = n2820 ^ n2815 ;
  assign n2822 = n2816 & n2821 ;
  assign n2823 = n2822 ^ n2819 ;
  assign n2824 = n2823 ^ n2815 ;
  assign n2826 = n146 & n148 ;
  assign n2825 = n137 & n169 ;
  assign n2827 = n2826 ^ n2825 ;
  assign n2829 = n171 & n207 ;
  assign n2828 = n160 & n180 ;
  assign n2830 = n2829 ^ n2828 ;
  assign n2831 = n2827 & n2830 ;
  assign n2832 = n2831 ^ n2827 ;
  assign n2833 = n2832 ^ n2830 ;
  assign n2834 = n188 & ~n2833 ;
  assign n2835 = n2834 ^ n188 ;
  assign n2836 = n2824 & n2835 ;
  assign n2837 = n2836 ^ n2824 ;
  assign n2838 = n2837 ^ n2835 ;
  assign n2839 = n2807 & n2838 ;
  assign n2840 = n2839 ^ n2807 ;
  assign n2841 = n2840 ^ n2838 ;
  assign n2889 = n2888 ^ n2841 ;
  assign n2890 = x134 & n2889 ;
  assign n2891 = n2890 ^ n2889 ;
  assign n2892 = n2891 ^ n2841 ;
  assign n2978 = n148 & n863 ;
  assign n2975 = n137 & n900 ;
  assign n2976 = n2975 ^ n137 ;
  assign n2977 = n2976 ^ n137 ;
  assign n2979 = n2978 ^ n2977 ;
  assign n2983 = n171 & n961 ;
  assign n2980 = n160 & n919 ;
  assign n2981 = n2980 ^ n160 ;
  assign n2982 = n2981 ^ n160 ;
  assign n2984 = n2983 ^ n2982 ;
  assign n2985 = n2979 & n2984 ;
  assign n2986 = n2985 ^ n2979 ;
  assign n2987 = n2986 ^ n2984 ;
  assign n2988 = n188 & n2987 ;
  assign n2963 = n148 & n1021 ;
  assign n2960 = n137 & n1058 ;
  assign n2961 = n2960 ^ n137 ;
  assign n2962 = n2961 ^ n137 ;
  assign n2964 = n2963 ^ n2962 ;
  assign n2968 = n171 & n882 ;
  assign n2965 = n160 & n1077 ;
  assign n2966 = n2965 ^ n160 ;
  assign n2967 = n2966 ^ n160 ;
  assign n2969 = n2968 ^ n2967 ;
  assign n2970 = n2964 & n2969 ;
  assign n2971 = n2970 ^ n2964 ;
  assign n2972 = n2971 ^ n2969 ;
  assign n2973 = n136 & ~n2972 ;
  assign n2974 = n2973 ^ n136 ;
  assign n2989 = n2988 ^ n2974 ;
  assign n3008 = n148 & n558 ;
  assign n3005 = n137 & n595 ;
  assign n3006 = n3005 ^ n137 ;
  assign n3007 = n3006 ^ n137 ;
  assign n3009 = n3008 ^ n3007 ;
  assign n3013 = n171 & n1119 ;
  assign n3010 = n160 & n614 ;
  assign n3011 = n3010 ^ n160 ;
  assign n3012 = n3011 ^ n160 ;
  assign n3014 = n3013 ^ n3012 ;
  assign n3015 = n3009 & n3014 ;
  assign n3016 = n3015 ^ n3009 ;
  assign n3017 = n3016 ^ n3014 ;
  assign n3018 = n236 & n3017 ;
  assign n2993 = n148 & n1100 ;
  assign n2990 = n137 & n1137 ;
  assign n2991 = n2990 ^ n137 ;
  assign n2992 = n2991 ^ n137 ;
  assign n2994 = n2993 ^ n2992 ;
  assign n2998 = n171 & n1040 ;
  assign n2995 = n160 & n1156 ;
  assign n2996 = n2995 ^ n160 ;
  assign n2997 = n2996 ^ n160 ;
  assign n2999 = n2998 ^ n2997 ;
  assign n3000 = n2994 & n2999 ;
  assign n3001 = n3000 ^ n2994 ;
  assign n3002 = n3001 ^ n2999 ;
  assign n3003 = n314 & ~n3002 ;
  assign n3004 = n3003 ^ n314 ;
  assign n3019 = n3018 ^ n3004 ;
  assign n3020 = n2989 & n3019 ;
  assign n3021 = n3020 ^ n2989 ;
  assign n3022 = n3021 ^ n3019 ;
  assign n2911 = n148 & n637 ;
  assign n2908 = n137 & n674 ;
  assign n2909 = n2908 ^ n137 ;
  assign n2910 = n2909 ^ n137 ;
  assign n2912 = n2911 ^ n2910 ;
  assign n2916 = n171 & n808 ;
  assign n2913 = n160 & n693 ;
  assign n2914 = n2913 ^ n160 ;
  assign n2915 = n2914 ^ n160 ;
  assign n2917 = n2916 ^ n2915 ;
  assign n2918 = n2912 & n2917 ;
  assign n2919 = n2918 ^ n2912 ;
  assign n2920 = n2919 ^ n2917 ;
  assign n2921 = n314 & n2920 ;
  assign n2896 = n148 & n942 ;
  assign n2893 = n137 & n979 ;
  assign n2894 = n2893 ^ n137 ;
  assign n2895 = n2894 ^ n137 ;
  assign n2897 = n2896 ^ n2895 ;
  assign n2901 = n171 & n656 ;
  assign n2898 = n160 & n998 ;
  assign n2899 = n2898 ^ n160 ;
  assign n2900 = n2899 ^ n160 ;
  assign n2902 = n2901 ^ n2900 ;
  assign n2903 = n2897 & n2902 ;
  assign n2904 = n2903 ^ n2897 ;
  assign n2905 = n2904 ^ n2902 ;
  assign n2906 = n236 & ~n2905 ;
  assign n2907 = n2906 ^ n236 ;
  assign n2922 = n2921 ^ n2907 ;
  assign n2926 = n171 & n735 ;
  assign n2923 = n160 & n837 ;
  assign n2924 = n2923 ^ n160 ;
  assign n2925 = n2924 ^ n160 ;
  assign n2927 = n2926 ^ n2925 ;
  assign n2931 = n148 & n790 ;
  assign n2928 = n137 & n820 ;
  assign n2929 = n2928 ^ n137 ;
  assign n2930 = n2929 ^ n137 ;
  assign n2932 = n2931 ^ n2930 ;
  assign n2933 = n136 & n2932 ;
  assign n2934 = n2933 ^ n136 ;
  assign n2935 = n2927 & n2934 ;
  assign n2936 = n2935 ^ n2934 ;
  assign n2937 = n2936 ^ n136 ;
  assign n2941 = n148 & n716 ;
  assign n2938 = n137 & n753 ;
  assign n2939 = n2938 ^ n137 ;
  assign n2940 = n2939 ^ n137 ;
  assign n2942 = n2941 ^ n2940 ;
  assign n2946 = n171 & n577 ;
  assign n2943 = n160 & n772 ;
  assign n2944 = n2943 ^ n160 ;
  assign n2945 = n2944 ^ n160 ;
  assign n2947 = n2946 ^ n2945 ;
  assign n2948 = n2942 & n2947 ;
  assign n2949 = n2948 ^ n2942 ;
  assign n2950 = n2949 ^ n2947 ;
  assign n2951 = n188 & n2950 ;
  assign n2952 = n2951 ^ n188 ;
  assign n2953 = n2952 ^ n188 ;
  assign n2954 = n2937 & n2953 ;
  assign n2955 = n2954 ^ n2937 ;
  assign n2956 = n2955 ^ n2953 ;
  assign n2957 = n2922 & n2956 ;
  assign n2958 = n2957 ^ n2922 ;
  assign n2959 = n2958 ^ n2956 ;
  assign n3023 = n3022 ^ n2959 ;
  assign n3024 = x134 & n3023 ;
  assign n3025 = n3024 ^ n3023 ;
  assign n3026 = n3025 ^ n2959 ;
  assign n3090 = n148 & n1291 ;
  assign n3089 = n137 & n1301 ;
  assign n3091 = n3090 ^ n3089 ;
  assign n3093 = n171 & n1320 ;
  assign n3092 = n160 & n1305 ;
  assign n3094 = n3093 ^ n3092 ;
  assign n3095 = n3091 & n3094 ;
  assign n3096 = n3095 ^ n3091 ;
  assign n3097 = n3096 ^ n3094 ;
  assign n3098 = n188 & n3097 ;
  assign n3079 = n148 & n1341 ;
  assign n3078 = n137 & n1352 ;
  assign n3080 = n3079 ^ n3078 ;
  assign n3082 = n171 & n1295 ;
  assign n3081 = n160 & n1356 ;
  assign n3083 = n3082 ^ n3081 ;
  assign n3084 = n3080 & n3083 ;
  assign n3085 = n3084 ^ n3080 ;
  assign n3086 = n3085 ^ n3083 ;
  assign n3087 = n136 & ~n3086 ;
  assign n3088 = n3087 ^ n136 ;
  assign n3099 = n3098 ^ n3088 ;
  assign n3112 = n148 & n1174 ;
  assign n3111 = n137 & n1184 ;
  assign n3113 = n3112 ^ n3111 ;
  assign n3115 = n171 & n1371 ;
  assign n3114 = n160 & n1188 ;
  assign n3116 = n3115 ^ n3114 ;
  assign n3117 = n3113 & n3116 ;
  assign n3118 = n3117 ^ n3113 ;
  assign n3119 = n3118 ^ n3116 ;
  assign n3120 = n236 & n3119 ;
  assign n3101 = n148 & n1367 ;
  assign n3100 = n137 & n1377 ;
  assign n3102 = n3101 ^ n3100 ;
  assign n3104 = n171 & n1346 ;
  assign n3103 = n160 & n1381 ;
  assign n3105 = n3104 ^ n3103 ;
  assign n3106 = n3102 & n3105 ;
  assign n3107 = n3106 ^ n3102 ;
  assign n3108 = n3107 ^ n3105 ;
  assign n3109 = n314 & ~n3108 ;
  assign n3110 = n3109 ^ n314 ;
  assign n3121 = n3120 ^ n3110 ;
  assign n3122 = n3099 & n3121 ;
  assign n3123 = n3122 ^ n3099 ;
  assign n3124 = n3123 ^ n3121 ;
  assign n3039 = n148 & n1199 ;
  assign n3038 = n137 & n1210 ;
  assign n3040 = n3039 ^ n3038 ;
  assign n3042 = n171 & n1255 ;
  assign n3041 = n160 & n1214 ;
  assign n3043 = n3042 ^ n3041 ;
  assign n3044 = n3040 & n3043 ;
  assign n3045 = n3044 ^ n3040 ;
  assign n3046 = n3045 ^ n3043 ;
  assign n3047 = n314 & n3046 ;
  assign n3028 = n148 & n1316 ;
  assign n3027 = n137 & n1326 ;
  assign n3029 = n3028 ^ n3027 ;
  assign n3031 = n171 & n1204 ;
  assign n3030 = n160 & n1330 ;
  assign n3032 = n3031 ^ n3030 ;
  assign n3033 = n3029 & n3032 ;
  assign n3034 = n3033 ^ n3029 ;
  assign n3035 = n3034 ^ n3032 ;
  assign n3036 = n236 & ~n3035 ;
  assign n3037 = n3036 ^ n236 ;
  assign n3048 = n3047 ^ n3037 ;
  assign n3063 = n148 & n1250 ;
  assign n3060 = n137 & n1266 ;
  assign n3061 = n3060 ^ n137 ;
  assign n3062 = n3061 ^ n137 ;
  assign n3064 = n3063 ^ n3062 ;
  assign n3068 = n171 & n1229 ;
  assign n3065 = n160 & n1277 ;
  assign n3066 = n3065 ^ n160 ;
  assign n3067 = n3066 ^ n160 ;
  assign n3069 = n3068 ^ n3067 ;
  assign n3070 = n3064 & n3069 ;
  assign n3071 = n3070 ^ n3064 ;
  assign n3072 = n3071 ^ n3069 ;
  assign n3073 = n136 & n3072 ;
  assign n3050 = n148 & n1225 ;
  assign n3049 = n137 & n1235 ;
  assign n3051 = n3050 ^ n3049 ;
  assign n3053 = n171 & n1178 ;
  assign n3052 = n160 & n1239 ;
  assign n3054 = n3053 ^ n3052 ;
  assign n3055 = n3051 & n3054 ;
  assign n3056 = n3055 ^ n3051 ;
  assign n3057 = n3056 ^ n3054 ;
  assign n3058 = n188 & ~n3057 ;
  assign n3059 = n3058 ^ n188 ;
  assign n3074 = n3073 ^ n3059 ;
  assign n3075 = n3048 & n3074 ;
  assign n3076 = n3075 ^ n3048 ;
  assign n3077 = n3076 ^ n3074 ;
  assign n3125 = n3124 ^ n3077 ;
  assign n3126 = x134 & n3125 ;
  assign n3127 = n3126 ^ n3125 ;
  assign n3128 = n3127 ^ n3077 ;
  assign n3210 = n148 & n1636 ;
  assign n3207 = n137 & n1661 ;
  assign n3208 = n3207 ^ n137 ;
  assign n3209 = n3208 ^ n137 ;
  assign n3211 = n3210 ^ n3209 ;
  assign n3215 = n171 & n1760 ;
  assign n3212 = n160 & n1673 ;
  assign n3213 = n3212 ^ n160 ;
  assign n3214 = n3213 ^ n160 ;
  assign n3216 = n3215 ^ n3214 ;
  assign n3217 = n3211 & n3216 ;
  assign n3218 = n3217 ^ n3211 ;
  assign n3219 = n3218 ^ n3216 ;
  assign n3220 = n188 & n3219 ;
  assign n3195 = n148 & n1691 ;
  assign n3192 = n137 & n1718 ;
  assign n3193 = n3192 ^ n137 ;
  assign n3194 = n3193 ^ n137 ;
  assign n3196 = n3195 ^ n3194 ;
  assign n3200 = n171 & n1648 ;
  assign n3197 = n160 & n1730 ;
  assign n3198 = n3197 ^ n160 ;
  assign n3199 = n3198 ^ n160 ;
  assign n3201 = n3200 ^ n3199 ;
  assign n3202 = n3196 & n3201 ;
  assign n3203 = n3202 ^ n3196 ;
  assign n3204 = n3203 ^ n3201 ;
  assign n3205 = n136 & ~n3204 ;
  assign n3206 = n3205 ^ n136 ;
  assign n3221 = n3220 ^ n3206 ;
  assign n3240 = n148 & n1578 ;
  assign n3237 = n137 & n1603 ;
  assign n3238 = n3237 ^ n137 ;
  assign n3239 = n3238 ^ n137 ;
  assign n3241 = n3240 ^ n3239 ;
  assign n3245 = n171 & n1815 ;
  assign n3242 = n160 & n1615 ;
  assign n3243 = n3242 ^ n160 ;
  assign n3244 = n3243 ^ n160 ;
  assign n3246 = n3245 ^ n3244 ;
  assign n3247 = n3241 & n3246 ;
  assign n3248 = n3247 ^ n3241 ;
  assign n3249 = n3248 ^ n3246 ;
  assign n3250 = n236 & n3249 ;
  assign n3225 = n148 & n1803 ;
  assign n3222 = n137 & n1828 ;
  assign n3223 = n3222 ^ n137 ;
  assign n3224 = n3223 ^ n137 ;
  assign n3226 = n3225 ^ n3224 ;
  assign n3230 = n171 & n1705 ;
  assign n3227 = n160 & n1840 ;
  assign n3228 = n3227 ^ n160 ;
  assign n3229 = n3228 ^ n160 ;
  assign n3231 = n3230 ^ n3229 ;
  assign n3232 = n3226 & n3231 ;
  assign n3233 = n3232 ^ n3226 ;
  assign n3234 = n3233 ^ n3231 ;
  assign n3235 = n314 & ~n3234 ;
  assign n3236 = n3235 ^ n314 ;
  assign n3251 = n3250 ^ n3236 ;
  assign n3252 = n3221 & n3251 ;
  assign n3253 = n3252 ^ n3221 ;
  assign n3254 = n3253 ^ n3251 ;
  assign n3147 = n148 & n1464 ;
  assign n3144 = n137 & n1491 ;
  assign n3145 = n3144 ^ n137 ;
  assign n3146 = n3145 ^ n137 ;
  assign n3148 = n3147 ^ n3146 ;
  assign n3152 = n171 & n1415 ;
  assign n3149 = n160 & n1503 ;
  assign n3150 = n3149 ^ n160 ;
  assign n3151 = n3150 ^ n160 ;
  assign n3153 = n3152 ^ n3151 ;
  assign n3154 = n3148 & n3153 ;
  assign n3155 = n3154 ^ n3148 ;
  assign n3156 = n3155 ^ n3153 ;
  assign n3157 = n314 & n3156 ;
  assign n3132 = n148 & n1748 ;
  assign n3129 = n137 & n1773 ;
  assign n3130 = n3129 ^ n137 ;
  assign n3131 = n3130 ^ n137 ;
  assign n3133 = n3132 ^ n3131 ;
  assign n3137 = n171 & n1478 ;
  assign n3134 = n160 & n1785 ;
  assign n3135 = n3134 ^ n160 ;
  assign n3136 = n3135 ^ n160 ;
  assign n3138 = n3137 ^ n3136 ;
  assign n3139 = n3133 & n3138 ;
  assign n3140 = n3139 ^ n3133 ;
  assign n3141 = n3140 ^ n3138 ;
  assign n3142 = n236 & ~n3141 ;
  assign n3143 = n3142 ^ n236 ;
  assign n3158 = n3157 ^ n3143 ;
  assign n3175 = n137 & n1433 ;
  assign n3176 = n3175 ^ n137 ;
  assign n3177 = n3176 ^ n137 ;
  assign n3174 = n148 & n1402 ;
  assign n3178 = n3177 ^ n3174 ;
  assign n3182 = n171 & n1535 ;
  assign n3179 = n160 & n1446 ;
  assign n3180 = n3179 ^ n160 ;
  assign n3181 = n3180 ^ n160 ;
  assign n3183 = n3182 ^ n3181 ;
  assign n3184 = n3178 & n3183 ;
  assign n3185 = n3184 ^ n3178 ;
  assign n3186 = n3185 ^ n3183 ;
  assign n3187 = n136 & n3186 ;
  assign n3162 = n148 & n1521 ;
  assign n3159 = n137 & n1548 ;
  assign n3160 = n3159 ^ n137 ;
  assign n3161 = n3160 ^ n137 ;
  assign n3163 = n3162 ^ n3161 ;
  assign n3167 = n171 & n1590 ;
  assign n3164 = n160 & n1560 ;
  assign n3165 = n3164 ^ n160 ;
  assign n3166 = n3165 ^ n160 ;
  assign n3168 = n3167 ^ n3166 ;
  assign n3169 = n3163 & n3168 ;
  assign n3170 = n3169 ^ n3163 ;
  assign n3171 = n3170 ^ n3168 ;
  assign n3172 = n188 & ~n3171 ;
  assign n3173 = n3172 ^ n188 ;
  assign n3188 = n3187 ^ n3173 ;
  assign n3189 = n3158 & n3188 ;
  assign n3190 = n3189 ^ n3158 ;
  assign n3191 = n3190 ^ n3188 ;
  assign n3255 = n3254 ^ n3191 ;
  assign n3256 = x134 & n3255 ;
  assign n3257 = n3256 ^ n3255 ;
  assign n3258 = n3257 ^ n3191 ;
  assign n3278 = n188 & n391 ;
  assign n3276 = n136 & ~n485 ;
  assign n3277 = n3276 ^ n136 ;
  assign n3279 = n3278 ^ n3277 ;
  assign n3282 = n233 & n236 ;
  assign n3280 = n314 & ~n533 ;
  assign n3281 = n3280 ^ n314 ;
  assign n3283 = n3282 ^ n3281 ;
  assign n3284 = n3279 & n3283 ;
  assign n3285 = n3284 ^ n3279 ;
  assign n3286 = n3285 ^ n3283 ;
  assign n3261 = n236 & n438 ;
  assign n3259 = ~n185 & n188 ;
  assign n3260 = n3259 ^ n188 ;
  assign n3262 = n3261 ^ n3260 ;
  assign n3263 = ~n281 & n314 ;
  assign n3264 = n3263 ^ n314 ;
  assign n3265 = n136 & n335 ;
  assign n3266 = n3265 ^ n136 ;
  assign n3267 = n313 & n3266 ;
  assign n3268 = n3267 ^ n3266 ;
  assign n3269 = n3268 ^ n136 ;
  assign n3270 = n3264 & n3269 ;
  assign n3271 = n3270 ^ n3264 ;
  assign n3272 = n3271 ^ n3269 ;
  assign n3273 = n3262 & n3272 ;
  assign n3274 = n3273 ^ n3262 ;
  assign n3275 = n3274 ^ n3272 ;
  assign n3287 = n3286 ^ n3275 ;
  assign n3288 = x134 & n3287 ;
  assign n3289 = n3288 ^ n3287 ;
  assign n3290 = n3289 ^ n3275 ;
  assign n3304 = n188 & n924 ;
  assign n3302 = n136 & ~n1082 ;
  assign n3303 = n3302 ^ n136 ;
  assign n3305 = n3304 ^ n3303 ;
  assign n3308 = n236 & n619 ;
  assign n3306 = n314 & ~n1161 ;
  assign n3307 = n3306 ^ n314 ;
  assign n3309 = n3308 ^ n3307 ;
  assign n3310 = n3305 & n3309 ;
  assign n3311 = n3310 ^ n3305 ;
  assign n3312 = n3311 ^ n3309 ;
  assign n3293 = n314 & n698 ;
  assign n3291 = n236 & ~n1003 ;
  assign n3292 = n3291 ^ n236 ;
  assign n3294 = n3293 ^ n3292 ;
  assign n3297 = n136 & n842 ;
  assign n3295 = n188 & ~n777 ;
  assign n3296 = n3295 ^ n188 ;
  assign n3298 = n3297 ^ n3296 ;
  assign n3299 = n3294 & n3298 ;
  assign n3300 = n3299 ^ n3294 ;
  assign n3301 = n3300 ^ n3298 ;
  assign n3313 = n3312 ^ n3301 ;
  assign n3314 = x134 & n3313 ;
  assign n3315 = n3314 ^ n3313 ;
  assign n3316 = n3315 ^ n3301 ;
  assign n3330 = n188 & n1310 ;
  assign n3328 = n136 & ~n1361 ;
  assign n3329 = n3328 ^ n136 ;
  assign n3331 = n3330 ^ n3329 ;
  assign n3334 = n236 & n1193 ;
  assign n3332 = n314 & ~n1386 ;
  assign n3333 = n3332 ^ n314 ;
  assign n3335 = n3334 ^ n3333 ;
  assign n3336 = n3331 & n3335 ;
  assign n3337 = n3336 ^ n3331 ;
  assign n3338 = n3337 ^ n3335 ;
  assign n3319 = n314 & n1219 ;
  assign n3317 = n236 & ~n1335 ;
  assign n3318 = n3317 ^ n236 ;
  assign n3320 = n3319 ^ n3318 ;
  assign n3323 = n136 & n1282 ;
  assign n3321 = n188 & ~n1244 ;
  assign n3322 = n3321 ^ n188 ;
  assign n3324 = n3323 ^ n3322 ;
  assign n3325 = n3320 & n3324 ;
  assign n3326 = n3325 ^ n3320 ;
  assign n3327 = n3326 ^ n3324 ;
  assign n3339 = n3338 ^ n3327 ;
  assign n3340 = x134 & n3339 ;
  assign n3341 = n3340 ^ n3339 ;
  assign n3342 = n3341 ^ n3327 ;
  assign n3356 = n136 & n1735 ;
  assign n3354 = n188 & ~n1678 ;
  assign n3355 = n3354 ^ n188 ;
  assign n3357 = n3356 ^ n3355 ;
  assign n3360 = n314 & n1845 ;
  assign n3358 = n236 & ~n1620 ;
  assign n3359 = n3358 ^ n236 ;
  assign n3361 = n3360 ^ n3359 ;
  assign n3362 = n3357 & n3361 ;
  assign n3363 = n3362 ^ n3357 ;
  assign n3364 = n3363 ^ n3361 ;
  assign n3345 = n314 & n1508 ;
  assign n3343 = n236 & ~n1790 ;
  assign n3344 = n3343 ^ n236 ;
  assign n3346 = n3345 ^ n3344 ;
  assign n3349 = n188 & n1565 ;
  assign n3347 = n136 & ~n1451 ;
  assign n3348 = n3347 ^ n136 ;
  assign n3350 = n3349 ^ n3348 ;
  assign n3351 = n3346 & n3350 ;
  assign n3352 = n3351 ^ n3346 ;
  assign n3353 = n3352 ^ n3350 ;
  assign n3365 = n3364 ^ n3353 ;
  assign n3366 = x134 & n3365 ;
  assign n3367 = n3366 ^ n3365 ;
  assign n3368 = n3367 ^ n3353 ;
  assign n3388 = n188 & n1913 ;
  assign n3386 = n136 & ~n1935 ;
  assign n3387 = n3386 ^ n136 ;
  assign n3389 = n3388 ^ n3387 ;
  assign n3392 = n236 & n1888 ;
  assign n3390 = n314 & ~n1946 ;
  assign n3391 = n3390 ^ n314 ;
  assign n3393 = n3392 ^ n3391 ;
  assign n3394 = n3389 & n3393 ;
  assign n3395 = n3394 ^ n3389 ;
  assign n3396 = n3395 ^ n3393 ;
  assign n3369 = n236 & ~n1924 ;
  assign n3370 = n3369 ^ n236 ;
  assign n3371 = n136 & n1860 ;
  assign n3372 = n3371 ^ n136 ;
  assign n3373 = n1857 & n3372 ;
  assign n3374 = n3373 ^ n3372 ;
  assign n3375 = n3374 ^ n136 ;
  assign n3376 = n3370 & n3375 ;
  assign n3377 = n3376 ^ n3370 ;
  assign n3378 = n3377 ^ n3375 ;
  assign n3381 = n188 & n1899 ;
  assign n3379 = n314 & ~n1874 ;
  assign n3380 = n3379 ^ n314 ;
  assign n3382 = n3381 ^ n3380 ;
  assign n3383 = n3378 & n3382 ;
  assign n3384 = n3383 ^ n3378 ;
  assign n3385 = n3384 ^ n3382 ;
  assign n3397 = n3396 ^ n3385 ;
  assign n3398 = x134 & n3397 ;
  assign n3399 = n3398 ^ n3397 ;
  assign n3400 = n3399 ^ n3385 ;
  assign n3424 = n188 & n2039 ;
  assign n3422 = n136 & ~n2069 ;
  assign n3423 = n3422 ^ n136 ;
  assign n3425 = n3424 ^ n3423 ;
  assign n3428 = n236 & n2006 ;
  assign n3426 = n314 & ~n2084 ;
  assign n3427 = n3426 ^ n314 ;
  assign n3429 = n3428 ^ n3427 ;
  assign n3430 = n3425 & n3429 ;
  assign n3431 = n3430 ^ n3425 ;
  assign n3432 = n3431 ^ n3429 ;
  assign n3401 = n236 & n2054 ;
  assign n3402 = n3401 ^ n236 ;
  assign n3403 = n3402 ^ n236 ;
  assign n3404 = n1960 ^ n136 ;
  assign n3405 = n136 & n3404 ;
  assign n3406 = n3405 ^ n3404 ;
  assign n3407 = n3406 ^ n136 ;
  assign n3408 = n3407 ^ n1965 ;
  assign n3409 = n1966 & n3408 ;
  assign n3410 = n3409 ^ n3406 ;
  assign n3411 = n3410 ^ n1965 ;
  assign n3412 = n3403 & n3411 ;
  assign n3413 = n3412 ^ n3403 ;
  assign n3414 = n3413 ^ n3411 ;
  assign n3417 = n188 & n2021 ;
  assign n3415 = n314 & ~n1987 ;
  assign n3416 = n3415 ^ n314 ;
  assign n3418 = n3417 ^ n3416 ;
  assign n3419 = n3414 & n3418 ;
  assign n3420 = n3419 ^ n3414 ;
  assign n3421 = n3420 ^ n3418 ;
  assign n3433 = n3432 ^ n3421 ;
  assign n3434 = x134 & n3433 ;
  assign n3435 = n3434 ^ n3433 ;
  assign n3436 = n3435 ^ n3421 ;
  assign n3450 = n188 & n2149 ;
  assign n3448 = n136 & ~n2171 ;
  assign n3449 = n3448 ^ n136 ;
  assign n3451 = n3450 ^ n3449 ;
  assign n3454 = n236 & n2124 ;
  assign n3452 = n314 & ~n2182 ;
  assign n3453 = n3452 ^ n314 ;
  assign n3455 = n3454 ^ n3453 ;
  assign n3456 = n3451 & n3455 ;
  assign n3457 = n3456 ^ n3451 ;
  assign n3458 = n3457 ^ n3455 ;
  assign n3439 = n236 & n2160 ;
  assign n3437 = n136 & ~n2113 ;
  assign n3438 = n3437 ^ n136 ;
  assign n3440 = n3439 ^ n3438 ;
  assign n3443 = n188 & n2135 ;
  assign n3441 = n314 & ~n2102 ;
  assign n3442 = n3441 ^ n314 ;
  assign n3444 = n3443 ^ n3442 ;
  assign n3445 = n3440 & n3444 ;
  assign n3446 = n3445 ^ n3440 ;
  assign n3447 = n3446 ^ n3444 ;
  assign n3459 = n3458 ^ n3447 ;
  assign n3460 = x134 & n3459 ;
  assign n3461 = n3460 ^ n3459 ;
  assign n3462 = n3461 ^ n3447 ;
  assign n3476 = n188 & n2266 ;
  assign n3474 = n236 & ~n2233 ;
  assign n3475 = n3474 ^ n236 ;
  assign n3477 = n3476 ^ n3475 ;
  assign n3480 = n314 & n2311 ;
  assign n3478 = n136 & ~n2296 ;
  assign n3479 = n3478 ^ n136 ;
  assign n3481 = n3480 ^ n3479 ;
  assign n3482 = n3477 & n3481 ;
  assign n3483 = n3482 ^ n3477 ;
  assign n3484 = n3483 ^ n3481 ;
  assign n3465 = n136 & n2218 ;
  assign n3463 = n314 & ~n2204 ;
  assign n3464 = n3463 ^ n314 ;
  assign n3466 = n3465 ^ n3464 ;
  assign n3469 = n188 & n2248 ;
  assign n3467 = n236 & ~n2281 ;
  assign n3468 = n3467 ^ n236 ;
  assign n3470 = n3469 ^ n3468 ;
  assign n3471 = n3466 & n3470 ;
  assign n3472 = n3471 ^ n3466 ;
  assign n3473 = n3472 ^ n3470 ;
  assign n3485 = n3484 ^ n3473 ;
  assign n3486 = x134 & n3485 ;
  assign n3487 = n3486 ^ n3485 ;
  assign n3488 = n3487 ^ n3473 ;
  assign n3511 = n188 & n2383 ;
  assign n3509 = n236 & ~n2366 ;
  assign n3510 = n3509 ^ n236 ;
  assign n3512 = n3511 ^ n3510 ;
  assign n3515 = n314 & n2416 ;
  assign n3513 = n136 & ~n2405 ;
  assign n3514 = n3513 ^ n136 ;
  assign n3516 = n3515 ^ n3514 ;
  assign n3517 = n3512 & n3516 ;
  assign n3518 = n3517 ^ n3512 ;
  assign n3519 = n3518 ^ n3516 ;
  assign n3491 = n136 & n2340 ;
  assign n3489 = n314 & ~n2329 ;
  assign n3490 = n3489 ^ n314 ;
  assign n3492 = n3491 ^ n3490 ;
  assign n3493 = n2345 ^ n188 ;
  assign n3494 = n188 & n3493 ;
  assign n3495 = n3494 ^ n3493 ;
  assign n3496 = n3495 ^ n188 ;
  assign n3497 = n3496 ^ n2348 ;
  assign n3498 = n2349 & n3497 ;
  assign n3499 = n3498 ^ n3495 ;
  assign n3500 = n3499 ^ n2348 ;
  assign n3501 = n236 & ~n2394 ;
  assign n3502 = n3501 ^ n236 ;
  assign n3503 = n3500 & n3502 ;
  assign n3504 = n3503 ^ n3500 ;
  assign n3505 = n3504 ^ n3502 ;
  assign n3506 = n3492 & n3505 ;
  assign n3507 = n3506 ^ n3492 ;
  assign n3508 = n3507 ^ n3505 ;
  assign n3520 = n3519 ^ n3508 ;
  assign n3521 = x134 & n3520 ;
  assign n3522 = n3521 ^ n3520 ;
  assign n3523 = n3522 ^ n3508 ;
  assign n3537 = n188 & n2501 ;
  assign n3535 = n236 & ~n2468 ;
  assign n3536 = n3535 ^ n236 ;
  assign n3538 = n3537 ^ n3536 ;
  assign n3541 = n314 & n2546 ;
  assign n3539 = n136 & ~n2531 ;
  assign n3540 = n3539 ^ n136 ;
  assign n3542 = n3541 ^ n3540 ;
  assign n3543 = n3538 & n3542 ;
  assign n3544 = n3543 ^ n3538 ;
  assign n3545 = n3544 ^ n3542 ;
  assign n3526 = n136 & n2453 ;
  assign n3524 = n314 & ~n2438 ;
  assign n3525 = n3524 ^ n314 ;
  assign n3527 = n3526 ^ n3525 ;
  assign n3530 = n188 & n2483 ;
  assign n3528 = n236 & ~n2516 ;
  assign n3529 = n3528 ^ n236 ;
  assign n3531 = n3530 ^ n3529 ;
  assign n3532 = n3527 & n3531 ;
  assign n3533 = n3532 ^ n3527 ;
  assign n3534 = n3533 ^ n3531 ;
  assign n3546 = n3545 ^ n3534 ;
  assign n3547 = x134 & n3546 ;
  assign n3548 = n3547 ^ n3546 ;
  assign n3549 = n3548 ^ n3534 ;
  assign n3563 = n188 & n2613 ;
  assign n3561 = n136 & ~n2635 ;
  assign n3562 = n3561 ^ n136 ;
  assign n3564 = n3563 ^ n3562 ;
  assign n3567 = n236 & n2586 ;
  assign n3565 = n314 & ~n2646 ;
  assign n3566 = n3565 ^ n314 ;
  assign n3568 = n3567 ^ n3566 ;
  assign n3569 = n3564 & n3568 ;
  assign n3570 = n3569 ^ n3564 ;
  assign n3571 = n3570 ^ n3568 ;
  assign n3552 = n136 & n2575 ;
  assign n3550 = n314 & ~n2564 ;
  assign n3551 = n3550 ^ n314 ;
  assign n3553 = n3552 ^ n3551 ;
  assign n3556 = n188 & n2599 ;
  assign n3554 = n236 & ~n2624 ;
  assign n3555 = n3554 ^ n236 ;
  assign n3557 = n3556 ^ n3555 ;
  assign n3558 = n3553 & n3557 ;
  assign n3559 = n3558 ^ n3553 ;
  assign n3560 = n3559 ^ n3557 ;
  assign n3572 = n3571 ^ n3560 ;
  assign n3573 = x134 & n3572 ;
  assign n3574 = n3573 ^ n3572 ;
  assign n3575 = n3574 ^ n3560 ;
  assign n3589 = n188 & n2731 ;
  assign n3587 = n136 & ~n2761 ;
  assign n3588 = n3587 ^ n136 ;
  assign n3590 = n3589 ^ n3588 ;
  assign n3593 = n236 & n2698 ;
  assign n3591 = n314 & ~n2776 ;
  assign n3592 = n3591 ^ n314 ;
  assign n3594 = n3593 ^ n3592 ;
  assign n3595 = n3590 & n3594 ;
  assign n3596 = n3595 ^ n3590 ;
  assign n3597 = n3596 ^ n3594 ;
  assign n3578 = n136 & n2683 ;
  assign n3576 = n314 & ~n2668 ;
  assign n3577 = n3576 ^ n314 ;
  assign n3579 = n3578 ^ n3577 ;
  assign n3582 = n188 & n2713 ;
  assign n3580 = n236 & ~n2746 ;
  assign n3581 = n3580 ^ n236 ;
  assign n3583 = n3582 ^ n3581 ;
  assign n3584 = n3579 & n3583 ;
  assign n3585 = n3584 ^ n3579 ;
  assign n3586 = n3585 ^ n3583 ;
  assign n3598 = n3597 ^ n3586 ;
  assign n3599 = x134 & n3598 ;
  assign n3600 = n3599 ^ n3598 ;
  assign n3601 = n3600 ^ n3586 ;
  assign n3624 = n188 & n2850 ;
  assign n3622 = n136 & ~n2872 ;
  assign n3623 = n3622 ^ n136 ;
  assign n3625 = n3624 ^ n3623 ;
  assign n3628 = n236 & n2833 ;
  assign n3626 = n314 & ~n2883 ;
  assign n3627 = n3626 ^ n314 ;
  assign n3629 = n3628 ^ n3627 ;
  assign n3630 = n3625 & n3629 ;
  assign n3631 = n3630 ^ n3625 ;
  assign n3632 = n3631 ^ n3629 ;
  assign n3604 = n136 & n2805 ;
  assign n3602 = n314 & ~n2794 ;
  assign n3603 = n3602 ^ n314 ;
  assign n3605 = n3604 ^ n3603 ;
  assign n3606 = n2810 ^ n188 ;
  assign n3607 = n188 & n3606 ;
  assign n3608 = n3607 ^ n3606 ;
  assign n3609 = n3608 ^ n188 ;
  assign n3610 = n3609 ^ n2815 ;
  assign n3611 = n2816 & n3610 ;
  assign n3612 = n3611 ^ n3608 ;
  assign n3613 = n3612 ^ n2815 ;
  assign n3614 = n236 & ~n2861 ;
  assign n3615 = n3614 ^ n236 ;
  assign n3616 = n3613 & n3615 ;
  assign n3617 = n3616 ^ n3613 ;
  assign n3618 = n3617 ^ n3615 ;
  assign n3619 = n3605 & n3618 ;
  assign n3620 = n3619 ^ n3605 ;
  assign n3621 = n3620 ^ n3618 ;
  assign n3633 = n3632 ^ n3621 ;
  assign n3634 = x134 & n3633 ;
  assign n3635 = n3634 ^ n3633 ;
  assign n3636 = n3635 ^ n3621 ;
  assign n3657 = n188 & n2972 ;
  assign n3655 = n136 & ~n3002 ;
  assign n3656 = n3655 ^ n136 ;
  assign n3658 = n3657 ^ n3656 ;
  assign n3661 = n236 & n2950 ;
  assign n3659 = n314 & ~n3017 ;
  assign n3660 = n3659 ^ n314 ;
  assign n3662 = n3661 ^ n3660 ;
  assign n3663 = n3658 & n3662 ;
  assign n3664 = n3663 ^ n3658 ;
  assign n3665 = n3664 ^ n3662 ;
  assign n3639 = n136 & n2920 ;
  assign n3637 = n314 & ~n2905 ;
  assign n3638 = n3637 ^ n314 ;
  assign n3640 = n3639 ^ n3638 ;
  assign n3641 = n188 & n2932 ;
  assign n3642 = n3641 ^ n188 ;
  assign n3643 = n2927 & n3642 ;
  assign n3644 = n3643 ^ n3642 ;
  assign n3645 = n3644 ^ n188 ;
  assign n3646 = n236 & n2987 ;
  assign n3647 = n3646 ^ n236 ;
  assign n3648 = n3647 ^ n236 ;
  assign n3649 = n3645 & n3648 ;
  assign n3650 = n3649 ^ n3645 ;
  assign n3651 = n3650 ^ n3648 ;
  assign n3652 = n3640 & n3651 ;
  assign n3653 = n3652 ^ n3640 ;
  assign n3654 = n3653 ^ n3651 ;
  assign n3666 = n3665 ^ n3654 ;
  assign n3667 = x134 & n3666 ;
  assign n3668 = n3667 ^ n3666 ;
  assign n3669 = n3668 ^ n3654 ;
  assign n3683 = n188 & n3086 ;
  assign n3681 = n136 & ~n3108 ;
  assign n3682 = n3681 ^ n136 ;
  assign n3684 = n3683 ^ n3682 ;
  assign n3687 = n236 & n3057 ;
  assign n3685 = n314 & ~n3119 ;
  assign n3686 = n3685 ^ n314 ;
  assign n3688 = n3687 ^ n3686 ;
  assign n3689 = n3684 & n3688 ;
  assign n3690 = n3689 ^ n3684 ;
  assign n3691 = n3690 ^ n3688 ;
  assign n3672 = n136 & n3046 ;
  assign n3670 = n314 & ~n3035 ;
  assign n3671 = n3670 ^ n314 ;
  assign n3673 = n3672 ^ n3671 ;
  assign n3676 = n188 & n3072 ;
  assign n3674 = n236 & ~n3097 ;
  assign n3675 = n3674 ^ n236 ;
  assign n3677 = n3676 ^ n3675 ;
  assign n3678 = n3673 & n3677 ;
  assign n3679 = n3678 ^ n3673 ;
  assign n3680 = n3679 ^ n3677 ;
  assign n3692 = n3691 ^ n3680 ;
  assign n3693 = x134 & n3692 ;
  assign n3694 = n3693 ^ n3692 ;
  assign n3695 = n3694 ^ n3680 ;
  assign n3709 = n188 & n3204 ;
  assign n3707 = n136 & ~n3234 ;
  assign n3708 = n3707 ^ n136 ;
  assign n3710 = n3709 ^ n3708 ;
  assign n3713 = n236 & n3171 ;
  assign n3711 = n314 & ~n3249 ;
  assign n3712 = n3711 ^ n314 ;
  assign n3714 = n3713 ^ n3712 ;
  assign n3715 = n3710 & n3714 ;
  assign n3716 = n3715 ^ n3710 ;
  assign n3717 = n3716 ^ n3714 ;
  assign n3698 = n136 & n3156 ;
  assign n3696 = n314 & ~n3141 ;
  assign n3697 = n3696 ^ n314 ;
  assign n3699 = n3698 ^ n3697 ;
  assign n3702 = n188 & n3186 ;
  assign n3700 = n236 & ~n3219 ;
  assign n3701 = n3700 ^ n236 ;
  assign n3703 = n3702 ^ n3701 ;
  assign n3704 = n3699 & n3703 ;
  assign n3705 = n3704 ^ n3699 ;
  assign n3706 = n3705 ^ n3703 ;
  assign n3718 = n3717 ^ n3706 ;
  assign n3719 = x134 & n3718 ;
  assign n3720 = n3719 ^ n3718 ;
  assign n3721 = n3720 ^ n3706 ;
  assign n3741 = n188 & n485 ;
  assign n3739 = n136 & ~n533 ;
  assign n3740 = n3739 ^ n136 ;
  assign n3742 = n3741 ^ n3740 ;
  assign n3745 = n185 & n236 ;
  assign n3743 = ~n233 & n314 ;
  assign n3744 = n3743 ^ n314 ;
  assign n3746 = n3745 ^ n3744 ;
  assign n3747 = n3742 & n3746 ;
  assign n3748 = n3747 ^ n3742 ;
  assign n3749 = n3748 ^ n3746 ;
  assign n3724 = n314 & n438 ;
  assign n3722 = n236 & ~n391 ;
  assign n3723 = n3722 ^ n236 ;
  assign n3725 = n3724 ^ n3723 ;
  assign n3726 = n136 & ~n281 ;
  assign n3727 = n3726 ^ n136 ;
  assign n3728 = n188 & n335 ;
  assign n3729 = n3728 ^ n188 ;
  assign n3730 = n313 & n3729 ;
  assign n3731 = n3730 ^ n3729 ;
  assign n3732 = n3731 ^ n188 ;
  assign n3733 = n3727 & n3732 ;
  assign n3734 = n3733 ^ n3727 ;
  assign n3735 = n3734 ^ n3732 ;
  assign n3736 = n3725 & n3735 ;
  assign n3737 = n3736 ^ n3725 ;
  assign n3738 = n3737 ^ n3735 ;
  assign n3750 = n3749 ^ n3738 ;
  assign n3751 = x134 & n3750 ;
  assign n3752 = n3751 ^ n3750 ;
  assign n3753 = n3752 ^ n3738 ;
  assign n3767 = n188 & n1082 ;
  assign n3765 = n136 & ~n1161 ;
  assign n3766 = n3765 ^ n136 ;
  assign n3768 = n3767 ^ n3766 ;
  assign n3771 = n236 & n777 ;
  assign n3769 = n314 & ~n619 ;
  assign n3770 = n3769 ^ n314 ;
  assign n3772 = n3771 ^ n3770 ;
  assign n3773 = n3768 & n3772 ;
  assign n3774 = n3773 ^ n3768 ;
  assign n3775 = n3774 ^ n3772 ;
  assign n3756 = n136 & n698 ;
  assign n3754 = n314 & ~n1003 ;
  assign n3755 = n3754 ^ n314 ;
  assign n3757 = n3756 ^ n3755 ;
  assign n3760 = n188 & n842 ;
  assign n3758 = n236 & ~n924 ;
  assign n3759 = n3758 ^ n236 ;
  assign n3761 = n3760 ^ n3759 ;
  assign n3762 = n3757 & n3761 ;
  assign n3763 = n3762 ^ n3757 ;
  assign n3764 = n3763 ^ n3761 ;
  assign n3776 = n3775 ^ n3764 ;
  assign n3777 = x134 & n3776 ;
  assign n3778 = n3777 ^ n3776 ;
  assign n3779 = n3778 ^ n3764 ;
  assign n3793 = n188 & n1361 ;
  assign n3791 = n136 & ~n1386 ;
  assign n3792 = n3791 ^ n136 ;
  assign n3794 = n3793 ^ n3792 ;
  assign n3797 = n236 & n1244 ;
  assign n3795 = n314 & ~n1193 ;
  assign n3796 = n3795 ^ n314 ;
  assign n3798 = n3797 ^ n3796 ;
  assign n3799 = n3794 & n3798 ;
  assign n3800 = n3799 ^ n3794 ;
  assign n3801 = n3800 ^ n3798 ;
  assign n3782 = n136 & n1219 ;
  assign n3780 = n314 & ~n1335 ;
  assign n3781 = n3780 ^ n314 ;
  assign n3783 = n3782 ^ n3781 ;
  assign n3786 = n188 & n1282 ;
  assign n3784 = n236 & ~n1310 ;
  assign n3785 = n3784 ^ n236 ;
  assign n3787 = n3786 ^ n3785 ;
  assign n3788 = n3783 & n3787 ;
  assign n3789 = n3788 ^ n3783 ;
  assign n3790 = n3789 ^ n3787 ;
  assign n3802 = n3801 ^ n3790 ;
  assign n3803 = x134 & n3802 ;
  assign n3804 = n3803 ^ n3802 ;
  assign n3805 = n3804 ^ n3790 ;
  assign n3819 = n188 & n1735 ;
  assign n3817 = n236 & ~n1565 ;
  assign n3818 = n3817 ^ n236 ;
  assign n3820 = n3819 ^ n3818 ;
  assign n3823 = n136 & n1845 ;
  assign n3821 = n314 & ~n1620 ;
  assign n3822 = n3821 ^ n314 ;
  assign n3824 = n3823 ^ n3822 ;
  assign n3825 = n3820 & n3824 ;
  assign n3826 = n3825 ^ n3820 ;
  assign n3827 = n3826 ^ n3824 ;
  assign n3808 = n136 & n1508 ;
  assign n3806 = n236 & ~n1678 ;
  assign n3807 = n3806 ^ n236 ;
  assign n3809 = n3808 ^ n3807 ;
  assign n3812 = n188 & n1451 ;
  assign n3810 = n314 & ~n1790 ;
  assign n3811 = n3810 ^ n314 ;
  assign n3813 = n3812 ^ n3811 ;
  assign n3814 = n3809 & n3813 ;
  assign n3815 = n3814 ^ n3809 ;
  assign n3816 = n3815 ^ n3813 ;
  assign n3828 = n3827 ^ n3816 ;
  assign n3829 = x134 & n3828 ;
  assign n3830 = n3829 ^ n3828 ;
  assign n3831 = n3830 ^ n3816 ;
  assign n3851 = n188 & n1935 ;
  assign n3849 = n136 & ~n1946 ;
  assign n3850 = n3849 ^ n136 ;
  assign n3852 = n3851 ^ n3850 ;
  assign n3855 = n236 & n1899 ;
  assign n3853 = n314 & ~n1888 ;
  assign n3854 = n3853 ^ n314 ;
  assign n3856 = n3855 ^ n3854 ;
  assign n3857 = n3852 & n3856 ;
  assign n3858 = n3857 ^ n3852 ;
  assign n3859 = n3858 ^ n3856 ;
  assign n3834 = n314 & n1924 ;
  assign n3832 = n236 & ~n1913 ;
  assign n3833 = n3832 ^ n236 ;
  assign n3835 = n3834 ^ n3833 ;
  assign n3836 = n136 & ~n1874 ;
  assign n3837 = n3836 ^ n136 ;
  assign n3838 = n188 & n1860 ;
  assign n3839 = n3838 ^ n188 ;
  assign n3840 = n1857 & n3839 ;
  assign n3841 = n3840 ^ n3839 ;
  assign n3842 = n3841 ^ n188 ;
  assign n3843 = n3837 & n3842 ;
  assign n3844 = n3843 ^ n3837 ;
  assign n3845 = n3844 ^ n3842 ;
  assign n3846 = n3835 & n3845 ;
  assign n3847 = n3846 ^ n3835 ;
  assign n3848 = n3847 ^ n3845 ;
  assign n3860 = n3859 ^ n3848 ;
  assign n3861 = x134 & n3860 ;
  assign n3862 = n3861 ^ n3860 ;
  assign n3863 = n3862 ^ n3848 ;
  assign n3887 = n188 & n2069 ;
  assign n3885 = n136 & ~n2084 ;
  assign n3886 = n3885 ^ n136 ;
  assign n3888 = n3887 ^ n3886 ;
  assign n3891 = n236 & n2021 ;
  assign n3889 = n314 & ~n2006 ;
  assign n3890 = n3889 ^ n314 ;
  assign n3892 = n3891 ^ n3890 ;
  assign n3893 = n3888 & n3892 ;
  assign n3894 = n3893 ^ n3888 ;
  assign n3895 = n3894 ^ n3892 ;
  assign n3866 = n314 & n2054 ;
  assign n3864 = n236 & ~n2039 ;
  assign n3865 = n3864 ^ n236 ;
  assign n3867 = n3866 ^ n3865 ;
  assign n3868 = n136 & n1987 ;
  assign n3869 = n3868 ^ n136 ;
  assign n3870 = n3869 ^ n136 ;
  assign n3871 = n1960 ^ n188 ;
  assign n3872 = n188 & n3871 ;
  assign n3873 = n3872 ^ n3871 ;
  assign n3874 = n3873 ^ n188 ;
  assign n3875 = n3874 ^ n1965 ;
  assign n3876 = n1966 & n3875 ;
  assign n3877 = n3876 ^ n3873 ;
  assign n3878 = n3877 ^ n1965 ;
  assign n3879 = n3870 & n3878 ;
  assign n3880 = n3879 ^ n3870 ;
  assign n3881 = n3880 ^ n3878 ;
  assign n3882 = n3867 & n3881 ;
  assign n3883 = n3882 ^ n3867 ;
  assign n3884 = n3883 ^ n3881 ;
  assign n3896 = n3895 ^ n3884 ;
  assign n3897 = x134 & n3896 ;
  assign n3898 = n3897 ^ n3896 ;
  assign n3899 = n3898 ^ n3884 ;
  assign n3913 = n188 & n2171 ;
  assign n3911 = n136 & ~n2182 ;
  assign n3912 = n3911 ^ n136 ;
  assign n3914 = n3913 ^ n3912 ;
  assign n3917 = n236 & n2135 ;
  assign n3915 = n314 & ~n2124 ;
  assign n3916 = n3915 ^ n314 ;
  assign n3918 = n3917 ^ n3916 ;
  assign n3919 = n3914 & n3918 ;
  assign n3920 = n3919 ^ n3914 ;
  assign n3921 = n3920 ^ n3918 ;
  assign n3902 = n314 & n2160 ;
  assign n3900 = n236 & ~n2149 ;
  assign n3901 = n3900 ^ n236 ;
  assign n3903 = n3902 ^ n3901 ;
  assign n3906 = n136 & n2102 ;
  assign n3904 = n188 & ~n2113 ;
  assign n3905 = n3904 ^ n188 ;
  assign n3907 = n3906 ^ n3905 ;
  assign n3908 = n3903 & n3907 ;
  assign n3909 = n3908 ^ n3903 ;
  assign n3910 = n3909 ^ n3907 ;
  assign n3922 = n3921 ^ n3910 ;
  assign n3923 = x134 & n3922 ;
  assign n3924 = n3923 ^ n3922 ;
  assign n3925 = n3924 ^ n3910 ;
  assign n3939 = n314 & n2233 ;
  assign n3937 = n236 & ~n2248 ;
  assign n3938 = n3937 ^ n236 ;
  assign n3940 = n3939 ^ n3938 ;
  assign n3943 = n136 & n2311 ;
  assign n3941 = n188 & ~n2296 ;
  assign n3942 = n3941 ^ n188 ;
  assign n3944 = n3943 ^ n3942 ;
  assign n3945 = n3940 & n3944 ;
  assign n3946 = n3945 ^ n3940 ;
  assign n3947 = n3946 ^ n3944 ;
  assign n3928 = n188 & n2218 ;
  assign n3926 = n136 & ~n2204 ;
  assign n3927 = n3926 ^ n136 ;
  assign n3929 = n3928 ^ n3927 ;
  assign n3932 = n236 & n2266 ;
  assign n3930 = n314 & ~n2281 ;
  assign n3931 = n3930 ^ n314 ;
  assign n3933 = n3932 ^ n3931 ;
  assign n3934 = n3929 & n3933 ;
  assign n3935 = n3934 ^ n3929 ;
  assign n3936 = n3935 ^ n3933 ;
  assign n3948 = n3947 ^ n3936 ;
  assign n3949 = x134 & n3948 ;
  assign n3950 = n3949 ^ n3948 ;
  assign n3951 = n3950 ^ n3936 ;
  assign n3963 = n314 & ~n2366 ;
  assign n3964 = n3963 ^ n314 ;
  assign n3965 = n2345 ^ n236 ;
  assign n3966 = n236 & n3965 ;
  assign n3967 = n3966 ^ n3965 ;
  assign n3968 = n3967 ^ n236 ;
  assign n3969 = n3968 ^ n2348 ;
  assign n3970 = n2349 & n3969 ;
  assign n3971 = n3970 ^ n3967 ;
  assign n3972 = n3971 ^ n2348 ;
  assign n3973 = n3964 & n3972 ;
  assign n3974 = n3973 ^ n3964 ;
  assign n3975 = n3974 ^ n3972 ;
  assign n3978 = n136 & n2416 ;
  assign n3976 = n188 & ~n2405 ;
  assign n3977 = n3976 ^ n188 ;
  assign n3979 = n3978 ^ n3977 ;
  assign n3980 = n3975 & n3979 ;
  assign n3981 = n3980 ^ n3975 ;
  assign n3982 = n3981 ^ n3979 ;
  assign n3954 = n188 & n2340 ;
  assign n3952 = n136 & ~n2329 ;
  assign n3953 = n3952 ^ n136 ;
  assign n3955 = n3954 ^ n3953 ;
  assign n3958 = n236 & n2383 ;
  assign n3956 = n314 & ~n2394 ;
  assign n3957 = n3956 ^ n314 ;
  assign n3959 = n3958 ^ n3957 ;
  assign n3960 = n3955 & n3959 ;
  assign n3961 = n3960 ^ n3955 ;
  assign n3962 = n3961 ^ n3959 ;
  assign n3983 = n3982 ^ n3962 ;
  assign n3984 = x134 & n3983 ;
  assign n3985 = n3984 ^ n3983 ;
  assign n3986 = n3985 ^ n3962 ;
  assign n4000 = n314 & n2468 ;
  assign n3998 = n236 & ~n2483 ;
  assign n3999 = n3998 ^ n236 ;
  assign n4001 = n4000 ^ n3999 ;
  assign n4004 = n136 & n2546 ;
  assign n4002 = n188 & ~n2531 ;
  assign n4003 = n4002 ^ n188 ;
  assign n4005 = n4004 ^ n4003 ;
  assign n4006 = n4001 & n4005 ;
  assign n4007 = n4006 ^ n4001 ;
  assign n4008 = n4007 ^ n4005 ;
  assign n3989 = n188 & n2453 ;
  assign n3987 = n136 & ~n2438 ;
  assign n3988 = n3987 ^ n136 ;
  assign n3990 = n3989 ^ n3988 ;
  assign n3993 = n236 & n2501 ;
  assign n3991 = n314 & ~n2516 ;
  assign n3992 = n3991 ^ n314 ;
  assign n3994 = n3993 ^ n3992 ;
  assign n3995 = n3990 & n3994 ;
  assign n3996 = n3995 ^ n3990 ;
  assign n3997 = n3996 ^ n3994 ;
  assign n4009 = n4008 ^ n3997 ;
  assign n4010 = x134 & n4009 ;
  assign n4011 = n4010 ^ n4009 ;
  assign n4012 = n4011 ^ n3997 ;
  assign n4026 = n188 & n2635 ;
  assign n4024 = n136 & ~n2646 ;
  assign n4025 = n4024 ^ n136 ;
  assign n4027 = n4026 ^ n4025 ;
  assign n4030 = n236 & n2599 ;
  assign n4028 = n314 & ~n2586 ;
  assign n4029 = n4028 ^ n314 ;
  assign n4031 = n4030 ^ n4029 ;
  assign n4032 = n4027 & n4031 ;
  assign n4033 = n4032 ^ n4027 ;
  assign n4034 = n4033 ^ n4031 ;
  assign n4015 = n188 & n2575 ;
  assign n4013 = n136 & ~n2564 ;
  assign n4014 = n4013 ^ n136 ;
  assign n4016 = n4015 ^ n4014 ;
  assign n4019 = n236 & n2613 ;
  assign n4017 = n314 & ~n2624 ;
  assign n4018 = n4017 ^ n314 ;
  assign n4020 = n4019 ^ n4018 ;
  assign n4021 = n4016 & n4020 ;
  assign n4022 = n4021 ^ n4016 ;
  assign n4023 = n4022 ^ n4020 ;
  assign n4035 = n4034 ^ n4023 ;
  assign n4036 = x134 & n4035 ;
  assign n4037 = n4036 ^ n4035 ;
  assign n4038 = n4037 ^ n4023 ;
  assign n4052 = n188 & n2761 ;
  assign n4050 = n136 & ~n2776 ;
  assign n4051 = n4050 ^ n136 ;
  assign n4053 = n4052 ^ n4051 ;
  assign n4056 = n236 & n2713 ;
  assign n4054 = n314 & ~n2698 ;
  assign n4055 = n4054 ^ n314 ;
  assign n4057 = n4056 ^ n4055 ;
  assign n4058 = n4053 & n4057 ;
  assign n4059 = n4058 ^ n4053 ;
  assign n4060 = n4059 ^ n4057 ;
  assign n4041 = n188 & n2683 ;
  assign n4039 = n136 & ~n2668 ;
  assign n4040 = n4039 ^ n136 ;
  assign n4042 = n4041 ^ n4040 ;
  assign n4045 = n236 & n2731 ;
  assign n4043 = n314 & ~n2746 ;
  assign n4044 = n4043 ^ n314 ;
  assign n4046 = n4045 ^ n4044 ;
  assign n4047 = n4042 & n4046 ;
  assign n4048 = n4047 ^ n4042 ;
  assign n4049 = n4048 ^ n4046 ;
  assign n4061 = n4060 ^ n4049 ;
  assign n4062 = x134 & n4061 ;
  assign n4063 = n4062 ^ n4061 ;
  assign n4064 = n4063 ^ n4049 ;
  assign n4078 = n188 & n2872 ;
  assign n4076 = n136 & ~n2883 ;
  assign n4077 = n4076 ^ n136 ;
  assign n4079 = n4078 ^ n4077 ;
  assign n4080 = n2810 ^ n236 ;
  assign n4081 = n236 & n4080 ;
  assign n4082 = n4081 ^ n4080 ;
  assign n4083 = n4082 ^ n236 ;
  assign n4084 = n4083 ^ n2815 ;
  assign n4085 = n2816 & n4084 ;
  assign n4086 = n4085 ^ n4082 ;
  assign n4087 = n4086 ^ n2815 ;
  assign n4088 = n314 & ~n2833 ;
  assign n4089 = n4088 ^ n314 ;
  assign n4090 = n4087 & n4089 ;
  assign n4091 = n4090 ^ n4087 ;
  assign n4092 = n4091 ^ n4089 ;
  assign n4093 = n4079 & n4092 ;
  assign n4094 = n4093 ^ n4079 ;
  assign n4095 = n4094 ^ n4092 ;
  assign n4067 = n188 & n2805 ;
  assign n4065 = n136 & ~n2794 ;
  assign n4066 = n4065 ^ n136 ;
  assign n4068 = n4067 ^ n4066 ;
  assign n4071 = n236 & n2850 ;
  assign n4069 = n314 & ~n2861 ;
  assign n4070 = n4069 ^ n314 ;
  assign n4072 = n4071 ^ n4070 ;
  assign n4073 = n4068 & n4072 ;
  assign n4074 = n4073 ^ n4068 ;
  assign n4075 = n4074 ^ n4072 ;
  assign n4096 = n4095 ^ n4075 ;
  assign n4097 = x134 & n4096 ;
  assign n4098 = n4097 ^ n4096 ;
  assign n4099 = n4098 ^ n4075 ;
  assign n4113 = n188 & n3002 ;
  assign n4111 = n136 & ~n3017 ;
  assign n4112 = n4111 ^ n136 ;
  assign n4114 = n4113 ^ n4112 ;
  assign n4115 = n236 & n2932 ;
  assign n4116 = n4115 ^ n236 ;
  assign n4117 = n2927 & n4116 ;
  assign n4118 = n4117 ^ n4116 ;
  assign n4119 = n4118 ^ n236 ;
  assign n4120 = n314 & n2950 ;
  assign n4121 = n4120 ^ n314 ;
  assign n4122 = n4121 ^ n314 ;
  assign n4123 = n4119 & n4122 ;
  assign n4124 = n4123 ^ n4119 ;
  assign n4125 = n4124 ^ n4122 ;
  assign n4126 = n4114 & n4125 ;
  assign n4127 = n4126 ^ n4114 ;
  assign n4128 = n4127 ^ n4125 ;
  assign n4102 = n188 & n2920 ;
  assign n4100 = n136 & ~n2905 ;
  assign n4101 = n4100 ^ n136 ;
  assign n4103 = n4102 ^ n4101 ;
  assign n4106 = n236 & n2972 ;
  assign n4104 = n314 & ~n2987 ;
  assign n4105 = n4104 ^ n314 ;
  assign n4107 = n4106 ^ n4105 ;
  assign n4108 = n4103 & n4107 ;
  assign n4109 = n4108 ^ n4103 ;
  assign n4110 = n4109 ^ n4107 ;
  assign n4129 = n4128 ^ n4110 ;
  assign n4130 = x134 & n4129 ;
  assign n4131 = n4130 ^ n4129 ;
  assign n4132 = n4131 ^ n4110 ;
  assign n4146 = n188 & n3108 ;
  assign n4144 = n136 & ~n3119 ;
  assign n4145 = n4144 ^ n136 ;
  assign n4147 = n4146 ^ n4145 ;
  assign n4150 = n236 & n3072 ;
  assign n4148 = n314 & ~n3057 ;
  assign n4149 = n4148 ^ n314 ;
  assign n4151 = n4150 ^ n4149 ;
  assign n4152 = n4147 & n4151 ;
  assign n4153 = n4152 ^ n4147 ;
  assign n4154 = n4153 ^ n4151 ;
  assign n4135 = n188 & n3046 ;
  assign n4133 = n136 & ~n3035 ;
  assign n4134 = n4133 ^ n136 ;
  assign n4136 = n4135 ^ n4134 ;
  assign n4139 = n236 & n3086 ;
  assign n4137 = n314 & ~n3097 ;
  assign n4138 = n4137 ^ n314 ;
  assign n4140 = n4139 ^ n4138 ;
  assign n4141 = n4136 & n4140 ;
  assign n4142 = n4141 ^ n4136 ;
  assign n4143 = n4142 ^ n4140 ;
  assign n4155 = n4154 ^ n4143 ;
  assign n4156 = x134 & n4155 ;
  assign n4157 = n4156 ^ n4155 ;
  assign n4158 = n4157 ^ n4143 ;
  assign n4172 = n188 & n3234 ;
  assign n4170 = n136 & ~n3249 ;
  assign n4171 = n4170 ^ n136 ;
  assign n4173 = n4172 ^ n4171 ;
  assign n4176 = n236 & n3186 ;
  assign n4174 = n314 & ~n3171 ;
  assign n4175 = n4174 ^ n314 ;
  assign n4177 = n4176 ^ n4175 ;
  assign n4178 = n4173 & n4177 ;
  assign n4179 = n4178 ^ n4173 ;
  assign n4180 = n4179 ^ n4177 ;
  assign n4161 = n188 & n3156 ;
  assign n4159 = n136 & ~n3141 ;
  assign n4160 = n4159 ^ n136 ;
  assign n4162 = n4161 ^ n4160 ;
  assign n4165 = n236 & n3204 ;
  assign n4163 = n314 & ~n3219 ;
  assign n4164 = n4163 ^ n314 ;
  assign n4166 = n4165 ^ n4164 ;
  assign n4167 = n4162 & n4166 ;
  assign n4168 = n4167 ^ n4162 ;
  assign n4169 = n4168 ^ n4166 ;
  assign n4181 = n4180 ^ n4169 ;
  assign n4182 = x134 & n4181 ;
  assign n4183 = n4182 ^ n4181 ;
  assign n4184 = n4183 ^ n4169 ;
  assign n4198 = n188 & n533 ;
  assign n4196 = n136 & ~n233 ;
  assign n4197 = n4196 ^ n136 ;
  assign n4199 = n4198 ^ n4197 ;
  assign n4200 = n236 & n335 ;
  assign n4201 = n4200 ^ n236 ;
  assign n4202 = n313 & n4201 ;
  assign n4203 = n4202 ^ n4201 ;
  assign n4204 = n4203 ^ n236 ;
  assign n4205 = ~n185 & n314 ;
  assign n4206 = n4205 ^ n314 ;
  assign n4207 = n4204 & n4206 ;
  assign n4208 = n4207 ^ n4204 ;
  assign n4209 = n4208 ^ n4206 ;
  assign n4210 = n4199 & n4209 ;
  assign n4211 = n4210 ^ n4199 ;
  assign n4212 = n4211 ^ n4209 ;
  assign n4187 = n136 & n438 ;
  assign n4185 = n314 & ~n391 ;
  assign n4186 = n4185 ^ n314 ;
  assign n4188 = n4187 ^ n4186 ;
  assign n4191 = n188 & n281 ;
  assign n4189 = n236 & ~n485 ;
  assign n4190 = n4189 ^ n236 ;
  assign n4192 = n4191 ^ n4190 ;
  assign n4193 = n4188 & n4192 ;
  assign n4194 = n4193 ^ n4188 ;
  assign n4195 = n4194 ^ n4192 ;
  assign n4213 = n4212 ^ n4195 ;
  assign n4214 = x134 & n4213 ;
  assign n4215 = n4214 ^ n4213 ;
  assign n4216 = n4215 ^ n4195 ;
  assign n4230 = n188 & n1161 ;
  assign n4228 = n136 & ~n619 ;
  assign n4229 = n4228 ^ n136 ;
  assign n4231 = n4230 ^ n4229 ;
  assign n4234 = n236 & n842 ;
  assign n4232 = n314 & ~n777 ;
  assign n4233 = n4232 ^ n314 ;
  assign n4235 = n4234 ^ n4233 ;
  assign n4236 = n4231 & n4235 ;
  assign n4237 = n4236 ^ n4231 ;
  assign n4238 = n4237 ^ n4235 ;
  assign n4219 = n188 & n698 ;
  assign n4217 = n136 & ~n1003 ;
  assign n4218 = n4217 ^ n136 ;
  assign n4220 = n4219 ^ n4218 ;
  assign n4223 = n236 & n1082 ;
  assign n4221 = n314 & ~n924 ;
  assign n4222 = n4221 ^ n314 ;
  assign n4224 = n4223 ^ n4222 ;
  assign n4225 = n4220 & n4224 ;
  assign n4226 = n4225 ^ n4220 ;
  assign n4227 = n4226 ^ n4224 ;
  assign n4239 = n4238 ^ n4227 ;
  assign n4240 = x134 & n4239 ;
  assign n4241 = n4240 ^ n4239 ;
  assign n4242 = n4241 ^ n4227 ;
  assign n4256 = n188 & n1386 ;
  assign n4254 = n136 & ~n1193 ;
  assign n4255 = n4254 ^ n136 ;
  assign n4257 = n4256 ^ n4255 ;
  assign n4260 = n236 & n1282 ;
  assign n4258 = n314 & ~n1244 ;
  assign n4259 = n4258 ^ n314 ;
  assign n4261 = n4260 ^ n4259 ;
  assign n4262 = n4257 & n4261 ;
  assign n4263 = n4262 ^ n4257 ;
  assign n4264 = n4263 ^ n4261 ;
  assign n4245 = n188 & n1219 ;
  assign n4243 = n136 & ~n1335 ;
  assign n4244 = n4243 ^ n136 ;
  assign n4246 = n4245 ^ n4244 ;
  assign n4249 = n236 & n1361 ;
  assign n4247 = n314 & ~n1310 ;
  assign n4248 = n4247 ^ n314 ;
  assign n4250 = n4249 ^ n4248 ;
  assign n4251 = n4246 & n4250 ;
  assign n4252 = n4251 ^ n4246 ;
  assign n4253 = n4252 ^ n4250 ;
  assign n4265 = n4264 ^ n4253 ;
  assign n4266 = x134 & n4265 ;
  assign n4267 = n4266 ^ n4265 ;
  assign n4268 = n4267 ^ n4253 ;
  assign n4282 = n236 & n1451 ;
  assign n4280 = n314 & ~n1565 ;
  assign n4281 = n4280 ^ n314 ;
  assign n4283 = n4282 ^ n4281 ;
  assign n4286 = n188 & n1845 ;
  assign n4284 = n136 & ~n1620 ;
  assign n4285 = n4284 ^ n136 ;
  assign n4287 = n4286 ^ n4285 ;
  assign n4288 = n4283 & n4287 ;
  assign n4289 = n4288 ^ n4283 ;
  assign n4290 = n4289 ^ n4287 ;
  assign n4271 = n188 & n1508 ;
  assign n4269 = n236 & ~n1735 ;
  assign n4270 = n4269 ^ n236 ;
  assign n4272 = n4271 ^ n4270 ;
  assign n4275 = n136 & n1790 ;
  assign n4273 = n314 & ~n1678 ;
  assign n4274 = n4273 ^ n314 ;
  assign n4276 = n4275 ^ n4274 ;
  assign n4277 = n4272 & n4276 ;
  assign n4278 = n4277 ^ n4272 ;
  assign n4279 = n4278 ^ n4276 ;
  assign n4291 = n4290 ^ n4279 ;
  assign n4292 = x134 & n4291 ;
  assign n4293 = n4292 ^ n4291 ;
  assign n4294 = n4293 ^ n4279 ;
  assign n4306 = n236 & n1860 ;
  assign n4307 = n4306 ^ n236 ;
  assign n4308 = n1857 & n4307 ;
  assign n4309 = n4308 ^ n4307 ;
  assign n4310 = n4309 ^ n236 ;
  assign n4311 = n188 & ~n1946 ;
  assign n4312 = n4311 ^ n188 ;
  assign n4313 = n4310 & n4312 ;
  assign n4314 = n4313 ^ n4310 ;
  assign n4315 = n4314 ^ n4312 ;
  assign n4318 = n314 & n1899 ;
  assign n4316 = n136 & ~n1888 ;
  assign n4317 = n4316 ^ n136 ;
  assign n4319 = n4318 ^ n4317 ;
  assign n4320 = n4315 & n4319 ;
  assign n4321 = n4320 ^ n4315 ;
  assign n4322 = n4321 ^ n4319 ;
  assign n4297 = n136 & n1924 ;
  assign n4295 = n314 & ~n1913 ;
  assign n4296 = n4295 ^ n314 ;
  assign n4298 = n4297 ^ n4296 ;
  assign n4301 = n236 & n1935 ;
  assign n4299 = n188 & ~n1874 ;
  assign n4300 = n4299 ^ n188 ;
  assign n4302 = n4301 ^ n4300 ;
  assign n4303 = n4298 & n4302 ;
  assign n4304 = n4303 ^ n4298 ;
  assign n4305 = n4304 ^ n4302 ;
  assign n4323 = n4322 ^ n4305 ;
  assign n4324 = x134 & n4323 ;
  assign n4325 = n4324 ^ n4323 ;
  assign n4326 = n4325 ^ n4305 ;
  assign n4338 = n1960 ^ n236 ;
  assign n4339 = n236 & n4338 ;
  assign n4340 = n4339 ^ n4338 ;
  assign n4341 = n4340 ^ n236 ;
  assign n4342 = n4341 ^ n1965 ;
  assign n4343 = n1966 & n4342 ;
  assign n4344 = n4343 ^ n4340 ;
  assign n4345 = n4344 ^ n1965 ;
  assign n4346 = n188 & n2084 ;
  assign n4347 = n4346 ^ n188 ;
  assign n4348 = n4347 ^ n188 ;
  assign n4349 = n4345 & n4348 ;
  assign n4350 = n4349 ^ n4345 ;
  assign n4351 = n4350 ^ n4348 ;
  assign n4354 = n314 & n2021 ;
  assign n4352 = n136 & ~n2006 ;
  assign n4353 = n4352 ^ n136 ;
  assign n4355 = n4354 ^ n4353 ;
  assign n4356 = n4351 & n4355 ;
  assign n4357 = n4356 ^ n4351 ;
  assign n4358 = n4357 ^ n4355 ;
  assign n4329 = n136 & n2054 ;
  assign n4327 = n314 & ~n2039 ;
  assign n4328 = n4327 ^ n314 ;
  assign n4330 = n4329 ^ n4328 ;
  assign n4333 = n236 & n2069 ;
  assign n4331 = n188 & ~n1987 ;
  assign n4332 = n4331 ^ n188 ;
  assign n4334 = n4333 ^ n4332 ;
  assign n4335 = n4330 & n4334 ;
  assign n4336 = n4335 ^ n4330 ;
  assign n4337 = n4336 ^ n4334 ;
  assign n4359 = n4358 ^ n4337 ;
  assign n4360 = x134 & n4359 ;
  assign n4361 = n4360 ^ n4359 ;
  assign n4362 = n4361 ^ n4337 ;
  assign n4376 = n236 & n2113 ;
  assign n4374 = n188 & ~n2182 ;
  assign n4375 = n4374 ^ n188 ;
  assign n4377 = n4376 ^ n4375 ;
  assign n4380 = n314 & n2135 ;
  assign n4378 = n136 & ~n2124 ;
  assign n4379 = n4378 ^ n136 ;
  assign n4381 = n4380 ^ n4379 ;
  assign n4382 = n4377 & n4381 ;
  assign n4383 = n4382 ^ n4377 ;
  assign n4384 = n4383 ^ n4381 ;
  assign n4365 = n136 & n2160 ;
  assign n4363 = n314 & ~n2149 ;
  assign n4364 = n4363 ^ n314 ;
  assign n4366 = n4365 ^ n4364 ;
  assign n4369 = n236 & n2171 ;
  assign n4367 = n188 & ~n2102 ;
  assign n4368 = n4367 ^ n188 ;
  assign n4370 = n4369 ^ n4368 ;
  assign n4371 = n4366 & n4370 ;
  assign n4372 = n4371 ^ n4366 ;
  assign n4373 = n4372 ^ n4370 ;
  assign n4385 = n4384 ^ n4373 ;
  assign n4386 = x134 & n4385 ;
  assign n4387 = n4386 ^ n4385 ;
  assign n4388 = n4387 ^ n4373 ;
  assign n4402 = n236 & n2218 ;
  assign n4400 = n136 & ~n2233 ;
  assign n4401 = n4400 ^ n136 ;
  assign n4403 = n4402 ^ n4401 ;
  assign n4406 = n188 & n2311 ;
  assign n4404 = n314 & ~n2248 ;
  assign n4405 = n4404 ^ n314 ;
  assign n4407 = n4406 ^ n4405 ;
  assign n4408 = n4403 & n4407 ;
  assign n4409 = n4408 ^ n4403 ;
  assign n4410 = n4409 ^ n4407 ;
  assign n4391 = n188 & n2204 ;
  assign n4389 = n136 & ~n2281 ;
  assign n4390 = n4389 ^ n136 ;
  assign n4392 = n4391 ^ n4390 ;
  assign n4395 = n236 & n2296 ;
  assign n4393 = n314 & ~n2266 ;
  assign n4394 = n4393 ^ n314 ;
  assign n4396 = n4395 ^ n4394 ;
  assign n4397 = n4392 & n4396 ;
  assign n4398 = n4397 ^ n4392 ;
  assign n4399 = n4398 ^ n4396 ;
  assign n4411 = n4410 ^ n4399 ;
  assign n4412 = x134 & n4411 ;
  assign n4413 = n4412 ^ n4411 ;
  assign n4414 = n4413 ^ n4399 ;
  assign n4428 = n236 & n2340 ;
  assign n4426 = n136 & ~n2366 ;
  assign n4427 = n4426 ^ n136 ;
  assign n4429 = n4428 ^ n4427 ;
  assign n4430 = n188 & ~n2416 ;
  assign n4431 = n4430 ^ n188 ;
  assign n4432 = n2345 ^ n314 ;
  assign n4433 = n314 & n4432 ;
  assign n4434 = n4433 ^ n4432 ;
  assign n4435 = n4434 ^ n314 ;
  assign n4436 = n4435 ^ n2348 ;
  assign n4437 = n2349 & n4436 ;
  assign n4438 = n4437 ^ n4434 ;
  assign n4439 = n4438 ^ n2348 ;
  assign n4440 = n4431 & n4439 ;
  assign n4441 = n4440 ^ n4431 ;
  assign n4442 = n4441 ^ n4439 ;
  assign n4443 = n4429 & n4442 ;
  assign n4444 = n4443 ^ n4429 ;
  assign n4445 = n4444 ^ n4442 ;
  assign n4417 = n188 & n2329 ;
  assign n4415 = n136 & ~n2394 ;
  assign n4416 = n4415 ^ n136 ;
  assign n4418 = n4417 ^ n4416 ;
  assign n4421 = n236 & n2405 ;
  assign n4419 = n314 & ~n2383 ;
  assign n4420 = n4419 ^ n314 ;
  assign n4422 = n4421 ^ n4420 ;
  assign n4423 = n4418 & n4422 ;
  assign n4424 = n4423 ^ n4418 ;
  assign n4425 = n4424 ^ n4422 ;
  assign n4446 = n4445 ^ n4425 ;
  assign n4447 = x134 & n4446 ;
  assign n4448 = n4447 ^ n4446 ;
  assign n4449 = n4448 ^ n4425 ;
  assign n4463 = n236 & n2453 ;
  assign n4461 = n136 & ~n2468 ;
  assign n4462 = n4461 ^ n136 ;
  assign n4464 = n4463 ^ n4462 ;
  assign n4467 = n188 & n2546 ;
  assign n4465 = n314 & ~n2483 ;
  assign n4466 = n4465 ^ n314 ;
  assign n4468 = n4467 ^ n4466 ;
  assign n4469 = n4464 & n4468 ;
  assign n4470 = n4469 ^ n4464 ;
  assign n4471 = n4470 ^ n4468 ;
  assign n4452 = n188 & n2438 ;
  assign n4450 = n136 & ~n2516 ;
  assign n4451 = n4450 ^ n136 ;
  assign n4453 = n4452 ^ n4451 ;
  assign n4456 = n236 & n2531 ;
  assign n4454 = n314 & ~n2501 ;
  assign n4455 = n4454 ^ n314 ;
  assign n4457 = n4456 ^ n4455 ;
  assign n4458 = n4453 & n4457 ;
  assign n4459 = n4458 ^ n4453 ;
  assign n4460 = n4459 ^ n4457 ;
  assign n4472 = n4471 ^ n4460 ;
  assign n4473 = x134 & n4472 ;
  assign n4474 = n4473 ^ n4472 ;
  assign n4475 = n4474 ^ n4460 ;
  assign n4489 = n236 & n2575 ;
  assign n4487 = n188 & ~n2646 ;
  assign n4488 = n4487 ^ n188 ;
  assign n4490 = n4489 ^ n4488 ;
  assign n4493 = n314 & n2599 ;
  assign n4491 = n136 & ~n2586 ;
  assign n4492 = n4491 ^ n136 ;
  assign n4494 = n4493 ^ n4492 ;
  assign n4495 = n4490 & n4494 ;
  assign n4496 = n4495 ^ n4490 ;
  assign n4497 = n4496 ^ n4494 ;
  assign n4478 = n188 & n2564 ;
  assign n4476 = n136 & ~n2624 ;
  assign n4477 = n4476 ^ n136 ;
  assign n4479 = n4478 ^ n4477 ;
  assign n4482 = n236 & n2635 ;
  assign n4480 = n314 & ~n2613 ;
  assign n4481 = n4480 ^ n314 ;
  assign n4483 = n4482 ^ n4481 ;
  assign n4484 = n4479 & n4483 ;
  assign n4485 = n4484 ^ n4479 ;
  assign n4486 = n4485 ^ n4483 ;
  assign n4498 = n4497 ^ n4486 ;
  assign n4499 = x134 & n4498 ;
  assign n4500 = n4499 ^ n4498 ;
  assign n4501 = n4500 ^ n4486 ;
  assign n4515 = n236 & n2683 ;
  assign n4513 = n188 & ~n2776 ;
  assign n4514 = n4513 ^ n188 ;
  assign n4516 = n4515 ^ n4514 ;
  assign n4519 = n314 & n2713 ;
  assign n4517 = n136 & ~n2698 ;
  assign n4518 = n4517 ^ n136 ;
  assign n4520 = n4519 ^ n4518 ;
  assign n4521 = n4516 & n4520 ;
  assign n4522 = n4521 ^ n4516 ;
  assign n4523 = n4522 ^ n4520 ;
  assign n4504 = n188 & n2668 ;
  assign n4502 = n136 & ~n2746 ;
  assign n4503 = n4502 ^ n136 ;
  assign n4505 = n4504 ^ n4503 ;
  assign n4508 = n236 & n2761 ;
  assign n4506 = n314 & ~n2731 ;
  assign n4507 = n4506 ^ n314 ;
  assign n4509 = n4508 ^ n4507 ;
  assign n4510 = n4505 & n4509 ;
  assign n4511 = n4510 ^ n4505 ;
  assign n4512 = n4511 ^ n4509 ;
  assign n4524 = n4523 ^ n4512 ;
  assign n4525 = x134 & n4524 ;
  assign n4526 = n4525 ^ n4524 ;
  assign n4527 = n4526 ^ n4512 ;
  assign n4541 = n236 & n2805 ;
  assign n4539 = n188 & ~n2883 ;
  assign n4540 = n4539 ^ n188 ;
  assign n4542 = n4541 ^ n4540 ;
  assign n4543 = n2810 ^ n314 ;
  assign n4544 = n314 & n4543 ;
  assign n4545 = n4544 ^ n4543 ;
  assign n4546 = n4545 ^ n314 ;
  assign n4547 = n4546 ^ n2815 ;
  assign n4548 = n2816 & n4547 ;
  assign n4549 = n4548 ^ n4545 ;
  assign n4550 = n4549 ^ n2815 ;
  assign n4551 = n136 & ~n2833 ;
  assign n4552 = n4551 ^ n136 ;
  assign n4553 = n4550 & n4552 ;
  assign n4554 = n4553 ^ n4550 ;
  assign n4555 = n4554 ^ n4552 ;
  assign n4556 = n4542 & n4555 ;
  assign n4557 = n4556 ^ n4542 ;
  assign n4558 = n4557 ^ n4555 ;
  assign n4530 = n188 & n2794 ;
  assign n4528 = n136 & ~n2861 ;
  assign n4529 = n4528 ^ n136 ;
  assign n4531 = n4530 ^ n4529 ;
  assign n4534 = n236 & n2872 ;
  assign n4532 = n314 & ~n2850 ;
  assign n4533 = n4532 ^ n314 ;
  assign n4535 = n4534 ^ n4533 ;
  assign n4536 = n4531 & n4535 ;
  assign n4537 = n4536 ^ n4531 ;
  assign n4538 = n4537 ^ n4535 ;
  assign n4559 = n4558 ^ n4538 ;
  assign n4560 = x134 & n4559 ;
  assign n4561 = n4560 ^ n4559 ;
  assign n4562 = n4561 ^ n4538 ;
  assign n4576 = n236 & n2920 ;
  assign n4574 = n188 & ~n3017 ;
  assign n4575 = n4574 ^ n188 ;
  assign n4577 = n4576 ^ n4575 ;
  assign n4578 = n314 & n2932 ;
  assign n4579 = n4578 ^ n314 ;
  assign n4580 = n2927 & n4579 ;
  assign n4581 = n4580 ^ n4579 ;
  assign n4582 = n4581 ^ n314 ;
  assign n4583 = n136 & n2950 ;
  assign n4584 = n4583 ^ n136 ;
  assign n4585 = n4584 ^ n136 ;
  assign n4586 = n4582 & n4585 ;
  assign n4587 = n4586 ^ n4582 ;
  assign n4588 = n4587 ^ n4585 ;
  assign n4589 = n4577 & n4588 ;
  assign n4590 = n4589 ^ n4577 ;
  assign n4591 = n4590 ^ n4588 ;
  assign n4565 = n188 & n2905 ;
  assign n4563 = n136 & ~n2987 ;
  assign n4564 = n4563 ^ n136 ;
  assign n4566 = n4565 ^ n4564 ;
  assign n4569 = n236 & n3002 ;
  assign n4567 = n314 & ~n2972 ;
  assign n4568 = n4567 ^ n314 ;
  assign n4570 = n4569 ^ n4568 ;
  assign n4571 = n4566 & n4570 ;
  assign n4572 = n4571 ^ n4566 ;
  assign n4573 = n4572 ^ n4570 ;
  assign n4592 = n4591 ^ n4573 ;
  assign n4593 = x134 & n4592 ;
  assign n4594 = n4593 ^ n4592 ;
  assign n4595 = n4594 ^ n4573 ;
  assign n4609 = n236 & n3046 ;
  assign n4607 = n188 & ~n3119 ;
  assign n4608 = n4607 ^ n188 ;
  assign n4610 = n4609 ^ n4608 ;
  assign n4613 = n314 & n3072 ;
  assign n4611 = n136 & ~n3057 ;
  assign n4612 = n4611 ^ n136 ;
  assign n4614 = n4613 ^ n4612 ;
  assign n4615 = n4610 & n4614 ;
  assign n4616 = n4615 ^ n4610 ;
  assign n4617 = n4616 ^ n4614 ;
  assign n4598 = n188 & n3035 ;
  assign n4596 = n136 & ~n3097 ;
  assign n4597 = n4596 ^ n136 ;
  assign n4599 = n4598 ^ n4597 ;
  assign n4602 = n236 & n3108 ;
  assign n4600 = n314 & ~n3086 ;
  assign n4601 = n4600 ^ n314 ;
  assign n4603 = n4602 ^ n4601 ;
  assign n4604 = n4599 & n4603 ;
  assign n4605 = n4604 ^ n4599 ;
  assign n4606 = n4605 ^ n4603 ;
  assign n4618 = n4617 ^ n4606 ;
  assign n4619 = x134 & n4618 ;
  assign n4620 = n4619 ^ n4618 ;
  assign n4621 = n4620 ^ n4606 ;
  assign n4635 = n236 & n3156 ;
  assign n4633 = n188 & ~n3249 ;
  assign n4634 = n4633 ^ n188 ;
  assign n4636 = n4635 ^ n4634 ;
  assign n4639 = n314 & n3186 ;
  assign n4637 = n136 & ~n3171 ;
  assign n4638 = n4637 ^ n136 ;
  assign n4640 = n4639 ^ n4638 ;
  assign n4641 = n4636 & n4640 ;
  assign n4642 = n4641 ^ n4636 ;
  assign n4643 = n4642 ^ n4640 ;
  assign n4624 = n188 & n3141 ;
  assign n4622 = n136 & ~n3219 ;
  assign n4623 = n4622 ^ n136 ;
  assign n4625 = n4624 ^ n4623 ;
  assign n4628 = n236 & n3234 ;
  assign n4626 = n314 & ~n3204 ;
  assign n4627 = n4626 ^ n314 ;
  assign n4629 = n4628 ^ n4627 ;
  assign n4630 = n4625 & n4629 ;
  assign n4631 = n4630 ^ n4625 ;
  assign n4632 = n4631 ^ n4629 ;
  assign n4644 = n4643 ^ n4632 ;
  assign n4645 = x134 & n4644 ;
  assign n4646 = n4645 ^ n4644 ;
  assign n4647 = n4646 ^ n4632 ;
  assign n4648 = n540 ^ n346 ;
  assign n4649 = n1168 ^ n847 ;
  assign n4650 = n1393 ^ n1287 ;
  assign n4651 = n1852 ^ n1625 ;
  assign n4652 = n1953 ^ n1904 ;
  assign n4653 = n2091 ^ n2026 ;
  assign n4654 = n2189 ^ n2140 ;
  assign n4655 = n2318 ^ n2253 ;
  assign n4656 = n2423 ^ n2374 ;
  assign n4657 = n2553 ^ n2488 ;
  assign n4658 = n2653 ^ n2604 ;
  assign n4659 = n2783 ^ n2718 ;
  assign n4660 = n2890 ^ n2841 ;
  assign n4661 = n3024 ^ n2959 ;
  assign n4662 = n3126 ^ n3077 ;
  assign n4663 = n3256 ^ n3191 ;
  assign n4664 = n3288 ^ n3275 ;
  assign n4665 = n3314 ^ n3301 ;
  assign n4666 = n3340 ^ n3327 ;
  assign n4667 = n3366 ^ n3353 ;
  assign n4668 = n3398 ^ n3385 ;
  assign n4669 = n3434 ^ n3421 ;
  assign n4670 = n3460 ^ n3447 ;
  assign n4671 = n3486 ^ n3473 ;
  assign n4672 = n3521 ^ n3508 ;
  assign n4673 = n3547 ^ n3534 ;
  assign n4674 = n3573 ^ n3560 ;
  assign n4675 = n3599 ^ n3586 ;
  assign n4676 = n3634 ^ n3621 ;
  assign n4677 = n3667 ^ n3654 ;
  assign n4678 = n3693 ^ n3680 ;
  assign n4679 = n3719 ^ n3706 ;
  assign n4680 = n3751 ^ n3738 ;
  assign n4681 = n3777 ^ n3764 ;
  assign n4682 = n3803 ^ n3790 ;
  assign n4683 = n3829 ^ n3816 ;
  assign n4684 = n3861 ^ n3848 ;
  assign n4685 = n3897 ^ n3884 ;
  assign n4686 = n3923 ^ n3910 ;
  assign n4687 = n3949 ^ n3936 ;
  assign n4688 = n3984 ^ n3962 ;
  assign n4689 = n4010 ^ n3997 ;
  assign n4690 = n4036 ^ n4023 ;
  assign n4691 = n4062 ^ n4049 ;
  assign n4692 = n4097 ^ n4075 ;
  assign n4693 = n4130 ^ n4110 ;
  assign n4694 = n4156 ^ n4143 ;
  assign n4695 = n4182 ^ n4169 ;
  assign n4696 = n4214 ^ n4195 ;
  assign n4697 = n4240 ^ n4227 ;
  assign n4698 = n4266 ^ n4253 ;
  assign n4699 = n4292 ^ n4279 ;
  assign n4700 = n4324 ^ n4305 ;
  assign n4701 = n4360 ^ n4337 ;
  assign n4702 = n4386 ^ n4373 ;
  assign n4703 = n4412 ^ n4399 ;
  assign n4704 = n4447 ^ n4425 ;
  assign n4705 = n4473 ^ n4460 ;
  assign n4706 = n4499 ^ n4486 ;
  assign n4707 = n4525 ^ n4512 ;
  assign n4708 = n4560 ^ n4538 ;
  assign n4709 = n4593 ^ n4573 ;
  assign n4710 = n4619 ^ n4606 ;
  assign n4711 = n4645 ^ n4632 ;
  assign y0 = n542 ;
  assign y1 = n1170 ;
  assign y2 = n1395 ;
  assign y3 = n1854 ;
  assign y4 = n1955 ;
  assign y5 = n2093 ;
  assign y6 = n2191 ;
  assign y7 = n2320 ;
  assign y8 = n2425 ;
  assign y9 = n2555 ;
  assign y10 = n2655 ;
  assign y11 = n2785 ;
  assign y12 = n2892 ;
  assign y13 = n3026 ;
  assign y14 = n3128 ;
  assign y15 = n3258 ;
  assign y16 = n3290 ;
  assign y17 = n3316 ;
  assign y18 = n3342 ;
  assign y19 = n3368 ;
  assign y20 = n3400 ;
  assign y21 = n3436 ;
  assign y22 = n3462 ;
  assign y23 = n3488 ;
  assign y24 = n3523 ;
  assign y25 = n3549 ;
  assign y26 = n3575 ;
  assign y27 = n3601 ;
  assign y28 = n3636 ;
  assign y29 = n3669 ;
  assign y30 = n3695 ;
  assign y31 = n3721 ;
  assign y32 = n3753 ;
  assign y33 = n3779 ;
  assign y34 = n3805 ;
  assign y35 = n3831 ;
  assign y36 = n3863 ;
  assign y37 = n3899 ;
  assign y38 = n3925 ;
  assign y39 = n3951 ;
  assign y40 = n3986 ;
  assign y41 = n4012 ;
  assign y42 = n4038 ;
  assign y43 = n4064 ;
  assign y44 = n4099 ;
  assign y45 = n4132 ;
  assign y46 = n4158 ;
  assign y47 = n4184 ;
  assign y48 = n4216 ;
  assign y49 = n4242 ;
  assign y50 = n4268 ;
  assign y51 = n4294 ;
  assign y52 = n4326 ;
  assign y53 = n4362 ;
  assign y54 = n4388 ;
  assign y55 = n4414 ;
  assign y56 = n4449 ;
  assign y57 = n4475 ;
  assign y58 = n4501 ;
  assign y59 = n4527 ;
  assign y60 = n4562 ;
  assign y61 = n4595 ;
  assign y62 = n4621 ;
  assign y63 = n4647 ;
  assign y64 = n4648 ;
  assign y65 = n4649 ;
  assign y66 = n4650 ;
  assign y67 = n4651 ;
  assign y68 = n4652 ;
  assign y69 = n4653 ;
  assign y70 = n4654 ;
  assign y71 = n4655 ;
  assign y72 = n4656 ;
  assign y73 = n4657 ;
  assign y74 = n4658 ;
  assign y75 = n4659 ;
  assign y76 = n4660 ;
  assign y77 = n4661 ;
  assign y78 = n4662 ;
  assign y79 = n4663 ;
  assign y80 = n4664 ;
  assign y81 = n4665 ;
  assign y82 = n4666 ;
  assign y83 = n4667 ;
  assign y84 = n4668 ;
  assign y85 = n4669 ;
  assign y86 = n4670 ;
  assign y87 = n4671 ;
  assign y88 = n4672 ;
  assign y89 = n4673 ;
  assign y90 = n4674 ;
  assign y91 = n4675 ;
  assign y92 = n4676 ;
  assign y93 = n4677 ;
  assign y94 = n4678 ;
  assign y95 = n4679 ;
  assign y96 = n4680 ;
  assign y97 = n4681 ;
  assign y98 = n4682 ;
  assign y99 = n4683 ;
  assign y100 = n4684 ;
  assign y101 = n4685 ;
  assign y102 = n4686 ;
  assign y103 = n4687 ;
  assign y104 = n4688 ;
  assign y105 = n4689 ;
  assign y106 = n4690 ;
  assign y107 = n4691 ;
  assign y108 = n4692 ;
  assign y109 = n4693 ;
  assign y110 = n4694 ;
  assign y111 = n4695 ;
  assign y112 = n4696 ;
  assign y113 = n4697 ;
  assign y114 = n4698 ;
  assign y115 = n4699 ;
  assign y116 = n4700 ;
  assign y117 = n4701 ;
  assign y118 = n4702 ;
  assign y119 = n4703 ;
  assign y120 = n4704 ;
  assign y121 = n4705 ;
  assign y122 = n4706 ;
  assign y123 = n4707 ;
  assign y124 = n4708 ;
  assign y125 = n4709 ;
  assign y126 = n4710 ;
  assign y127 = n4711 ;
endmodule
