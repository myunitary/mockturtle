// Benchmark "/tmp/tmp" written by ABC on Wed Nov 12 17:23:41 2025

module adder_opt ( 
    n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
    n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127, po128  );
  input  n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
    n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
    n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127, po128;
  wire new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933;
  assign new_n257 = n129 ^ n1;
  assign new_n258 = n1 & n129;
  assign new_n259 = n130 ^ n2;
  assign new_n260 = new_n259 ^ new_n258;
  assign new_n261 = n131 ^ n3;
  assign new_n262 = new_n258 ^ n130;
  assign new_n263 = ~new_n262 & new_n259;
  assign new_n264 = new_n263 ^ n2;
  assign new_n265 = new_n264 ^ new_n261;
  assign new_n266 = n132 ^ n4;
  assign new_n267 = new_n264 ^ n131;
  assign new_n268 = ~new_n267 & new_n261;
  assign new_n269 = new_n268 ^ n3;
  assign new_n270 = new_n269 ^ new_n266;
  assign new_n271 = n133 ^ n5;
  assign new_n272 = new_n269 ^ n132;
  assign new_n273 = ~new_n272 & new_n266;
  assign new_n274 = new_n273 ^ n4;
  assign new_n275 = new_n274 ^ new_n271;
  assign new_n276 = n134 ^ n6;
  assign new_n277 = n133 ^ n4;
  assign new_n278 = new_n277 ^ new_n273;
  assign new_n279 = ~new_n278 & new_n271;
  assign new_n280 = new_n279 ^ n5;
  assign new_n281 = new_n280 ^ new_n276;
  assign new_n282 = n135 ^ n7;
  assign new_n283 = new_n280 ^ n134;
  assign new_n284 = ~new_n283 & new_n276;
  assign new_n285 = new_n284 ^ n6;
  assign new_n286 = new_n285 ^ new_n282;
  assign new_n287 = n136 ^ n8;
  assign new_n288 = n135 ^ n6;
  assign new_n289 = new_n288 ^ new_n284;
  assign new_n290 = ~new_n289 & new_n282;
  assign new_n291 = new_n290 ^ n7;
  assign new_n292 = new_n291 ^ new_n287;
  assign new_n293 = n137 ^ n9;
  assign new_n294 = new_n291 ^ n136;
  assign new_n295 = ~new_n294 & new_n287;
  assign new_n296 = new_n295 ^ n8;
  assign new_n297 = new_n296 ^ new_n293;
  assign new_n298 = n138 ^ n10;
  assign new_n299 = n137 ^ n8;
  assign new_n300 = new_n299 ^ new_n295;
  assign new_n301 = ~new_n300 & new_n293;
  assign new_n302 = new_n301 ^ n9;
  assign new_n303 = new_n302 ^ new_n298;
  assign new_n304 = new_n302 ^ n138;
  assign new_n305 = ~new_n304 & new_n298;
  assign new_n306 = new_n305 ^ n10;
  assign new_n307 = n139 ^ n11;
  assign new_n308 = new_n307 ^ new_n306;
  assign new_n309 = n140 ^ n12;
  assign new_n310 = new_n306 ^ n139;
  assign new_n311 = ~new_n310 & new_n307;
  assign new_n312 = new_n311 ^ n11;
  assign new_n313 = new_n312 ^ new_n309;
  assign new_n314 = n141 ^ n13;
  assign new_n315 = new_n312 ^ n140;
  assign new_n316 = ~new_n315 & new_n309;
  assign new_n317 = new_n316 ^ n12;
  assign new_n318 = new_n317 ^ new_n314;
  assign new_n319 = n142 ^ n14;
  assign new_n320 = n141 ^ n12;
  assign new_n321 = new_n320 ^ new_n316;
  assign new_n322 = ~new_n321 & new_n314;
  assign new_n323 = new_n322 ^ n13;
  assign new_n324 = new_n323 ^ new_n319;
  assign new_n325 = n143 ^ n15;
  assign new_n326 = new_n323 ^ n142;
  assign new_n327 = ~new_n326 & new_n319;
  assign new_n328 = new_n327 ^ n14;
  assign new_n329 = new_n328 ^ new_n325;
  assign new_n330 = n144 ^ n16;
  assign new_n331 = n143 ^ n14;
  assign new_n332 = new_n331 ^ new_n327;
  assign new_n333 = ~new_n332 & new_n325;
  assign new_n334 = new_n333 ^ n15;
  assign new_n335 = new_n334 ^ new_n330;
  assign new_n336 = n145 ^ n17;
  assign new_n337 = new_n334 ^ n144;
  assign new_n338 = ~new_n337 & new_n330;
  assign new_n339 = new_n338 ^ n16;
  assign new_n340 = new_n339 ^ new_n336;
  assign new_n341 = n146 ^ n18;
  assign new_n342 = n145 ^ n16;
  assign new_n343 = new_n342 ^ new_n338;
  assign new_n344 = ~new_n343 & new_n336;
  assign new_n345 = new_n344 ^ n17;
  assign new_n346 = new_n345 ^ new_n341;
  assign new_n347 = n147 ^ n19;
  assign new_n348 = new_n345 ^ n146;
  assign new_n349 = ~new_n348 & new_n341;
  assign new_n350 = new_n349 ^ n18;
  assign new_n351 = new_n350 ^ new_n347;
  assign new_n352 = n148 ^ n20;
  assign new_n353 = n147 ^ n18;
  assign new_n354 = new_n353 ^ new_n349;
  assign new_n355 = ~new_n354 & new_n347;
  assign new_n356 = new_n355 ^ n19;
  assign new_n357 = new_n356 ^ new_n352;
  assign new_n358 = new_n356 ^ n148;
  assign new_n359 = ~new_n358 & new_n352;
  assign new_n360 = new_n359 ^ n20;
  assign new_n361 = n149 ^ n21;
  assign new_n362 = new_n361 ^ new_n360;
  assign new_n363 = n150 ^ n22;
  assign new_n364 = new_n360 ^ n149;
  assign new_n365 = ~new_n364 & new_n361;
  assign new_n366 = new_n365 ^ n21;
  assign new_n367 = new_n366 ^ new_n363;
  assign new_n368 = n151 ^ n23;
  assign new_n369 = new_n366 ^ n150;
  assign new_n370 = ~new_n369 & new_n363;
  assign new_n371 = new_n370 ^ n22;
  assign new_n372 = new_n371 ^ new_n368;
  assign new_n373 = n152 ^ n24;
  assign new_n374 = n151 ^ n22;
  assign new_n375 = new_n374 ^ new_n370;
  assign new_n376 = ~new_n375 & new_n368;
  assign new_n377 = new_n376 ^ n23;
  assign new_n378 = new_n377 ^ new_n373;
  assign new_n379 = n153 ^ n25;
  assign new_n380 = new_n377 ^ n152;
  assign new_n381 = ~new_n380 & new_n373;
  assign new_n382 = new_n381 ^ n24;
  assign new_n383 = new_n382 ^ new_n379;
  assign new_n384 = n154 ^ n26;
  assign new_n385 = n153 ^ n24;
  assign new_n386 = new_n385 ^ new_n381;
  assign new_n387 = ~new_n386 & new_n379;
  assign new_n388 = new_n387 ^ n25;
  assign new_n389 = new_n388 ^ new_n384;
  assign new_n390 = n155 ^ n27;
  assign new_n391 = new_n388 ^ n154;
  assign new_n392 = ~new_n391 & new_n384;
  assign new_n393 = new_n392 ^ n26;
  assign new_n394 = new_n393 ^ new_n390;
  assign new_n395 = n156 ^ n28;
  assign new_n396 = n155 ^ n26;
  assign new_n397 = new_n396 ^ new_n392;
  assign new_n398 = ~new_n397 & new_n390;
  assign new_n399 = new_n398 ^ n27;
  assign new_n400 = new_n399 ^ new_n395;
  assign new_n401 = n157 ^ n29;
  assign new_n402 = new_n399 ^ n156;
  assign new_n403 = ~new_n402 & new_n395;
  assign new_n404 = new_n403 ^ n28;
  assign new_n405 = new_n404 ^ new_n401;
  assign new_n406 = n158 ^ n30;
  assign new_n407 = n157 ^ n28;
  assign new_n408 = new_n407 ^ new_n403;
  assign new_n409 = ~new_n408 & new_n401;
  assign new_n410 = new_n409 ^ n29;
  assign new_n411 = new_n410 ^ new_n406;
  assign new_n412 = new_n410 ^ n158;
  assign new_n413 = ~new_n412 & new_n406;
  assign new_n414 = new_n413 ^ n30;
  assign new_n415 = n159 ^ n31;
  assign new_n416 = new_n415 ^ new_n414;
  assign new_n417 = n160 ^ n32;
  assign new_n418 = new_n414 ^ n159;
  assign new_n419 = ~new_n418 & new_n415;
  assign new_n420 = new_n419 ^ n31;
  assign new_n421 = new_n420 ^ new_n417;
  assign new_n422 = n161 ^ n33;
  assign new_n423 = new_n420 ^ n160;
  assign new_n424 = ~new_n423 & new_n417;
  assign new_n425 = new_n424 ^ n32;
  assign new_n426 = new_n425 ^ new_n422;
  assign new_n427 = n162 ^ n34;
  assign new_n428 = n161 ^ n32;
  assign new_n429 = new_n428 ^ new_n424;
  assign new_n430 = ~new_n429 & new_n422;
  assign new_n431 = new_n430 ^ n33;
  assign new_n432 = new_n431 ^ new_n427;
  assign new_n433 = n163 ^ n35;
  assign new_n434 = new_n431 ^ n162;
  assign new_n435 = ~new_n434 & new_n427;
  assign new_n436 = new_n435 ^ n34;
  assign new_n437 = new_n436 ^ new_n433;
  assign new_n438 = n164 ^ n36;
  assign new_n439 = n163 ^ n34;
  assign new_n440 = new_n439 ^ new_n435;
  assign new_n441 = ~new_n440 & new_n433;
  assign new_n442 = new_n441 ^ n35;
  assign new_n443 = new_n442 ^ new_n438;
  assign new_n444 = n165 ^ n37;
  assign new_n445 = new_n442 ^ n164;
  assign new_n446 = ~new_n445 & new_n438;
  assign new_n447 = new_n446 ^ n36;
  assign new_n448 = new_n447 ^ new_n444;
  assign new_n449 = n166 ^ n38;
  assign new_n450 = n165 ^ n36;
  assign new_n451 = new_n450 ^ new_n446;
  assign new_n452 = ~new_n451 & new_n444;
  assign new_n453 = new_n452 ^ n37;
  assign new_n454 = new_n453 ^ new_n449;
  assign new_n455 = n167 ^ n39;
  assign new_n456 = new_n453 ^ n166;
  assign new_n457 = ~new_n456 & new_n449;
  assign new_n458 = new_n457 ^ n38;
  assign new_n459 = new_n458 ^ new_n455;
  assign new_n460 = n168 ^ n40;
  assign new_n461 = n167 ^ n38;
  assign new_n462 = new_n461 ^ new_n457;
  assign new_n463 = ~new_n462 & new_n455;
  assign new_n464 = new_n463 ^ n39;
  assign new_n465 = new_n464 ^ new_n460;
  assign new_n466 = new_n464 ^ n168;
  assign new_n467 = ~new_n466 & new_n460;
  assign new_n468 = new_n467 ^ n40;
  assign new_n469 = n169 ^ n41;
  assign new_n470 = new_n469 ^ new_n468;
  assign new_n471 = n170 ^ n42;
  assign new_n472 = new_n468 ^ n169;
  assign new_n473 = ~new_n472 & new_n469;
  assign new_n474 = new_n473 ^ n41;
  assign new_n475 = new_n474 ^ new_n471;
  assign new_n476 = n171 ^ n43;
  assign new_n477 = new_n474 ^ n170;
  assign new_n478 = ~new_n477 & new_n471;
  assign new_n479 = new_n478 ^ n42;
  assign new_n480 = new_n479 ^ new_n476;
  assign new_n481 = n172 ^ n44;
  assign new_n482 = n171 ^ n42;
  assign new_n483 = new_n482 ^ new_n478;
  assign new_n484 = ~new_n483 & new_n476;
  assign new_n485 = new_n484 ^ n43;
  assign new_n486 = new_n485 ^ new_n481;
  assign new_n487 = n173 ^ n45;
  assign new_n488 = new_n485 ^ n172;
  assign new_n489 = ~new_n488 & new_n481;
  assign new_n490 = new_n489 ^ n44;
  assign new_n491 = new_n490 ^ new_n487;
  assign new_n492 = n174 ^ n46;
  assign new_n493 = n173 ^ n44;
  assign new_n494 = new_n493 ^ new_n489;
  assign new_n495 = ~new_n494 & new_n487;
  assign new_n496 = new_n495 ^ n45;
  assign new_n497 = new_n496 ^ new_n492;
  assign new_n498 = n175 ^ n47;
  assign new_n499 = new_n496 ^ n174;
  assign new_n500 = ~new_n499 & new_n492;
  assign new_n501 = new_n500 ^ n46;
  assign new_n502 = new_n501 ^ new_n498;
  assign new_n503 = n176 ^ n48;
  assign new_n504 = n175 ^ n46;
  assign new_n505 = new_n504 ^ new_n500;
  assign new_n506 = ~new_n505 & new_n498;
  assign new_n507 = new_n506 ^ n47;
  assign new_n508 = new_n507 ^ new_n503;
  assign new_n509 = n177 ^ n49;
  assign new_n510 = new_n507 ^ n176;
  assign new_n511 = ~new_n510 & new_n503;
  assign new_n512 = new_n511 ^ n48;
  assign new_n513 = new_n512 ^ new_n509;
  assign new_n514 = n178 ^ n50;
  assign new_n515 = n177 ^ n48;
  assign new_n516 = new_n515 ^ new_n511;
  assign new_n517 = ~new_n516 & new_n509;
  assign new_n518 = new_n517 ^ n49;
  assign new_n519 = new_n518 ^ new_n514;
  assign new_n520 = new_n518 ^ n178;
  assign new_n521 = ~new_n520 & new_n514;
  assign new_n522 = new_n521 ^ n50;
  assign new_n523 = n179 ^ n51;
  assign new_n524 = new_n523 ^ new_n522;
  assign new_n525 = n180 ^ n52;
  assign new_n526 = new_n522 ^ n179;
  assign new_n527 = ~new_n526 & new_n523;
  assign new_n528 = new_n527 ^ n51;
  assign new_n529 = new_n528 ^ new_n525;
  assign new_n530 = n181 ^ n53;
  assign new_n531 = new_n528 ^ n180;
  assign new_n532 = ~new_n531 & new_n525;
  assign new_n533 = new_n532 ^ n52;
  assign new_n534 = new_n533 ^ new_n530;
  assign new_n535 = n182 ^ n54;
  assign new_n536 = n181 ^ n52;
  assign new_n537 = new_n536 ^ new_n532;
  assign new_n538 = ~new_n537 & new_n530;
  assign new_n539 = new_n538 ^ n53;
  assign new_n540 = new_n539 ^ new_n535;
  assign new_n541 = n183 ^ n55;
  assign new_n542 = new_n539 ^ n182;
  assign new_n543 = ~new_n542 & new_n535;
  assign new_n544 = new_n543 ^ n54;
  assign new_n545 = new_n544 ^ new_n541;
  assign new_n546 = n184 ^ n56;
  assign new_n547 = n183 ^ n54;
  assign new_n548 = new_n547 ^ new_n543;
  assign new_n549 = ~new_n548 & new_n541;
  assign new_n550 = new_n549 ^ n55;
  assign new_n551 = new_n550 ^ new_n546;
  assign new_n552 = n185 ^ n57;
  assign new_n553 = new_n550 ^ n184;
  assign new_n554 = ~new_n553 & new_n546;
  assign new_n555 = new_n554 ^ n56;
  assign new_n556 = new_n555 ^ new_n552;
  assign new_n557 = n186 ^ n58;
  assign new_n558 = n185 ^ n56;
  assign new_n559 = new_n558 ^ new_n554;
  assign new_n560 = ~new_n559 & new_n552;
  assign new_n561 = new_n560 ^ n57;
  assign new_n562 = new_n561 ^ new_n557;
  assign new_n563 = n187 ^ n59;
  assign new_n564 = new_n561 ^ n186;
  assign new_n565 = ~new_n564 & new_n557;
  assign new_n566 = new_n565 ^ n58;
  assign new_n567 = new_n566 ^ new_n563;
  assign new_n568 = n188 ^ n60;
  assign new_n569 = n187 ^ n58;
  assign new_n570 = new_n569 ^ new_n565;
  assign new_n571 = ~new_n570 & new_n563;
  assign new_n572 = new_n571 ^ n59;
  assign new_n573 = new_n572 ^ new_n568;
  assign new_n574 = new_n572 ^ n188;
  assign new_n575 = ~new_n574 & new_n568;
  assign new_n576 = new_n575 ^ n60;
  assign new_n577 = n189 ^ n61;
  assign new_n578 = new_n577 ^ new_n576;
  assign new_n579 = n190 ^ n62;
  assign new_n580 = new_n576 ^ n189;
  assign new_n581 = ~new_n580 & new_n577;
  assign new_n582 = new_n581 ^ n61;
  assign new_n583 = new_n582 ^ new_n579;
  assign new_n584 = n191 ^ n63;
  assign new_n585 = new_n582 ^ n190;
  assign new_n586 = ~new_n585 & new_n579;
  assign new_n587 = new_n586 ^ n62;
  assign new_n588 = new_n587 ^ new_n584;
  assign new_n589 = n192 ^ n64;
  assign new_n590 = n191 ^ n62;
  assign new_n591 = new_n590 ^ new_n586;
  assign new_n592 = ~new_n591 & new_n584;
  assign new_n593 = new_n592 ^ n63;
  assign new_n594 = new_n593 ^ new_n589;
  assign new_n595 = n193 ^ n65;
  assign new_n596 = new_n593 ^ n192;
  assign new_n597 = ~new_n596 & new_n589;
  assign new_n598 = new_n597 ^ n64;
  assign new_n599 = new_n598 ^ new_n595;
  assign new_n600 = n194 ^ n66;
  assign new_n601 = n193 ^ n64;
  assign new_n602 = new_n601 ^ new_n597;
  assign new_n603 = ~new_n602 & new_n595;
  assign new_n604 = new_n603 ^ n65;
  assign new_n605 = new_n604 ^ new_n600;
  assign new_n606 = n195 ^ n67;
  assign new_n607 = new_n604 ^ n194;
  assign new_n608 = ~new_n607 & new_n600;
  assign new_n609 = new_n608 ^ n66;
  assign new_n610 = new_n609 ^ new_n606;
  assign new_n611 = n196 ^ n68;
  assign new_n612 = n195 ^ n66;
  assign new_n613 = new_n612 ^ new_n608;
  assign new_n614 = ~new_n613 & new_n606;
  assign new_n615 = new_n614 ^ n67;
  assign new_n616 = new_n615 ^ new_n611;
  assign new_n617 = n197 ^ n69;
  assign new_n618 = new_n615 ^ n196;
  assign new_n619 = ~new_n618 & new_n611;
  assign new_n620 = new_n619 ^ n68;
  assign new_n621 = new_n620 ^ new_n617;
  assign new_n622 = n198 ^ n70;
  assign new_n623 = n197 ^ n68;
  assign new_n624 = new_n623 ^ new_n619;
  assign new_n625 = ~new_n624 & new_n617;
  assign new_n626 = new_n625 ^ n69;
  assign new_n627 = new_n626 ^ new_n622;
  assign new_n628 = new_n626 ^ n198;
  assign new_n629 = ~new_n628 & new_n622;
  assign new_n630 = new_n629 ^ n70;
  assign new_n631 = n199 ^ n71;
  assign new_n632 = new_n631 ^ new_n630;
  assign new_n633 = n200 ^ n72;
  assign new_n634 = new_n630 ^ n199;
  assign new_n635 = ~new_n634 & new_n631;
  assign new_n636 = new_n635 ^ n71;
  assign new_n637 = new_n636 ^ new_n633;
  assign new_n638 = n201 ^ n73;
  assign new_n639 = new_n636 ^ n200;
  assign new_n640 = ~new_n639 & new_n633;
  assign new_n641 = new_n640 ^ n72;
  assign new_n642 = new_n641 ^ new_n638;
  assign new_n643 = n202 ^ n74;
  assign new_n644 = n201 ^ n72;
  assign new_n645 = new_n644 ^ new_n640;
  assign new_n646 = ~new_n645 & new_n638;
  assign new_n647 = new_n646 ^ n73;
  assign new_n648 = new_n647 ^ new_n643;
  assign new_n649 = n203 ^ n75;
  assign new_n650 = new_n647 ^ n202;
  assign new_n651 = ~new_n650 & new_n643;
  assign new_n652 = new_n651 ^ n74;
  assign new_n653 = new_n652 ^ new_n649;
  assign new_n654 = n204 ^ n76;
  assign new_n655 = n203 ^ n74;
  assign new_n656 = new_n655 ^ new_n651;
  assign new_n657 = ~new_n656 & new_n649;
  assign new_n658 = new_n657 ^ n75;
  assign new_n659 = new_n658 ^ new_n654;
  assign new_n660 = n205 ^ n77;
  assign new_n661 = new_n658 ^ n204;
  assign new_n662 = ~new_n661 & new_n654;
  assign new_n663 = new_n662 ^ n76;
  assign new_n664 = new_n663 ^ new_n660;
  assign new_n665 = n206 ^ n78;
  assign new_n666 = n205 ^ n76;
  assign new_n667 = new_n666 ^ new_n662;
  assign new_n668 = ~new_n667 & new_n660;
  assign new_n669 = new_n668 ^ n77;
  assign new_n670 = new_n669 ^ new_n665;
  assign new_n671 = n207 ^ n79;
  assign new_n672 = new_n669 ^ n206;
  assign new_n673 = ~new_n672 & new_n665;
  assign new_n674 = new_n673 ^ n78;
  assign new_n675 = new_n674 ^ new_n671;
  assign new_n676 = n208 ^ n80;
  assign new_n677 = n207 ^ n78;
  assign new_n678 = new_n677 ^ new_n673;
  assign new_n679 = ~new_n678 & new_n671;
  assign new_n680 = new_n679 ^ n79;
  assign new_n681 = new_n680 ^ new_n676;
  assign new_n682 = new_n680 ^ n208;
  assign new_n683 = ~new_n682 & new_n676;
  assign new_n684 = new_n683 ^ n80;
  assign new_n685 = n209 ^ n81;
  assign new_n686 = new_n685 ^ new_n684;
  assign new_n687 = n210 ^ n82;
  assign new_n688 = new_n684 ^ n209;
  assign new_n689 = ~new_n688 & new_n685;
  assign new_n690 = new_n689 ^ n81;
  assign new_n691 = new_n690 ^ new_n687;
  assign new_n692 = n211 ^ n83;
  assign new_n693 = new_n690 ^ n210;
  assign new_n694 = ~new_n693 & new_n687;
  assign new_n695 = new_n694 ^ n82;
  assign new_n696 = new_n695 ^ new_n692;
  assign new_n697 = n212 ^ n84;
  assign new_n698 = n211 ^ n82;
  assign new_n699 = new_n698 ^ new_n694;
  assign new_n700 = ~new_n699 & new_n692;
  assign new_n701 = new_n700 ^ n83;
  assign new_n702 = new_n701 ^ new_n697;
  assign new_n703 = n213 ^ n85;
  assign new_n704 = new_n701 ^ n212;
  assign new_n705 = ~new_n704 & new_n697;
  assign new_n706 = new_n705 ^ n84;
  assign new_n707 = new_n706 ^ new_n703;
  assign new_n708 = n214 ^ n86;
  assign new_n709 = n213 ^ n84;
  assign new_n710 = new_n709 ^ new_n705;
  assign new_n711 = ~new_n710 & new_n703;
  assign new_n712 = new_n711 ^ n85;
  assign new_n713 = new_n712 ^ new_n708;
  assign new_n714 = n215 ^ n87;
  assign new_n715 = new_n712 ^ n214;
  assign new_n716 = ~new_n715 & new_n708;
  assign new_n717 = new_n716 ^ n86;
  assign new_n718 = new_n717 ^ new_n714;
  assign new_n719 = n216 ^ n88;
  assign new_n720 = n215 ^ n86;
  assign new_n721 = new_n720 ^ new_n716;
  assign new_n722 = ~new_n721 & new_n714;
  assign new_n723 = new_n722 ^ n87;
  assign new_n724 = new_n723 ^ new_n719;
  assign new_n725 = n217 ^ n89;
  assign new_n726 = new_n723 ^ n216;
  assign new_n727 = ~new_n726 & new_n719;
  assign new_n728 = new_n727 ^ n88;
  assign new_n729 = new_n728 ^ new_n725;
  assign new_n730 = n218 ^ n90;
  assign new_n731 = n217 ^ n88;
  assign new_n732 = new_n731 ^ new_n727;
  assign new_n733 = ~new_n732 & new_n725;
  assign new_n734 = new_n733 ^ n89;
  assign new_n735 = new_n734 ^ new_n730;
  assign new_n736 = new_n734 ^ n218;
  assign new_n737 = ~new_n736 & new_n730;
  assign new_n738 = new_n737 ^ n90;
  assign new_n739 = n219 ^ n91;
  assign new_n740 = new_n739 ^ new_n738;
  assign new_n741 = n220 ^ n92;
  assign new_n742 = new_n738 ^ n219;
  assign new_n743 = ~new_n742 & new_n739;
  assign new_n744 = new_n743 ^ n91;
  assign new_n745 = new_n744 ^ new_n741;
  assign new_n746 = new_n744 ^ n220;
  assign new_n747 = ~new_n746 & new_n741;
  assign new_n748 = new_n747 ^ n92;
  assign new_n749 = n221 ^ n93;
  assign new_n750 = new_n749 ^ new_n748;
  assign new_n751 = n222 ^ n94;
  assign new_n752 = new_n748 ^ n221;
  assign new_n753 = ~new_n752 & new_n749;
  assign new_n754 = new_n753 ^ n93;
  assign new_n755 = new_n754 ^ new_n751;
  assign new_n756 = n223 ^ n95;
  assign new_n757 = new_n754 ^ n222;
  assign new_n758 = ~new_n757 & new_n751;
  assign new_n759 = new_n758 ^ n94;
  assign new_n760 = new_n759 ^ new_n756;
  assign new_n761 = n224 ^ n96;
  assign new_n762 = new_n759 ^ n223;
  assign new_n763 = ~new_n762 & new_n756;
  assign new_n764 = new_n763 ^ n95;
  assign new_n765 = new_n764 ^ new_n761;
  assign new_n766 = n225 ^ n97;
  assign new_n767 = new_n764 ^ n224;
  assign new_n768 = ~new_n767 & new_n761;
  assign new_n769 = new_n768 ^ n96;
  assign new_n770 = new_n769 ^ new_n766;
  assign new_n771 = n226 ^ n98;
  assign new_n772 = new_n769 ^ n225;
  assign new_n773 = ~new_n772 & new_n766;
  assign new_n774 = new_n773 ^ n97;
  assign new_n775 = new_n774 ^ new_n771;
  assign new_n776 = n227 ^ n99;
  assign new_n777 = new_n774 ^ n226;
  assign new_n778 = ~new_n777 & new_n771;
  assign new_n779 = new_n778 ^ n98;
  assign new_n780 = new_n779 ^ new_n776;
  assign new_n781 = n228 ^ n100;
  assign new_n782 = n227 ^ n98;
  assign new_n783 = new_n782 ^ new_n778;
  assign new_n784 = ~new_n783 & new_n776;
  assign new_n785 = new_n784 ^ n99;
  assign new_n786 = new_n785 ^ new_n781;
  assign new_n787 = n229 ^ n101;
  assign new_n788 = new_n785 ^ n228;
  assign new_n789 = ~new_n788 & new_n781;
  assign new_n790 = new_n789 ^ n100;
  assign new_n791 = new_n790 ^ new_n787;
  assign new_n792 = n230 ^ n102;
  assign new_n793 = n229 ^ n100;
  assign new_n794 = new_n793 ^ new_n789;
  assign new_n795 = ~new_n794 & new_n787;
  assign new_n796 = new_n795 ^ n101;
  assign new_n797 = new_n796 ^ new_n792;
  assign new_n798 = n231 ^ n103;
  assign new_n799 = new_n796 ^ n230;
  assign new_n800 = ~new_n799 & new_n792;
  assign new_n801 = new_n800 ^ n102;
  assign new_n802 = new_n801 ^ new_n798;
  assign new_n803 = n232 ^ n104;
  assign new_n804 = n231 ^ n102;
  assign new_n805 = new_n804 ^ new_n800;
  assign new_n806 = ~new_n805 & new_n798;
  assign new_n807 = new_n806 ^ n103;
  assign new_n808 = new_n807 ^ new_n803;
  assign new_n809 = n233 ^ n105;
  assign new_n810 = new_n807 ^ n232;
  assign new_n811 = ~new_n810 & new_n803;
  assign new_n812 = new_n811 ^ n104;
  assign new_n813 = new_n812 ^ new_n809;
  assign new_n814 = n234 ^ n106;
  assign new_n815 = new_n812 ^ n233;
  assign new_n816 = ~new_n815 & new_n809;
  assign new_n817 = new_n816 ^ n105;
  assign new_n818 = new_n817 ^ new_n814;
  assign new_n819 = n235 ^ n107;
  assign new_n820 = new_n817 ^ n234;
  assign new_n821 = ~new_n820 & new_n814;
  assign new_n822 = new_n821 ^ n106;
  assign new_n823 = new_n822 ^ new_n819;
  assign new_n824 = n236 ^ n108;
  assign new_n825 = n235 ^ n106;
  assign new_n826 = new_n825 ^ new_n821;
  assign new_n827 = ~new_n826 & new_n819;
  assign new_n828 = new_n827 ^ n107;
  assign new_n829 = new_n828 ^ new_n824;
  assign new_n830 = n237 ^ n109;
  assign new_n831 = new_n828 ^ n236;
  assign new_n832 = ~new_n831 & new_n824;
  assign new_n833 = new_n832 ^ n108;
  assign new_n834 = new_n833 ^ new_n830;
  assign new_n835 = n238 ^ n110;
  assign new_n836 = new_n833 ^ n237;
  assign new_n837 = ~new_n836 & new_n830;
  assign new_n838 = new_n837 ^ n109;
  assign new_n839 = new_n838 ^ new_n835;
  assign new_n840 = n239 ^ n111;
  assign new_n841 = new_n838 ^ n238;
  assign new_n842 = ~new_n841 & new_n835;
  assign new_n843 = new_n842 ^ n110;
  assign new_n844 = new_n843 ^ new_n840;
  assign new_n845 = n240 ^ n112;
  assign new_n846 = n239 ^ n110;
  assign new_n847 = new_n846 ^ new_n842;
  assign new_n848 = ~new_n847 & new_n840;
  assign new_n849 = new_n848 ^ n111;
  assign new_n850 = new_n849 ^ new_n845;
  assign new_n851 = n241 ^ n113;
  assign new_n852 = new_n849 ^ n240;
  assign new_n853 = ~new_n852 & new_n845;
  assign new_n854 = new_n853 ^ n112;
  assign new_n855 = new_n854 ^ new_n851;
  assign new_n856 = n242 ^ n114;
  assign new_n857 = new_n854 ^ n241;
  assign new_n858 = ~new_n857 & new_n851;
  assign new_n859 = new_n858 ^ n113;
  assign new_n860 = new_n859 ^ new_n856;
  assign new_n861 = n243 ^ n115;
  assign new_n862 = new_n859 ^ n242;
  assign new_n863 = ~new_n862 & new_n856;
  assign new_n864 = new_n863 ^ n114;
  assign new_n865 = new_n864 ^ new_n861;
  assign new_n866 = n244 ^ n116;
  assign new_n867 = new_n864 ^ n243;
  assign new_n868 = ~new_n867 & new_n861;
  assign new_n869 = new_n868 ^ n115;
  assign new_n870 = new_n869 ^ new_n866;
  assign new_n871 = n245 ^ n117;
  assign new_n872 = new_n869 ^ n244;
  assign new_n873 = ~new_n872 & new_n866;
  assign new_n874 = new_n873 ^ n116;
  assign new_n875 = new_n874 ^ new_n871;
  assign new_n876 = n246 ^ n118;
  assign new_n877 = new_n874 ^ n245;
  assign new_n878 = ~new_n877 & new_n871;
  assign new_n879 = new_n878 ^ n117;
  assign new_n880 = new_n879 ^ new_n876;
  assign new_n881 = n247 ^ n119;
  assign new_n882 = new_n879 ^ n246;
  assign new_n883 = ~new_n882 & new_n876;
  assign new_n884 = new_n883 ^ n118;
  assign new_n885 = new_n884 ^ new_n881;
  assign new_n886 = n248 ^ n120;
  assign new_n887 = new_n884 ^ n247;
  assign new_n888 = ~new_n887 & new_n881;
  assign new_n889 = new_n888 ^ n119;
  assign new_n890 = new_n889 ^ new_n886;
  assign new_n891 = n249 ^ n121;
  assign new_n892 = new_n889 ^ n248;
  assign new_n893 = ~new_n892 & new_n886;
  assign new_n894 = new_n893 ^ n120;
  assign new_n895 = new_n894 ^ new_n891;
  assign new_n896 = n250 ^ n122;
  assign new_n897 = new_n894 ^ n249;
  assign new_n898 = ~new_n897 & new_n891;
  assign new_n899 = new_n898 ^ n121;
  assign new_n900 = new_n899 ^ new_n896;
  assign new_n901 = n251 ^ n123;
  assign new_n902 = new_n899 ^ n250;
  assign new_n903 = ~new_n902 & new_n896;
  assign new_n904 = new_n903 ^ n122;
  assign new_n905 = new_n904 ^ new_n901;
  assign new_n906 = n252 ^ n124;
  assign new_n907 = new_n904 ^ n251;
  assign new_n908 = ~new_n907 & new_n901;
  assign new_n909 = new_n908 ^ n123;
  assign new_n910 = new_n909 ^ new_n906;
  assign new_n911 = n253 ^ n125;
  assign new_n912 = new_n909 ^ n252;
  assign new_n913 = ~new_n912 & new_n906;
  assign new_n914 = new_n913 ^ n124;
  assign new_n915 = new_n914 ^ new_n911;
  assign new_n916 = n254 ^ n126;
  assign new_n917 = new_n914 ^ n253;
  assign new_n918 = ~new_n917 & new_n911;
  assign new_n919 = new_n918 ^ n125;
  assign new_n920 = new_n919 ^ new_n916;
  assign new_n921 = n255 ^ n127;
  assign new_n922 = new_n919 ^ n254;
  assign new_n923 = ~new_n922 & new_n916;
  assign new_n924 = new_n923 ^ n126;
  assign new_n925 = new_n924 ^ new_n921;
  assign new_n926 = n256 ^ n128;
  assign new_n927 = new_n924 ^ n255;
  assign new_n928 = ~new_n927 & new_n921;
  assign new_n929 = new_n928 ^ n127;
  assign new_n930 = new_n929 ^ new_n926;
  assign new_n931 = new_n929 ^ n256;
  assign new_n932 = ~new_n931 & new_n926;
  assign new_n933 = new_n932 ^ n128;
  assign po0 = new_n257;
  assign po1 = new_n260;
  assign po2 = new_n265;
  assign po3 = new_n270;
  assign po4 = new_n275;
  assign po5 = new_n281;
  assign po6 = new_n286;
  assign po7 = new_n292;
  assign po8 = new_n297;
  assign po9 = new_n303;
  assign po10 = new_n308;
  assign po11 = new_n313;
  assign po12 = new_n318;
  assign po13 = new_n324;
  assign po14 = new_n329;
  assign po15 = new_n335;
  assign po16 = new_n340;
  assign po17 = new_n346;
  assign po18 = new_n351;
  assign po19 = new_n357;
  assign po20 = new_n362;
  assign po21 = new_n367;
  assign po22 = new_n372;
  assign po23 = new_n378;
  assign po24 = new_n383;
  assign po25 = new_n389;
  assign po26 = new_n394;
  assign po27 = new_n400;
  assign po28 = new_n405;
  assign po29 = new_n411;
  assign po30 = new_n416;
  assign po31 = new_n421;
  assign po32 = new_n426;
  assign po33 = new_n432;
  assign po34 = new_n437;
  assign po35 = new_n443;
  assign po36 = new_n448;
  assign po37 = new_n454;
  assign po38 = new_n459;
  assign po39 = new_n465;
  assign po40 = new_n470;
  assign po41 = new_n475;
  assign po42 = new_n480;
  assign po43 = new_n486;
  assign po44 = new_n491;
  assign po45 = new_n497;
  assign po46 = new_n502;
  assign po47 = new_n508;
  assign po48 = new_n513;
  assign po49 = new_n519;
  assign po50 = new_n524;
  assign po51 = new_n529;
  assign po52 = new_n534;
  assign po53 = new_n540;
  assign po54 = new_n545;
  assign po55 = new_n551;
  assign po56 = new_n556;
  assign po57 = new_n562;
  assign po58 = new_n567;
  assign po59 = new_n573;
  assign po60 = new_n578;
  assign po61 = new_n583;
  assign po62 = new_n588;
  assign po63 = new_n594;
  assign po64 = new_n599;
  assign po65 = new_n605;
  assign po66 = new_n610;
  assign po67 = new_n616;
  assign po68 = new_n621;
  assign po69 = new_n627;
  assign po70 = new_n632;
  assign po71 = new_n637;
  assign po72 = new_n642;
  assign po73 = new_n648;
  assign po74 = new_n653;
  assign po75 = new_n659;
  assign po76 = new_n664;
  assign po77 = new_n670;
  assign po78 = new_n675;
  assign po79 = new_n681;
  assign po80 = new_n686;
  assign po81 = new_n691;
  assign po82 = new_n696;
  assign po83 = new_n702;
  assign po84 = new_n707;
  assign po85 = new_n713;
  assign po86 = new_n718;
  assign po87 = new_n724;
  assign po88 = new_n729;
  assign po89 = new_n735;
  assign po90 = new_n740;
  assign po91 = new_n745;
  assign po92 = new_n750;
  assign po93 = new_n755;
  assign po94 = new_n760;
  assign po95 = new_n765;
  assign po96 = new_n770;
  assign po97 = new_n775;
  assign po98 = new_n780;
  assign po99 = new_n786;
  assign po100 = new_n791;
  assign po101 = new_n797;
  assign po102 = new_n802;
  assign po103 = new_n808;
  assign po104 = new_n813;
  assign po105 = new_n818;
  assign po106 = new_n823;
  assign po107 = new_n829;
  assign po108 = new_n834;
  assign po109 = new_n839;
  assign po110 = new_n844;
  assign po111 = new_n850;
  assign po112 = new_n855;
  assign po113 = new_n860;
  assign po114 = new_n865;
  assign po115 = new_n870;
  assign po116 = new_n875;
  assign po117 = new_n880;
  assign po118 = new_n885;
  assign po119 = new_n890;
  assign po120 = new_n895;
  assign po121 = new_n900;
  assign po122 = new_n905;
  assign po123 = new_n910;
  assign po124 = new_n915;
  assign po125 = new_n920;
  assign po126 = new_n925;
  assign po127 = new_n930;
  assign po128 = new_n933;
endmodule


