module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 ;
  assign n150 = x3 ^ x2 ;
  assign n136 = x10 ^ x8 ;
  assign n135 = x9 ^ x8 ;
  assign n137 = n136 ^ n135 ;
  assign n138 = n137 ^ x10 ;
  assign n139 = n138 ^ x7 ;
  assign n143 = ~x2 & ~n139 ;
  assign n141 = ~n136 & ~n139 ;
  assign n140 = x3 & ~n139 ;
  assign n142 = n141 ^ n140 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = n144 ^ x3 ;
  assign n146 = n145 ^ x2 ;
  assign n147 = n146 ^ n137 ;
  assign n148 = n137 & ~n147 ;
  assign n149 = n148 ^ n144 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = n151 ^ x9 ;
  assign n157 = x10 ^ x7 ;
  assign n158 = n157 ^ n136 ;
  assign n156 = n150 ^ n135 ;
  assign n159 = n158 ^ n156 ;
  assign n160 = x10 & n159 ;
  assign n161 = ~n152 & n160 ;
  assign n154 = ~n144 & ~n152 ;
  assign n153 = ~n148 & ~n152 ;
  assign n155 = n154 ^ n153 ;
  assign n162 = n161 ^ n155 ;
  assign n163 = n162 ^ n157 ;
  assign n164 = n163 ^ x10 ;
  assign n165 = n164 ^ n157 ;
  assign n199 = x6 & x10 ;
  assign n200 = ~n165 & n199 ;
  assign n69 = ~x6 & ~x7 ;
  assign n197 = x10 & n69 ;
  assign n64 = x4 & x5 ;
  assign n81 = n64 ^ x4 ;
  assign n82 = x8 & n81 ;
  assign n73 = x1 & x4 ;
  assign n70 = x8 ^ x1 ;
  assign n71 = x4 & n70 ;
  assign n72 = n71 ^ x8 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ x0 ;
  assign n76 = x0 & n75 ;
  assign n77 = n76 ^ n75 ;
  assign n78 = n77 ^ n72 ;
  assign n79 = n78 ^ x0 ;
  assign n80 = n69 & n79 ;
  assign n110 = n82 ^ n80 ;
  assign n111 = n110 ^ x5 ;
  assign n114 = x5 & n111 ;
  assign n115 = n114 ^ x5 ;
  assign n116 = n115 ^ n111 ;
  assign n112 = n82 & n111 ;
  assign n113 = n112 ^ n82 ;
  assign n117 = n116 ^ n113 ;
  assign n107 = ~x4 & x5 ;
  assign n108 = x8 & n107 ;
  assign n109 = n108 ^ x5 ;
  assign n118 = n117 ^ n109 ;
  assign n54 = x3 & ~x8 ;
  assign n190 = ~x9 & n54 ;
  assign n191 = ~n118 & n190 ;
  assign n55 = x2 & x7 ;
  assign n56 = n55 ^ x2 ;
  assign n57 = n56 ^ x7 ;
  assign n58 = x1 & x5 ;
  assign n59 = n57 & n58 ;
  assign n60 = n59 ^ n58 ;
  assign n23 = x4 & x7 ;
  assign n24 = n23 ^ x7 ;
  assign n61 = n60 ^ n24 ;
  assign n166 = x6 & ~x10 ;
  assign n172 = ~n165 & n166 ;
  assign n173 = n172 ^ n166 ;
  assign n192 = n61 & n173 ;
  assign n193 = n191 & n192 ;
  assign n185 = x9 & ~n118 ;
  assign n186 = n185 ^ n118 ;
  assign n50 = x7 & ~x8 ;
  assign n28 = x3 & x4 ;
  assign n104 = n28 ^ x4 ;
  assign n105 = n50 & n104 ;
  assign n187 = ~n105 & n173 ;
  assign n188 = ~n186 & n187 ;
  assign n189 = n188 ^ n173 ;
  assign n194 = n193 ^ n189 ;
  assign n12 = x7 & x8 ;
  assign n13 = n12 ^ x7 ;
  assign n14 = n13 ^ x8 ;
  assign n19 = x2 & n14 ;
  assign n20 = n19 ^ x2 ;
  assign n21 = n20 ^ n14 ;
  assign n15 = x1 & x2 ;
  assign n16 = n14 & n15 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n17 ^ n15 ;
  assign n22 = n21 ^ n18 ;
  assign n40 = x9 & n22 ;
  assign n41 = n40 ^ x9 ;
  assign n42 = n41 ^ n22 ;
  assign n35 = x1 & ~x2 ;
  assign n36 = ~x9 & n35 ;
  assign n37 = ~n24 & ~n28 ;
  assign n38 = n36 & n37 ;
  assign n25 = ~x9 & ~n24 ;
  assign n26 = ~n22 & n25 ;
  assign n27 = n15 ^ x1 ;
  assign n29 = x4 & x8 ;
  assign n30 = n28 & n29 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n27 & ~n31 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n26 & n33 ;
  assign n39 = n38 ^ n34 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = x5 & ~x6 ;
  assign n45 = ~x5 & x6 ;
  assign n46 = x9 & ~n45 ;
  assign n47 = n44 & n46 ;
  assign n180 = n43 & n47 ;
  assign n181 = n173 & n180 ;
  assign n96 = ~x9 & n44 ;
  assign n169 = n43 & n96 ;
  assign n170 = n169 ^ n96 ;
  assign n171 = n170 ^ n96 ;
  assign n90 = n82 ^ x5 ;
  assign n52 = ~x4 & n50 ;
  assign n51 = ~n28 & n50 ;
  assign n53 = n52 ^ n51 ;
  assign n86 = x5 & n53 ;
  assign n84 = x5 & n54 ;
  assign n85 = n61 & n84 ;
  assign n87 = n86 ^ n85 ;
  assign n62 = n54 & n61 ;
  assign n63 = n62 ^ n53 ;
  assign n88 = n87 ^ n63 ;
  assign n83 = n53 & n82 ;
  assign n89 = n88 ^ n83 ;
  assign n91 = n90 ^ n89 ;
  assign n92 = n80 & ~n91 ;
  assign n93 = n92 ^ n91 ;
  assign n176 = ~n93 & n173 ;
  assign n177 = n176 ^ n173 ;
  assign n178 = n171 & n177 ;
  assign n65 = n64 ^ x5 ;
  assign n66 = x8 & n65 ;
  assign n67 = x5 & ~n66 ;
  assign n68 = ~n63 & n67 ;
  assign n174 = ~n68 & n173 ;
  assign n175 = n171 & n174 ;
  assign n179 = n178 ^ n175 ;
  assign n182 = n181 ^ n179 ;
  assign n183 = n182 ^ n173 ;
  assign n167 = n46 & n166 ;
  assign n168 = n165 & n167 ;
  assign n184 = n183 ^ n168 ;
  assign n195 = n194 ^ n184 ;
  assign n125 = ~x9 & n61 ;
  assign n126 = n54 & n125 ;
  assign n127 = ~n118 & n126 ;
  assign n119 = n118 ^ n105 ;
  assign n120 = x9 & n105 ;
  assign n121 = n120 ^ n118 ;
  assign n122 = n121 ^ x9 ;
  assign n123 = n119 & n122 ;
  assign n124 = n123 ^ n120 ;
  assign n128 = n127 ^ n124 ;
  assign n106 = n105 ^ x9 ;
  assign n129 = n128 ^ n106 ;
  assign n130 = n129 ^ n46 ;
  assign n131 = x10 & ~n130 ;
  assign n132 = n131 ^ n130 ;
  assign n94 = n93 ^ n68 ;
  assign n95 = n94 ^ n43 ;
  assign n97 = ~x10 & n96 ;
  assign n98 = n97 ^ n43 ;
  assign n99 = ~n97 & n98 ;
  assign n100 = n99 ^ n43 ;
  assign n101 = ~n95 & ~n100 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = n102 ^ n94 ;
  assign n133 = n132 ^ n103 ;
  assign n48 = ~x10 & n47 ;
  assign n49 = n43 & n48 ;
  assign n134 = n133 ^ n49 ;
  assign n196 = n195 ^ n134 ;
  assign n198 = n197 ^ n196 ;
  assign n201 = n200 ^ n198 ;
  assign n244 = n29 ^ x8 ;
  assign n245 = n244 ^ x7 ;
  assign n251 = x9 & ~n245 ;
  assign n252 = n251 ^ n244 ;
  assign n351 = n252 ^ x6 ;
  assign n352 = ~x5 & ~x10 ;
  assign n353 = n352 ^ x6 ;
  assign n354 = ~x6 & ~n353 ;
  assign n355 = n354 ^ n252 ;
  assign n356 = ~n351 & n355 ;
  assign n357 = n356 ^ n354 ;
  assign n358 = n357 ^ n352 ;
  assign n359 = n358 ^ n252 ;
  assign n259 = x8 & x9 ;
  assign n260 = n259 ^ x8 ;
  assign n261 = n260 ^ x9 ;
  assign n360 = x7 & ~n261 ;
  assign n361 = x7 & x9 ;
  assign n362 = n361 ^ x9 ;
  assign n363 = ~n28 & ~n362 ;
  assign n364 = n360 & n363 ;
  assign n365 = n364 ^ n362 ;
  assign n372 = n365 ^ n359 ;
  assign n373 = n359 & n372 ;
  assign n374 = n373 ^ n359 ;
  assign n375 = n374 ^ n372 ;
  assign n313 = x4 & x9 ;
  assign n314 = n313 ^ x4 ;
  assign n315 = n314 ^ x9 ;
  assign n316 = n57 & n315 ;
  assign n317 = n316 ^ n57 ;
  assign n318 = n317 ^ n315 ;
  assign n319 = n318 ^ n57 ;
  assign n320 = n319 ^ n315 ;
  assign n325 = n320 ^ x1 ;
  assign n326 = ~n320 & ~n325 ;
  assign n327 = n326 ^ n320 ;
  assign n328 = n327 ^ n325 ;
  assign n321 = n260 ^ x1 ;
  assign n322 = ~x1 & n321 ;
  assign n323 = ~n320 & n322 ;
  assign n324 = n323 ^ n321 ;
  assign n329 = n328 ^ n324 ;
  assign n330 = n329 ^ n260 ;
  assign n331 = n330 ^ n260 ;
  assign n305 = n23 ^ x4 ;
  assign n306 = x0 & x2 ;
  assign n307 = n306 ^ x2 ;
  assign n308 = ~n305 & ~n307 ;
  assign n343 = n308 ^ n305 ;
  assign n344 = n343 ^ n307 ;
  assign n345 = n344 ^ n305 ;
  assign n346 = ~x6 & n345 ;
  assign n347 = ~n331 & n346 ;
  assign n348 = n347 ^ n346 ;
  assign n309 = n308 ^ n307 ;
  assign n332 = x0 & x6 ;
  assign n333 = n332 ^ x0 ;
  assign n334 = n15 & ~n333 ;
  assign n335 = n334 ^ n15 ;
  assign n336 = n335 ^ n333 ;
  assign n337 = n309 & ~n336 ;
  assign n338 = n337 ^ n309 ;
  assign n339 = n338 ^ n336 ;
  assign n340 = ~n331 & n339 ;
  assign n341 = n340 ^ n339 ;
  assign n310 = x6 & n309 ;
  assign n311 = n310 ^ x6 ;
  assign n312 = n311 ^ n309 ;
  assign n342 = n341 ^ n312 ;
  assign n349 = n348 ^ n342 ;
  assign n350 = n349 ^ n339 ;
  assign n366 = n359 & ~n365 ;
  assign n367 = n366 ^ n350 ;
  assign n368 = n350 & n367 ;
  assign n369 = n368 ^ n350 ;
  assign n370 = n369 ^ n350 ;
  assign n371 = n370 ^ n367 ;
  assign n376 = n375 ^ n371 ;
  assign n377 = n376 ^ n365 ;
  assign n243 = x5 & ~x10 ;
  assign n248 = x6 & ~n244 ;
  assign n246 = x6 & x9 ;
  assign n247 = ~n245 & n246 ;
  assign n249 = n248 ^ n247 ;
  assign n250 = n249 ^ x6 ;
  assign n253 = n252 ^ n250 ;
  assign n300 = n253 ^ n243 ;
  assign n301 = ~n243 & ~n300 ;
  assign n254 = n243 & ~n253 ;
  assign n270 = x7 ^ x4 ;
  assign n271 = x9 & n270 ;
  assign n272 = n271 ^ n270 ;
  assign n273 = n272 ^ x7 ;
  assign n293 = ~x3 & x6 ;
  assign n294 = n261 & n293 ;
  assign n295 = n273 & n294 ;
  assign n269 = x3 & x6 ;
  assign n277 = n261 & n269 ;
  assign n289 = n273 & n277 ;
  assign n284 = ~n261 & n269 ;
  assign n285 = n269 & ~n284 ;
  assign n286 = ~n269 & n284 ;
  assign n287 = ~n285 & ~n286 ;
  assign n262 = x4 & ~n261 ;
  assign n256 = x7 & n15 ;
  assign n263 = n256 ^ x7 ;
  assign n264 = n263 ^ n15 ;
  assign n265 = n262 & ~n264 ;
  assign n266 = n265 ^ n262 ;
  assign n255 = ~x4 & ~x6 ;
  assign n257 = n256 ^ n15 ;
  assign n258 = n255 & n257 ;
  assign n267 = n266 ^ n258 ;
  assign n281 = n273 ^ n267 ;
  assign n282 = ~n267 & n281 ;
  assign n279 = ~n267 & n273 ;
  assign n274 = n261 & n273 ;
  assign n275 = n269 & n274 ;
  assign n276 = n267 & n275 ;
  assign n278 = n277 ^ n276 ;
  assign n280 = n279 ^ n278 ;
  assign n283 = n282 ^ n280 ;
  assign n288 = n287 ^ n283 ;
  assign n290 = n289 ^ n288 ;
  assign n268 = x3 & ~n267 ;
  assign n291 = n290 ^ n268 ;
  assign n292 = n291 ^ x3 ;
  assign n296 = n295 ^ n292 ;
  assign n297 = n296 ^ n253 ;
  assign n298 = n254 & ~n297 ;
  assign n299 = n298 ^ n297 ;
  assign n302 = n301 ^ n299 ;
  assign n303 = n302 ^ n296 ;
  assign n304 = n303 ^ x10 ;
  assign n378 = n377 ^ n304 ;
  assign n202 = x8 & x10 ;
  assign n203 = x6 & x7 ;
  assign n204 = ~x9 & n203 ;
  assign n205 = n202 & n204 ;
  assign n206 = ~x8 & ~n203 ;
  assign n212 = ~x7 & ~x10 ;
  assign n213 = n206 & n212 ;
  assign n214 = ~n205 & n213 ;
  assign n207 = x10 & n206 ;
  assign n380 = n213 ^ n207 ;
  assign n381 = n205 & n380 ;
  assign n382 = n381 ^ n205 ;
  assign n383 = n382 ^ n380 ;
  assign n227 = x6 & ~x9 ;
  assign n228 = x2 & n28 ;
  assign n229 = n227 & n228 ;
  assign n219 = x3 & x5 ;
  assign n220 = n219 ^ x5 ;
  assign n221 = x6 & n220 ;
  assign n222 = n221 ^ n220 ;
  assign n215 = x4 & x6 ;
  assign n216 = n215 ^ x6 ;
  assign n217 = x9 & n216 ;
  assign n218 = n217 ^ n216 ;
  assign n223 = n222 ^ n218 ;
  assign n224 = x2 & ~n223 ;
  assign n225 = n224 ^ x2 ;
  assign n226 = n225 ^ n223 ;
  assign n230 = n229 ^ n226 ;
  assign n231 = ~x4 & n227 ;
  assign n236 = ~x3 & n231 ;
  assign n237 = ~n230 & n236 ;
  assign n238 = n237 ^ n230 ;
  assign n232 = ~x1 & ~x3 ;
  assign n233 = n44 & n232 ;
  assign n234 = ~n231 & n233 ;
  assign n235 = ~n230 & n234 ;
  assign n239 = n238 ^ n235 ;
  assign n384 = n383 ^ n239 ;
  assign n208 = ~n205 & n207 ;
  assign n379 = n208 ^ n205 ;
  assign n385 = n384 ^ n379 ;
  assign n386 = n214 & ~n385 ;
  assign n387 = n386 ^ n379 ;
  assign n388 = n378 & n387 ;
  assign n389 = n388 ^ n378 ;
  assign n390 = n389 ^ n387 ;
  assign n391 = n390 ^ n387 ;
  assign n240 = n214 & ~n239 ;
  assign n209 = n205 & ~n208 ;
  assign n210 = ~n205 & n208 ;
  assign n211 = ~n209 & ~n210 ;
  assign n241 = n240 ^ n211 ;
  assign n242 = n241 ^ n214 ;
  assign n392 = n391 ^ n242 ;
  assign n474 = x5 & x7 ;
  assign n475 = x8 & ~x10 ;
  assign n476 = ~n474 & n475 ;
  assign n477 = n476 ^ x10 ;
  assign n478 = x9 & ~n477 ;
  assign n479 = n478 ^ x9 ;
  assign n493 = n203 ^ x6 ;
  assign n494 = n64 & n493 ;
  assign n495 = n494 ^ n493 ;
  assign n496 = n495 ^ x6 ;
  assign n497 = n496 ^ x7 ;
  assign n519 = x9 & ~x10 ;
  assign n520 = x8 & n519 ;
  assign n521 = n497 & n520 ;
  assign n522 = n521 ^ n519 ;
  assign n523 = n522 ^ x10 ;
  assign n526 = x5 & x8 ;
  assign n527 = n526 ^ x5 ;
  assign n528 = x9 & n527 ;
  assign n529 = ~n202 & n203 ;
  assign n530 = ~n528 & n529 ;
  assign n531 = n523 & n530 ;
  assign n532 = ~n479 & n531 ;
  assign n524 = ~n203 & n523 ;
  assign n525 = ~n479 & n524 ;
  assign n533 = n532 ^ n525 ;
  assign n431 = x5 & x6 ;
  assign n450 = ~x8 & ~n28 ;
  assign n451 = n431 & n450 ;
  assign n452 = n451 ^ x8 ;
  assign n396 = x2 & x5 ;
  assign n397 = n396 ^ x2 ;
  assign n398 = x6 & n397 ;
  assign n393 = n58 ^ x5 ;
  assign n394 = x6 & n393 ;
  assign n395 = n394 ^ n393 ;
  assign n399 = n398 ^ n395 ;
  assign n402 = ~n28 & n399 ;
  assign n400 = x8 & n28 ;
  assign n401 = n399 & ~n400 ;
  assign n403 = n402 ^ n401 ;
  assign n453 = n452 ^ n403 ;
  assign n460 = ~n220 & n305 ;
  assign n461 = ~n453 & n460 ;
  assign n454 = x2 & x3 ;
  assign n455 = n454 ^ x3 ;
  assign n456 = x6 & n455 ;
  assign n457 = n456 ^ n455 ;
  assign n458 = n305 & ~n457 ;
  assign n459 = ~n453 & n458 ;
  assign n462 = n461 ^ n459 ;
  assign n412 = x0 & x1 ;
  assign n413 = n28 & n412 ;
  assign n414 = n413 ^ n28 ;
  assign n415 = n414 ^ n255 ;
  assign n468 = n397 & n415 ;
  assign n469 = n462 & n468 ;
  assign n407 = x3 & ~n65 ;
  assign n408 = n407 ^ x3 ;
  assign n404 = ~n104 & ~n333 ;
  assign n405 = n404 ^ n104 ;
  assign n406 = n405 ^ n333 ;
  assign n409 = n408 ^ n406 ;
  assign n463 = ~x5 & n15 ;
  assign n464 = n415 & n463 ;
  assign n465 = n464 ^ n15 ;
  assign n466 = ~n409 & n465 ;
  assign n467 = n462 & n466 ;
  assign n470 = n469 ^ n467 ;
  assign n440 = n28 & ~n400 ;
  assign n441 = ~n28 & n400 ;
  assign n442 = ~n440 & ~n441 ;
  assign n432 = n400 ^ x8 ;
  assign n433 = n432 ^ n28 ;
  assign n434 = n431 & ~n433 ;
  assign n435 = n434 ^ n433 ;
  assign n448 = n442 ^ n435 ;
  assign n422 = n415 ^ x7 ;
  assign n423 = n397 ^ x7 ;
  assign n424 = ~n397 & ~n423 ;
  assign n425 = n424 ^ x7 ;
  assign n426 = ~n422 & n425 ;
  assign n427 = n426 ^ n424 ;
  assign n410 = n257 & n409 ;
  assign n411 = n410 ^ n257 ;
  assign n418 = n411 & n415 ;
  assign n419 = n418 ^ n415 ;
  assign n420 = n419 ^ n411 ;
  assign n416 = x5 & n415 ;
  assign n417 = n411 & n416 ;
  assign n421 = n420 ^ n417 ;
  assign n428 = n427 ^ n421 ;
  assign n443 = ~n428 & n442 ;
  assign n444 = n443 ^ n442 ;
  assign n445 = n444 ^ n428 ;
  assign n436 = ~n428 & n435 ;
  assign n437 = n436 ^ n435 ;
  assign n438 = n437 ^ n428 ;
  assign n429 = n403 & ~n428 ;
  assign n430 = n429 ^ n403 ;
  assign n439 = n438 ^ n430 ;
  assign n446 = n445 ^ n439 ;
  assign n447 = n446 ^ n403 ;
  assign n449 = n448 ^ n447 ;
  assign n471 = n470 ^ n449 ;
  assign n472 = n471 ^ n462 ;
  assign n473 = n472 ^ x8 ;
  assign n481 = x10 ^ x9 ;
  assign n480 = x10 ^ x5 ;
  assign n482 = n481 ^ n480 ;
  assign n483 = n480 ^ x10 ;
  assign n484 = n482 & n483 ;
  assign n485 = n484 ^ n480 ;
  assign n486 = ~x8 & n485 ;
  assign n487 = n486 ^ x10 ;
  assign n488 = n203 & ~n487 ;
  assign n489 = n488 ^ n203 ;
  assign n490 = n479 & n489 ;
  assign n491 = n490 ^ n479 ;
  assign n492 = n491 ^ n489 ;
  assign n498 = x9 & x10 ;
  assign n499 = n498 ^ x9 ;
  assign n500 = n499 ^ x10 ;
  assign n501 = x8 & ~n500 ;
  assign n502 = n497 & n501 ;
  assign n503 = n502 ^ n500 ;
  assign n514 = ~n64 & ~n203 ;
  assign n515 = ~n503 & n514 ;
  assign n516 = ~n492 & n515 ;
  assign n506 = x2 & x6 ;
  assign n507 = n506 ^ x6 ;
  assign n508 = x7 & n507 ;
  assign n509 = n508 ^ n507 ;
  assign n504 = n269 ^ x3 ;
  assign n505 = x7 & n504 ;
  assign n510 = n509 ^ n505 ;
  assign n511 = n64 & ~n510 ;
  assign n512 = ~n503 & n511 ;
  assign n513 = ~n492 & n512 ;
  assign n517 = n516 ^ n513 ;
  assign n518 = n473 & n517 ;
  assign n534 = n533 ^ n518 ;
  assign n535 = x7 & n431 ;
  assign n536 = ~x2 & n29 ;
  assign n537 = n535 & n536 ;
  assign n538 = ~x5 & ~x6 ;
  assign n539 = ~x4 & ~x7 ;
  assign n540 = ~x8 & n539 ;
  assign n541 = n538 & n540 ;
  assign n542 = ~n537 & ~n541 ;
  assign n543 = ~x3 & ~n500 ;
  assign n544 = ~n542 & n543 ;
  assign n545 = x3 & ~x7 ;
  assign n546 = n15 & n545 ;
  assign n558 = ~x5 & x7 ;
  assign n559 = n546 & n558 ;
  assign n557 = n44 & n546 ;
  assign n560 = n559 ^ n557 ;
  assign n550 = x6 & n219 ;
  assign n547 = ~x5 & ~x7 ;
  assign n551 = n550 ^ n547 ;
  assign n555 = n493 & ~n551 ;
  assign n556 = n555 ^ n551 ;
  assign n561 = n560 ^ n556 ;
  assign n570 = ~x8 & ~n561 ;
  assign n548 = ~n431 & ~n547 ;
  assign n549 = n546 & n548 ;
  assign n552 = n551 ^ n549 ;
  assign n553 = ~x4 & ~n493 ;
  assign n568 = ~x8 & n553 ;
  assign n569 = n552 & n568 ;
  assign n571 = n570 ^ n569 ;
  assign n554 = n552 & n553 ;
  assign n562 = n561 ^ n554 ;
  assign n563 = n412 & n538 ;
  assign n564 = ~n494 & ~n563 ;
  assign n565 = ~x8 & n454 ;
  assign n566 = ~n564 & n565 ;
  assign n567 = n562 & n566 ;
  assign n572 = n571 ^ n567 ;
  assign n573 = n12 & n431 ;
  assign n574 = x9 & ~n573 ;
  assign n577 = n64 & n204 ;
  assign n578 = x2 & ~x3 ;
  assign n579 = x3 & x8 ;
  assign n580 = ~n578 & ~n579 ;
  assign n581 = ~x10 & ~n580 ;
  assign n582 = n577 & n581 ;
  assign n583 = ~n574 & n582 ;
  assign n584 = ~n572 & n583 ;
  assign n575 = ~x10 & ~n574 ;
  assign n576 = ~n572 & n575 ;
  assign n585 = n584 ^ n576 ;
  assign n586 = n585 ^ x10 ;
  assign n589 = n54 & n412 ;
  assign n595 = n547 & n589 ;
  assign n596 = n595 ^ n573 ;
  assign n590 = x2 & x4 ;
  assign n597 = n579 & n590 ;
  assign n598 = n535 & n597 ;
  assign n599 = n596 & n598 ;
  assign n593 = n573 & n590 ;
  assign n591 = n547 & n590 ;
  assign n592 = n589 & n591 ;
  assign n594 = n593 ^ n592 ;
  assign n600 = n599 ^ n594 ;
  assign n587 = x4 & n579 ;
  assign n588 = n535 & n587 ;
  assign n601 = n600 ^ n588 ;
  assign n603 = n228 & n431 ;
  assign n604 = ~n14 & ~n538 ;
  assign n605 = ~n500 & n604 ;
  assign n606 = ~n603 & n605 ;
  assign n607 = ~n601 & n606 ;
  assign n602 = ~n500 & ~n601 ;
  assign n608 = n607 ^ n602 ;
  assign n609 = ~n14 & ~n500 ;
  assign n610 = ~n603 & n609 ;
  assign y0 = ~n201 ;
  assign y1 = n392 ;
  assign y2 = ~n534 ;
  assign y3 = ~n544 ;
  assign y4 = n586 ;
  assign y5 = ~n608 ;
  assign y6 = ~n610 ;
endmodule
