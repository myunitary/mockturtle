// Benchmark "/tmp/tmp" written by ABC on Sun Nov  9 12:39:31 2025

module sha3_24cc_firstframe ( 
    n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
    n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127, po128, po129, po130, po131, po132, po133, po134, po135, po136,
    po137, po138, po139, po140, po141, po142, po143, po144, po145, po146,
    po147, po148, po149, po150, po151, po152, po153, po154, po155, po156,
    po157, po158, po159, po160, po161, po162, po163, po164, po165, po166,
    po167, po168, po169, po170, po171, po172, po173, po174, po175, po176,
    po177, po178, po179, po180, po181, po182, po183, po184, po185, po186,
    po187, po188, po189, po190, po191, po192, po193, po194, po195, po196,
    po197, po198, po199, po200, po201, po202, po203, po204, po205, po206,
    po207, po208, po209, po210, po211, po212, po213, po214, po215, po216,
    po217, po218, po219, po220, po221, po222, po223, po224, po225, po226,
    po227, po228, po229, po230, po231, po232, po233, po234, po235, po236,
    po237, po238, po239, po240, po241, po242, po243, po244, po245, po246,
    po247, po248, po249, po250, po251, po252, po253, po254, po255, po256,
    po257, po258, po259, po260, po261, po262, po263, po264, po265, po266,
    po267, po268, po269, po270, po271, po272, po273, po274, po275, po276,
    po277, po278, po279, po280, po281, po282, po283, po284, po285, po286,
    po287, po288, po289, po290, po291, po292, po293, po294, po295, po296,
    po297, po298, po299, po300, po301, po302, po303, po304, po305, po306,
    po307, po308, po309, po310, po311, po312, po313, po314, po315, po316,
    po317, po318, po319, po320, po321, po322, po323, po324, po325, po326,
    po327, po328, po329, po330, po331, po332, po333, po334, po335, po336,
    po337, po338, po339, po340, po341, po342, po343, po344, po345, po346,
    po347, po348, po349, po350, po351, po352, po353, po354, po355, po356,
    po357, po358, po359, po360, po361, po362, po363, po364, po365, po366,
    po367, po368, po369, po370, po371, po372, po373, po374, po375, po376,
    po377, po378, po379, po380, po381, po382, po383, po384, po385, po386,
    po387, po388, po389, po390, po391, po392, po393, po394, po395, po396,
    po397, po398, po399, po400, po401, po402, po403, po404, po405, po406,
    po407, po408, po409, po410, po411, po412, po413, po414, po415, po416,
    po417, po418, po419, po420, po421, po422, po423, po424, po425, po426,
    po427, po428, po429, po430, po431, po432, po433, po434, po435, po436,
    po437, po438, po439, po440, po441, po442, po443, po444, po445, po446,
    po447, po448, po449, po450, po451, po452, po453, po454, po455, po456,
    po457, po458, po459, po460, po461, po462, po463, po464, po465, po466,
    po467, po468, po469, po470, po471, po472, po473, po474, po475, po476,
    po477, po478, po479, po480, po481, po482, po483, po484, po485, po486,
    po487, po488, po489, po490, po491, po492, po493, po494, po495, po496,
    po497, po498, po499, po500, po501, po502, po503, po504, po505, po506,
    po507, po508, po509, po510, po511, po512, po513, po514, po515, po516,
    po517, po518, po519, po520, po521, po522, po523, po524, po525, po526,
    po527, po528, po529, po530, po531, po532, po533, po534, po535, po536,
    po537, po538, po539, po540, po541, po542, po543, po544, po545, po546,
    po547, po548, po549, po550, po551, po552, po553, po554, po555, po556,
    po557, po558, po559, po560, po561, po562, po563, po564, po565, po566,
    po567, po568, po569, po570, po571, po572, po573, po574, po575, po576,
    po577, po578, po579, po580, po581, po582, po583, po584, po585, po586,
    po587, po588, po589, po590, po591, po592, po593, po594, po595, po596,
    po597, po598, po599, po600, po601, po602, po603, po604, po605, po606,
    po607, po608, po609, po610, po611, po612, po613, po614, po615, po616,
    po617, po618, po619, po620, po621, po622, po623, po624, po625, po626,
    po627, po628, po629, po630, po631, po632, po633, po634, po635, po636,
    po637, po638, po639, po640, po641, po642, po643, po644, po645, po646,
    po647, po648, po649, po650, po651, po652, po653, po654, po655, po656,
    po657, po658, po659, po660, po661, po662, po663, po664, po665, po666,
    po667, po668, po669, po670, po671, po672, po673, po674, po675, po676,
    po677, po678, po679, po680, po681, po682, po683, po684, po685, po686,
    po687, po688, po689, po690, po691, po692, po693, po694, po695, po696,
    po697, po698, po699, po700, po701, po702, po703, po704, po705, po706,
    po707, po708, po709, po710, po711, po712, po713, po714, po715, po716,
    po717, po718, po719, po720, po721, po722, po723, po724, po725, po726,
    po727, po728, po729, po730, po731, po732, po733, po734, po735, po736,
    po737, po738, po739, po740, po741, po742, po743, po744, po745, po746,
    po747, po748, po749, po750, po751, po752, po753, po754, po755, po756,
    po757, po758, po759, po760, po761, po762, po763, po764, po765, po766,
    po767, po768, po769, po770, po771, po772, po773, po774, po775, po776,
    po777, po778, po779, po780, po781, po782, po783, po784, po785, po786,
    po787, po788, po789, po790, po791, po792, po793, po794, po795, po796,
    po797, po798, po799, po800, po801, po802, po803, po804, po805, po806,
    po807, po808, po809, po810, po811, po812, po813, po814, po815, po816,
    po817, po818, po819, po820, po821, po822, po823, po824, po825, po826,
    po827, po828, po829, po830, po831, po832, po833, po834, po835, po836,
    po837, po838, po839, po840, po841, po842, po843, po844, po845, po846,
    po847, po848, po849, po850, po851, po852, po853, po854, po855, po856,
    po857, po858, po859, po860, po861, po862, po863, po864, po865, po866,
    po867, po868, po869, po870, po871, po872, po873, po874, po875, po876,
    po877, po878, po879, po880, po881, po882, po883, po884, po885, po886,
    po887, po888, po889, po890, po891, po892, po893, po894, po895, po896,
    po897, po898, po899, po900, po901, po902, po903, po904, po905, po906,
    po907, po908, po909, po910, po911, po912, po913, po914, po915, po916,
    po917, po918, po919, po920, po921, po922, po923, po924, po925, po926,
    po927, po928, po929, po930, po931, po932, po933, po934, po935, po936,
    po937, po938, po939, po940, po941, po942, po943, po944, po945, po946,
    po947, po948, po949, po950, po951, po952, po953, po954, po955, po956,
    po957, po958, po959, po960, po961, po962, po963, po964, po965, po966,
    po967, po968, po969, po970, po971, po972, po973, po974, po975, po976,
    po977, po978, po979, po980, po981, po982, po983, po984, po985, po986,
    po987, po988, po989, po990, po991, po992, po993, po994, po995, po996,
    po997, po998, po999, po1000, po1001, po1002, po1003, po1004, po1005,
    po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014,
    po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023,
    po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032,
    po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041,
    po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050,
    po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059,
    po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068,
    po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077,
    po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086,
    po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095,
    po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104,
    po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113,
    po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122,
    po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131,
    po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140,
    po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149,
    po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158,
    po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167,
    po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176,
    po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185,
    po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194,
    po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203,
    po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212,
    po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221,
    po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230,
    po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239,
    po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248,
    po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257,
    po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266,
    po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275,
    po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284,
    po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293,
    po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302,
    po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311,
    po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320,
    po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329,
    po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338,
    po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347,
    po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356,
    po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365,
    po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374,
    po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383,
    po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392,
    po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401,
    po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410,
    po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419,
    po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428,
    po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437,
    po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446,
    po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455,
    po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464,
    po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473,
    po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482,
    po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491,
    po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500,
    po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509,
    po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518,
    po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527,
    po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536,
    po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545,
    po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554,
    po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563,
    po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572,
    po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581,
    po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590,
    po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599,
    po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608,
    po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617,
    po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626,
    po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635,
    po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644,
    po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653,
    po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662,
    po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671,
    po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680,
    po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689,
    po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698,
    po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707,
    po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716,
    po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725,
    po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734,
    po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743,
    po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752,
    po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761,
    po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770,
    po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779,
    po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788,
    po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797,
    po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806,
    po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815,
    po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824,
    po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833,
    po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842,
    po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851,
    po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860,
    po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869,
    po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878,
    po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887,
    po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896,
    po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905,
    po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914,
    po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923,
    po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932,
    po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941,
    po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950,
    po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959,
    po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968,
    po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977,
    po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986,
    po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995,
    po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004,
    po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013,
    po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022,
    po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031,
    po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040,
    po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049,
    po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058,
    po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067,
    po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076,
    po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085,
    po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094,
    po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103,
    po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112,
    po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121,
    po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130,
    po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139,
    po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148,
    po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157,
    po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166,
    po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175,
    po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184,
    po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193,
    po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202,
    po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211,
    po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220,
    po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229,
    po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238,
    po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247,
    po2248, po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256,
    po2257, po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265,
    po2266, po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274,
    po2275, po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283,
    po2284, po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292,
    po2293, po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301,
    po2302, po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310,
    po2311, po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319,
    po2320, po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328,
    po2329, po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337,
    po2338, po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346,
    po2347, po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355,
    po2356, po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364,
    po2365, po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373,
    po2374, po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382,
    po2383, po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391,
    po2392, po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400,
    po2401, po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409,
    po2410, po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418,
    po2419, po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427,
    po2428, po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436,
    po2437, po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445,
    po2446, po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454,
    po2455, po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463,
    po2464, po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472,
    po2473, po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481,
    po2482, po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490,
    po2491, po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499,
    po2500, po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508,
    po2509, po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517,
    po2518, po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526,
    po2527, po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535,
    po2536, po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544,
    po2545, po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553,
    po2554, po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562,
    po2563, po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571,
    po2572, po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580,
    po2581, po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589,
    po2590, po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598,
    po2599, po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607,
    po2608, po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616,
    po2617, po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625,
    po2626, po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634,
    po2635, po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643,
    po2644, po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652,
    po2653, po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661,
    po2662, po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670,
    po2671, po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679,
    po2680, po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688,
    po2689, po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697,
    po2698, po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706,
    po2707, po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715,
    po2716, po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724,
    po2725, po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733,
    po2734, po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742,
    po2743, po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751,
    po2752, po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760,
    po2761, po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769,
    po2770, po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778,
    po2779, po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787,
    po2788, po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796,
    po2797, po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805,
    po2806, po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814,
    po2815, po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823,
    po2824, po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832,
    po2833, po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841,
    po2842, po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850,
    po2851, po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859,
    po2860, po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868,
    po2869, po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877,
    po2878, po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886,
    po2887, po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895,
    po2896, po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904,
    po2905, po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913,
    po2914, po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922,
    po2923, po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931,
    po2932, po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940,
    po2941, po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949,
    po2950, po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958,
    po2959, po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967,
    po2968, po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976,
    po2977, po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985,
    po2986, po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994,
    po2995, po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003,
    po3004, po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012,
    po3013, po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021,
    po3022, po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030,
    po3031, po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039,
    po3040, po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048,
    po3049, po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057,
    po3058, po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066,
    po3067, po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075,
    po3076, po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084,
    po3085, po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093,
    po3094, po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102,
    po3103, po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111,
    po3112, po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120,
    po3121, po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129,
    po3130, po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138,
    po3139, po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147,
    po3148, po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156,
    po3157, po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165,
    po3166, po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174,
    po3175, po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183,
    po3184, po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192,
    po3193, po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201,
    po3202, po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210,
    po3211, po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219,
    po3220, po3221, po3222, po3223, po3224  );
  input  n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
    n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
    n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127, po128, po129, po130, po131, po132, po133, po134, po135, po136,
    po137, po138, po139, po140, po141, po142, po143, po144, po145, po146,
    po147, po148, po149, po150, po151, po152, po153, po154, po155, po156,
    po157, po158, po159, po160, po161, po162, po163, po164, po165, po166,
    po167, po168, po169, po170, po171, po172, po173, po174, po175, po176,
    po177, po178, po179, po180, po181, po182, po183, po184, po185, po186,
    po187, po188, po189, po190, po191, po192, po193, po194, po195, po196,
    po197, po198, po199, po200, po201, po202, po203, po204, po205, po206,
    po207, po208, po209, po210, po211, po212, po213, po214, po215, po216,
    po217, po218, po219, po220, po221, po222, po223, po224, po225, po226,
    po227, po228, po229, po230, po231, po232, po233, po234, po235, po236,
    po237, po238, po239, po240, po241, po242, po243, po244, po245, po246,
    po247, po248, po249, po250, po251, po252, po253, po254, po255, po256,
    po257, po258, po259, po260, po261, po262, po263, po264, po265, po266,
    po267, po268, po269, po270, po271, po272, po273, po274, po275, po276,
    po277, po278, po279, po280, po281, po282, po283, po284, po285, po286,
    po287, po288, po289, po290, po291, po292, po293, po294, po295, po296,
    po297, po298, po299, po300, po301, po302, po303, po304, po305, po306,
    po307, po308, po309, po310, po311, po312, po313, po314, po315, po316,
    po317, po318, po319, po320, po321, po322, po323, po324, po325, po326,
    po327, po328, po329, po330, po331, po332, po333, po334, po335, po336,
    po337, po338, po339, po340, po341, po342, po343, po344, po345, po346,
    po347, po348, po349, po350, po351, po352, po353, po354, po355, po356,
    po357, po358, po359, po360, po361, po362, po363, po364, po365, po366,
    po367, po368, po369, po370, po371, po372, po373, po374, po375, po376,
    po377, po378, po379, po380, po381, po382, po383, po384, po385, po386,
    po387, po388, po389, po390, po391, po392, po393, po394, po395, po396,
    po397, po398, po399, po400, po401, po402, po403, po404, po405, po406,
    po407, po408, po409, po410, po411, po412, po413, po414, po415, po416,
    po417, po418, po419, po420, po421, po422, po423, po424, po425, po426,
    po427, po428, po429, po430, po431, po432, po433, po434, po435, po436,
    po437, po438, po439, po440, po441, po442, po443, po444, po445, po446,
    po447, po448, po449, po450, po451, po452, po453, po454, po455, po456,
    po457, po458, po459, po460, po461, po462, po463, po464, po465, po466,
    po467, po468, po469, po470, po471, po472, po473, po474, po475, po476,
    po477, po478, po479, po480, po481, po482, po483, po484, po485, po486,
    po487, po488, po489, po490, po491, po492, po493, po494, po495, po496,
    po497, po498, po499, po500, po501, po502, po503, po504, po505, po506,
    po507, po508, po509, po510, po511, po512, po513, po514, po515, po516,
    po517, po518, po519, po520, po521, po522, po523, po524, po525, po526,
    po527, po528, po529, po530, po531, po532, po533, po534, po535, po536,
    po537, po538, po539, po540, po541, po542, po543, po544, po545, po546,
    po547, po548, po549, po550, po551, po552, po553, po554, po555, po556,
    po557, po558, po559, po560, po561, po562, po563, po564, po565, po566,
    po567, po568, po569, po570, po571, po572, po573, po574, po575, po576,
    po577, po578, po579, po580, po581, po582, po583, po584, po585, po586,
    po587, po588, po589, po590, po591, po592, po593, po594, po595, po596,
    po597, po598, po599, po600, po601, po602, po603, po604, po605, po606,
    po607, po608, po609, po610, po611, po612, po613, po614, po615, po616,
    po617, po618, po619, po620, po621, po622, po623, po624, po625, po626,
    po627, po628, po629, po630, po631, po632, po633, po634, po635, po636,
    po637, po638, po639, po640, po641, po642, po643, po644, po645, po646,
    po647, po648, po649, po650, po651, po652, po653, po654, po655, po656,
    po657, po658, po659, po660, po661, po662, po663, po664, po665, po666,
    po667, po668, po669, po670, po671, po672, po673, po674, po675, po676,
    po677, po678, po679, po680, po681, po682, po683, po684, po685, po686,
    po687, po688, po689, po690, po691, po692, po693, po694, po695, po696,
    po697, po698, po699, po700, po701, po702, po703, po704, po705, po706,
    po707, po708, po709, po710, po711, po712, po713, po714, po715, po716,
    po717, po718, po719, po720, po721, po722, po723, po724, po725, po726,
    po727, po728, po729, po730, po731, po732, po733, po734, po735, po736,
    po737, po738, po739, po740, po741, po742, po743, po744, po745, po746,
    po747, po748, po749, po750, po751, po752, po753, po754, po755, po756,
    po757, po758, po759, po760, po761, po762, po763, po764, po765, po766,
    po767, po768, po769, po770, po771, po772, po773, po774, po775, po776,
    po777, po778, po779, po780, po781, po782, po783, po784, po785, po786,
    po787, po788, po789, po790, po791, po792, po793, po794, po795, po796,
    po797, po798, po799, po800, po801, po802, po803, po804, po805, po806,
    po807, po808, po809, po810, po811, po812, po813, po814, po815, po816,
    po817, po818, po819, po820, po821, po822, po823, po824, po825, po826,
    po827, po828, po829, po830, po831, po832, po833, po834, po835, po836,
    po837, po838, po839, po840, po841, po842, po843, po844, po845, po846,
    po847, po848, po849, po850, po851, po852, po853, po854, po855, po856,
    po857, po858, po859, po860, po861, po862, po863, po864, po865, po866,
    po867, po868, po869, po870, po871, po872, po873, po874, po875, po876,
    po877, po878, po879, po880, po881, po882, po883, po884, po885, po886,
    po887, po888, po889, po890, po891, po892, po893, po894, po895, po896,
    po897, po898, po899, po900, po901, po902, po903, po904, po905, po906,
    po907, po908, po909, po910, po911, po912, po913, po914, po915, po916,
    po917, po918, po919, po920, po921, po922, po923, po924, po925, po926,
    po927, po928, po929, po930, po931, po932, po933, po934, po935, po936,
    po937, po938, po939, po940, po941, po942, po943, po944, po945, po946,
    po947, po948, po949, po950, po951, po952, po953, po954, po955, po956,
    po957, po958, po959, po960, po961, po962, po963, po964, po965, po966,
    po967, po968, po969, po970, po971, po972, po973, po974, po975, po976,
    po977, po978, po979, po980, po981, po982, po983, po984, po985, po986,
    po987, po988, po989, po990, po991, po992, po993, po994, po995, po996,
    po997, po998, po999, po1000, po1001, po1002, po1003, po1004, po1005,
    po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014,
    po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023,
    po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032,
    po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041,
    po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050,
    po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059,
    po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068,
    po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077,
    po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086,
    po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095,
    po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104,
    po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113,
    po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122,
    po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131,
    po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140,
    po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149,
    po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158,
    po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167,
    po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176,
    po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185,
    po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194,
    po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203,
    po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212,
    po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221,
    po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230,
    po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239,
    po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248,
    po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257,
    po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266,
    po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275,
    po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284,
    po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293,
    po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302,
    po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311,
    po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320,
    po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329,
    po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338,
    po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347,
    po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356,
    po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365,
    po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374,
    po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383,
    po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392,
    po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401,
    po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410,
    po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419,
    po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428,
    po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437,
    po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446,
    po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455,
    po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464,
    po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473,
    po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482,
    po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491,
    po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500,
    po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509,
    po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518,
    po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527,
    po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536,
    po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545,
    po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554,
    po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563,
    po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572,
    po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581,
    po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590,
    po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599,
    po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608,
    po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617,
    po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626,
    po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635,
    po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644,
    po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653,
    po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662,
    po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671,
    po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680,
    po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689,
    po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698,
    po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707,
    po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716,
    po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725,
    po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734,
    po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743,
    po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752,
    po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761,
    po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770,
    po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779,
    po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788,
    po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797,
    po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806,
    po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815,
    po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824,
    po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833,
    po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842,
    po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851,
    po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860,
    po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869,
    po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878,
    po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887,
    po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896,
    po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905,
    po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914,
    po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923,
    po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932,
    po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941,
    po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950,
    po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959,
    po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968,
    po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977,
    po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986,
    po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995,
    po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004,
    po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013,
    po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022,
    po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031,
    po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040,
    po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049,
    po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058,
    po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067,
    po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076,
    po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085,
    po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094,
    po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103,
    po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112,
    po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121,
    po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130,
    po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139,
    po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148,
    po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157,
    po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166,
    po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175,
    po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184,
    po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193,
    po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202,
    po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211,
    po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220,
    po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229,
    po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238,
    po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247,
    po2248, po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256,
    po2257, po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265,
    po2266, po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274,
    po2275, po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283,
    po2284, po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292,
    po2293, po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301,
    po2302, po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310,
    po2311, po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319,
    po2320, po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328,
    po2329, po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337,
    po2338, po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346,
    po2347, po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355,
    po2356, po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364,
    po2365, po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373,
    po2374, po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382,
    po2383, po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391,
    po2392, po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400,
    po2401, po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409,
    po2410, po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418,
    po2419, po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427,
    po2428, po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436,
    po2437, po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445,
    po2446, po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454,
    po2455, po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463,
    po2464, po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472,
    po2473, po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481,
    po2482, po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490,
    po2491, po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499,
    po2500, po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508,
    po2509, po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517,
    po2518, po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526,
    po2527, po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535,
    po2536, po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544,
    po2545, po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553,
    po2554, po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562,
    po2563, po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571,
    po2572, po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580,
    po2581, po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589,
    po2590, po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598,
    po2599, po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607,
    po2608, po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616,
    po2617, po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625,
    po2626, po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634,
    po2635, po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643,
    po2644, po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652,
    po2653, po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661,
    po2662, po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670,
    po2671, po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679,
    po2680, po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688,
    po2689, po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697,
    po2698, po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706,
    po2707, po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715,
    po2716, po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724,
    po2725, po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733,
    po2734, po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742,
    po2743, po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751,
    po2752, po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760,
    po2761, po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769,
    po2770, po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778,
    po2779, po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787,
    po2788, po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796,
    po2797, po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805,
    po2806, po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814,
    po2815, po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823,
    po2824, po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832,
    po2833, po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841,
    po2842, po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850,
    po2851, po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859,
    po2860, po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868,
    po2869, po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877,
    po2878, po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886,
    po2887, po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895,
    po2896, po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904,
    po2905, po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913,
    po2914, po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922,
    po2923, po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931,
    po2932, po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940,
    po2941, po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949,
    po2950, po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958,
    po2959, po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967,
    po2968, po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976,
    po2977, po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985,
    po2986, po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994,
    po2995, po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003,
    po3004, po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012,
    po3013, po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021,
    po3022, po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030,
    po3031, po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039,
    po3040, po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048,
    po3049, po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057,
    po3058, po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066,
    po3067, po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075,
    po3076, po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084,
    po3085, po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093,
    po3094, po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102,
    po3103, po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111,
    po3112, po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120,
    po3121, po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129,
    po3130, po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138,
    po3139, po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147,
    po3148, po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156,
    po3157, po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165,
    po3166, po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174,
    po3175, po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183,
    po3184, po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192,
    po3193, po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201,
    po3202, po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210,
    po3211, po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219,
    po3220, po3221, po3222, po3223, po3224;
  wire new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510, new_n1511, new_n1512,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1564, new_n1565, new_n1566,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1584,
    new_n1585, new_n1586, new_n1587, new_n1588, new_n1589, new_n1590,
    new_n1591, new_n1592, new_n1593, new_n1594, new_n1595, new_n1596,
    new_n1597, new_n1598, new_n1599, new_n1600, new_n1601, new_n1602,
    new_n1603, new_n1604, new_n1605, new_n1606, new_n1607, new_n1608,
    new_n1609, new_n1610, new_n1611, new_n1612, new_n1613, new_n1614,
    new_n1615, new_n1616, new_n1617, new_n1618, new_n1619, new_n1620,
    new_n1621, new_n1622, new_n1623, new_n1624, new_n1625, new_n1626,
    new_n1627, new_n1628, new_n1629, new_n1630, new_n1631, new_n1632,
    new_n1633, new_n1634, new_n1635, new_n1636, new_n1637, new_n1638,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1644,
    new_n1645, new_n1646, new_n1647, new_n1648, new_n1649, new_n1650,
    new_n1651, new_n1652, new_n1653, new_n1654, new_n1655, new_n1656,
    new_n1657, new_n1658, new_n1659, new_n1660, new_n1661, new_n1662,
    new_n1663, new_n1664, new_n1665, new_n1666, new_n1667, new_n1668,
    new_n1669, new_n1670, new_n1671, new_n1672, new_n1673, new_n1674,
    new_n1675, new_n1676, new_n1677, new_n1678, new_n1679, new_n1680,
    new_n1681, new_n1682, new_n1683, new_n1684, new_n1685, new_n1686,
    new_n1687, new_n1688, new_n1689, new_n1690, new_n1691, new_n1692,
    new_n1693, new_n1694, new_n1695, new_n1696, new_n1697, new_n1698,
    new_n1699, new_n1700, new_n1701, new_n1702, new_n1703, new_n1704,
    new_n1705, new_n1706, new_n1707, new_n1708, new_n1709, new_n1710,
    new_n1711, new_n1712, new_n1713, new_n1714, new_n1715, new_n1716,
    new_n1717, new_n1718, new_n1719, new_n1720, new_n1721, new_n1722,
    new_n1723, new_n1724, new_n1725, new_n1726, new_n1727, new_n1728,
    new_n1729, new_n1730, new_n1731, new_n1732, new_n1733, new_n1734,
    new_n1735, new_n1736, new_n1737, new_n1738, new_n1739, new_n1740,
    new_n1741, new_n1742, new_n1743, new_n1744, new_n1745, new_n1746,
    new_n1747, new_n1748, new_n1749, new_n1750, new_n1751, new_n1752,
    new_n1753, new_n1754, new_n1755, new_n1756, new_n1757, new_n1758,
    new_n1759, new_n1760, new_n1761, new_n1762, new_n1763, new_n1764,
    new_n1765, new_n1766, new_n1767, new_n1768, new_n1769, new_n1770,
    new_n1771, new_n1772, new_n1773, new_n1774, new_n1775, new_n1776,
    new_n1777, new_n1778, new_n1779, new_n1780, new_n1781, new_n1782,
    new_n1783, new_n1784, new_n1785, new_n1786, new_n1787, new_n1788,
    new_n1789, new_n1790, new_n1791, new_n1792, new_n1793, new_n1794,
    new_n1795, new_n1796, new_n1797, new_n1798, new_n1799, new_n1800,
    new_n1801, new_n1802, new_n1803, new_n1804, new_n1805, new_n1806,
    new_n1807, new_n1808, new_n1809, new_n1810, new_n1811, new_n1812,
    new_n1813, new_n1814, new_n1815, new_n1816, new_n1817, new_n1818,
    new_n1819, new_n1820, new_n1821, new_n1822, new_n1823, new_n1824,
    new_n1825, new_n1826, new_n1827, new_n1828, new_n1829, new_n1830,
    new_n1831, new_n1832, new_n1833, new_n1834, new_n1835, new_n1836,
    new_n1837, new_n1838, new_n1839, new_n1840, new_n1841, new_n1842,
    new_n1843, new_n1844, new_n1845, new_n1846, new_n1847, new_n1848,
    new_n1849, new_n1850, new_n1851, new_n1852, new_n1853, new_n1854,
    new_n1855, new_n1856, new_n1857, new_n1858, new_n1859, new_n1860,
    new_n1861, new_n1862, new_n1863, new_n1864, new_n1865, new_n1866,
    new_n1867, new_n1868, new_n1869, new_n1870, new_n1871, new_n1872,
    new_n1873, new_n1874, new_n1875, new_n1876, new_n1877, new_n1878,
    new_n1879, new_n1880, new_n1881, new_n1882, new_n1883, new_n1884,
    new_n1885, new_n1886, new_n1887, new_n1888, new_n1889, new_n1890,
    new_n1891, new_n1892, new_n1893, new_n1894, new_n1895, new_n1896,
    new_n1897, new_n1898, new_n1899, new_n1900, new_n1901, new_n1902,
    new_n1903, new_n1904, new_n1905, new_n1906, new_n1907, new_n1908,
    new_n1909, new_n1910, new_n1911, new_n1912, new_n1913, new_n1914,
    new_n1915, new_n1916, new_n1917, new_n1918, new_n1919, new_n1920,
    new_n1921, new_n1922, new_n1923, new_n1924, new_n1925, new_n1926,
    new_n1927, new_n1928, new_n1929, new_n1930, new_n1931, new_n1932,
    new_n1933, new_n1934, new_n1935, new_n1936, new_n1937, new_n1938,
    new_n1939, new_n1940, new_n1941, new_n1942, new_n1943, new_n1944,
    new_n1945, new_n1946, new_n1947, new_n1948, new_n1949, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986,
    new_n1987, new_n1988, new_n1989, new_n1990, new_n1991, new_n1992,
    new_n1993, new_n1994, new_n1995, new_n1996, new_n1997, new_n1998,
    new_n1999, new_n2000, new_n2001, new_n2002, new_n2003, new_n2004,
    new_n2005, new_n2006, new_n2007, new_n2008, new_n2009, new_n2010,
    new_n2011, new_n2012, new_n2013, new_n2014, new_n2015, new_n2016,
    new_n2017, new_n2018, new_n2019, new_n2020, new_n2021, new_n2022,
    new_n2023, new_n2024, new_n2025, new_n2026, new_n2027, new_n2028,
    new_n2029, new_n2030, new_n2031, new_n2032, new_n2033, new_n2034,
    new_n2035, new_n2036, new_n2037, new_n2038, new_n2039, new_n2040,
    new_n2041, new_n2042, new_n2043, new_n2044, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058,
    new_n2059, new_n2060, new_n2061, new_n2062, new_n2063, new_n2064,
    new_n2065, new_n2066, new_n2067, new_n2068, new_n2069, new_n2070,
    new_n2071, new_n2072, new_n2073, new_n2074, new_n2075, new_n2076,
    new_n2077, new_n2078, new_n2079, new_n2080, new_n2081, new_n2082,
    new_n2083, new_n2084, new_n2085, new_n2086, new_n2087, new_n2088,
    new_n2089, new_n2090, new_n2091, new_n2092, new_n2093, new_n2094,
    new_n2095, new_n2096, new_n2097, new_n2098, new_n2099, new_n2100,
    new_n2101, new_n2102, new_n2103, new_n2104, new_n2105, new_n2106,
    new_n2107, new_n2108, new_n2109, new_n2110, new_n2111, new_n2112,
    new_n2113, new_n2114, new_n2115, new_n2116, new_n2117, new_n2118,
    new_n2119, new_n2120, new_n2121, new_n2122, new_n2123, new_n2124,
    new_n2125, new_n2126, new_n2127, new_n2128, new_n2129, new_n2130,
    new_n2131, new_n2132, new_n2133, new_n2134, new_n2135, new_n2136,
    new_n2137, new_n2138, new_n2139, new_n2140, new_n2141, new_n2142,
    new_n2143, new_n2144, new_n2145, new_n2146, new_n2147, new_n2148,
    new_n2149, new_n2150, new_n2151, new_n2152, new_n2153, new_n2154,
    new_n2155, new_n2156, new_n2157, new_n2158, new_n2159, new_n2160,
    new_n2161, new_n2162, new_n2163, new_n2164, new_n2165, new_n2166,
    new_n2167, new_n2168, new_n2169, new_n2170, new_n2171, new_n2172,
    new_n2173, new_n2174, new_n2175, new_n2176, new_n2177, new_n2178,
    new_n2179, new_n2180, new_n2181, new_n2182, new_n2183, new_n2184,
    new_n2185, new_n2186, new_n2187, new_n2188, new_n2189, new_n2190,
    new_n2191, new_n2192, new_n2193, new_n2194, new_n2195, new_n2196,
    new_n2197, new_n2198, new_n2199, new_n2200, new_n2201, new_n2202,
    new_n2203, new_n2204, new_n2205, new_n2206, new_n2207, new_n2208,
    new_n2209, new_n2210, new_n2211, new_n2212, new_n2213, new_n2214,
    new_n2215, new_n2216, new_n2217, new_n2218, new_n2219, new_n2220,
    new_n2221, new_n2222, new_n2223, new_n2224, new_n2225, new_n2226,
    new_n2227, new_n2228, new_n2229, new_n2230, new_n2231, new_n2232,
    new_n2233, new_n2234, new_n2235, new_n2236, new_n2237, new_n2238,
    new_n2239, new_n2240, new_n2241, new_n2242, new_n2243, new_n2244,
    new_n2245, new_n2246, new_n2247, new_n2248, new_n2249, new_n2250,
    new_n2251, new_n2252, new_n2253, new_n2254, new_n2255, new_n2256,
    new_n2257, new_n2258, new_n2259, new_n2260, new_n2261, new_n2262,
    new_n2263, new_n2264, new_n2265, new_n2266, new_n2267, new_n2268,
    new_n2269, new_n2270, new_n2271, new_n2272, new_n2273, new_n2274,
    new_n2275, new_n2276, new_n2277, new_n2278, new_n2279, new_n2280,
    new_n2281, new_n2282, new_n2283, new_n2284, new_n2285, new_n2286,
    new_n2287, new_n2288, new_n2289, new_n2290, new_n2291, new_n2292,
    new_n2293, new_n2294, new_n2295, new_n2296, new_n2297, new_n2298,
    new_n2299, new_n2300, new_n2301, new_n2302, new_n2303, new_n2304,
    new_n2305, new_n2306, new_n2307, new_n2308, new_n2309, new_n2310,
    new_n2311, new_n2312, new_n2313, new_n2314, new_n2315, new_n2316,
    new_n2317, new_n2318, new_n2319, new_n2320, new_n2321, new_n2322,
    new_n2323, new_n2324, new_n2325, new_n2326, new_n2327, new_n2328,
    new_n2329, new_n2330, new_n2331, new_n2332, new_n2333, new_n2334,
    new_n2335, new_n2336, new_n2337, new_n2338, new_n2339, new_n2340,
    new_n2341, new_n2342, new_n2343, new_n2344, new_n2345, new_n2346,
    new_n2347, new_n2348, new_n2349, new_n2350, new_n2351, new_n2352,
    new_n2353, new_n2354, new_n2355, new_n2356, new_n2357, new_n2358,
    new_n2359, new_n2360, new_n2361, new_n2362, new_n2363, new_n2364,
    new_n2365, new_n2366, new_n2367, new_n2368, new_n2369, new_n2370,
    new_n2371, new_n2372, new_n2373, new_n2374, new_n2375, new_n2376,
    new_n2377, new_n2378, new_n2379, new_n2380, new_n2381, new_n2382,
    new_n2383, new_n2384, new_n2385, new_n2386, new_n2387, new_n2388,
    new_n2389, new_n2390, new_n2391, new_n2392, new_n2393, new_n2394,
    new_n2395, new_n2396, new_n2397, new_n2398, new_n2399, new_n2400,
    new_n2401, new_n2402, new_n2403, new_n2404, new_n2405, new_n2406,
    new_n2407, new_n2408, new_n2409, new_n2410, new_n2411, new_n2412,
    new_n2413, new_n2414, new_n2415, new_n2416, new_n2417, new_n2418,
    new_n2419, new_n2420, new_n2421, new_n2422, new_n2423, new_n2424,
    new_n2425, new_n2426, new_n2427, new_n2428, new_n2429, new_n2430,
    new_n2431, new_n2432, new_n2433, new_n2434, new_n2435, new_n2436,
    new_n2437, new_n2438, new_n2439, new_n2440, new_n2441, new_n2442,
    new_n2443, new_n2444, new_n2445, new_n2446, new_n2447, new_n2448,
    new_n2449, new_n2450, new_n2451, new_n2452, new_n2453, new_n2454,
    new_n2455, new_n2456, new_n2457, new_n2458, new_n2459, new_n2460,
    new_n2461, new_n2462, new_n2463, new_n2464, new_n2465, new_n2466,
    new_n2467, new_n2468, new_n2469, new_n2470, new_n2471, new_n2472,
    new_n2473, new_n2474, new_n2475, new_n2476, new_n2477, new_n2478,
    new_n2479, new_n2480, new_n2481, new_n2482, new_n2483, new_n2484,
    new_n2485, new_n2486, new_n2487, new_n2488, new_n2489, new_n2490,
    new_n2491, new_n2492, new_n2493, new_n2494, new_n2495, new_n2496,
    new_n2497, new_n2498, new_n2499, new_n2500, new_n2501, new_n2502,
    new_n2503, new_n2504, new_n2505, new_n2506, new_n2507, new_n2508,
    new_n2509, new_n2510, new_n2511, new_n2512, new_n2513, new_n2514,
    new_n2515, new_n2516, new_n2517, new_n2518, new_n2519, new_n2520,
    new_n2521, new_n2522, new_n2523, new_n2524, new_n2525, new_n2526,
    new_n2527, new_n2528, new_n2529, new_n2530, new_n2531, new_n2532,
    new_n2533, new_n2534, new_n2535, new_n2536, new_n2537, new_n2538,
    new_n2539, new_n2540, new_n2541, new_n2542, new_n2543, new_n2544,
    new_n2545, new_n2546, new_n2547, new_n2548, new_n2549, new_n2550,
    new_n2551, new_n2552, new_n2553, new_n2554, new_n2555, new_n2556,
    new_n2557, new_n2558, new_n2559, new_n2560, new_n2561, new_n2562,
    new_n2563, new_n2564, new_n2565, new_n2566, new_n2567, new_n2568,
    new_n2569, new_n2570, new_n2571, new_n2572, new_n2573, new_n2574,
    new_n2575, new_n2576, new_n2577, new_n2578, new_n2579, new_n2580,
    new_n2581, new_n2582, new_n2583, new_n2584, new_n2585, new_n2586,
    new_n2587, new_n2588, new_n2589, new_n2590, new_n2591, new_n2592,
    new_n2593, new_n2594, new_n2595, new_n2596, new_n2597, new_n2598,
    new_n2599, new_n2600, new_n2601, new_n2602, new_n2603, new_n2604,
    new_n2605, new_n2606, new_n2607, new_n2608, new_n2609, new_n2610,
    new_n2611, new_n2612, new_n2613, new_n2614, new_n2615, new_n2616,
    new_n2617, new_n2618, new_n2619, new_n2620, new_n2621, new_n2622,
    new_n2623, new_n2624, new_n2625, new_n2626, new_n2627, new_n2628,
    new_n2629, new_n2630, new_n2631, new_n2632, new_n2633, new_n2634,
    new_n2635, new_n2636, new_n2637, new_n2638, new_n2639, new_n2640,
    new_n2641, new_n2642, new_n2643, new_n2644, new_n2645, new_n2646,
    new_n2647, new_n2648, new_n2649, new_n2650, new_n2651, new_n2652,
    new_n2653, new_n2654, new_n2655, new_n2656, new_n2657, new_n2658,
    new_n2659, new_n2660, new_n2661, new_n2662, new_n2663, new_n2664,
    new_n2665, new_n2666, new_n2667, new_n2668, new_n2669, new_n2670,
    new_n2671, new_n2672, new_n2673, new_n2674, new_n2675, new_n2676,
    new_n2677, new_n2678, new_n2679, new_n2680, new_n2681, new_n2682,
    new_n2683, new_n2684, new_n2685, new_n2686, new_n2687, new_n2688,
    new_n2689, new_n2690, new_n2691, new_n2692, new_n2693, new_n2694,
    new_n2695, new_n2696, new_n2697, new_n2698, new_n2699, new_n2700,
    new_n2701, new_n2702, new_n2703, new_n2704, new_n2705, new_n2706,
    new_n2707, new_n2708, new_n2709, new_n2710, new_n2711, new_n2712,
    new_n2713, new_n2714, new_n2715, new_n2716, new_n2717, new_n2718,
    new_n2719, new_n2720, new_n2721, new_n2722, new_n2723, new_n2724,
    new_n2725, new_n2726, new_n2727, new_n2728, new_n2729, new_n2730,
    new_n2731, new_n2732, new_n2733, new_n2734, new_n2735, new_n2736,
    new_n2737, new_n2738, new_n2739, new_n2740, new_n2741, new_n2742,
    new_n2743, new_n2744, new_n2745, new_n2746, new_n2747, new_n2748,
    new_n2749, new_n2750, new_n2751, new_n2752, new_n2753, new_n2754,
    new_n2755, new_n2756, new_n2757, new_n2758, new_n2759, new_n2760,
    new_n2761, new_n2762, new_n2763, new_n2764, new_n2765, new_n2766,
    new_n2767, new_n2768, new_n2769, new_n2770, new_n2771, new_n2772,
    new_n2773, new_n2774, new_n2775, new_n2776, new_n2777, new_n2778,
    new_n2779, new_n2780, new_n2781, new_n2782, new_n2783, new_n2784,
    new_n2785, new_n2786, new_n2787, new_n2788, new_n2789, new_n2790,
    new_n2791, new_n2792, new_n2793, new_n2794, new_n2795, new_n2796,
    new_n2797, new_n2798, new_n2799, new_n2800, new_n2801, new_n2802,
    new_n2803, new_n2804, new_n2805, new_n2806, new_n2807, new_n2808,
    new_n2809, new_n2810, new_n2811, new_n2812, new_n2813, new_n2814,
    new_n2815, new_n2816, new_n2817, new_n2818, new_n2819, new_n2820,
    new_n2821, new_n2822, new_n2823, new_n2824, new_n2825, new_n2826,
    new_n2827, new_n2828, new_n2829, new_n2830, new_n2831, new_n2832,
    new_n2833, new_n2834, new_n2835, new_n2836, new_n2837, new_n2838,
    new_n2839, new_n2840, new_n2841, new_n2842, new_n2843, new_n2844,
    new_n2845, new_n2846, new_n2847, new_n2848, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2853, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858, new_n2859, new_n2860, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874,
    new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886,
    new_n2887, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944, new_n2945, new_n2946,
    new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978, new_n2979, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017, new_n3018,
    new_n3019, new_n3020, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125, new_n3126,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156,
    new_n3157, new_n3158, new_n3159, new_n3160, new_n3161, new_n3162,
    new_n3163, new_n3164, new_n3165, new_n3166, new_n3167, new_n3168,
    new_n3169, new_n3170, new_n3171, new_n3172, new_n3173, new_n3174,
    new_n3175, new_n3176, new_n3177, new_n3178, new_n3179, new_n3180,
    new_n3181, new_n3182, new_n3183, new_n3184, new_n3185, new_n3186,
    new_n3187, new_n3188, new_n3189, new_n3190, new_n3191, new_n3192,
    new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198,
    new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204,
    new_n3205, new_n3206, new_n3207, new_n3208, new_n3209, new_n3210,
    new_n3211, new_n3212, new_n3213, new_n3214, new_n3215, new_n3216,
    new_n3217, new_n3218, new_n3219, new_n3220, new_n3221, new_n3222,
    new_n3223, new_n3224, new_n3225, new_n3226, new_n3227, new_n3228,
    new_n3229, new_n3230, new_n3231, new_n3232, new_n3233, new_n3234,
    new_n3235, new_n3236, new_n3237, new_n3238, new_n3239, new_n3240,
    new_n3241, new_n3242, new_n3243, new_n3244, new_n3245, new_n3246,
    new_n3247, new_n3248, new_n3249, new_n3250, new_n3251, new_n3252,
    new_n3253, new_n3254, new_n3255, new_n3256, new_n3257, new_n3258,
    new_n3259, new_n3260, new_n3261, new_n3262, new_n3263, new_n3264,
    new_n3265, new_n3266, new_n3267, new_n3268, new_n3269, new_n3270,
    new_n3271, new_n3272, new_n3273, new_n3274, new_n3275, new_n3276,
    new_n3277, new_n3278, new_n3279, new_n3280, new_n3281, new_n3282,
    new_n3283, new_n3284, new_n3285, new_n3286, new_n3287, new_n3288,
    new_n3289, new_n3290, new_n3291, new_n3292, new_n3293, new_n3294,
    new_n3295, new_n3296, new_n3297, new_n3298, new_n3299, new_n3300,
    new_n3301, new_n3302, new_n3303, new_n3304, new_n3305, new_n3306,
    new_n3307, new_n3308, new_n3309, new_n3310, new_n3311, new_n3312,
    new_n3313, new_n3314, new_n3315, new_n3316, new_n3317, new_n3318,
    new_n3319, new_n3320, new_n3321, new_n3322, new_n3323, new_n3324,
    new_n3325, new_n3326, new_n3327, new_n3328, new_n3329, new_n3330,
    new_n3331, new_n3332, new_n3333, new_n3334, new_n3335, new_n3336,
    new_n3337, new_n3338, new_n3339, new_n3340, new_n3341, new_n3342,
    new_n3343, new_n3344, new_n3345, new_n3346, new_n3347, new_n3348,
    new_n3349, new_n3350, new_n3351, new_n3352, new_n3353, new_n3354,
    new_n3355, new_n3356, new_n3357, new_n3358, new_n3359, new_n3360,
    new_n3361, new_n3362, new_n3363, new_n3364, new_n3365, new_n3366,
    new_n3367, new_n3368, new_n3369, new_n3370, new_n3371, new_n3372,
    new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378,
    new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384,
    new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390,
    new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396,
    new_n3397, new_n3398, new_n3399, new_n3400, new_n3401, new_n3402,
    new_n3403, new_n3404, new_n3405, new_n3406, new_n3407, new_n3408,
    new_n3409, new_n3410, new_n3411, new_n3412, new_n3413, new_n3414,
    new_n3415, new_n3416, new_n3417, new_n3418, new_n3419, new_n3420,
    new_n3421, new_n3422, new_n3423, new_n3424, new_n3425, new_n3426,
    new_n3427, new_n3428, new_n3429, new_n3430, new_n3431, new_n3432,
    new_n3433, new_n3434, new_n3435, new_n3436, new_n3437, new_n3438,
    new_n3439, new_n3440, new_n3441, new_n3442, new_n3443, new_n3444,
    new_n3445, new_n3446, new_n3447, new_n3448, new_n3449, new_n3450,
    new_n3451, new_n3452, new_n3453, new_n3454, new_n3455, new_n3456,
    new_n3457, new_n3458, new_n3459, new_n3460, new_n3461, new_n3462,
    new_n3463, new_n3464, new_n3465, new_n3466, new_n3467, new_n3468,
    new_n3469, new_n3470, new_n3471, new_n3472, new_n3473, new_n3474,
    new_n3475, new_n3476, new_n3477, new_n3478, new_n3479, new_n3480,
    new_n3481, new_n3482, new_n3483, new_n3484, new_n3485, new_n3486,
    new_n3487, new_n3488, new_n3489, new_n3490, new_n3491, new_n3492,
    new_n3493, new_n3494, new_n3495, new_n3496, new_n3497, new_n3498,
    new_n3499, new_n3500, new_n3501, new_n3502, new_n3503, new_n3504,
    new_n3505, new_n3506, new_n3507, new_n3508, new_n3509, new_n3510,
    new_n3511, new_n3512, new_n3513, new_n3514, new_n3515, new_n3516,
    new_n3517, new_n3518, new_n3519, new_n3520, new_n3521, new_n3522,
    new_n3523, new_n3524, new_n3525, new_n3526, new_n3527, new_n3528,
    new_n3529, new_n3530, new_n3531, new_n3532, new_n3533, new_n3534,
    new_n3535, new_n3536, new_n3537, new_n3538, new_n3539, new_n3540,
    new_n3541, new_n3542, new_n3543, new_n3544, new_n3545, new_n3546,
    new_n3547, new_n3548, new_n3549, new_n3550, new_n3551, new_n3552,
    new_n3553, new_n3554, new_n3555, new_n3556, new_n3557, new_n3558,
    new_n3559, new_n3560, new_n3561, new_n3562, new_n3563, new_n3564,
    new_n3565, new_n3566, new_n3567, new_n3568, new_n3569, new_n3570,
    new_n3571, new_n3572, new_n3573, new_n3574, new_n3575, new_n3576,
    new_n3577, new_n3578, new_n3579, new_n3580, new_n3581, new_n3582,
    new_n3583, new_n3584, new_n3585, new_n3586, new_n3587, new_n3588,
    new_n3589, new_n3590, new_n3591, new_n3592, new_n3593, new_n3594,
    new_n3595, new_n3596, new_n3597, new_n3598, new_n3599, new_n3600,
    new_n3601, new_n3602, new_n3603, new_n3604, new_n3605, new_n3606,
    new_n3607, new_n3608, new_n3609, new_n3610, new_n3611, new_n3612,
    new_n3613, new_n3614, new_n3615, new_n3616, new_n3617, new_n3618,
    new_n3619, new_n3620, new_n3621, new_n3622, new_n3623, new_n3624,
    new_n3625, new_n3626, new_n3627, new_n3628, new_n3629, new_n3630,
    new_n3631, new_n3632, new_n3633, new_n3634, new_n3635, new_n3636,
    new_n3637, new_n3638, new_n3639, new_n3640, new_n3641, new_n3642,
    new_n3643, new_n3644, new_n3645, new_n3646, new_n3647, new_n3648,
    new_n3649, new_n3650, new_n3651, new_n3652, new_n3653, new_n3654,
    new_n3655, new_n3656, new_n3657, new_n3658, new_n3659, new_n3660,
    new_n3661, new_n3662, new_n3663, new_n3664, new_n3665, new_n3666,
    new_n3667, new_n3668, new_n3669, new_n3670, new_n3671, new_n3672,
    new_n3673, new_n3674, new_n3675, new_n3676, new_n3677, new_n3678,
    new_n3679, new_n3680, new_n3681, new_n3682, new_n3683, new_n3684,
    new_n3685, new_n3686, new_n3687, new_n3688, new_n3689, new_n3690,
    new_n3691, new_n3692, new_n3693, new_n3694, new_n3695, new_n3696,
    new_n3697, new_n3698, new_n3699, new_n3700, new_n3701, new_n3702,
    new_n3703, new_n3704, new_n3705, new_n3706, new_n3707, new_n3708,
    new_n3709, new_n3710, new_n3711, new_n3712, new_n3713, new_n3714,
    new_n3715, new_n3716, new_n3717, new_n3718, new_n3719, new_n3720,
    new_n3721, new_n3722, new_n3723, new_n3724, new_n3725, new_n3726,
    new_n3727, new_n3728, new_n3729, new_n3730, new_n3731, new_n3732,
    new_n3733, new_n3734, new_n3735, new_n3736, new_n3737, new_n3738,
    new_n3739, new_n3740, new_n3741, new_n3742, new_n3743, new_n3744,
    new_n3745, new_n3746, new_n3747, new_n3748, new_n3749, new_n3750,
    new_n3751, new_n3752, new_n3753, new_n3754, new_n3755, new_n3756,
    new_n3757, new_n3758, new_n3759, new_n3760, new_n3761, new_n3762,
    new_n3763, new_n3764, new_n3765, new_n3766, new_n3767, new_n3768,
    new_n3769, new_n3770, new_n3771, new_n3772, new_n3773, new_n3774,
    new_n3775, new_n3776, new_n3777, new_n3778, new_n3779, new_n3780,
    new_n3781, new_n3782, new_n3783, new_n3784, new_n3785, new_n3786,
    new_n3787, new_n3788, new_n3789, new_n3790, new_n3791, new_n3792,
    new_n3793, new_n3794, new_n3795, new_n3796, new_n3797, new_n3798,
    new_n3799, new_n3800, new_n3801, new_n3802, new_n3803, new_n3804,
    new_n3805, new_n3806, new_n3807, new_n3808, new_n3809, new_n3810,
    new_n3811, new_n3812, new_n3813, new_n3814, new_n3815, new_n3816,
    new_n3817, new_n3818, new_n3819, new_n3820, new_n3821, new_n3822,
    new_n3823, new_n3824, new_n3825, new_n3826, new_n3827, new_n3828,
    new_n3829, new_n3830, new_n3831, new_n3832, new_n3833, new_n3834,
    new_n3835, new_n3836, new_n3837, new_n3838, new_n3839, new_n3840,
    new_n3841, new_n3842, new_n3843, new_n3844, new_n3845, new_n3846,
    new_n3847, new_n3848, new_n3849, new_n3850, new_n3851, new_n3852,
    new_n3853, new_n3854, new_n3855, new_n3856, new_n3857, new_n3858,
    new_n3859, new_n3860, new_n3861, new_n3862, new_n3863, new_n3864,
    new_n3865, new_n3866, new_n3867, new_n3868, new_n3869, new_n3870,
    new_n3871, new_n3872, new_n3873, new_n3874, new_n3875, new_n3876,
    new_n3877, new_n3878, new_n3879, new_n3880, new_n3881, new_n3882,
    new_n3883, new_n3884, new_n3885, new_n3886, new_n3887, new_n3888,
    new_n3889, new_n3890, new_n3891, new_n3892, new_n3893, new_n3894,
    new_n3895, new_n3896, new_n3897, new_n3898, new_n3899, new_n3900,
    new_n3901, new_n3902, new_n3903, new_n3904, new_n3905, new_n3906,
    new_n3907, new_n3908, new_n3909, new_n3910, new_n3911, new_n3912,
    new_n3913, new_n3914, new_n3915, new_n3916, new_n3917, new_n3918,
    new_n3919, new_n3920, new_n3921, new_n3922, new_n3923, new_n3924,
    new_n3925, new_n3926, new_n3927, new_n3928, new_n3929, new_n3930,
    new_n3931, new_n3932, new_n3933, new_n3934, new_n3935, new_n3936,
    new_n3937, new_n3938, new_n3939, new_n3940, new_n3941, new_n3942,
    new_n3943, new_n3944, new_n3945, new_n3946, new_n3947, new_n3948,
    new_n3949, new_n3950, new_n3951, new_n3952, new_n3953, new_n3954,
    new_n3955, new_n3956, new_n3957, new_n3958, new_n3959, new_n3960,
    new_n3961, new_n3962, new_n3963, new_n3964, new_n3965, new_n3966,
    new_n3967, new_n3968, new_n3969, new_n3970, new_n3971, new_n3972,
    new_n3973, new_n3974, new_n3975, new_n3976, new_n3977, new_n3978,
    new_n3979, new_n3980, new_n3981, new_n3982, new_n3983, new_n3984,
    new_n3985, new_n3986, new_n3987, new_n3988, new_n3989, new_n3990,
    new_n3991, new_n3992, new_n3993, new_n3994, new_n3995, new_n3996,
    new_n3997, new_n3998, new_n3999, new_n4000, new_n4001, new_n4002,
    new_n4003, new_n4004, new_n4005, new_n4006, new_n4007, new_n4008,
    new_n4009, new_n4010, new_n4011, new_n4012, new_n4013, new_n4014,
    new_n4015, new_n4016, new_n4017, new_n4018, new_n4019, new_n4020,
    new_n4021, new_n4022, new_n4023, new_n4024, new_n4025, new_n4026,
    new_n4027, new_n4028, new_n4029, new_n4030, new_n4031, new_n4032,
    new_n4033, new_n4034, new_n4035, new_n4036, new_n4037, new_n4038,
    new_n4039, new_n4040, new_n4041, new_n4042, new_n4043, new_n4044,
    new_n4045, new_n4046, new_n4047, new_n4048, new_n4049, new_n4050,
    new_n4051, new_n4052, new_n4053, new_n4054, new_n4055, new_n4056,
    new_n4057, new_n4058, new_n4059, new_n4060, new_n4061, new_n4062,
    new_n4063, new_n4064, new_n4065, new_n4066, new_n4067, new_n4068,
    new_n4069, new_n4070, new_n4071, new_n4072, new_n4073, new_n4074,
    new_n4075, new_n4076, new_n4077, new_n4078, new_n4079, new_n4080,
    new_n4081, new_n4082, new_n4083, new_n4084, new_n4085, new_n4086,
    new_n4087, new_n4088, new_n4089, new_n4090, new_n4091, new_n4092,
    new_n4093, new_n4094, new_n4095, new_n4096, new_n4097, new_n4098,
    new_n4099, new_n4100, new_n4101, new_n4102, new_n4103, new_n4104,
    new_n4105, new_n4106, new_n4107, new_n4108, new_n4109, new_n4110,
    new_n4111, new_n4112, new_n4113, new_n4114, new_n4115, new_n4116,
    new_n4117, new_n4118, new_n4119, new_n4120, new_n4121, new_n4122,
    new_n4123, new_n4124, new_n4125, new_n4126, new_n4127, new_n4128,
    new_n4129, new_n4130, new_n4131, new_n4132, new_n4133, new_n4134,
    new_n4135, new_n4136, new_n4137, new_n4138, new_n4139, new_n4140,
    new_n4141, new_n4142, new_n4143, new_n4144, new_n4145, new_n4146,
    new_n4147, new_n4148, new_n4149, new_n4150, new_n4151, new_n4152,
    new_n4153, new_n4154, new_n4155, new_n4156, new_n4157, new_n4158,
    new_n4159, new_n4160, new_n4161, new_n4162, new_n4163, new_n4164,
    new_n4165, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170,
    new_n4171, new_n4172, new_n4173, new_n4174, new_n4175, new_n4176,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200,
    new_n4201, new_n4202, new_n4203, new_n4204, new_n4205, new_n4206,
    new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221, new_n4222, new_n4223, new_n4224,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230,
    new_n4231, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254,
    new_n4255, new_n4256, new_n4257, new_n4258, new_n4259, new_n4260,
    new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266,
    new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272,
    new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278,
    new_n4279, new_n4280, new_n4281, new_n4282, new_n4283, new_n4284,
    new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290,
    new_n4291, new_n4292, new_n4293, new_n4294, new_n4295, new_n4296,
    new_n4297, new_n4298, new_n4299, new_n4300, new_n4301, new_n4302,
    new_n4303, new_n4304, new_n4305, new_n4306, new_n4307, new_n4308,
    new_n4309, new_n4310, new_n4311, new_n4312, new_n4313, new_n4314,
    new_n4315, new_n4316, new_n4317, new_n4318, new_n4319, new_n4320,
    new_n4321, new_n4322, new_n4323, new_n4324, new_n4325, new_n4326,
    new_n4327, new_n4328, new_n4329, new_n4330, new_n4331, new_n4332,
    new_n4333, new_n4334, new_n4335, new_n4336, new_n4337, new_n4338,
    new_n4339, new_n4340, new_n4341, new_n4342, new_n4343, new_n4344,
    new_n4345, new_n4346, new_n4347, new_n4348, new_n4349, new_n4350,
    new_n4351, new_n4352, new_n4353, new_n4354, new_n4355, new_n4356,
    new_n4357, new_n4358, new_n4359, new_n4360, new_n4361, new_n4362,
    new_n4363, new_n4364, new_n4365, new_n4366, new_n4367, new_n4368,
    new_n4369, new_n4370, new_n4371, new_n4372, new_n4373, new_n4374,
    new_n4375, new_n4376, new_n4377, new_n4378, new_n4379, new_n4380,
    new_n4381, new_n4382, new_n4383, new_n4384, new_n4385, new_n4386,
    new_n4387, new_n4388, new_n4389, new_n4390, new_n4391, new_n4392,
    new_n4393, new_n4394, new_n4395, new_n4396, new_n4397, new_n4398,
    new_n4399, new_n4400, new_n4401, new_n4402, new_n4403, new_n4404,
    new_n4405, new_n4406, new_n4407, new_n4408, new_n4409, new_n4410,
    new_n4411, new_n4412, new_n4413, new_n4414, new_n4415, new_n4416,
    new_n4417, new_n4418, new_n4419, new_n4420, new_n4421, new_n4422,
    new_n4423, new_n4424, new_n4425, new_n4426, new_n4427, new_n4428,
    new_n4429, new_n4430, new_n4431, new_n4432, new_n4433, new_n4434,
    new_n4435, new_n4436, new_n4437, new_n4438, new_n4439, new_n4440,
    new_n4441, new_n4442, new_n4443, new_n4444, new_n4445, new_n4446,
    new_n4447, new_n4448, new_n4449, new_n4450, new_n4451, new_n4452,
    new_n4453, new_n4454, new_n4455, new_n4456, new_n4457, new_n4458,
    new_n4459, new_n4460, new_n4461, new_n4462, new_n4463, new_n4464,
    new_n4465, new_n4466, new_n4467, new_n4468, new_n4469, new_n4470,
    new_n4471, new_n4472, new_n4473, new_n4474, new_n4475, new_n4476,
    new_n4477, new_n4478, new_n4479, new_n4480, new_n4481, new_n4482,
    new_n4483, new_n4484, new_n4485, new_n4486, new_n4487, new_n4488,
    new_n4489, new_n4490, new_n4491, new_n4492, new_n4493, new_n4494,
    new_n4495, new_n4496, new_n4497, new_n4498, new_n4499, new_n4500,
    new_n4501, new_n4502, new_n4503, new_n4504, new_n4505, new_n4506,
    new_n4507, new_n4508, new_n4509, new_n4510, new_n4511, new_n4512,
    new_n4513, new_n4514, new_n4515, new_n4516, new_n4517, new_n4518,
    new_n4519, new_n4520, new_n4521, new_n4522, new_n4523, new_n4524,
    new_n4525, new_n4526, new_n4527, new_n4528, new_n4529, new_n4530,
    new_n4531, new_n4532, new_n4533, new_n4534, new_n4535, new_n4536,
    new_n4537, new_n4538, new_n4539, new_n4540, new_n4541, new_n4542,
    new_n4543, new_n4544, new_n4545, new_n4546, new_n4547, new_n4548,
    new_n4549, new_n4550, new_n4551, new_n4552, new_n4553, new_n4554,
    new_n4555, new_n4556, new_n4557, new_n4558, new_n4559, new_n4560,
    new_n4561, new_n4562, new_n4563, new_n4564, new_n4565, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4574, new_n4575, new_n4576, new_n4577, new_n4578,
    new_n4579, new_n4580, new_n4581, new_n4582, new_n4583, new_n4584,
    new_n4585, new_n4586, new_n4587, new_n4588, new_n4589, new_n4590,
    new_n4591, new_n4592, new_n4593, new_n4594, new_n4595, new_n4596,
    new_n4597, new_n4598, new_n4599, new_n4600, new_n4601, new_n4602,
    new_n4603, new_n4604, new_n4605, new_n4606, new_n4607, new_n4608,
    new_n4609, new_n4610, new_n4611, new_n4612, new_n4613, new_n4614,
    new_n4615, new_n4616, new_n4617, new_n4618, new_n4619, new_n4620,
    new_n4621, new_n4622, new_n4623, new_n4624, new_n4625, new_n4626,
    new_n4627, new_n4628, new_n4629, new_n4630, new_n4631, new_n4632,
    new_n4633, new_n4634, new_n4635, new_n4636, new_n4637, new_n4638,
    new_n4639, new_n4640, new_n4641, new_n4642, new_n4643, new_n4644,
    new_n4645, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650,
    new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656,
    new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662,
    new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668,
    new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674,
    new_n4675, new_n4676, new_n4677, new_n4678, new_n4679, new_n4680,
    new_n4681, new_n4682, new_n4683, new_n4684, new_n4685, new_n4686,
    new_n4687, new_n4688, new_n4689, new_n4690, new_n4691, new_n4692,
    new_n4693, new_n4694, new_n4695, new_n4696, new_n4697, new_n4698,
    new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704,
    new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710,
    new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716,
    new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722,
    new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728,
    new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743, new_n4744, new_n4745, new_n4746,
    new_n4747, new_n4748, new_n4749, new_n4750, new_n4751, new_n4752,
    new_n4753, new_n4754, new_n4755, new_n4756, new_n4757, new_n4758,
    new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764,
    new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770,
    new_n4771, new_n4772, new_n4773, new_n4774, new_n4775, new_n4776,
    new_n4777, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782,
    new_n4783, new_n4784, new_n4785, new_n4786, new_n4787, new_n4788,
    new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794,
    new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800,
    new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806,
    new_n4807, new_n4808, new_n4809, new_n4810, new_n4811, new_n4812,
    new_n4813, new_n4814, new_n4815, new_n4816, new_n4817, new_n4818,
    new_n4819, new_n4820, new_n4821, new_n4822, new_n4823, new_n4824,
    new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4830,
    new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836,
    new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842,
    new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848,
    new_n4849, new_n4850, new_n4851, new_n4852, new_n4853, new_n4854,
    new_n4855, new_n4856, new_n4857, new_n4858, new_n4859, new_n4860,
    new_n4861, new_n4862, new_n4863, new_n4864, new_n4865, new_n4866,
    new_n4867, new_n4868, new_n4869, new_n4870, new_n4871, new_n4872,
    new_n4873, new_n4874, new_n4875, new_n4876, new_n4877, new_n4878,
    new_n4879, new_n4880, new_n4881, new_n4882, new_n4883, new_n4884,
    new_n4885, new_n4886, new_n4887, new_n4888, new_n4889, new_n4890,
    new_n4891, new_n4892, new_n4893, new_n4894, new_n4895, new_n4896,
    new_n4897, new_n4898, new_n4899, new_n4900, new_n4901, new_n4902,
    new_n4903, new_n4904, new_n4905, new_n4906, new_n4907, new_n4908,
    new_n4909, new_n4910, new_n4911, new_n4912, new_n4913, new_n4914,
    new_n4915, new_n4916, new_n4917, new_n4918, new_n4919, new_n4920,
    new_n4921, new_n4922, new_n4923, new_n4924, new_n4925, new_n4926,
    new_n4927, new_n4928;
  assign new_n577 = n481 ^ n225;
  assign new_n578 = n290 ^ n34;
  assign new_n579 = new_n578 ^ new_n577;
  assign new_n580 = n461 ^ n205;
  assign new_n581 = n332 ^ n76;
  assign new_n582 = new_n581 ^ new_n580;
  assign new_n583 = n398 ^ n142;
  assign new_n584 = new_n583 ^ n13;
  assign new_n585 = ~new_n584 & new_n582;
  assign new_n586 = new_n585 ^ new_n579;
  assign new_n587 = n482 ^ n226;
  assign new_n588 = n291 ^ n35;
  assign new_n589 = new_n588 ^ new_n587;
  assign new_n590 = n462 ^ n206;
  assign new_n591 = n333 ^ n77;
  assign new_n592 = new_n591 ^ new_n590;
  assign new_n593 = n399 ^ n143;
  assign new_n594 = new_n593 ^ n14;
  assign new_n595 = ~new_n594 & new_n592;
  assign new_n596 = new_n595 ^ new_n589;
  assign new_n597 = n483 ^ n227;
  assign new_n598 = n292 ^ n36;
  assign new_n599 = new_n598 ^ new_n597;
  assign new_n600 = n463 ^ n207;
  assign new_n601 = n334 ^ n78;
  assign new_n602 = new_n601 ^ new_n600;
  assign new_n603 = n400 ^ n144;
  assign new_n604 = new_n603 ^ n15;
  assign new_n605 = ~new_n604 & new_n602;
  assign new_n606 = new_n605 ^ new_n599;
  assign new_n607 = n484 ^ n228;
  assign new_n608 = n293 ^ n37;
  assign new_n609 = new_n608 ^ new_n607;
  assign new_n610 = n464 ^ n208;
  assign new_n611 = n335 ^ n79;
  assign new_n612 = new_n611 ^ new_n610;
  assign new_n613 = n401 ^ n145;
  assign new_n614 = new_n613 ^ n16;
  assign new_n615 = ~new_n614 & new_n612;
  assign new_n616 = new_n615 ^ new_n609;
  assign new_n617 = n485 ^ n229;
  assign new_n618 = n294 ^ n38;
  assign new_n619 = new_n618 ^ new_n617;
  assign new_n620 = n465 ^ n209;
  assign new_n621 = n336 ^ n80;
  assign new_n622 = new_n621 ^ new_n620;
  assign new_n623 = n402 ^ n146;
  assign new_n624 = new_n623 ^ n17;
  assign new_n625 = ~new_n624 & new_n622;
  assign new_n626 = new_n625 ^ new_n619;
  assign new_n627 = n486 ^ n230;
  assign new_n628 = n295 ^ n39;
  assign new_n629 = new_n628 ^ new_n627;
  assign new_n630 = n466 ^ n210;
  assign new_n631 = n337 ^ n81;
  assign new_n632 = new_n631 ^ new_n630;
  assign new_n633 = n403 ^ n147;
  assign new_n634 = new_n633 ^ n18;
  assign new_n635 = ~new_n634 & new_n632;
  assign new_n636 = new_n635 ^ new_n629;
  assign new_n637 = n487 ^ n231;
  assign new_n638 = n296 ^ n40;
  assign new_n639 = new_n638 ^ new_n637;
  assign new_n640 = n467 ^ n211;
  assign new_n641 = n338 ^ n82;
  assign new_n642 = new_n641 ^ new_n640;
  assign new_n643 = n404 ^ n148;
  assign new_n644 = new_n643 ^ n19;
  assign new_n645 = ~new_n644 & new_n642;
  assign new_n646 = new_n645 ^ new_n639;
  assign new_n647 = n488 ^ n232;
  assign new_n648 = n297 ^ n41;
  assign new_n649 = new_n648 ^ new_n647;
  assign new_n650 = n468 ^ n212;
  assign new_n651 = n339 ^ n83;
  assign new_n652 = new_n651 ^ new_n650;
  assign new_n653 = n405 ^ n149;
  assign new_n654 = new_n653 ^ n20;
  assign new_n655 = ~new_n654 & new_n652;
  assign new_n656 = new_n655 ^ new_n649;
  assign new_n657 = n489 ^ n233;
  assign new_n658 = n298 ^ n42;
  assign new_n659 = new_n658 ^ new_n657;
  assign new_n660 = n469 ^ n213;
  assign new_n661 = n340 ^ n84;
  assign new_n662 = new_n661 ^ new_n660;
  assign new_n663 = n406 ^ n150;
  assign new_n664 = new_n663 ^ n21;
  assign new_n665 = ~new_n664 & new_n662;
  assign new_n666 = new_n665 ^ new_n659;
  assign new_n667 = n490 ^ n234;
  assign new_n668 = n299 ^ n43;
  assign new_n669 = new_n668 ^ new_n667;
  assign new_n670 = n470 ^ n214;
  assign new_n671 = n341 ^ n85;
  assign new_n672 = new_n671 ^ new_n670;
  assign new_n673 = n407 ^ n151;
  assign new_n674 = new_n673 ^ n22;
  assign new_n675 = ~new_n674 & new_n672;
  assign new_n676 = new_n675 ^ new_n669;
  assign new_n677 = n491 ^ n235;
  assign new_n678 = n300 ^ n44;
  assign new_n679 = new_n678 ^ new_n677;
  assign new_n680 = n471 ^ n215;
  assign new_n681 = n342 ^ n86;
  assign new_n682 = new_n681 ^ new_n680;
  assign new_n683 = n408 ^ n152;
  assign new_n684 = new_n683 ^ n23;
  assign new_n685 = ~new_n684 & new_n682;
  assign new_n686 = new_n685 ^ new_n679;
  assign new_n687 = n492 ^ n236;
  assign new_n688 = n301 ^ n45;
  assign new_n689 = new_n688 ^ new_n687;
  assign new_n690 = n472 ^ n216;
  assign new_n691 = n343 ^ n87;
  assign new_n692 = new_n691 ^ new_n690;
  assign new_n693 = n409 ^ n153;
  assign new_n694 = new_n693 ^ n24;
  assign new_n695 = ~new_n694 & new_n692;
  assign new_n696 = new_n695 ^ new_n689;
  assign new_n697 = n493 ^ n237;
  assign new_n698 = n302 ^ n46;
  assign new_n699 = new_n698 ^ new_n697;
  assign new_n700 = n473 ^ n217;
  assign new_n701 = n344 ^ n88;
  assign new_n702 = new_n701 ^ new_n700;
  assign new_n703 = n410 ^ n154;
  assign new_n704 = new_n703 ^ n25;
  assign new_n705 = ~new_n704 & new_n702;
  assign new_n706 = new_n705 ^ new_n699;
  assign new_n707 = n494 ^ n238;
  assign new_n708 = n303 ^ n47;
  assign new_n709 = new_n708 ^ new_n707;
  assign new_n710 = n474 ^ n218;
  assign new_n711 = n345 ^ n89;
  assign new_n712 = new_n711 ^ new_n710;
  assign new_n713 = n411 ^ n155;
  assign new_n714 = new_n713 ^ n26;
  assign new_n715 = ~new_n714 & new_n712;
  assign new_n716 = new_n715 ^ new_n709;
  assign new_n717 = n495 ^ n239;
  assign new_n718 = n304 ^ n48;
  assign new_n719 = new_n718 ^ new_n717;
  assign new_n720 = n475 ^ n219;
  assign new_n721 = n346 ^ n90;
  assign new_n722 = new_n721 ^ new_n720;
  assign new_n723 = n412 ^ n156;
  assign new_n724 = new_n723 ^ n27;
  assign new_n725 = ~new_n724 & new_n722;
  assign new_n726 = new_n725 ^ new_n719;
  assign new_n727 = n496 ^ n240;
  assign new_n728 = n305 ^ n49;
  assign new_n729 = new_n728 ^ new_n727;
  assign new_n730 = n476 ^ n220;
  assign new_n731 = n347 ^ n91;
  assign new_n732 = new_n731 ^ new_n730;
  assign new_n733 = n413 ^ n157;
  assign new_n734 = new_n733 ^ n28;
  assign new_n735 = ~new_n734 & new_n732;
  assign new_n736 = new_n735 ^ new_n729;
  assign new_n737 = n497 ^ n241;
  assign new_n738 = n306 ^ n50;
  assign new_n739 = new_n738 ^ new_n737;
  assign new_n740 = n477 ^ n221;
  assign new_n741 = n348 ^ n92;
  assign new_n742 = new_n741 ^ new_n740;
  assign new_n743 = n414 ^ n158;
  assign new_n744 = new_n743 ^ n29;
  assign new_n745 = ~new_n744 & new_n742;
  assign new_n746 = new_n745 ^ new_n739;
  assign new_n747 = n498 ^ n242;
  assign new_n748 = n307 ^ n51;
  assign new_n749 = new_n748 ^ new_n747;
  assign new_n750 = n478 ^ n222;
  assign new_n751 = n349 ^ n93;
  assign new_n752 = new_n751 ^ new_n750;
  assign new_n753 = n415 ^ n159;
  assign new_n754 = new_n753 ^ n30;
  assign new_n755 = ~new_n754 & new_n752;
  assign new_n756 = new_n755 ^ new_n749;
  assign new_n757 = n499 ^ n243;
  assign new_n758 = n308 ^ n52;
  assign new_n759 = new_n758 ^ new_n757;
  assign new_n760 = n479 ^ n223;
  assign new_n761 = n350 ^ n94;
  assign new_n762 = new_n761 ^ new_n760;
  assign new_n763 = n416 ^ n160;
  assign new_n764 = new_n763 ^ n31;
  assign new_n765 = ~new_n764 & new_n762;
  assign new_n766 = new_n765 ^ new_n759;
  assign new_n767 = n500 ^ n244;
  assign new_n768 = n309 ^ n53;
  assign new_n769 = new_n768 ^ new_n767;
  assign new_n770 = n480 ^ n224;
  assign new_n771 = n351 ^ n95;
  assign new_n772 = new_n771 ^ new_n770;
  assign new_n773 = n353 ^ n97;
  assign new_n774 = new_n773 ^ n32;
  assign new_n775 = ~new_n774 & new_n772;
  assign new_n776 = new_n775 ^ new_n769;
  assign new_n777 = n310 ^ n54;
  assign new_n778 = n501 ^ n245;
  assign new_n779 = new_n778 ^ new_n777;
  assign new_n780 = n417 ^ n161;
  assign new_n781 = n352 ^ n96;
  assign new_n782 = new_n781 ^ new_n780;
  assign new_n783 = n354 ^ n98;
  assign new_n784 = new_n783 ^ n545;
  assign new_n785 = ~new_n784 & new_n782;
  assign new_n786 = new_n785 ^ new_n779;
  assign new_n787 = n311 ^ n55;
  assign new_n788 = n502 ^ n246;
  assign new_n789 = new_n788 ^ new_n787;
  assign new_n790 = n418 ^ n162;
  assign new_n791 = n289 ^ n33;
  assign new_n792 = new_n791 ^ new_n790;
  assign new_n793 = n355 ^ n99;
  assign new_n794 = new_n793 ^ n546;
  assign new_n795 = ~new_n794 & new_n792;
  assign new_n796 = new_n795 ^ new_n789;
  assign new_n797 = n312 ^ n56;
  assign new_n798 = n503 ^ n247;
  assign new_n799 = new_n798 ^ new_n797;
  assign new_n800 = n419 ^ n163;
  assign new_n801 = new_n800 ^ new_n578;
  assign new_n802 = n356 ^ n100;
  assign new_n803 = new_n802 ^ n547;
  assign new_n804 = ~new_n803 & new_n801;
  assign new_n805 = new_n804 ^ new_n799;
  assign new_n806 = n313 ^ n57;
  assign new_n807 = n504 ^ n248;
  assign new_n808 = new_n807 ^ new_n806;
  assign new_n809 = n420 ^ n164;
  assign new_n810 = new_n809 ^ new_n588;
  assign new_n811 = n357 ^ n101;
  assign new_n812 = new_n811 ^ n548;
  assign new_n813 = ~new_n812 & new_n810;
  assign new_n814 = new_n813 ^ new_n808;
  assign new_n815 = n314 ^ n58;
  assign new_n816 = n505 ^ n249;
  assign new_n817 = new_n816 ^ new_n815;
  assign new_n818 = n421 ^ n165;
  assign new_n819 = new_n818 ^ new_n598;
  assign new_n820 = n358 ^ n102;
  assign new_n821 = new_n820 ^ n549;
  assign new_n822 = ~new_n821 & new_n819;
  assign new_n823 = new_n822 ^ new_n817;
  assign new_n824 = n315 ^ n59;
  assign new_n825 = n506 ^ n250;
  assign new_n826 = new_n825 ^ new_n824;
  assign new_n827 = n422 ^ n166;
  assign new_n828 = new_n827 ^ new_n608;
  assign new_n829 = n359 ^ n103;
  assign new_n830 = new_n829 ^ n550;
  assign new_n831 = ~new_n830 & new_n828;
  assign new_n832 = new_n831 ^ new_n826;
  assign new_n833 = n316 ^ n60;
  assign new_n834 = n507 ^ n251;
  assign new_n835 = new_n834 ^ new_n833;
  assign new_n836 = n423 ^ n167;
  assign new_n837 = new_n836 ^ new_n618;
  assign new_n838 = n360 ^ n104;
  assign new_n839 = new_n838 ^ n551;
  assign new_n840 = ~new_n839 & new_n837;
  assign new_n841 = new_n840 ^ new_n835;
  assign new_n842 = n317 ^ n61;
  assign new_n843 = n508 ^ n252;
  assign new_n844 = new_n843 ^ new_n842;
  assign new_n845 = n424 ^ n168;
  assign new_n846 = new_n845 ^ new_n628;
  assign new_n847 = n361 ^ n105;
  assign new_n848 = new_n847 ^ n552;
  assign new_n849 = ~new_n848 & new_n846;
  assign new_n850 = new_n849 ^ new_n844;
  assign new_n851 = n318 ^ n62;
  assign new_n852 = n509 ^ n253;
  assign new_n853 = new_n852 ^ new_n851;
  assign new_n854 = n425 ^ n169;
  assign new_n855 = new_n854 ^ new_n638;
  assign new_n856 = n362 ^ n106;
  assign new_n857 = new_n856 ^ n553;
  assign new_n858 = ~new_n857 & new_n855;
  assign new_n859 = new_n858 ^ new_n853;
  assign new_n860 = n319 ^ n63;
  assign new_n861 = n510 ^ n254;
  assign new_n862 = new_n861 ^ new_n860;
  assign new_n863 = n426 ^ n170;
  assign new_n864 = new_n863 ^ new_n648;
  assign new_n865 = n363 ^ n107;
  assign new_n866 = new_n865 ^ n554;
  assign new_n867 = ~new_n866 & new_n864;
  assign new_n868 = new_n867 ^ new_n862;
  assign new_n869 = n320 ^ n64;
  assign new_n870 = n511 ^ n255;
  assign new_n871 = new_n870 ^ new_n869;
  assign new_n872 = n427 ^ n171;
  assign new_n873 = new_n872 ^ new_n658;
  assign new_n874 = n364 ^ n108;
  assign new_n875 = new_n874 ^ n555;
  assign new_n876 = ~new_n875 & new_n873;
  assign new_n877 = new_n876 ^ new_n871;
  assign new_n878 = n321 ^ n65;
  assign new_n879 = n512 ^ n256;
  assign new_n880 = new_n879 ^ new_n878;
  assign new_n881 = n428 ^ n172;
  assign new_n882 = new_n881 ^ new_n668;
  assign new_n883 = n365 ^ n109;
  assign new_n884 = new_n883 ^ n556;
  assign new_n885 = ~new_n884 & new_n882;
  assign new_n886 = new_n885 ^ new_n880;
  assign new_n887 = n322 ^ n66;
  assign new_n888 = n513 ^ n257;
  assign new_n889 = new_n888 ^ new_n887;
  assign new_n890 = n429 ^ n173;
  assign new_n891 = new_n890 ^ new_n678;
  assign new_n892 = n366 ^ n110;
  assign new_n893 = new_n892 ^ n557;
  assign new_n894 = ~new_n893 & new_n891;
  assign new_n895 = new_n894 ^ new_n889;
  assign new_n896 = n323 ^ n67;
  assign new_n897 = n514 ^ n258;
  assign new_n898 = new_n897 ^ new_n896;
  assign new_n899 = n430 ^ n174;
  assign new_n900 = new_n899 ^ new_n688;
  assign new_n901 = n367 ^ n111;
  assign new_n902 = new_n901 ^ n558;
  assign new_n903 = ~new_n902 & new_n900;
  assign new_n904 = new_n903 ^ new_n898;
  assign new_n905 = n324 ^ n68;
  assign new_n906 = n515 ^ n259;
  assign new_n907 = new_n906 ^ new_n905;
  assign new_n908 = n431 ^ n175;
  assign new_n909 = new_n908 ^ new_n698;
  assign new_n910 = n368 ^ n112;
  assign new_n911 = new_n910 ^ n559;
  assign new_n912 = ~new_n911 & new_n909;
  assign new_n913 = new_n912 ^ new_n907;
  assign new_n914 = n325 ^ n69;
  assign new_n915 = n516 ^ n260;
  assign new_n916 = new_n915 ^ new_n914;
  assign new_n917 = n432 ^ n176;
  assign new_n918 = new_n917 ^ new_n708;
  assign new_n919 = n369 ^ n113;
  assign new_n920 = new_n919 ^ n560;
  assign new_n921 = ~new_n920 & new_n918;
  assign new_n922 = new_n921 ^ new_n916;
  assign new_n923 = n326 ^ n70;
  assign new_n924 = n517 ^ n261;
  assign new_n925 = new_n924 ^ new_n923;
  assign new_n926 = n433 ^ n177;
  assign new_n927 = new_n926 ^ new_n718;
  assign new_n928 = n370 ^ n114;
  assign new_n929 = new_n928 ^ n561;
  assign new_n930 = ~new_n929 & new_n927;
  assign new_n931 = new_n930 ^ new_n925;
  assign new_n932 = n327 ^ n71;
  assign new_n933 = n518 ^ n262;
  assign new_n934 = new_n933 ^ new_n932;
  assign new_n935 = n434 ^ n178;
  assign new_n936 = new_n935 ^ new_n728;
  assign new_n937 = n371 ^ n115;
  assign new_n938 = new_n937 ^ n562;
  assign new_n939 = ~new_n938 & new_n936;
  assign new_n940 = new_n939 ^ new_n934;
  assign new_n941 = n328 ^ n72;
  assign new_n942 = n519 ^ n263;
  assign new_n943 = new_n942 ^ new_n941;
  assign new_n944 = n435 ^ n179;
  assign new_n945 = new_n944 ^ new_n738;
  assign new_n946 = n372 ^ n116;
  assign new_n947 = new_n946 ^ n563;
  assign new_n948 = ~new_n947 & new_n945;
  assign new_n949 = new_n948 ^ new_n943;
  assign new_n950 = n329 ^ n73;
  assign new_n951 = n520 ^ n264;
  assign new_n952 = new_n951 ^ new_n950;
  assign new_n953 = n436 ^ n180;
  assign new_n954 = new_n953 ^ new_n748;
  assign new_n955 = n373 ^ n117;
  assign new_n956 = new_n955 ^ n564;
  assign new_n957 = ~new_n956 & new_n954;
  assign new_n958 = new_n957 ^ new_n952;
  assign new_n959 = n330 ^ n74;
  assign new_n960 = n521 ^ n265;
  assign new_n961 = new_n960 ^ new_n959;
  assign new_n962 = n437 ^ n181;
  assign new_n963 = new_n962 ^ new_n758;
  assign new_n964 = n374 ^ n118;
  assign new_n965 = new_n964 ^ n565;
  assign new_n966 = ~new_n965 & new_n963;
  assign new_n967 = new_n966 ^ new_n961;
  assign new_n968 = n331 ^ n75;
  assign new_n969 = n522 ^ n266;
  assign new_n970 = new_n969 ^ new_n968;
  assign new_n971 = n438 ^ n182;
  assign new_n972 = new_n971 ^ new_n768;
  assign new_n973 = n375 ^ n119;
  assign new_n974 = new_n973 ^ n566;
  assign new_n975 = ~new_n974 & new_n972;
  assign new_n976 = new_n975 ^ new_n970;
  assign new_n977 = n523 ^ n267;
  assign new_n978 = new_n977 ^ new_n581;
  assign new_n979 = n439 ^ n183;
  assign new_n980 = new_n979 ^ new_n777;
  assign new_n981 = n376 ^ n120;
  assign new_n982 = new_n981 ^ n567;
  assign new_n983 = ~new_n982 & new_n980;
  assign new_n984 = new_n983 ^ new_n978;
  assign new_n985 = n524 ^ n268;
  assign new_n986 = new_n985 ^ new_n591;
  assign new_n987 = n440 ^ n184;
  assign new_n988 = new_n987 ^ new_n787;
  assign new_n989 = n377 ^ n121;
  assign new_n990 = new_n989 ^ n568;
  assign new_n991 = ~new_n990 & new_n988;
  assign new_n992 = new_n991 ^ new_n986;
  assign new_n993 = n525 ^ n269;
  assign new_n994 = new_n993 ^ new_n601;
  assign new_n995 = n441 ^ n185;
  assign new_n996 = new_n995 ^ new_n797;
  assign new_n997 = n378 ^ n122;
  assign new_n998 = new_n997 ^ n569;
  assign new_n999 = ~new_n998 & new_n996;
  assign new_n1000 = new_n999 ^ new_n994;
  assign new_n1001 = n526 ^ n270;
  assign new_n1002 = new_n1001 ^ new_n611;
  assign new_n1003 = n442 ^ n186;
  assign new_n1004 = new_n1003 ^ new_n806;
  assign new_n1005 = n379 ^ n123;
  assign new_n1006 = new_n1005 ^ n570;
  assign new_n1007 = ~new_n1006 & new_n1004;
  assign new_n1008 = new_n1007 ^ new_n1002;
  assign new_n1009 = n527 ^ n271;
  assign new_n1010 = new_n1009 ^ new_n621;
  assign new_n1011 = n443 ^ n187;
  assign new_n1012 = new_n1011 ^ new_n815;
  assign new_n1013 = n380 ^ n124;
  assign new_n1014 = new_n1013 ^ n571;
  assign new_n1015 = ~new_n1014 & new_n1012;
  assign new_n1016 = new_n1015 ^ new_n1010;
  assign new_n1017 = n528 ^ n272;
  assign new_n1018 = new_n1017 ^ new_n631;
  assign new_n1019 = n444 ^ n188;
  assign new_n1020 = new_n1019 ^ new_n824;
  assign new_n1021 = n381 ^ n125;
  assign new_n1022 = new_n1021 ^ n572;
  assign new_n1023 = ~new_n1022 & new_n1020;
  assign new_n1024 = new_n1023 ^ new_n1018;
  assign new_n1025 = n529 ^ n273;
  assign new_n1026 = new_n1025 ^ new_n641;
  assign new_n1027 = n445 ^ n189;
  assign new_n1028 = new_n1027 ^ new_n833;
  assign new_n1029 = n382 ^ n126;
  assign new_n1030 = new_n1029 ^ n573;
  assign new_n1031 = ~new_n1030 & new_n1028;
  assign new_n1032 = new_n1031 ^ new_n1026;
  assign new_n1033 = n530 ^ n274;
  assign new_n1034 = new_n1033 ^ new_n651;
  assign new_n1035 = n446 ^ n190;
  assign new_n1036 = new_n1035 ^ new_n842;
  assign new_n1037 = n383 ^ n127;
  assign new_n1038 = new_n1037 ^ n574;
  assign new_n1039 = ~new_n1038 & new_n1036;
  assign new_n1040 = new_n1039 ^ new_n1034;
  assign new_n1041 = n531 ^ n275;
  assign new_n1042 = new_n1041 ^ new_n661;
  assign new_n1043 = n447 ^ n191;
  assign new_n1044 = new_n1043 ^ new_n851;
  assign new_n1045 = n384 ^ n128;
  assign new_n1046 = new_n1045 ^ n575;
  assign new_n1047 = ~new_n1046 & new_n1044;
  assign new_n1048 = new_n1047 ^ new_n1042;
  assign new_n1049 = n532 ^ n276;
  assign new_n1050 = new_n1049 ^ new_n671;
  assign new_n1051 = n448 ^ n192;
  assign new_n1052 = new_n1051 ^ new_n860;
  assign new_n1053 = n385 ^ n129;
  assign new_n1054 = new_n1053 ^ n576;
  assign new_n1055 = ~new_n1054 & new_n1052;
  assign new_n1056 = new_n1055 ^ new_n1050;
  assign new_n1057 = n533 ^ n277;
  assign new_n1058 = new_n1057 ^ new_n681;
  assign new_n1059 = n449 ^ n193;
  assign new_n1060 = new_n1059 ^ new_n869;
  assign new_n1061 = n386 ^ n130;
  assign new_n1062 = new_n1061 ^ n1;
  assign new_n1063 = ~new_n1062 & new_n1060;
  assign new_n1064 = new_n1063 ^ new_n1058;
  assign new_n1065 = n534 ^ n278;
  assign new_n1066 = new_n1065 ^ new_n691;
  assign new_n1067 = n450 ^ n194;
  assign new_n1068 = new_n1067 ^ new_n878;
  assign new_n1069 = n387 ^ n131;
  assign new_n1070 = new_n1069 ^ n2;
  assign new_n1071 = ~new_n1070 & new_n1068;
  assign new_n1072 = new_n1071 ^ new_n1066;
  assign new_n1073 = n535 ^ n279;
  assign new_n1074 = new_n1073 ^ new_n701;
  assign new_n1075 = n451 ^ n195;
  assign new_n1076 = new_n1075 ^ new_n887;
  assign new_n1077 = n388 ^ n132;
  assign new_n1078 = new_n1077 ^ n3;
  assign new_n1079 = ~new_n1078 & new_n1076;
  assign new_n1080 = new_n1079 ^ new_n1074;
  assign new_n1081 = n536 ^ n280;
  assign new_n1082 = new_n1081 ^ new_n711;
  assign new_n1083 = n452 ^ n196;
  assign new_n1084 = new_n1083 ^ new_n896;
  assign new_n1085 = n389 ^ n133;
  assign new_n1086 = new_n1085 ^ n4;
  assign new_n1087 = ~new_n1086 & new_n1084;
  assign new_n1088 = new_n1087 ^ new_n1082;
  assign new_n1089 = n537 ^ n281;
  assign new_n1090 = new_n1089 ^ new_n721;
  assign new_n1091 = n453 ^ n197;
  assign new_n1092 = new_n1091 ^ new_n905;
  assign new_n1093 = n390 ^ n134;
  assign new_n1094 = new_n1093 ^ n5;
  assign new_n1095 = ~new_n1094 & new_n1092;
  assign new_n1096 = new_n1095 ^ new_n1090;
  assign new_n1097 = n538 ^ n282;
  assign new_n1098 = new_n1097 ^ new_n731;
  assign new_n1099 = n454 ^ n198;
  assign new_n1100 = new_n1099 ^ new_n914;
  assign new_n1101 = n391 ^ n135;
  assign new_n1102 = new_n1101 ^ n6;
  assign new_n1103 = ~new_n1102 & new_n1100;
  assign new_n1104 = new_n1103 ^ new_n1098;
  assign new_n1105 = n539 ^ n283;
  assign new_n1106 = new_n1105 ^ new_n741;
  assign new_n1107 = n455 ^ n199;
  assign new_n1108 = new_n1107 ^ new_n923;
  assign new_n1109 = n392 ^ n136;
  assign new_n1110 = new_n1109 ^ n7;
  assign new_n1111 = ~new_n1110 & new_n1108;
  assign new_n1112 = new_n1111 ^ new_n1106;
  assign new_n1113 = n540 ^ n284;
  assign new_n1114 = new_n1113 ^ new_n751;
  assign new_n1115 = n456 ^ n200;
  assign new_n1116 = new_n1115 ^ new_n932;
  assign new_n1117 = n393 ^ n137;
  assign new_n1118 = new_n1117 ^ n8;
  assign new_n1119 = ~new_n1118 & new_n1116;
  assign new_n1120 = new_n1119 ^ new_n1114;
  assign new_n1121 = n541 ^ n285;
  assign new_n1122 = new_n1121 ^ new_n761;
  assign new_n1123 = n457 ^ n201;
  assign new_n1124 = new_n1123 ^ new_n941;
  assign new_n1125 = n394 ^ n138;
  assign new_n1126 = new_n1125 ^ n9;
  assign new_n1127 = ~new_n1126 & new_n1124;
  assign new_n1128 = new_n1127 ^ new_n1122;
  assign new_n1129 = n542 ^ n286;
  assign new_n1130 = new_n1129 ^ new_n771;
  assign new_n1131 = n458 ^ n202;
  assign new_n1132 = new_n1131 ^ new_n950;
  assign new_n1133 = n395 ^ n139;
  assign new_n1134 = new_n1133 ^ n10;
  assign new_n1135 = ~new_n1134 & new_n1132;
  assign new_n1136 = new_n1135 ^ new_n1130;
  assign new_n1137 = n543 ^ n287;
  assign new_n1138 = new_n1137 ^ new_n781;
  assign new_n1139 = n459 ^ n203;
  assign new_n1140 = new_n1139 ^ new_n959;
  assign new_n1141 = n396 ^ n140;
  assign new_n1142 = new_n1141 ^ n11;
  assign new_n1143 = ~new_n1142 & new_n1140;
  assign new_n1144 = new_n1143 ^ new_n1138;
  assign new_n1145 = n544 ^ n288;
  assign new_n1146 = new_n1145 ^ new_n791;
  assign new_n1147 = n460 ^ n204;
  assign new_n1148 = new_n1147 ^ new_n968;
  assign new_n1149 = n397 ^ n141;
  assign new_n1150 = new_n1149 ^ n12;
  assign new_n1151 = ~new_n1150 & new_n1148;
  assign new_n1152 = new_n1151 ^ new_n1146;
  assign new_n1153 = new_n964 ^ new_n798;
  assign new_n1154 = new_n1153 ^ n438;
  assign new_n1155 = ~new_n582 & new_n1154;
  assign new_n1156 = new_n1155 ^ new_n584;
  assign new_n1157 = new_n973 ^ new_n807;
  assign new_n1158 = new_n1157 ^ n439;
  assign new_n1159 = ~new_n592 & new_n1158;
  assign new_n1160 = new_n1159 ^ new_n594;
  assign new_n1161 = new_n981 ^ new_n816;
  assign new_n1162 = new_n1161 ^ n440;
  assign new_n1163 = ~new_n602 & new_n1162;
  assign new_n1164 = new_n1163 ^ new_n604;
  assign new_n1165 = new_n989 ^ new_n825;
  assign new_n1166 = new_n1165 ^ n441;
  assign new_n1167 = ~new_n612 & new_n1166;
  assign new_n1168 = new_n1167 ^ new_n614;
  assign new_n1169 = new_n997 ^ new_n834;
  assign new_n1170 = new_n1169 ^ n442;
  assign new_n1171 = ~new_n622 & new_n1170;
  assign new_n1172 = new_n1171 ^ new_n624;
  assign new_n1173 = new_n1005 ^ new_n843;
  assign new_n1174 = new_n1173 ^ n443;
  assign new_n1175 = ~new_n632 & new_n1174;
  assign new_n1176 = new_n1175 ^ new_n634;
  assign new_n1177 = new_n1013 ^ new_n852;
  assign new_n1178 = new_n1177 ^ n444;
  assign new_n1179 = ~new_n642 & new_n1178;
  assign new_n1180 = new_n1179 ^ new_n644;
  assign new_n1181 = new_n1021 ^ new_n861;
  assign new_n1182 = new_n1181 ^ n445;
  assign new_n1183 = ~new_n652 & new_n1182;
  assign new_n1184 = new_n1183 ^ new_n654;
  assign new_n1185 = new_n1029 ^ new_n870;
  assign new_n1186 = new_n1185 ^ n446;
  assign new_n1187 = ~new_n662 & new_n1186;
  assign new_n1188 = new_n1187 ^ new_n664;
  assign new_n1189 = new_n1037 ^ new_n879;
  assign new_n1190 = new_n1189 ^ n447;
  assign new_n1191 = ~new_n672 & new_n1190;
  assign new_n1192 = new_n1191 ^ new_n674;
  assign new_n1193 = new_n1045 ^ new_n888;
  assign new_n1194 = new_n1193 ^ n448;
  assign new_n1195 = ~new_n682 & new_n1194;
  assign new_n1196 = new_n1195 ^ new_n684;
  assign new_n1197 = new_n1053 ^ new_n897;
  assign new_n1198 = new_n1197 ^ n449;
  assign new_n1199 = ~new_n692 & new_n1198;
  assign new_n1200 = new_n1199 ^ new_n694;
  assign new_n1201 = new_n1061 ^ new_n906;
  assign new_n1202 = new_n1201 ^ n450;
  assign new_n1203 = ~new_n702 & new_n1202;
  assign new_n1204 = new_n1203 ^ new_n704;
  assign new_n1205 = new_n1069 ^ new_n915;
  assign new_n1206 = new_n1205 ^ n451;
  assign new_n1207 = ~new_n712 & new_n1206;
  assign new_n1208 = new_n1207 ^ new_n714;
  assign new_n1209 = new_n1077 ^ new_n924;
  assign new_n1210 = new_n1209 ^ n452;
  assign new_n1211 = ~new_n722 & new_n1210;
  assign new_n1212 = new_n1211 ^ new_n724;
  assign new_n1213 = new_n1085 ^ new_n933;
  assign new_n1214 = new_n1213 ^ n453;
  assign new_n1215 = ~new_n732 & new_n1214;
  assign new_n1216 = new_n1215 ^ new_n734;
  assign new_n1217 = new_n1093 ^ new_n942;
  assign new_n1218 = new_n1217 ^ n454;
  assign new_n1219 = ~new_n742 & new_n1218;
  assign new_n1220 = new_n1219 ^ new_n744;
  assign new_n1221 = new_n1101 ^ new_n951;
  assign new_n1222 = new_n1221 ^ n455;
  assign new_n1223 = ~new_n752 & new_n1222;
  assign new_n1224 = new_n1223 ^ new_n754;
  assign new_n1225 = new_n1109 ^ new_n960;
  assign new_n1226 = new_n1225 ^ n456;
  assign new_n1227 = ~new_n762 & new_n1226;
  assign new_n1228 = new_n1227 ^ new_n764;
  assign new_n1229 = new_n1117 ^ new_n969;
  assign new_n1230 = new_n1229 ^ n457;
  assign new_n1231 = ~new_n772 & new_n1230;
  assign new_n1232 = new_n1231 ^ new_n774;
  assign new_n1233 = new_n1125 ^ new_n977;
  assign new_n1234 = new_n1233 ^ n458;
  assign new_n1235 = ~new_n782 & new_n1234;
  assign new_n1236 = new_n1235 ^ new_n784;
  assign new_n1237 = new_n1133 ^ new_n985;
  assign new_n1238 = new_n1237 ^ n459;
  assign new_n1239 = ~new_n792 & new_n1238;
  assign new_n1240 = new_n1239 ^ new_n794;
  assign new_n1241 = new_n1141 ^ new_n993;
  assign new_n1242 = new_n1241 ^ n460;
  assign new_n1243 = ~new_n801 & new_n1242;
  assign new_n1244 = new_n1243 ^ new_n803;
  assign new_n1245 = new_n1149 ^ new_n1001;
  assign new_n1246 = new_n1245 ^ n461;
  assign new_n1247 = ~new_n810 & new_n1246;
  assign new_n1248 = new_n1247 ^ new_n812;
  assign new_n1249 = new_n1009 ^ new_n583;
  assign new_n1250 = new_n1249 ^ n462;
  assign new_n1251 = ~new_n819 & new_n1250;
  assign new_n1252 = new_n1251 ^ new_n821;
  assign new_n1253 = new_n1017 ^ new_n593;
  assign new_n1254 = new_n1253 ^ n463;
  assign new_n1255 = ~new_n828 & new_n1254;
  assign new_n1256 = new_n1255 ^ new_n830;
  assign new_n1257 = new_n1025 ^ new_n603;
  assign new_n1258 = new_n1257 ^ n464;
  assign new_n1259 = ~new_n837 & new_n1258;
  assign new_n1260 = new_n1259 ^ new_n839;
  assign new_n1261 = new_n1033 ^ new_n613;
  assign new_n1262 = new_n1261 ^ n465;
  assign new_n1263 = ~new_n846 & new_n1262;
  assign new_n1264 = new_n1263 ^ new_n848;
  assign new_n1265 = new_n1041 ^ new_n623;
  assign new_n1266 = new_n1265 ^ n466;
  assign new_n1267 = ~new_n855 & new_n1266;
  assign new_n1268 = new_n1267 ^ new_n857;
  assign new_n1269 = new_n1049 ^ new_n633;
  assign new_n1270 = new_n1269 ^ n467;
  assign new_n1271 = ~new_n864 & new_n1270;
  assign new_n1272 = new_n1271 ^ new_n866;
  assign new_n1273 = new_n1057 ^ new_n643;
  assign new_n1274 = new_n1273 ^ n468;
  assign new_n1275 = ~new_n873 & new_n1274;
  assign new_n1276 = new_n1275 ^ new_n875;
  assign new_n1277 = new_n1065 ^ new_n653;
  assign new_n1278 = new_n1277 ^ n469;
  assign new_n1279 = ~new_n882 & new_n1278;
  assign new_n1280 = new_n1279 ^ new_n884;
  assign new_n1281 = new_n1073 ^ new_n663;
  assign new_n1282 = new_n1281 ^ n470;
  assign new_n1283 = ~new_n891 & new_n1282;
  assign new_n1284 = new_n1283 ^ new_n893;
  assign new_n1285 = new_n1081 ^ new_n673;
  assign new_n1286 = new_n1285 ^ n471;
  assign new_n1287 = ~new_n900 & new_n1286;
  assign new_n1288 = new_n1287 ^ new_n902;
  assign new_n1289 = new_n1089 ^ new_n683;
  assign new_n1290 = new_n1289 ^ n472;
  assign new_n1291 = ~new_n909 & new_n1290;
  assign new_n1292 = new_n1291 ^ new_n911;
  assign new_n1293 = new_n1097 ^ new_n693;
  assign new_n1294 = new_n1293 ^ n473;
  assign new_n1295 = ~new_n918 & new_n1294;
  assign new_n1296 = new_n1295 ^ new_n920;
  assign new_n1297 = new_n1105 ^ new_n703;
  assign new_n1298 = new_n1297 ^ n474;
  assign new_n1299 = ~new_n927 & new_n1298;
  assign new_n1300 = new_n1299 ^ new_n929;
  assign new_n1301 = new_n1113 ^ new_n713;
  assign new_n1302 = new_n1301 ^ n475;
  assign new_n1303 = ~new_n936 & new_n1302;
  assign new_n1304 = new_n1303 ^ new_n938;
  assign new_n1305 = new_n1121 ^ new_n723;
  assign new_n1306 = new_n1305 ^ n476;
  assign new_n1307 = ~new_n945 & new_n1306;
  assign new_n1308 = new_n1307 ^ new_n947;
  assign new_n1309 = new_n1129 ^ new_n733;
  assign new_n1310 = new_n1309 ^ n477;
  assign new_n1311 = ~new_n954 & new_n1310;
  assign new_n1312 = new_n1311 ^ new_n956;
  assign new_n1313 = new_n1137 ^ new_n743;
  assign new_n1314 = new_n1313 ^ n478;
  assign new_n1315 = ~new_n963 & new_n1314;
  assign new_n1316 = new_n1315 ^ new_n965;
  assign new_n1317 = new_n1145 ^ new_n753;
  assign new_n1318 = new_n1317 ^ n479;
  assign new_n1319 = ~new_n972 & new_n1318;
  assign new_n1320 = new_n1319 ^ new_n974;
  assign new_n1321 = new_n763 ^ new_n577;
  assign new_n1322 = new_n1321 ^ n480;
  assign new_n1323 = ~new_n980 & new_n1322;
  assign new_n1324 = new_n1323 ^ new_n982;
  assign new_n1325 = new_n773 ^ new_n587;
  assign new_n1326 = new_n1325 ^ n417;
  assign new_n1327 = ~new_n988 & new_n1326;
  assign new_n1328 = new_n1327 ^ new_n990;
  assign new_n1329 = new_n783 ^ new_n597;
  assign new_n1330 = new_n1329 ^ n418;
  assign new_n1331 = ~new_n996 & new_n1330;
  assign new_n1332 = new_n1331 ^ new_n998;
  assign new_n1333 = new_n793 ^ new_n607;
  assign new_n1334 = new_n1333 ^ n419;
  assign new_n1335 = ~new_n1004 & new_n1334;
  assign new_n1336 = new_n1335 ^ new_n1006;
  assign new_n1337 = new_n802 ^ new_n617;
  assign new_n1338 = new_n1337 ^ n420;
  assign new_n1339 = ~new_n1012 & new_n1338;
  assign new_n1340 = new_n1339 ^ new_n1014;
  assign new_n1341 = new_n811 ^ new_n627;
  assign new_n1342 = new_n1341 ^ n421;
  assign new_n1343 = ~new_n1020 & new_n1342;
  assign new_n1344 = new_n1343 ^ new_n1022;
  assign new_n1345 = new_n820 ^ new_n637;
  assign new_n1346 = new_n1345 ^ n422;
  assign new_n1347 = ~new_n1028 & new_n1346;
  assign new_n1348 = new_n1347 ^ new_n1030;
  assign new_n1349 = new_n829 ^ new_n647;
  assign new_n1350 = new_n1349 ^ n423;
  assign new_n1351 = ~new_n1036 & new_n1350;
  assign new_n1352 = new_n1351 ^ new_n1038;
  assign new_n1353 = new_n838 ^ new_n657;
  assign new_n1354 = new_n1353 ^ n424;
  assign new_n1355 = ~new_n1044 & new_n1354;
  assign new_n1356 = new_n1355 ^ new_n1046;
  assign new_n1357 = new_n847 ^ new_n667;
  assign new_n1358 = new_n1357 ^ n425;
  assign new_n1359 = ~new_n1052 & new_n1358;
  assign new_n1360 = new_n1359 ^ new_n1054;
  assign new_n1361 = new_n856 ^ new_n677;
  assign new_n1362 = new_n1361 ^ n426;
  assign new_n1363 = ~new_n1060 & new_n1362;
  assign new_n1364 = new_n1363 ^ new_n1062;
  assign new_n1365 = new_n865 ^ new_n687;
  assign new_n1366 = new_n1365 ^ n427;
  assign new_n1367 = ~new_n1068 & new_n1366;
  assign new_n1368 = new_n1367 ^ new_n1070;
  assign new_n1369 = new_n874 ^ new_n697;
  assign new_n1370 = new_n1369 ^ n428;
  assign new_n1371 = ~new_n1076 & new_n1370;
  assign new_n1372 = new_n1371 ^ new_n1078;
  assign new_n1373 = new_n883 ^ new_n707;
  assign new_n1374 = new_n1373 ^ n429;
  assign new_n1375 = ~new_n1084 & new_n1374;
  assign new_n1376 = new_n1375 ^ new_n1086;
  assign new_n1377 = new_n892 ^ new_n717;
  assign new_n1378 = new_n1377 ^ n430;
  assign new_n1379 = ~new_n1092 & new_n1378;
  assign new_n1380 = new_n1379 ^ new_n1094;
  assign new_n1381 = new_n901 ^ new_n727;
  assign new_n1382 = new_n1381 ^ n431;
  assign new_n1383 = ~new_n1100 & new_n1382;
  assign new_n1384 = new_n1383 ^ new_n1102;
  assign new_n1385 = new_n910 ^ new_n737;
  assign new_n1386 = new_n1385 ^ n432;
  assign new_n1387 = ~new_n1108 & new_n1386;
  assign new_n1388 = new_n1387 ^ new_n1110;
  assign new_n1389 = new_n919 ^ new_n747;
  assign new_n1390 = new_n1389 ^ n433;
  assign new_n1391 = ~new_n1116 & new_n1390;
  assign new_n1392 = new_n1391 ^ new_n1118;
  assign new_n1393 = new_n928 ^ new_n757;
  assign new_n1394 = new_n1393 ^ n434;
  assign new_n1395 = ~new_n1124 & new_n1394;
  assign new_n1396 = new_n1395 ^ new_n1126;
  assign new_n1397 = new_n937 ^ new_n767;
  assign new_n1398 = new_n1397 ^ n435;
  assign new_n1399 = ~new_n1132 & new_n1398;
  assign new_n1400 = new_n1399 ^ new_n1134;
  assign new_n1401 = new_n946 ^ new_n778;
  assign new_n1402 = new_n1401 ^ n436;
  assign new_n1403 = ~new_n1140 & new_n1402;
  assign new_n1404 = new_n1403 ^ new_n1142;
  assign new_n1405 = new_n955 ^ new_n788;
  assign new_n1406 = new_n1405 ^ n437;
  assign new_n1407 = ~new_n1148 & new_n1406;
  assign new_n1408 = new_n1407 ^ new_n1150;
  assign new_n1409 = new_n908 ^ n560;
  assign new_n1410 = new_n1409 ^ n239;
  assign new_n1411 = ~new_n1154 & new_n1410;
  assign new_n1412 = new_n1411 ^ new_n582;
  assign new_n1413 = new_n917 ^ n561;
  assign new_n1414 = new_n1413 ^ n240;
  assign new_n1415 = ~new_n1158 & new_n1414;
  assign new_n1416 = new_n1415 ^ new_n592;
  assign new_n1417 = new_n926 ^ n562;
  assign new_n1418 = new_n1417 ^ n241;
  assign new_n1419 = ~new_n1162 & new_n1418;
  assign new_n1420 = new_n1419 ^ new_n602;
  assign new_n1421 = new_n935 ^ n563;
  assign new_n1422 = new_n1421 ^ n242;
  assign new_n1423 = ~new_n1166 & new_n1422;
  assign new_n1424 = new_n1423 ^ new_n612;
  assign new_n1425 = new_n944 ^ n564;
  assign new_n1426 = new_n1425 ^ n243;
  assign new_n1427 = ~new_n1170 & new_n1426;
  assign new_n1428 = new_n1427 ^ new_n622;
  assign new_n1429 = new_n953 ^ n565;
  assign new_n1430 = new_n1429 ^ n244;
  assign new_n1431 = ~new_n1174 & new_n1430;
  assign new_n1432 = new_n1431 ^ new_n632;
  assign new_n1433 = new_n962 ^ n566;
  assign new_n1434 = new_n1433 ^ n245;
  assign new_n1435 = ~new_n1178 & new_n1434;
  assign new_n1436 = new_n1435 ^ new_n642;
  assign new_n1437 = new_n971 ^ n567;
  assign new_n1438 = new_n1437 ^ n246;
  assign new_n1439 = ~new_n1182 & new_n1438;
  assign new_n1440 = new_n1439 ^ new_n652;
  assign new_n1441 = new_n979 ^ n568;
  assign new_n1442 = new_n1441 ^ n247;
  assign new_n1443 = ~new_n1186 & new_n1442;
  assign new_n1444 = new_n1443 ^ new_n662;
  assign new_n1445 = new_n987 ^ n569;
  assign new_n1446 = new_n1445 ^ n248;
  assign new_n1447 = ~new_n1190 & new_n1446;
  assign new_n1448 = new_n1447 ^ new_n672;
  assign new_n1449 = new_n995 ^ n570;
  assign new_n1450 = new_n1449 ^ n249;
  assign new_n1451 = ~new_n1194 & new_n1450;
  assign new_n1452 = new_n1451 ^ new_n682;
  assign new_n1453 = new_n1003 ^ n571;
  assign new_n1454 = new_n1453 ^ n250;
  assign new_n1455 = ~new_n1198 & new_n1454;
  assign new_n1456 = new_n1455 ^ new_n692;
  assign new_n1457 = new_n1011 ^ n572;
  assign new_n1458 = new_n1457 ^ n251;
  assign new_n1459 = ~new_n1202 & new_n1458;
  assign new_n1460 = new_n1459 ^ new_n702;
  assign new_n1461 = new_n1019 ^ n573;
  assign new_n1462 = new_n1461 ^ n252;
  assign new_n1463 = ~new_n1206 & new_n1462;
  assign new_n1464 = new_n1463 ^ new_n712;
  assign new_n1465 = new_n1027 ^ n574;
  assign new_n1466 = new_n1465 ^ n253;
  assign new_n1467 = ~new_n1210 & new_n1466;
  assign new_n1468 = new_n1467 ^ new_n722;
  assign new_n1469 = new_n1035 ^ n575;
  assign new_n1470 = new_n1469 ^ n254;
  assign new_n1471 = ~new_n1214 & new_n1470;
  assign new_n1472 = new_n1471 ^ new_n732;
  assign new_n1473 = new_n1043 ^ n576;
  assign new_n1474 = new_n1473 ^ n255;
  assign new_n1475 = ~new_n1218 & new_n1474;
  assign new_n1476 = new_n1475 ^ new_n742;
  assign new_n1477 = new_n1051 ^ n1;
  assign new_n1478 = new_n1477 ^ n256;
  assign new_n1479 = ~new_n1222 & new_n1478;
  assign new_n1480 = new_n1479 ^ new_n752;
  assign new_n1481 = new_n1059 ^ n2;
  assign new_n1482 = new_n1481 ^ n257;
  assign new_n1483 = ~new_n1226 & new_n1482;
  assign new_n1484 = new_n1483 ^ new_n762;
  assign new_n1485 = new_n1067 ^ n3;
  assign new_n1486 = new_n1485 ^ n258;
  assign new_n1487 = ~new_n1230 & new_n1486;
  assign new_n1488 = new_n1487 ^ new_n772;
  assign new_n1489 = new_n1075 ^ n4;
  assign new_n1490 = new_n1489 ^ n259;
  assign new_n1491 = ~new_n1234 & new_n1490;
  assign new_n1492 = new_n1491 ^ new_n782;
  assign new_n1493 = new_n1083 ^ n5;
  assign new_n1494 = new_n1493 ^ n260;
  assign new_n1495 = ~new_n1238 & new_n1494;
  assign new_n1496 = new_n1495 ^ new_n792;
  assign new_n1497 = new_n1091 ^ n6;
  assign new_n1498 = new_n1497 ^ n261;
  assign new_n1499 = ~new_n1242 & new_n1498;
  assign new_n1500 = new_n1499 ^ new_n801;
  assign new_n1501 = new_n1099 ^ n7;
  assign new_n1502 = new_n1501 ^ n262;
  assign new_n1503 = ~new_n1246 & new_n1502;
  assign new_n1504 = new_n1503 ^ new_n810;
  assign new_n1505 = new_n1107 ^ n8;
  assign new_n1506 = new_n1505 ^ n263;
  assign new_n1507 = ~new_n1250 & new_n1506;
  assign new_n1508 = new_n1507 ^ new_n819;
  assign new_n1509 = new_n1115 ^ n9;
  assign new_n1510 = new_n1509 ^ n264;
  assign new_n1511 = ~new_n1254 & new_n1510;
  assign new_n1512 = new_n1511 ^ new_n828;
  assign new_n1513 = new_n1123 ^ n10;
  assign new_n1514 = new_n1513 ^ n265;
  assign new_n1515 = ~new_n1258 & new_n1514;
  assign new_n1516 = new_n1515 ^ new_n837;
  assign new_n1517 = new_n1131 ^ n11;
  assign new_n1518 = new_n1517 ^ n266;
  assign new_n1519 = ~new_n1262 & new_n1518;
  assign new_n1520 = new_n1519 ^ new_n846;
  assign new_n1521 = new_n1139 ^ n12;
  assign new_n1522 = new_n1521 ^ n267;
  assign new_n1523 = ~new_n1266 & new_n1522;
  assign new_n1524 = new_n1523 ^ new_n855;
  assign new_n1525 = new_n1147 ^ n13;
  assign new_n1526 = new_n1525 ^ n268;
  assign new_n1527 = ~new_n1270 & new_n1526;
  assign new_n1528 = new_n1527 ^ new_n864;
  assign new_n1529 = new_n580 ^ n14;
  assign new_n1530 = new_n1529 ^ n269;
  assign new_n1531 = ~new_n1274 & new_n1530;
  assign new_n1532 = new_n1531 ^ new_n873;
  assign new_n1533 = new_n590 ^ n15;
  assign new_n1534 = new_n1533 ^ n270;
  assign new_n1535 = ~new_n1278 & new_n1534;
  assign new_n1536 = new_n1535 ^ new_n882;
  assign new_n1537 = new_n600 ^ n16;
  assign new_n1538 = new_n1537 ^ n271;
  assign new_n1539 = ~new_n1282 & new_n1538;
  assign new_n1540 = new_n1539 ^ new_n891;
  assign new_n1541 = new_n610 ^ n17;
  assign new_n1542 = new_n1541 ^ n272;
  assign new_n1543 = ~new_n1286 & new_n1542;
  assign new_n1544 = new_n1543 ^ new_n900;
  assign new_n1545 = new_n620 ^ n18;
  assign new_n1546 = new_n1545 ^ n273;
  assign new_n1547 = ~new_n1290 & new_n1546;
  assign new_n1548 = new_n1547 ^ new_n909;
  assign new_n1549 = new_n630 ^ n19;
  assign new_n1550 = new_n1549 ^ n274;
  assign new_n1551 = ~new_n1294 & new_n1550;
  assign new_n1552 = new_n1551 ^ new_n918;
  assign new_n1553 = new_n640 ^ n20;
  assign new_n1554 = new_n1553 ^ n275;
  assign new_n1555 = ~new_n1298 & new_n1554;
  assign new_n1556 = new_n1555 ^ new_n927;
  assign new_n1557 = new_n650 ^ n21;
  assign new_n1558 = new_n1557 ^ n276;
  assign new_n1559 = ~new_n1302 & new_n1558;
  assign new_n1560 = new_n1559 ^ new_n936;
  assign new_n1561 = new_n660 ^ n22;
  assign new_n1562 = new_n1561 ^ n277;
  assign new_n1563 = ~new_n1306 & new_n1562;
  assign new_n1564 = new_n1563 ^ new_n945;
  assign new_n1565 = new_n670 ^ n23;
  assign new_n1566 = new_n1565 ^ n278;
  assign new_n1567 = ~new_n1310 & new_n1566;
  assign new_n1568 = new_n1567 ^ new_n954;
  assign new_n1569 = new_n680 ^ n24;
  assign new_n1570 = new_n1569 ^ n279;
  assign new_n1571 = ~new_n1314 & new_n1570;
  assign new_n1572 = new_n1571 ^ new_n963;
  assign new_n1573 = new_n690 ^ n25;
  assign new_n1574 = new_n1573 ^ n280;
  assign new_n1575 = ~new_n1318 & new_n1574;
  assign new_n1576 = new_n1575 ^ new_n972;
  assign new_n1577 = new_n700 ^ n26;
  assign new_n1578 = new_n1577 ^ n281;
  assign new_n1579 = ~new_n1322 & new_n1578;
  assign new_n1580 = new_n1579 ^ new_n980;
  assign new_n1581 = new_n710 ^ n27;
  assign new_n1582 = new_n1581 ^ n282;
  assign new_n1583 = ~new_n1326 & new_n1582;
  assign new_n1584 = new_n1583 ^ new_n988;
  assign new_n1585 = new_n720 ^ n28;
  assign new_n1586 = new_n1585 ^ n283;
  assign new_n1587 = ~new_n1330 & new_n1586;
  assign new_n1588 = new_n1587 ^ new_n996;
  assign new_n1589 = new_n730 ^ n29;
  assign new_n1590 = new_n1589 ^ n284;
  assign new_n1591 = ~new_n1334 & new_n1590;
  assign new_n1592 = new_n1591 ^ new_n1004;
  assign new_n1593 = new_n740 ^ n30;
  assign new_n1594 = new_n1593 ^ n285;
  assign new_n1595 = ~new_n1338 & new_n1594;
  assign new_n1596 = new_n1595 ^ new_n1012;
  assign new_n1597 = new_n750 ^ n31;
  assign new_n1598 = new_n1597 ^ n286;
  assign new_n1599 = ~new_n1342 & new_n1598;
  assign new_n1600 = new_n1599 ^ new_n1020;
  assign new_n1601 = new_n760 ^ n32;
  assign new_n1602 = new_n1601 ^ n287;
  assign new_n1603 = ~new_n1346 & new_n1602;
  assign new_n1604 = new_n1603 ^ new_n1028;
  assign new_n1605 = new_n770 ^ n545;
  assign new_n1606 = new_n1605 ^ n288;
  assign new_n1607 = ~new_n1350 & new_n1606;
  assign new_n1608 = new_n1607 ^ new_n1036;
  assign new_n1609 = new_n780 ^ n546;
  assign new_n1610 = new_n1609 ^ n225;
  assign new_n1611 = ~new_n1354 & new_n1610;
  assign new_n1612 = new_n1611 ^ new_n1044;
  assign new_n1613 = new_n790 ^ n547;
  assign new_n1614 = new_n1613 ^ n226;
  assign new_n1615 = ~new_n1358 & new_n1614;
  assign new_n1616 = new_n1615 ^ new_n1052;
  assign new_n1617 = new_n800 ^ n548;
  assign new_n1618 = new_n1617 ^ n227;
  assign new_n1619 = ~new_n1362 & new_n1618;
  assign new_n1620 = new_n1619 ^ new_n1060;
  assign new_n1621 = new_n809 ^ n549;
  assign new_n1622 = new_n1621 ^ n228;
  assign new_n1623 = ~new_n1366 & new_n1622;
  assign new_n1624 = new_n1623 ^ new_n1068;
  assign new_n1625 = new_n818 ^ n550;
  assign new_n1626 = new_n1625 ^ n229;
  assign new_n1627 = ~new_n1370 & new_n1626;
  assign new_n1628 = new_n1627 ^ new_n1076;
  assign new_n1629 = new_n827 ^ n551;
  assign new_n1630 = new_n1629 ^ n230;
  assign new_n1631 = ~new_n1374 & new_n1630;
  assign new_n1632 = new_n1631 ^ new_n1084;
  assign new_n1633 = new_n836 ^ n552;
  assign new_n1634 = new_n1633 ^ n231;
  assign new_n1635 = ~new_n1378 & new_n1634;
  assign new_n1636 = new_n1635 ^ new_n1092;
  assign new_n1637 = new_n845 ^ n553;
  assign new_n1638 = new_n1637 ^ n232;
  assign new_n1639 = ~new_n1382 & new_n1638;
  assign new_n1640 = new_n1639 ^ new_n1100;
  assign new_n1641 = new_n854 ^ n554;
  assign new_n1642 = new_n1641 ^ n233;
  assign new_n1643 = ~new_n1386 & new_n1642;
  assign new_n1644 = new_n1643 ^ new_n1108;
  assign new_n1645 = new_n863 ^ n555;
  assign new_n1646 = new_n1645 ^ n234;
  assign new_n1647 = ~new_n1390 & new_n1646;
  assign new_n1648 = new_n1647 ^ new_n1116;
  assign new_n1649 = new_n872 ^ n556;
  assign new_n1650 = new_n1649 ^ n235;
  assign new_n1651 = ~new_n1394 & new_n1650;
  assign new_n1652 = new_n1651 ^ new_n1124;
  assign new_n1653 = new_n881 ^ n557;
  assign new_n1654 = new_n1653 ^ n236;
  assign new_n1655 = ~new_n1398 & new_n1654;
  assign new_n1656 = new_n1655 ^ new_n1132;
  assign new_n1657 = new_n890 ^ n558;
  assign new_n1658 = new_n1657 ^ n237;
  assign new_n1659 = ~new_n1402 & new_n1658;
  assign new_n1660 = new_n1659 ^ new_n1140;
  assign new_n1661 = new_n899 ^ n559;
  assign new_n1662 = new_n1661 ^ n238;
  assign new_n1663 = ~new_n1406 & new_n1662;
  assign new_n1664 = new_n1663 ^ new_n1148;
  assign new_n1665 = ~new_n1410 & new_n579;
  assign new_n1666 = new_n1665 ^ new_n1154;
  assign new_n1667 = ~new_n1414 & new_n589;
  assign new_n1668 = new_n1667 ^ new_n1158;
  assign new_n1669 = ~new_n1418 & new_n599;
  assign new_n1670 = new_n1669 ^ new_n1162;
  assign new_n1671 = ~new_n1422 & new_n609;
  assign new_n1672 = new_n1671 ^ new_n1166;
  assign new_n1673 = ~new_n1426 & new_n619;
  assign new_n1674 = new_n1673 ^ new_n1170;
  assign new_n1675 = ~new_n1430 & new_n629;
  assign new_n1676 = new_n1675 ^ new_n1174;
  assign new_n1677 = ~new_n1434 & new_n639;
  assign new_n1678 = new_n1677 ^ new_n1178;
  assign new_n1679 = ~new_n1438 & new_n649;
  assign new_n1680 = new_n1679 ^ new_n1182;
  assign new_n1681 = ~new_n1442 & new_n659;
  assign new_n1682 = new_n1681 ^ new_n1186;
  assign new_n1683 = ~new_n1446 & new_n669;
  assign new_n1684 = new_n1683 ^ new_n1190;
  assign new_n1685 = ~new_n1450 & new_n679;
  assign new_n1686 = new_n1685 ^ new_n1194;
  assign new_n1687 = ~new_n1454 & new_n689;
  assign new_n1688 = new_n1687 ^ new_n1198;
  assign new_n1689 = ~new_n1458 & new_n699;
  assign new_n1690 = new_n1689 ^ new_n1202;
  assign new_n1691 = ~new_n1462 & new_n709;
  assign new_n1692 = new_n1691 ^ new_n1206;
  assign new_n1693 = ~new_n1466 & new_n719;
  assign new_n1694 = new_n1693 ^ new_n1210;
  assign new_n1695 = ~new_n1470 & new_n729;
  assign new_n1696 = new_n1695 ^ new_n1214;
  assign new_n1697 = ~new_n1474 & new_n739;
  assign new_n1698 = new_n1697 ^ new_n1218;
  assign new_n1699 = ~new_n1478 & new_n749;
  assign new_n1700 = new_n1699 ^ new_n1222;
  assign new_n1701 = ~new_n1482 & new_n759;
  assign new_n1702 = new_n1701 ^ new_n1226;
  assign new_n1703 = ~new_n1486 & new_n769;
  assign new_n1704 = new_n1703 ^ new_n1230;
  assign new_n1705 = ~new_n1490 & new_n779;
  assign new_n1706 = new_n1705 ^ new_n1234;
  assign new_n1707 = ~new_n1494 & new_n789;
  assign new_n1708 = new_n1707 ^ new_n1238;
  assign new_n1709 = ~new_n1498 & new_n799;
  assign new_n1710 = new_n1709 ^ new_n1242;
  assign new_n1711 = ~new_n1502 & new_n808;
  assign new_n1712 = new_n1711 ^ new_n1246;
  assign new_n1713 = ~new_n1506 & new_n817;
  assign new_n1714 = new_n1713 ^ new_n1250;
  assign new_n1715 = ~new_n1510 & new_n826;
  assign new_n1716 = new_n1715 ^ new_n1254;
  assign new_n1717 = ~new_n1514 & new_n835;
  assign new_n1718 = new_n1717 ^ new_n1258;
  assign new_n1719 = ~new_n1518 & new_n844;
  assign new_n1720 = new_n1719 ^ new_n1262;
  assign new_n1721 = ~new_n1522 & new_n853;
  assign new_n1722 = new_n1721 ^ new_n1266;
  assign new_n1723 = ~new_n1526 & new_n862;
  assign new_n1724 = new_n1723 ^ new_n1270;
  assign new_n1725 = ~new_n1530 & new_n871;
  assign new_n1726 = new_n1725 ^ new_n1274;
  assign new_n1727 = ~new_n1534 & new_n880;
  assign new_n1728 = new_n1727 ^ new_n1278;
  assign new_n1729 = ~new_n1538 & new_n889;
  assign new_n1730 = new_n1729 ^ new_n1282;
  assign new_n1731 = ~new_n1542 & new_n898;
  assign new_n1732 = new_n1731 ^ new_n1286;
  assign new_n1733 = ~new_n1546 & new_n907;
  assign new_n1734 = new_n1733 ^ new_n1290;
  assign new_n1735 = ~new_n1550 & new_n916;
  assign new_n1736 = new_n1735 ^ new_n1294;
  assign new_n1737 = ~new_n1554 & new_n925;
  assign new_n1738 = new_n1737 ^ new_n1298;
  assign new_n1739 = ~new_n1558 & new_n934;
  assign new_n1740 = new_n1739 ^ new_n1302;
  assign new_n1741 = ~new_n1562 & new_n943;
  assign new_n1742 = new_n1741 ^ new_n1306;
  assign new_n1743 = ~new_n1566 & new_n952;
  assign new_n1744 = new_n1743 ^ new_n1310;
  assign new_n1745 = ~new_n1570 & new_n961;
  assign new_n1746 = new_n1745 ^ new_n1314;
  assign new_n1747 = ~new_n1574 & new_n970;
  assign new_n1748 = new_n1747 ^ new_n1318;
  assign new_n1749 = ~new_n1578 & new_n978;
  assign new_n1750 = new_n1749 ^ new_n1322;
  assign new_n1751 = ~new_n1582 & new_n986;
  assign new_n1752 = new_n1751 ^ new_n1326;
  assign new_n1753 = ~new_n1586 & new_n994;
  assign new_n1754 = new_n1753 ^ new_n1330;
  assign new_n1755 = ~new_n1590 & new_n1002;
  assign new_n1756 = new_n1755 ^ new_n1334;
  assign new_n1757 = ~new_n1594 & new_n1010;
  assign new_n1758 = new_n1757 ^ new_n1338;
  assign new_n1759 = ~new_n1598 & new_n1018;
  assign new_n1760 = new_n1759 ^ new_n1342;
  assign new_n1761 = ~new_n1602 & new_n1026;
  assign new_n1762 = new_n1761 ^ new_n1346;
  assign new_n1763 = ~new_n1606 & new_n1034;
  assign new_n1764 = new_n1763 ^ new_n1350;
  assign new_n1765 = ~new_n1610 & new_n1042;
  assign new_n1766 = new_n1765 ^ new_n1354;
  assign new_n1767 = ~new_n1614 & new_n1050;
  assign new_n1768 = new_n1767 ^ new_n1358;
  assign new_n1769 = ~new_n1618 & new_n1058;
  assign new_n1770 = new_n1769 ^ new_n1362;
  assign new_n1771 = ~new_n1622 & new_n1066;
  assign new_n1772 = new_n1771 ^ new_n1366;
  assign new_n1773 = ~new_n1626 & new_n1074;
  assign new_n1774 = new_n1773 ^ new_n1370;
  assign new_n1775 = ~new_n1630 & new_n1082;
  assign new_n1776 = new_n1775 ^ new_n1374;
  assign new_n1777 = ~new_n1634 & new_n1090;
  assign new_n1778 = new_n1777 ^ new_n1378;
  assign new_n1779 = ~new_n1638 & new_n1098;
  assign new_n1780 = new_n1779 ^ new_n1382;
  assign new_n1781 = ~new_n1642 & new_n1106;
  assign new_n1782 = new_n1781 ^ new_n1386;
  assign new_n1783 = ~new_n1646 & new_n1114;
  assign new_n1784 = new_n1783 ^ new_n1390;
  assign new_n1785 = ~new_n1650 & new_n1122;
  assign new_n1786 = new_n1785 ^ new_n1394;
  assign new_n1787 = ~new_n1654 & new_n1130;
  assign new_n1788 = new_n1787 ^ new_n1398;
  assign new_n1789 = ~new_n1658 & new_n1138;
  assign new_n1790 = new_n1789 ^ new_n1402;
  assign new_n1791 = ~new_n1662 & new_n1146;
  assign new_n1792 = new_n1791 ^ new_n1406;
  assign new_n1793 = ~new_n579 & new_n584;
  assign new_n1794 = new_n1793 ^ new_n1410;
  assign new_n1795 = ~new_n589 & new_n594;
  assign new_n1796 = new_n1795 ^ new_n1414;
  assign new_n1797 = ~new_n599 & new_n604;
  assign new_n1798 = new_n1797 ^ new_n1418;
  assign new_n1799 = ~new_n609 & new_n614;
  assign new_n1800 = new_n1799 ^ new_n1422;
  assign new_n1801 = ~new_n619 & new_n624;
  assign new_n1802 = new_n1801 ^ new_n1426;
  assign new_n1803 = ~new_n629 & new_n634;
  assign new_n1804 = new_n1803 ^ new_n1430;
  assign new_n1805 = ~new_n639 & new_n644;
  assign new_n1806 = new_n1805 ^ new_n1434;
  assign new_n1807 = ~new_n649 & new_n654;
  assign new_n1808 = new_n1807 ^ new_n1438;
  assign new_n1809 = ~new_n659 & new_n664;
  assign new_n1810 = new_n1809 ^ new_n1442;
  assign new_n1811 = ~new_n669 & new_n674;
  assign new_n1812 = new_n1811 ^ new_n1446;
  assign new_n1813 = ~new_n679 & new_n684;
  assign new_n1814 = new_n1813 ^ new_n1450;
  assign new_n1815 = ~new_n689 & new_n694;
  assign new_n1816 = new_n1815 ^ new_n1454;
  assign new_n1817 = ~new_n699 & new_n704;
  assign new_n1818 = new_n1817 ^ new_n1458;
  assign new_n1819 = ~new_n709 & new_n714;
  assign new_n1820 = new_n1819 ^ new_n1462;
  assign new_n1821 = ~new_n719 & new_n724;
  assign new_n1822 = new_n1821 ^ new_n1466;
  assign new_n1823 = ~new_n729 & new_n734;
  assign new_n1824 = new_n1823 ^ new_n1470;
  assign new_n1825 = ~new_n739 & new_n744;
  assign new_n1826 = new_n1825 ^ new_n1474;
  assign new_n1827 = ~new_n749 & new_n754;
  assign new_n1828 = new_n1827 ^ new_n1478;
  assign new_n1829 = ~new_n759 & new_n764;
  assign new_n1830 = new_n1829 ^ new_n1482;
  assign new_n1831 = ~new_n769 & new_n774;
  assign new_n1832 = new_n1831 ^ new_n1486;
  assign new_n1833 = ~new_n779 & new_n784;
  assign new_n1834 = new_n1833 ^ new_n1490;
  assign new_n1835 = ~new_n789 & new_n794;
  assign new_n1836 = new_n1835 ^ new_n1494;
  assign new_n1837 = ~new_n799 & new_n803;
  assign new_n1838 = new_n1837 ^ new_n1498;
  assign new_n1839 = ~new_n808 & new_n812;
  assign new_n1840 = new_n1839 ^ new_n1502;
  assign new_n1841 = ~new_n817 & new_n821;
  assign new_n1842 = new_n1841 ^ new_n1506;
  assign new_n1843 = ~new_n826 & new_n830;
  assign new_n1844 = new_n1843 ^ new_n1510;
  assign new_n1845 = ~new_n835 & new_n839;
  assign new_n1846 = new_n1845 ^ new_n1514;
  assign new_n1847 = ~new_n844 & new_n848;
  assign new_n1848 = new_n1847 ^ new_n1518;
  assign new_n1849 = ~new_n853 & new_n857;
  assign new_n1850 = new_n1849 ^ new_n1522;
  assign new_n1851 = ~new_n862 & new_n866;
  assign new_n1852 = new_n1851 ^ new_n1526;
  assign new_n1853 = ~new_n871 & new_n875;
  assign new_n1854 = new_n1853 ^ new_n1530;
  assign new_n1855 = ~new_n880 & new_n884;
  assign new_n1856 = new_n1855 ^ new_n1534;
  assign new_n1857 = ~new_n889 & new_n893;
  assign new_n1858 = new_n1857 ^ new_n1538;
  assign new_n1859 = ~new_n898 & new_n902;
  assign new_n1860 = new_n1859 ^ new_n1542;
  assign new_n1861 = ~new_n907 & new_n911;
  assign new_n1862 = new_n1861 ^ new_n1546;
  assign new_n1863 = ~new_n916 & new_n920;
  assign new_n1864 = new_n1863 ^ new_n1550;
  assign new_n1865 = ~new_n925 & new_n929;
  assign new_n1866 = new_n1865 ^ new_n1554;
  assign new_n1867 = ~new_n934 & new_n938;
  assign new_n1868 = new_n1867 ^ new_n1558;
  assign new_n1869 = ~new_n943 & new_n947;
  assign new_n1870 = new_n1869 ^ new_n1562;
  assign new_n1871 = ~new_n952 & new_n956;
  assign new_n1872 = new_n1871 ^ new_n1566;
  assign new_n1873 = ~new_n961 & new_n965;
  assign new_n1874 = new_n1873 ^ new_n1570;
  assign new_n1875 = ~new_n970 & new_n974;
  assign new_n1876 = new_n1875 ^ new_n1574;
  assign new_n1877 = ~new_n978 & new_n982;
  assign new_n1878 = new_n1877 ^ new_n1578;
  assign new_n1879 = ~new_n986 & new_n990;
  assign new_n1880 = new_n1879 ^ new_n1582;
  assign new_n1881 = ~new_n994 & new_n998;
  assign new_n1882 = new_n1881 ^ new_n1586;
  assign new_n1883 = ~new_n1002 & new_n1006;
  assign new_n1884 = new_n1883 ^ new_n1590;
  assign new_n1885 = ~new_n1010 & new_n1014;
  assign new_n1886 = new_n1885 ^ new_n1594;
  assign new_n1887 = ~new_n1018 & new_n1022;
  assign new_n1888 = new_n1887 ^ new_n1598;
  assign new_n1889 = ~new_n1026 & new_n1030;
  assign new_n1890 = new_n1889 ^ new_n1602;
  assign new_n1891 = ~new_n1034 & new_n1038;
  assign new_n1892 = new_n1891 ^ new_n1606;
  assign new_n1893 = ~new_n1042 & new_n1046;
  assign new_n1894 = new_n1893 ^ new_n1610;
  assign new_n1895 = ~new_n1050 & new_n1054;
  assign new_n1896 = new_n1895 ^ new_n1614;
  assign new_n1897 = ~new_n1058 & new_n1062;
  assign new_n1898 = new_n1897 ^ new_n1618;
  assign new_n1899 = ~new_n1066 & new_n1070;
  assign new_n1900 = new_n1899 ^ new_n1622;
  assign new_n1901 = ~new_n1074 & new_n1078;
  assign new_n1902 = new_n1901 ^ new_n1626;
  assign new_n1903 = ~new_n1082 & new_n1086;
  assign new_n1904 = new_n1903 ^ new_n1630;
  assign new_n1905 = ~new_n1090 & new_n1094;
  assign new_n1906 = new_n1905 ^ new_n1634;
  assign new_n1907 = ~new_n1098 & new_n1102;
  assign new_n1908 = new_n1907 ^ new_n1638;
  assign new_n1909 = ~new_n1106 & new_n1110;
  assign new_n1910 = new_n1909 ^ new_n1642;
  assign new_n1911 = ~new_n1114 & new_n1118;
  assign new_n1912 = new_n1911 ^ new_n1646;
  assign new_n1913 = ~new_n1122 & new_n1126;
  assign new_n1914 = new_n1913 ^ new_n1650;
  assign new_n1915 = ~new_n1130 & new_n1134;
  assign new_n1916 = new_n1915 ^ new_n1654;
  assign new_n1917 = ~new_n1138 & new_n1142;
  assign new_n1918 = new_n1917 ^ new_n1658;
  assign new_n1919 = ~new_n1146 & new_n1150;
  assign new_n1920 = new_n1919 ^ new_n1662;
  assign new_n1921 = ~new_n1433 & new_n609;
  assign new_n1922 = new_n1921 ^ new_n1181;
  assign new_n1923 = ~new_n1437 & new_n619;
  assign new_n1924 = new_n1923 ^ new_n1185;
  assign new_n1925 = ~new_n1441 & new_n629;
  assign new_n1926 = new_n1925 ^ new_n1189;
  assign new_n1927 = ~new_n1445 & new_n639;
  assign new_n1928 = new_n1927 ^ new_n1193;
  assign new_n1929 = ~new_n1449 & new_n649;
  assign new_n1930 = new_n1929 ^ new_n1197;
  assign new_n1931 = ~new_n1453 & new_n659;
  assign new_n1932 = new_n1931 ^ new_n1201;
  assign new_n1933 = ~new_n1457 & new_n669;
  assign new_n1934 = new_n1933 ^ new_n1205;
  assign new_n1935 = ~new_n1461 & new_n679;
  assign new_n1936 = new_n1935 ^ new_n1209;
  assign new_n1937 = ~new_n1465 & new_n689;
  assign new_n1938 = new_n1937 ^ new_n1213;
  assign new_n1939 = ~new_n1469 & new_n699;
  assign new_n1940 = new_n1939 ^ new_n1217;
  assign new_n1941 = ~new_n1473 & new_n709;
  assign new_n1942 = new_n1941 ^ new_n1221;
  assign new_n1943 = ~new_n1477 & new_n719;
  assign new_n1944 = new_n1943 ^ new_n1225;
  assign new_n1945 = ~new_n1481 & new_n729;
  assign new_n1946 = new_n1945 ^ new_n1229;
  assign new_n1947 = ~new_n1485 & new_n739;
  assign new_n1948 = new_n1947 ^ new_n1233;
  assign new_n1949 = ~new_n1489 & new_n749;
  assign new_n1950 = new_n1949 ^ new_n1237;
  assign new_n1951 = ~new_n1493 & new_n759;
  assign new_n1952 = new_n1951 ^ new_n1241;
  assign new_n1953 = ~new_n1497 & new_n769;
  assign new_n1954 = new_n1953 ^ new_n1245;
  assign new_n1955 = ~new_n1501 & new_n779;
  assign new_n1956 = new_n1955 ^ new_n1249;
  assign new_n1957 = ~new_n1505 & new_n789;
  assign new_n1958 = new_n1957 ^ new_n1253;
  assign new_n1959 = ~new_n1509 & new_n799;
  assign new_n1960 = new_n1959 ^ new_n1257;
  assign new_n1961 = ~new_n1513 & new_n808;
  assign new_n1962 = new_n1961 ^ new_n1261;
  assign new_n1963 = ~new_n1517 & new_n817;
  assign new_n1964 = new_n1963 ^ new_n1265;
  assign new_n1965 = ~new_n1521 & new_n826;
  assign new_n1966 = new_n1965 ^ new_n1269;
  assign new_n1967 = ~new_n1525 & new_n835;
  assign new_n1968 = new_n1967 ^ new_n1273;
  assign new_n1969 = ~new_n1529 & new_n844;
  assign new_n1970 = new_n1969 ^ new_n1277;
  assign new_n1971 = ~new_n1533 & new_n853;
  assign new_n1972 = new_n1971 ^ new_n1281;
  assign new_n1973 = ~new_n1537 & new_n862;
  assign new_n1974 = new_n1973 ^ new_n1285;
  assign new_n1975 = ~new_n1541 & new_n871;
  assign new_n1976 = new_n1975 ^ new_n1289;
  assign new_n1977 = ~new_n1545 & new_n880;
  assign new_n1978 = new_n1977 ^ new_n1293;
  assign new_n1979 = ~new_n1549 & new_n889;
  assign new_n1980 = new_n1979 ^ new_n1297;
  assign new_n1981 = ~new_n1553 & new_n898;
  assign new_n1982 = new_n1981 ^ new_n1301;
  assign new_n1983 = ~new_n1557 & new_n907;
  assign new_n1984 = new_n1983 ^ new_n1305;
  assign new_n1985 = ~new_n1561 & new_n916;
  assign new_n1986 = new_n1985 ^ new_n1309;
  assign new_n1987 = ~new_n1565 & new_n925;
  assign new_n1988 = new_n1987 ^ new_n1313;
  assign new_n1989 = ~new_n1569 & new_n934;
  assign new_n1990 = new_n1989 ^ new_n1317;
  assign new_n1991 = ~new_n1573 & new_n943;
  assign new_n1992 = new_n1991 ^ new_n1321;
  assign new_n1993 = ~new_n1577 & new_n952;
  assign new_n1994 = new_n1993 ^ new_n1325;
  assign new_n1995 = ~new_n1581 & new_n961;
  assign new_n1996 = new_n1995 ^ new_n1329;
  assign new_n1997 = ~new_n1585 & new_n970;
  assign new_n1998 = new_n1997 ^ new_n1333;
  assign new_n1999 = ~new_n1589 & new_n978;
  assign new_n2000 = new_n1999 ^ new_n1337;
  assign new_n2001 = ~new_n1593 & new_n986;
  assign new_n2002 = new_n2001 ^ new_n1341;
  assign new_n2003 = ~new_n1597 & new_n994;
  assign new_n2004 = new_n2003 ^ new_n1345;
  assign new_n2005 = ~new_n1601 & new_n1002;
  assign new_n2006 = new_n2005 ^ new_n1349;
  assign new_n2007 = ~new_n1605 & new_n1010;
  assign new_n2008 = new_n2007 ^ new_n1353;
  assign new_n2009 = ~new_n1609 & new_n1018;
  assign new_n2010 = new_n2009 ^ new_n1357;
  assign new_n2011 = ~new_n1613 & new_n1026;
  assign new_n2012 = new_n2011 ^ new_n1361;
  assign new_n2013 = ~new_n1617 & new_n1034;
  assign new_n2014 = new_n2013 ^ new_n1365;
  assign new_n2015 = ~new_n1621 & new_n1042;
  assign new_n2016 = new_n2015 ^ new_n1369;
  assign new_n2017 = ~new_n1625 & new_n1050;
  assign new_n2018 = new_n2017 ^ new_n1373;
  assign new_n2019 = ~new_n1629 & new_n1058;
  assign new_n2020 = new_n2019 ^ new_n1377;
  assign new_n2021 = ~new_n1633 & new_n1066;
  assign new_n2022 = new_n2021 ^ new_n1381;
  assign new_n2023 = ~new_n1637 & new_n1074;
  assign new_n2024 = new_n2023 ^ new_n1385;
  assign new_n2025 = ~new_n1641 & new_n1082;
  assign new_n2026 = new_n2025 ^ new_n1389;
  assign new_n2027 = ~new_n1645 & new_n1090;
  assign new_n2028 = new_n2027 ^ new_n1393;
  assign new_n2029 = ~new_n1649 & new_n1098;
  assign new_n2030 = new_n2029 ^ new_n1397;
  assign new_n2031 = ~new_n1653 & new_n1106;
  assign new_n2032 = new_n2031 ^ new_n1401;
  assign new_n2033 = ~new_n1657 & new_n1114;
  assign new_n2034 = new_n2033 ^ new_n1405;
  assign new_n2035 = ~new_n1661 & new_n1122;
  assign new_n2036 = new_n2035 ^ new_n1153;
  assign new_n2037 = ~new_n1409 & new_n1130;
  assign new_n2038 = new_n2037 ^ new_n1157;
  assign new_n2039 = ~new_n1413 & new_n1138;
  assign new_n2040 = new_n2039 ^ new_n1161;
  assign new_n2041 = ~new_n1417 & new_n1146;
  assign new_n2042 = new_n2041 ^ new_n1165;
  assign new_n2043 = ~new_n1421 & new_n579;
  assign new_n2044 = new_n2043 ^ new_n1169;
  assign new_n2045 = ~new_n1425 & new_n589;
  assign new_n2046 = new_n2045 ^ new_n1173;
  assign new_n2047 = ~new_n1429 & new_n599;
  assign new_n2048 = new_n2047 ^ new_n1177;
  assign new_n2049 = new_n594 ^ n334;
  assign new_n2050 = ~new_n609 & new_n2049;
  assign new_n2051 = new_n2050 ^ new_n1433;
  assign new_n2052 = new_n604 ^ n335;
  assign new_n2053 = ~new_n619 & new_n2052;
  assign new_n2054 = new_n2053 ^ new_n1437;
  assign new_n2055 = new_n614 ^ n336;
  assign new_n2056 = ~new_n629 & new_n2055;
  assign new_n2057 = new_n2056 ^ new_n1441;
  assign new_n2058 = new_n624 ^ n337;
  assign new_n2059 = ~new_n639 & new_n2058;
  assign new_n2060 = new_n2059 ^ new_n1445;
  assign new_n2061 = new_n634 ^ n338;
  assign new_n2062 = ~new_n649 & new_n2061;
  assign new_n2063 = new_n2062 ^ new_n1449;
  assign new_n2064 = new_n644 ^ n339;
  assign new_n2065 = ~new_n659 & new_n2064;
  assign new_n2066 = new_n2065 ^ new_n1453;
  assign new_n2067 = new_n654 ^ n340;
  assign new_n2068 = ~new_n669 & new_n2067;
  assign new_n2069 = new_n2068 ^ new_n1457;
  assign new_n2070 = new_n664 ^ n341;
  assign new_n2071 = ~new_n679 & new_n2070;
  assign new_n2072 = new_n2071 ^ new_n1461;
  assign new_n2073 = new_n674 ^ n342;
  assign new_n2074 = ~new_n689 & new_n2073;
  assign new_n2075 = new_n2074 ^ new_n1465;
  assign new_n2076 = new_n684 ^ n343;
  assign new_n2077 = ~new_n699 & new_n2076;
  assign new_n2078 = new_n2077 ^ new_n1469;
  assign new_n2079 = new_n694 ^ n344;
  assign new_n2080 = ~new_n709 & new_n2079;
  assign new_n2081 = new_n2080 ^ new_n1473;
  assign new_n2082 = new_n704 ^ n345;
  assign new_n2083 = ~new_n719 & new_n2082;
  assign new_n2084 = new_n2083 ^ new_n1477;
  assign new_n2085 = new_n714 ^ n346;
  assign new_n2086 = ~new_n729 & new_n2085;
  assign new_n2087 = new_n2086 ^ new_n1481;
  assign new_n2088 = new_n724 ^ n347;
  assign new_n2089 = ~new_n739 & new_n2088;
  assign new_n2090 = new_n2089 ^ new_n1485;
  assign new_n2091 = new_n734 ^ n348;
  assign new_n2092 = ~new_n749 & new_n2091;
  assign new_n2093 = new_n2092 ^ new_n1489;
  assign new_n2094 = new_n744 ^ n349;
  assign new_n2095 = ~new_n759 & new_n2094;
  assign new_n2096 = new_n2095 ^ new_n1493;
  assign new_n2097 = new_n754 ^ n350;
  assign new_n2098 = ~new_n769 & new_n2097;
  assign new_n2099 = new_n2098 ^ new_n1497;
  assign new_n2100 = new_n764 ^ n351;
  assign new_n2101 = ~new_n779 & new_n2100;
  assign new_n2102 = new_n2101 ^ new_n1501;
  assign new_n2103 = new_n774 ^ n352;
  assign new_n2104 = ~new_n789 & new_n2103;
  assign new_n2105 = new_n2104 ^ new_n1505;
  assign new_n2106 = new_n784 ^ n289;
  assign new_n2107 = ~new_n799 & new_n2106;
  assign new_n2108 = new_n2107 ^ new_n1509;
  assign new_n2109 = new_n794 ^ n290;
  assign new_n2110 = ~new_n808 & new_n2109;
  assign new_n2111 = new_n2110 ^ new_n1513;
  assign new_n2112 = new_n803 ^ n291;
  assign new_n2113 = ~new_n817 & new_n2112;
  assign new_n2114 = new_n2113 ^ new_n1517;
  assign new_n2115 = new_n812 ^ n292;
  assign new_n2116 = ~new_n826 & new_n2115;
  assign new_n2117 = new_n2116 ^ new_n1521;
  assign new_n2118 = new_n821 ^ n293;
  assign new_n2119 = ~new_n835 & new_n2118;
  assign new_n2120 = new_n2119 ^ new_n1525;
  assign new_n2121 = new_n830 ^ n294;
  assign new_n2122 = ~new_n844 & new_n2121;
  assign new_n2123 = new_n2122 ^ new_n1529;
  assign new_n2124 = new_n839 ^ n295;
  assign new_n2125 = ~new_n853 & new_n2124;
  assign new_n2126 = new_n2125 ^ new_n1533;
  assign new_n2127 = new_n848 ^ n296;
  assign new_n2128 = ~new_n862 & new_n2127;
  assign new_n2129 = new_n2128 ^ new_n1537;
  assign new_n2130 = new_n857 ^ n297;
  assign new_n2131 = ~new_n871 & new_n2130;
  assign new_n2132 = new_n2131 ^ new_n1541;
  assign new_n2133 = new_n866 ^ n298;
  assign new_n2134 = ~new_n880 & new_n2133;
  assign new_n2135 = new_n2134 ^ new_n1545;
  assign new_n2136 = new_n875 ^ n299;
  assign new_n2137 = ~new_n889 & new_n2136;
  assign new_n2138 = new_n2137 ^ new_n1549;
  assign new_n2139 = new_n884 ^ n300;
  assign new_n2140 = ~new_n898 & new_n2139;
  assign new_n2141 = new_n2140 ^ new_n1553;
  assign new_n2142 = new_n893 ^ n301;
  assign new_n2143 = ~new_n907 & new_n2142;
  assign new_n2144 = new_n2143 ^ new_n1557;
  assign new_n2145 = new_n902 ^ n302;
  assign new_n2146 = ~new_n916 & new_n2145;
  assign new_n2147 = new_n2146 ^ new_n1561;
  assign new_n2148 = new_n911 ^ n303;
  assign new_n2149 = ~new_n925 & new_n2148;
  assign new_n2150 = new_n2149 ^ new_n1565;
  assign new_n2151 = new_n920 ^ n304;
  assign new_n2152 = ~new_n934 & new_n2151;
  assign new_n2153 = new_n2152 ^ new_n1569;
  assign new_n2154 = new_n929 ^ n305;
  assign new_n2155 = ~new_n943 & new_n2154;
  assign new_n2156 = new_n2155 ^ new_n1573;
  assign new_n2157 = new_n938 ^ n306;
  assign new_n2158 = ~new_n952 & new_n2157;
  assign new_n2159 = new_n2158 ^ new_n1577;
  assign new_n2160 = new_n947 ^ n307;
  assign new_n2161 = ~new_n961 & new_n2160;
  assign new_n2162 = new_n2161 ^ new_n1581;
  assign new_n2163 = new_n956 ^ n308;
  assign new_n2164 = ~new_n970 & new_n2163;
  assign new_n2165 = new_n2164 ^ new_n1585;
  assign new_n2166 = new_n965 ^ n309;
  assign new_n2167 = ~new_n978 & new_n2166;
  assign new_n2168 = new_n2167 ^ new_n1589;
  assign new_n2169 = new_n974 ^ n310;
  assign new_n2170 = ~new_n986 & new_n2169;
  assign new_n2171 = new_n2170 ^ new_n1593;
  assign new_n2172 = new_n982 ^ n311;
  assign new_n2173 = ~new_n994 & new_n2172;
  assign new_n2174 = new_n2173 ^ new_n1597;
  assign new_n2175 = new_n990 ^ n312;
  assign new_n2176 = ~new_n1002 & new_n2175;
  assign new_n2177 = new_n2176 ^ new_n1601;
  assign new_n2178 = new_n998 ^ n313;
  assign new_n2179 = ~new_n1010 & new_n2178;
  assign new_n2180 = new_n2179 ^ new_n1605;
  assign new_n2181 = new_n1006 ^ n314;
  assign new_n2182 = ~new_n1018 & new_n2181;
  assign new_n2183 = new_n2182 ^ new_n1609;
  assign new_n2184 = new_n1014 ^ n315;
  assign new_n2185 = ~new_n1026 & new_n2184;
  assign new_n2186 = new_n2185 ^ new_n1613;
  assign new_n2187 = new_n1022 ^ n316;
  assign new_n2188 = ~new_n1034 & new_n2187;
  assign new_n2189 = new_n2188 ^ new_n1617;
  assign new_n2190 = new_n1030 ^ n317;
  assign new_n2191 = ~new_n1042 & new_n2190;
  assign new_n2192 = new_n2191 ^ new_n1621;
  assign new_n2193 = new_n1038 ^ n318;
  assign new_n2194 = ~new_n1050 & new_n2193;
  assign new_n2195 = new_n2194 ^ new_n1625;
  assign new_n2196 = new_n1046 ^ n319;
  assign new_n2197 = ~new_n1058 & new_n2196;
  assign new_n2198 = new_n2197 ^ new_n1629;
  assign new_n2199 = new_n1054 ^ n320;
  assign new_n2200 = ~new_n1066 & new_n2199;
  assign new_n2201 = new_n2200 ^ new_n1633;
  assign new_n2202 = new_n1062 ^ n321;
  assign new_n2203 = ~new_n1074 & new_n2202;
  assign new_n2204 = new_n2203 ^ new_n1637;
  assign new_n2205 = new_n1070 ^ n322;
  assign new_n2206 = ~new_n1082 & new_n2205;
  assign new_n2207 = new_n2206 ^ new_n1641;
  assign new_n2208 = new_n1078 ^ n323;
  assign new_n2209 = ~new_n1090 & new_n2208;
  assign new_n2210 = new_n2209 ^ new_n1645;
  assign new_n2211 = new_n1086 ^ n324;
  assign new_n2212 = ~new_n1098 & new_n2211;
  assign new_n2213 = new_n2212 ^ new_n1649;
  assign new_n2214 = new_n1094 ^ n325;
  assign new_n2215 = ~new_n1106 & new_n2214;
  assign new_n2216 = new_n2215 ^ new_n1653;
  assign new_n2217 = new_n1102 ^ n326;
  assign new_n2218 = ~new_n1114 & new_n2217;
  assign new_n2219 = new_n2218 ^ new_n1657;
  assign new_n2220 = new_n1110 ^ n327;
  assign new_n2221 = ~new_n1122 & new_n2220;
  assign new_n2222 = new_n2221 ^ new_n1661;
  assign new_n2223 = new_n1118 ^ n328;
  assign new_n2224 = ~new_n1130 & new_n2223;
  assign new_n2225 = new_n2224 ^ new_n1409;
  assign new_n2226 = new_n1126 ^ n329;
  assign new_n2227 = ~new_n1138 & new_n2226;
  assign new_n2228 = new_n2227 ^ new_n1413;
  assign new_n2229 = new_n1134 ^ n330;
  assign new_n2230 = ~new_n1146 & new_n2229;
  assign new_n2231 = new_n2230 ^ new_n1417;
  assign new_n2232 = new_n1142 ^ n331;
  assign new_n2233 = ~new_n579 & new_n2232;
  assign new_n2234 = new_n2233 ^ new_n1421;
  assign new_n2235 = new_n1150 ^ n332;
  assign new_n2236 = ~new_n589 & new_n2235;
  assign new_n2237 = new_n2236 ^ new_n1425;
  assign new_n2238 = new_n584 ^ n333;
  assign new_n2239 = ~new_n599 & new_n2238;
  assign new_n2240 = new_n2239 ^ new_n1429;
  assign new_n2241 = new_n762 ^ n158;
  assign new_n2242 = ~new_n2049 & new_n2241;
  assign new_n2243 = new_n2242 ^ new_n609;
  assign new_n2244 = new_n772 ^ n159;
  assign new_n2245 = ~new_n2052 & new_n2244;
  assign new_n2246 = new_n2245 ^ new_n619;
  assign new_n2247 = new_n782 ^ n160;
  assign new_n2248 = ~new_n2055 & new_n2247;
  assign new_n2249 = new_n2248 ^ new_n629;
  assign new_n2250 = new_n792 ^ n97;
  assign new_n2251 = ~new_n2058 & new_n2250;
  assign new_n2252 = new_n2251 ^ new_n639;
  assign new_n2253 = new_n801 ^ n98;
  assign new_n2254 = ~new_n2061 & new_n2253;
  assign new_n2255 = new_n2254 ^ new_n649;
  assign new_n2256 = new_n810 ^ n99;
  assign new_n2257 = ~new_n2064 & new_n2256;
  assign new_n2258 = new_n2257 ^ new_n659;
  assign new_n2259 = new_n819 ^ n100;
  assign new_n2260 = ~new_n2067 & new_n2259;
  assign new_n2261 = new_n2260 ^ new_n669;
  assign new_n2262 = new_n828 ^ n101;
  assign new_n2263 = ~new_n2070 & new_n2262;
  assign new_n2264 = new_n2263 ^ new_n679;
  assign new_n2265 = new_n837 ^ n102;
  assign new_n2266 = ~new_n2073 & new_n2265;
  assign new_n2267 = new_n2266 ^ new_n689;
  assign new_n2268 = new_n846 ^ n103;
  assign new_n2269 = ~new_n2076 & new_n2268;
  assign new_n2270 = new_n2269 ^ new_n699;
  assign new_n2271 = new_n855 ^ n104;
  assign new_n2272 = ~new_n2079 & new_n2271;
  assign new_n2273 = new_n2272 ^ new_n709;
  assign new_n2274 = new_n864 ^ n105;
  assign new_n2275 = ~new_n2082 & new_n2274;
  assign new_n2276 = new_n2275 ^ new_n719;
  assign new_n2277 = new_n873 ^ n106;
  assign new_n2278 = ~new_n2085 & new_n2277;
  assign new_n2279 = new_n2278 ^ new_n729;
  assign new_n2280 = new_n882 ^ n107;
  assign new_n2281 = ~new_n2088 & new_n2280;
  assign new_n2282 = new_n2281 ^ new_n739;
  assign new_n2283 = new_n891 ^ n108;
  assign new_n2284 = ~new_n2091 & new_n2283;
  assign new_n2285 = new_n2284 ^ new_n749;
  assign new_n2286 = new_n900 ^ n109;
  assign new_n2287 = ~new_n2094 & new_n2286;
  assign new_n2288 = new_n2287 ^ new_n759;
  assign new_n2289 = new_n909 ^ n110;
  assign new_n2290 = ~new_n2097 & new_n2289;
  assign new_n2291 = new_n2290 ^ new_n769;
  assign new_n2292 = new_n918 ^ n111;
  assign new_n2293 = ~new_n2100 & new_n2292;
  assign new_n2294 = new_n2293 ^ new_n779;
  assign new_n2295 = new_n927 ^ n112;
  assign new_n2296 = ~new_n2103 & new_n2295;
  assign new_n2297 = new_n2296 ^ new_n789;
  assign new_n2298 = new_n936 ^ n113;
  assign new_n2299 = ~new_n2106 & new_n2298;
  assign new_n2300 = new_n2299 ^ new_n799;
  assign new_n2301 = new_n945 ^ n114;
  assign new_n2302 = ~new_n2109 & new_n2301;
  assign new_n2303 = new_n2302 ^ new_n808;
  assign new_n2304 = new_n954 ^ n115;
  assign new_n2305 = ~new_n2112 & new_n2304;
  assign new_n2306 = new_n2305 ^ new_n817;
  assign new_n2307 = new_n963 ^ n116;
  assign new_n2308 = ~new_n2115 & new_n2307;
  assign new_n2309 = new_n2308 ^ new_n826;
  assign new_n2310 = new_n972 ^ n117;
  assign new_n2311 = ~new_n2118 & new_n2310;
  assign new_n2312 = new_n2311 ^ new_n835;
  assign new_n2313 = new_n980 ^ n118;
  assign new_n2314 = ~new_n2121 & new_n2313;
  assign new_n2315 = new_n2314 ^ new_n844;
  assign new_n2316 = new_n988 ^ n119;
  assign new_n2317 = ~new_n2124 & new_n2316;
  assign new_n2318 = new_n2317 ^ new_n853;
  assign new_n2319 = new_n996 ^ n120;
  assign new_n2320 = ~new_n2127 & new_n2319;
  assign new_n2321 = new_n2320 ^ new_n862;
  assign new_n2322 = new_n1004 ^ n121;
  assign new_n2323 = ~new_n2130 & new_n2322;
  assign new_n2324 = new_n2323 ^ new_n871;
  assign new_n2325 = new_n1012 ^ n122;
  assign new_n2326 = ~new_n2133 & new_n2325;
  assign new_n2327 = new_n2326 ^ new_n880;
  assign new_n2328 = new_n1020 ^ n123;
  assign new_n2329 = ~new_n2136 & new_n2328;
  assign new_n2330 = new_n2329 ^ new_n889;
  assign new_n2331 = new_n1028 ^ n124;
  assign new_n2332 = ~new_n2139 & new_n2331;
  assign new_n2333 = new_n2332 ^ new_n898;
  assign new_n2334 = new_n1036 ^ n125;
  assign new_n2335 = ~new_n2142 & new_n2334;
  assign new_n2336 = new_n2335 ^ new_n907;
  assign new_n2337 = new_n1044 ^ n126;
  assign new_n2338 = ~new_n2145 & new_n2337;
  assign new_n2339 = new_n2338 ^ new_n916;
  assign new_n2340 = new_n1052 ^ n127;
  assign new_n2341 = ~new_n2148 & new_n2340;
  assign new_n2342 = new_n2341 ^ new_n925;
  assign new_n2343 = new_n1060 ^ n128;
  assign new_n2344 = ~new_n2151 & new_n2343;
  assign new_n2345 = new_n2344 ^ new_n934;
  assign new_n2346 = new_n1068 ^ n129;
  assign new_n2347 = ~new_n2154 & new_n2346;
  assign new_n2348 = new_n2347 ^ new_n943;
  assign new_n2349 = new_n1076 ^ n130;
  assign new_n2350 = ~new_n2157 & new_n2349;
  assign new_n2351 = new_n2350 ^ new_n952;
  assign new_n2352 = new_n1084 ^ n131;
  assign new_n2353 = ~new_n2160 & new_n2352;
  assign new_n2354 = new_n2353 ^ new_n961;
  assign new_n2355 = new_n1092 ^ n132;
  assign new_n2356 = ~new_n2163 & new_n2355;
  assign new_n2357 = new_n2356 ^ new_n970;
  assign new_n2358 = new_n1100 ^ n133;
  assign new_n2359 = ~new_n2166 & new_n2358;
  assign new_n2360 = new_n2359 ^ new_n978;
  assign new_n2361 = new_n1108 ^ n134;
  assign new_n2362 = ~new_n2169 & new_n2361;
  assign new_n2363 = new_n2362 ^ new_n986;
  assign new_n2364 = new_n1116 ^ n135;
  assign new_n2365 = ~new_n2172 & new_n2364;
  assign new_n2366 = new_n2365 ^ new_n994;
  assign new_n2367 = new_n1124 ^ n136;
  assign new_n2368 = ~new_n2175 & new_n2367;
  assign new_n2369 = new_n2368 ^ new_n1002;
  assign new_n2370 = new_n1132 ^ n137;
  assign new_n2371 = ~new_n2178 & new_n2370;
  assign new_n2372 = new_n2371 ^ new_n1010;
  assign new_n2373 = new_n1140 ^ n138;
  assign new_n2374 = ~new_n2181 & new_n2373;
  assign new_n2375 = new_n2374 ^ new_n1018;
  assign new_n2376 = new_n1148 ^ n139;
  assign new_n2377 = ~new_n2184 & new_n2376;
  assign new_n2378 = new_n2377 ^ new_n1026;
  assign new_n2379 = new_n582 ^ n140;
  assign new_n2380 = ~new_n2187 & new_n2379;
  assign new_n2381 = new_n2380 ^ new_n1034;
  assign new_n2382 = new_n592 ^ n141;
  assign new_n2383 = ~new_n2190 & new_n2382;
  assign new_n2384 = new_n2383 ^ new_n1042;
  assign new_n2385 = new_n602 ^ n142;
  assign new_n2386 = ~new_n2193 & new_n2385;
  assign new_n2387 = new_n2386 ^ new_n1050;
  assign new_n2388 = new_n612 ^ n143;
  assign new_n2389 = ~new_n2196 & new_n2388;
  assign new_n2390 = new_n2389 ^ new_n1058;
  assign new_n2391 = new_n622 ^ n144;
  assign new_n2392 = ~new_n2199 & new_n2391;
  assign new_n2393 = new_n2392 ^ new_n1066;
  assign new_n2394 = new_n632 ^ n145;
  assign new_n2395 = ~new_n2202 & new_n2394;
  assign new_n2396 = new_n2395 ^ new_n1074;
  assign new_n2397 = new_n642 ^ n146;
  assign new_n2398 = ~new_n2205 & new_n2397;
  assign new_n2399 = new_n2398 ^ new_n1082;
  assign new_n2400 = new_n652 ^ n147;
  assign new_n2401 = ~new_n2208 & new_n2400;
  assign new_n2402 = new_n2401 ^ new_n1090;
  assign new_n2403 = new_n662 ^ n148;
  assign new_n2404 = ~new_n2211 & new_n2403;
  assign new_n2405 = new_n2404 ^ new_n1098;
  assign new_n2406 = new_n672 ^ n149;
  assign new_n2407 = ~new_n2214 & new_n2406;
  assign new_n2408 = new_n2407 ^ new_n1106;
  assign new_n2409 = new_n682 ^ n150;
  assign new_n2410 = ~new_n2217 & new_n2409;
  assign new_n2411 = new_n2410 ^ new_n1114;
  assign new_n2412 = new_n692 ^ n151;
  assign new_n2413 = ~new_n2220 & new_n2412;
  assign new_n2414 = new_n2413 ^ new_n1122;
  assign new_n2415 = new_n702 ^ n152;
  assign new_n2416 = ~new_n2223 & new_n2415;
  assign new_n2417 = new_n2416 ^ new_n1130;
  assign new_n2418 = new_n712 ^ n153;
  assign new_n2419 = ~new_n2226 & new_n2418;
  assign new_n2420 = new_n2419 ^ new_n1138;
  assign new_n2421 = new_n722 ^ n154;
  assign new_n2422 = ~new_n2229 & new_n2421;
  assign new_n2423 = new_n2422 ^ new_n1146;
  assign new_n2424 = new_n732 ^ n155;
  assign new_n2425 = ~new_n2232 & new_n2424;
  assign new_n2426 = new_n2425 ^ new_n579;
  assign new_n2427 = new_n742 ^ n156;
  assign new_n2428 = ~new_n2235 & new_n2427;
  assign new_n2429 = new_n2428 ^ new_n589;
  assign new_n2430 = new_n752 ^ n157;
  assign new_n2431 = ~new_n2238 & new_n2430;
  assign new_n2432 = new_n2431 ^ new_n599;
  assign new_n2433 = ~new_n2241 & new_n1181;
  assign new_n2434 = new_n2433 ^ new_n2049;
  assign new_n2435 = ~new_n2244 & new_n1185;
  assign new_n2436 = new_n2435 ^ new_n2052;
  assign new_n2437 = ~new_n2247 & new_n1189;
  assign new_n2438 = new_n2437 ^ new_n2055;
  assign new_n2439 = ~new_n2250 & new_n1193;
  assign new_n2440 = new_n2439 ^ new_n2058;
  assign new_n2441 = ~new_n2253 & new_n1197;
  assign new_n2442 = new_n2441 ^ new_n2061;
  assign new_n2443 = ~new_n2256 & new_n1201;
  assign new_n2444 = new_n2443 ^ new_n2064;
  assign new_n2445 = ~new_n2259 & new_n1205;
  assign new_n2446 = new_n2445 ^ new_n2067;
  assign new_n2447 = ~new_n2262 & new_n1209;
  assign new_n2448 = new_n2447 ^ new_n2070;
  assign new_n2449 = ~new_n2265 & new_n1213;
  assign new_n2450 = new_n2449 ^ new_n2073;
  assign new_n2451 = ~new_n2268 & new_n1217;
  assign new_n2452 = new_n2451 ^ new_n2076;
  assign new_n2453 = ~new_n2271 & new_n1221;
  assign new_n2454 = new_n2453 ^ new_n2079;
  assign new_n2455 = ~new_n2274 & new_n1225;
  assign new_n2456 = new_n2455 ^ new_n2082;
  assign new_n2457 = ~new_n2277 & new_n1229;
  assign new_n2458 = new_n2457 ^ new_n2085;
  assign new_n2459 = ~new_n2280 & new_n1233;
  assign new_n2460 = new_n2459 ^ new_n2088;
  assign new_n2461 = ~new_n2283 & new_n1237;
  assign new_n2462 = new_n2461 ^ new_n2091;
  assign new_n2463 = ~new_n2286 & new_n1241;
  assign new_n2464 = new_n2463 ^ new_n2094;
  assign new_n2465 = ~new_n2289 & new_n1245;
  assign new_n2466 = new_n2465 ^ new_n2097;
  assign new_n2467 = ~new_n2292 & new_n1249;
  assign new_n2468 = new_n2467 ^ new_n2100;
  assign new_n2469 = ~new_n2295 & new_n1253;
  assign new_n2470 = new_n2469 ^ new_n2103;
  assign new_n2471 = ~new_n2298 & new_n1257;
  assign new_n2472 = new_n2471 ^ new_n2106;
  assign new_n2473 = ~new_n2301 & new_n1261;
  assign new_n2474 = new_n2473 ^ new_n2109;
  assign new_n2475 = ~new_n2304 & new_n1265;
  assign new_n2476 = new_n2475 ^ new_n2112;
  assign new_n2477 = ~new_n2307 & new_n1269;
  assign new_n2478 = new_n2477 ^ new_n2115;
  assign new_n2479 = ~new_n2310 & new_n1273;
  assign new_n2480 = new_n2479 ^ new_n2118;
  assign new_n2481 = ~new_n2313 & new_n1277;
  assign new_n2482 = new_n2481 ^ new_n2121;
  assign new_n2483 = ~new_n2316 & new_n1281;
  assign new_n2484 = new_n2483 ^ new_n2124;
  assign new_n2485 = ~new_n2319 & new_n1285;
  assign new_n2486 = new_n2485 ^ new_n2127;
  assign new_n2487 = ~new_n2322 & new_n1289;
  assign new_n2488 = new_n2487 ^ new_n2130;
  assign new_n2489 = ~new_n2325 & new_n1293;
  assign new_n2490 = new_n2489 ^ new_n2133;
  assign new_n2491 = ~new_n2328 & new_n1297;
  assign new_n2492 = new_n2491 ^ new_n2136;
  assign new_n2493 = ~new_n2331 & new_n1301;
  assign new_n2494 = new_n2493 ^ new_n2139;
  assign new_n2495 = ~new_n2334 & new_n1305;
  assign new_n2496 = new_n2495 ^ new_n2142;
  assign new_n2497 = ~new_n2337 & new_n1309;
  assign new_n2498 = new_n2497 ^ new_n2145;
  assign new_n2499 = ~new_n2340 & new_n1313;
  assign new_n2500 = new_n2499 ^ new_n2148;
  assign new_n2501 = ~new_n2343 & new_n1317;
  assign new_n2502 = new_n2501 ^ new_n2151;
  assign new_n2503 = ~new_n2346 & new_n1321;
  assign new_n2504 = new_n2503 ^ new_n2154;
  assign new_n2505 = ~new_n2349 & new_n1325;
  assign new_n2506 = new_n2505 ^ new_n2157;
  assign new_n2507 = ~new_n2352 & new_n1329;
  assign new_n2508 = new_n2507 ^ new_n2160;
  assign new_n2509 = ~new_n2355 & new_n1333;
  assign new_n2510 = new_n2509 ^ new_n2163;
  assign new_n2511 = ~new_n2358 & new_n1337;
  assign new_n2512 = new_n2511 ^ new_n2166;
  assign new_n2513 = ~new_n2361 & new_n1341;
  assign new_n2514 = new_n2513 ^ new_n2169;
  assign new_n2515 = ~new_n2364 & new_n1345;
  assign new_n2516 = new_n2515 ^ new_n2172;
  assign new_n2517 = ~new_n2367 & new_n1349;
  assign new_n2518 = new_n2517 ^ new_n2175;
  assign new_n2519 = ~new_n2370 & new_n1353;
  assign new_n2520 = new_n2519 ^ new_n2178;
  assign new_n2521 = ~new_n2373 & new_n1357;
  assign new_n2522 = new_n2521 ^ new_n2181;
  assign new_n2523 = ~new_n2376 & new_n1361;
  assign new_n2524 = new_n2523 ^ new_n2184;
  assign new_n2525 = ~new_n2379 & new_n1365;
  assign new_n2526 = new_n2525 ^ new_n2187;
  assign new_n2527 = ~new_n2382 & new_n1369;
  assign new_n2528 = new_n2527 ^ new_n2190;
  assign new_n2529 = ~new_n2385 & new_n1373;
  assign new_n2530 = new_n2529 ^ new_n2193;
  assign new_n2531 = ~new_n2388 & new_n1377;
  assign new_n2532 = new_n2531 ^ new_n2196;
  assign new_n2533 = ~new_n2391 & new_n1381;
  assign new_n2534 = new_n2533 ^ new_n2199;
  assign new_n2535 = ~new_n2394 & new_n1385;
  assign new_n2536 = new_n2535 ^ new_n2202;
  assign new_n2537 = ~new_n2397 & new_n1389;
  assign new_n2538 = new_n2537 ^ new_n2205;
  assign new_n2539 = ~new_n2400 & new_n1393;
  assign new_n2540 = new_n2539 ^ new_n2208;
  assign new_n2541 = ~new_n2403 & new_n1397;
  assign new_n2542 = new_n2541 ^ new_n2211;
  assign new_n2543 = ~new_n2406 & new_n1401;
  assign new_n2544 = new_n2543 ^ new_n2214;
  assign new_n2545 = ~new_n2409 & new_n1405;
  assign new_n2546 = new_n2545 ^ new_n2217;
  assign new_n2547 = ~new_n2412 & new_n1153;
  assign new_n2548 = new_n2547 ^ new_n2220;
  assign new_n2549 = ~new_n2415 & new_n1157;
  assign new_n2550 = new_n2549 ^ new_n2223;
  assign new_n2551 = ~new_n2418 & new_n1161;
  assign new_n2552 = new_n2551 ^ new_n2226;
  assign new_n2553 = ~new_n2421 & new_n1165;
  assign new_n2554 = new_n2553 ^ new_n2229;
  assign new_n2555 = ~new_n2424 & new_n1169;
  assign new_n2556 = new_n2555 ^ new_n2232;
  assign new_n2557 = ~new_n2427 & new_n1173;
  assign new_n2558 = new_n2557 ^ new_n2235;
  assign new_n2559 = ~new_n2430 & new_n1177;
  assign new_n2560 = new_n2559 ^ new_n2238;
  assign new_n2561 = ~new_n1181 & new_n1433;
  assign new_n2562 = new_n2561 ^ new_n2241;
  assign new_n2563 = ~new_n1185 & new_n1437;
  assign new_n2564 = new_n2563 ^ new_n2244;
  assign new_n2565 = ~new_n1189 & new_n1441;
  assign new_n2566 = new_n2565 ^ new_n2247;
  assign new_n2567 = ~new_n1193 & new_n1445;
  assign new_n2568 = new_n2567 ^ new_n2250;
  assign new_n2569 = ~new_n1197 & new_n1449;
  assign new_n2570 = new_n2569 ^ new_n2253;
  assign new_n2571 = ~new_n1201 & new_n1453;
  assign new_n2572 = new_n2571 ^ new_n2256;
  assign new_n2573 = ~new_n1205 & new_n1457;
  assign new_n2574 = new_n2573 ^ new_n2259;
  assign new_n2575 = ~new_n1209 & new_n1461;
  assign new_n2576 = new_n2575 ^ new_n2262;
  assign new_n2577 = ~new_n1213 & new_n1465;
  assign new_n2578 = new_n2577 ^ new_n2265;
  assign new_n2579 = ~new_n1217 & new_n1469;
  assign new_n2580 = new_n2579 ^ new_n2268;
  assign new_n2581 = ~new_n1221 & new_n1473;
  assign new_n2582 = new_n2581 ^ new_n2271;
  assign new_n2583 = ~new_n1225 & new_n1477;
  assign new_n2584 = new_n2583 ^ new_n2274;
  assign new_n2585 = ~new_n1229 & new_n1481;
  assign new_n2586 = new_n2585 ^ new_n2277;
  assign new_n2587 = ~new_n1233 & new_n1485;
  assign new_n2588 = new_n2587 ^ new_n2280;
  assign new_n2589 = ~new_n1237 & new_n1489;
  assign new_n2590 = new_n2589 ^ new_n2283;
  assign new_n2591 = ~new_n1241 & new_n1493;
  assign new_n2592 = new_n2591 ^ new_n2286;
  assign new_n2593 = ~new_n1245 & new_n1497;
  assign new_n2594 = new_n2593 ^ new_n2289;
  assign new_n2595 = ~new_n1249 & new_n1501;
  assign new_n2596 = new_n2595 ^ new_n2292;
  assign new_n2597 = ~new_n1253 & new_n1505;
  assign new_n2598 = new_n2597 ^ new_n2295;
  assign new_n2599 = ~new_n1257 & new_n1509;
  assign new_n2600 = new_n2599 ^ new_n2298;
  assign new_n2601 = ~new_n1261 & new_n1513;
  assign new_n2602 = new_n2601 ^ new_n2301;
  assign new_n2603 = ~new_n1265 & new_n1517;
  assign new_n2604 = new_n2603 ^ new_n2304;
  assign new_n2605 = ~new_n1269 & new_n1521;
  assign new_n2606 = new_n2605 ^ new_n2307;
  assign new_n2607 = ~new_n1273 & new_n1525;
  assign new_n2608 = new_n2607 ^ new_n2310;
  assign new_n2609 = ~new_n1277 & new_n1529;
  assign new_n2610 = new_n2609 ^ new_n2313;
  assign new_n2611 = ~new_n1281 & new_n1533;
  assign new_n2612 = new_n2611 ^ new_n2316;
  assign new_n2613 = ~new_n1285 & new_n1537;
  assign new_n2614 = new_n2613 ^ new_n2319;
  assign new_n2615 = ~new_n1289 & new_n1541;
  assign new_n2616 = new_n2615 ^ new_n2322;
  assign new_n2617 = ~new_n1293 & new_n1545;
  assign new_n2618 = new_n2617 ^ new_n2325;
  assign new_n2619 = ~new_n1297 & new_n1549;
  assign new_n2620 = new_n2619 ^ new_n2328;
  assign new_n2621 = ~new_n1301 & new_n1553;
  assign new_n2622 = new_n2621 ^ new_n2331;
  assign new_n2623 = ~new_n1305 & new_n1557;
  assign new_n2624 = new_n2623 ^ new_n2334;
  assign new_n2625 = ~new_n1309 & new_n1561;
  assign new_n2626 = new_n2625 ^ new_n2337;
  assign new_n2627 = ~new_n1313 & new_n1565;
  assign new_n2628 = new_n2627 ^ new_n2340;
  assign new_n2629 = ~new_n1317 & new_n1569;
  assign new_n2630 = new_n2629 ^ new_n2343;
  assign new_n2631 = ~new_n1321 & new_n1573;
  assign new_n2632 = new_n2631 ^ new_n2346;
  assign new_n2633 = ~new_n1325 & new_n1577;
  assign new_n2634 = new_n2633 ^ new_n2349;
  assign new_n2635 = ~new_n1329 & new_n1581;
  assign new_n2636 = new_n2635 ^ new_n2352;
  assign new_n2637 = ~new_n1333 & new_n1585;
  assign new_n2638 = new_n2637 ^ new_n2355;
  assign new_n2639 = ~new_n1337 & new_n1589;
  assign new_n2640 = new_n2639 ^ new_n2358;
  assign new_n2641 = ~new_n1341 & new_n1593;
  assign new_n2642 = new_n2641 ^ new_n2361;
  assign new_n2643 = ~new_n1345 & new_n1597;
  assign new_n2644 = new_n2643 ^ new_n2364;
  assign new_n2645 = ~new_n1349 & new_n1601;
  assign new_n2646 = new_n2645 ^ new_n2367;
  assign new_n2647 = ~new_n1353 & new_n1605;
  assign new_n2648 = new_n2647 ^ new_n2370;
  assign new_n2649 = ~new_n1357 & new_n1609;
  assign new_n2650 = new_n2649 ^ new_n2373;
  assign new_n2651 = ~new_n1361 & new_n1613;
  assign new_n2652 = new_n2651 ^ new_n2376;
  assign new_n2653 = ~new_n1365 & new_n1617;
  assign new_n2654 = new_n2653 ^ new_n2379;
  assign new_n2655 = ~new_n1369 & new_n1621;
  assign new_n2656 = new_n2655 ^ new_n2382;
  assign new_n2657 = ~new_n1373 & new_n1625;
  assign new_n2658 = new_n2657 ^ new_n2385;
  assign new_n2659 = ~new_n1377 & new_n1629;
  assign new_n2660 = new_n2659 ^ new_n2388;
  assign new_n2661 = ~new_n1381 & new_n1633;
  assign new_n2662 = new_n2661 ^ new_n2391;
  assign new_n2663 = ~new_n1385 & new_n1637;
  assign new_n2664 = new_n2663 ^ new_n2394;
  assign new_n2665 = ~new_n1389 & new_n1641;
  assign new_n2666 = new_n2665 ^ new_n2397;
  assign new_n2667 = ~new_n1393 & new_n1645;
  assign new_n2668 = new_n2667 ^ new_n2400;
  assign new_n2669 = ~new_n1397 & new_n1649;
  assign new_n2670 = new_n2669 ^ new_n2403;
  assign new_n2671 = ~new_n1401 & new_n1653;
  assign new_n2672 = new_n2671 ^ new_n2406;
  assign new_n2673 = ~new_n1405 & new_n1657;
  assign new_n2674 = new_n2673 ^ new_n2409;
  assign new_n2675 = ~new_n1153 & new_n1661;
  assign new_n2676 = new_n2675 ^ new_n2412;
  assign new_n2677 = ~new_n1157 & new_n1409;
  assign new_n2678 = new_n2677 ^ new_n2415;
  assign new_n2679 = ~new_n1161 & new_n1413;
  assign new_n2680 = new_n2679 ^ new_n2418;
  assign new_n2681 = ~new_n1165 & new_n1417;
  assign new_n2682 = new_n2681 ^ new_n2421;
  assign new_n2683 = ~new_n1169 & new_n1421;
  assign new_n2684 = new_n2683 ^ new_n2424;
  assign new_n2685 = ~new_n1173 & new_n1425;
  assign new_n2686 = new_n2685 ^ new_n2427;
  assign new_n2687 = ~new_n1177 & new_n1429;
  assign new_n2688 = new_n2687 ^ new_n2430;
  assign new_n2689 = ~new_n846 & new_n1169;
  assign new_n2690 = new_n2689 ^ new_n794;
  assign new_n2691 = ~new_n855 & new_n1173;
  assign new_n2692 = new_n2691 ^ new_n803;
  assign new_n2693 = ~new_n864 & new_n1177;
  assign new_n2694 = new_n2693 ^ new_n812;
  assign new_n2695 = ~new_n873 & new_n1181;
  assign new_n2696 = new_n2695 ^ new_n821;
  assign new_n2697 = ~new_n882 & new_n1185;
  assign new_n2698 = new_n2697 ^ new_n830;
  assign new_n2699 = ~new_n891 & new_n1189;
  assign new_n2700 = new_n2699 ^ new_n839;
  assign new_n2701 = ~new_n900 & new_n1193;
  assign new_n2702 = new_n2701 ^ new_n848;
  assign new_n2703 = ~new_n909 & new_n1197;
  assign new_n2704 = new_n2703 ^ new_n857;
  assign new_n2705 = ~new_n918 & new_n1201;
  assign new_n2706 = new_n2705 ^ new_n866;
  assign new_n2707 = ~new_n927 & new_n1205;
  assign new_n2708 = new_n2707 ^ new_n875;
  assign new_n2709 = ~new_n936 & new_n1209;
  assign new_n2710 = new_n2709 ^ new_n884;
  assign new_n2711 = ~new_n945 & new_n1213;
  assign new_n2712 = new_n2711 ^ new_n893;
  assign new_n2713 = ~new_n954 & new_n1217;
  assign new_n2714 = new_n2713 ^ new_n902;
  assign new_n2715 = ~new_n963 & new_n1221;
  assign new_n2716 = new_n2715 ^ new_n911;
  assign new_n2717 = ~new_n972 & new_n1225;
  assign new_n2718 = new_n2717 ^ new_n920;
  assign new_n2719 = ~new_n980 & new_n1229;
  assign new_n2720 = new_n2719 ^ new_n929;
  assign new_n2721 = ~new_n988 & new_n1233;
  assign new_n2722 = new_n2721 ^ new_n938;
  assign new_n2723 = ~new_n996 & new_n1237;
  assign new_n2724 = new_n2723 ^ new_n947;
  assign new_n2725 = ~new_n1004 & new_n1241;
  assign new_n2726 = new_n2725 ^ new_n956;
  assign new_n2727 = ~new_n1012 & new_n1245;
  assign new_n2728 = new_n2727 ^ new_n965;
  assign new_n2729 = ~new_n1020 & new_n1249;
  assign new_n2730 = new_n2729 ^ new_n974;
  assign new_n2731 = ~new_n1028 & new_n1253;
  assign new_n2732 = new_n2731 ^ new_n982;
  assign new_n2733 = ~new_n1036 & new_n1257;
  assign new_n2734 = new_n2733 ^ new_n990;
  assign new_n2735 = ~new_n1044 & new_n1261;
  assign new_n2736 = new_n2735 ^ new_n998;
  assign new_n2737 = ~new_n1052 & new_n1265;
  assign new_n2738 = new_n2737 ^ new_n1006;
  assign new_n2739 = ~new_n1060 & new_n1269;
  assign new_n2740 = new_n2739 ^ new_n1014;
  assign new_n2741 = ~new_n1068 & new_n1273;
  assign new_n2742 = new_n2741 ^ new_n1022;
  assign new_n2743 = ~new_n1076 & new_n1277;
  assign new_n2744 = new_n2743 ^ new_n1030;
  assign new_n2745 = ~new_n1084 & new_n1281;
  assign new_n2746 = new_n2745 ^ new_n1038;
  assign new_n2747 = ~new_n1092 & new_n1285;
  assign new_n2748 = new_n2747 ^ new_n1046;
  assign new_n2749 = ~new_n1100 & new_n1289;
  assign new_n2750 = new_n2749 ^ new_n1054;
  assign new_n2751 = ~new_n1108 & new_n1293;
  assign new_n2752 = new_n2751 ^ new_n1062;
  assign new_n2753 = ~new_n1116 & new_n1297;
  assign new_n2754 = new_n2753 ^ new_n1070;
  assign new_n2755 = ~new_n1124 & new_n1301;
  assign new_n2756 = new_n2755 ^ new_n1078;
  assign new_n2757 = ~new_n1132 & new_n1305;
  assign new_n2758 = new_n2757 ^ new_n1086;
  assign new_n2759 = ~new_n1140 & new_n1309;
  assign new_n2760 = new_n2759 ^ new_n1094;
  assign new_n2761 = ~new_n1148 & new_n1313;
  assign new_n2762 = new_n2761 ^ new_n1102;
  assign new_n2763 = ~new_n582 & new_n1317;
  assign new_n2764 = new_n2763 ^ new_n1110;
  assign new_n2765 = ~new_n592 & new_n1321;
  assign new_n2766 = new_n2765 ^ new_n1118;
  assign new_n2767 = ~new_n602 & new_n1325;
  assign new_n2768 = new_n2767 ^ new_n1126;
  assign new_n2769 = ~new_n612 & new_n1329;
  assign new_n2770 = new_n2769 ^ new_n1134;
  assign new_n2771 = ~new_n622 & new_n1333;
  assign new_n2772 = new_n2771 ^ new_n1142;
  assign new_n2773 = ~new_n632 & new_n1337;
  assign new_n2774 = new_n2773 ^ new_n1150;
  assign new_n2775 = ~new_n642 & new_n1341;
  assign new_n2776 = new_n2775 ^ new_n584;
  assign new_n2777 = ~new_n652 & new_n1345;
  assign new_n2778 = new_n2777 ^ new_n594;
  assign new_n2779 = ~new_n662 & new_n1349;
  assign new_n2780 = new_n2779 ^ new_n604;
  assign new_n2781 = ~new_n672 & new_n1353;
  assign new_n2782 = new_n2781 ^ new_n614;
  assign new_n2783 = ~new_n682 & new_n1357;
  assign new_n2784 = new_n2783 ^ new_n624;
  assign new_n2785 = ~new_n692 & new_n1361;
  assign new_n2786 = new_n2785 ^ new_n634;
  assign new_n2787 = ~new_n702 & new_n1365;
  assign new_n2788 = new_n2787 ^ new_n644;
  assign new_n2789 = ~new_n712 & new_n1369;
  assign new_n2790 = new_n2789 ^ new_n654;
  assign new_n2791 = ~new_n722 & new_n1373;
  assign new_n2792 = new_n2791 ^ new_n664;
  assign new_n2793 = ~new_n732 & new_n1377;
  assign new_n2794 = new_n2793 ^ new_n674;
  assign new_n2795 = ~new_n742 & new_n1381;
  assign new_n2796 = new_n2795 ^ new_n684;
  assign new_n2797 = ~new_n752 & new_n1385;
  assign new_n2798 = new_n2797 ^ new_n694;
  assign new_n2799 = ~new_n762 & new_n1389;
  assign new_n2800 = new_n2799 ^ new_n704;
  assign new_n2801 = ~new_n772 & new_n1393;
  assign new_n2802 = new_n2801 ^ new_n714;
  assign new_n2803 = ~new_n782 & new_n1397;
  assign new_n2804 = new_n2803 ^ new_n724;
  assign new_n2805 = ~new_n792 & new_n1401;
  assign new_n2806 = new_n2805 ^ new_n734;
  assign new_n2807 = ~new_n801 & new_n1405;
  assign new_n2808 = new_n2807 ^ new_n744;
  assign new_n2809 = ~new_n810 & new_n1153;
  assign new_n2810 = new_n2809 ^ new_n754;
  assign new_n2811 = ~new_n819 & new_n1157;
  assign new_n2812 = new_n2811 ^ new_n764;
  assign new_n2813 = ~new_n828 & new_n1161;
  assign new_n2814 = new_n2813 ^ new_n774;
  assign new_n2815 = ~new_n837 & new_n1165;
  assign new_n2816 = new_n2815 ^ new_n784;
  assign new_n2817 = new_n1641 ^ n489;
  assign new_n2818 = ~new_n1169 & new_n2817;
  assign new_n2819 = new_n2818 ^ new_n846;
  assign new_n2820 = new_n1645 ^ n490;
  assign new_n2821 = ~new_n1173 & new_n2820;
  assign new_n2822 = new_n2821 ^ new_n855;
  assign new_n2823 = new_n1649 ^ n491;
  assign new_n2824 = ~new_n1177 & new_n2823;
  assign new_n2825 = new_n2824 ^ new_n864;
  assign new_n2826 = new_n1653 ^ n492;
  assign new_n2827 = ~new_n1181 & new_n2826;
  assign new_n2828 = new_n2827 ^ new_n873;
  assign new_n2829 = new_n1657 ^ n493;
  assign new_n2830 = ~new_n1185 & new_n2829;
  assign new_n2831 = new_n2830 ^ new_n882;
  assign new_n2832 = new_n1661 ^ n494;
  assign new_n2833 = ~new_n1189 & new_n2832;
  assign new_n2834 = new_n2833 ^ new_n891;
  assign new_n2835 = new_n1409 ^ n495;
  assign new_n2836 = ~new_n1193 & new_n2835;
  assign new_n2837 = new_n2836 ^ new_n900;
  assign new_n2838 = new_n1413 ^ n496;
  assign new_n2839 = ~new_n1197 & new_n2838;
  assign new_n2840 = new_n2839 ^ new_n909;
  assign new_n2841 = new_n1417 ^ n497;
  assign new_n2842 = ~new_n1201 & new_n2841;
  assign new_n2843 = new_n2842 ^ new_n918;
  assign new_n2844 = new_n1421 ^ n498;
  assign new_n2845 = ~new_n1205 & new_n2844;
  assign new_n2846 = new_n2845 ^ new_n927;
  assign new_n2847 = new_n1425 ^ n499;
  assign new_n2848 = ~new_n1209 & new_n2847;
  assign new_n2849 = new_n2848 ^ new_n936;
  assign new_n2850 = new_n1429 ^ n500;
  assign new_n2851 = ~new_n1213 & new_n2850;
  assign new_n2852 = new_n2851 ^ new_n945;
  assign new_n2853 = new_n1433 ^ n501;
  assign new_n2854 = ~new_n1217 & new_n2853;
  assign new_n2855 = new_n2854 ^ new_n954;
  assign new_n2856 = new_n1437 ^ n502;
  assign new_n2857 = ~new_n1221 & new_n2856;
  assign new_n2858 = new_n2857 ^ new_n963;
  assign new_n2859 = new_n1441 ^ n503;
  assign new_n2860 = ~new_n1225 & new_n2859;
  assign new_n2861 = new_n2860 ^ new_n972;
  assign new_n2862 = new_n1445 ^ n504;
  assign new_n2863 = ~new_n1229 & new_n2862;
  assign new_n2864 = new_n2863 ^ new_n980;
  assign new_n2865 = new_n1449 ^ n505;
  assign new_n2866 = ~new_n1233 & new_n2865;
  assign new_n2867 = new_n2866 ^ new_n988;
  assign new_n2868 = new_n1453 ^ n506;
  assign new_n2869 = ~new_n1237 & new_n2868;
  assign new_n2870 = new_n2869 ^ new_n996;
  assign new_n2871 = new_n1457 ^ n507;
  assign new_n2872 = ~new_n1241 & new_n2871;
  assign new_n2873 = new_n2872 ^ new_n1004;
  assign new_n2874 = new_n1461 ^ n508;
  assign new_n2875 = ~new_n1245 & new_n2874;
  assign new_n2876 = new_n2875 ^ new_n1012;
  assign new_n2877 = new_n1465 ^ n509;
  assign new_n2878 = ~new_n1249 & new_n2877;
  assign new_n2879 = new_n2878 ^ new_n1020;
  assign new_n2880 = new_n1469 ^ n510;
  assign new_n2881 = ~new_n1253 & new_n2880;
  assign new_n2882 = new_n2881 ^ new_n1028;
  assign new_n2883 = new_n1473 ^ n511;
  assign new_n2884 = ~new_n1257 & new_n2883;
  assign new_n2885 = new_n2884 ^ new_n1036;
  assign new_n2886 = new_n1477 ^ n512;
  assign new_n2887 = ~new_n1261 & new_n2886;
  assign new_n2888 = new_n2887 ^ new_n1044;
  assign new_n2889 = new_n1481 ^ n513;
  assign new_n2890 = ~new_n1265 & new_n2889;
  assign new_n2891 = new_n2890 ^ new_n1052;
  assign new_n2892 = new_n1485 ^ n514;
  assign new_n2893 = ~new_n1269 & new_n2892;
  assign new_n2894 = new_n2893 ^ new_n1060;
  assign new_n2895 = new_n1489 ^ n515;
  assign new_n2896 = ~new_n1273 & new_n2895;
  assign new_n2897 = new_n2896 ^ new_n1068;
  assign new_n2898 = new_n1493 ^ n516;
  assign new_n2899 = ~new_n1277 & new_n2898;
  assign new_n2900 = new_n2899 ^ new_n1076;
  assign new_n2901 = new_n1497 ^ n517;
  assign new_n2902 = ~new_n1281 & new_n2901;
  assign new_n2903 = new_n2902 ^ new_n1084;
  assign new_n2904 = new_n1501 ^ n518;
  assign new_n2905 = ~new_n1285 & new_n2904;
  assign new_n2906 = new_n2905 ^ new_n1092;
  assign new_n2907 = new_n1505 ^ n519;
  assign new_n2908 = ~new_n1289 & new_n2907;
  assign new_n2909 = new_n2908 ^ new_n1100;
  assign new_n2910 = new_n1509 ^ n520;
  assign new_n2911 = ~new_n1293 & new_n2910;
  assign new_n2912 = new_n2911 ^ new_n1108;
  assign new_n2913 = new_n1513 ^ n521;
  assign new_n2914 = ~new_n1297 & new_n2913;
  assign new_n2915 = new_n2914 ^ new_n1116;
  assign new_n2916 = new_n1517 ^ n522;
  assign new_n2917 = ~new_n1301 & new_n2916;
  assign new_n2918 = new_n2917 ^ new_n1124;
  assign new_n2919 = new_n1521 ^ n523;
  assign new_n2920 = ~new_n1305 & new_n2919;
  assign new_n2921 = new_n2920 ^ new_n1132;
  assign new_n2922 = new_n1525 ^ n524;
  assign new_n2923 = ~new_n1309 & new_n2922;
  assign new_n2924 = new_n2923 ^ new_n1140;
  assign new_n2925 = new_n1529 ^ n525;
  assign new_n2926 = ~new_n1313 & new_n2925;
  assign new_n2927 = new_n2926 ^ new_n1148;
  assign new_n2928 = new_n1533 ^ n526;
  assign new_n2929 = ~new_n1317 & new_n2928;
  assign new_n2930 = new_n2929 ^ new_n582;
  assign new_n2931 = new_n1537 ^ n527;
  assign new_n2932 = ~new_n1321 & new_n2931;
  assign new_n2933 = new_n2932 ^ new_n592;
  assign new_n2934 = new_n1541 ^ n528;
  assign new_n2935 = ~new_n1325 & new_n2934;
  assign new_n2936 = new_n2935 ^ new_n602;
  assign new_n2937 = new_n1545 ^ n529;
  assign new_n2938 = ~new_n1329 & new_n2937;
  assign new_n2939 = new_n2938 ^ new_n612;
  assign new_n2940 = new_n1549 ^ n530;
  assign new_n2941 = ~new_n1333 & new_n2940;
  assign new_n2942 = new_n2941 ^ new_n622;
  assign new_n2943 = new_n1553 ^ n531;
  assign new_n2944 = ~new_n1337 & new_n2943;
  assign new_n2945 = new_n2944 ^ new_n632;
  assign new_n2946 = new_n1557 ^ n532;
  assign new_n2947 = ~new_n1341 & new_n2946;
  assign new_n2948 = new_n2947 ^ new_n642;
  assign new_n2949 = new_n1561 ^ n533;
  assign new_n2950 = ~new_n1345 & new_n2949;
  assign new_n2951 = new_n2950 ^ new_n652;
  assign new_n2952 = new_n1565 ^ n534;
  assign new_n2953 = ~new_n1349 & new_n2952;
  assign new_n2954 = new_n2953 ^ new_n662;
  assign new_n2955 = new_n1569 ^ n535;
  assign new_n2956 = ~new_n1353 & new_n2955;
  assign new_n2957 = new_n2956 ^ new_n672;
  assign new_n2958 = new_n1573 ^ n536;
  assign new_n2959 = ~new_n1357 & new_n2958;
  assign new_n2960 = new_n2959 ^ new_n682;
  assign new_n2961 = new_n1577 ^ n537;
  assign new_n2962 = ~new_n1361 & new_n2961;
  assign new_n2963 = new_n2962 ^ new_n692;
  assign new_n2964 = new_n1581 ^ n538;
  assign new_n2965 = ~new_n1365 & new_n2964;
  assign new_n2966 = new_n2965 ^ new_n702;
  assign new_n2967 = new_n1585 ^ n539;
  assign new_n2968 = ~new_n1369 & new_n2967;
  assign new_n2969 = new_n2968 ^ new_n712;
  assign new_n2970 = new_n1589 ^ n540;
  assign new_n2971 = ~new_n1373 & new_n2970;
  assign new_n2972 = new_n2971 ^ new_n722;
  assign new_n2973 = new_n1593 ^ n541;
  assign new_n2974 = ~new_n1377 & new_n2973;
  assign new_n2975 = new_n2974 ^ new_n732;
  assign new_n2976 = new_n1597 ^ n542;
  assign new_n2977 = ~new_n1381 & new_n2976;
  assign new_n2978 = new_n2977 ^ new_n742;
  assign new_n2979 = new_n1601 ^ n543;
  assign new_n2980 = ~new_n1385 & new_n2979;
  assign new_n2981 = new_n2980 ^ new_n752;
  assign new_n2982 = new_n1605 ^ n544;
  assign new_n2983 = ~new_n1389 & new_n2982;
  assign new_n2984 = new_n2983 ^ new_n762;
  assign new_n2985 = new_n1609 ^ n481;
  assign new_n2986 = ~new_n1393 & new_n2985;
  assign new_n2987 = new_n2986 ^ new_n772;
  assign new_n2988 = new_n1613 ^ n482;
  assign new_n2989 = ~new_n1397 & new_n2988;
  assign new_n2990 = new_n2989 ^ new_n782;
  assign new_n2991 = new_n1617 ^ n483;
  assign new_n2992 = ~new_n1401 & new_n2991;
  assign new_n2993 = new_n2992 ^ new_n792;
  assign new_n2994 = new_n1621 ^ n484;
  assign new_n2995 = ~new_n1405 & new_n2994;
  assign new_n2996 = new_n2995 ^ new_n801;
  assign new_n2997 = new_n1625 ^ n485;
  assign new_n2998 = ~new_n1153 & new_n2997;
  assign new_n2999 = new_n2998 ^ new_n810;
  assign new_n3000 = new_n1629 ^ n486;
  assign new_n3001 = ~new_n1157 & new_n3000;
  assign new_n3002 = new_n3001 ^ new_n819;
  assign new_n3003 = new_n1633 ^ n487;
  assign new_n3004 = ~new_n1161 & new_n3003;
  assign new_n3005 = new_n3004 ^ new_n828;
  assign new_n3006 = new_n1637 ^ n488;
  assign new_n3007 = ~new_n1165 & new_n3006;
  assign new_n3008 = new_n3007 ^ new_n837;
  assign new_n3009 = new_n759 ^ n563;
  assign new_n3010 = ~new_n2817 & new_n3009;
  assign new_n3011 = new_n3010 ^ new_n1169;
  assign new_n3012 = new_n769 ^ n564;
  assign new_n3013 = ~new_n2820 & new_n3012;
  assign new_n3014 = new_n3013 ^ new_n1173;
  assign new_n3015 = new_n779 ^ n565;
  assign new_n3016 = ~new_n2823 & new_n3015;
  assign new_n3017 = new_n3016 ^ new_n1177;
  assign new_n3018 = new_n789 ^ n566;
  assign new_n3019 = ~new_n2826 & new_n3018;
  assign new_n3020 = new_n3019 ^ new_n1181;
  assign new_n3021 = new_n799 ^ n567;
  assign new_n3022 = ~new_n2829 & new_n3021;
  assign new_n3023 = new_n3022 ^ new_n1185;
  assign new_n3024 = new_n808 ^ n568;
  assign new_n3025 = ~new_n2832 & new_n3024;
  assign new_n3026 = new_n3025 ^ new_n1189;
  assign new_n3027 = new_n817 ^ n569;
  assign new_n3028 = ~new_n2835 & new_n3027;
  assign new_n3029 = new_n3028 ^ new_n1193;
  assign new_n3030 = new_n826 ^ n570;
  assign new_n3031 = ~new_n2838 & new_n3030;
  assign new_n3032 = new_n3031 ^ new_n1197;
  assign new_n3033 = new_n835 ^ n571;
  assign new_n3034 = ~new_n2841 & new_n3033;
  assign new_n3035 = new_n3034 ^ new_n1201;
  assign new_n3036 = new_n844 ^ n572;
  assign new_n3037 = ~new_n2844 & new_n3036;
  assign new_n3038 = new_n3037 ^ new_n1205;
  assign new_n3039 = new_n853 ^ n573;
  assign new_n3040 = ~new_n2847 & new_n3039;
  assign new_n3041 = new_n3040 ^ new_n1209;
  assign new_n3042 = new_n862 ^ n574;
  assign new_n3043 = ~new_n2850 & new_n3042;
  assign new_n3044 = new_n3043 ^ new_n1213;
  assign new_n3045 = new_n871 ^ n575;
  assign new_n3046 = ~new_n2853 & new_n3045;
  assign new_n3047 = new_n3046 ^ new_n1217;
  assign new_n3048 = new_n880 ^ n576;
  assign new_n3049 = ~new_n2856 & new_n3048;
  assign new_n3050 = new_n3049 ^ new_n1221;
  assign new_n3051 = new_n889 ^ n1;
  assign new_n3052 = ~new_n2859 & new_n3051;
  assign new_n3053 = new_n3052 ^ new_n1225;
  assign new_n3054 = new_n898 ^ n2;
  assign new_n3055 = ~new_n2862 & new_n3054;
  assign new_n3056 = new_n3055 ^ new_n1229;
  assign new_n3057 = new_n907 ^ n3;
  assign new_n3058 = ~new_n2865 & new_n3057;
  assign new_n3059 = new_n3058 ^ new_n1233;
  assign new_n3060 = new_n916 ^ n4;
  assign new_n3061 = ~new_n2868 & new_n3060;
  assign new_n3062 = new_n3061 ^ new_n1237;
  assign new_n3063 = new_n925 ^ n5;
  assign new_n3064 = ~new_n2871 & new_n3063;
  assign new_n3065 = new_n3064 ^ new_n1241;
  assign new_n3066 = new_n934 ^ n6;
  assign new_n3067 = ~new_n2874 & new_n3066;
  assign new_n3068 = new_n3067 ^ new_n1245;
  assign new_n3069 = new_n943 ^ n7;
  assign new_n3070 = ~new_n2877 & new_n3069;
  assign new_n3071 = new_n3070 ^ new_n1249;
  assign new_n3072 = new_n952 ^ n8;
  assign new_n3073 = ~new_n2880 & new_n3072;
  assign new_n3074 = new_n3073 ^ new_n1253;
  assign new_n3075 = new_n961 ^ n9;
  assign new_n3076 = ~new_n2883 & new_n3075;
  assign new_n3077 = new_n3076 ^ new_n1257;
  assign new_n3078 = new_n970 ^ n10;
  assign new_n3079 = ~new_n2886 & new_n3078;
  assign new_n3080 = new_n3079 ^ new_n1261;
  assign new_n3081 = new_n978 ^ n11;
  assign new_n3082 = ~new_n2889 & new_n3081;
  assign new_n3083 = new_n3082 ^ new_n1265;
  assign new_n3084 = new_n986 ^ n12;
  assign new_n3085 = ~new_n2892 & new_n3084;
  assign new_n3086 = new_n3085 ^ new_n1269;
  assign new_n3087 = new_n994 ^ n13;
  assign new_n3088 = ~new_n2895 & new_n3087;
  assign new_n3089 = new_n3088 ^ new_n1273;
  assign new_n3090 = new_n1002 ^ n14;
  assign new_n3091 = ~new_n2898 & new_n3090;
  assign new_n3092 = new_n3091 ^ new_n1277;
  assign new_n3093 = new_n1010 ^ n15;
  assign new_n3094 = ~new_n2901 & new_n3093;
  assign new_n3095 = new_n3094 ^ new_n1281;
  assign new_n3096 = new_n1018 ^ n16;
  assign new_n3097 = ~new_n2904 & new_n3096;
  assign new_n3098 = new_n3097 ^ new_n1285;
  assign new_n3099 = new_n1026 ^ n17;
  assign new_n3100 = ~new_n2907 & new_n3099;
  assign new_n3101 = new_n3100 ^ new_n1289;
  assign new_n3102 = new_n1034 ^ n18;
  assign new_n3103 = ~new_n2910 & new_n3102;
  assign new_n3104 = new_n3103 ^ new_n1293;
  assign new_n3105 = new_n1042 ^ n19;
  assign new_n3106 = ~new_n2913 & new_n3105;
  assign new_n3107 = new_n3106 ^ new_n1297;
  assign new_n3108 = new_n1050 ^ n20;
  assign new_n3109 = ~new_n2916 & new_n3108;
  assign new_n3110 = new_n3109 ^ new_n1301;
  assign new_n3111 = new_n1058 ^ n21;
  assign new_n3112 = ~new_n2919 & new_n3111;
  assign new_n3113 = new_n3112 ^ new_n1305;
  assign new_n3114 = new_n1066 ^ n22;
  assign new_n3115 = ~new_n2922 & new_n3114;
  assign new_n3116 = new_n3115 ^ new_n1309;
  assign new_n3117 = new_n1074 ^ n23;
  assign new_n3118 = ~new_n2925 & new_n3117;
  assign new_n3119 = new_n3118 ^ new_n1313;
  assign new_n3120 = new_n1082 ^ n24;
  assign new_n3121 = ~new_n2928 & new_n3120;
  assign new_n3122 = new_n3121 ^ new_n1317;
  assign new_n3123 = new_n1090 ^ n25;
  assign new_n3124 = ~new_n2931 & new_n3123;
  assign new_n3125 = new_n3124 ^ new_n1321;
  assign new_n3126 = new_n1098 ^ n26;
  assign new_n3127 = ~new_n2934 & new_n3126;
  assign new_n3128 = new_n3127 ^ new_n1325;
  assign new_n3129 = new_n1106 ^ n27;
  assign new_n3130 = ~new_n2937 & new_n3129;
  assign new_n3131 = new_n3130 ^ new_n1329;
  assign new_n3132 = new_n1114 ^ n28;
  assign new_n3133 = ~new_n2940 & new_n3132;
  assign new_n3134 = new_n3133 ^ new_n1333;
  assign new_n3135 = new_n1122 ^ n29;
  assign new_n3136 = ~new_n2943 & new_n3135;
  assign new_n3137 = new_n3136 ^ new_n1337;
  assign new_n3138 = new_n1130 ^ n30;
  assign new_n3139 = ~new_n2946 & new_n3138;
  assign new_n3140 = new_n3139 ^ new_n1341;
  assign new_n3141 = new_n1138 ^ n31;
  assign new_n3142 = ~new_n2949 & new_n3141;
  assign new_n3143 = new_n3142 ^ new_n1345;
  assign new_n3144 = new_n1146 ^ n32;
  assign new_n3145 = ~new_n2952 & new_n3144;
  assign new_n3146 = new_n3145 ^ new_n1349;
  assign new_n3147 = new_n579 ^ n545;
  assign new_n3148 = ~new_n2955 & new_n3147;
  assign new_n3149 = new_n3148 ^ new_n1353;
  assign new_n3150 = new_n589 ^ n546;
  assign new_n3151 = ~new_n2958 & new_n3150;
  assign new_n3152 = new_n3151 ^ new_n1357;
  assign new_n3153 = new_n599 ^ n547;
  assign new_n3154 = ~new_n2961 & new_n3153;
  assign new_n3155 = new_n3154 ^ new_n1361;
  assign new_n3156 = new_n609 ^ n548;
  assign new_n3157 = ~new_n2964 & new_n3156;
  assign new_n3158 = new_n3157 ^ new_n1365;
  assign new_n3159 = new_n619 ^ n549;
  assign new_n3160 = ~new_n2967 & new_n3159;
  assign new_n3161 = new_n3160 ^ new_n1369;
  assign new_n3162 = new_n629 ^ n550;
  assign new_n3163 = ~new_n2970 & new_n3162;
  assign new_n3164 = new_n3163 ^ new_n1373;
  assign new_n3165 = new_n639 ^ n551;
  assign new_n3166 = ~new_n2973 & new_n3165;
  assign new_n3167 = new_n3166 ^ new_n1377;
  assign new_n3168 = new_n649 ^ n552;
  assign new_n3169 = ~new_n2976 & new_n3168;
  assign new_n3170 = new_n3169 ^ new_n1381;
  assign new_n3171 = new_n659 ^ n553;
  assign new_n3172 = ~new_n2979 & new_n3171;
  assign new_n3173 = new_n3172 ^ new_n1385;
  assign new_n3174 = new_n669 ^ n554;
  assign new_n3175 = ~new_n2982 & new_n3174;
  assign new_n3176 = new_n3175 ^ new_n1389;
  assign new_n3177 = new_n679 ^ n555;
  assign new_n3178 = ~new_n2985 & new_n3177;
  assign new_n3179 = new_n3178 ^ new_n1393;
  assign new_n3180 = new_n689 ^ n556;
  assign new_n3181 = ~new_n2988 & new_n3180;
  assign new_n3182 = new_n3181 ^ new_n1397;
  assign new_n3183 = new_n699 ^ n557;
  assign new_n3184 = ~new_n2991 & new_n3183;
  assign new_n3185 = new_n3184 ^ new_n1401;
  assign new_n3186 = new_n709 ^ n558;
  assign new_n3187 = ~new_n2994 & new_n3186;
  assign new_n3188 = new_n3187 ^ new_n1405;
  assign new_n3189 = new_n719 ^ n559;
  assign new_n3190 = ~new_n2997 & new_n3189;
  assign new_n3191 = new_n3190 ^ new_n1153;
  assign new_n3192 = new_n729 ^ n560;
  assign new_n3193 = ~new_n3000 & new_n3192;
  assign new_n3194 = new_n3193 ^ new_n1157;
  assign new_n3195 = new_n739 ^ n561;
  assign new_n3196 = ~new_n3003 & new_n3195;
  assign new_n3197 = new_n3196 ^ new_n1161;
  assign new_n3198 = new_n749 ^ n562;
  assign new_n3199 = ~new_n3006 & new_n3198;
  assign new_n3200 = new_n3199 ^ new_n1165;
  assign new_n3201 = ~new_n3009 & new_n794;
  assign new_n3202 = new_n3201 ^ new_n2817;
  assign new_n3203 = ~new_n3012 & new_n803;
  assign new_n3204 = new_n3203 ^ new_n2820;
  assign new_n3205 = ~new_n3015 & new_n812;
  assign new_n3206 = new_n3205 ^ new_n2823;
  assign new_n3207 = ~new_n3018 & new_n821;
  assign new_n3208 = new_n3207 ^ new_n2826;
  assign new_n3209 = ~new_n3021 & new_n830;
  assign new_n3210 = new_n3209 ^ new_n2829;
  assign new_n3211 = ~new_n3024 & new_n839;
  assign new_n3212 = new_n3211 ^ new_n2832;
  assign new_n3213 = ~new_n3027 & new_n848;
  assign new_n3214 = new_n3213 ^ new_n2835;
  assign new_n3215 = ~new_n3030 & new_n857;
  assign new_n3216 = new_n3215 ^ new_n2838;
  assign new_n3217 = ~new_n3033 & new_n866;
  assign new_n3218 = new_n3217 ^ new_n2841;
  assign new_n3219 = ~new_n3036 & new_n875;
  assign new_n3220 = new_n3219 ^ new_n2844;
  assign new_n3221 = ~new_n3039 & new_n884;
  assign new_n3222 = new_n3221 ^ new_n2847;
  assign new_n3223 = ~new_n3042 & new_n893;
  assign new_n3224 = new_n3223 ^ new_n2850;
  assign new_n3225 = ~new_n3045 & new_n902;
  assign new_n3226 = new_n3225 ^ new_n2853;
  assign new_n3227 = ~new_n3048 & new_n911;
  assign new_n3228 = new_n3227 ^ new_n2856;
  assign new_n3229 = ~new_n3051 & new_n920;
  assign new_n3230 = new_n3229 ^ new_n2859;
  assign new_n3231 = ~new_n3054 & new_n929;
  assign new_n3232 = new_n3231 ^ new_n2862;
  assign new_n3233 = ~new_n3057 & new_n938;
  assign new_n3234 = new_n3233 ^ new_n2865;
  assign new_n3235 = ~new_n3060 & new_n947;
  assign new_n3236 = new_n3235 ^ new_n2868;
  assign new_n3237 = ~new_n3063 & new_n956;
  assign new_n3238 = new_n3237 ^ new_n2871;
  assign new_n3239 = ~new_n3066 & new_n965;
  assign new_n3240 = new_n3239 ^ new_n2874;
  assign new_n3241 = ~new_n3069 & new_n974;
  assign new_n3242 = new_n3241 ^ new_n2877;
  assign new_n3243 = ~new_n3072 & new_n982;
  assign new_n3244 = new_n3243 ^ new_n2880;
  assign new_n3245 = ~new_n3075 & new_n990;
  assign new_n3246 = new_n3245 ^ new_n2883;
  assign new_n3247 = ~new_n3078 & new_n998;
  assign new_n3248 = new_n3247 ^ new_n2886;
  assign new_n3249 = ~new_n3081 & new_n1006;
  assign new_n3250 = new_n3249 ^ new_n2889;
  assign new_n3251 = ~new_n3084 & new_n1014;
  assign new_n3252 = new_n3251 ^ new_n2892;
  assign new_n3253 = ~new_n3087 & new_n1022;
  assign new_n3254 = new_n3253 ^ new_n2895;
  assign new_n3255 = ~new_n3090 & new_n1030;
  assign new_n3256 = new_n3255 ^ new_n2898;
  assign new_n3257 = ~new_n3093 & new_n1038;
  assign new_n3258 = new_n3257 ^ new_n2901;
  assign new_n3259 = ~new_n3096 & new_n1046;
  assign new_n3260 = new_n3259 ^ new_n2904;
  assign new_n3261 = ~new_n3099 & new_n1054;
  assign new_n3262 = new_n3261 ^ new_n2907;
  assign new_n3263 = ~new_n3102 & new_n1062;
  assign new_n3264 = new_n3263 ^ new_n2910;
  assign new_n3265 = ~new_n3105 & new_n1070;
  assign new_n3266 = new_n3265 ^ new_n2913;
  assign new_n3267 = ~new_n3108 & new_n1078;
  assign new_n3268 = new_n3267 ^ new_n2916;
  assign new_n3269 = ~new_n3111 & new_n1086;
  assign new_n3270 = new_n3269 ^ new_n2919;
  assign new_n3271 = ~new_n3114 & new_n1094;
  assign new_n3272 = new_n3271 ^ new_n2922;
  assign new_n3273 = ~new_n3117 & new_n1102;
  assign new_n3274 = new_n3273 ^ new_n2925;
  assign new_n3275 = ~new_n3120 & new_n1110;
  assign new_n3276 = new_n3275 ^ new_n2928;
  assign new_n3277 = ~new_n3123 & new_n1118;
  assign new_n3278 = new_n3277 ^ new_n2931;
  assign new_n3279 = ~new_n3126 & new_n1126;
  assign new_n3280 = new_n3279 ^ new_n2934;
  assign new_n3281 = ~new_n3129 & new_n1134;
  assign new_n3282 = new_n3281 ^ new_n2937;
  assign new_n3283 = ~new_n3132 & new_n1142;
  assign new_n3284 = new_n3283 ^ new_n2940;
  assign new_n3285 = ~new_n3135 & new_n1150;
  assign new_n3286 = new_n3285 ^ new_n2943;
  assign new_n3287 = ~new_n3138 & new_n584;
  assign new_n3288 = new_n3287 ^ new_n2946;
  assign new_n3289 = ~new_n3141 & new_n594;
  assign new_n3290 = new_n3289 ^ new_n2949;
  assign new_n3291 = ~new_n3144 & new_n604;
  assign new_n3292 = new_n3291 ^ new_n2952;
  assign new_n3293 = ~new_n3147 & new_n614;
  assign new_n3294 = new_n3293 ^ new_n2955;
  assign new_n3295 = ~new_n3150 & new_n624;
  assign new_n3296 = new_n3295 ^ new_n2958;
  assign new_n3297 = ~new_n3153 & new_n634;
  assign new_n3298 = new_n3297 ^ new_n2961;
  assign new_n3299 = ~new_n3156 & new_n644;
  assign new_n3300 = new_n3299 ^ new_n2964;
  assign new_n3301 = ~new_n3159 & new_n654;
  assign new_n3302 = new_n3301 ^ new_n2967;
  assign new_n3303 = ~new_n3162 & new_n664;
  assign new_n3304 = new_n3303 ^ new_n2970;
  assign new_n3305 = ~new_n3165 & new_n674;
  assign new_n3306 = new_n3305 ^ new_n2973;
  assign new_n3307 = ~new_n3168 & new_n684;
  assign new_n3308 = new_n3307 ^ new_n2976;
  assign new_n3309 = ~new_n3171 & new_n694;
  assign new_n3310 = new_n3309 ^ new_n2979;
  assign new_n3311 = ~new_n3174 & new_n704;
  assign new_n3312 = new_n3311 ^ new_n2982;
  assign new_n3313 = ~new_n3177 & new_n714;
  assign new_n3314 = new_n3313 ^ new_n2985;
  assign new_n3315 = ~new_n3180 & new_n724;
  assign new_n3316 = new_n3315 ^ new_n2988;
  assign new_n3317 = ~new_n3183 & new_n734;
  assign new_n3318 = new_n3317 ^ new_n2991;
  assign new_n3319 = ~new_n3186 & new_n744;
  assign new_n3320 = new_n3319 ^ new_n2994;
  assign new_n3321 = ~new_n3189 & new_n754;
  assign new_n3322 = new_n3321 ^ new_n2997;
  assign new_n3323 = ~new_n3192 & new_n764;
  assign new_n3324 = new_n3323 ^ new_n3000;
  assign new_n3325 = ~new_n3195 & new_n774;
  assign new_n3326 = new_n3325 ^ new_n3003;
  assign new_n3327 = ~new_n3198 & new_n784;
  assign new_n3328 = new_n3327 ^ new_n3006;
  assign new_n3329 = ~new_n794 & new_n846;
  assign new_n3330 = new_n3329 ^ new_n3009;
  assign new_n3331 = ~new_n803 & new_n855;
  assign new_n3332 = new_n3331 ^ new_n3012;
  assign new_n3333 = ~new_n812 & new_n864;
  assign new_n3334 = new_n3333 ^ new_n3015;
  assign new_n3335 = ~new_n821 & new_n873;
  assign new_n3336 = new_n3335 ^ new_n3018;
  assign new_n3337 = ~new_n830 & new_n882;
  assign new_n3338 = new_n3337 ^ new_n3021;
  assign new_n3339 = ~new_n839 & new_n891;
  assign new_n3340 = new_n3339 ^ new_n3024;
  assign new_n3341 = ~new_n848 & new_n900;
  assign new_n3342 = new_n3341 ^ new_n3027;
  assign new_n3343 = ~new_n857 & new_n909;
  assign new_n3344 = new_n3343 ^ new_n3030;
  assign new_n3345 = ~new_n866 & new_n918;
  assign new_n3346 = new_n3345 ^ new_n3033;
  assign new_n3347 = ~new_n875 & new_n927;
  assign new_n3348 = new_n3347 ^ new_n3036;
  assign new_n3349 = ~new_n884 & new_n936;
  assign new_n3350 = new_n3349 ^ new_n3039;
  assign new_n3351 = ~new_n893 & new_n945;
  assign new_n3352 = new_n3351 ^ new_n3042;
  assign new_n3353 = ~new_n902 & new_n954;
  assign new_n3354 = new_n3353 ^ new_n3045;
  assign new_n3355 = ~new_n911 & new_n963;
  assign new_n3356 = new_n3355 ^ new_n3048;
  assign new_n3357 = ~new_n920 & new_n972;
  assign new_n3358 = new_n3357 ^ new_n3051;
  assign new_n3359 = ~new_n929 & new_n980;
  assign new_n3360 = new_n3359 ^ new_n3054;
  assign new_n3361 = ~new_n938 & new_n988;
  assign new_n3362 = new_n3361 ^ new_n3057;
  assign new_n3363 = ~new_n947 & new_n996;
  assign new_n3364 = new_n3363 ^ new_n3060;
  assign new_n3365 = ~new_n956 & new_n1004;
  assign new_n3366 = new_n3365 ^ new_n3063;
  assign new_n3367 = ~new_n965 & new_n1012;
  assign new_n3368 = new_n3367 ^ new_n3066;
  assign new_n3369 = ~new_n974 & new_n1020;
  assign new_n3370 = new_n3369 ^ new_n3069;
  assign new_n3371 = ~new_n982 & new_n1028;
  assign new_n3372 = new_n3371 ^ new_n3072;
  assign new_n3373 = ~new_n990 & new_n1036;
  assign new_n3374 = new_n3373 ^ new_n3075;
  assign new_n3375 = ~new_n998 & new_n1044;
  assign new_n3376 = new_n3375 ^ new_n3078;
  assign new_n3377 = ~new_n1006 & new_n1052;
  assign new_n3378 = new_n3377 ^ new_n3081;
  assign new_n3379 = ~new_n1014 & new_n1060;
  assign new_n3380 = new_n3379 ^ new_n3084;
  assign new_n3381 = ~new_n1022 & new_n1068;
  assign new_n3382 = new_n3381 ^ new_n3087;
  assign new_n3383 = ~new_n1030 & new_n1076;
  assign new_n3384 = new_n3383 ^ new_n3090;
  assign new_n3385 = ~new_n1038 & new_n1084;
  assign new_n3386 = new_n3385 ^ new_n3093;
  assign new_n3387 = ~new_n1046 & new_n1092;
  assign new_n3388 = new_n3387 ^ new_n3096;
  assign new_n3389 = ~new_n1054 & new_n1100;
  assign new_n3390 = new_n3389 ^ new_n3099;
  assign new_n3391 = ~new_n1062 & new_n1108;
  assign new_n3392 = new_n3391 ^ new_n3102;
  assign new_n3393 = ~new_n1070 & new_n1116;
  assign new_n3394 = new_n3393 ^ new_n3105;
  assign new_n3395 = ~new_n1078 & new_n1124;
  assign new_n3396 = new_n3395 ^ new_n3108;
  assign new_n3397 = ~new_n1086 & new_n1132;
  assign new_n3398 = new_n3397 ^ new_n3111;
  assign new_n3399 = ~new_n1094 & new_n1140;
  assign new_n3400 = new_n3399 ^ new_n3114;
  assign new_n3401 = ~new_n1102 & new_n1148;
  assign new_n3402 = new_n3401 ^ new_n3117;
  assign new_n3403 = ~new_n1110 & new_n582;
  assign new_n3404 = new_n3403 ^ new_n3120;
  assign new_n3405 = ~new_n1118 & new_n592;
  assign new_n3406 = new_n3405 ^ new_n3123;
  assign new_n3407 = ~new_n1126 & new_n602;
  assign new_n3408 = new_n3407 ^ new_n3126;
  assign new_n3409 = ~new_n1134 & new_n612;
  assign new_n3410 = new_n3409 ^ new_n3129;
  assign new_n3411 = ~new_n1142 & new_n622;
  assign new_n3412 = new_n3411 ^ new_n3132;
  assign new_n3413 = ~new_n1150 & new_n632;
  assign new_n3414 = new_n3413 ^ new_n3135;
  assign new_n3415 = ~new_n584 & new_n642;
  assign new_n3416 = new_n3415 ^ new_n3138;
  assign new_n3417 = ~new_n594 & new_n652;
  assign new_n3418 = new_n3417 ^ new_n3141;
  assign new_n3419 = ~new_n604 & new_n662;
  assign new_n3420 = new_n3419 ^ new_n3144;
  assign new_n3421 = ~new_n614 & new_n672;
  assign new_n3422 = new_n3421 ^ new_n3147;
  assign new_n3423 = ~new_n624 & new_n682;
  assign new_n3424 = new_n3423 ^ new_n3150;
  assign new_n3425 = ~new_n634 & new_n692;
  assign new_n3426 = new_n3425 ^ new_n3153;
  assign new_n3427 = ~new_n644 & new_n702;
  assign new_n3428 = new_n3427 ^ new_n3156;
  assign new_n3429 = ~new_n654 & new_n712;
  assign new_n3430 = new_n3429 ^ new_n3159;
  assign new_n3431 = ~new_n664 & new_n722;
  assign new_n3432 = new_n3431 ^ new_n3162;
  assign new_n3433 = ~new_n674 & new_n732;
  assign new_n3434 = new_n3433 ^ new_n3165;
  assign new_n3435 = ~new_n684 & new_n742;
  assign new_n3436 = new_n3435 ^ new_n3168;
  assign new_n3437 = ~new_n694 & new_n752;
  assign new_n3438 = new_n3437 ^ new_n3171;
  assign new_n3439 = ~new_n704 & new_n762;
  assign new_n3440 = new_n3439 ^ new_n3174;
  assign new_n3441 = ~new_n714 & new_n772;
  assign new_n3442 = new_n3441 ^ new_n3177;
  assign new_n3443 = ~new_n724 & new_n782;
  assign new_n3444 = new_n3443 ^ new_n3180;
  assign new_n3445 = ~new_n734 & new_n792;
  assign new_n3446 = new_n3445 ^ new_n3183;
  assign new_n3447 = ~new_n744 & new_n801;
  assign new_n3448 = new_n3447 ^ new_n3186;
  assign new_n3449 = ~new_n754 & new_n810;
  assign new_n3450 = new_n3449 ^ new_n3189;
  assign new_n3451 = ~new_n764 & new_n819;
  assign new_n3452 = new_n3451 ^ new_n3192;
  assign new_n3453 = ~new_n774 & new_n828;
  assign new_n3454 = new_n3453 ^ new_n3195;
  assign new_n3455 = ~new_n784 & new_n837;
  assign new_n3456 = new_n3455 ^ new_n3198;
  assign new_n3457 = ~new_n925 & new_n875;
  assign new_n3458 = new_n3457 ^ new_n1461;
  assign new_n3459 = ~new_n934 & new_n884;
  assign new_n3460 = new_n3459 ^ new_n1465;
  assign new_n3461 = ~new_n943 & new_n893;
  assign new_n3462 = new_n3461 ^ new_n1469;
  assign new_n3463 = ~new_n952 & new_n902;
  assign new_n3464 = new_n3463 ^ new_n1473;
  assign new_n3465 = ~new_n961 & new_n911;
  assign new_n3466 = new_n3465 ^ new_n1477;
  assign new_n3467 = ~new_n970 & new_n920;
  assign new_n3468 = new_n3467 ^ new_n1481;
  assign new_n3469 = ~new_n978 & new_n929;
  assign new_n3470 = new_n3469 ^ new_n1485;
  assign new_n3471 = ~new_n986 & new_n938;
  assign new_n3472 = new_n3471 ^ new_n1489;
  assign new_n3473 = ~new_n994 & new_n947;
  assign new_n3474 = new_n3473 ^ new_n1493;
  assign new_n3475 = ~new_n1002 & new_n956;
  assign new_n3476 = new_n3475 ^ new_n1497;
  assign new_n3477 = ~new_n1010 & new_n965;
  assign new_n3478 = new_n3477 ^ new_n1501;
  assign new_n3479 = ~new_n1018 & new_n974;
  assign new_n3480 = new_n3479 ^ new_n1505;
  assign new_n3481 = ~new_n1026 & new_n982;
  assign new_n3482 = new_n3481 ^ new_n1509;
  assign new_n3483 = ~new_n1034 & new_n990;
  assign new_n3484 = new_n3483 ^ new_n1513;
  assign new_n3485 = ~new_n1042 & new_n998;
  assign new_n3486 = new_n3485 ^ new_n1517;
  assign new_n3487 = ~new_n1050 & new_n1006;
  assign new_n3488 = new_n3487 ^ new_n1521;
  assign new_n3489 = ~new_n1058 & new_n1014;
  assign new_n3490 = new_n3489 ^ new_n1525;
  assign new_n3491 = ~new_n1066 & new_n1022;
  assign new_n3492 = new_n3491 ^ new_n1529;
  assign new_n3493 = ~new_n1074 & new_n1030;
  assign new_n3494 = new_n3493 ^ new_n1533;
  assign new_n3495 = ~new_n1082 & new_n1038;
  assign new_n3496 = new_n3495 ^ new_n1537;
  assign new_n3497 = ~new_n1090 & new_n1046;
  assign new_n3498 = new_n3497 ^ new_n1541;
  assign new_n3499 = ~new_n1098 & new_n1054;
  assign new_n3500 = new_n3499 ^ new_n1545;
  assign new_n3501 = ~new_n1106 & new_n1062;
  assign new_n3502 = new_n3501 ^ new_n1549;
  assign new_n3503 = ~new_n1114 & new_n1070;
  assign new_n3504 = new_n3503 ^ new_n1553;
  assign new_n3505 = ~new_n1122 & new_n1078;
  assign new_n3506 = new_n3505 ^ new_n1557;
  assign new_n3507 = ~new_n1130 & new_n1086;
  assign new_n3508 = new_n3507 ^ new_n1561;
  assign new_n3509 = ~new_n1138 & new_n1094;
  assign new_n3510 = new_n3509 ^ new_n1565;
  assign new_n3511 = ~new_n1146 & new_n1102;
  assign new_n3512 = new_n3511 ^ new_n1569;
  assign new_n3513 = ~new_n579 & new_n1110;
  assign new_n3514 = new_n3513 ^ new_n1573;
  assign new_n3515 = ~new_n589 & new_n1118;
  assign new_n3516 = new_n3515 ^ new_n1577;
  assign new_n3517 = ~new_n599 & new_n1126;
  assign new_n3518 = new_n3517 ^ new_n1581;
  assign new_n3519 = ~new_n609 & new_n1134;
  assign new_n3520 = new_n3519 ^ new_n1585;
  assign new_n3521 = ~new_n619 & new_n1142;
  assign new_n3522 = new_n3521 ^ new_n1589;
  assign new_n3523 = ~new_n629 & new_n1150;
  assign new_n3524 = new_n3523 ^ new_n1593;
  assign new_n3525 = ~new_n639 & new_n584;
  assign new_n3526 = new_n3525 ^ new_n1597;
  assign new_n3527 = ~new_n649 & new_n594;
  assign new_n3528 = new_n3527 ^ new_n1601;
  assign new_n3529 = ~new_n659 & new_n604;
  assign new_n3530 = new_n3529 ^ new_n1605;
  assign new_n3531 = ~new_n669 & new_n614;
  assign new_n3532 = new_n3531 ^ new_n1609;
  assign new_n3533 = ~new_n679 & new_n624;
  assign new_n3534 = new_n3533 ^ new_n1613;
  assign new_n3535 = ~new_n689 & new_n634;
  assign new_n3536 = new_n3535 ^ new_n1617;
  assign new_n3537 = ~new_n699 & new_n644;
  assign new_n3538 = new_n3537 ^ new_n1621;
  assign new_n3539 = ~new_n709 & new_n654;
  assign new_n3540 = new_n3539 ^ new_n1625;
  assign new_n3541 = ~new_n719 & new_n664;
  assign new_n3542 = new_n3541 ^ new_n1629;
  assign new_n3543 = ~new_n729 & new_n674;
  assign new_n3544 = new_n3543 ^ new_n1633;
  assign new_n3545 = ~new_n739 & new_n684;
  assign new_n3546 = new_n3545 ^ new_n1637;
  assign new_n3547 = ~new_n749 & new_n694;
  assign new_n3548 = new_n3547 ^ new_n1641;
  assign new_n3549 = ~new_n759 & new_n704;
  assign new_n3550 = new_n3549 ^ new_n1645;
  assign new_n3551 = ~new_n769 & new_n714;
  assign new_n3552 = new_n3551 ^ new_n1649;
  assign new_n3553 = ~new_n779 & new_n724;
  assign new_n3554 = new_n3553 ^ new_n1653;
  assign new_n3555 = ~new_n789 & new_n734;
  assign new_n3556 = new_n3555 ^ new_n1657;
  assign new_n3557 = ~new_n799 & new_n744;
  assign new_n3558 = new_n3557 ^ new_n1661;
  assign new_n3559 = ~new_n808 & new_n754;
  assign new_n3560 = new_n3559 ^ new_n1409;
  assign new_n3561 = ~new_n817 & new_n764;
  assign new_n3562 = new_n3561 ^ new_n1413;
  assign new_n3563 = ~new_n826 & new_n774;
  assign new_n3564 = new_n3563 ^ new_n1417;
  assign new_n3565 = ~new_n835 & new_n784;
  assign new_n3566 = new_n3565 ^ new_n1421;
  assign new_n3567 = ~new_n844 & new_n794;
  assign new_n3568 = new_n3567 ^ new_n1425;
  assign new_n3569 = ~new_n853 & new_n803;
  assign new_n3570 = new_n3569 ^ new_n1429;
  assign new_n3571 = ~new_n862 & new_n812;
  assign new_n3572 = new_n3571 ^ new_n1433;
  assign new_n3573 = ~new_n871 & new_n821;
  assign new_n3574 = new_n3573 ^ new_n1437;
  assign new_n3575 = ~new_n880 & new_n830;
  assign new_n3576 = new_n3575 ^ new_n1441;
  assign new_n3577 = ~new_n889 & new_n839;
  assign new_n3578 = new_n3577 ^ new_n1445;
  assign new_n3579 = ~new_n898 & new_n848;
  assign new_n3580 = new_n3579 ^ new_n1449;
  assign new_n3581 = ~new_n907 & new_n857;
  assign new_n3582 = new_n3581 ^ new_n1453;
  assign new_n3583 = ~new_n916 & new_n866;
  assign new_n3584 = new_n3583 ^ new_n1457;
  assign new_n3585 = new_n927 ^ n368;
  assign new_n3586 = ~new_n875 & new_n3585;
  assign new_n3587 = new_n3586 ^ new_n925;
  assign new_n3588 = new_n936 ^ n369;
  assign new_n3589 = ~new_n884 & new_n3588;
  assign new_n3590 = new_n3589 ^ new_n934;
  assign new_n3591 = new_n945 ^ n370;
  assign new_n3592 = ~new_n893 & new_n3591;
  assign new_n3593 = new_n3592 ^ new_n943;
  assign new_n3594 = new_n954 ^ n371;
  assign new_n3595 = ~new_n902 & new_n3594;
  assign new_n3596 = new_n3595 ^ new_n952;
  assign new_n3597 = new_n963 ^ n372;
  assign new_n3598 = ~new_n911 & new_n3597;
  assign new_n3599 = new_n3598 ^ new_n961;
  assign new_n3600 = new_n972 ^ n373;
  assign new_n3601 = ~new_n920 & new_n3600;
  assign new_n3602 = new_n3601 ^ new_n970;
  assign new_n3603 = new_n980 ^ n374;
  assign new_n3604 = ~new_n929 & new_n3603;
  assign new_n3605 = new_n3604 ^ new_n978;
  assign new_n3606 = new_n988 ^ n375;
  assign new_n3607 = ~new_n938 & new_n3606;
  assign new_n3608 = new_n3607 ^ new_n986;
  assign new_n3609 = new_n996 ^ n376;
  assign new_n3610 = ~new_n947 & new_n3609;
  assign new_n3611 = new_n3610 ^ new_n994;
  assign new_n3612 = new_n1004 ^ n377;
  assign new_n3613 = ~new_n956 & new_n3612;
  assign new_n3614 = new_n3613 ^ new_n1002;
  assign new_n3615 = new_n1012 ^ n378;
  assign new_n3616 = ~new_n965 & new_n3615;
  assign new_n3617 = new_n3616 ^ new_n1010;
  assign new_n3618 = new_n1020 ^ n379;
  assign new_n3619 = ~new_n974 & new_n3618;
  assign new_n3620 = new_n3619 ^ new_n1018;
  assign new_n3621 = new_n1028 ^ n380;
  assign new_n3622 = ~new_n982 & new_n3621;
  assign new_n3623 = new_n3622 ^ new_n1026;
  assign new_n3624 = new_n1036 ^ n381;
  assign new_n3625 = ~new_n990 & new_n3624;
  assign new_n3626 = new_n3625 ^ new_n1034;
  assign new_n3627 = new_n1044 ^ n382;
  assign new_n3628 = ~new_n998 & new_n3627;
  assign new_n3629 = new_n3628 ^ new_n1042;
  assign new_n3630 = new_n1052 ^ n383;
  assign new_n3631 = ~new_n1006 & new_n3630;
  assign new_n3632 = new_n3631 ^ new_n1050;
  assign new_n3633 = new_n1060 ^ n384;
  assign new_n3634 = ~new_n1014 & new_n3633;
  assign new_n3635 = new_n3634 ^ new_n1058;
  assign new_n3636 = new_n1068 ^ n385;
  assign new_n3637 = ~new_n1022 & new_n3636;
  assign new_n3638 = new_n3637 ^ new_n1066;
  assign new_n3639 = new_n1076 ^ n386;
  assign new_n3640 = ~new_n1030 & new_n3639;
  assign new_n3641 = new_n3640 ^ new_n1074;
  assign new_n3642 = new_n1084 ^ n387;
  assign new_n3643 = ~new_n1038 & new_n3642;
  assign new_n3644 = new_n3643 ^ new_n1082;
  assign new_n3645 = new_n1092 ^ n388;
  assign new_n3646 = ~new_n1046 & new_n3645;
  assign new_n3647 = new_n3646 ^ new_n1090;
  assign new_n3648 = new_n1100 ^ n389;
  assign new_n3649 = ~new_n1054 & new_n3648;
  assign new_n3650 = new_n3649 ^ new_n1098;
  assign new_n3651 = new_n1108 ^ n390;
  assign new_n3652 = ~new_n1062 & new_n3651;
  assign new_n3653 = new_n3652 ^ new_n1106;
  assign new_n3654 = new_n1116 ^ n391;
  assign new_n3655 = ~new_n1070 & new_n3654;
  assign new_n3656 = new_n3655 ^ new_n1114;
  assign new_n3657 = new_n1124 ^ n392;
  assign new_n3658 = ~new_n1078 & new_n3657;
  assign new_n3659 = new_n3658 ^ new_n1122;
  assign new_n3660 = new_n1132 ^ n393;
  assign new_n3661 = ~new_n1086 & new_n3660;
  assign new_n3662 = new_n3661 ^ new_n1130;
  assign new_n3663 = new_n1140 ^ n394;
  assign new_n3664 = ~new_n1094 & new_n3663;
  assign new_n3665 = new_n3664 ^ new_n1138;
  assign new_n3666 = new_n1148 ^ n395;
  assign new_n3667 = ~new_n1102 & new_n3666;
  assign new_n3668 = new_n3667 ^ new_n1146;
  assign new_n3669 = new_n582 ^ n396;
  assign new_n3670 = ~new_n1110 & new_n3669;
  assign new_n3671 = new_n3670 ^ new_n579;
  assign new_n3672 = new_n592 ^ n397;
  assign new_n3673 = ~new_n1118 & new_n3672;
  assign new_n3674 = new_n3673 ^ new_n589;
  assign new_n3675 = new_n602 ^ n398;
  assign new_n3676 = ~new_n1126 & new_n3675;
  assign new_n3677 = new_n3676 ^ new_n599;
  assign new_n3678 = new_n612 ^ n399;
  assign new_n3679 = ~new_n1134 & new_n3678;
  assign new_n3680 = new_n3679 ^ new_n609;
  assign new_n3681 = new_n622 ^ n400;
  assign new_n3682 = ~new_n1142 & new_n3681;
  assign new_n3683 = new_n3682 ^ new_n619;
  assign new_n3684 = new_n632 ^ n401;
  assign new_n3685 = ~new_n1150 & new_n3684;
  assign new_n3686 = new_n3685 ^ new_n629;
  assign new_n3687 = new_n642 ^ n402;
  assign new_n3688 = ~new_n584 & new_n3687;
  assign new_n3689 = new_n3688 ^ new_n639;
  assign new_n3690 = new_n652 ^ n403;
  assign new_n3691 = ~new_n594 & new_n3690;
  assign new_n3692 = new_n3691 ^ new_n649;
  assign new_n3693 = new_n662 ^ n404;
  assign new_n3694 = ~new_n604 & new_n3693;
  assign new_n3695 = new_n3694 ^ new_n659;
  assign new_n3696 = new_n672 ^ n405;
  assign new_n3697 = ~new_n614 & new_n3696;
  assign new_n3698 = new_n3697 ^ new_n669;
  assign new_n3699 = new_n682 ^ n406;
  assign new_n3700 = ~new_n624 & new_n3699;
  assign new_n3701 = new_n3700 ^ new_n679;
  assign new_n3702 = new_n692 ^ n407;
  assign new_n3703 = ~new_n634 & new_n3702;
  assign new_n3704 = new_n3703 ^ new_n689;
  assign new_n3705 = new_n702 ^ n408;
  assign new_n3706 = ~new_n644 & new_n3705;
  assign new_n3707 = new_n3706 ^ new_n699;
  assign new_n3708 = new_n712 ^ n409;
  assign new_n3709 = ~new_n654 & new_n3708;
  assign new_n3710 = new_n3709 ^ new_n709;
  assign new_n3711 = new_n722 ^ n410;
  assign new_n3712 = ~new_n664 & new_n3711;
  assign new_n3713 = new_n3712 ^ new_n719;
  assign new_n3714 = new_n732 ^ n411;
  assign new_n3715 = ~new_n674 & new_n3714;
  assign new_n3716 = new_n3715 ^ new_n729;
  assign new_n3717 = new_n742 ^ n412;
  assign new_n3718 = ~new_n684 & new_n3717;
  assign new_n3719 = new_n3718 ^ new_n739;
  assign new_n3720 = new_n752 ^ n413;
  assign new_n3721 = ~new_n694 & new_n3720;
  assign new_n3722 = new_n3721 ^ new_n749;
  assign new_n3723 = new_n762 ^ n414;
  assign new_n3724 = ~new_n704 & new_n3723;
  assign new_n3725 = new_n3724 ^ new_n759;
  assign new_n3726 = new_n772 ^ n415;
  assign new_n3727 = ~new_n714 & new_n3726;
  assign new_n3728 = new_n3727 ^ new_n769;
  assign new_n3729 = new_n782 ^ n416;
  assign new_n3730 = ~new_n724 & new_n3729;
  assign new_n3731 = new_n3730 ^ new_n779;
  assign new_n3732 = new_n792 ^ n353;
  assign new_n3733 = ~new_n734 & new_n3732;
  assign new_n3734 = new_n3733 ^ new_n789;
  assign new_n3735 = new_n801 ^ n354;
  assign new_n3736 = ~new_n744 & new_n3735;
  assign new_n3737 = new_n3736 ^ new_n799;
  assign new_n3738 = new_n810 ^ n355;
  assign new_n3739 = ~new_n754 & new_n3738;
  assign new_n3740 = new_n3739 ^ new_n808;
  assign new_n3741 = new_n819 ^ n356;
  assign new_n3742 = ~new_n764 & new_n3741;
  assign new_n3743 = new_n3742 ^ new_n817;
  assign new_n3744 = new_n828 ^ n357;
  assign new_n3745 = ~new_n774 & new_n3744;
  assign new_n3746 = new_n3745 ^ new_n826;
  assign new_n3747 = new_n837 ^ n358;
  assign new_n3748 = ~new_n784 & new_n3747;
  assign new_n3749 = new_n3748 ^ new_n835;
  assign new_n3750 = new_n846 ^ n359;
  assign new_n3751 = ~new_n794 & new_n3750;
  assign new_n3752 = new_n3751 ^ new_n844;
  assign new_n3753 = new_n855 ^ n360;
  assign new_n3754 = ~new_n803 & new_n3753;
  assign new_n3755 = new_n3754 ^ new_n853;
  assign new_n3756 = new_n864 ^ n361;
  assign new_n3757 = ~new_n812 & new_n3756;
  assign new_n3758 = new_n3757 ^ new_n862;
  assign new_n3759 = new_n873 ^ n362;
  assign new_n3760 = ~new_n821 & new_n3759;
  assign new_n3761 = new_n3760 ^ new_n871;
  assign new_n3762 = new_n882 ^ n363;
  assign new_n3763 = ~new_n830 & new_n3762;
  assign new_n3764 = new_n3763 ^ new_n880;
  assign new_n3765 = new_n891 ^ n364;
  assign new_n3766 = ~new_n839 & new_n3765;
  assign new_n3767 = new_n3766 ^ new_n889;
  assign new_n3768 = new_n900 ^ n365;
  assign new_n3769 = ~new_n848 & new_n3768;
  assign new_n3770 = new_n3769 ^ new_n898;
  assign new_n3771 = new_n909 ^ n366;
  assign new_n3772 = ~new_n857 & new_n3771;
  assign new_n3773 = new_n3772 ^ new_n907;
  assign new_n3774 = new_n918 ^ n367;
  assign new_n3775 = ~new_n866 & new_n3774;
  assign new_n3776 = new_n3775 ^ new_n916;
  assign new_n3777 = new_n1293 ^ n217;
  assign new_n3778 = ~new_n3585 & new_n3777;
  assign new_n3779 = new_n3778 ^ new_n875;
  assign new_n3780 = new_n1297 ^ n218;
  assign new_n3781 = ~new_n3588 & new_n3780;
  assign new_n3782 = new_n3781 ^ new_n884;
  assign new_n3783 = new_n1301 ^ n219;
  assign new_n3784 = ~new_n3591 & new_n3783;
  assign new_n3785 = new_n3784 ^ new_n893;
  assign new_n3786 = new_n1305 ^ n220;
  assign new_n3787 = ~new_n3594 & new_n3786;
  assign new_n3788 = new_n3787 ^ new_n902;
  assign new_n3789 = new_n1309 ^ n221;
  assign new_n3790 = ~new_n3597 & new_n3789;
  assign new_n3791 = new_n3790 ^ new_n911;
  assign new_n3792 = new_n1313 ^ n222;
  assign new_n3793 = ~new_n3600 & new_n3792;
  assign new_n3794 = new_n3793 ^ new_n920;
  assign new_n3795 = new_n1317 ^ n223;
  assign new_n3796 = ~new_n3603 & new_n3795;
  assign new_n3797 = new_n3796 ^ new_n929;
  assign new_n3798 = new_n1321 ^ n224;
  assign new_n3799 = ~new_n3606 & new_n3798;
  assign new_n3800 = new_n3799 ^ new_n938;
  assign new_n3801 = new_n1325 ^ n161;
  assign new_n3802 = ~new_n3609 & new_n3801;
  assign new_n3803 = new_n3802 ^ new_n947;
  assign new_n3804 = new_n1329 ^ n162;
  assign new_n3805 = ~new_n3612 & new_n3804;
  assign new_n3806 = new_n3805 ^ new_n956;
  assign new_n3807 = new_n1333 ^ n163;
  assign new_n3808 = ~new_n3615 & new_n3807;
  assign new_n3809 = new_n3808 ^ new_n965;
  assign new_n3810 = new_n1337 ^ n164;
  assign new_n3811 = ~new_n3618 & new_n3810;
  assign new_n3812 = new_n3811 ^ new_n974;
  assign new_n3813 = new_n1341 ^ n165;
  assign new_n3814 = ~new_n3621 & new_n3813;
  assign new_n3815 = new_n3814 ^ new_n982;
  assign new_n3816 = new_n1345 ^ n166;
  assign new_n3817 = ~new_n3624 & new_n3816;
  assign new_n3818 = new_n3817 ^ new_n990;
  assign new_n3819 = new_n1349 ^ n167;
  assign new_n3820 = ~new_n3627 & new_n3819;
  assign new_n3821 = new_n3820 ^ new_n998;
  assign new_n3822 = new_n1353 ^ n168;
  assign new_n3823 = ~new_n3630 & new_n3822;
  assign new_n3824 = new_n3823 ^ new_n1006;
  assign new_n3825 = new_n1357 ^ n169;
  assign new_n3826 = ~new_n3633 & new_n3825;
  assign new_n3827 = new_n3826 ^ new_n1014;
  assign new_n3828 = new_n1361 ^ n170;
  assign new_n3829 = ~new_n3636 & new_n3828;
  assign new_n3830 = new_n3829 ^ new_n1022;
  assign new_n3831 = new_n1365 ^ n171;
  assign new_n3832 = ~new_n3639 & new_n3831;
  assign new_n3833 = new_n3832 ^ new_n1030;
  assign new_n3834 = new_n1369 ^ n172;
  assign new_n3835 = ~new_n3642 & new_n3834;
  assign new_n3836 = new_n3835 ^ new_n1038;
  assign new_n3837 = new_n1373 ^ n173;
  assign new_n3838 = ~new_n3645 & new_n3837;
  assign new_n3839 = new_n3838 ^ new_n1046;
  assign new_n3840 = new_n1377 ^ n174;
  assign new_n3841 = ~new_n3648 & new_n3840;
  assign new_n3842 = new_n3841 ^ new_n1054;
  assign new_n3843 = new_n1381 ^ n175;
  assign new_n3844 = ~new_n3651 & new_n3843;
  assign new_n3845 = new_n3844 ^ new_n1062;
  assign new_n3846 = new_n1385 ^ n176;
  assign new_n3847 = ~new_n3654 & new_n3846;
  assign new_n3848 = new_n3847 ^ new_n1070;
  assign new_n3849 = new_n1389 ^ n177;
  assign new_n3850 = ~new_n3657 & new_n3849;
  assign new_n3851 = new_n3850 ^ new_n1078;
  assign new_n3852 = new_n1393 ^ n178;
  assign new_n3853 = ~new_n3660 & new_n3852;
  assign new_n3854 = new_n3853 ^ new_n1086;
  assign new_n3855 = new_n1397 ^ n179;
  assign new_n3856 = ~new_n3663 & new_n3855;
  assign new_n3857 = new_n3856 ^ new_n1094;
  assign new_n3858 = new_n1401 ^ n180;
  assign new_n3859 = ~new_n3666 & new_n3858;
  assign new_n3860 = new_n3859 ^ new_n1102;
  assign new_n3861 = new_n1405 ^ n181;
  assign new_n3862 = ~new_n3669 & new_n3861;
  assign new_n3863 = new_n3862 ^ new_n1110;
  assign new_n3864 = new_n1153 ^ n182;
  assign new_n3865 = ~new_n3672 & new_n3864;
  assign new_n3866 = new_n3865 ^ new_n1118;
  assign new_n3867 = new_n1157 ^ n183;
  assign new_n3868 = ~new_n3675 & new_n3867;
  assign new_n3869 = new_n3868 ^ new_n1126;
  assign new_n3870 = new_n1161 ^ n184;
  assign new_n3871 = ~new_n3678 & new_n3870;
  assign new_n3872 = new_n3871 ^ new_n1134;
  assign new_n3873 = new_n1165 ^ n185;
  assign new_n3874 = ~new_n3681 & new_n3873;
  assign new_n3875 = new_n3874 ^ new_n1142;
  assign new_n3876 = new_n1169 ^ n186;
  assign new_n3877 = ~new_n3684 & new_n3876;
  assign new_n3878 = new_n3877 ^ new_n1150;
  assign new_n3879 = new_n1173 ^ n187;
  assign new_n3880 = ~new_n3687 & new_n3879;
  assign new_n3881 = new_n3880 ^ new_n584;
  assign new_n3882 = new_n1177 ^ n188;
  assign new_n3883 = ~new_n3690 & new_n3882;
  assign new_n3884 = new_n3883 ^ new_n594;
  assign new_n3885 = new_n1181 ^ n189;
  assign new_n3886 = ~new_n3693 & new_n3885;
  assign new_n3887 = new_n3886 ^ new_n604;
  assign new_n3888 = new_n1185 ^ n190;
  assign new_n3889 = ~new_n3696 & new_n3888;
  assign new_n3890 = new_n3889 ^ new_n614;
  assign new_n3891 = new_n1189 ^ n191;
  assign new_n3892 = ~new_n3699 & new_n3891;
  assign new_n3893 = new_n3892 ^ new_n624;
  assign new_n3894 = new_n1193 ^ n192;
  assign new_n3895 = ~new_n3702 & new_n3894;
  assign new_n3896 = new_n3895 ^ new_n634;
  assign new_n3897 = new_n1197 ^ n193;
  assign new_n3898 = ~new_n3705 & new_n3897;
  assign new_n3899 = new_n3898 ^ new_n644;
  assign new_n3900 = new_n1201 ^ n194;
  assign new_n3901 = ~new_n3708 & new_n3900;
  assign new_n3902 = new_n3901 ^ new_n654;
  assign new_n3903 = new_n1205 ^ n195;
  assign new_n3904 = ~new_n3711 & new_n3903;
  assign new_n3905 = new_n3904 ^ new_n664;
  assign new_n3906 = new_n1209 ^ n196;
  assign new_n3907 = ~new_n3714 & new_n3906;
  assign new_n3908 = new_n3907 ^ new_n674;
  assign new_n3909 = new_n1213 ^ n197;
  assign new_n3910 = ~new_n3717 & new_n3909;
  assign new_n3911 = new_n3910 ^ new_n684;
  assign new_n3912 = new_n1217 ^ n198;
  assign new_n3913 = ~new_n3720 & new_n3912;
  assign new_n3914 = new_n3913 ^ new_n694;
  assign new_n3915 = new_n1221 ^ n199;
  assign new_n3916 = ~new_n3723 & new_n3915;
  assign new_n3917 = new_n3916 ^ new_n704;
  assign new_n3918 = new_n1225 ^ n200;
  assign new_n3919 = ~new_n3726 & new_n3918;
  assign new_n3920 = new_n3919 ^ new_n714;
  assign new_n3921 = new_n1229 ^ n201;
  assign new_n3922 = ~new_n3729 & new_n3921;
  assign new_n3923 = new_n3922 ^ new_n724;
  assign new_n3924 = new_n1233 ^ n202;
  assign new_n3925 = ~new_n3732 & new_n3924;
  assign new_n3926 = new_n3925 ^ new_n734;
  assign new_n3927 = new_n1237 ^ n203;
  assign new_n3928 = ~new_n3735 & new_n3927;
  assign new_n3929 = new_n3928 ^ new_n744;
  assign new_n3930 = new_n1241 ^ n204;
  assign new_n3931 = ~new_n3738 & new_n3930;
  assign new_n3932 = new_n3931 ^ new_n754;
  assign new_n3933 = new_n1245 ^ n205;
  assign new_n3934 = ~new_n3741 & new_n3933;
  assign new_n3935 = new_n3934 ^ new_n764;
  assign new_n3936 = new_n1249 ^ n206;
  assign new_n3937 = ~new_n3744 & new_n3936;
  assign new_n3938 = new_n3937 ^ new_n774;
  assign new_n3939 = new_n1253 ^ n207;
  assign new_n3940 = ~new_n3747 & new_n3939;
  assign new_n3941 = new_n3940 ^ new_n784;
  assign new_n3942 = new_n1257 ^ n208;
  assign new_n3943 = ~new_n3750 & new_n3942;
  assign new_n3944 = new_n3943 ^ new_n794;
  assign new_n3945 = new_n1261 ^ n209;
  assign new_n3946 = ~new_n3753 & new_n3945;
  assign new_n3947 = new_n3946 ^ new_n803;
  assign new_n3948 = new_n1265 ^ n210;
  assign new_n3949 = ~new_n3756 & new_n3948;
  assign new_n3950 = new_n3949 ^ new_n812;
  assign new_n3951 = new_n1269 ^ n211;
  assign new_n3952 = ~new_n3759 & new_n3951;
  assign new_n3953 = new_n3952 ^ new_n821;
  assign new_n3954 = new_n1273 ^ n212;
  assign new_n3955 = ~new_n3762 & new_n3954;
  assign new_n3956 = new_n3955 ^ new_n830;
  assign new_n3957 = new_n1277 ^ n213;
  assign new_n3958 = ~new_n3765 & new_n3957;
  assign new_n3959 = new_n3958 ^ new_n839;
  assign new_n3960 = new_n1281 ^ n214;
  assign new_n3961 = ~new_n3768 & new_n3960;
  assign new_n3962 = new_n3961 ^ new_n848;
  assign new_n3963 = new_n1285 ^ n215;
  assign new_n3964 = ~new_n3771 & new_n3963;
  assign new_n3965 = new_n3964 ^ new_n857;
  assign new_n3966 = new_n1289 ^ n216;
  assign new_n3967 = ~new_n3774 & new_n3966;
  assign new_n3968 = new_n3967 ^ new_n866;
  assign new_n3969 = ~new_n3777 & new_n1461;
  assign new_n3970 = new_n3969 ^ new_n3585;
  assign new_n3971 = ~new_n3780 & new_n1465;
  assign new_n3972 = new_n3971 ^ new_n3588;
  assign new_n3973 = ~new_n3783 & new_n1469;
  assign new_n3974 = new_n3973 ^ new_n3591;
  assign new_n3975 = ~new_n3786 & new_n1473;
  assign new_n3976 = new_n3975 ^ new_n3594;
  assign new_n3977 = ~new_n3789 & new_n1477;
  assign new_n3978 = new_n3977 ^ new_n3597;
  assign new_n3979 = ~new_n3792 & new_n1481;
  assign new_n3980 = new_n3979 ^ new_n3600;
  assign new_n3981 = ~new_n3795 & new_n1485;
  assign new_n3982 = new_n3981 ^ new_n3603;
  assign new_n3983 = ~new_n3798 & new_n1489;
  assign new_n3984 = new_n3983 ^ new_n3606;
  assign new_n3985 = ~new_n3801 & new_n1493;
  assign new_n3986 = new_n3985 ^ new_n3609;
  assign new_n3987 = ~new_n3804 & new_n1497;
  assign new_n3988 = new_n3987 ^ new_n3612;
  assign new_n3989 = ~new_n3807 & new_n1501;
  assign new_n3990 = new_n3989 ^ new_n3615;
  assign new_n3991 = ~new_n3810 & new_n1505;
  assign new_n3992 = new_n3991 ^ new_n3618;
  assign new_n3993 = ~new_n3813 & new_n1509;
  assign new_n3994 = new_n3993 ^ new_n3621;
  assign new_n3995 = ~new_n3816 & new_n1513;
  assign new_n3996 = new_n3995 ^ new_n3624;
  assign new_n3997 = ~new_n3819 & new_n1517;
  assign new_n3998 = new_n3997 ^ new_n3627;
  assign new_n3999 = ~new_n3822 & new_n1521;
  assign new_n4000 = new_n3999 ^ new_n3630;
  assign new_n4001 = ~new_n3825 & new_n1525;
  assign new_n4002 = new_n4001 ^ new_n3633;
  assign new_n4003 = ~new_n3828 & new_n1529;
  assign new_n4004 = new_n4003 ^ new_n3636;
  assign new_n4005 = ~new_n3831 & new_n1533;
  assign new_n4006 = new_n4005 ^ new_n3639;
  assign new_n4007 = ~new_n3834 & new_n1537;
  assign new_n4008 = new_n4007 ^ new_n3642;
  assign new_n4009 = ~new_n3837 & new_n1541;
  assign new_n4010 = new_n4009 ^ new_n3645;
  assign new_n4011 = ~new_n3840 & new_n1545;
  assign new_n4012 = new_n4011 ^ new_n3648;
  assign new_n4013 = ~new_n3843 & new_n1549;
  assign new_n4014 = new_n4013 ^ new_n3651;
  assign new_n4015 = ~new_n3846 & new_n1553;
  assign new_n4016 = new_n4015 ^ new_n3654;
  assign new_n4017 = ~new_n3849 & new_n1557;
  assign new_n4018 = new_n4017 ^ new_n3657;
  assign new_n4019 = ~new_n3852 & new_n1561;
  assign new_n4020 = new_n4019 ^ new_n3660;
  assign new_n4021 = ~new_n3855 & new_n1565;
  assign new_n4022 = new_n4021 ^ new_n3663;
  assign new_n4023 = ~new_n3858 & new_n1569;
  assign new_n4024 = new_n4023 ^ new_n3666;
  assign new_n4025 = ~new_n3861 & new_n1573;
  assign new_n4026 = new_n4025 ^ new_n3669;
  assign new_n4027 = ~new_n3864 & new_n1577;
  assign new_n4028 = new_n4027 ^ new_n3672;
  assign new_n4029 = ~new_n3867 & new_n1581;
  assign new_n4030 = new_n4029 ^ new_n3675;
  assign new_n4031 = ~new_n3870 & new_n1585;
  assign new_n4032 = new_n4031 ^ new_n3678;
  assign new_n4033 = ~new_n3873 & new_n1589;
  assign new_n4034 = new_n4033 ^ new_n3681;
  assign new_n4035 = ~new_n3876 & new_n1593;
  assign new_n4036 = new_n4035 ^ new_n3684;
  assign new_n4037 = ~new_n3879 & new_n1597;
  assign new_n4038 = new_n4037 ^ new_n3687;
  assign new_n4039 = ~new_n3882 & new_n1601;
  assign new_n4040 = new_n4039 ^ new_n3690;
  assign new_n4041 = ~new_n3885 & new_n1605;
  assign new_n4042 = new_n4041 ^ new_n3693;
  assign new_n4043 = ~new_n3888 & new_n1609;
  assign new_n4044 = new_n4043 ^ new_n3696;
  assign new_n4045 = ~new_n3891 & new_n1613;
  assign new_n4046 = new_n4045 ^ new_n3699;
  assign new_n4047 = ~new_n3894 & new_n1617;
  assign new_n4048 = new_n4047 ^ new_n3702;
  assign new_n4049 = ~new_n3897 & new_n1621;
  assign new_n4050 = new_n4049 ^ new_n3705;
  assign new_n4051 = ~new_n3900 & new_n1625;
  assign new_n4052 = new_n4051 ^ new_n3708;
  assign new_n4053 = ~new_n3903 & new_n1629;
  assign new_n4054 = new_n4053 ^ new_n3711;
  assign new_n4055 = ~new_n3906 & new_n1633;
  assign new_n4056 = new_n4055 ^ new_n3714;
  assign new_n4057 = ~new_n3909 & new_n1637;
  assign new_n4058 = new_n4057 ^ new_n3717;
  assign new_n4059 = ~new_n3912 & new_n1641;
  assign new_n4060 = new_n4059 ^ new_n3720;
  assign new_n4061 = ~new_n3915 & new_n1645;
  assign new_n4062 = new_n4061 ^ new_n3723;
  assign new_n4063 = ~new_n3918 & new_n1649;
  assign new_n4064 = new_n4063 ^ new_n3726;
  assign new_n4065 = ~new_n3921 & new_n1653;
  assign new_n4066 = new_n4065 ^ new_n3729;
  assign new_n4067 = ~new_n3924 & new_n1657;
  assign new_n4068 = new_n4067 ^ new_n3732;
  assign new_n4069 = ~new_n3927 & new_n1661;
  assign new_n4070 = new_n4069 ^ new_n3735;
  assign new_n4071 = ~new_n3930 & new_n1409;
  assign new_n4072 = new_n4071 ^ new_n3738;
  assign new_n4073 = ~new_n3933 & new_n1413;
  assign new_n4074 = new_n4073 ^ new_n3741;
  assign new_n4075 = ~new_n3936 & new_n1417;
  assign new_n4076 = new_n4075 ^ new_n3744;
  assign new_n4077 = ~new_n3939 & new_n1421;
  assign new_n4078 = new_n4077 ^ new_n3747;
  assign new_n4079 = ~new_n3942 & new_n1425;
  assign new_n4080 = new_n4079 ^ new_n3750;
  assign new_n4081 = ~new_n3945 & new_n1429;
  assign new_n4082 = new_n4081 ^ new_n3753;
  assign new_n4083 = ~new_n3948 & new_n1433;
  assign new_n4084 = new_n4083 ^ new_n3756;
  assign new_n4085 = ~new_n3951 & new_n1437;
  assign new_n4086 = new_n4085 ^ new_n3759;
  assign new_n4087 = ~new_n3954 & new_n1441;
  assign new_n4088 = new_n4087 ^ new_n3762;
  assign new_n4089 = ~new_n3957 & new_n1445;
  assign new_n4090 = new_n4089 ^ new_n3765;
  assign new_n4091 = ~new_n3960 & new_n1449;
  assign new_n4092 = new_n4091 ^ new_n3768;
  assign new_n4093 = ~new_n3963 & new_n1453;
  assign new_n4094 = new_n4093 ^ new_n3771;
  assign new_n4095 = ~new_n3966 & new_n1457;
  assign new_n4096 = new_n4095 ^ new_n3774;
  assign new_n4097 = ~new_n1461 & new_n925;
  assign new_n4098 = new_n4097 ^ new_n3777;
  assign new_n4099 = ~new_n1465 & new_n934;
  assign new_n4100 = new_n4099 ^ new_n3780;
  assign new_n4101 = ~new_n1469 & new_n943;
  assign new_n4102 = new_n4101 ^ new_n3783;
  assign new_n4103 = ~new_n1473 & new_n952;
  assign new_n4104 = new_n4103 ^ new_n3786;
  assign new_n4105 = ~new_n1477 & new_n961;
  assign new_n4106 = new_n4105 ^ new_n3789;
  assign new_n4107 = ~new_n1481 & new_n970;
  assign new_n4108 = new_n4107 ^ new_n3792;
  assign new_n4109 = ~new_n1485 & new_n978;
  assign new_n4110 = new_n4109 ^ new_n3795;
  assign new_n4111 = ~new_n1489 & new_n986;
  assign new_n4112 = new_n4111 ^ new_n3798;
  assign new_n4113 = ~new_n1493 & new_n994;
  assign new_n4114 = new_n4113 ^ new_n3801;
  assign new_n4115 = ~new_n1497 & new_n1002;
  assign new_n4116 = new_n4115 ^ new_n3804;
  assign new_n4117 = ~new_n1501 & new_n1010;
  assign new_n4118 = new_n4117 ^ new_n3807;
  assign new_n4119 = ~new_n1505 & new_n1018;
  assign new_n4120 = new_n4119 ^ new_n3810;
  assign new_n4121 = ~new_n1509 & new_n1026;
  assign new_n4122 = new_n4121 ^ new_n3813;
  assign new_n4123 = ~new_n1513 & new_n1034;
  assign new_n4124 = new_n4123 ^ new_n3816;
  assign new_n4125 = ~new_n1517 & new_n1042;
  assign new_n4126 = new_n4125 ^ new_n3819;
  assign new_n4127 = ~new_n1521 & new_n1050;
  assign new_n4128 = new_n4127 ^ new_n3822;
  assign new_n4129 = ~new_n1525 & new_n1058;
  assign new_n4130 = new_n4129 ^ new_n3825;
  assign new_n4131 = ~new_n1529 & new_n1066;
  assign new_n4132 = new_n4131 ^ new_n3828;
  assign new_n4133 = ~new_n1533 & new_n1074;
  assign new_n4134 = new_n4133 ^ new_n3831;
  assign new_n4135 = ~new_n1537 & new_n1082;
  assign new_n4136 = new_n4135 ^ new_n3834;
  assign new_n4137 = ~new_n1541 & new_n1090;
  assign new_n4138 = new_n4137 ^ new_n3837;
  assign new_n4139 = ~new_n1545 & new_n1098;
  assign new_n4140 = new_n4139 ^ new_n3840;
  assign new_n4141 = ~new_n1549 & new_n1106;
  assign new_n4142 = new_n4141 ^ new_n3843;
  assign new_n4143 = ~new_n1553 & new_n1114;
  assign new_n4144 = new_n4143 ^ new_n3846;
  assign new_n4145 = ~new_n1557 & new_n1122;
  assign new_n4146 = new_n4145 ^ new_n3849;
  assign new_n4147 = ~new_n1561 & new_n1130;
  assign new_n4148 = new_n4147 ^ new_n3852;
  assign new_n4149 = ~new_n1565 & new_n1138;
  assign new_n4150 = new_n4149 ^ new_n3855;
  assign new_n4151 = ~new_n1569 & new_n1146;
  assign new_n4152 = new_n4151 ^ new_n3858;
  assign new_n4153 = ~new_n1573 & new_n579;
  assign new_n4154 = new_n4153 ^ new_n3861;
  assign new_n4155 = ~new_n1577 & new_n589;
  assign new_n4156 = new_n4155 ^ new_n3864;
  assign new_n4157 = ~new_n1581 & new_n599;
  assign new_n4158 = new_n4157 ^ new_n3867;
  assign new_n4159 = ~new_n1585 & new_n609;
  assign new_n4160 = new_n4159 ^ new_n3870;
  assign new_n4161 = ~new_n1589 & new_n619;
  assign new_n4162 = new_n4161 ^ new_n3873;
  assign new_n4163 = ~new_n1593 & new_n629;
  assign new_n4164 = new_n4163 ^ new_n3876;
  assign new_n4165 = ~new_n1597 & new_n639;
  assign new_n4166 = new_n4165 ^ new_n3879;
  assign new_n4167 = ~new_n1601 & new_n649;
  assign new_n4168 = new_n4167 ^ new_n3882;
  assign new_n4169 = ~new_n1605 & new_n659;
  assign new_n4170 = new_n4169 ^ new_n3885;
  assign new_n4171 = ~new_n1609 & new_n669;
  assign new_n4172 = new_n4171 ^ new_n3888;
  assign new_n4173 = ~new_n1613 & new_n679;
  assign new_n4174 = new_n4173 ^ new_n3891;
  assign new_n4175 = ~new_n1617 & new_n689;
  assign new_n4176 = new_n4175 ^ new_n3894;
  assign new_n4177 = ~new_n1621 & new_n699;
  assign new_n4178 = new_n4177 ^ new_n3897;
  assign new_n4179 = ~new_n1625 & new_n709;
  assign new_n4180 = new_n4179 ^ new_n3900;
  assign new_n4181 = ~new_n1629 & new_n719;
  assign new_n4182 = new_n4181 ^ new_n3903;
  assign new_n4183 = ~new_n1633 & new_n729;
  assign new_n4184 = new_n4183 ^ new_n3906;
  assign new_n4185 = ~new_n1637 & new_n739;
  assign new_n4186 = new_n4185 ^ new_n3909;
  assign new_n4187 = ~new_n1641 & new_n749;
  assign new_n4188 = new_n4187 ^ new_n3912;
  assign new_n4189 = ~new_n1645 & new_n759;
  assign new_n4190 = new_n4189 ^ new_n3915;
  assign new_n4191 = ~new_n1649 & new_n769;
  assign new_n4192 = new_n4191 ^ new_n3918;
  assign new_n4193 = ~new_n1653 & new_n779;
  assign new_n4194 = new_n4193 ^ new_n3921;
  assign new_n4195 = ~new_n1657 & new_n789;
  assign new_n4196 = new_n4195 ^ new_n3924;
  assign new_n4197 = ~new_n1661 & new_n799;
  assign new_n4198 = new_n4197 ^ new_n3927;
  assign new_n4199 = ~new_n1409 & new_n808;
  assign new_n4200 = new_n4199 ^ new_n3930;
  assign new_n4201 = ~new_n1413 & new_n817;
  assign new_n4202 = new_n4201 ^ new_n3933;
  assign new_n4203 = ~new_n1417 & new_n826;
  assign new_n4204 = new_n4203 ^ new_n3936;
  assign new_n4205 = ~new_n1421 & new_n835;
  assign new_n4206 = new_n4205 ^ new_n3939;
  assign new_n4207 = ~new_n1425 & new_n844;
  assign new_n4208 = new_n4207 ^ new_n3942;
  assign new_n4209 = ~new_n1429 & new_n853;
  assign new_n4210 = new_n4209 ^ new_n3945;
  assign new_n4211 = ~new_n1433 & new_n862;
  assign new_n4212 = new_n4211 ^ new_n3948;
  assign new_n4213 = ~new_n1437 & new_n871;
  assign new_n4214 = new_n4213 ^ new_n3951;
  assign new_n4215 = ~new_n1441 & new_n880;
  assign new_n4216 = new_n4215 ^ new_n3954;
  assign new_n4217 = ~new_n1445 & new_n889;
  assign new_n4218 = new_n4217 ^ new_n3957;
  assign new_n4219 = ~new_n1449 & new_n898;
  assign new_n4220 = new_n4219 ^ new_n3960;
  assign new_n4221 = ~new_n1453 & new_n907;
  assign new_n4222 = new_n4221 ^ new_n3963;
  assign new_n4223 = ~new_n1457 & new_n916;
  assign new_n4224 = new_n4223 ^ new_n3966;
  assign new_n4225 = ~new_n1289 & new_n1509;
  assign new_n4226 = new_n4225 ^ new_n772;
  assign new_n4227 = ~new_n1293 & new_n1513;
  assign new_n4228 = new_n4227 ^ new_n782;
  assign new_n4229 = ~new_n1297 & new_n1517;
  assign new_n4230 = new_n4229 ^ new_n792;
  assign new_n4231 = ~new_n1301 & new_n1521;
  assign new_n4232 = new_n4231 ^ new_n801;
  assign new_n4233 = ~new_n1305 & new_n1525;
  assign new_n4234 = new_n4233 ^ new_n810;
  assign new_n4235 = ~new_n1309 & new_n1529;
  assign new_n4236 = new_n4235 ^ new_n819;
  assign new_n4237 = ~new_n1313 & new_n1533;
  assign new_n4238 = new_n4237 ^ new_n828;
  assign new_n4239 = ~new_n1317 & new_n1537;
  assign new_n4240 = new_n4239 ^ new_n837;
  assign new_n4241 = ~new_n1321 & new_n1541;
  assign new_n4242 = new_n4241 ^ new_n846;
  assign new_n4243 = ~new_n1325 & new_n1545;
  assign new_n4244 = new_n4243 ^ new_n855;
  assign new_n4245 = ~new_n1329 & new_n1549;
  assign new_n4246 = new_n4245 ^ new_n864;
  assign new_n4247 = ~new_n1333 & new_n1553;
  assign new_n4248 = new_n4247 ^ new_n873;
  assign new_n4249 = ~new_n1337 & new_n1557;
  assign new_n4250 = new_n4249 ^ new_n882;
  assign new_n4251 = ~new_n1341 & new_n1561;
  assign new_n4252 = new_n4251 ^ new_n891;
  assign new_n4253 = ~new_n1345 & new_n1565;
  assign new_n4254 = new_n4253 ^ new_n900;
  assign new_n4255 = ~new_n1349 & new_n1569;
  assign new_n4256 = new_n4255 ^ new_n909;
  assign new_n4257 = ~new_n1353 & new_n1573;
  assign new_n4258 = new_n4257 ^ new_n918;
  assign new_n4259 = ~new_n1357 & new_n1577;
  assign new_n4260 = new_n4259 ^ new_n927;
  assign new_n4261 = ~new_n1361 & new_n1581;
  assign new_n4262 = new_n4261 ^ new_n936;
  assign new_n4263 = ~new_n1365 & new_n1585;
  assign new_n4264 = new_n4263 ^ new_n945;
  assign new_n4265 = ~new_n1369 & new_n1589;
  assign new_n4266 = new_n4265 ^ new_n954;
  assign new_n4267 = ~new_n1373 & new_n1593;
  assign new_n4268 = new_n4267 ^ new_n963;
  assign new_n4269 = ~new_n1377 & new_n1597;
  assign new_n4270 = new_n4269 ^ new_n972;
  assign new_n4271 = ~new_n1381 & new_n1601;
  assign new_n4272 = new_n4271 ^ new_n980;
  assign new_n4273 = ~new_n1385 & new_n1605;
  assign new_n4274 = new_n4273 ^ new_n988;
  assign new_n4275 = ~new_n1389 & new_n1609;
  assign new_n4276 = new_n4275 ^ new_n996;
  assign new_n4277 = ~new_n1393 & new_n1613;
  assign new_n4278 = new_n4277 ^ new_n1004;
  assign new_n4279 = ~new_n1397 & new_n1617;
  assign new_n4280 = new_n4279 ^ new_n1012;
  assign new_n4281 = ~new_n1401 & new_n1621;
  assign new_n4282 = new_n4281 ^ new_n1020;
  assign new_n4283 = ~new_n1405 & new_n1625;
  assign new_n4284 = new_n4283 ^ new_n1028;
  assign new_n4285 = ~new_n1153 & new_n1629;
  assign new_n4286 = new_n4285 ^ new_n1036;
  assign new_n4287 = ~new_n1157 & new_n1633;
  assign new_n4288 = new_n4287 ^ new_n1044;
  assign new_n4289 = ~new_n1161 & new_n1637;
  assign new_n4290 = new_n4289 ^ new_n1052;
  assign new_n4291 = ~new_n1165 & new_n1641;
  assign new_n4292 = new_n4291 ^ new_n1060;
  assign new_n4293 = ~new_n1169 & new_n1645;
  assign new_n4294 = new_n4293 ^ new_n1068;
  assign new_n4295 = ~new_n1173 & new_n1649;
  assign new_n4296 = new_n4295 ^ new_n1076;
  assign new_n4297 = ~new_n1177 & new_n1653;
  assign new_n4298 = new_n4297 ^ new_n1084;
  assign new_n4299 = ~new_n1181 & new_n1657;
  assign new_n4300 = new_n4299 ^ new_n1092;
  assign new_n4301 = ~new_n1185 & new_n1661;
  assign new_n4302 = new_n4301 ^ new_n1100;
  assign new_n4303 = ~new_n1189 & new_n1409;
  assign new_n4304 = new_n4303 ^ new_n1108;
  assign new_n4305 = ~new_n1193 & new_n1413;
  assign new_n4306 = new_n4305 ^ new_n1116;
  assign new_n4307 = ~new_n1197 & new_n1417;
  assign new_n4308 = new_n4307 ^ new_n1124;
  assign new_n4309 = ~new_n1201 & new_n1421;
  assign new_n4310 = new_n4309 ^ new_n1132;
  assign new_n4311 = ~new_n1205 & new_n1425;
  assign new_n4312 = new_n4311 ^ new_n1140;
  assign new_n4313 = ~new_n1209 & new_n1429;
  assign new_n4314 = new_n4313 ^ new_n1148;
  assign new_n4315 = ~new_n1213 & new_n1433;
  assign new_n4316 = new_n4315 ^ new_n582;
  assign new_n4317 = ~new_n1217 & new_n1437;
  assign new_n4318 = new_n4317 ^ new_n592;
  assign new_n4319 = ~new_n1221 & new_n1441;
  assign new_n4320 = new_n4319 ^ new_n602;
  assign new_n4321 = ~new_n1225 & new_n1445;
  assign new_n4322 = new_n4321 ^ new_n612;
  assign new_n4323 = ~new_n1229 & new_n1449;
  assign new_n4324 = new_n4323 ^ new_n622;
  assign new_n4325 = ~new_n1233 & new_n1453;
  assign new_n4326 = new_n4325 ^ new_n632;
  assign new_n4327 = ~new_n1237 & new_n1457;
  assign new_n4328 = new_n4327 ^ new_n642;
  assign new_n4329 = ~new_n1241 & new_n1461;
  assign new_n4330 = new_n4329 ^ new_n652;
  assign new_n4331 = ~new_n1245 & new_n1465;
  assign new_n4332 = new_n4331 ^ new_n662;
  assign new_n4333 = ~new_n1249 & new_n1469;
  assign new_n4334 = new_n4333 ^ new_n672;
  assign new_n4335 = ~new_n1253 & new_n1473;
  assign new_n4336 = new_n4335 ^ new_n682;
  assign new_n4337 = ~new_n1257 & new_n1477;
  assign new_n4338 = new_n4337 ^ new_n692;
  assign new_n4339 = ~new_n1261 & new_n1481;
  assign new_n4340 = new_n4339 ^ new_n702;
  assign new_n4341 = ~new_n1265 & new_n1485;
  assign new_n4342 = new_n4341 ^ new_n712;
  assign new_n4343 = ~new_n1269 & new_n1489;
  assign new_n4344 = new_n4343 ^ new_n722;
  assign new_n4345 = ~new_n1273 & new_n1493;
  assign new_n4346 = new_n4345 ^ new_n732;
  assign new_n4347 = ~new_n1277 & new_n1497;
  assign new_n4348 = new_n4347 ^ new_n742;
  assign new_n4349 = ~new_n1281 & new_n1501;
  assign new_n4350 = new_n4349 ^ new_n752;
  assign new_n4351 = ~new_n1285 & new_n1505;
  assign new_n4352 = new_n4351 ^ new_n762;
  assign new_n4353 = ~new_n1509 & new_n970;
  assign new_n4354 = new_n4353 ^ new_n1289;
  assign new_n4355 = ~new_n1513 & new_n978;
  assign new_n4356 = new_n4355 ^ new_n1293;
  assign new_n4357 = ~new_n1517 & new_n986;
  assign new_n4358 = new_n4357 ^ new_n1297;
  assign new_n4359 = ~new_n1521 & new_n994;
  assign new_n4360 = new_n4359 ^ new_n1301;
  assign new_n4361 = ~new_n1525 & new_n1002;
  assign new_n4362 = new_n4361 ^ new_n1305;
  assign new_n4363 = ~new_n1529 & new_n1010;
  assign new_n4364 = new_n4363 ^ new_n1309;
  assign new_n4365 = ~new_n1533 & new_n1018;
  assign new_n4366 = new_n4365 ^ new_n1313;
  assign new_n4367 = ~new_n1537 & new_n1026;
  assign new_n4368 = new_n4367 ^ new_n1317;
  assign new_n4369 = ~new_n1541 & new_n1034;
  assign new_n4370 = new_n4369 ^ new_n1321;
  assign new_n4371 = ~new_n1545 & new_n1042;
  assign new_n4372 = new_n4371 ^ new_n1325;
  assign new_n4373 = ~new_n1549 & new_n1050;
  assign new_n4374 = new_n4373 ^ new_n1329;
  assign new_n4375 = ~new_n1553 & new_n1058;
  assign new_n4376 = new_n4375 ^ new_n1333;
  assign new_n4377 = ~new_n1557 & new_n1066;
  assign new_n4378 = new_n4377 ^ new_n1337;
  assign new_n4379 = ~new_n1561 & new_n1074;
  assign new_n4380 = new_n4379 ^ new_n1341;
  assign new_n4381 = ~new_n1565 & new_n1082;
  assign new_n4382 = new_n4381 ^ new_n1345;
  assign new_n4383 = ~new_n1569 & new_n1090;
  assign new_n4384 = new_n4383 ^ new_n1349;
  assign new_n4385 = ~new_n1573 & new_n1098;
  assign new_n4386 = new_n4385 ^ new_n1353;
  assign new_n4387 = ~new_n1577 & new_n1106;
  assign new_n4388 = new_n4387 ^ new_n1357;
  assign new_n4389 = ~new_n1581 & new_n1114;
  assign new_n4390 = new_n4389 ^ new_n1361;
  assign new_n4391 = ~new_n1585 & new_n1122;
  assign new_n4392 = new_n4391 ^ new_n1365;
  assign new_n4393 = ~new_n1589 & new_n1130;
  assign new_n4394 = new_n4393 ^ new_n1369;
  assign new_n4395 = ~new_n1593 & new_n1138;
  assign new_n4396 = new_n4395 ^ new_n1373;
  assign new_n4397 = ~new_n1597 & new_n1146;
  assign new_n4398 = new_n4397 ^ new_n1377;
  assign new_n4399 = ~new_n1601 & new_n579;
  assign new_n4400 = new_n4399 ^ new_n1381;
  assign new_n4401 = ~new_n1605 & new_n589;
  assign new_n4402 = new_n4401 ^ new_n1385;
  assign new_n4403 = ~new_n1609 & new_n599;
  assign new_n4404 = new_n4403 ^ new_n1389;
  assign new_n4405 = ~new_n1613 & new_n609;
  assign new_n4406 = new_n4405 ^ new_n1393;
  assign new_n4407 = ~new_n1617 & new_n619;
  assign new_n4408 = new_n4407 ^ new_n1397;
  assign new_n4409 = ~new_n1621 & new_n629;
  assign new_n4410 = new_n4409 ^ new_n1401;
  assign new_n4411 = ~new_n1625 & new_n639;
  assign new_n4412 = new_n4411 ^ new_n1405;
  assign new_n4413 = ~new_n1629 & new_n649;
  assign new_n4414 = new_n4413 ^ new_n1153;
  assign new_n4415 = ~new_n1633 & new_n659;
  assign new_n4416 = new_n4415 ^ new_n1157;
  assign new_n4417 = ~new_n1637 & new_n669;
  assign new_n4418 = new_n4417 ^ new_n1161;
  assign new_n4419 = ~new_n1641 & new_n679;
  assign new_n4420 = new_n4419 ^ new_n1165;
  assign new_n4421 = ~new_n1645 & new_n689;
  assign new_n4422 = new_n4421 ^ new_n1169;
  assign new_n4423 = ~new_n1649 & new_n699;
  assign new_n4424 = new_n4423 ^ new_n1173;
  assign new_n4425 = ~new_n1653 & new_n709;
  assign new_n4426 = new_n4425 ^ new_n1177;
  assign new_n4427 = ~new_n1657 & new_n719;
  assign new_n4428 = new_n4427 ^ new_n1181;
  assign new_n4429 = ~new_n1661 & new_n729;
  assign new_n4430 = new_n4429 ^ new_n1185;
  assign new_n4431 = ~new_n1409 & new_n739;
  assign new_n4432 = new_n4431 ^ new_n1189;
  assign new_n4433 = ~new_n1413 & new_n749;
  assign new_n4434 = new_n4433 ^ new_n1193;
  assign new_n4435 = ~new_n1417 & new_n759;
  assign new_n4436 = new_n4435 ^ new_n1197;
  assign new_n4437 = ~new_n1421 & new_n769;
  assign new_n4438 = new_n4437 ^ new_n1201;
  assign new_n4439 = ~new_n1425 & new_n779;
  assign new_n4440 = new_n4439 ^ new_n1205;
  assign new_n4441 = ~new_n1429 & new_n789;
  assign new_n4442 = new_n4441 ^ new_n1209;
  assign new_n4443 = ~new_n1433 & new_n799;
  assign new_n4444 = new_n4443 ^ new_n1213;
  assign new_n4445 = ~new_n1437 & new_n808;
  assign new_n4446 = new_n4445 ^ new_n1217;
  assign new_n4447 = ~new_n1441 & new_n817;
  assign new_n4448 = new_n4447 ^ new_n1221;
  assign new_n4449 = ~new_n1445 & new_n826;
  assign new_n4450 = new_n4449 ^ new_n1225;
  assign new_n4451 = ~new_n1449 & new_n835;
  assign new_n4452 = new_n4451 ^ new_n1229;
  assign new_n4453 = ~new_n1453 & new_n844;
  assign new_n4454 = new_n4453 ^ new_n1233;
  assign new_n4455 = ~new_n1457 & new_n853;
  assign new_n4456 = new_n4455 ^ new_n1237;
  assign new_n4457 = ~new_n1461 & new_n862;
  assign new_n4458 = new_n4457 ^ new_n1241;
  assign new_n4459 = ~new_n1465 & new_n871;
  assign new_n4460 = new_n4459 ^ new_n1245;
  assign new_n4461 = ~new_n1469 & new_n880;
  assign new_n4462 = new_n4461 ^ new_n1249;
  assign new_n4463 = ~new_n1473 & new_n889;
  assign new_n4464 = new_n4463 ^ new_n1253;
  assign new_n4465 = ~new_n1477 & new_n898;
  assign new_n4466 = new_n4465 ^ new_n1257;
  assign new_n4467 = ~new_n1481 & new_n907;
  assign new_n4468 = new_n4467 ^ new_n1261;
  assign new_n4469 = ~new_n1485 & new_n916;
  assign new_n4470 = new_n4469 ^ new_n1265;
  assign new_n4471 = ~new_n1489 & new_n925;
  assign new_n4472 = new_n4471 ^ new_n1269;
  assign new_n4473 = ~new_n1493 & new_n934;
  assign new_n4474 = new_n4473 ^ new_n1273;
  assign new_n4475 = ~new_n1497 & new_n943;
  assign new_n4476 = new_n4475 ^ new_n1277;
  assign new_n4477 = ~new_n1501 & new_n952;
  assign new_n4478 = new_n4477 ^ new_n1281;
  assign new_n4479 = ~new_n1505 & new_n961;
  assign new_n4480 = new_n4479 ^ new_n1285;
  assign new_n4481 = new_n803 ^ n35;
  assign new_n4482 = ~new_n970 & new_n4481;
  assign new_n4483 = new_n4482 ^ new_n1509;
  assign new_n4484 = new_n812 ^ n36;
  assign new_n4485 = ~new_n978 & new_n4484;
  assign new_n4486 = new_n4485 ^ new_n1513;
  assign new_n4487 = new_n821 ^ n37;
  assign new_n4488 = ~new_n986 & new_n4487;
  assign new_n4489 = new_n4488 ^ new_n1517;
  assign new_n4490 = new_n830 ^ n38;
  assign new_n4491 = ~new_n994 & new_n4490;
  assign new_n4492 = new_n4491 ^ new_n1521;
  assign new_n4493 = new_n839 ^ n39;
  assign new_n4494 = ~new_n1002 & new_n4493;
  assign new_n4495 = new_n4494 ^ new_n1525;
  assign new_n4496 = new_n848 ^ n40;
  assign new_n4497 = ~new_n1010 & new_n4496;
  assign new_n4498 = new_n4497 ^ new_n1529;
  assign new_n4499 = new_n857 ^ n41;
  assign new_n4500 = ~new_n1018 & new_n4499;
  assign new_n4501 = new_n4500 ^ new_n1533;
  assign new_n4502 = new_n866 ^ n42;
  assign new_n4503 = ~new_n1026 & new_n4502;
  assign new_n4504 = new_n4503 ^ new_n1537;
  assign new_n4505 = new_n875 ^ n43;
  assign new_n4506 = ~new_n1034 & new_n4505;
  assign new_n4507 = new_n4506 ^ new_n1541;
  assign new_n4508 = new_n884 ^ n44;
  assign new_n4509 = ~new_n1042 & new_n4508;
  assign new_n4510 = new_n4509 ^ new_n1545;
  assign new_n4511 = new_n893 ^ n45;
  assign new_n4512 = ~new_n1050 & new_n4511;
  assign new_n4513 = new_n4512 ^ new_n1549;
  assign new_n4514 = new_n902 ^ n46;
  assign new_n4515 = ~new_n1058 & new_n4514;
  assign new_n4516 = new_n4515 ^ new_n1553;
  assign new_n4517 = new_n911 ^ n47;
  assign new_n4518 = ~new_n1066 & new_n4517;
  assign new_n4519 = new_n4518 ^ new_n1557;
  assign new_n4520 = new_n920 ^ n48;
  assign new_n4521 = ~new_n1074 & new_n4520;
  assign new_n4522 = new_n4521 ^ new_n1561;
  assign new_n4523 = new_n929 ^ n49;
  assign new_n4524 = ~new_n1082 & new_n4523;
  assign new_n4525 = new_n4524 ^ new_n1565;
  assign new_n4526 = new_n938 ^ n50;
  assign new_n4527 = ~new_n1090 & new_n4526;
  assign new_n4528 = new_n4527 ^ new_n1569;
  assign new_n4529 = new_n947 ^ n51;
  assign new_n4530 = ~new_n1098 & new_n4529;
  assign new_n4531 = new_n4530 ^ new_n1573;
  assign new_n4532 = new_n956 ^ n52;
  assign new_n4533 = ~new_n1106 & new_n4532;
  assign new_n4534 = new_n4533 ^ new_n1577;
  assign new_n4535 = new_n965 ^ n53;
  assign new_n4536 = ~new_n1114 & new_n4535;
  assign new_n4537 = new_n4536 ^ new_n1581;
  assign new_n4538 = new_n974 ^ n54;
  assign new_n4539 = ~new_n1122 & new_n4538;
  assign new_n4540 = new_n4539 ^ new_n1585;
  assign new_n4541 = new_n982 ^ n55;
  assign new_n4542 = ~new_n1130 & new_n4541;
  assign new_n4543 = new_n4542 ^ new_n1589;
  assign new_n4544 = new_n990 ^ n56;
  assign new_n4545 = ~new_n1138 & new_n4544;
  assign new_n4546 = new_n4545 ^ new_n1593;
  assign new_n4547 = new_n998 ^ n57;
  assign new_n4548 = ~new_n1146 & new_n4547;
  assign new_n4549 = new_n4548 ^ new_n1597;
  assign new_n4550 = new_n1006 ^ n58;
  assign new_n4551 = ~new_n579 & new_n4550;
  assign new_n4552 = new_n4551 ^ new_n1601;
  assign new_n4553 = new_n1014 ^ n59;
  assign new_n4554 = ~new_n589 & new_n4553;
  assign new_n4555 = new_n4554 ^ new_n1605;
  assign new_n4556 = new_n1022 ^ n60;
  assign new_n4557 = ~new_n599 & new_n4556;
  assign new_n4558 = new_n4557 ^ new_n1609;
  assign new_n4559 = new_n1030 ^ n61;
  assign new_n4560 = ~new_n609 & new_n4559;
  assign new_n4561 = new_n4560 ^ new_n1613;
  assign new_n4562 = new_n1038 ^ n62;
  assign new_n4563 = ~new_n619 & new_n4562;
  assign new_n4564 = new_n4563 ^ new_n1617;
  assign new_n4565 = new_n1046 ^ n63;
  assign new_n4566 = ~new_n629 & new_n4565;
  assign new_n4567 = new_n4566 ^ new_n1621;
  assign new_n4568 = new_n1054 ^ n64;
  assign new_n4569 = ~new_n639 & new_n4568;
  assign new_n4570 = new_n4569 ^ new_n1625;
  assign new_n4571 = new_n1062 ^ n65;
  assign new_n4572 = ~new_n649 & new_n4571;
  assign new_n4573 = new_n4572 ^ new_n1629;
  assign new_n4574 = new_n1070 ^ n66;
  assign new_n4575 = ~new_n659 & new_n4574;
  assign new_n4576 = new_n4575 ^ new_n1633;
  assign new_n4577 = new_n1078 ^ n67;
  assign new_n4578 = ~new_n669 & new_n4577;
  assign new_n4579 = new_n4578 ^ new_n1637;
  assign new_n4580 = new_n1086 ^ n68;
  assign new_n4581 = ~new_n679 & new_n4580;
  assign new_n4582 = new_n4581 ^ new_n1641;
  assign new_n4583 = new_n1094 ^ n69;
  assign new_n4584 = ~new_n689 & new_n4583;
  assign new_n4585 = new_n4584 ^ new_n1645;
  assign new_n4586 = new_n1102 ^ n70;
  assign new_n4587 = ~new_n699 & new_n4586;
  assign new_n4588 = new_n4587 ^ new_n1649;
  assign new_n4589 = new_n1110 ^ n71;
  assign new_n4590 = ~new_n709 & new_n4589;
  assign new_n4591 = new_n4590 ^ new_n1653;
  assign new_n4592 = new_n1118 ^ n72;
  assign new_n4593 = ~new_n719 & new_n4592;
  assign new_n4594 = new_n4593 ^ new_n1657;
  assign new_n4595 = new_n1126 ^ n73;
  assign new_n4596 = ~new_n729 & new_n4595;
  assign new_n4597 = new_n4596 ^ new_n1661;
  assign new_n4598 = new_n1134 ^ n74;
  assign new_n4599 = ~new_n739 & new_n4598;
  assign new_n4600 = new_n4599 ^ new_n1409;
  assign new_n4601 = new_n1142 ^ n75;
  assign new_n4602 = ~new_n749 & new_n4601;
  assign new_n4603 = new_n4602 ^ new_n1413;
  assign new_n4604 = new_n1150 ^ n76;
  assign new_n4605 = ~new_n759 & new_n4604;
  assign new_n4606 = new_n4605 ^ new_n1417;
  assign new_n4607 = new_n584 ^ n77;
  assign new_n4608 = ~new_n769 & new_n4607;
  assign new_n4609 = new_n4608 ^ new_n1421;
  assign new_n4610 = new_n594 ^ n78;
  assign new_n4611 = ~new_n779 & new_n4610;
  assign new_n4612 = new_n4611 ^ new_n1425;
  assign new_n4613 = new_n604 ^ n79;
  assign new_n4614 = ~new_n789 & new_n4613;
  assign new_n4615 = new_n4614 ^ new_n1429;
  assign new_n4616 = new_n614 ^ n80;
  assign new_n4617 = ~new_n799 & new_n4616;
  assign new_n4618 = new_n4617 ^ new_n1433;
  assign new_n4619 = new_n624 ^ n81;
  assign new_n4620 = ~new_n808 & new_n4619;
  assign new_n4621 = new_n4620 ^ new_n1437;
  assign new_n4622 = new_n634 ^ n82;
  assign new_n4623 = ~new_n817 & new_n4622;
  assign new_n4624 = new_n4623 ^ new_n1441;
  assign new_n4625 = new_n644 ^ n83;
  assign new_n4626 = ~new_n826 & new_n4625;
  assign new_n4627 = new_n4626 ^ new_n1445;
  assign new_n4628 = new_n654 ^ n84;
  assign new_n4629 = ~new_n835 & new_n4628;
  assign new_n4630 = new_n4629 ^ new_n1449;
  assign new_n4631 = new_n664 ^ n85;
  assign new_n4632 = ~new_n844 & new_n4631;
  assign new_n4633 = new_n4632 ^ new_n1453;
  assign new_n4634 = new_n674 ^ n86;
  assign new_n4635 = ~new_n853 & new_n4634;
  assign new_n4636 = new_n4635 ^ new_n1457;
  assign new_n4637 = new_n684 ^ n87;
  assign new_n4638 = ~new_n862 & new_n4637;
  assign new_n4639 = new_n4638 ^ new_n1461;
  assign new_n4640 = new_n694 ^ n88;
  assign new_n4641 = ~new_n871 & new_n4640;
  assign new_n4642 = new_n4641 ^ new_n1465;
  assign new_n4643 = new_n704 ^ n89;
  assign new_n4644 = ~new_n880 & new_n4643;
  assign new_n4645 = new_n4644 ^ new_n1469;
  assign new_n4646 = new_n714 ^ n90;
  assign new_n4647 = ~new_n889 & new_n4646;
  assign new_n4648 = new_n4647 ^ new_n1473;
  assign new_n4649 = new_n724 ^ n91;
  assign new_n4650 = ~new_n898 & new_n4649;
  assign new_n4651 = new_n4650 ^ new_n1477;
  assign new_n4652 = new_n734 ^ n92;
  assign new_n4653 = ~new_n907 & new_n4652;
  assign new_n4654 = new_n4653 ^ new_n1481;
  assign new_n4655 = new_n744 ^ n93;
  assign new_n4656 = ~new_n916 & new_n4655;
  assign new_n4657 = new_n4656 ^ new_n1485;
  assign new_n4658 = new_n754 ^ n94;
  assign new_n4659 = ~new_n925 & new_n4658;
  assign new_n4660 = new_n4659 ^ new_n1489;
  assign new_n4661 = new_n764 ^ n95;
  assign new_n4662 = ~new_n934 & new_n4661;
  assign new_n4663 = new_n4662 ^ new_n1493;
  assign new_n4664 = new_n774 ^ n96;
  assign new_n4665 = ~new_n943 & new_n4664;
  assign new_n4666 = new_n4665 ^ new_n1497;
  assign new_n4667 = new_n784 ^ n33;
  assign new_n4668 = ~new_n952 & new_n4667;
  assign new_n4669 = new_n4668 ^ new_n1501;
  assign new_n4670 = new_n794 ^ n34;
  assign new_n4671 = ~new_n961 & new_n4670;
  assign new_n4672 = new_n4671 ^ new_n1505;
  assign new_n4673 = ~new_n4481 & new_n772;
  assign new_n4674 = new_n4673 ^ new_n970;
  assign new_n4675 = ~new_n4484 & new_n782;
  assign new_n4676 = new_n4675 ^ new_n978;
  assign new_n4677 = ~new_n4487 & new_n792;
  assign new_n4678 = new_n4677 ^ new_n986;
  assign new_n4679 = ~new_n4490 & new_n801;
  assign new_n4680 = new_n4679 ^ new_n994;
  assign new_n4681 = ~new_n4493 & new_n810;
  assign new_n4682 = new_n4681 ^ new_n1002;
  assign new_n4683 = ~new_n4496 & new_n819;
  assign new_n4684 = new_n4683 ^ new_n1010;
  assign new_n4685 = ~new_n4499 & new_n828;
  assign new_n4686 = new_n4685 ^ new_n1018;
  assign new_n4687 = ~new_n4502 & new_n837;
  assign new_n4688 = new_n4687 ^ new_n1026;
  assign new_n4689 = ~new_n4505 & new_n846;
  assign new_n4690 = new_n4689 ^ new_n1034;
  assign new_n4691 = ~new_n4508 & new_n855;
  assign new_n4692 = new_n4691 ^ new_n1042;
  assign new_n4693 = ~new_n4511 & new_n864;
  assign new_n4694 = new_n4693 ^ new_n1050;
  assign new_n4695 = ~new_n4514 & new_n873;
  assign new_n4696 = new_n4695 ^ new_n1058;
  assign new_n4697 = ~new_n4517 & new_n882;
  assign new_n4698 = new_n4697 ^ new_n1066;
  assign new_n4699 = ~new_n4520 & new_n891;
  assign new_n4700 = new_n4699 ^ new_n1074;
  assign new_n4701 = ~new_n4523 & new_n900;
  assign new_n4702 = new_n4701 ^ new_n1082;
  assign new_n4703 = ~new_n4526 & new_n909;
  assign new_n4704 = new_n4703 ^ new_n1090;
  assign new_n4705 = ~new_n4529 & new_n918;
  assign new_n4706 = new_n4705 ^ new_n1098;
  assign new_n4707 = ~new_n4532 & new_n927;
  assign new_n4708 = new_n4707 ^ new_n1106;
  assign new_n4709 = ~new_n4535 & new_n936;
  assign new_n4710 = new_n4709 ^ new_n1114;
  assign new_n4711 = ~new_n4538 & new_n945;
  assign new_n4712 = new_n4711 ^ new_n1122;
  assign new_n4713 = ~new_n4541 & new_n954;
  assign new_n4714 = new_n4713 ^ new_n1130;
  assign new_n4715 = ~new_n4544 & new_n963;
  assign new_n4716 = new_n4715 ^ new_n1138;
  assign new_n4717 = ~new_n4547 & new_n972;
  assign new_n4718 = new_n4717 ^ new_n1146;
  assign new_n4719 = ~new_n4550 & new_n980;
  assign new_n4720 = new_n4719 ^ new_n579;
  assign new_n4721 = ~new_n4553 & new_n988;
  assign new_n4722 = new_n4721 ^ new_n589;
  assign new_n4723 = ~new_n4556 & new_n996;
  assign new_n4724 = new_n4723 ^ new_n599;
  assign new_n4725 = ~new_n4559 & new_n1004;
  assign new_n4726 = new_n4725 ^ new_n609;
  assign new_n4727 = ~new_n4562 & new_n1012;
  assign new_n4728 = new_n4727 ^ new_n619;
  assign new_n4729 = ~new_n4565 & new_n1020;
  assign new_n4730 = new_n4729 ^ new_n629;
  assign new_n4731 = ~new_n4568 & new_n1028;
  assign new_n4732 = new_n4731 ^ new_n639;
  assign new_n4733 = ~new_n4571 & new_n1036;
  assign new_n4734 = new_n4733 ^ new_n649;
  assign new_n4735 = ~new_n4574 & new_n1044;
  assign new_n4736 = new_n4735 ^ new_n659;
  assign new_n4737 = ~new_n4577 & new_n1052;
  assign new_n4738 = new_n4737 ^ new_n669;
  assign new_n4739 = ~new_n4580 & new_n1060;
  assign new_n4740 = new_n4739 ^ new_n679;
  assign new_n4741 = ~new_n4583 & new_n1068;
  assign new_n4742 = new_n4741 ^ new_n689;
  assign new_n4743 = ~new_n4586 & new_n1076;
  assign new_n4744 = new_n4743 ^ new_n699;
  assign new_n4745 = ~new_n4589 & new_n1084;
  assign new_n4746 = new_n4745 ^ new_n709;
  assign new_n4747 = ~new_n4592 & new_n1092;
  assign new_n4748 = new_n4747 ^ new_n719;
  assign new_n4749 = ~new_n4595 & new_n1100;
  assign new_n4750 = new_n4749 ^ new_n729;
  assign new_n4751 = ~new_n4598 & new_n1108;
  assign new_n4752 = new_n4751 ^ new_n739;
  assign new_n4753 = ~new_n4601 & new_n1116;
  assign new_n4754 = new_n4753 ^ new_n749;
  assign new_n4755 = ~new_n4604 & new_n1124;
  assign new_n4756 = new_n4755 ^ new_n759;
  assign new_n4757 = ~new_n4607 & new_n1132;
  assign new_n4758 = new_n4757 ^ new_n769;
  assign new_n4759 = ~new_n4610 & new_n1140;
  assign new_n4760 = new_n4759 ^ new_n779;
  assign new_n4761 = ~new_n4613 & new_n1148;
  assign new_n4762 = new_n4761 ^ new_n789;
  assign new_n4763 = ~new_n4616 & new_n582;
  assign new_n4764 = new_n4763 ^ new_n799;
  assign new_n4765 = ~new_n4619 & new_n592;
  assign new_n4766 = new_n4765 ^ new_n808;
  assign new_n4767 = ~new_n4622 & new_n602;
  assign new_n4768 = new_n4767 ^ new_n817;
  assign new_n4769 = ~new_n4625 & new_n612;
  assign new_n4770 = new_n4769 ^ new_n826;
  assign new_n4771 = ~new_n4628 & new_n622;
  assign new_n4772 = new_n4771 ^ new_n835;
  assign new_n4773 = ~new_n4631 & new_n632;
  assign new_n4774 = new_n4773 ^ new_n844;
  assign new_n4775 = ~new_n4634 & new_n642;
  assign new_n4776 = new_n4775 ^ new_n853;
  assign new_n4777 = ~new_n4637 & new_n652;
  assign new_n4778 = new_n4777 ^ new_n862;
  assign new_n4779 = ~new_n4640 & new_n662;
  assign new_n4780 = new_n4779 ^ new_n871;
  assign new_n4781 = ~new_n4643 & new_n672;
  assign new_n4782 = new_n4781 ^ new_n880;
  assign new_n4783 = ~new_n4646 & new_n682;
  assign new_n4784 = new_n4783 ^ new_n889;
  assign new_n4785 = ~new_n4649 & new_n692;
  assign new_n4786 = new_n4785 ^ new_n898;
  assign new_n4787 = ~new_n4652 & new_n702;
  assign new_n4788 = new_n4787 ^ new_n907;
  assign new_n4789 = ~new_n4655 & new_n712;
  assign new_n4790 = new_n4789 ^ new_n916;
  assign new_n4791 = ~new_n4658 & new_n722;
  assign new_n4792 = new_n4791 ^ new_n925;
  assign new_n4793 = ~new_n4661 & new_n732;
  assign new_n4794 = new_n4793 ^ new_n934;
  assign new_n4795 = ~new_n4664 & new_n742;
  assign new_n4796 = new_n4795 ^ new_n943;
  assign new_n4797 = ~new_n4667 & new_n752;
  assign new_n4798 = new_n4797 ^ new_n952;
  assign new_n4799 = ~new_n4670 & new_n762;
  assign new_n4800 = new_n4799 ^ new_n961;
  assign new_n4801 = ~new_n772 & new_n1289;
  assign new_n4802 = new_n4801 ^ new_n4481;
  assign new_n4803 = ~new_n782 & new_n1293;
  assign new_n4804 = new_n4803 ^ new_n4484;
  assign new_n4805 = ~new_n792 & new_n1297;
  assign new_n4806 = new_n4805 ^ new_n4487;
  assign new_n4807 = ~new_n801 & new_n1301;
  assign new_n4808 = new_n4807 ^ new_n4490;
  assign new_n4809 = ~new_n810 & new_n1305;
  assign new_n4810 = new_n4809 ^ new_n4493;
  assign new_n4811 = ~new_n819 & new_n1309;
  assign new_n4812 = new_n4811 ^ new_n4496;
  assign new_n4813 = ~new_n828 & new_n1313;
  assign new_n4814 = new_n4813 ^ new_n4499;
  assign new_n4815 = ~new_n837 & new_n1317;
  assign new_n4816 = new_n4815 ^ new_n4502;
  assign new_n4817 = ~new_n846 & new_n1321;
  assign new_n4818 = new_n4817 ^ new_n4505;
  assign new_n4819 = ~new_n855 & new_n1325;
  assign new_n4820 = new_n4819 ^ new_n4508;
  assign new_n4821 = ~new_n864 & new_n1329;
  assign new_n4822 = new_n4821 ^ new_n4511;
  assign new_n4823 = ~new_n873 & new_n1333;
  assign new_n4824 = new_n4823 ^ new_n4514;
  assign new_n4825 = ~new_n882 & new_n1337;
  assign new_n4826 = new_n4825 ^ new_n4517;
  assign new_n4827 = ~new_n891 & new_n1341;
  assign new_n4828 = new_n4827 ^ new_n4520;
  assign new_n4829 = ~new_n900 & new_n1345;
  assign new_n4830 = new_n4829 ^ new_n4523;
  assign new_n4831 = ~new_n909 & new_n1349;
  assign new_n4832 = new_n4831 ^ new_n4526;
  assign new_n4833 = ~new_n918 & new_n1353;
  assign new_n4834 = new_n4833 ^ new_n4529;
  assign new_n4835 = ~new_n927 & new_n1357;
  assign new_n4836 = new_n4835 ^ new_n4532;
  assign new_n4837 = ~new_n936 & new_n1361;
  assign new_n4838 = new_n4837 ^ new_n4535;
  assign new_n4839 = ~new_n945 & new_n1365;
  assign new_n4840 = new_n4839 ^ new_n4538;
  assign new_n4841 = ~new_n954 & new_n1369;
  assign new_n4842 = new_n4841 ^ new_n4541;
  assign new_n4843 = ~new_n963 & new_n1373;
  assign new_n4844 = new_n4843 ^ new_n4544;
  assign new_n4845 = ~new_n972 & new_n1377;
  assign new_n4846 = new_n4845 ^ new_n4547;
  assign new_n4847 = ~new_n980 & new_n1381;
  assign new_n4848 = new_n4847 ^ new_n4550;
  assign new_n4849 = ~new_n988 & new_n1385;
  assign new_n4850 = new_n4849 ^ new_n4553;
  assign new_n4851 = ~new_n996 & new_n1389;
  assign new_n4852 = new_n4851 ^ new_n4556;
  assign new_n4853 = ~new_n1004 & new_n1393;
  assign new_n4854 = new_n4853 ^ new_n4559;
  assign new_n4855 = ~new_n1012 & new_n1397;
  assign new_n4856 = new_n4855 ^ new_n4562;
  assign new_n4857 = ~new_n1020 & new_n1401;
  assign new_n4858 = new_n4857 ^ new_n4565;
  assign new_n4859 = ~new_n1028 & new_n1405;
  assign new_n4860 = new_n4859 ^ new_n4568;
  assign new_n4861 = ~new_n1036 & new_n1153;
  assign new_n4862 = new_n4861 ^ new_n4571;
  assign new_n4863 = ~new_n1044 & new_n1157;
  assign new_n4864 = new_n4863 ^ new_n4574;
  assign new_n4865 = ~new_n1052 & new_n1161;
  assign new_n4866 = new_n4865 ^ new_n4577;
  assign new_n4867 = ~new_n1060 & new_n1165;
  assign new_n4868 = new_n4867 ^ new_n4580;
  assign new_n4869 = ~new_n1068 & new_n1169;
  assign new_n4870 = new_n4869 ^ new_n4583;
  assign new_n4871 = ~new_n1076 & new_n1173;
  assign new_n4872 = new_n4871 ^ new_n4586;
  assign new_n4873 = ~new_n1084 & new_n1177;
  assign new_n4874 = new_n4873 ^ new_n4589;
  assign new_n4875 = ~new_n1092 & new_n1181;
  assign new_n4876 = new_n4875 ^ new_n4592;
  assign new_n4877 = ~new_n1100 & new_n1185;
  assign new_n4878 = new_n4877 ^ new_n4595;
  assign new_n4879 = ~new_n1108 & new_n1189;
  assign new_n4880 = new_n4879 ^ new_n4598;
  assign new_n4881 = ~new_n1116 & new_n1193;
  assign new_n4882 = new_n4881 ^ new_n4601;
  assign new_n4883 = ~new_n1124 & new_n1197;
  assign new_n4884 = new_n4883 ^ new_n4604;
  assign new_n4885 = ~new_n1132 & new_n1201;
  assign new_n4886 = new_n4885 ^ new_n4607;
  assign new_n4887 = ~new_n1140 & new_n1205;
  assign new_n4888 = new_n4887 ^ new_n4610;
  assign new_n4889 = ~new_n1148 & new_n1209;
  assign new_n4890 = new_n4889 ^ new_n4613;
  assign new_n4891 = ~new_n582 & new_n1213;
  assign new_n4892 = new_n4891 ^ new_n4616;
  assign new_n4893 = ~new_n592 & new_n1217;
  assign new_n4894 = new_n4893 ^ new_n4619;
  assign new_n4895 = ~new_n602 & new_n1221;
  assign new_n4896 = new_n4895 ^ new_n4622;
  assign new_n4897 = ~new_n612 & new_n1225;
  assign new_n4898 = new_n4897 ^ new_n4625;
  assign new_n4899 = ~new_n622 & new_n1229;
  assign new_n4900 = new_n4899 ^ new_n4628;
  assign new_n4901 = ~new_n632 & new_n1233;
  assign new_n4902 = new_n4901 ^ new_n4631;
  assign new_n4903 = ~new_n642 & new_n1237;
  assign new_n4904 = new_n4903 ^ new_n4634;
  assign new_n4905 = ~new_n652 & new_n1241;
  assign new_n4906 = new_n4905 ^ new_n4637;
  assign new_n4907 = ~new_n662 & new_n1245;
  assign new_n4908 = new_n4907 ^ new_n4640;
  assign new_n4909 = ~new_n672 & new_n1249;
  assign new_n4910 = new_n4909 ^ new_n4643;
  assign new_n4911 = ~new_n682 & new_n1253;
  assign new_n4912 = new_n4911 ^ new_n4646;
  assign new_n4913 = ~new_n692 & new_n1257;
  assign new_n4914 = new_n4913 ^ new_n4649;
  assign new_n4915 = ~new_n702 & new_n1261;
  assign new_n4916 = new_n4915 ^ new_n4652;
  assign new_n4917 = ~new_n712 & new_n1265;
  assign new_n4918 = new_n4917 ^ new_n4655;
  assign new_n4919 = ~new_n722 & new_n1269;
  assign new_n4920 = new_n4919 ^ new_n4658;
  assign new_n4921 = ~new_n732 & new_n1273;
  assign new_n4922 = new_n4921 ^ new_n4661;
  assign new_n4923 = ~new_n742 & new_n1277;
  assign new_n4924 = new_n4923 ^ new_n4664;
  assign new_n4925 = ~new_n752 & new_n1281;
  assign new_n4926 = new_n4925 ^ new_n4667;
  assign new_n4927 = ~new_n762 & new_n1285;
  assign new_n4928 = new_n4927 ^ new_n4670;
  assign po0 = new_n586;
  assign po1 = new_n596;
  assign po2 = new_n606;
  assign po3 = new_n616;
  assign po4 = new_n626;
  assign po5 = new_n636;
  assign po6 = new_n646;
  assign po7 = new_n656;
  assign po8 = new_n666;
  assign po9 = new_n676;
  assign po10 = new_n686;
  assign po11 = new_n696;
  assign po12 = new_n706;
  assign po13 = new_n716;
  assign po14 = new_n726;
  assign po15 = new_n736;
  assign po16 = new_n746;
  assign po17 = new_n756;
  assign po18 = new_n766;
  assign po19 = new_n776;
  assign po20 = new_n786;
  assign po21 = new_n796;
  assign po22 = new_n805;
  assign po23 = new_n814;
  assign po24 = new_n823;
  assign po25 = new_n832;
  assign po26 = new_n841;
  assign po27 = new_n850;
  assign po28 = new_n859;
  assign po29 = new_n868;
  assign po30 = new_n877;
  assign po31 = new_n886;
  assign po32 = new_n895;
  assign po33 = new_n904;
  assign po34 = new_n913;
  assign po35 = new_n922;
  assign po36 = new_n931;
  assign po37 = new_n940;
  assign po38 = new_n949;
  assign po39 = new_n958;
  assign po40 = new_n967;
  assign po41 = new_n976;
  assign po42 = new_n984;
  assign po43 = new_n992;
  assign po44 = new_n1000;
  assign po45 = new_n1008;
  assign po46 = new_n1016;
  assign po47 = new_n1024;
  assign po48 = new_n1032;
  assign po49 = new_n1040;
  assign po50 = new_n1048;
  assign po51 = new_n1056;
  assign po52 = new_n1064;
  assign po53 = new_n1072;
  assign po54 = new_n1080;
  assign po55 = new_n1088;
  assign po56 = new_n1096;
  assign po57 = new_n1104;
  assign po58 = new_n1112;
  assign po59 = new_n1120;
  assign po60 = new_n1128;
  assign po61 = new_n1136;
  assign po62 = new_n1144;
  assign po63 = new_n1152;
  assign po64 = new_n1156;
  assign po65 = new_n1160;
  assign po66 = new_n1164;
  assign po67 = new_n1168;
  assign po68 = new_n1172;
  assign po69 = new_n1176;
  assign po70 = new_n1180;
  assign po71 = new_n1184;
  assign po72 = new_n1188;
  assign po73 = new_n1192;
  assign po74 = new_n1196;
  assign po75 = new_n1200;
  assign po76 = new_n1204;
  assign po77 = new_n1208;
  assign po78 = new_n1212;
  assign po79 = new_n1216;
  assign po80 = new_n1220;
  assign po81 = new_n1224;
  assign po82 = new_n1228;
  assign po83 = new_n1232;
  assign po84 = new_n1236;
  assign po85 = new_n1240;
  assign po86 = new_n1244;
  assign po87 = new_n1248;
  assign po88 = new_n1252;
  assign po89 = new_n1256;
  assign po90 = new_n1260;
  assign po91 = new_n1264;
  assign po92 = new_n1268;
  assign po93 = new_n1272;
  assign po94 = new_n1276;
  assign po95 = new_n1280;
  assign po96 = new_n1284;
  assign po97 = new_n1288;
  assign po98 = new_n1292;
  assign po99 = new_n1296;
  assign po100 = new_n1300;
  assign po101 = new_n1304;
  assign po102 = new_n1308;
  assign po103 = new_n1312;
  assign po104 = new_n1316;
  assign po105 = new_n1320;
  assign po106 = new_n1324;
  assign po107 = new_n1328;
  assign po108 = new_n1332;
  assign po109 = new_n1336;
  assign po110 = new_n1340;
  assign po111 = new_n1344;
  assign po112 = new_n1348;
  assign po113 = new_n1352;
  assign po114 = new_n1356;
  assign po115 = new_n1360;
  assign po116 = new_n1364;
  assign po117 = new_n1368;
  assign po118 = new_n1372;
  assign po119 = new_n1376;
  assign po120 = new_n1380;
  assign po121 = new_n1384;
  assign po122 = new_n1388;
  assign po123 = new_n1392;
  assign po124 = new_n1396;
  assign po125 = new_n1400;
  assign po126 = new_n1404;
  assign po127 = new_n1408;
  assign po128 = new_n1412;
  assign po129 = new_n1416;
  assign po130 = new_n1420;
  assign po131 = new_n1424;
  assign po132 = new_n1428;
  assign po133 = new_n1432;
  assign po134 = new_n1436;
  assign po135 = new_n1440;
  assign po136 = new_n1444;
  assign po137 = new_n1448;
  assign po138 = new_n1452;
  assign po139 = new_n1456;
  assign po140 = new_n1460;
  assign po141 = new_n1464;
  assign po142 = new_n1468;
  assign po143 = new_n1472;
  assign po144 = new_n1476;
  assign po145 = new_n1480;
  assign po146 = new_n1484;
  assign po147 = new_n1488;
  assign po148 = new_n1492;
  assign po149 = new_n1496;
  assign po150 = new_n1500;
  assign po151 = new_n1504;
  assign po152 = new_n1508;
  assign po153 = new_n1512;
  assign po154 = new_n1516;
  assign po155 = new_n1520;
  assign po156 = new_n1524;
  assign po157 = new_n1528;
  assign po158 = new_n1532;
  assign po159 = new_n1536;
  assign po160 = new_n1540;
  assign po161 = new_n1544;
  assign po162 = new_n1548;
  assign po163 = new_n1552;
  assign po164 = new_n1556;
  assign po165 = new_n1560;
  assign po166 = new_n1564;
  assign po167 = new_n1568;
  assign po168 = new_n1572;
  assign po169 = new_n1576;
  assign po170 = new_n1580;
  assign po171 = new_n1584;
  assign po172 = new_n1588;
  assign po173 = new_n1592;
  assign po174 = new_n1596;
  assign po175 = new_n1600;
  assign po176 = new_n1604;
  assign po177 = new_n1608;
  assign po178 = new_n1612;
  assign po179 = new_n1616;
  assign po180 = new_n1620;
  assign po181 = new_n1624;
  assign po182 = new_n1628;
  assign po183 = new_n1632;
  assign po184 = new_n1636;
  assign po185 = new_n1640;
  assign po186 = new_n1644;
  assign po187 = new_n1648;
  assign po188 = new_n1652;
  assign po189 = new_n1656;
  assign po190 = new_n1660;
  assign po191 = new_n1664;
  assign po192 = new_n1666;
  assign po193 = new_n1668;
  assign po194 = new_n1670;
  assign po195 = new_n1672;
  assign po196 = new_n1674;
  assign po197 = new_n1676;
  assign po198 = new_n1678;
  assign po199 = new_n1680;
  assign po200 = new_n1682;
  assign po201 = new_n1684;
  assign po202 = new_n1686;
  assign po203 = new_n1688;
  assign po204 = new_n1690;
  assign po205 = new_n1692;
  assign po206 = new_n1694;
  assign po207 = new_n1696;
  assign po208 = new_n1698;
  assign po209 = new_n1700;
  assign po210 = new_n1702;
  assign po211 = new_n1704;
  assign po212 = new_n1706;
  assign po213 = new_n1708;
  assign po214 = new_n1710;
  assign po215 = new_n1712;
  assign po216 = new_n1714;
  assign po217 = new_n1716;
  assign po218 = new_n1718;
  assign po219 = new_n1720;
  assign po220 = new_n1722;
  assign po221 = new_n1724;
  assign po222 = new_n1726;
  assign po223 = new_n1728;
  assign po224 = new_n1730;
  assign po225 = new_n1732;
  assign po226 = new_n1734;
  assign po227 = new_n1736;
  assign po228 = new_n1738;
  assign po229 = new_n1740;
  assign po230 = new_n1742;
  assign po231 = new_n1744;
  assign po232 = new_n1746;
  assign po233 = new_n1748;
  assign po234 = new_n1750;
  assign po235 = new_n1752;
  assign po236 = new_n1754;
  assign po237 = new_n1756;
  assign po238 = new_n1758;
  assign po239 = new_n1760;
  assign po240 = new_n1762;
  assign po241 = new_n1764;
  assign po242 = new_n1766;
  assign po243 = new_n1768;
  assign po244 = new_n1770;
  assign po245 = new_n1772;
  assign po246 = new_n1774;
  assign po247 = new_n1776;
  assign po248 = new_n1778;
  assign po249 = new_n1780;
  assign po250 = new_n1782;
  assign po251 = new_n1784;
  assign po252 = new_n1786;
  assign po253 = new_n1788;
  assign po254 = new_n1790;
  assign po255 = new_n1792;
  assign po256 = new_n1794;
  assign po257 = new_n1796;
  assign po258 = new_n1798;
  assign po259 = new_n1800;
  assign po260 = new_n1802;
  assign po261 = new_n1804;
  assign po262 = new_n1806;
  assign po263 = new_n1808;
  assign po264 = new_n1810;
  assign po265 = new_n1812;
  assign po266 = new_n1814;
  assign po267 = new_n1816;
  assign po268 = new_n1818;
  assign po269 = new_n1820;
  assign po270 = new_n1822;
  assign po271 = new_n1824;
  assign po272 = new_n1826;
  assign po273 = new_n1828;
  assign po274 = new_n1830;
  assign po275 = new_n1832;
  assign po276 = new_n1834;
  assign po277 = new_n1836;
  assign po278 = new_n1838;
  assign po279 = new_n1840;
  assign po280 = new_n1842;
  assign po281 = new_n1844;
  assign po282 = new_n1846;
  assign po283 = new_n1848;
  assign po284 = new_n1850;
  assign po285 = new_n1852;
  assign po286 = new_n1854;
  assign po287 = new_n1856;
  assign po288 = new_n1858;
  assign po289 = new_n1860;
  assign po290 = new_n1862;
  assign po291 = new_n1864;
  assign po292 = new_n1866;
  assign po293 = new_n1868;
  assign po294 = new_n1870;
  assign po295 = new_n1872;
  assign po296 = new_n1874;
  assign po297 = new_n1876;
  assign po298 = new_n1878;
  assign po299 = new_n1880;
  assign po300 = new_n1882;
  assign po301 = new_n1884;
  assign po302 = new_n1886;
  assign po303 = new_n1888;
  assign po304 = new_n1890;
  assign po305 = new_n1892;
  assign po306 = new_n1894;
  assign po307 = new_n1896;
  assign po308 = new_n1898;
  assign po309 = new_n1900;
  assign po310 = new_n1902;
  assign po311 = new_n1904;
  assign po312 = new_n1906;
  assign po313 = new_n1908;
  assign po314 = new_n1910;
  assign po315 = new_n1912;
  assign po316 = new_n1914;
  assign po317 = new_n1916;
  assign po318 = new_n1918;
  assign po319 = new_n1920;
  assign po320 = new_n1922;
  assign po321 = new_n1924;
  assign po322 = new_n1926;
  assign po323 = new_n1928;
  assign po324 = new_n1930;
  assign po325 = new_n1932;
  assign po326 = new_n1934;
  assign po327 = new_n1936;
  assign po328 = new_n1938;
  assign po329 = new_n1940;
  assign po330 = new_n1942;
  assign po331 = new_n1944;
  assign po332 = new_n1946;
  assign po333 = new_n1948;
  assign po334 = new_n1950;
  assign po335 = new_n1952;
  assign po336 = new_n1954;
  assign po337 = new_n1956;
  assign po338 = new_n1958;
  assign po339 = new_n1960;
  assign po340 = new_n1962;
  assign po341 = new_n1964;
  assign po342 = new_n1966;
  assign po343 = new_n1968;
  assign po344 = new_n1970;
  assign po345 = new_n1972;
  assign po346 = new_n1974;
  assign po347 = new_n1976;
  assign po348 = new_n1978;
  assign po349 = new_n1980;
  assign po350 = new_n1982;
  assign po351 = new_n1984;
  assign po352 = new_n1986;
  assign po353 = new_n1988;
  assign po354 = new_n1990;
  assign po355 = new_n1992;
  assign po356 = new_n1994;
  assign po357 = new_n1996;
  assign po358 = new_n1998;
  assign po359 = new_n2000;
  assign po360 = new_n2002;
  assign po361 = new_n2004;
  assign po362 = new_n2006;
  assign po363 = new_n2008;
  assign po364 = new_n2010;
  assign po365 = new_n2012;
  assign po366 = new_n2014;
  assign po367 = new_n2016;
  assign po368 = new_n2018;
  assign po369 = new_n2020;
  assign po370 = new_n2022;
  assign po371 = new_n2024;
  assign po372 = new_n2026;
  assign po373 = new_n2028;
  assign po374 = new_n2030;
  assign po375 = new_n2032;
  assign po376 = new_n2034;
  assign po377 = new_n2036;
  assign po378 = new_n2038;
  assign po379 = new_n2040;
  assign po380 = new_n2042;
  assign po381 = new_n2044;
  assign po382 = new_n2046;
  assign po383 = new_n2048;
  assign po384 = new_n2051;
  assign po385 = new_n2054;
  assign po386 = new_n2057;
  assign po387 = new_n2060;
  assign po388 = new_n2063;
  assign po389 = new_n2066;
  assign po390 = new_n2069;
  assign po391 = new_n2072;
  assign po392 = new_n2075;
  assign po393 = new_n2078;
  assign po394 = new_n2081;
  assign po395 = new_n2084;
  assign po396 = new_n2087;
  assign po397 = new_n2090;
  assign po398 = new_n2093;
  assign po399 = new_n2096;
  assign po400 = new_n2099;
  assign po401 = new_n2102;
  assign po402 = new_n2105;
  assign po403 = new_n2108;
  assign po404 = new_n2111;
  assign po405 = new_n2114;
  assign po406 = new_n2117;
  assign po407 = new_n2120;
  assign po408 = new_n2123;
  assign po409 = new_n2126;
  assign po410 = new_n2129;
  assign po411 = new_n2132;
  assign po412 = new_n2135;
  assign po413 = new_n2138;
  assign po414 = new_n2141;
  assign po415 = new_n2144;
  assign po416 = new_n2147;
  assign po417 = new_n2150;
  assign po418 = new_n2153;
  assign po419 = new_n2156;
  assign po420 = new_n2159;
  assign po421 = new_n2162;
  assign po422 = new_n2165;
  assign po423 = new_n2168;
  assign po424 = new_n2171;
  assign po425 = new_n2174;
  assign po426 = new_n2177;
  assign po427 = new_n2180;
  assign po428 = new_n2183;
  assign po429 = new_n2186;
  assign po430 = new_n2189;
  assign po431 = new_n2192;
  assign po432 = new_n2195;
  assign po433 = new_n2198;
  assign po434 = new_n2201;
  assign po435 = new_n2204;
  assign po436 = new_n2207;
  assign po437 = new_n2210;
  assign po438 = new_n2213;
  assign po439 = new_n2216;
  assign po440 = new_n2219;
  assign po441 = new_n2222;
  assign po442 = new_n2225;
  assign po443 = new_n2228;
  assign po444 = new_n2231;
  assign po445 = new_n2234;
  assign po446 = new_n2237;
  assign po447 = new_n2240;
  assign po448 = new_n2243;
  assign po449 = new_n2246;
  assign po450 = new_n2249;
  assign po451 = new_n2252;
  assign po452 = new_n2255;
  assign po453 = new_n2258;
  assign po454 = new_n2261;
  assign po455 = new_n2264;
  assign po456 = new_n2267;
  assign po457 = new_n2270;
  assign po458 = new_n2273;
  assign po459 = new_n2276;
  assign po460 = new_n2279;
  assign po461 = new_n2282;
  assign po462 = new_n2285;
  assign po463 = new_n2288;
  assign po464 = new_n2291;
  assign po465 = new_n2294;
  assign po466 = new_n2297;
  assign po467 = new_n2300;
  assign po468 = new_n2303;
  assign po469 = new_n2306;
  assign po470 = new_n2309;
  assign po471 = new_n2312;
  assign po472 = new_n2315;
  assign po473 = new_n2318;
  assign po474 = new_n2321;
  assign po475 = new_n2324;
  assign po476 = new_n2327;
  assign po477 = new_n2330;
  assign po478 = new_n2333;
  assign po479 = new_n2336;
  assign po480 = new_n2339;
  assign po481 = new_n2342;
  assign po482 = new_n2345;
  assign po483 = new_n2348;
  assign po484 = new_n2351;
  assign po485 = new_n2354;
  assign po486 = new_n2357;
  assign po487 = new_n2360;
  assign po488 = new_n2363;
  assign po489 = new_n2366;
  assign po490 = new_n2369;
  assign po491 = new_n2372;
  assign po492 = new_n2375;
  assign po493 = new_n2378;
  assign po494 = new_n2381;
  assign po495 = new_n2384;
  assign po496 = new_n2387;
  assign po497 = new_n2390;
  assign po498 = new_n2393;
  assign po499 = new_n2396;
  assign po500 = new_n2399;
  assign po501 = new_n2402;
  assign po502 = new_n2405;
  assign po503 = new_n2408;
  assign po504 = new_n2411;
  assign po505 = new_n2414;
  assign po506 = new_n2417;
  assign po507 = new_n2420;
  assign po508 = new_n2423;
  assign po509 = new_n2426;
  assign po510 = new_n2429;
  assign po511 = new_n2432;
  assign po512 = new_n2434;
  assign po513 = new_n2436;
  assign po514 = new_n2438;
  assign po515 = new_n2440;
  assign po516 = new_n2442;
  assign po517 = new_n2444;
  assign po518 = new_n2446;
  assign po519 = new_n2448;
  assign po520 = new_n2450;
  assign po521 = new_n2452;
  assign po522 = new_n2454;
  assign po523 = new_n2456;
  assign po524 = new_n2458;
  assign po525 = new_n2460;
  assign po526 = new_n2462;
  assign po527 = new_n2464;
  assign po528 = new_n2466;
  assign po529 = new_n2468;
  assign po530 = new_n2470;
  assign po531 = new_n2472;
  assign po532 = new_n2474;
  assign po533 = new_n2476;
  assign po534 = new_n2478;
  assign po535 = new_n2480;
  assign po536 = new_n2482;
  assign po537 = new_n2484;
  assign po538 = new_n2486;
  assign po539 = new_n2488;
  assign po540 = new_n2490;
  assign po541 = new_n2492;
  assign po542 = new_n2494;
  assign po543 = new_n2496;
  assign po544 = new_n2498;
  assign po545 = new_n2500;
  assign po546 = new_n2502;
  assign po547 = new_n2504;
  assign po548 = new_n2506;
  assign po549 = new_n2508;
  assign po550 = new_n2510;
  assign po551 = new_n2512;
  assign po552 = new_n2514;
  assign po553 = new_n2516;
  assign po554 = new_n2518;
  assign po555 = new_n2520;
  assign po556 = new_n2522;
  assign po557 = new_n2524;
  assign po558 = new_n2526;
  assign po559 = new_n2528;
  assign po560 = new_n2530;
  assign po561 = new_n2532;
  assign po562 = new_n2534;
  assign po563 = new_n2536;
  assign po564 = new_n2538;
  assign po565 = new_n2540;
  assign po566 = new_n2542;
  assign po567 = new_n2544;
  assign po568 = new_n2546;
  assign po569 = new_n2548;
  assign po570 = new_n2550;
  assign po571 = new_n2552;
  assign po572 = new_n2554;
  assign po573 = new_n2556;
  assign po574 = new_n2558;
  assign po575 = new_n2560;
  assign po576 = new_n2562;
  assign po577 = new_n2564;
  assign po578 = new_n2566;
  assign po579 = new_n2568;
  assign po580 = new_n2570;
  assign po581 = new_n2572;
  assign po582 = new_n2574;
  assign po583 = new_n2576;
  assign po584 = new_n2578;
  assign po585 = new_n2580;
  assign po586 = new_n2582;
  assign po587 = new_n2584;
  assign po588 = new_n2586;
  assign po589 = new_n2588;
  assign po590 = new_n2590;
  assign po591 = new_n2592;
  assign po592 = new_n2594;
  assign po593 = new_n2596;
  assign po594 = new_n2598;
  assign po595 = new_n2600;
  assign po596 = new_n2602;
  assign po597 = new_n2604;
  assign po598 = new_n2606;
  assign po599 = new_n2608;
  assign po600 = new_n2610;
  assign po601 = new_n2612;
  assign po602 = new_n2614;
  assign po603 = new_n2616;
  assign po604 = new_n2618;
  assign po605 = new_n2620;
  assign po606 = new_n2622;
  assign po607 = new_n2624;
  assign po608 = new_n2626;
  assign po609 = new_n2628;
  assign po610 = new_n2630;
  assign po611 = new_n2632;
  assign po612 = new_n2634;
  assign po613 = new_n2636;
  assign po614 = new_n2638;
  assign po615 = new_n2640;
  assign po616 = new_n2642;
  assign po617 = new_n2644;
  assign po618 = new_n2646;
  assign po619 = new_n2648;
  assign po620 = new_n2650;
  assign po621 = new_n2652;
  assign po622 = new_n2654;
  assign po623 = new_n2656;
  assign po624 = new_n2658;
  assign po625 = new_n2660;
  assign po626 = new_n2662;
  assign po627 = new_n2664;
  assign po628 = new_n2666;
  assign po629 = new_n2668;
  assign po630 = new_n2670;
  assign po631 = new_n2672;
  assign po632 = new_n2674;
  assign po633 = new_n2676;
  assign po634 = new_n2678;
  assign po635 = new_n2680;
  assign po636 = new_n2682;
  assign po637 = new_n2684;
  assign po638 = new_n2686;
  assign po639 = new_n2688;
  assign po640 = new_n2690;
  assign po641 = new_n2692;
  assign po642 = new_n2694;
  assign po643 = new_n2696;
  assign po644 = new_n2698;
  assign po645 = new_n2700;
  assign po646 = new_n2702;
  assign po647 = new_n2704;
  assign po648 = new_n2706;
  assign po649 = new_n2708;
  assign po650 = new_n2710;
  assign po651 = new_n2712;
  assign po652 = new_n2714;
  assign po653 = new_n2716;
  assign po654 = new_n2718;
  assign po655 = new_n2720;
  assign po656 = new_n2722;
  assign po657 = new_n2724;
  assign po658 = new_n2726;
  assign po659 = new_n2728;
  assign po660 = new_n2730;
  assign po661 = new_n2732;
  assign po662 = new_n2734;
  assign po663 = new_n2736;
  assign po664 = new_n2738;
  assign po665 = new_n2740;
  assign po666 = new_n2742;
  assign po667 = new_n2744;
  assign po668 = new_n2746;
  assign po669 = new_n2748;
  assign po670 = new_n2750;
  assign po671 = new_n2752;
  assign po672 = new_n2754;
  assign po673 = new_n2756;
  assign po674 = new_n2758;
  assign po675 = new_n2760;
  assign po676 = new_n2762;
  assign po677 = new_n2764;
  assign po678 = new_n2766;
  assign po679 = new_n2768;
  assign po680 = new_n2770;
  assign po681 = new_n2772;
  assign po682 = new_n2774;
  assign po683 = new_n2776;
  assign po684 = new_n2778;
  assign po685 = new_n2780;
  assign po686 = new_n2782;
  assign po687 = new_n2784;
  assign po688 = new_n2786;
  assign po689 = new_n2788;
  assign po690 = new_n2790;
  assign po691 = new_n2792;
  assign po692 = new_n2794;
  assign po693 = new_n2796;
  assign po694 = new_n2798;
  assign po695 = new_n2800;
  assign po696 = new_n2802;
  assign po697 = new_n2804;
  assign po698 = new_n2806;
  assign po699 = new_n2808;
  assign po700 = new_n2810;
  assign po701 = new_n2812;
  assign po702 = new_n2814;
  assign po703 = new_n2816;
  assign po704 = new_n2819;
  assign po705 = new_n2822;
  assign po706 = new_n2825;
  assign po707 = new_n2828;
  assign po708 = new_n2831;
  assign po709 = new_n2834;
  assign po710 = new_n2837;
  assign po711 = new_n2840;
  assign po712 = new_n2843;
  assign po713 = new_n2846;
  assign po714 = new_n2849;
  assign po715 = new_n2852;
  assign po716 = new_n2855;
  assign po717 = new_n2858;
  assign po718 = new_n2861;
  assign po719 = new_n2864;
  assign po720 = new_n2867;
  assign po721 = new_n2870;
  assign po722 = new_n2873;
  assign po723 = new_n2876;
  assign po724 = new_n2879;
  assign po725 = new_n2882;
  assign po726 = new_n2885;
  assign po727 = new_n2888;
  assign po728 = new_n2891;
  assign po729 = new_n2894;
  assign po730 = new_n2897;
  assign po731 = new_n2900;
  assign po732 = new_n2903;
  assign po733 = new_n2906;
  assign po734 = new_n2909;
  assign po735 = new_n2912;
  assign po736 = new_n2915;
  assign po737 = new_n2918;
  assign po738 = new_n2921;
  assign po739 = new_n2924;
  assign po740 = new_n2927;
  assign po741 = new_n2930;
  assign po742 = new_n2933;
  assign po743 = new_n2936;
  assign po744 = new_n2939;
  assign po745 = new_n2942;
  assign po746 = new_n2945;
  assign po747 = new_n2948;
  assign po748 = new_n2951;
  assign po749 = new_n2954;
  assign po750 = new_n2957;
  assign po751 = new_n2960;
  assign po752 = new_n2963;
  assign po753 = new_n2966;
  assign po754 = new_n2969;
  assign po755 = new_n2972;
  assign po756 = new_n2975;
  assign po757 = new_n2978;
  assign po758 = new_n2981;
  assign po759 = new_n2984;
  assign po760 = new_n2987;
  assign po761 = new_n2990;
  assign po762 = new_n2993;
  assign po763 = new_n2996;
  assign po764 = new_n2999;
  assign po765 = new_n3002;
  assign po766 = new_n3005;
  assign po767 = new_n3008;
  assign po768 = new_n3011;
  assign po769 = new_n3014;
  assign po770 = new_n3017;
  assign po771 = new_n3020;
  assign po772 = new_n3023;
  assign po773 = new_n3026;
  assign po774 = new_n3029;
  assign po775 = new_n3032;
  assign po776 = new_n3035;
  assign po777 = new_n3038;
  assign po778 = new_n3041;
  assign po779 = new_n3044;
  assign po780 = new_n3047;
  assign po781 = new_n3050;
  assign po782 = new_n3053;
  assign po783 = new_n3056;
  assign po784 = new_n3059;
  assign po785 = new_n3062;
  assign po786 = new_n3065;
  assign po787 = new_n3068;
  assign po788 = new_n3071;
  assign po789 = new_n3074;
  assign po790 = new_n3077;
  assign po791 = new_n3080;
  assign po792 = new_n3083;
  assign po793 = new_n3086;
  assign po794 = new_n3089;
  assign po795 = new_n3092;
  assign po796 = new_n3095;
  assign po797 = new_n3098;
  assign po798 = new_n3101;
  assign po799 = new_n3104;
  assign po800 = new_n3107;
  assign po801 = new_n3110;
  assign po802 = new_n3113;
  assign po803 = new_n3116;
  assign po804 = new_n3119;
  assign po805 = new_n3122;
  assign po806 = new_n3125;
  assign po807 = new_n3128;
  assign po808 = new_n3131;
  assign po809 = new_n3134;
  assign po810 = new_n3137;
  assign po811 = new_n3140;
  assign po812 = new_n3143;
  assign po813 = new_n3146;
  assign po814 = new_n3149;
  assign po815 = new_n3152;
  assign po816 = new_n3155;
  assign po817 = new_n3158;
  assign po818 = new_n3161;
  assign po819 = new_n3164;
  assign po820 = new_n3167;
  assign po821 = new_n3170;
  assign po822 = new_n3173;
  assign po823 = new_n3176;
  assign po824 = new_n3179;
  assign po825 = new_n3182;
  assign po826 = new_n3185;
  assign po827 = new_n3188;
  assign po828 = new_n3191;
  assign po829 = new_n3194;
  assign po830 = new_n3197;
  assign po831 = new_n3200;
  assign po832 = new_n3202;
  assign po833 = new_n3204;
  assign po834 = new_n3206;
  assign po835 = new_n3208;
  assign po836 = new_n3210;
  assign po837 = new_n3212;
  assign po838 = new_n3214;
  assign po839 = new_n3216;
  assign po840 = new_n3218;
  assign po841 = new_n3220;
  assign po842 = new_n3222;
  assign po843 = new_n3224;
  assign po844 = new_n3226;
  assign po845 = new_n3228;
  assign po846 = new_n3230;
  assign po847 = new_n3232;
  assign po848 = new_n3234;
  assign po849 = new_n3236;
  assign po850 = new_n3238;
  assign po851 = new_n3240;
  assign po852 = new_n3242;
  assign po853 = new_n3244;
  assign po854 = new_n3246;
  assign po855 = new_n3248;
  assign po856 = new_n3250;
  assign po857 = new_n3252;
  assign po858 = new_n3254;
  assign po859 = new_n3256;
  assign po860 = new_n3258;
  assign po861 = new_n3260;
  assign po862 = new_n3262;
  assign po863 = new_n3264;
  assign po864 = new_n3266;
  assign po865 = new_n3268;
  assign po866 = new_n3270;
  assign po867 = new_n3272;
  assign po868 = new_n3274;
  assign po869 = new_n3276;
  assign po870 = new_n3278;
  assign po871 = new_n3280;
  assign po872 = new_n3282;
  assign po873 = new_n3284;
  assign po874 = new_n3286;
  assign po875 = new_n3288;
  assign po876 = new_n3290;
  assign po877 = new_n3292;
  assign po878 = new_n3294;
  assign po879 = new_n3296;
  assign po880 = new_n3298;
  assign po881 = new_n3300;
  assign po882 = new_n3302;
  assign po883 = new_n3304;
  assign po884 = new_n3306;
  assign po885 = new_n3308;
  assign po886 = new_n3310;
  assign po887 = new_n3312;
  assign po888 = new_n3314;
  assign po889 = new_n3316;
  assign po890 = new_n3318;
  assign po891 = new_n3320;
  assign po892 = new_n3322;
  assign po893 = new_n3324;
  assign po894 = new_n3326;
  assign po895 = new_n3328;
  assign po896 = new_n3330;
  assign po897 = new_n3332;
  assign po898 = new_n3334;
  assign po899 = new_n3336;
  assign po900 = new_n3338;
  assign po901 = new_n3340;
  assign po902 = new_n3342;
  assign po903 = new_n3344;
  assign po904 = new_n3346;
  assign po905 = new_n3348;
  assign po906 = new_n3350;
  assign po907 = new_n3352;
  assign po908 = new_n3354;
  assign po909 = new_n3356;
  assign po910 = new_n3358;
  assign po911 = new_n3360;
  assign po912 = new_n3362;
  assign po913 = new_n3364;
  assign po914 = new_n3366;
  assign po915 = new_n3368;
  assign po916 = new_n3370;
  assign po917 = new_n3372;
  assign po918 = new_n3374;
  assign po919 = new_n3376;
  assign po920 = new_n3378;
  assign po921 = new_n3380;
  assign po922 = new_n3382;
  assign po923 = new_n3384;
  assign po924 = new_n3386;
  assign po925 = new_n3388;
  assign po926 = new_n3390;
  assign po927 = new_n3392;
  assign po928 = new_n3394;
  assign po929 = new_n3396;
  assign po930 = new_n3398;
  assign po931 = new_n3400;
  assign po932 = new_n3402;
  assign po933 = new_n3404;
  assign po934 = new_n3406;
  assign po935 = new_n3408;
  assign po936 = new_n3410;
  assign po937 = new_n3412;
  assign po938 = new_n3414;
  assign po939 = new_n3416;
  assign po940 = new_n3418;
  assign po941 = new_n3420;
  assign po942 = new_n3422;
  assign po943 = new_n3424;
  assign po944 = new_n3426;
  assign po945 = new_n3428;
  assign po946 = new_n3430;
  assign po947 = new_n3432;
  assign po948 = new_n3434;
  assign po949 = new_n3436;
  assign po950 = new_n3438;
  assign po951 = new_n3440;
  assign po952 = new_n3442;
  assign po953 = new_n3444;
  assign po954 = new_n3446;
  assign po955 = new_n3448;
  assign po956 = new_n3450;
  assign po957 = new_n3452;
  assign po958 = new_n3454;
  assign po959 = new_n3456;
  assign po960 = new_n3458;
  assign po961 = new_n3460;
  assign po962 = new_n3462;
  assign po963 = new_n3464;
  assign po964 = new_n3466;
  assign po965 = new_n3468;
  assign po966 = new_n3470;
  assign po967 = new_n3472;
  assign po968 = new_n3474;
  assign po969 = new_n3476;
  assign po970 = new_n3478;
  assign po971 = new_n3480;
  assign po972 = new_n3482;
  assign po973 = new_n3484;
  assign po974 = new_n3486;
  assign po975 = new_n3488;
  assign po976 = new_n3490;
  assign po977 = new_n3492;
  assign po978 = new_n3494;
  assign po979 = new_n3496;
  assign po980 = new_n3498;
  assign po981 = new_n3500;
  assign po982 = new_n3502;
  assign po983 = new_n3504;
  assign po984 = new_n3506;
  assign po985 = new_n3508;
  assign po986 = new_n3510;
  assign po987 = new_n3512;
  assign po988 = new_n3514;
  assign po989 = new_n3516;
  assign po990 = new_n3518;
  assign po991 = new_n3520;
  assign po992 = new_n3522;
  assign po993 = new_n3524;
  assign po994 = new_n3526;
  assign po995 = new_n3528;
  assign po996 = new_n3530;
  assign po997 = new_n3532;
  assign po998 = new_n3534;
  assign po999 = new_n3536;
  assign po1000 = new_n3538;
  assign po1001 = new_n3540;
  assign po1002 = new_n3542;
  assign po1003 = new_n3544;
  assign po1004 = new_n3546;
  assign po1005 = new_n3548;
  assign po1006 = new_n3550;
  assign po1007 = new_n3552;
  assign po1008 = new_n3554;
  assign po1009 = new_n3556;
  assign po1010 = new_n3558;
  assign po1011 = new_n3560;
  assign po1012 = new_n3562;
  assign po1013 = new_n3564;
  assign po1014 = new_n3566;
  assign po1015 = new_n3568;
  assign po1016 = new_n3570;
  assign po1017 = new_n3572;
  assign po1018 = new_n3574;
  assign po1019 = new_n3576;
  assign po1020 = new_n3578;
  assign po1021 = new_n3580;
  assign po1022 = new_n3582;
  assign po1023 = new_n3584;
  assign po1024 = new_n3587;
  assign po1025 = new_n3590;
  assign po1026 = new_n3593;
  assign po1027 = new_n3596;
  assign po1028 = new_n3599;
  assign po1029 = new_n3602;
  assign po1030 = new_n3605;
  assign po1031 = new_n3608;
  assign po1032 = new_n3611;
  assign po1033 = new_n3614;
  assign po1034 = new_n3617;
  assign po1035 = new_n3620;
  assign po1036 = new_n3623;
  assign po1037 = new_n3626;
  assign po1038 = new_n3629;
  assign po1039 = new_n3632;
  assign po1040 = new_n3635;
  assign po1041 = new_n3638;
  assign po1042 = new_n3641;
  assign po1043 = new_n3644;
  assign po1044 = new_n3647;
  assign po1045 = new_n3650;
  assign po1046 = new_n3653;
  assign po1047 = new_n3656;
  assign po1048 = new_n3659;
  assign po1049 = new_n3662;
  assign po1050 = new_n3665;
  assign po1051 = new_n3668;
  assign po1052 = new_n3671;
  assign po1053 = new_n3674;
  assign po1054 = new_n3677;
  assign po1055 = new_n3680;
  assign po1056 = new_n3683;
  assign po1057 = new_n3686;
  assign po1058 = new_n3689;
  assign po1059 = new_n3692;
  assign po1060 = new_n3695;
  assign po1061 = new_n3698;
  assign po1062 = new_n3701;
  assign po1063 = new_n3704;
  assign po1064 = new_n3707;
  assign po1065 = new_n3710;
  assign po1066 = new_n3713;
  assign po1067 = new_n3716;
  assign po1068 = new_n3719;
  assign po1069 = new_n3722;
  assign po1070 = new_n3725;
  assign po1071 = new_n3728;
  assign po1072 = new_n3731;
  assign po1073 = new_n3734;
  assign po1074 = new_n3737;
  assign po1075 = new_n3740;
  assign po1076 = new_n3743;
  assign po1077 = new_n3746;
  assign po1078 = new_n3749;
  assign po1079 = new_n3752;
  assign po1080 = new_n3755;
  assign po1081 = new_n3758;
  assign po1082 = new_n3761;
  assign po1083 = new_n3764;
  assign po1084 = new_n3767;
  assign po1085 = new_n3770;
  assign po1086 = new_n3773;
  assign po1087 = new_n3776;
  assign po1088 = new_n3779;
  assign po1089 = new_n3782;
  assign po1090 = new_n3785;
  assign po1091 = new_n3788;
  assign po1092 = new_n3791;
  assign po1093 = new_n3794;
  assign po1094 = new_n3797;
  assign po1095 = new_n3800;
  assign po1096 = new_n3803;
  assign po1097 = new_n3806;
  assign po1098 = new_n3809;
  assign po1099 = new_n3812;
  assign po1100 = new_n3815;
  assign po1101 = new_n3818;
  assign po1102 = new_n3821;
  assign po1103 = new_n3824;
  assign po1104 = new_n3827;
  assign po1105 = new_n3830;
  assign po1106 = new_n3833;
  assign po1107 = new_n3836;
  assign po1108 = new_n3839;
  assign po1109 = new_n3842;
  assign po1110 = new_n3845;
  assign po1111 = new_n3848;
  assign po1112 = new_n3851;
  assign po1113 = new_n3854;
  assign po1114 = new_n3857;
  assign po1115 = new_n3860;
  assign po1116 = new_n3863;
  assign po1117 = new_n3866;
  assign po1118 = new_n3869;
  assign po1119 = new_n3872;
  assign po1120 = new_n3875;
  assign po1121 = new_n3878;
  assign po1122 = new_n3881;
  assign po1123 = new_n3884;
  assign po1124 = new_n3887;
  assign po1125 = new_n3890;
  assign po1126 = new_n3893;
  assign po1127 = new_n3896;
  assign po1128 = new_n3899;
  assign po1129 = new_n3902;
  assign po1130 = new_n3905;
  assign po1131 = new_n3908;
  assign po1132 = new_n3911;
  assign po1133 = new_n3914;
  assign po1134 = new_n3917;
  assign po1135 = new_n3920;
  assign po1136 = new_n3923;
  assign po1137 = new_n3926;
  assign po1138 = new_n3929;
  assign po1139 = new_n3932;
  assign po1140 = new_n3935;
  assign po1141 = new_n3938;
  assign po1142 = new_n3941;
  assign po1143 = new_n3944;
  assign po1144 = new_n3947;
  assign po1145 = new_n3950;
  assign po1146 = new_n3953;
  assign po1147 = new_n3956;
  assign po1148 = new_n3959;
  assign po1149 = new_n3962;
  assign po1150 = new_n3965;
  assign po1151 = new_n3968;
  assign po1152 = new_n3970;
  assign po1153 = new_n3972;
  assign po1154 = new_n3974;
  assign po1155 = new_n3976;
  assign po1156 = new_n3978;
  assign po1157 = new_n3980;
  assign po1158 = new_n3982;
  assign po1159 = new_n3984;
  assign po1160 = new_n3986;
  assign po1161 = new_n3988;
  assign po1162 = new_n3990;
  assign po1163 = new_n3992;
  assign po1164 = new_n3994;
  assign po1165 = new_n3996;
  assign po1166 = new_n3998;
  assign po1167 = new_n4000;
  assign po1168 = new_n4002;
  assign po1169 = new_n4004;
  assign po1170 = new_n4006;
  assign po1171 = new_n4008;
  assign po1172 = new_n4010;
  assign po1173 = new_n4012;
  assign po1174 = new_n4014;
  assign po1175 = new_n4016;
  assign po1176 = new_n4018;
  assign po1177 = new_n4020;
  assign po1178 = new_n4022;
  assign po1179 = new_n4024;
  assign po1180 = new_n4026;
  assign po1181 = new_n4028;
  assign po1182 = new_n4030;
  assign po1183 = new_n4032;
  assign po1184 = new_n4034;
  assign po1185 = new_n4036;
  assign po1186 = new_n4038;
  assign po1187 = new_n4040;
  assign po1188 = new_n4042;
  assign po1189 = new_n4044;
  assign po1190 = new_n4046;
  assign po1191 = new_n4048;
  assign po1192 = new_n4050;
  assign po1193 = new_n4052;
  assign po1194 = new_n4054;
  assign po1195 = new_n4056;
  assign po1196 = new_n4058;
  assign po1197 = new_n4060;
  assign po1198 = new_n4062;
  assign po1199 = new_n4064;
  assign po1200 = new_n4066;
  assign po1201 = new_n4068;
  assign po1202 = new_n4070;
  assign po1203 = new_n4072;
  assign po1204 = new_n4074;
  assign po1205 = new_n4076;
  assign po1206 = new_n4078;
  assign po1207 = new_n4080;
  assign po1208 = new_n4082;
  assign po1209 = new_n4084;
  assign po1210 = new_n4086;
  assign po1211 = new_n4088;
  assign po1212 = new_n4090;
  assign po1213 = new_n4092;
  assign po1214 = new_n4094;
  assign po1215 = new_n4096;
  assign po1216 = new_n4098;
  assign po1217 = new_n4100;
  assign po1218 = new_n4102;
  assign po1219 = new_n4104;
  assign po1220 = new_n4106;
  assign po1221 = new_n4108;
  assign po1222 = new_n4110;
  assign po1223 = new_n4112;
  assign po1224 = new_n4114;
  assign po1225 = new_n4116;
  assign po1226 = new_n4118;
  assign po1227 = new_n4120;
  assign po1228 = new_n4122;
  assign po1229 = new_n4124;
  assign po1230 = new_n4126;
  assign po1231 = new_n4128;
  assign po1232 = new_n4130;
  assign po1233 = new_n4132;
  assign po1234 = new_n4134;
  assign po1235 = new_n4136;
  assign po1236 = new_n4138;
  assign po1237 = new_n4140;
  assign po1238 = new_n4142;
  assign po1239 = new_n4144;
  assign po1240 = new_n4146;
  assign po1241 = new_n4148;
  assign po1242 = new_n4150;
  assign po1243 = new_n4152;
  assign po1244 = new_n4154;
  assign po1245 = new_n4156;
  assign po1246 = new_n4158;
  assign po1247 = new_n4160;
  assign po1248 = new_n4162;
  assign po1249 = new_n4164;
  assign po1250 = new_n4166;
  assign po1251 = new_n4168;
  assign po1252 = new_n4170;
  assign po1253 = new_n4172;
  assign po1254 = new_n4174;
  assign po1255 = new_n4176;
  assign po1256 = new_n4178;
  assign po1257 = new_n4180;
  assign po1258 = new_n4182;
  assign po1259 = new_n4184;
  assign po1260 = new_n4186;
  assign po1261 = new_n4188;
  assign po1262 = new_n4190;
  assign po1263 = new_n4192;
  assign po1264 = new_n4194;
  assign po1265 = new_n4196;
  assign po1266 = new_n4198;
  assign po1267 = new_n4200;
  assign po1268 = new_n4202;
  assign po1269 = new_n4204;
  assign po1270 = new_n4206;
  assign po1271 = new_n4208;
  assign po1272 = new_n4210;
  assign po1273 = new_n4212;
  assign po1274 = new_n4214;
  assign po1275 = new_n4216;
  assign po1276 = new_n4218;
  assign po1277 = new_n4220;
  assign po1278 = new_n4222;
  assign po1279 = new_n4224;
  assign po1280 = new_n4226;
  assign po1281 = new_n4228;
  assign po1282 = new_n4230;
  assign po1283 = new_n4232;
  assign po1284 = new_n4234;
  assign po1285 = new_n4236;
  assign po1286 = new_n4238;
  assign po1287 = new_n4240;
  assign po1288 = new_n4242;
  assign po1289 = new_n4244;
  assign po1290 = new_n4246;
  assign po1291 = new_n4248;
  assign po1292 = new_n4250;
  assign po1293 = new_n4252;
  assign po1294 = new_n4254;
  assign po1295 = new_n4256;
  assign po1296 = new_n4258;
  assign po1297 = new_n4260;
  assign po1298 = new_n4262;
  assign po1299 = new_n4264;
  assign po1300 = new_n4266;
  assign po1301 = new_n4268;
  assign po1302 = new_n4270;
  assign po1303 = new_n4272;
  assign po1304 = new_n4274;
  assign po1305 = new_n4276;
  assign po1306 = new_n4278;
  assign po1307 = new_n4280;
  assign po1308 = new_n4282;
  assign po1309 = new_n4284;
  assign po1310 = new_n4286;
  assign po1311 = new_n4288;
  assign po1312 = new_n4290;
  assign po1313 = new_n4292;
  assign po1314 = new_n4294;
  assign po1315 = new_n4296;
  assign po1316 = new_n4298;
  assign po1317 = new_n4300;
  assign po1318 = new_n4302;
  assign po1319 = new_n4304;
  assign po1320 = new_n4306;
  assign po1321 = new_n4308;
  assign po1322 = new_n4310;
  assign po1323 = new_n4312;
  assign po1324 = new_n4314;
  assign po1325 = new_n4316;
  assign po1326 = new_n4318;
  assign po1327 = new_n4320;
  assign po1328 = new_n4322;
  assign po1329 = new_n4324;
  assign po1330 = new_n4326;
  assign po1331 = new_n4328;
  assign po1332 = new_n4330;
  assign po1333 = new_n4332;
  assign po1334 = new_n4334;
  assign po1335 = new_n4336;
  assign po1336 = new_n4338;
  assign po1337 = new_n4340;
  assign po1338 = new_n4342;
  assign po1339 = new_n4344;
  assign po1340 = new_n4346;
  assign po1341 = new_n4348;
  assign po1342 = new_n4350;
  assign po1343 = new_n4352;
  assign po1344 = new_n4354;
  assign po1345 = new_n4356;
  assign po1346 = new_n4358;
  assign po1347 = new_n4360;
  assign po1348 = new_n4362;
  assign po1349 = new_n4364;
  assign po1350 = new_n4366;
  assign po1351 = new_n4368;
  assign po1352 = new_n4370;
  assign po1353 = new_n4372;
  assign po1354 = new_n4374;
  assign po1355 = new_n4376;
  assign po1356 = new_n4378;
  assign po1357 = new_n4380;
  assign po1358 = new_n4382;
  assign po1359 = new_n4384;
  assign po1360 = new_n4386;
  assign po1361 = new_n4388;
  assign po1362 = new_n4390;
  assign po1363 = new_n4392;
  assign po1364 = new_n4394;
  assign po1365 = new_n4396;
  assign po1366 = new_n4398;
  assign po1367 = new_n4400;
  assign po1368 = new_n4402;
  assign po1369 = new_n4404;
  assign po1370 = new_n4406;
  assign po1371 = new_n4408;
  assign po1372 = new_n4410;
  assign po1373 = new_n4412;
  assign po1374 = new_n4414;
  assign po1375 = new_n4416;
  assign po1376 = new_n4418;
  assign po1377 = new_n4420;
  assign po1378 = new_n4422;
  assign po1379 = new_n4424;
  assign po1380 = new_n4426;
  assign po1381 = new_n4428;
  assign po1382 = new_n4430;
  assign po1383 = new_n4432;
  assign po1384 = new_n4434;
  assign po1385 = new_n4436;
  assign po1386 = new_n4438;
  assign po1387 = new_n4440;
  assign po1388 = new_n4442;
  assign po1389 = new_n4444;
  assign po1390 = new_n4446;
  assign po1391 = new_n4448;
  assign po1392 = new_n4450;
  assign po1393 = new_n4452;
  assign po1394 = new_n4454;
  assign po1395 = new_n4456;
  assign po1396 = new_n4458;
  assign po1397 = new_n4460;
  assign po1398 = new_n4462;
  assign po1399 = new_n4464;
  assign po1400 = new_n4466;
  assign po1401 = new_n4468;
  assign po1402 = new_n4470;
  assign po1403 = new_n4472;
  assign po1404 = new_n4474;
  assign po1405 = new_n4476;
  assign po1406 = new_n4478;
  assign po1407 = new_n4480;
  assign po1408 = new_n4483;
  assign po1409 = new_n4486;
  assign po1410 = new_n4489;
  assign po1411 = new_n4492;
  assign po1412 = new_n4495;
  assign po1413 = new_n4498;
  assign po1414 = new_n4501;
  assign po1415 = new_n4504;
  assign po1416 = new_n4507;
  assign po1417 = new_n4510;
  assign po1418 = new_n4513;
  assign po1419 = new_n4516;
  assign po1420 = new_n4519;
  assign po1421 = new_n4522;
  assign po1422 = new_n4525;
  assign po1423 = new_n4528;
  assign po1424 = new_n4531;
  assign po1425 = new_n4534;
  assign po1426 = new_n4537;
  assign po1427 = new_n4540;
  assign po1428 = new_n4543;
  assign po1429 = new_n4546;
  assign po1430 = new_n4549;
  assign po1431 = new_n4552;
  assign po1432 = new_n4555;
  assign po1433 = new_n4558;
  assign po1434 = new_n4561;
  assign po1435 = new_n4564;
  assign po1436 = new_n4567;
  assign po1437 = new_n4570;
  assign po1438 = new_n4573;
  assign po1439 = new_n4576;
  assign po1440 = new_n4579;
  assign po1441 = new_n4582;
  assign po1442 = new_n4585;
  assign po1443 = new_n4588;
  assign po1444 = new_n4591;
  assign po1445 = new_n4594;
  assign po1446 = new_n4597;
  assign po1447 = new_n4600;
  assign po1448 = new_n4603;
  assign po1449 = new_n4606;
  assign po1450 = new_n4609;
  assign po1451 = new_n4612;
  assign po1452 = new_n4615;
  assign po1453 = new_n4618;
  assign po1454 = new_n4621;
  assign po1455 = new_n4624;
  assign po1456 = new_n4627;
  assign po1457 = new_n4630;
  assign po1458 = new_n4633;
  assign po1459 = new_n4636;
  assign po1460 = new_n4639;
  assign po1461 = new_n4642;
  assign po1462 = new_n4645;
  assign po1463 = new_n4648;
  assign po1464 = new_n4651;
  assign po1465 = new_n4654;
  assign po1466 = new_n4657;
  assign po1467 = new_n4660;
  assign po1468 = new_n4663;
  assign po1469 = new_n4666;
  assign po1470 = new_n4669;
  assign po1471 = new_n4672;
  assign po1472 = new_n4674;
  assign po1473 = new_n4676;
  assign po1474 = new_n4678;
  assign po1475 = new_n4680;
  assign po1476 = new_n4682;
  assign po1477 = new_n4684;
  assign po1478 = new_n4686;
  assign po1479 = new_n4688;
  assign po1480 = new_n4690;
  assign po1481 = new_n4692;
  assign po1482 = new_n4694;
  assign po1483 = new_n4696;
  assign po1484 = new_n4698;
  assign po1485 = new_n4700;
  assign po1486 = new_n4702;
  assign po1487 = new_n4704;
  assign po1488 = new_n4706;
  assign po1489 = new_n4708;
  assign po1490 = new_n4710;
  assign po1491 = new_n4712;
  assign po1492 = new_n4714;
  assign po1493 = new_n4716;
  assign po1494 = new_n4718;
  assign po1495 = new_n4720;
  assign po1496 = new_n4722;
  assign po1497 = new_n4724;
  assign po1498 = new_n4726;
  assign po1499 = new_n4728;
  assign po1500 = new_n4730;
  assign po1501 = new_n4732;
  assign po1502 = new_n4734;
  assign po1503 = new_n4736;
  assign po1504 = new_n4738;
  assign po1505 = new_n4740;
  assign po1506 = new_n4742;
  assign po1507 = new_n4744;
  assign po1508 = new_n4746;
  assign po1509 = new_n4748;
  assign po1510 = new_n4750;
  assign po1511 = new_n4752;
  assign po1512 = new_n4754;
  assign po1513 = new_n4756;
  assign po1514 = new_n4758;
  assign po1515 = new_n4760;
  assign po1516 = new_n4762;
  assign po1517 = new_n4764;
  assign po1518 = new_n4766;
  assign po1519 = new_n4768;
  assign po1520 = new_n4770;
  assign po1521 = new_n4772;
  assign po1522 = new_n4774;
  assign po1523 = new_n4776;
  assign po1524 = new_n4778;
  assign po1525 = new_n4780;
  assign po1526 = new_n4782;
  assign po1527 = new_n4784;
  assign po1528 = new_n4786;
  assign po1529 = new_n4788;
  assign po1530 = new_n4790;
  assign po1531 = new_n4792;
  assign po1532 = new_n4794;
  assign po1533 = new_n4796;
  assign po1534 = new_n4798;
  assign po1535 = new_n4800;
  assign po1536 = new_n4802;
  assign po1537 = new_n4804;
  assign po1538 = new_n4806;
  assign po1539 = new_n4808;
  assign po1540 = new_n4810;
  assign po1541 = new_n4812;
  assign po1542 = new_n4814;
  assign po1543 = new_n4816;
  assign po1544 = new_n4818;
  assign po1545 = new_n4820;
  assign po1546 = new_n4822;
  assign po1547 = new_n4824;
  assign po1548 = new_n4826;
  assign po1549 = new_n4828;
  assign po1550 = new_n4830;
  assign po1551 = new_n4832;
  assign po1552 = new_n4834;
  assign po1553 = new_n4836;
  assign po1554 = new_n4838;
  assign po1555 = new_n4840;
  assign po1556 = new_n4842;
  assign po1557 = new_n4844;
  assign po1558 = new_n4846;
  assign po1559 = new_n4848;
  assign po1560 = new_n4850;
  assign po1561 = new_n4852;
  assign po1562 = new_n4854;
  assign po1563 = new_n4856;
  assign po1564 = new_n4858;
  assign po1565 = new_n4860;
  assign po1566 = new_n4862;
  assign po1567 = new_n4864;
  assign po1568 = new_n4866;
  assign po1569 = new_n4868;
  assign po1570 = new_n4870;
  assign po1571 = new_n4872;
  assign po1572 = new_n4874;
  assign po1573 = new_n4876;
  assign po1574 = new_n4878;
  assign po1575 = new_n4880;
  assign po1576 = new_n4882;
  assign po1577 = new_n4884;
  assign po1578 = new_n4886;
  assign po1579 = new_n4888;
  assign po1580 = new_n4890;
  assign po1581 = new_n4892;
  assign po1582 = new_n4894;
  assign po1583 = new_n4896;
  assign po1584 = new_n4898;
  assign po1585 = new_n4900;
  assign po1586 = new_n4902;
  assign po1587 = new_n4904;
  assign po1588 = new_n4906;
  assign po1589 = new_n4908;
  assign po1590 = new_n4910;
  assign po1591 = new_n4912;
  assign po1592 = new_n4914;
  assign po1593 = new_n4916;
  assign po1594 = new_n4918;
  assign po1595 = new_n4920;
  assign po1596 = new_n4922;
  assign po1597 = new_n4924;
  assign po1598 = new_n4926;
  assign po1599 = new_n4928;
  assign po1625 = new_n4928;
  assign po1626 = new_n4926;
  assign po1627 = new_n4924;
  assign po1628 = new_n4922;
  assign po1629 = new_n4920;
  assign po1630 = new_n4918;
  assign po1631 = new_n4916;
  assign po1632 = new_n4914;
  assign po1633 = new_n4912;
  assign po1634 = new_n4910;
  assign po1635 = new_n4908;
  assign po1636 = new_n4906;
  assign po1637 = new_n4904;
  assign po1638 = new_n4902;
  assign po1639 = new_n4900;
  assign po1640 = new_n4898;
  assign po1641 = new_n4896;
  assign po1642 = new_n4894;
  assign po1643 = new_n4892;
  assign po1644 = new_n4890;
  assign po1645 = new_n4888;
  assign po1646 = new_n4886;
  assign po1647 = new_n4884;
  assign po1648 = new_n4882;
  assign po1649 = new_n4880;
  assign po1650 = new_n4878;
  assign po1651 = new_n4876;
  assign po1652 = new_n4874;
  assign po1653 = new_n4872;
  assign po1654 = new_n4870;
  assign po1655 = new_n4868;
  assign po1656 = new_n4866;
  assign po1657 = new_n4864;
  assign po1658 = new_n4862;
  assign po1659 = new_n4860;
  assign po1660 = new_n4858;
  assign po1661 = new_n4856;
  assign po1662 = new_n4854;
  assign po1663 = new_n4852;
  assign po1664 = new_n4850;
  assign po1665 = new_n4848;
  assign po1666 = new_n4846;
  assign po1667 = new_n4844;
  assign po1668 = new_n4842;
  assign po1669 = new_n4840;
  assign po1670 = new_n4838;
  assign po1671 = new_n4836;
  assign po1672 = new_n4834;
  assign po1673 = new_n4832;
  assign po1674 = new_n4830;
  assign po1675 = new_n4828;
  assign po1676 = new_n4826;
  assign po1677 = new_n4824;
  assign po1678 = new_n4822;
  assign po1679 = new_n4820;
  assign po1680 = new_n4818;
  assign po1681 = new_n4816;
  assign po1682 = new_n4814;
  assign po1683 = new_n4812;
  assign po1684 = new_n4810;
  assign po1685 = new_n4808;
  assign po1686 = new_n4806;
  assign po1687 = new_n4804;
  assign po1688 = new_n4802;
  assign po1689 = new_n4800;
  assign po1690 = new_n4798;
  assign po1691 = new_n4796;
  assign po1692 = new_n4794;
  assign po1693 = new_n4792;
  assign po1694 = new_n4790;
  assign po1695 = new_n4788;
  assign po1696 = new_n4786;
  assign po1697 = new_n4784;
  assign po1698 = new_n4782;
  assign po1699 = new_n4780;
  assign po1700 = new_n4778;
  assign po1701 = new_n4776;
  assign po1702 = new_n4774;
  assign po1703 = new_n4772;
  assign po1704 = new_n4770;
  assign po1705 = new_n4768;
  assign po1706 = new_n4766;
  assign po1707 = new_n4764;
  assign po1708 = new_n4762;
  assign po1709 = new_n4760;
  assign po1710 = new_n4758;
  assign po1711 = new_n4756;
  assign po1712 = new_n4754;
  assign po1713 = new_n4752;
  assign po1714 = new_n4750;
  assign po1715 = new_n4748;
  assign po1716 = new_n4746;
  assign po1717 = new_n4744;
  assign po1718 = new_n4742;
  assign po1719 = new_n4740;
  assign po1720 = new_n4738;
  assign po1721 = new_n4736;
  assign po1722 = new_n4734;
  assign po1723 = new_n4732;
  assign po1724 = new_n4730;
  assign po1725 = new_n4728;
  assign po1726 = new_n4726;
  assign po1727 = new_n4724;
  assign po1728 = new_n4722;
  assign po1729 = new_n4720;
  assign po1730 = new_n4718;
  assign po1731 = new_n4716;
  assign po1732 = new_n4714;
  assign po1733 = new_n4712;
  assign po1734 = new_n4710;
  assign po1735 = new_n4708;
  assign po1736 = new_n4706;
  assign po1737 = new_n4704;
  assign po1738 = new_n4702;
  assign po1739 = new_n4700;
  assign po1740 = new_n4698;
  assign po1741 = new_n4696;
  assign po1742 = new_n4694;
  assign po1743 = new_n4692;
  assign po1744 = new_n4690;
  assign po1745 = new_n4688;
  assign po1746 = new_n4686;
  assign po1747 = new_n4684;
  assign po1748 = new_n4682;
  assign po1749 = new_n4680;
  assign po1750 = new_n4678;
  assign po1751 = new_n4676;
  assign po1752 = new_n4674;
  assign po1753 = new_n4672;
  assign po1754 = new_n4669;
  assign po1755 = new_n4666;
  assign po1756 = new_n4663;
  assign po1757 = new_n4660;
  assign po1758 = new_n4657;
  assign po1759 = new_n4654;
  assign po1760 = new_n4651;
  assign po1761 = new_n4648;
  assign po1762 = new_n4645;
  assign po1763 = new_n4642;
  assign po1764 = new_n4639;
  assign po1765 = new_n4636;
  assign po1766 = new_n4633;
  assign po1767 = new_n4630;
  assign po1768 = new_n4627;
  assign po1769 = new_n4624;
  assign po1770 = new_n4621;
  assign po1771 = new_n4618;
  assign po1772 = new_n4615;
  assign po1773 = new_n4612;
  assign po1774 = new_n4609;
  assign po1775 = new_n4606;
  assign po1776 = new_n4603;
  assign po1777 = new_n4600;
  assign po1778 = new_n4597;
  assign po1779 = new_n4594;
  assign po1780 = new_n4591;
  assign po1781 = new_n4588;
  assign po1782 = new_n4585;
  assign po1783 = new_n4582;
  assign po1784 = new_n4579;
  assign po1785 = new_n4576;
  assign po1786 = new_n4573;
  assign po1787 = new_n4570;
  assign po1788 = new_n4567;
  assign po1789 = new_n4564;
  assign po1790 = new_n4561;
  assign po1791 = new_n4558;
  assign po1792 = new_n4555;
  assign po1793 = new_n4552;
  assign po1794 = new_n4549;
  assign po1795 = new_n4546;
  assign po1796 = new_n4543;
  assign po1797 = new_n4540;
  assign po1798 = new_n4537;
  assign po1799 = new_n4534;
  assign po1800 = new_n4531;
  assign po1801 = new_n4528;
  assign po1802 = new_n4525;
  assign po1803 = new_n4522;
  assign po1804 = new_n4519;
  assign po1805 = new_n4516;
  assign po1806 = new_n4513;
  assign po1807 = new_n4510;
  assign po1808 = new_n4507;
  assign po1809 = new_n4504;
  assign po1810 = new_n4501;
  assign po1811 = new_n4498;
  assign po1812 = new_n4495;
  assign po1813 = new_n4492;
  assign po1814 = new_n4489;
  assign po1815 = new_n4486;
  assign po1816 = new_n4483;
  assign po1817 = new_n4480;
  assign po1818 = new_n4478;
  assign po1819 = new_n4476;
  assign po1820 = new_n4474;
  assign po1821 = new_n4472;
  assign po1822 = new_n4470;
  assign po1823 = new_n4468;
  assign po1824 = new_n4466;
  assign po1825 = new_n4464;
  assign po1826 = new_n4462;
  assign po1827 = new_n4460;
  assign po1828 = new_n4458;
  assign po1829 = new_n4456;
  assign po1830 = new_n4454;
  assign po1831 = new_n4452;
  assign po1832 = new_n4450;
  assign po1833 = new_n4448;
  assign po1834 = new_n4446;
  assign po1835 = new_n4444;
  assign po1836 = new_n4442;
  assign po1837 = new_n4440;
  assign po1838 = new_n4438;
  assign po1839 = new_n4436;
  assign po1840 = new_n4434;
  assign po1841 = new_n4432;
  assign po1842 = new_n4430;
  assign po1843 = new_n4428;
  assign po1844 = new_n4426;
  assign po1845 = new_n4424;
  assign po1846 = new_n4422;
  assign po1847 = new_n4420;
  assign po1848 = new_n4418;
  assign po1849 = new_n4416;
  assign po1850 = new_n4414;
  assign po1851 = new_n4412;
  assign po1852 = new_n4410;
  assign po1853 = new_n4408;
  assign po1854 = new_n4406;
  assign po1855 = new_n4404;
  assign po1856 = new_n4402;
  assign po1857 = new_n4400;
  assign po1858 = new_n4398;
  assign po1859 = new_n4396;
  assign po1860 = new_n4394;
  assign po1861 = new_n4392;
  assign po1862 = new_n4390;
  assign po1863 = new_n4388;
  assign po1864 = new_n4386;
  assign po1865 = new_n4384;
  assign po1866 = new_n4382;
  assign po1867 = new_n4380;
  assign po1868 = new_n4378;
  assign po1869 = new_n4376;
  assign po1870 = new_n4374;
  assign po1871 = new_n4372;
  assign po1872 = new_n4370;
  assign po1873 = new_n4368;
  assign po1874 = new_n4366;
  assign po1875 = new_n4364;
  assign po1876 = new_n4362;
  assign po1877 = new_n4360;
  assign po1878 = new_n4358;
  assign po1879 = new_n4356;
  assign po1880 = new_n4354;
  assign po1881 = new_n4352;
  assign po1882 = new_n4350;
  assign po1883 = new_n4348;
  assign po1884 = new_n4346;
  assign po1885 = new_n4344;
  assign po1886 = new_n4342;
  assign po1887 = new_n4340;
  assign po1888 = new_n4338;
  assign po1889 = new_n4336;
  assign po1890 = new_n4334;
  assign po1891 = new_n4332;
  assign po1892 = new_n4330;
  assign po1893 = new_n4328;
  assign po1894 = new_n4326;
  assign po1895 = new_n4324;
  assign po1896 = new_n4322;
  assign po1897 = new_n4320;
  assign po1898 = new_n4318;
  assign po1899 = new_n4316;
  assign po1900 = new_n4314;
  assign po1901 = new_n4312;
  assign po1902 = new_n4310;
  assign po1903 = new_n4308;
  assign po1904 = new_n4306;
  assign po1905 = new_n4304;
  assign po1906 = new_n4302;
  assign po1907 = new_n4300;
  assign po1908 = new_n4298;
  assign po1909 = new_n4296;
  assign po1910 = new_n4294;
  assign po1911 = new_n4292;
  assign po1912 = new_n4290;
  assign po1913 = new_n4288;
  assign po1914 = new_n4286;
  assign po1915 = new_n4284;
  assign po1916 = new_n4282;
  assign po1917 = new_n4280;
  assign po1918 = new_n4278;
  assign po1919 = new_n4276;
  assign po1920 = new_n4274;
  assign po1921 = new_n4272;
  assign po1922 = new_n4270;
  assign po1923 = new_n4268;
  assign po1924 = new_n4266;
  assign po1925 = new_n4264;
  assign po1926 = new_n4262;
  assign po1927 = new_n4260;
  assign po1928 = new_n4258;
  assign po1929 = new_n4256;
  assign po1930 = new_n4254;
  assign po1931 = new_n4252;
  assign po1932 = new_n4250;
  assign po1933 = new_n4248;
  assign po1934 = new_n4246;
  assign po1935 = new_n4244;
  assign po1936 = new_n4242;
  assign po1937 = new_n4240;
  assign po1938 = new_n4238;
  assign po1939 = new_n4236;
  assign po1940 = new_n4234;
  assign po1941 = new_n4232;
  assign po1942 = new_n4230;
  assign po1943 = new_n4228;
  assign po1944 = new_n4226;
  assign po1945 = new_n4224;
  assign po1946 = new_n4222;
  assign po1947 = new_n4220;
  assign po1948 = new_n4218;
  assign po1949 = new_n4216;
  assign po1950 = new_n4214;
  assign po1951 = new_n4212;
  assign po1952 = new_n4210;
  assign po1953 = new_n4208;
  assign po1954 = new_n4206;
  assign po1955 = new_n4204;
  assign po1956 = new_n4202;
  assign po1957 = new_n4200;
  assign po1958 = new_n4198;
  assign po1959 = new_n4196;
  assign po1960 = new_n4194;
  assign po1961 = new_n4192;
  assign po1962 = new_n4190;
  assign po1963 = new_n4188;
  assign po1964 = new_n4186;
  assign po1965 = new_n4184;
  assign po1966 = new_n4182;
  assign po1967 = new_n4180;
  assign po1968 = new_n4178;
  assign po1969 = new_n4176;
  assign po1970 = new_n4174;
  assign po1971 = new_n4172;
  assign po1972 = new_n4170;
  assign po1973 = new_n4168;
  assign po1974 = new_n4166;
  assign po1975 = new_n4164;
  assign po1976 = new_n4162;
  assign po1977 = new_n4160;
  assign po1978 = new_n4158;
  assign po1979 = new_n4156;
  assign po1980 = new_n4154;
  assign po1981 = new_n4152;
  assign po1982 = new_n4150;
  assign po1983 = new_n4148;
  assign po1984 = new_n4146;
  assign po1985 = new_n4144;
  assign po1986 = new_n4142;
  assign po1987 = new_n4140;
  assign po1988 = new_n4138;
  assign po1989 = new_n4136;
  assign po1990 = new_n4134;
  assign po1991 = new_n4132;
  assign po1992 = new_n4130;
  assign po1993 = new_n4128;
  assign po1994 = new_n4126;
  assign po1995 = new_n4124;
  assign po1996 = new_n4122;
  assign po1997 = new_n4120;
  assign po1998 = new_n4118;
  assign po1999 = new_n4116;
  assign po2000 = new_n4114;
  assign po2001 = new_n4112;
  assign po2002 = new_n4110;
  assign po2003 = new_n4108;
  assign po2004 = new_n4106;
  assign po2005 = new_n4104;
  assign po2006 = new_n4102;
  assign po2007 = new_n4100;
  assign po2008 = new_n4098;
  assign po2009 = new_n4096;
  assign po2010 = new_n4094;
  assign po2011 = new_n4092;
  assign po2012 = new_n4090;
  assign po2013 = new_n4088;
  assign po2014 = new_n4086;
  assign po2015 = new_n4084;
  assign po2016 = new_n4082;
  assign po2017 = new_n4080;
  assign po2018 = new_n4078;
  assign po2019 = new_n4076;
  assign po2020 = new_n4074;
  assign po2021 = new_n4072;
  assign po2022 = new_n4070;
  assign po2023 = new_n4068;
  assign po2024 = new_n4066;
  assign po2025 = new_n4064;
  assign po2026 = new_n4062;
  assign po2027 = new_n4060;
  assign po2028 = new_n4058;
  assign po2029 = new_n4056;
  assign po2030 = new_n4054;
  assign po2031 = new_n4052;
  assign po2032 = new_n4050;
  assign po2033 = new_n4048;
  assign po2034 = new_n4046;
  assign po2035 = new_n4044;
  assign po2036 = new_n4042;
  assign po2037 = new_n4040;
  assign po2038 = new_n4038;
  assign po2039 = new_n4036;
  assign po2040 = new_n4034;
  assign po2041 = new_n4032;
  assign po2042 = new_n4030;
  assign po2043 = new_n4028;
  assign po2044 = new_n4026;
  assign po2045 = new_n4024;
  assign po2046 = new_n4022;
  assign po2047 = new_n4020;
  assign po2048 = new_n4018;
  assign po2049 = new_n4016;
  assign po2050 = new_n4014;
  assign po2051 = new_n4012;
  assign po2052 = new_n4010;
  assign po2053 = new_n4008;
  assign po2054 = new_n4006;
  assign po2055 = new_n4004;
  assign po2056 = new_n4002;
  assign po2057 = new_n4000;
  assign po2058 = new_n3998;
  assign po2059 = new_n3996;
  assign po2060 = new_n3994;
  assign po2061 = new_n3992;
  assign po2062 = new_n3990;
  assign po2063 = new_n3988;
  assign po2064 = new_n3986;
  assign po2065 = new_n3984;
  assign po2066 = new_n3982;
  assign po2067 = new_n3980;
  assign po2068 = new_n3978;
  assign po2069 = new_n3976;
  assign po2070 = new_n3974;
  assign po2071 = new_n3972;
  assign po2072 = new_n3970;
  assign po2073 = new_n3968;
  assign po2074 = new_n3965;
  assign po2075 = new_n3962;
  assign po2076 = new_n3959;
  assign po2077 = new_n3956;
  assign po2078 = new_n3953;
  assign po2079 = new_n3950;
  assign po2080 = new_n3947;
  assign po2081 = new_n3944;
  assign po2082 = new_n3941;
  assign po2083 = new_n3938;
  assign po2084 = new_n3935;
  assign po2085 = new_n3932;
  assign po2086 = new_n3929;
  assign po2087 = new_n3926;
  assign po2088 = new_n3923;
  assign po2089 = new_n3920;
  assign po2090 = new_n3917;
  assign po2091 = new_n3914;
  assign po2092 = new_n3911;
  assign po2093 = new_n3908;
  assign po2094 = new_n3905;
  assign po2095 = new_n3902;
  assign po2096 = new_n3899;
  assign po2097 = new_n3896;
  assign po2098 = new_n3893;
  assign po2099 = new_n3890;
  assign po2100 = new_n3887;
  assign po2101 = new_n3884;
  assign po2102 = new_n3881;
  assign po2103 = new_n3878;
  assign po2104 = new_n3875;
  assign po2105 = new_n3872;
  assign po2106 = new_n3869;
  assign po2107 = new_n3866;
  assign po2108 = new_n3863;
  assign po2109 = new_n3860;
  assign po2110 = new_n3857;
  assign po2111 = new_n3854;
  assign po2112 = new_n3851;
  assign po2113 = new_n3848;
  assign po2114 = new_n3845;
  assign po2115 = new_n3842;
  assign po2116 = new_n3839;
  assign po2117 = new_n3836;
  assign po2118 = new_n3833;
  assign po2119 = new_n3830;
  assign po2120 = new_n3827;
  assign po2121 = new_n3824;
  assign po2122 = new_n3821;
  assign po2123 = new_n3818;
  assign po2124 = new_n3815;
  assign po2125 = new_n3812;
  assign po2126 = new_n3809;
  assign po2127 = new_n3806;
  assign po2128 = new_n3803;
  assign po2129 = new_n3800;
  assign po2130 = new_n3797;
  assign po2131 = new_n3794;
  assign po2132 = new_n3791;
  assign po2133 = new_n3788;
  assign po2134 = new_n3785;
  assign po2135 = new_n3782;
  assign po2136 = new_n3779;
  assign po2137 = new_n3776;
  assign po2138 = new_n3773;
  assign po2139 = new_n3770;
  assign po2140 = new_n3767;
  assign po2141 = new_n3764;
  assign po2142 = new_n3761;
  assign po2143 = new_n3758;
  assign po2144 = new_n3755;
  assign po2145 = new_n3752;
  assign po2146 = new_n3749;
  assign po2147 = new_n3746;
  assign po2148 = new_n3743;
  assign po2149 = new_n3740;
  assign po2150 = new_n3737;
  assign po2151 = new_n3734;
  assign po2152 = new_n3731;
  assign po2153 = new_n3728;
  assign po2154 = new_n3725;
  assign po2155 = new_n3722;
  assign po2156 = new_n3719;
  assign po2157 = new_n3716;
  assign po2158 = new_n3713;
  assign po2159 = new_n3710;
  assign po2160 = new_n3707;
  assign po2161 = new_n3704;
  assign po2162 = new_n3701;
  assign po2163 = new_n3698;
  assign po2164 = new_n3695;
  assign po2165 = new_n3692;
  assign po2166 = new_n3689;
  assign po2167 = new_n3686;
  assign po2168 = new_n3683;
  assign po2169 = new_n3680;
  assign po2170 = new_n3677;
  assign po2171 = new_n3674;
  assign po2172 = new_n3671;
  assign po2173 = new_n3668;
  assign po2174 = new_n3665;
  assign po2175 = new_n3662;
  assign po2176 = new_n3659;
  assign po2177 = new_n3656;
  assign po2178 = new_n3653;
  assign po2179 = new_n3650;
  assign po2180 = new_n3647;
  assign po2181 = new_n3644;
  assign po2182 = new_n3641;
  assign po2183 = new_n3638;
  assign po2184 = new_n3635;
  assign po2185 = new_n3632;
  assign po2186 = new_n3629;
  assign po2187 = new_n3626;
  assign po2188 = new_n3623;
  assign po2189 = new_n3620;
  assign po2190 = new_n3617;
  assign po2191 = new_n3614;
  assign po2192 = new_n3611;
  assign po2193 = new_n3608;
  assign po2194 = new_n3605;
  assign po2195 = new_n3602;
  assign po2196 = new_n3599;
  assign po2197 = new_n3596;
  assign po2198 = new_n3593;
  assign po2199 = new_n3590;
  assign po2200 = new_n3587;
  assign po2201 = new_n3584;
  assign po2202 = new_n3582;
  assign po2203 = new_n3580;
  assign po2204 = new_n3578;
  assign po2205 = new_n3576;
  assign po2206 = new_n3574;
  assign po2207 = new_n3572;
  assign po2208 = new_n3570;
  assign po2209 = new_n3568;
  assign po2210 = new_n3566;
  assign po2211 = new_n3564;
  assign po2212 = new_n3562;
  assign po2213 = new_n3560;
  assign po2214 = new_n3558;
  assign po2215 = new_n3556;
  assign po2216 = new_n3554;
  assign po2217 = new_n3552;
  assign po2218 = new_n3550;
  assign po2219 = new_n3548;
  assign po2220 = new_n3546;
  assign po2221 = new_n3544;
  assign po2222 = new_n3542;
  assign po2223 = new_n3540;
  assign po2224 = new_n3538;
  assign po2225 = new_n3536;
  assign po2226 = new_n3534;
  assign po2227 = new_n3532;
  assign po2228 = new_n3530;
  assign po2229 = new_n3528;
  assign po2230 = new_n3526;
  assign po2231 = new_n3524;
  assign po2232 = new_n3522;
  assign po2233 = new_n3520;
  assign po2234 = new_n3518;
  assign po2235 = new_n3516;
  assign po2236 = new_n3514;
  assign po2237 = new_n3512;
  assign po2238 = new_n3510;
  assign po2239 = new_n3508;
  assign po2240 = new_n3506;
  assign po2241 = new_n3504;
  assign po2242 = new_n3502;
  assign po2243 = new_n3500;
  assign po2244 = new_n3498;
  assign po2245 = new_n3496;
  assign po2246 = new_n3494;
  assign po2247 = new_n3492;
  assign po2248 = new_n3490;
  assign po2249 = new_n3488;
  assign po2250 = new_n3486;
  assign po2251 = new_n3484;
  assign po2252 = new_n3482;
  assign po2253 = new_n3480;
  assign po2254 = new_n3478;
  assign po2255 = new_n3476;
  assign po2256 = new_n3474;
  assign po2257 = new_n3472;
  assign po2258 = new_n3470;
  assign po2259 = new_n3468;
  assign po2260 = new_n3466;
  assign po2261 = new_n3464;
  assign po2262 = new_n3462;
  assign po2263 = new_n3460;
  assign po2264 = new_n3458;
  assign po2265 = new_n3456;
  assign po2266 = new_n3454;
  assign po2267 = new_n3452;
  assign po2268 = new_n3450;
  assign po2269 = new_n3448;
  assign po2270 = new_n3446;
  assign po2271 = new_n3444;
  assign po2272 = new_n3442;
  assign po2273 = new_n3440;
  assign po2274 = new_n3438;
  assign po2275 = new_n3436;
  assign po2276 = new_n3434;
  assign po2277 = new_n3432;
  assign po2278 = new_n3430;
  assign po2279 = new_n3428;
  assign po2280 = new_n3426;
  assign po2281 = new_n3424;
  assign po2282 = new_n3422;
  assign po2283 = new_n3420;
  assign po2284 = new_n3418;
  assign po2285 = new_n3416;
  assign po2286 = new_n3414;
  assign po2287 = new_n3412;
  assign po2288 = new_n3410;
  assign po2289 = new_n3408;
  assign po2290 = new_n3406;
  assign po2291 = new_n3404;
  assign po2292 = new_n3402;
  assign po2293 = new_n3400;
  assign po2294 = new_n3398;
  assign po2295 = new_n3396;
  assign po2296 = new_n3394;
  assign po2297 = new_n3392;
  assign po2298 = new_n3390;
  assign po2299 = new_n3388;
  assign po2300 = new_n3386;
  assign po2301 = new_n3384;
  assign po2302 = new_n3382;
  assign po2303 = new_n3380;
  assign po2304 = new_n3378;
  assign po2305 = new_n3376;
  assign po2306 = new_n3374;
  assign po2307 = new_n3372;
  assign po2308 = new_n3370;
  assign po2309 = new_n3368;
  assign po2310 = new_n3366;
  assign po2311 = new_n3364;
  assign po2312 = new_n3362;
  assign po2313 = new_n3360;
  assign po2314 = new_n3358;
  assign po2315 = new_n3356;
  assign po2316 = new_n3354;
  assign po2317 = new_n3352;
  assign po2318 = new_n3350;
  assign po2319 = new_n3348;
  assign po2320 = new_n3346;
  assign po2321 = new_n3344;
  assign po2322 = new_n3342;
  assign po2323 = new_n3340;
  assign po2324 = new_n3338;
  assign po2325 = new_n3336;
  assign po2326 = new_n3334;
  assign po2327 = new_n3332;
  assign po2328 = new_n3330;
  assign po2329 = new_n3328;
  assign po2330 = new_n3326;
  assign po2331 = new_n3324;
  assign po2332 = new_n3322;
  assign po2333 = new_n3320;
  assign po2334 = new_n3318;
  assign po2335 = new_n3316;
  assign po2336 = new_n3314;
  assign po2337 = new_n3312;
  assign po2338 = new_n3310;
  assign po2339 = new_n3308;
  assign po2340 = new_n3306;
  assign po2341 = new_n3304;
  assign po2342 = new_n3302;
  assign po2343 = new_n3300;
  assign po2344 = new_n3298;
  assign po2345 = new_n3296;
  assign po2346 = new_n3294;
  assign po2347 = new_n3292;
  assign po2348 = new_n3290;
  assign po2349 = new_n3288;
  assign po2350 = new_n3286;
  assign po2351 = new_n3284;
  assign po2352 = new_n3282;
  assign po2353 = new_n3280;
  assign po2354 = new_n3278;
  assign po2355 = new_n3276;
  assign po2356 = new_n3274;
  assign po2357 = new_n3272;
  assign po2358 = new_n3270;
  assign po2359 = new_n3268;
  assign po2360 = new_n3266;
  assign po2361 = new_n3264;
  assign po2362 = new_n3262;
  assign po2363 = new_n3260;
  assign po2364 = new_n3258;
  assign po2365 = new_n3256;
  assign po2366 = new_n3254;
  assign po2367 = new_n3252;
  assign po2368 = new_n3250;
  assign po2369 = new_n3248;
  assign po2370 = new_n3246;
  assign po2371 = new_n3244;
  assign po2372 = new_n3242;
  assign po2373 = new_n3240;
  assign po2374 = new_n3238;
  assign po2375 = new_n3236;
  assign po2376 = new_n3234;
  assign po2377 = new_n3232;
  assign po2378 = new_n3230;
  assign po2379 = new_n3228;
  assign po2380 = new_n3226;
  assign po2381 = new_n3224;
  assign po2382 = new_n3222;
  assign po2383 = new_n3220;
  assign po2384 = new_n3218;
  assign po2385 = new_n3216;
  assign po2386 = new_n3214;
  assign po2387 = new_n3212;
  assign po2388 = new_n3210;
  assign po2389 = new_n3208;
  assign po2390 = new_n3206;
  assign po2391 = new_n3204;
  assign po2392 = new_n3202;
  assign po2393 = new_n3200;
  assign po2394 = new_n3197;
  assign po2395 = new_n3194;
  assign po2396 = new_n3191;
  assign po2397 = new_n3188;
  assign po2398 = new_n3185;
  assign po2399 = new_n3182;
  assign po2400 = new_n3179;
  assign po2401 = new_n3176;
  assign po2402 = new_n3173;
  assign po2403 = new_n3170;
  assign po2404 = new_n3167;
  assign po2405 = new_n3164;
  assign po2406 = new_n3161;
  assign po2407 = new_n3158;
  assign po2408 = new_n3155;
  assign po2409 = new_n3152;
  assign po2410 = new_n3149;
  assign po2411 = new_n3146;
  assign po2412 = new_n3143;
  assign po2413 = new_n3140;
  assign po2414 = new_n3137;
  assign po2415 = new_n3134;
  assign po2416 = new_n3131;
  assign po2417 = new_n3128;
  assign po2418 = new_n3125;
  assign po2419 = new_n3122;
  assign po2420 = new_n3119;
  assign po2421 = new_n3116;
  assign po2422 = new_n3113;
  assign po2423 = new_n3110;
  assign po2424 = new_n3107;
  assign po2425 = new_n3104;
  assign po2426 = new_n3101;
  assign po2427 = new_n3098;
  assign po2428 = new_n3095;
  assign po2429 = new_n3092;
  assign po2430 = new_n3089;
  assign po2431 = new_n3086;
  assign po2432 = new_n3083;
  assign po2433 = new_n3080;
  assign po2434 = new_n3077;
  assign po2435 = new_n3074;
  assign po2436 = new_n3071;
  assign po2437 = new_n3068;
  assign po2438 = new_n3065;
  assign po2439 = new_n3062;
  assign po2440 = new_n3059;
  assign po2441 = new_n3056;
  assign po2442 = new_n3053;
  assign po2443 = new_n3050;
  assign po2444 = new_n3047;
  assign po2445 = new_n3044;
  assign po2446 = new_n3041;
  assign po2447 = new_n3038;
  assign po2448 = new_n3035;
  assign po2449 = new_n3032;
  assign po2450 = new_n3029;
  assign po2451 = new_n3026;
  assign po2452 = new_n3023;
  assign po2453 = new_n3020;
  assign po2454 = new_n3017;
  assign po2455 = new_n3014;
  assign po2456 = new_n3011;
  assign po2457 = new_n3008;
  assign po2458 = new_n3005;
  assign po2459 = new_n3002;
  assign po2460 = new_n2999;
  assign po2461 = new_n2996;
  assign po2462 = new_n2993;
  assign po2463 = new_n2990;
  assign po2464 = new_n2987;
  assign po2465 = new_n2984;
  assign po2466 = new_n2981;
  assign po2467 = new_n2978;
  assign po2468 = new_n2975;
  assign po2469 = new_n2972;
  assign po2470 = new_n2969;
  assign po2471 = new_n2966;
  assign po2472 = new_n2963;
  assign po2473 = new_n2960;
  assign po2474 = new_n2957;
  assign po2475 = new_n2954;
  assign po2476 = new_n2951;
  assign po2477 = new_n2948;
  assign po2478 = new_n2945;
  assign po2479 = new_n2942;
  assign po2480 = new_n2939;
  assign po2481 = new_n2936;
  assign po2482 = new_n2933;
  assign po2483 = new_n2930;
  assign po2484 = new_n2927;
  assign po2485 = new_n2924;
  assign po2486 = new_n2921;
  assign po2487 = new_n2918;
  assign po2488 = new_n2915;
  assign po2489 = new_n2912;
  assign po2490 = new_n2909;
  assign po2491 = new_n2906;
  assign po2492 = new_n2903;
  assign po2493 = new_n2900;
  assign po2494 = new_n2897;
  assign po2495 = new_n2894;
  assign po2496 = new_n2891;
  assign po2497 = new_n2888;
  assign po2498 = new_n2885;
  assign po2499 = new_n2882;
  assign po2500 = new_n2879;
  assign po2501 = new_n2876;
  assign po2502 = new_n2873;
  assign po2503 = new_n2870;
  assign po2504 = new_n2867;
  assign po2505 = new_n2864;
  assign po2506 = new_n2861;
  assign po2507 = new_n2858;
  assign po2508 = new_n2855;
  assign po2509 = new_n2852;
  assign po2510 = new_n2849;
  assign po2511 = new_n2846;
  assign po2512 = new_n2843;
  assign po2513 = new_n2840;
  assign po2514 = new_n2837;
  assign po2515 = new_n2834;
  assign po2516 = new_n2831;
  assign po2517 = new_n2828;
  assign po2518 = new_n2825;
  assign po2519 = new_n2822;
  assign po2520 = new_n2819;
  assign po2521 = new_n2816;
  assign po2522 = new_n2814;
  assign po2523 = new_n2812;
  assign po2524 = new_n2810;
  assign po2525 = new_n2808;
  assign po2526 = new_n2806;
  assign po2527 = new_n2804;
  assign po2528 = new_n2802;
  assign po2529 = new_n2800;
  assign po2530 = new_n2798;
  assign po2531 = new_n2796;
  assign po2532 = new_n2794;
  assign po2533 = new_n2792;
  assign po2534 = new_n2790;
  assign po2535 = new_n2788;
  assign po2536 = new_n2786;
  assign po2537 = new_n2784;
  assign po2538 = new_n2782;
  assign po2539 = new_n2780;
  assign po2540 = new_n2778;
  assign po2541 = new_n2776;
  assign po2542 = new_n2774;
  assign po2543 = new_n2772;
  assign po2544 = new_n2770;
  assign po2545 = new_n2768;
  assign po2546 = new_n2766;
  assign po2547 = new_n2764;
  assign po2548 = new_n2762;
  assign po2549 = new_n2760;
  assign po2550 = new_n2758;
  assign po2551 = new_n2756;
  assign po2552 = new_n2754;
  assign po2553 = new_n2752;
  assign po2554 = new_n2750;
  assign po2555 = new_n2748;
  assign po2556 = new_n2746;
  assign po2557 = new_n2744;
  assign po2558 = new_n2742;
  assign po2559 = new_n2740;
  assign po2560 = new_n2738;
  assign po2561 = new_n2736;
  assign po2562 = new_n2734;
  assign po2563 = new_n2732;
  assign po2564 = new_n2730;
  assign po2565 = new_n2728;
  assign po2566 = new_n2726;
  assign po2567 = new_n2724;
  assign po2568 = new_n2722;
  assign po2569 = new_n2720;
  assign po2570 = new_n2718;
  assign po2571 = new_n2716;
  assign po2572 = new_n2714;
  assign po2573 = new_n2712;
  assign po2574 = new_n2710;
  assign po2575 = new_n2708;
  assign po2576 = new_n2706;
  assign po2577 = new_n2704;
  assign po2578 = new_n2702;
  assign po2579 = new_n2700;
  assign po2580 = new_n2698;
  assign po2581 = new_n2696;
  assign po2582 = new_n2694;
  assign po2583 = new_n2692;
  assign po2584 = new_n2690;
  assign po2585 = new_n2688;
  assign po2586 = new_n2686;
  assign po2587 = new_n2684;
  assign po2588 = new_n2682;
  assign po2589 = new_n2680;
  assign po2590 = new_n2678;
  assign po2591 = new_n2676;
  assign po2592 = new_n2674;
  assign po2593 = new_n2672;
  assign po2594 = new_n2670;
  assign po2595 = new_n2668;
  assign po2596 = new_n2666;
  assign po2597 = new_n2664;
  assign po2598 = new_n2662;
  assign po2599 = new_n2660;
  assign po2600 = new_n2658;
  assign po2601 = new_n2656;
  assign po2602 = new_n2654;
  assign po2603 = new_n2652;
  assign po2604 = new_n2650;
  assign po2605 = new_n2648;
  assign po2606 = new_n2646;
  assign po2607 = new_n2644;
  assign po2608 = new_n2642;
  assign po2609 = new_n2640;
  assign po2610 = new_n2638;
  assign po2611 = new_n2636;
  assign po2612 = new_n2634;
  assign po2613 = new_n2632;
  assign po2614 = new_n2630;
  assign po2615 = new_n2628;
  assign po2616 = new_n2626;
  assign po2617 = new_n2624;
  assign po2618 = new_n2622;
  assign po2619 = new_n2620;
  assign po2620 = new_n2618;
  assign po2621 = new_n2616;
  assign po2622 = new_n2614;
  assign po2623 = new_n2612;
  assign po2624 = new_n2610;
  assign po2625 = new_n2608;
  assign po2626 = new_n2606;
  assign po2627 = new_n2604;
  assign po2628 = new_n2602;
  assign po2629 = new_n2600;
  assign po2630 = new_n2598;
  assign po2631 = new_n2596;
  assign po2632 = new_n2594;
  assign po2633 = new_n2592;
  assign po2634 = new_n2590;
  assign po2635 = new_n2588;
  assign po2636 = new_n2586;
  assign po2637 = new_n2584;
  assign po2638 = new_n2582;
  assign po2639 = new_n2580;
  assign po2640 = new_n2578;
  assign po2641 = new_n2576;
  assign po2642 = new_n2574;
  assign po2643 = new_n2572;
  assign po2644 = new_n2570;
  assign po2645 = new_n2568;
  assign po2646 = new_n2566;
  assign po2647 = new_n2564;
  assign po2648 = new_n2562;
  assign po2649 = new_n2560;
  assign po2650 = new_n2558;
  assign po2651 = new_n2556;
  assign po2652 = new_n2554;
  assign po2653 = new_n2552;
  assign po2654 = new_n2550;
  assign po2655 = new_n2548;
  assign po2656 = new_n2546;
  assign po2657 = new_n2544;
  assign po2658 = new_n2542;
  assign po2659 = new_n2540;
  assign po2660 = new_n2538;
  assign po2661 = new_n2536;
  assign po2662 = new_n2534;
  assign po2663 = new_n2532;
  assign po2664 = new_n2530;
  assign po2665 = new_n2528;
  assign po2666 = new_n2526;
  assign po2667 = new_n2524;
  assign po2668 = new_n2522;
  assign po2669 = new_n2520;
  assign po2670 = new_n2518;
  assign po2671 = new_n2516;
  assign po2672 = new_n2514;
  assign po2673 = new_n2512;
  assign po2674 = new_n2510;
  assign po2675 = new_n2508;
  assign po2676 = new_n2506;
  assign po2677 = new_n2504;
  assign po2678 = new_n2502;
  assign po2679 = new_n2500;
  assign po2680 = new_n2498;
  assign po2681 = new_n2496;
  assign po2682 = new_n2494;
  assign po2683 = new_n2492;
  assign po2684 = new_n2490;
  assign po2685 = new_n2488;
  assign po2686 = new_n2486;
  assign po2687 = new_n2484;
  assign po2688 = new_n2482;
  assign po2689 = new_n2480;
  assign po2690 = new_n2478;
  assign po2691 = new_n2476;
  assign po2692 = new_n2474;
  assign po2693 = new_n2472;
  assign po2694 = new_n2470;
  assign po2695 = new_n2468;
  assign po2696 = new_n2466;
  assign po2697 = new_n2464;
  assign po2698 = new_n2462;
  assign po2699 = new_n2460;
  assign po2700 = new_n2458;
  assign po2701 = new_n2456;
  assign po2702 = new_n2454;
  assign po2703 = new_n2452;
  assign po2704 = new_n2450;
  assign po2705 = new_n2448;
  assign po2706 = new_n2446;
  assign po2707 = new_n2444;
  assign po2708 = new_n2442;
  assign po2709 = new_n2440;
  assign po2710 = new_n2438;
  assign po2711 = new_n2436;
  assign po2712 = new_n2434;
  assign po2713 = new_n2432;
  assign po2714 = new_n2429;
  assign po2715 = new_n2426;
  assign po2716 = new_n2423;
  assign po2717 = new_n2420;
  assign po2718 = new_n2417;
  assign po2719 = new_n2414;
  assign po2720 = new_n2411;
  assign po2721 = new_n2408;
  assign po2722 = new_n2405;
  assign po2723 = new_n2402;
  assign po2724 = new_n2399;
  assign po2725 = new_n2396;
  assign po2726 = new_n2393;
  assign po2727 = new_n2390;
  assign po2728 = new_n2387;
  assign po2729 = new_n2384;
  assign po2730 = new_n2381;
  assign po2731 = new_n2378;
  assign po2732 = new_n2375;
  assign po2733 = new_n2372;
  assign po2734 = new_n2369;
  assign po2735 = new_n2366;
  assign po2736 = new_n2363;
  assign po2737 = new_n2360;
  assign po2738 = new_n2357;
  assign po2739 = new_n2354;
  assign po2740 = new_n2351;
  assign po2741 = new_n2348;
  assign po2742 = new_n2345;
  assign po2743 = new_n2342;
  assign po2744 = new_n2339;
  assign po2745 = new_n2336;
  assign po2746 = new_n2333;
  assign po2747 = new_n2330;
  assign po2748 = new_n2327;
  assign po2749 = new_n2324;
  assign po2750 = new_n2321;
  assign po2751 = new_n2318;
  assign po2752 = new_n2315;
  assign po2753 = new_n2312;
  assign po2754 = new_n2309;
  assign po2755 = new_n2306;
  assign po2756 = new_n2303;
  assign po2757 = new_n2300;
  assign po2758 = new_n2297;
  assign po2759 = new_n2294;
  assign po2760 = new_n2291;
  assign po2761 = new_n2288;
  assign po2762 = new_n2285;
  assign po2763 = new_n2282;
  assign po2764 = new_n2279;
  assign po2765 = new_n2276;
  assign po2766 = new_n2273;
  assign po2767 = new_n2270;
  assign po2768 = new_n2267;
  assign po2769 = new_n2264;
  assign po2770 = new_n2261;
  assign po2771 = new_n2258;
  assign po2772 = new_n2255;
  assign po2773 = new_n2252;
  assign po2774 = new_n2249;
  assign po2775 = new_n2246;
  assign po2776 = new_n2243;
  assign po2777 = new_n2240;
  assign po2778 = new_n2237;
  assign po2779 = new_n2234;
  assign po2780 = new_n2231;
  assign po2781 = new_n2228;
  assign po2782 = new_n2225;
  assign po2783 = new_n2222;
  assign po2784 = new_n2219;
  assign po2785 = new_n2216;
  assign po2786 = new_n2213;
  assign po2787 = new_n2210;
  assign po2788 = new_n2207;
  assign po2789 = new_n2204;
  assign po2790 = new_n2201;
  assign po2791 = new_n2198;
  assign po2792 = new_n2195;
  assign po2793 = new_n2192;
  assign po2794 = new_n2189;
  assign po2795 = new_n2186;
  assign po2796 = new_n2183;
  assign po2797 = new_n2180;
  assign po2798 = new_n2177;
  assign po2799 = new_n2174;
  assign po2800 = new_n2171;
  assign po2801 = new_n2168;
  assign po2802 = new_n2165;
  assign po2803 = new_n2162;
  assign po2804 = new_n2159;
  assign po2805 = new_n2156;
  assign po2806 = new_n2153;
  assign po2807 = new_n2150;
  assign po2808 = new_n2147;
  assign po2809 = new_n2144;
  assign po2810 = new_n2141;
  assign po2811 = new_n2138;
  assign po2812 = new_n2135;
  assign po2813 = new_n2132;
  assign po2814 = new_n2129;
  assign po2815 = new_n2126;
  assign po2816 = new_n2123;
  assign po2817 = new_n2120;
  assign po2818 = new_n2117;
  assign po2819 = new_n2114;
  assign po2820 = new_n2111;
  assign po2821 = new_n2108;
  assign po2822 = new_n2105;
  assign po2823 = new_n2102;
  assign po2824 = new_n2099;
  assign po2825 = new_n2096;
  assign po2826 = new_n2093;
  assign po2827 = new_n2090;
  assign po2828 = new_n2087;
  assign po2829 = new_n2084;
  assign po2830 = new_n2081;
  assign po2831 = new_n2078;
  assign po2832 = new_n2075;
  assign po2833 = new_n2072;
  assign po2834 = new_n2069;
  assign po2835 = new_n2066;
  assign po2836 = new_n2063;
  assign po2837 = new_n2060;
  assign po2838 = new_n2057;
  assign po2839 = new_n2054;
  assign po2840 = new_n2051;
  assign po2841 = new_n2048;
  assign po2842 = new_n2046;
  assign po2843 = new_n2044;
  assign po2844 = new_n2042;
  assign po2845 = new_n2040;
  assign po2846 = new_n2038;
  assign po2847 = new_n2036;
  assign po2848 = new_n2034;
  assign po2849 = new_n2032;
  assign po2850 = new_n2030;
  assign po2851 = new_n2028;
  assign po2852 = new_n2026;
  assign po2853 = new_n2024;
  assign po2854 = new_n2022;
  assign po2855 = new_n2020;
  assign po2856 = new_n2018;
  assign po2857 = new_n2016;
  assign po2858 = new_n2014;
  assign po2859 = new_n2012;
  assign po2860 = new_n2010;
  assign po2861 = new_n2008;
  assign po2862 = new_n2006;
  assign po2863 = new_n2004;
  assign po2864 = new_n2002;
  assign po2865 = new_n2000;
  assign po2866 = new_n1998;
  assign po2867 = new_n1996;
  assign po2868 = new_n1994;
  assign po2869 = new_n1992;
  assign po2870 = new_n1990;
  assign po2871 = new_n1988;
  assign po2872 = new_n1986;
  assign po2873 = new_n1984;
  assign po2874 = new_n1982;
  assign po2875 = new_n1980;
  assign po2876 = new_n1978;
  assign po2877 = new_n1976;
  assign po2878 = new_n1974;
  assign po2879 = new_n1972;
  assign po2880 = new_n1970;
  assign po2881 = new_n1968;
  assign po2882 = new_n1966;
  assign po2883 = new_n1964;
  assign po2884 = new_n1962;
  assign po2885 = new_n1960;
  assign po2886 = new_n1958;
  assign po2887 = new_n1956;
  assign po2888 = new_n1954;
  assign po2889 = new_n1952;
  assign po2890 = new_n1950;
  assign po2891 = new_n1948;
  assign po2892 = new_n1946;
  assign po2893 = new_n1944;
  assign po2894 = new_n1942;
  assign po2895 = new_n1940;
  assign po2896 = new_n1938;
  assign po2897 = new_n1936;
  assign po2898 = new_n1934;
  assign po2899 = new_n1932;
  assign po2900 = new_n1930;
  assign po2901 = new_n1928;
  assign po2902 = new_n1926;
  assign po2903 = new_n1924;
  assign po2904 = new_n1922;
  assign po2905 = new_n1920;
  assign po2906 = new_n1918;
  assign po2907 = new_n1916;
  assign po2908 = new_n1914;
  assign po2909 = new_n1912;
  assign po2910 = new_n1910;
  assign po2911 = new_n1908;
  assign po2912 = new_n1906;
  assign po2913 = new_n1904;
  assign po2914 = new_n1902;
  assign po2915 = new_n1900;
  assign po2916 = new_n1898;
  assign po2917 = new_n1896;
  assign po2918 = new_n1894;
  assign po2919 = new_n1892;
  assign po2920 = new_n1890;
  assign po2921 = new_n1888;
  assign po2922 = new_n1886;
  assign po2923 = new_n1884;
  assign po2924 = new_n1882;
  assign po2925 = new_n1880;
  assign po2926 = new_n1878;
  assign po2927 = new_n1876;
  assign po2928 = new_n1874;
  assign po2929 = new_n1872;
  assign po2930 = new_n1870;
  assign po2931 = new_n1868;
  assign po2932 = new_n1866;
  assign po2933 = new_n1864;
  assign po2934 = new_n1862;
  assign po2935 = new_n1860;
  assign po2936 = new_n1858;
  assign po2937 = new_n1856;
  assign po2938 = new_n1854;
  assign po2939 = new_n1852;
  assign po2940 = new_n1850;
  assign po2941 = new_n1848;
  assign po2942 = new_n1846;
  assign po2943 = new_n1844;
  assign po2944 = new_n1842;
  assign po2945 = new_n1840;
  assign po2946 = new_n1838;
  assign po2947 = new_n1836;
  assign po2948 = new_n1834;
  assign po2949 = new_n1832;
  assign po2950 = new_n1830;
  assign po2951 = new_n1828;
  assign po2952 = new_n1826;
  assign po2953 = new_n1824;
  assign po2954 = new_n1822;
  assign po2955 = new_n1820;
  assign po2956 = new_n1818;
  assign po2957 = new_n1816;
  assign po2958 = new_n1814;
  assign po2959 = new_n1812;
  assign po2960 = new_n1810;
  assign po2961 = new_n1808;
  assign po2962 = new_n1806;
  assign po2963 = new_n1804;
  assign po2964 = new_n1802;
  assign po2965 = new_n1800;
  assign po2966 = new_n1798;
  assign po2967 = new_n1796;
  assign po2968 = new_n1794;
  assign po2969 = new_n1792;
  assign po2970 = new_n1790;
  assign po2971 = new_n1788;
  assign po2972 = new_n1786;
  assign po2973 = new_n1784;
  assign po2974 = new_n1782;
  assign po2975 = new_n1780;
  assign po2976 = new_n1778;
  assign po2977 = new_n1776;
  assign po2978 = new_n1774;
  assign po2979 = new_n1772;
  assign po2980 = new_n1770;
  assign po2981 = new_n1768;
  assign po2982 = new_n1766;
  assign po2983 = new_n1764;
  assign po2984 = new_n1762;
  assign po2985 = new_n1760;
  assign po2986 = new_n1758;
  assign po2987 = new_n1756;
  assign po2988 = new_n1754;
  assign po2989 = new_n1752;
  assign po2990 = new_n1750;
  assign po2991 = new_n1748;
  assign po2992 = new_n1746;
  assign po2993 = new_n1744;
  assign po2994 = new_n1742;
  assign po2995 = new_n1740;
  assign po2996 = new_n1738;
  assign po2997 = new_n1736;
  assign po2998 = new_n1734;
  assign po2999 = new_n1732;
  assign po3000 = new_n1730;
  assign po3001 = new_n1728;
  assign po3002 = new_n1726;
  assign po3003 = new_n1724;
  assign po3004 = new_n1722;
  assign po3005 = new_n1720;
  assign po3006 = new_n1718;
  assign po3007 = new_n1716;
  assign po3008 = new_n1714;
  assign po3009 = new_n1712;
  assign po3010 = new_n1710;
  assign po3011 = new_n1708;
  assign po3012 = new_n1706;
  assign po3013 = new_n1704;
  assign po3014 = new_n1702;
  assign po3015 = new_n1700;
  assign po3016 = new_n1698;
  assign po3017 = new_n1696;
  assign po3018 = new_n1694;
  assign po3019 = new_n1692;
  assign po3020 = new_n1690;
  assign po3021 = new_n1688;
  assign po3022 = new_n1686;
  assign po3023 = new_n1684;
  assign po3024 = new_n1682;
  assign po3025 = new_n1680;
  assign po3026 = new_n1678;
  assign po3027 = new_n1676;
  assign po3028 = new_n1674;
  assign po3029 = new_n1672;
  assign po3030 = new_n1670;
  assign po3031 = new_n1668;
  assign po3032 = new_n1666;
  assign po3033 = new_n1664;
  assign po3034 = new_n1660;
  assign po3035 = new_n1656;
  assign po3036 = new_n1652;
  assign po3037 = new_n1648;
  assign po3038 = new_n1644;
  assign po3039 = new_n1640;
  assign po3040 = new_n1636;
  assign po3041 = new_n1632;
  assign po3042 = new_n1628;
  assign po3043 = new_n1624;
  assign po3044 = new_n1620;
  assign po3045 = new_n1616;
  assign po3046 = new_n1612;
  assign po3047 = new_n1608;
  assign po3048 = new_n1604;
  assign po3049 = new_n1600;
  assign po3050 = new_n1596;
  assign po3051 = new_n1592;
  assign po3052 = new_n1588;
  assign po3053 = new_n1584;
  assign po3054 = new_n1580;
  assign po3055 = new_n1576;
  assign po3056 = new_n1572;
  assign po3057 = new_n1568;
  assign po3058 = new_n1564;
  assign po3059 = new_n1560;
  assign po3060 = new_n1556;
  assign po3061 = new_n1552;
  assign po3062 = new_n1548;
  assign po3063 = new_n1544;
  assign po3064 = new_n1540;
  assign po3065 = new_n1536;
  assign po3066 = new_n1532;
  assign po3067 = new_n1528;
  assign po3068 = new_n1524;
  assign po3069 = new_n1520;
  assign po3070 = new_n1516;
  assign po3071 = new_n1512;
  assign po3072 = new_n1508;
  assign po3073 = new_n1504;
  assign po3074 = new_n1500;
  assign po3075 = new_n1496;
  assign po3076 = new_n1492;
  assign po3077 = new_n1488;
  assign po3078 = new_n1484;
  assign po3079 = new_n1480;
  assign po3080 = new_n1476;
  assign po3081 = new_n1472;
  assign po3082 = new_n1468;
  assign po3083 = new_n1464;
  assign po3084 = new_n1460;
  assign po3085 = new_n1456;
  assign po3086 = new_n1452;
  assign po3087 = new_n1448;
  assign po3088 = new_n1444;
  assign po3089 = new_n1440;
  assign po3090 = new_n1436;
  assign po3091 = new_n1432;
  assign po3092 = new_n1428;
  assign po3093 = new_n1424;
  assign po3094 = new_n1420;
  assign po3095 = new_n1416;
  assign po3096 = new_n1412;
  assign po3097 = new_n1408;
  assign po3098 = new_n1404;
  assign po3099 = new_n1400;
  assign po3100 = new_n1396;
  assign po3101 = new_n1392;
  assign po3102 = new_n1388;
  assign po3103 = new_n1384;
  assign po3104 = new_n1380;
  assign po3105 = new_n1376;
  assign po3106 = new_n1372;
  assign po3107 = new_n1368;
  assign po3108 = new_n1364;
  assign po3109 = new_n1360;
  assign po3110 = new_n1356;
  assign po3111 = new_n1352;
  assign po3112 = new_n1348;
  assign po3113 = new_n1344;
  assign po3114 = new_n1340;
  assign po3115 = new_n1336;
  assign po3116 = new_n1332;
  assign po3117 = new_n1328;
  assign po3118 = new_n1324;
  assign po3119 = new_n1320;
  assign po3120 = new_n1316;
  assign po3121 = new_n1312;
  assign po3122 = new_n1308;
  assign po3123 = new_n1304;
  assign po3124 = new_n1300;
  assign po3125 = new_n1296;
  assign po3126 = new_n1292;
  assign po3127 = new_n1288;
  assign po3128 = new_n1284;
  assign po3129 = new_n1280;
  assign po3130 = new_n1276;
  assign po3131 = new_n1272;
  assign po3132 = new_n1268;
  assign po3133 = new_n1264;
  assign po3134 = new_n1260;
  assign po3135 = new_n1256;
  assign po3136 = new_n1252;
  assign po3137 = new_n1248;
  assign po3138 = new_n1244;
  assign po3139 = new_n1240;
  assign po3140 = new_n1236;
  assign po3141 = new_n1232;
  assign po3142 = new_n1228;
  assign po3143 = new_n1224;
  assign po3144 = new_n1220;
  assign po3145 = new_n1216;
  assign po3146 = new_n1212;
  assign po3147 = new_n1208;
  assign po3148 = new_n1204;
  assign po3149 = new_n1200;
  assign po3150 = new_n1196;
  assign po3151 = new_n1192;
  assign po3152 = new_n1188;
  assign po3153 = new_n1184;
  assign po3154 = new_n1180;
  assign po3155 = new_n1176;
  assign po3156 = new_n1172;
  assign po3157 = new_n1168;
  assign po3158 = new_n1164;
  assign po3159 = new_n1160;
  assign po3160 = new_n1156;
  assign po3161 = new_n1152;
  assign po3162 = new_n1144;
  assign po3163 = new_n1136;
  assign po3164 = new_n1128;
  assign po3165 = new_n1120;
  assign po3166 = new_n1112;
  assign po3167 = new_n1104;
  assign po3168 = new_n1096;
  assign po3169 = new_n1088;
  assign po3170 = new_n1080;
  assign po3171 = new_n1072;
  assign po3172 = new_n1064;
  assign po3173 = new_n1056;
  assign po3174 = new_n1048;
  assign po3175 = new_n1040;
  assign po3176 = new_n1032;
  assign po3177 = new_n1024;
  assign po3178 = new_n1016;
  assign po3179 = new_n1008;
  assign po3180 = new_n1000;
  assign po3181 = new_n992;
  assign po3182 = new_n984;
  assign po3183 = new_n976;
  assign po3184 = new_n967;
  assign po3185 = new_n958;
  assign po3186 = new_n949;
  assign po3187 = new_n940;
  assign po3188 = new_n931;
  assign po3189 = new_n922;
  assign po3190 = new_n913;
  assign po3191 = new_n904;
  assign po3192 = new_n895;
  assign po3193 = new_n886;
  assign po3194 = new_n877;
  assign po3195 = new_n868;
  assign po3196 = new_n859;
  assign po3197 = new_n850;
  assign po3198 = new_n841;
  assign po3199 = new_n832;
  assign po3200 = new_n823;
  assign po3201 = new_n814;
  assign po3202 = new_n805;
  assign po3203 = new_n796;
  assign po3204 = new_n786;
  assign po3205 = new_n776;
  assign po3206 = new_n766;
  assign po3207 = new_n756;
  assign po3208 = new_n746;
  assign po3209 = new_n736;
  assign po3210 = new_n726;
  assign po3211 = new_n716;
  assign po3212 = new_n706;
  assign po3213 = new_n696;
  assign po3214 = new_n686;
  assign po3215 = new_n676;
  assign po3216 = new_n666;
  assign po3217 = new_n656;
  assign po3218 = new_n646;
  assign po3219 = new_n636;
  assign po3220 = new_n626;
  assign po3221 = new_n616;
  assign po3222 = new_n606;
  assign po3223 = new_n596;
  assign po3224 = new_n586;
  assign po1600 = 1'b1;
  assign po1601 = 1'b1;
  assign po1602 = 1'b0;
  assign po1603 = 1'b0;
  assign po1604 = 1'b0;
  assign po1605 = 1'b0;
  assign po1606 = 1'b0;
  assign po1607 = 1'b0;
  assign po1608 = 1'b0;
  assign po1609 = 1'b0;
  assign po1610 = 1'b0;
  assign po1611 = 1'b0;
  assign po1612 = 1'b0;
  assign po1613 = 1'b0;
  assign po1614 = 1'b0;
  assign po1615 = 1'b0;
  assign po1616 = 1'b0;
  assign po1617 = 1'b0;
  assign po1618 = 1'b0;
  assign po1619 = 1'b0;
  assign po1620 = 1'b0;
  assign po1621 = 1'b0;
  assign po1622 = 1'b0;
  assign po1623 = 1'b0;
  assign po1624 = 1'b0;
endmodule


