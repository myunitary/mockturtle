module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 ;
  assign n151 = ~x5 & ~x22 ;
  assign n184 = ~x56 & n151 ;
  assign n148 = ~x4 & ~x19 ;
  assign n149 = ~x16 & ~x18 ;
  assign n150 = n148 & n149 ;
  assign n152 = ~x6 & ~x12 ;
  assign n153 = ~x17 & n152 ;
  assign n154 = n151 & n153 ;
  assign n155 = n150 & n154 ;
  assign n156 = ~x8 & ~x21 ;
  assign n157 = ~x7 & ~x13 ;
  assign n172 = x10 & n157 ;
  assign n173 = n156 & n172 ;
  assign n164 = ~x7 & ~x8 ;
  assign n166 = x21 & n164 ;
  assign n165 = x13 & n164 ;
  assign n167 = n166 ^ n165 ;
  assign n162 = ~x21 & n157 ;
  assign n160 = ~x8 & ~x13 ;
  assign n161 = ~x21 & n160 ;
  assign n163 = n162 ^ n161 ;
  assign n168 = n167 ^ n163 ;
  assign n169 = ~x10 & ~x14 ;
  assign n170 = n168 & n169 ;
  assign n158 = x14 & n157 ;
  assign n159 = n156 & n158 ;
  assign n171 = n170 ^ n159 ;
  assign n174 = n173 ^ n171 ;
  assign n175 = ~x9 & ~x11 ;
  assign n178 = ~x56 & n175 ;
  assign n179 = ~n151 & n178 ;
  assign n180 = n174 & n179 ;
  assign n181 = n155 & n180 ;
  assign n176 = n174 & n175 ;
  assign n177 = n155 & n176 ;
  assign n182 = n181 ^ n177 ;
  assign n183 = n182 ^ n178 ;
  assign n185 = n184 ^ n183 ;
  assign n200 = x54 & ~n185 ;
  assign n198 = x0 & ~x54 ;
  assign n186 = ~x14 & ~x22 ;
  assign n187 = n157 & n186 ;
  assign n188 = n175 & n187 ;
  assign n189 = ~x17 & ~x21 ;
  assign n190 = ~x8 & n189 ;
  assign n191 = ~x5 & n152 ;
  assign n192 = n190 & n191 ;
  assign n193 = n188 & n192 ;
  assign n194 = ~x0 & x54 ;
  assign n195 = n150 & n194 ;
  assign n196 = n193 & n195 ;
  assign n197 = ~n185 & n196 ;
  assign n199 = n198 ^ n197 ;
  assign n201 = n200 ^ n199 ;
  assign n202 = ~x3 & ~x129 ;
  assign n203 = ~n201 & n202 ;
  assign n204 = ~x5 & ~x6 ;
  assign n205 = ~x7 & ~x12 ;
  assign n206 = ~n204 & ~n205 ;
  assign n207 = ~x13 & ~n206 ;
  assign n208 = ~x5 & ~x7 ;
  assign n209 = n208 ^ n152 ;
  assign n210 = n207 & n209 ;
  assign n211 = x13 & n152 ;
  assign n212 = n208 & n211 ;
  assign n213 = ~x9 & ~n212 ;
  assign n214 = ~n210 & n213 ;
  assign n215 = n157 & n191 ;
  assign n216 = x9 & ~n215 ;
  assign n217 = ~x10 & x54 ;
  assign n218 = n186 & n217 ;
  assign n219 = ~x8 & ~x11 ;
  assign n220 = n189 & n219 ;
  assign n221 = n218 & n220 ;
  assign n222 = n150 & n221 ;
  assign n223 = ~n216 & n222 ;
  assign n224 = ~n214 & n223 ;
  assign n225 = n157 & n204 ;
  assign n226 = n150 & n225 ;
  assign n227 = ~x14 & n156 ;
  assign n228 = ~x11 & ~x12 ;
  assign n229 = ~x10 & ~x22 ;
  assign n230 = n228 & n229 ;
  assign n231 = n227 & n230 ;
  assign n232 = n226 & n231 ;
  assign n233 = ~x17 & x54 ;
  assign n234 = ~x1 & n233 ;
  assign n235 = ~n232 & n234 ;
  assign n236 = n235 ^ x1 ;
  assign n237 = n202 & n236 ;
  assign n238 = ~n224 & n237 ;
  assign n239 = n238 ^ n202 ;
  assign n240 = ~x38 & ~x50 ;
  assign n241 = ~x40 & ~x46 ;
  assign n242 = n240 & n241 ;
  assign n243 = ~x41 & ~x43 ;
  assign n244 = ~x42 & ~x44 ;
  assign n245 = n243 & n244 ;
  assign n246 = n242 & n245 ;
  assign n247 = ~x47 & ~x48 ;
  assign n248 = n246 & n247 ;
  assign n249 = ~x15 & ~x20 ;
  assign n250 = ~x45 & n249 ;
  assign n251 = ~x24 & ~x49 ;
  assign n252 = x82 & n251 ;
  assign n253 = n250 & n252 ;
  assign n254 = x122 & x127 ;
  assign n255 = ~x82 & ~n254 ;
  assign n256 = x2 & ~n255 ;
  assign n257 = n253 & n256 ;
  assign n258 = n248 & n257 ;
  assign n259 = n258 ^ n256 ;
  assign n264 = n250 & n251 ;
  assign n265 = ~x41 & ~x46 ;
  assign n266 = n240 & n265 ;
  assign n267 = ~x43 & ~x47 ;
  assign n268 = ~x2 & ~x48 ;
  assign n269 = n267 & n268 ;
  assign n270 = n266 & n269 ;
  assign n271 = n264 & n270 ;
  assign n272 = ~x40 & n244 ;
  assign n260 = ~x65 & ~n254 ;
  assign n273 = x82 & n260 ;
  assign n274 = n272 & n273 ;
  assign n275 = n271 & n274 ;
  assign n276 = ~n259 & n275 ;
  assign n261 = ~x82 & n260 ;
  assign n262 = ~n259 & n261 ;
  assign n263 = n262 ^ n259 ;
  assign n277 = n276 ^ n263 ;
  assign n278 = ~x129 & n277 ;
  assign n285 = ~x9 & ~x14 ;
  assign n286 = n229 & n285 ;
  assign n287 = ~x12 & n220 ;
  assign n288 = n286 & n287 ;
  assign n279 = x0 & ~x113 ;
  assign n280 = ~x123 & n279 ;
  assign n281 = ~x61 & ~x118 ;
  assign n289 = ~x129 & n281 ;
  assign n290 = ~n280 & n289 ;
  assign n291 = n226 & n290 ;
  assign n292 = n288 & n291 ;
  assign n282 = ~x129 & ~n281 ;
  assign n283 = ~n280 & n282 ;
  assign n284 = n283 ^ x129 ;
  assign n293 = n292 ^ n284 ;
  assign n303 = x4 & ~x54 ;
  assign n307 = n202 & n303 ;
  assign n294 = ~x18 & n148 ;
  assign n295 = ~x16 & x54 ;
  assign n296 = n189 & n295 ;
  assign n297 = n294 & n296 ;
  assign n298 = x10 & ~x22 ;
  assign n299 = n219 & n298 ;
  assign n300 = n297 & n299 ;
  assign n301 = n157 & n285 ;
  assign n302 = n191 & n301 ;
  assign n304 = n202 & ~n303 ;
  assign n305 = n302 & n304 ;
  assign n306 = n300 & n305 ;
  assign n308 = n307 ^ n306 ;
  assign n309 = x5 & ~x54 ;
  assign n310 = ~x13 & n286 ;
  assign n311 = ~x59 & n220 ;
  assign n312 = n310 & n311 ;
  assign n313 = n152 & n208 ;
  assign n314 = n295 & n313 ;
  assign n315 = ~x25 & x28 ;
  assign n316 = ~x29 & n315 ;
  assign n317 = n294 & n316 ;
  assign n318 = n314 & n317 ;
  assign n319 = n312 & n318 ;
  assign n320 = ~n309 & ~n319 ;
  assign n321 = n202 & ~n320 ;
  assign n322 = x6 & ~x54 ;
  assign n323 = ~x28 & ~x29 ;
  assign n324 = x25 & n323 ;
  assign n325 = n294 & n324 ;
  assign n326 = n314 & n325 ;
  assign n327 = n312 & n326 ;
  assign n328 = ~n322 & ~n327 ;
  assign n329 = n202 & ~n328 ;
  assign n330 = x7 & ~x54 ;
  assign n331 = x8 & n297 ;
  assign n332 = ~x11 & n313 ;
  assign n333 = n310 & n332 ;
  assign n334 = n331 & n333 ;
  assign n335 = ~n330 & ~n334 ;
  assign n336 = n202 & ~n335 ;
  assign n337 = x8 & ~x54 ;
  assign n338 = ~x12 & n286 ;
  assign n339 = n225 & n338 ;
  assign n340 = n148 & n295 ;
  assign n341 = ~x17 & ~x18 ;
  assign n342 = n219 & n341 ;
  assign n343 = x21 & n342 ;
  assign n344 = n340 & n343 ;
  assign n345 = n339 & n344 ;
  assign n346 = ~n337 & ~n345 ;
  assign n347 = n202 & ~n346 ;
  assign n348 = x9 & ~x54 ;
  assign n349 = ~x8 & n297 ;
  assign n350 = x11 & n313 ;
  assign n351 = n310 & n350 ;
  assign n352 = n349 & n351 ;
  assign n353 = ~n348 & ~n352 ;
  assign n354 = n202 & ~n353 ;
  assign n355 = x10 & ~x54 ;
  assign n356 = ~x9 & ~x18 ;
  assign n357 = n190 & n356 ;
  assign n358 = n229 & n357 ;
  assign n359 = ~x13 & x14 ;
  assign n360 = n340 & n359 ;
  assign n361 = n332 & n360 ;
  assign n362 = n358 & n361 ;
  assign n363 = ~n355 & ~n362 ;
  assign n364 = n202 & ~n363 ;
  assign n367 = x11 & ~x54 ;
  assign n372 = n202 & n367 ;
  assign n365 = ~x10 & ~x11 ;
  assign n366 = x22 & n365 ;
  assign n368 = n202 & ~n367 ;
  assign n369 = n366 & n368 ;
  assign n370 = n302 & n369 ;
  assign n371 = n349 & n370 ;
  assign n373 = n372 ^ n371 ;
  assign n374 = x12 & ~x54 ;
  assign n375 = x18 & n225 ;
  assign n376 = n286 & n340 ;
  assign n377 = n375 & n376 ;
  assign n378 = n287 & n377 ;
  assign n379 = ~n374 & ~n378 ;
  assign n380 = n202 & ~n379 ;
  assign n381 = ~x25 & ~x28 ;
  assign n382 = x29 & n381 ;
  assign n383 = ~x59 & n229 ;
  assign n384 = n382 & n383 ;
  assign n385 = n297 & n384 ;
  assign n386 = x13 & ~x54 ;
  assign n387 = n219 & ~n386 ;
  assign n388 = n302 & n387 ;
  assign n389 = n385 & n388 ;
  assign n390 = n389 ^ n386 ;
  assign n391 = n202 & n390 ;
  assign n392 = x14 & ~x54 ;
  assign n393 = x13 & ~x16 ;
  assign n394 = n148 & n393 ;
  assign n395 = n218 & n394 ;
  assign n396 = n332 & n395 ;
  assign n397 = n357 & n396 ;
  assign n398 = ~n392 & ~n397 ;
  assign n399 = n202 & ~n398 ;
  assign n415 = n266 & n272 ;
  assign n416 = ~x45 & n251 ;
  assign n417 = ~x48 & n267 ;
  assign n418 = n416 & n417 ;
  assign n419 = n415 & n418 ;
  assign n420 = x15 & ~n419 ;
  assign n421 = ~x15 & n251 ;
  assign n422 = ~x45 & n247 ;
  assign n423 = ~x2 & ~x20 ;
  assign n424 = n422 & ~n423 ;
  assign n425 = n421 & n424 ;
  assign n426 = n246 & n425 ;
  assign n427 = ~n420 & ~n426 ;
  assign n400 = n247 & n251 ;
  assign n401 = ~x15 & ~x45 ;
  assign n402 = n243 & n401 ;
  assign n403 = n400 & n402 ;
  assign n404 = x82 & n244 ;
  assign n405 = n242 & n404 ;
  assign n406 = n403 & n405 ;
  assign n407 = n406 ^ x82 ;
  assign n408 = ~x82 & n254 ;
  assign n409 = x15 & n408 ;
  assign n410 = ~x70 & ~n254 ;
  assign n411 = ~n409 & n410 ;
  assign n412 = ~n407 & n411 ;
  assign n413 = n412 ^ n409 ;
  assign n428 = x82 & ~x129 ;
  assign n429 = ~n413 & n428 ;
  assign n430 = ~n427 & n429 ;
  assign n414 = ~x129 & n413 ;
  assign n431 = n430 ^ n414 ;
  assign n432 = x16 & ~x54 ;
  assign n433 = n219 & n297 ;
  assign n434 = x6 & ~x13 ;
  assign n435 = n208 & n434 ;
  assign n436 = n338 & n435 ;
  assign n437 = n433 & n436 ;
  assign n438 = ~n432 & ~n437 ;
  assign n439 = n202 & ~n438 ;
  assign n440 = x17 & ~x54 ;
  assign n441 = ~x25 & x59 ;
  assign n442 = n156 & n441 ;
  assign n443 = n233 & n323 ;
  assign n444 = n442 & n443 ;
  assign n445 = n150 & n444 ;
  assign n446 = n333 & n445 ;
  assign n447 = ~n440 & ~n446 ;
  assign n448 = n202 & ~n447 ;
  assign n453 = x18 & ~x54 ;
  assign n457 = n202 & n453 ;
  assign n449 = n225 & n294 ;
  assign n450 = n338 & n449 ;
  assign n451 = x16 & x54 ;
  assign n452 = n220 & n451 ;
  assign n454 = n202 & ~n453 ;
  assign n455 = n452 & n454 ;
  assign n456 = n450 & n455 ;
  assign n458 = n457 ^ n456 ;
  assign n462 = x19 & ~x54 ;
  assign n466 = n202 & n462 ;
  assign n459 = x17 & ~x21 ;
  assign n460 = n219 & n459 ;
  assign n461 = n295 & n460 ;
  assign n463 = n202 & ~n462 ;
  assign n464 = n461 & n463 ;
  assign n465 = n450 & n464 ;
  assign n467 = n466 ^ n465 ;
  assign n482 = x20 & x82 ;
  assign n468 = ~x46 & ~x50 ;
  assign n469 = ~x38 & ~x40 ;
  assign n470 = n244 & n469 ;
  assign n471 = n468 & n470 ;
  assign n472 = n243 & n251 ;
  assign n473 = n422 & n472 ;
  assign n474 = n471 & n473 ;
  assign n479 = ~x15 & x82 ;
  assign n480 = n474 & n479 ;
  assign n475 = ~x2 & ~x15 ;
  assign n476 = ~x20 & x82 ;
  assign n477 = n475 & n476 ;
  assign n478 = n474 & n477 ;
  assign n481 = n480 ^ n478 ;
  assign n483 = n482 ^ n481 ;
  assign n484 = x20 & n408 ;
  assign n485 = ~x71 & ~n254 ;
  assign n489 = x82 & n249 ;
  assign n490 = n485 & n489 ;
  assign n491 = ~n484 & n490 ;
  assign n492 = n474 & n491 ;
  assign n486 = ~x82 & n485 ;
  assign n487 = ~n484 & n486 ;
  assign n488 = n487 ^ n484 ;
  assign n493 = n492 ^ n488 ;
  assign n494 = ~n483 & ~n493 ;
  assign n495 = ~x129 & ~n494 ;
  assign n496 = x21 & ~x54 ;
  assign n497 = ~x4 & x19 ;
  assign n498 = ~x21 & n497 ;
  assign n499 = n295 & n498 ;
  assign n500 = n342 & n499 ;
  assign n501 = n339 & n500 ;
  assign n502 = ~n496 & ~n501 ;
  assign n503 = n202 & ~n502 ;
  assign n504 = x22 & ~x54 ;
  assign n505 = x5 & ~x6 ;
  assign n506 = ~x14 & n505 ;
  assign n507 = n157 & n228 ;
  assign n508 = n506 & n507 ;
  assign n509 = n340 & n508 ;
  assign n510 = n358 & n509 ;
  assign n511 = ~n504 & ~n510 ;
  assign n512 = n202 & ~n511 ;
  assign n513 = ~x23 & x55 ;
  assign n514 = x61 & ~x129 ;
  assign n515 = ~n513 & n514 ;
  assign n520 = n243 & n422 ;
  assign n525 = x24 & x82 ;
  assign n526 = n468 & n525 ;
  assign n527 = n470 & n526 ;
  assign n528 = n520 & n527 ;
  assign n529 = ~x129 & ~n528 ;
  assign n516 = ~x2 & n249 ;
  assign n530 = ~x45 & ~x49 ;
  assign n531 = n247 & n530 ;
  assign n532 = n516 & n531 ;
  assign n533 = n246 & n532 ;
  assign n534 = x63 & ~n254 ;
  assign n535 = x82 & n534 ;
  assign n542 = ~n533 & n535 ;
  assign n543 = n542 ^ n534 ;
  assign n544 = n529 & ~n543 ;
  assign n517 = ~x49 & n516 ;
  assign n518 = x82 & ~n517 ;
  assign n519 = n254 & ~n518 ;
  assign n521 = n242 & n244 ;
  assign n522 = n520 & n521 ;
  assign n523 = x82 & ~n522 ;
  assign n524 = ~n519 & ~n523 ;
  assign n538 = ~x24 & ~n534 ;
  assign n536 = ~x24 & n535 ;
  assign n537 = ~n533 & n536 ;
  assign n539 = n538 ^ n537 ;
  assign n540 = n529 & n539 ;
  assign n541 = ~n524 & n540 ;
  assign n545 = n544 ^ n541 ;
  assign n586 = ~x53 & ~x58 ;
  assign n587 = ~x27 & ~x85 ;
  assign n581 = x25 & ~x116 ;
  assign n588 = ~x26 & n581 ;
  assign n589 = n587 & n588 ;
  assign n590 = ~n586 & ~n589 ;
  assign n591 = n202 & ~n590 ;
  assign n592 = x58 ^ x53 ;
  assign n596 = n591 & n592 ;
  assign n566 = ~x51 & ~x52 ;
  assign n567 = ~x39 & n566 ;
  assign n568 = x27 & ~n567 ;
  assign n569 = ~x95 & ~x100 ;
  assign n570 = ~x97 & ~x110 ;
  assign n571 = n569 & n570 ;
  assign n572 = n571 ^ x110 ;
  assign n573 = x25 & n572 ;
  assign n574 = ~n568 & n573 ;
  assign n575 = ~x26 & ~x85 ;
  assign n579 = x27 & n575 ;
  assign n580 = ~n574 & n579 ;
  assign n557 = x85 & x100 ;
  assign n558 = x116 & n557 ;
  assign n554 = ~x85 & ~x96 ;
  assign n555 = x100 & ~x110 ;
  assign n556 = n554 & n555 ;
  assign n559 = n558 ^ n556 ;
  assign n560 = x85 & ~x116 ;
  assign n561 = x25 & n560 ;
  assign n562 = ~n559 & ~n561 ;
  assign n563 = ~x26 & ~x27 ;
  assign n564 = ~n562 & n563 ;
  assign n546 = ~x39 & ~x52 ;
  assign n547 = ~x51 & x116 ;
  assign n548 = n546 & n547 ;
  assign n549 = ~x85 & ~n548 ;
  assign n550 = ~x25 & ~x116 ;
  assign n551 = x26 & ~x27 ;
  assign n552 = ~n550 & n551 ;
  assign n553 = n549 & n552 ;
  assign n565 = n564 ^ n553 ;
  assign n582 = ~n548 & ~n581 ;
  assign n583 = ~n565 & ~n582 ;
  assign n584 = n580 & n583 ;
  assign n576 = n574 & n575 ;
  assign n577 = ~n565 & n576 ;
  assign n578 = n577 ^ n565 ;
  assign n585 = n584 ^ n578 ;
  assign n593 = ~x53 & ~n592 ;
  assign n594 = n591 & n593 ;
  assign n595 = n585 & n594 ;
  assign n597 = n596 ^ n595 ;
  assign n598 = x26 & ~x85 ;
  assign n599 = ~n548 & n598 ;
  assign n600 = x26 & x116 ;
  assign n601 = n559 & ~n600 ;
  assign n602 = ~n599 & ~n601 ;
  assign n603 = ~x27 & ~x53 ;
  assign n604 = ~x58 & n603 ;
  assign n605 = n202 & n604 ;
  assign n606 = ~n602 & n605 ;
  assign n607 = x27 & n549 ;
  assign n608 = x85 & x116 ;
  assign n609 = ~x85 & ~x110 ;
  assign n610 = x95 & ~x96 ;
  assign n611 = n609 & n610 ;
  assign n612 = ~n608 & ~n611 ;
  assign n613 = ~x27 & ~x100 ;
  assign n614 = ~n612 & n613 ;
  assign n615 = ~n607 & ~n614 ;
  assign n616 = ~x26 & n202 ;
  assign n617 = n586 & n616 ;
  assign n618 = ~n615 & n617 ;
  assign n628 = ~x51 & n546 ;
  assign n629 = n600 & n628 ;
  assign n632 = ~x26 & ~x100 ;
  assign n633 = ~x110 & n632 ;
  assign n634 = n587 & n610 ;
  assign n635 = n633 & n634 ;
  assign n636 = ~n629 & n635 ;
  assign n630 = n587 & n629 ;
  assign n631 = n630 ^ x85 ;
  assign n637 = n636 ^ n631 ;
  assign n638 = ~x26 & x116 ;
  assign n639 = n568 & n638 ;
  assign n640 = ~n637 & n639 ;
  assign n641 = n640 ^ n637 ;
  assign n645 = ~x26 & ~x39 ;
  assign n646 = n566 & n645 ;
  assign n642 = ~x27 & ~x39 ;
  assign n643 = n566 & n642 ;
  assign n644 = n643 ^ x26 ;
  assign n647 = n646 ^ n644 ;
  assign n648 = n572 & ~n647 ;
  assign n649 = x27 ^ x26 ;
  assign n650 = ~x116 & n649 ;
  assign n651 = x28 & ~n650 ;
  assign n652 = ~n648 & n651 ;
  assign n653 = n652 ^ x28 ;
  assign n654 = x100 & x116 ;
  assign n655 = ~x28 & ~x116 ;
  assign n656 = n563 & ~n655 ;
  assign n657 = ~n654 & n656 ;
  assign n662 = ~x53 & ~x85 ;
  assign n663 = ~n657 & n662 ;
  assign n664 = ~n653 & n663 ;
  assign n665 = ~n641 & n664 ;
  assign n666 = n665 ^ n663 ;
  assign n658 = ~x53 & n657 ;
  assign n659 = ~n653 & n658 ;
  assign n660 = ~n641 & n659 ;
  assign n661 = n660 ^ n658 ;
  assign n667 = n666 ^ n661 ;
  assign n619 = ~x26 & ~x53 ;
  assign n620 = ~x85 & n619 ;
  assign n621 = ~x27 & x28 ;
  assign n622 = ~x116 & n621 ;
  assign n623 = x58 & n622 ;
  assign n624 = n620 & n623 ;
  assign n668 = ~x58 & n202 ;
  assign n669 = x53 & n575 ;
  assign n670 = n622 & n669 ;
  assign n671 = n668 & ~n670 ;
  assign n672 = ~n624 & n671 ;
  assign n673 = ~n667 & n672 ;
  assign n625 = x58 & n202 ;
  assign n626 = ~n624 & n625 ;
  assign n627 = n626 ^ n202 ;
  assign n674 = n673 ^ n627 ;
  assign n675 = x29 & ~x116 ;
  assign n696 = x53 & ~x58 ;
  assign n697 = n675 & n696 ;
  assign n701 = ~x27 & n697 ;
  assign n682 = ~x96 & ~x110 ;
  assign n683 = x97 & ~n682 ;
  assign n684 = x29 & ~x110 ;
  assign n685 = n569 & n684 ;
  assign n686 = ~n683 & n685 ;
  assign n681 = x29 & x110 ;
  assign n687 = n686 ^ n681 ;
  assign n688 = ~x58 & x97 ;
  assign n689 = n569 & n688 ;
  assign n690 = ~n683 & n689 ;
  assign n691 = n690 ^ x58 ;
  assign n692 = ~n687 & ~n691 ;
  assign n693 = x97 & x116 ;
  assign n694 = x58 & ~n675 ;
  assign n695 = ~n693 & n694 ;
  assign n698 = n603 & ~n697 ;
  assign n699 = ~n695 & n698 ;
  assign n700 = ~n692 & n699 ;
  assign n702 = n701 ^ n700 ;
  assign n676 = x85 & n675 ;
  assign n677 = n604 & n676 ;
  assign n703 = x27 & n586 ;
  assign n704 = n675 & n703 ;
  assign n705 = n575 & ~n704 ;
  assign n706 = ~n677 & n705 ;
  assign n707 = ~n702 & n706 ;
  assign n678 = ~x26 & x85 ;
  assign n679 = ~n677 & n678 ;
  assign n680 = n679 ^ x26 ;
  assign n708 = n707 ^ n680 ;
  assign n709 = ~x85 & n586 ;
  assign n710 = n551 & n709 ;
  assign n711 = n675 & n710 ;
  assign n712 = n202 & ~n711 ;
  assign n713 = n708 & n712 ;
  assign n714 = n713 ^ n202 ;
  assign n715 = ~x30 & ~x109 ;
  assign n716 = ~x60 & x109 ;
  assign n717 = ~n715 & ~n716 ;
  assign n718 = ~x106 & ~n717 ;
  assign n719 = ~x88 & x106 ;
  assign n720 = ~x129 & ~n719 ;
  assign n721 = ~n718 & n720 ;
  assign n722 = ~x31 & ~x109 ;
  assign n723 = ~x30 & x109 ;
  assign n724 = ~n722 & ~n723 ;
  assign n725 = ~x106 & ~n724 ;
  assign n726 = ~x89 & x106 ;
  assign n727 = ~x129 & ~n726 ;
  assign n728 = ~n725 & n727 ;
  assign n729 = ~x32 & ~x109 ;
  assign n730 = ~x31 & x109 ;
  assign n731 = ~n729 & ~n730 ;
  assign n732 = ~x106 & ~n731 ;
  assign n733 = ~x99 & x106 ;
  assign n734 = ~x129 & ~n733 ;
  assign n735 = ~n732 & n734 ;
  assign n736 = ~x33 & ~x109 ;
  assign n737 = ~x32 & x109 ;
  assign n738 = ~n736 & ~n737 ;
  assign n739 = ~x106 & ~n738 ;
  assign n740 = ~x90 & x106 ;
  assign n741 = ~x129 & ~n740 ;
  assign n742 = ~n739 & n741 ;
  assign n743 = ~x34 & ~x109 ;
  assign n744 = ~x33 & x109 ;
  assign n745 = ~n743 & ~n744 ;
  assign n746 = ~x106 & ~n745 ;
  assign n747 = ~x91 & x106 ;
  assign n748 = ~x129 & ~n747 ;
  assign n749 = ~n746 & n748 ;
  assign n750 = ~x35 & ~x109 ;
  assign n751 = ~x34 & x109 ;
  assign n752 = ~n750 & ~n751 ;
  assign n753 = ~x106 & ~n752 ;
  assign n754 = ~x92 & x106 ;
  assign n755 = ~x129 & ~n754 ;
  assign n756 = ~n753 & n755 ;
  assign n757 = ~x36 & ~x109 ;
  assign n758 = ~x35 & x109 ;
  assign n759 = ~n757 & ~n758 ;
  assign n760 = ~x106 & ~n759 ;
  assign n761 = ~x98 & x106 ;
  assign n762 = ~x129 & ~n761 ;
  assign n763 = ~n760 & n762 ;
  assign n764 = ~x37 & ~x109 ;
  assign n765 = ~x36 & x109 ;
  assign n766 = ~n764 & ~n765 ;
  assign n767 = ~x106 & ~n766 ;
  assign n768 = ~x93 & x106 ;
  assign n769 = ~x129 & ~n768 ;
  assign n770 = ~n767 & n769 ;
  assign n773 = ~x45 & ~x50 ;
  assign n774 = n251 & n773 ;
  assign n775 = n516 & n774 ;
  assign n776 = x82 & n265 ;
  assign n777 = n417 & n776 ;
  assign n778 = n775 & n777 ;
  assign n779 = n778 ^ x82 ;
  assign n771 = x82 & ~n272 ;
  assign n780 = ~x38 & n254 ;
  assign n781 = ~n771 & n780 ;
  assign n782 = ~n779 & n781 ;
  assign n772 = ~x38 & n771 ;
  assign n783 = n782 ^ n772 ;
  assign n792 = ~x44 & x82 ;
  assign n793 = ~x40 & ~x42 ;
  assign n794 = x38 & n793 ;
  assign n795 = n792 & n794 ;
  assign n796 = x74 & ~n254 ;
  assign n800 = ~x129 & ~n796 ;
  assign n801 = ~n795 & n800 ;
  assign n784 = ~x45 & ~x48 ;
  assign n785 = n251 & n784 ;
  assign n786 = n516 & n785 ;
  assign n787 = n265 & n267 ;
  assign n788 = ~x40 & ~x50 ;
  assign n789 = n244 & n788 ;
  assign n790 = n787 & n789 ;
  assign n791 = n786 & n790 ;
  assign n797 = n428 & n796 ;
  assign n798 = ~n795 & n797 ;
  assign n799 = ~n791 & n798 ;
  assign n802 = n801 ^ n799 ;
  assign n803 = ~n783 & n802 ;
  assign n804 = x109 & n566 ;
  assign n805 = x39 & ~n804 ;
  assign n806 = ~x51 & x109 ;
  assign n807 = n546 & n806 ;
  assign n808 = ~x106 & ~n807 ;
  assign n809 = ~n805 & n808 ;
  assign n810 = ~x129 & ~n809 ;
  assign n813 = n253 & n270 ;
  assign n814 = n813 ^ x82 ;
  assign n811 = x82 & ~n244 ;
  assign n815 = ~x40 & n254 ;
  assign n816 = ~n811 & n815 ;
  assign n817 = ~n814 & n816 ;
  assign n812 = ~x40 & n811 ;
  assign n818 = n817 ^ n812 ;
  assign n819 = ~x42 & n792 ;
  assign n820 = x40 & n819 ;
  assign n821 = ~x129 & ~n820 ;
  assign n822 = ~n818 & n821 ;
  assign n825 = ~x46 & n240 ;
  assign n826 = n243 & n825 ;
  assign n827 = ~x2 & ~x45 ;
  assign n828 = n251 & n827 ;
  assign n829 = n247 & n249 ;
  assign n830 = n828 & n829 ;
  assign n831 = n826 & n830 ;
  assign n832 = n244 & n831 ;
  assign n823 = x73 & ~n254 ;
  assign n833 = x82 & n823 ;
  assign n834 = ~n832 & n833 ;
  assign n835 = n822 & n834 ;
  assign n824 = n822 & ~n823 ;
  assign n836 = n835 ^ n824 ;
  assign n837 = x82 & n254 ;
  assign n838 = n269 & n837 ;
  assign n839 = n264 & n838 ;
  assign n840 = n839 ^ n408 ;
  assign n842 = ~x41 & x82 ;
  assign n843 = ~n521 & n842 ;
  assign n844 = ~n840 & n843 ;
  assign n841 = ~x41 & n840 ;
  assign n845 = n844 ^ n841 ;
  assign n846 = x41 & n819 ;
  assign n847 = n242 & n846 ;
  assign n848 = ~x129 & ~n847 ;
  assign n849 = ~n845 & n848 ;
  assign n852 = n264 & n269 ;
  assign n853 = n471 & n852 ;
  assign n850 = x76 & ~n254 ;
  assign n854 = x82 & n850 ;
  assign n855 = ~n853 & n854 ;
  assign n856 = n849 & n855 ;
  assign n851 = n849 & ~n850 ;
  assign n857 = n856 ^ n851 ;
  assign n863 = ~x40 & x82 ;
  assign n864 = n243 & n863 ;
  assign n865 = n825 & n864 ;
  assign n866 = n830 & n865 ;
  assign n867 = n866 ^ x82 ;
  assign n861 = x44 & x82 ;
  assign n868 = ~x42 & n254 ;
  assign n869 = ~n861 & n868 ;
  assign n870 = ~n867 & n869 ;
  assign n862 = ~x42 & n861 ;
  assign n871 = n870 ^ n862 ;
  assign n872 = x42 & n792 ;
  assign n873 = ~x129 & ~n872 ;
  assign n878 = ~x72 & n873 ;
  assign n879 = ~n871 & n878 ;
  assign n858 = n243 & n793 ;
  assign n859 = n825 & n858 ;
  assign n860 = n830 & n859 ;
  assign n874 = x72 & ~n255 ;
  assign n875 = n873 & n874 ;
  assign n876 = ~n871 & n875 ;
  assign n877 = ~n860 & n876 ;
  assign n880 = n879 ^ n877 ;
  assign n881 = n415 & n830 ;
  assign n882 = x82 & ~n881 ;
  assign n883 = x77 & ~n254 ;
  assign n884 = ~n882 & n883 ;
  assign n885 = n251 & n423 ;
  assign n886 = n247 & n401 ;
  assign n887 = n885 & n886 ;
  assign n889 = n408 & ~n887 ;
  assign n888 = n254 & n887 ;
  assign n890 = n889 ^ n888 ;
  assign n892 = ~x43 & x82 ;
  assign n893 = ~n415 & n892 ;
  assign n894 = ~n890 & n893 ;
  assign n891 = ~x43 & n890 ;
  assign n895 = n894 ^ n891 ;
  assign n896 = n792 & n793 ;
  assign n897 = n266 & n896 ;
  assign n898 = x43 & n897 ;
  assign n899 = ~x129 & ~n898 ;
  assign n900 = ~n895 & n899 ;
  assign n901 = ~n884 & n900 ;
  assign n902 = ~x67 & ~n254 ;
  assign n903 = x44 & n254 ;
  assign n904 = ~n902 & ~n903 ;
  assign n905 = ~x129 & ~n861 ;
  assign n907 = x82 & n905 ;
  assign n908 = n904 & n907 ;
  assign n909 = ~n860 & n908 ;
  assign n906 = ~n904 & n905 ;
  assign n910 = n909 ^ n906 ;
  assign n911 = ~x50 & n470 ;
  assign n912 = n777 & n911 ;
  assign n913 = n912 ^ x82 ;
  assign n914 = n254 & n423 ;
  assign n915 = n251 & n479 ;
  assign n916 = n914 & n915 ;
  assign n917 = n916 ^ n408 ;
  assign n918 = ~x45 & ~n917 ;
  assign n919 = ~n913 & n918 ;
  assign n920 = n919 ^ x45 ;
  assign n921 = n247 & n423 ;
  assign n922 = n421 & n921 ;
  assign n923 = n246 & n922 ;
  assign n924 = x68 & ~n254 ;
  assign n925 = x82 & n924 ;
  assign n926 = ~n923 & n925 ;
  assign n927 = n926 ^ n924 ;
  assign n928 = n265 & n417 ;
  assign n929 = x45 & x82 ;
  assign n930 = ~x50 & ~x129 ;
  assign n931 = n929 & n930 ;
  assign n932 = n470 & n931 ;
  assign n933 = n928 & n932 ;
  assign n934 = n933 ^ x129 ;
  assign n935 = ~n927 & ~n934 ;
  assign n936 = n920 & n935 ;
  assign n938 = ~x75 & ~n254 ;
  assign n941 = ~x82 & ~n938 ;
  assign n937 = x82 & n243 ;
  assign n939 = n937 & ~n938 ;
  assign n940 = n830 & n939 ;
  assign n942 = n941 ^ n940 ;
  assign n943 = n471 & ~n942 ;
  assign n945 = ~x75 & n255 ;
  assign n950 = ~n943 & ~n945 ;
  assign n944 = x82 & n911 ;
  assign n946 = x46 & ~n255 ;
  assign n947 = ~n945 & n946 ;
  assign n948 = ~n944 & n947 ;
  assign n949 = ~n943 & n948 ;
  assign n951 = n950 ^ n949 ;
  assign n952 = ~x129 & ~n951 ;
  assign n954 = n408 & ~n786 ;
  assign n953 = n254 & n786 ;
  assign n955 = n954 ^ n953 ;
  assign n957 = ~x47 & x82 ;
  assign n958 = ~n246 & n957 ;
  assign n959 = ~n955 & n958 ;
  assign n956 = ~x47 & n955 ;
  assign n960 = n959 ^ n956 ;
  assign n961 = ~x43 & x47 ;
  assign n962 = n897 & n961 ;
  assign n963 = ~x129 & ~n962 ;
  assign n964 = ~n960 & n963 ;
  assign n967 = n246 & n786 ;
  assign n965 = x64 & ~n254 ;
  assign n968 = x82 & n965 ;
  assign n969 = ~n967 & n968 ;
  assign n970 = n964 & n969 ;
  assign n966 = n964 & ~n965 ;
  assign n971 = n970 ^ n966 ;
  assign n972 = x82 & n787 ;
  assign n973 = n911 & n972 ;
  assign n974 = n973 ^ x82 ;
  assign n976 = ~x45 & x82 ;
  assign n977 = n251 & n976 ;
  assign n978 = n516 & n977 ;
  assign n979 = n978 ^ x82 ;
  assign n980 = ~x48 & n254 ;
  assign n981 = ~n979 & n980 ;
  assign n982 = ~n974 & n981 ;
  assign n975 = ~x48 & n974 ;
  assign n983 = n982 ^ n975 ;
  assign n984 = x48 & n267 ;
  assign n985 = n897 & n984 ;
  assign n986 = ~x129 & ~n985 ;
  assign n987 = ~n983 & n986 ;
  assign n990 = n416 & n516 ;
  assign n991 = ~x47 & n246 ;
  assign n992 = n990 & n991 ;
  assign n988 = x62 & ~n254 ;
  assign n993 = x82 & n988 ;
  assign n994 = ~n992 & n993 ;
  assign n995 = n987 & n994 ;
  assign n989 = n987 & ~n988 ;
  assign n996 = n995 ^ n989 ;
  assign n997 = n474 & ~n516 ;
  assign n998 = ~x24 & ~x40 ;
  assign n999 = n244 & n998 ;
  assign n1000 = n825 & n999 ;
  assign n1001 = x49 & n243 ;
  assign n1002 = n422 & n1001 ;
  assign n1003 = n1000 & n1002 ;
  assign n1004 = n1003 ^ x49 ;
  assign n1005 = x82 & ~n1004 ;
  assign n1006 = ~n997 & n1005 ;
  assign n1007 = n1006 ^ x82 ;
  assign n1008 = x82 & n468 ;
  assign n1009 = n470 & n1008 ;
  assign n1010 = n473 & n1009 ;
  assign n1011 = n1010 ^ x82 ;
  assign n1012 = x49 & n408 ;
  assign n1013 = ~x69 & ~n254 ;
  assign n1014 = ~n1012 & n1013 ;
  assign n1015 = ~n1011 & n1014 ;
  assign n1016 = n1015 ^ n1012 ;
  assign n1017 = ~x129 & ~n1016 ;
  assign n1018 = ~n1007 & n1017 ;
  assign n1019 = n1018 ^ x129 ;
  assign n1025 = n269 & n776 ;
  assign n1026 = n264 & n1025 ;
  assign n1027 = n1026 ^ x82 ;
  assign n1023 = x82 & ~n470 ;
  assign n1028 = ~x50 & n254 ;
  assign n1029 = ~n1023 & n1028 ;
  assign n1030 = ~n1027 & n1029 ;
  assign n1024 = ~x50 & n1023 ;
  assign n1031 = n1030 ^ n1024 ;
  assign n1032 = x50 & x82 ;
  assign n1033 = n470 & n1032 ;
  assign n1034 = ~x129 & ~n1033 ;
  assign n1039 = ~n1031 & n1034 ;
  assign n1020 = ~x50 & n787 ;
  assign n1021 = n786 & n1020 ;
  assign n1022 = x82 & ~n1021 ;
  assign n1035 = x66 & ~n254 ;
  assign n1036 = n1034 & n1035 ;
  assign n1037 = ~n1031 & n1036 ;
  assign n1038 = ~n1022 & n1037 ;
  assign n1040 = n1039 ^ n1038 ;
  assign n1041 = x51 & ~x109 ;
  assign n1042 = ~x106 & ~n806 ;
  assign n1043 = ~n1041 & n1042 ;
  assign n1044 = ~x129 & ~n1043 ;
  assign n1045 = x52 & ~n806 ;
  assign n1046 = ~x106 & ~n804 ;
  assign n1047 = ~n1045 & n1046 ;
  assign n1048 = ~x129 & ~n1047 ;
  assign n1049 = ~x116 & n696 ;
  assign n1050 = ~x53 & x97 ;
  assign n1051 = x58 & x116 ;
  assign n1052 = ~x58 & n569 ;
  assign n1053 = n682 & n1052 ;
  assign n1054 = ~n1051 & ~n1053 ;
  assign n1055 = n1050 & ~n1054 ;
  assign n1056 = ~n1049 & ~n1055 ;
  assign n1057 = n587 & n616 ;
  assign n1058 = ~n1056 & n1057 ;
  assign n1059 = n421 & n423 ;
  assign n1060 = ~n254 & n1059 ;
  assign n1061 = n522 & n1060 ;
  assign n1062 = ~x129 & ~n255 ;
  assign n1063 = ~n1061 & n1062 ;
  assign n1064 = ~x123 & ~x129 ;
  assign n1065 = x114 & ~x122 ;
  assign n1066 = n1064 & n1065 ;
  assign n1078 = ~x26 & x37 ;
  assign n1092 = n703 & n1078 ;
  assign n1073 = ~x26 & x58 ;
  assign n1074 = ~x94 & ~x116 ;
  assign n1075 = n1073 & n1074 ;
  assign n1076 = n1075 ^ n1073 ;
  assign n1069 = x26 & ~x58 ;
  assign n1070 = x94 & x116 ;
  assign n1071 = n1069 & n1070 ;
  assign n1067 = x37 & ~x58 ;
  assign n1068 = ~x116 & n1067 ;
  assign n1072 = n1071 ^ n1068 ;
  assign n1077 = n1076 ^ n1072 ;
  assign n1083 = ~x53 & n1077 ;
  assign n1081 = ~x58 & n1078 ;
  assign n1079 = n586 & n1078 ;
  assign n1080 = n1077 & n1079 ;
  assign n1082 = n1081 ^ n1080 ;
  assign n1084 = n1083 ^ n1082 ;
  assign n1089 = n587 & n1078 ;
  assign n1090 = n586 & n1089 ;
  assign n1091 = ~n1084 & n1090 ;
  assign n1093 = n1092 ^ n1091 ;
  assign n1086 = x85 & n586 ;
  assign n1087 = n1078 & n1086 ;
  assign n1085 = n587 & n1084 ;
  assign n1088 = n1087 ^ n1085 ;
  assign n1094 = n1093 ^ n1088 ;
  assign n1095 = n202 & n1094 ;
  assign n1101 = x26 & ~x53 ;
  assign n1102 = ~x58 & n1101 ;
  assign n1099 = ~x26 & ~x58 ;
  assign n1100 = ~x85 & n1099 ;
  assign n1103 = n1102 ^ n1100 ;
  assign n1104 = n1103 ^ n1086 ;
  assign n1113 = x57 & ~n620 ;
  assign n1114 = n1104 & n1113 ;
  assign n1115 = n1114 ^ n620 ;
  assign n1107 = x60 & n1051 ;
  assign n1110 = ~x57 & n620 ;
  assign n1111 = ~n1107 & n1110 ;
  assign n1105 = x57 & x116 ;
  assign n1106 = ~n1104 & n1105 ;
  assign n1108 = n620 & ~n1107 ;
  assign n1109 = n1106 & n1108 ;
  assign n1112 = n1111 ^ n1109 ;
  assign n1116 = n1115 ^ n1112 ;
  assign n1096 = x57 & ~x58 ;
  assign n1097 = n620 & n1096 ;
  assign n1117 = ~x27 & n202 ;
  assign n1118 = ~n1097 & n1117 ;
  assign n1119 = n1116 & n1118 ;
  assign n1098 = n202 & n1097 ;
  assign n1120 = n1119 ^ n1098 ;
  assign n1121 = x58 & ~x116 ;
  assign n1122 = n563 & n1121 ;
  assign n1123 = ~x58 & n649 ;
  assign n1124 = n548 & n1123 ;
  assign n1125 = ~n1122 & ~n1124 ;
  assign n1126 = n202 & n662 ;
  assign n1127 = ~n1125 & n1126 ;
  assign n1128 = x59 & ~x116 ;
  assign n1144 = x27 & n1128 ;
  assign n1145 = n709 & n1144 ;
  assign n1135 = x96 & n586 ;
  assign n1136 = ~n572 & n1135 ;
  assign n1133 = x59 & n586 ;
  assign n1134 = n572 & n1133 ;
  assign n1137 = n1136 ^ n1134 ;
  assign n1138 = n592 & n1128 ;
  assign n1139 = ~x85 & ~n1138 ;
  assign n1140 = ~n1137 & n1139 ;
  assign n1131 = n1086 & n1128 ;
  assign n1132 = n1131 ^ x85 ;
  assign n1141 = n1140 ^ n1132 ;
  assign n1142 = n563 & ~n1141 ;
  assign n1129 = x26 & n1128 ;
  assign n1130 = n709 & n1129 ;
  assign n1143 = n1142 ^ n1130 ;
  assign n1146 = n1145 ^ n1143 ;
  assign n1147 = n202 & n1146 ;
  assign n1148 = ~x117 & ~x122 ;
  assign n1149 = x60 & ~n1148 ;
  assign n1150 = x123 & n1148 ;
  assign n1151 = ~n1149 & ~n1150 ;
  assign n1152 = ~x114 & ~x122 ;
  assign n1153 = x123 & ~x129 ;
  assign n1154 = n1152 & n1153 ;
  assign n1155 = x136 & ~x137 ;
  assign n1156 = x131 & x132 ;
  assign n1157 = x133 & n1156 ;
  assign n1158 = ~x138 & n1157 ;
  assign n1159 = n1155 & n1158 ;
  assign n1160 = x140 & n1159 ;
  assign n1161 = ~x62 & ~n1159 ;
  assign n1162 = ~x129 & ~n1161 ;
  assign n1163 = ~n1160 & n1162 ;
  assign n1164 = x142 & n1159 ;
  assign n1165 = ~x63 & ~n1159 ;
  assign n1166 = ~x129 & ~n1165 ;
  assign n1167 = ~n1164 & n1166 ;
  assign n1168 = x139 & n1159 ;
  assign n1169 = ~x64 & ~n1159 ;
  assign n1170 = ~x129 & ~n1169 ;
  assign n1171 = ~n1168 & n1170 ;
  assign n1172 = x146 & n1159 ;
  assign n1173 = ~x65 & ~n1159 ;
  assign n1174 = ~x129 & ~n1173 ;
  assign n1175 = ~n1172 & n1174 ;
  assign n1176 = ~x136 & ~x137 ;
  assign n1177 = n1158 & n1176 ;
  assign n1178 = x143 & n1177 ;
  assign n1179 = ~x66 & ~n1177 ;
  assign n1180 = ~x129 & ~n1179 ;
  assign n1181 = ~n1178 & n1180 ;
  assign n1182 = x139 & n1177 ;
  assign n1183 = ~x67 & ~n1177 ;
  assign n1184 = ~x129 & ~n1183 ;
  assign n1185 = ~n1182 & n1184 ;
  assign n1186 = x141 & n1159 ;
  assign n1187 = ~x68 & ~n1159 ;
  assign n1188 = ~x129 & ~n1187 ;
  assign n1189 = ~n1186 & n1188 ;
  assign n1190 = x143 & n1159 ;
  assign n1191 = ~x69 & ~n1159 ;
  assign n1192 = ~x129 & ~n1191 ;
  assign n1193 = ~n1190 & n1192 ;
  assign n1194 = x144 & n1159 ;
  assign n1195 = ~x70 & ~n1159 ;
  assign n1196 = ~x129 & ~n1195 ;
  assign n1197 = ~n1194 & n1196 ;
  assign n1198 = x145 & n1159 ;
  assign n1199 = ~x71 & ~n1159 ;
  assign n1200 = ~x129 & ~n1199 ;
  assign n1201 = ~n1198 & n1200 ;
  assign n1202 = x140 & n1177 ;
  assign n1203 = ~x72 & ~n1177 ;
  assign n1204 = ~x129 & ~n1203 ;
  assign n1205 = ~n1202 & n1204 ;
  assign n1206 = x141 & n1177 ;
  assign n1207 = ~x73 & ~n1177 ;
  assign n1208 = ~x129 & ~n1207 ;
  assign n1209 = ~n1206 & n1208 ;
  assign n1210 = x142 & n1177 ;
  assign n1211 = ~x74 & ~n1177 ;
  assign n1212 = ~x129 & ~n1211 ;
  assign n1213 = ~n1210 & n1212 ;
  assign n1214 = x144 & n1177 ;
  assign n1215 = ~x75 & ~n1177 ;
  assign n1216 = ~x129 & ~n1215 ;
  assign n1217 = ~n1214 & n1216 ;
  assign n1218 = x145 & n1177 ;
  assign n1219 = ~x76 & ~n1177 ;
  assign n1220 = ~x129 & ~n1219 ;
  assign n1221 = ~n1218 & n1220 ;
  assign n1222 = x146 & n1177 ;
  assign n1223 = ~x77 & ~n1177 ;
  assign n1224 = ~x129 & ~n1223 ;
  assign n1225 = ~n1222 & n1224 ;
  assign n1226 = ~x136 & x137 ;
  assign n1227 = n1158 & n1226 ;
  assign n1228 = ~x142 & n1227 ;
  assign n1229 = ~x78 & ~n1227 ;
  assign n1230 = ~x129 & ~n1229 ;
  assign n1231 = ~n1228 & n1230 ;
  assign n1232 = ~x143 & n1227 ;
  assign n1233 = ~x79 & ~n1227 ;
  assign n1234 = ~x129 & ~n1233 ;
  assign n1235 = ~n1232 & n1234 ;
  assign n1236 = ~x144 & n1227 ;
  assign n1237 = ~x80 & ~n1227 ;
  assign n1238 = ~x129 & ~n1237 ;
  assign n1239 = ~n1236 & n1238 ;
  assign n1240 = ~x145 & n1227 ;
  assign n1241 = ~x81 & ~n1227 ;
  assign n1242 = ~x129 & ~n1241 ;
  assign n1243 = ~n1240 & n1242 ;
  assign n1244 = ~x146 & n1227 ;
  assign n1245 = ~x82 & ~n1227 ;
  assign n1246 = ~x129 & ~n1245 ;
  assign n1247 = ~n1244 & n1246 ;
  assign n1248 = x136 & ~x138 ;
  assign n1249 = x31 & n1248 ;
  assign n1250 = x115 & x138 ;
  assign n1251 = ~x87 & ~x138 ;
  assign n1252 = ~x136 & ~n1251 ;
  assign n1253 = ~n1250 & n1252 ;
  assign n1254 = ~n1249 & ~n1253 ;
  assign n1255 = x137 & ~n1254 ;
  assign n1256 = x62 & ~x138 ;
  assign n1257 = ~x89 & x138 ;
  assign n1258 = x136 & ~n1257 ;
  assign n1259 = ~n1256 & n1258 ;
  assign n1260 = x72 & ~x138 ;
  assign n1261 = ~x119 & x138 ;
  assign n1262 = ~x136 & ~n1261 ;
  assign n1263 = ~n1260 & n1262 ;
  assign n1264 = ~n1259 & ~n1263 ;
  assign n1265 = ~x137 & ~n1264 ;
  assign n1266 = ~n1255 & ~n1265 ;
  assign n1267 = ~x141 & n1227 ;
  assign n1268 = ~x84 & ~n1227 ;
  assign n1269 = ~x129 & ~n1268 ;
  assign n1270 = ~n1267 & n1269 ;
  assign n1271 = ~x97 & n569 ;
  assign n1272 = n609 & ~n1271 ;
  assign n1273 = x96 & n1272 ;
  assign n1274 = ~n560 & ~n1273 ;
  assign n1275 = n604 & n616 ;
  assign n1276 = ~n1274 & n1275 ;
  assign n1277 = ~x139 & n1227 ;
  assign n1278 = ~x86 & ~n1227 ;
  assign n1279 = ~x129 & ~n1278 ;
  assign n1280 = ~n1277 & n1279 ;
  assign n1281 = ~x140 & n1227 ;
  assign n1282 = ~x87 & ~n1227 ;
  assign n1283 = ~x129 & ~n1282 ;
  assign n1284 = ~n1281 & n1283 ;
  assign n1285 = x137 & n1248 ;
  assign n1286 = n1157 & n1285 ;
  assign n1287 = ~x139 & n1286 ;
  assign n1288 = ~x88 & ~n1286 ;
  assign n1289 = ~x129 & ~n1288 ;
  assign n1290 = ~n1287 & n1289 ;
  assign n1291 = ~x140 & n1286 ;
  assign n1292 = ~x89 & ~n1286 ;
  assign n1293 = ~x129 & ~n1292 ;
  assign n1294 = ~n1291 & n1293 ;
  assign n1295 = ~x142 & n1286 ;
  assign n1296 = ~x90 & ~n1286 ;
  assign n1297 = ~x129 & ~n1296 ;
  assign n1298 = ~n1295 & n1297 ;
  assign n1299 = ~x143 & n1286 ;
  assign n1300 = ~x91 & ~n1286 ;
  assign n1301 = ~x129 & ~n1300 ;
  assign n1302 = ~n1299 & n1301 ;
  assign n1303 = ~x144 & n1286 ;
  assign n1304 = ~x92 & ~n1286 ;
  assign n1305 = ~x129 & ~n1304 ;
  assign n1306 = ~n1303 & n1305 ;
  assign n1307 = ~x146 & n1286 ;
  assign n1308 = ~x93 & ~n1286 ;
  assign n1309 = ~x129 & ~n1308 ;
  assign n1310 = ~n1307 & n1309 ;
  assign n1311 = x82 & x138 ;
  assign n1312 = n1176 & n1311 ;
  assign n1313 = n1157 & n1312 ;
  assign n1314 = ~x142 & n1313 ;
  assign n1315 = ~x94 & ~n1313 ;
  assign n1316 = ~x129 & ~n1315 ;
  assign n1317 = ~n1314 & n1316 ;
  assign n1318 = ~x3 & ~x110 ;
  assign n1319 = ~n1157 & ~n1318 ;
  assign n1320 = ~n1313 & ~n1319 ;
  assign n1321 = x95 & n1320 ;
  assign n1322 = x143 & n1313 ;
  assign n1323 = ~n1321 & ~n1322 ;
  assign n1324 = ~x129 & ~n1323 ;
  assign n1325 = x96 & n1320 ;
  assign n1326 = x146 & n1313 ;
  assign n1327 = ~n1325 & ~n1326 ;
  assign n1328 = ~x129 & ~n1327 ;
  assign n1329 = x97 & n1320 ;
  assign n1330 = x145 & n1313 ;
  assign n1331 = ~n1329 & ~n1330 ;
  assign n1332 = ~x129 & ~n1331 ;
  assign n1333 = ~x145 & n1286 ;
  assign n1334 = ~x98 & ~n1286 ;
  assign n1335 = ~x129 & ~n1334 ;
  assign n1336 = ~n1333 & n1335 ;
  assign n1337 = ~x141 & n1286 ;
  assign n1338 = ~x99 & ~n1286 ;
  assign n1339 = ~x129 & ~n1338 ;
  assign n1340 = ~n1337 & n1339 ;
  assign n1341 = x100 & n1320 ;
  assign n1342 = x144 & n1313 ;
  assign n1343 = ~n1341 & ~n1342 ;
  assign n1344 = ~x129 & ~n1343 ;
  assign n1345 = x37 & n1248 ;
  assign n1346 = ~x96 & x138 ;
  assign n1347 = ~x82 & ~x138 ;
  assign n1348 = ~x136 & ~n1347 ;
  assign n1349 = ~n1346 & n1348 ;
  assign n1350 = ~n1345 & ~n1349 ;
  assign n1351 = x137 & ~n1350 ;
  assign n1352 = x65 & ~x138 ;
  assign n1353 = ~x93 & x138 ;
  assign n1354 = x136 & ~n1353 ;
  assign n1355 = ~n1352 & n1354 ;
  assign n1356 = x77 & ~x138 ;
  assign n1357 = ~x124 & x138 ;
  assign n1358 = ~x136 & ~n1357 ;
  assign n1359 = ~n1356 & n1358 ;
  assign n1360 = ~n1355 & ~n1359 ;
  assign n1361 = ~x137 & ~n1360 ;
  assign n1362 = ~n1351 & ~n1361 ;
  assign n1363 = x91 & n1155 ;
  assign n1364 = x95 & n1226 ;
  assign n1365 = ~n1363 & ~n1364 ;
  assign n1366 = x138 & ~n1365 ;
  assign n1367 = ~x34 & x136 ;
  assign n1368 = ~x79 & ~x136 ;
  assign n1369 = x137 & ~n1368 ;
  assign n1370 = ~n1367 & n1369 ;
  assign n1371 = x69 & x136 ;
  assign n1372 = x66 & ~x136 ;
  assign n1373 = ~x137 & ~n1372 ;
  assign n1374 = ~n1371 & n1373 ;
  assign n1375 = ~n1370 & ~n1374 ;
  assign n1376 = ~x138 & ~n1375 ;
  assign n1377 = ~n1366 & ~n1376 ;
  assign n1378 = x90 & n1155 ;
  assign n1379 = x94 & n1226 ;
  assign n1380 = ~n1378 & ~n1379 ;
  assign n1381 = x138 & ~n1380 ;
  assign n1382 = ~x33 & x136 ;
  assign n1383 = ~x78 & ~x136 ;
  assign n1384 = x137 & ~n1383 ;
  assign n1385 = ~n1382 & n1384 ;
  assign n1386 = x63 & x136 ;
  assign n1387 = x74 & ~x136 ;
  assign n1388 = ~x137 & ~n1387 ;
  assign n1389 = ~n1386 & n1388 ;
  assign n1390 = ~n1385 & ~n1389 ;
  assign n1391 = ~x138 & ~n1390 ;
  assign n1392 = ~n1381 & ~n1391 ;
  assign n1393 = x99 & n1155 ;
  assign n1394 = ~x112 & n1226 ;
  assign n1395 = ~n1393 & ~n1394 ;
  assign n1396 = x138 & ~n1395 ;
  assign n1397 = ~x32 & x136 ;
  assign n1398 = ~x84 & ~x136 ;
  assign n1399 = x137 & ~n1398 ;
  assign n1400 = ~n1397 & n1399 ;
  assign n1401 = x68 & x136 ;
  assign n1402 = x73 & ~x136 ;
  assign n1403 = ~x137 & ~n1402 ;
  assign n1404 = ~n1401 & n1403 ;
  assign n1405 = ~n1400 & ~n1404 ;
  assign n1406 = ~x138 & ~n1405 ;
  assign n1407 = ~n1396 & ~n1406 ;
  assign n1408 = x35 & n1248 ;
  assign n1409 = ~x100 & x138 ;
  assign n1410 = ~x80 & ~x138 ;
  assign n1411 = ~x136 & ~n1410 ;
  assign n1412 = ~n1409 & n1411 ;
  assign n1413 = ~n1408 & ~n1412 ;
  assign n1414 = x137 & ~n1413 ;
  assign n1415 = x70 & ~x138 ;
  assign n1416 = ~x92 & x138 ;
  assign n1417 = x136 & ~n1416 ;
  assign n1418 = ~n1415 & n1417 ;
  assign n1419 = x75 & ~x138 ;
  assign n1420 = ~x125 & x138 ;
  assign n1421 = ~x136 & ~n1420 ;
  assign n1422 = ~n1419 & n1421 ;
  assign n1423 = ~n1418 & ~n1422 ;
  assign n1424 = ~x137 & ~n1423 ;
  assign n1425 = ~n1414 & ~n1424 ;
  assign n1426 = ~x26 & n604 ;
  assign n1427 = n1272 & n1426 ;
  assign n1428 = ~n608 & ~n1427 ;
  assign n1429 = n202 & ~n1428 ;
  assign n1430 = x36 & n1248 ;
  assign n1431 = ~x97 & x138 ;
  assign n1432 = ~x81 & ~x138 ;
  assign n1433 = ~x136 & ~n1432 ;
  assign n1434 = ~n1431 & n1433 ;
  assign n1435 = ~n1430 & ~n1434 ;
  assign n1436 = x137 & ~n1435 ;
  assign n1437 = x71 & ~x138 ;
  assign n1438 = ~x98 & x138 ;
  assign n1439 = x136 & ~n1438 ;
  assign n1440 = ~n1437 & n1439 ;
  assign n1441 = x76 & ~x138 ;
  assign n1442 = ~x23 & x138 ;
  assign n1443 = ~x136 & ~n1442 ;
  assign n1444 = ~n1441 & n1443 ;
  assign n1445 = ~n1440 & ~n1444 ;
  assign n1446 = ~x137 & ~n1445 ;
  assign n1447 = ~n1436 & ~n1446 ;
  assign n1448 = x30 & n1248 ;
  assign n1449 = ~x111 & x138 ;
  assign n1450 = ~x86 & ~x138 ;
  assign n1451 = ~x136 & ~n1450 ;
  assign n1452 = ~n1449 & n1451 ;
  assign n1453 = ~n1448 & ~n1452 ;
  assign n1454 = x137 & ~n1453 ;
  assign n1455 = x64 & ~x138 ;
  assign n1456 = ~x88 & x138 ;
  assign n1457 = x136 & ~n1456 ;
  assign n1458 = ~n1455 & n1457 ;
  assign n1459 = x67 & ~x138 ;
  assign n1460 = ~x120 & x138 ;
  assign n1461 = ~x136 & ~n1460 ;
  assign n1462 = ~n1459 & n1461 ;
  assign n1463 = ~n1458 & ~n1462 ;
  assign n1464 = ~x137 & ~n1463 ;
  assign n1465 = ~n1454 & ~n1464 ;
  assign n1466 = ~x26 & n568 ;
  assign n1467 = ~n551 & ~n1466 ;
  assign n1468 = x116 & n202 ;
  assign n1469 = ~n1467 & n1468 ;
  assign n1470 = ~x53 & x58 ;
  assign n1471 = ~x97 & n1470 ;
  assign n1472 = ~n696 & ~n1471 ;
  assign n1473 = n1468 & ~n1472 ;
  assign n1474 = ~x139 & n1312 ;
  assign n1475 = ~x129 & n1157 ;
  assign n1476 = ~x111 & ~n1312 ;
  assign n1477 = n1475 & ~n1476 ;
  assign n1478 = ~n1474 & n1477 ;
  assign n1479 = x112 & ~n1312 ;
  assign n1480 = ~x141 & n1312 ;
  assign n1481 = n1475 & ~n1480 ;
  assign n1482 = ~n1479 & n1481 ;
  assign n1483 = ~x11 & ~x22 ;
  assign n1484 = x54 & n1483 ;
  assign n1485 = ~x54 & x113 ;
  assign n1486 = n202 & ~n1485 ;
  assign n1487 = ~n1484 & n1486 ;
  assign n1488 = x115 & ~n1312 ;
  assign n1489 = ~x140 & n1312 ;
  assign n1490 = n1475 & ~n1489 ;
  assign n1491 = ~n1488 & n1490 ;
  assign n1492 = x54 & n202 ;
  assign n1493 = ~x4 & ~x9 ;
  assign n1494 = n205 & n1493 ;
  assign n1495 = n1492 & ~n1494 ;
  assign n1496 = x122 & ~x129 ;
  assign n1497 = ~x54 & x118 ;
  assign n1498 = x54 & ~x59 ;
  assign n1499 = n382 & n1498 ;
  assign n1500 = ~n1497 & ~n1499 ;
  assign n1501 = ~x129 & ~n1500 ;
  assign n1502 = ~x129 & ~n569 ;
  assign n1503 = ~x120 & n1318 ;
  assign n1504 = ~x111 & ~x129 ;
  assign n1505 = ~n1503 & n1504 ;
  assign n1506 = x81 & x120 ;
  assign n1507 = ~x129 & n1506 ;
  assign n1508 = ~x129 & ~x134 ;
  assign n1509 = ~x129 & ~x135 ;
  assign n1510 = x57 & ~x129 ;
  assign n1511 = ~x96 & x125 ;
  assign n1512 = ~x3 & ~n1511 ;
  assign n1513 = ~x129 & ~n1512 ;
  assign n1514 = ~x126 & x132 ;
  assign n1515 = x133 & n1514 ;
  assign y0 = x108 ;
  assign y1 = x83 ;
  assign y2 = x104 ;
  assign y3 = x103 ;
  assign y4 = x102 ;
  assign y5 = x105 ;
  assign y6 = x107 ;
  assign y7 = x101 ;
  assign y8 = x126 ;
  assign y9 = x121 ;
  assign y10 = x1 ;
  assign y11 = x0 ;
  assign y12 = ~1'b0 ;
  assign y13 = x130 ;
  assign y14 = x128 ;
  assign y15 = ~n203 ;
  assign y16 = ~n239 ;
  assign y17 = n278 ;
  assign y18 = ~n293 ;
  assign y19 = n308 ;
  assign y20 = n321 ;
  assign y21 = n329 ;
  assign y22 = n336 ;
  assign y23 = n347 ;
  assign y24 = n354 ;
  assign y25 = n364 ;
  assign y26 = n373 ;
  assign y27 = n380 ;
  assign y28 = n391 ;
  assign y29 = n399 ;
  assign y30 = n431 ;
  assign y31 = n439 ;
  assign y32 = n448 ;
  assign y33 = n458 ;
  assign y34 = n467 ;
  assign y35 = n495 ;
  assign y36 = n503 ;
  assign y37 = n512 ;
  assign y38 = n515 ;
  assign y39 = n545 ;
  assign y40 = n597 ;
  assign y41 = n606 ;
  assign y42 = n618 ;
  assign y43 = n674 ;
  assign y44 = n714 ;
  assign y45 = n721 ;
  assign y46 = n728 ;
  assign y47 = n735 ;
  assign y48 = n742 ;
  assign y49 = n749 ;
  assign y50 = n756 ;
  assign y51 = n763 ;
  assign y52 = n770 ;
  assign y53 = n803 ;
  assign y54 = n810 ;
  assign y55 = n836 ;
  assign y56 = n857 ;
  assign y57 = n880 ;
  assign y58 = n901 ;
  assign y59 = n910 ;
  assign y60 = n936 ;
  assign y61 = n952 ;
  assign y62 = n971 ;
  assign y63 = n996 ;
  assign y64 = ~n1019 ;
  assign y65 = n1040 ;
  assign y66 = n1044 ;
  assign y67 = n1048 ;
  assign y68 = n1058 ;
  assign y69 = ~n1063 ;
  assign y70 = n1066 ;
  assign y71 = n1095 ;
  assign y72 = n1120 ;
  assign y73 = n1127 ;
  assign y74 = n1147 ;
  assign y75 = ~n1151 ;
  assign y76 = n1154 ;
  assign y77 = ~n1163 ;
  assign y78 = ~n1167 ;
  assign y79 = ~n1171 ;
  assign y80 = ~n1175 ;
  assign y81 = ~n1181 ;
  assign y82 = ~n1185 ;
  assign y83 = ~n1189 ;
  assign y84 = ~n1193 ;
  assign y85 = ~n1197 ;
  assign y86 = ~n1201 ;
  assign y87 = ~n1205 ;
  assign y88 = ~n1209 ;
  assign y89 = ~n1213 ;
  assign y90 = ~n1217 ;
  assign y91 = ~n1221 ;
  assign y92 = ~n1225 ;
  assign y93 = n1231 ;
  assign y94 = n1235 ;
  assign y95 = n1239 ;
  assign y96 = n1243 ;
  assign y97 = n1247 ;
  assign y98 = ~n1266 ;
  assign y99 = n1270 ;
  assign y100 = n1276 ;
  assign y101 = n1280 ;
  assign y102 = n1284 ;
  assign y103 = n1290 ;
  assign y104 = n1294 ;
  assign y105 = n1298 ;
  assign y106 = n1302 ;
  assign y107 = n1306 ;
  assign y108 = n1310 ;
  assign y109 = n1317 ;
  assign y110 = n1324 ;
  assign y111 = n1328 ;
  assign y112 = n1332 ;
  assign y113 = n1336 ;
  assign y114 = n1340 ;
  assign y115 = n1344 ;
  assign y116 = ~n1362 ;
  assign y117 = ~n1377 ;
  assign y118 = ~n1392 ;
  assign y119 = ~n1407 ;
  assign y120 = ~n1425 ;
  assign y121 = n1429 ;
  assign y122 = ~n1447 ;
  assign y123 = ~n1465 ;
  assign y124 = n1469 ;
  assign y125 = n1473 ;
  assign y126 = n1478 ;
  assign y127 = n1482 ;
  assign y128 = n1487 ;
  assign y129 = ~n1064 ;
  assign y130 = n1491 ;
  assign y131 = n1495 ;
  assign y132 = ~n1496 ;
  assign y133 = n1501 ;
  assign y134 = n1502 ;
  assign y135 = n1505 ;
  assign y136 = n1507 ;
  assign y137 = ~n1508 ;
  assign y138 = ~n1509 ;
  assign y139 = n1510 ;
  assign y140 = n1513 ;
  assign y141 = n1515 ;
endmodule
