module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 ;
  assign n33 = x29 & x30 ;
  assign n34 = x27 & x28 ;
  assign n35 = n33 & n34 ;
  assign n36 = x26 & x27 ;
  assign n37 = n35 & n36 ;
  assign n38 = x22 & x23 ;
  assign n39 = x23 & x24 ;
  assign n40 = n38 & n39 ;
  assign n41 = x25 & x26 ;
  assign n42 = x24 & x25 ;
  assign n43 = n41 & n42 ;
  assign n44 = n40 & n43 ;
  assign n45 = ~n37 & ~n44 ;
  assign n46 = n34 & n36 ;
  assign n47 = n43 & n46 ;
  assign n48 = ~n45 & n47 ;
  assign n49 = x28 & x29 ;
  assign n50 = x30 & x31 ;
  assign n51 = n33 & n50 ;
  assign n52 = n49 & n51 ;
  assign n53 = n34 & n52 ;
  assign n54 = n36 & n41 ;
  assign n55 = n39 & n42 ;
  assign n56 = n54 & n55 ;
  assign n57 = ~n53 & ~n56 ;
  assign n58 = n34 & n49 ;
  assign n59 = n54 & n58 ;
  assign n60 = ~n57 & n59 ;
  assign n61 = n48 & n60 ;
  assign n62 = x10 & x11 ;
  assign n63 = x17 & x18 ;
  assign n64 = ~n62 & ~n63 ;
  assign n65 = x12 & x13 ;
  assign n66 = x13 & x14 ;
  assign n67 = n65 & n66 ;
  assign n68 = x14 & x15 ;
  assign n69 = x15 & x16 ;
  assign n70 = n68 & n69 ;
  assign n71 = n67 & n70 ;
  assign n72 = n64 & n71 ;
  assign n73 = n72 ^ n71 ;
  assign n74 = x19 & x20 ;
  assign n75 = x18 & x19 ;
  assign n76 = n74 & n75 ;
  assign n77 = n63 & n75 ;
  assign n78 = x16 & x17 ;
  assign n79 = n69 & n78 ;
  assign n80 = n77 & n79 ;
  assign n81 = n76 & n80 ;
  assign n82 = ~n73 & ~n81 ;
  assign n83 = x11 & x12 ;
  assign n84 = ~n75 & ~n83 ;
  assign n85 = n66 & n68 ;
  assign n86 = n79 & n85 ;
  assign n87 = n84 & n86 ;
  assign n88 = n87 ^ n86 ;
  assign n89 = ~n82 & n88 ;
  assign n90 = x21 & x22 ;
  assign n91 = ~n68 & ~n90 ;
  assign n92 = n63 & n78 ;
  assign n93 = n76 & n92 ;
  assign n94 = n91 & n93 ;
  assign n95 = n94 ^ n93 ;
  assign n96 = x20 & x21 ;
  assign n97 = n75 & n96 ;
  assign n98 = n92 & n97 ;
  assign n99 = n80 & n98 ;
  assign n100 = n95 & n99 ;
  assign n101 = ~n89 & ~n100 ;
  assign n102 = ~n61 & n101 ;
  assign n103 = n74 & n90 ;
  assign n104 = n76 & n103 ;
  assign n105 = n38 & n96 ;
  assign n106 = n104 & n105 ;
  assign n107 = n63 & n97 ;
  assign n108 = n106 & n107 ;
  assign n109 = ~n39 & ~n78 ;
  assign n110 = n108 & ~n109 ;
  assign n111 = ~n41 & ~n75 ;
  assign n112 = n39 & n90 ;
  assign n113 = n96 & n112 ;
  assign n114 = ~n111 & n113 ;
  assign n115 = n46 & n56 ;
  assign n116 = ~n114 & ~n115 ;
  assign n117 = ~n36 & ~n74 ;
  assign n118 = n38 & n90 ;
  assign n119 = n55 & n118 ;
  assign n120 = ~n117 & n119 ;
  assign n121 = ~n116 & n120 ;
  assign n122 = ~n110 & ~n121 ;
  assign n123 = n102 & n122 ;
  assign n124 = x8 & x9 ;
  assign n125 = x7 & n124 ;
  assign n126 = x9 & x10 ;
  assign n127 = n83 & n126 ;
  assign n128 = n125 & n127 ;
  assign n129 = x7 & x8 ;
  assign n130 = n126 & n129 ;
  assign n131 = x6 & x7 ;
  assign n132 = n129 & n131 ;
  assign n133 = n130 & n132 ;
  assign n134 = n128 & n133 ;
  assign n135 = n62 & n126 ;
  assign n136 = n66 & n83 ;
  assign n137 = n135 & n136 ;
  assign n138 = n124 & n126 ;
  assign n139 = n62 & n83 ;
  assign n140 = n138 & n139 ;
  assign n141 = n137 & n140 ;
  assign n142 = n134 & n141 ;
  assign n143 = n142 ^ n134 ;
  assign n144 = n143 ^ n141 ;
  assign n145 = n65 & n83 ;
  assign n146 = n85 & n145 ;
  assign n147 = n70 & n146 ;
  assign n148 = ~n144 & ~n147 ;
  assign n149 = n135 & n145 ;
  assign n150 = ~n68 & ~n129 ;
  assign n151 = n149 & n150 ;
  assign n152 = n151 ^ n149 ;
  assign n153 = ~n148 & n152 ;
  assign n154 = x4 & x5 ;
  assign n155 = x3 & x4 ;
  assign n156 = n154 & n155 ;
  assign n157 = x5 & x6 ;
  assign n158 = n129 & n157 ;
  assign n159 = n156 & n158 ;
  assign n160 = n154 & n157 ;
  assign n161 = x2 & x3 ;
  assign n162 = n155 & n161 ;
  assign n163 = n160 & n162 ;
  assign n164 = n159 & n163 ;
  assign n165 = n124 & n131 ;
  assign n166 = n157 & n165 ;
  assign n167 = n130 & n166 ;
  assign n168 = n154 & n161 ;
  assign n169 = x1 & x2 ;
  assign n170 = n155 & n169 ;
  assign n171 = x0 & x1 ;
  assign n172 = n170 & n171 ;
  assign n173 = n168 & n172 ;
  assign n174 = ~n167 & ~n173 ;
  assign n175 = ~n164 & n174 ;
  assign n176 = n131 & n157 ;
  assign n177 = n156 & n176 ;
  assign n178 = n160 & n165 ;
  assign n179 = n177 & n178 ;
  assign n180 = n131 & n154 ;
  assign n181 = n162 & n180 ;
  assign n182 = n161 & n169 ;
  assign n183 = n156 & n182 ;
  assign n184 = n181 & n183 ;
  assign n185 = n179 & n184 ;
  assign n186 = n185 ^ n179 ;
  assign n187 = n186 ^ n184 ;
  assign n188 = ~n175 & n187 ;
  assign n189 = n132 & n160 ;
  assign n190 = n167 & n189 ;
  assign n191 = ~n134 & ~n190 ;
  assign n192 = n62 & n124 ;
  assign n193 = n133 & n192 ;
  assign n194 = n166 & n193 ;
  assign n195 = ~n191 & n194 ;
  assign n196 = ~n188 & ~n195 ;
  assign n197 = ~n153 & n196 ;
  assign n198 = n123 & n197 ;
  assign n455 = ~n69 & ~n161 ;
  assign n456 = ~n33 & ~n49 ;
  assign n457 = n455 & n456 ;
  assign n458 = ~n62 & ~n83 ;
  assign n459 = ~n65 & ~n66 ;
  assign n460 = n458 & n459 ;
  assign n461 = n457 & n460 ;
  assign n462 = ~n50 & ~n90 ;
  assign n463 = ~n42 & n462 ;
  assign n464 = ~n34 & ~n36 ;
  assign n465 = n111 & n464 ;
  assign n466 = n463 & n465 ;
  assign n467 = n461 & n466 ;
  assign n468 = ~n131 & ~n157 ;
  assign n469 = n109 & n468 ;
  assign n397 = ~n38 & ~n96 ;
  assign n399 = n63 & n74 ;
  assign n400 = n399 ^ n63 ;
  assign n401 = n400 ^ n74 ;
  assign n470 = n397 & ~n401 ;
  assign n471 = n469 & n470 ;
  assign n472 = ~n124 & ~n126 ;
  assign n473 = ~n169 & ~n171 ;
  assign n474 = n472 & n473 ;
  assign n475 = ~n154 & ~n155 ;
  assign n476 = n150 & n475 ;
  assign n477 = n474 & n476 ;
  assign n478 = n471 & n477 ;
  assign n479 = n467 & n478 ;
  assign n426 = ~x18 & ~x19 ;
  assign n427 = ~x21 & ~x22 ;
  assign n428 = n426 & n427 ;
  assign n429 = ~x14 & ~x15 ;
  assign n430 = ~x16 & ~x17 ;
  assign n431 = n429 & n430 ;
  assign n432 = n428 & n431 ;
  assign n433 = ~x28 & ~x29 ;
  assign n434 = ~x30 & ~x31 ;
  assign n435 = n433 & n434 ;
  assign n436 = ~x23 & ~x24 ;
  assign n437 = ~x25 & ~x27 ;
  assign n438 = n436 & n437 ;
  assign n439 = n435 & n438 ;
  assign n440 = n432 & n439 ;
  assign n441 = ~x1 & ~x2 ;
  assign n442 = ~x4 & ~x5 ;
  assign n443 = n441 & n442 ;
  assign n234 = ~x20 & ~x26 ;
  assign n382 = ~x0 & ~x3 ;
  assign n444 = n234 & n382 ;
  assign n445 = n443 & n444 ;
  assign n446 = ~x10 & ~x11 ;
  assign n447 = ~x12 & ~x13 ;
  assign n448 = n446 & n447 ;
  assign n449 = ~x6 & ~x7 ;
  assign n450 = ~x8 & ~x9 ;
  assign n451 = n449 & n450 ;
  assign n452 = n448 & n451 ;
  assign n453 = n445 & n452 ;
  assign n454 = n440 & n453 ;
  assign n480 = n479 ^ n454 ;
  assign n368 = n44 ^ n40 ;
  assign n369 = n368 ^ n43 ;
  assign n370 = n46 & n51 ;
  assign n371 = n370 ^ n46 ;
  assign n372 = n371 ^ n51 ;
  assign n373 = ~n369 & ~n372 ;
  assign n374 = n85 & n138 ;
  assign n375 = n374 ^ n85 ;
  assign n376 = n375 ^ n138 ;
  assign n243 = n33 & n49 ;
  assign n377 = n70 & n243 ;
  assign n378 = n377 ^ n243 ;
  assign n379 = n378 ^ n70 ;
  assign n380 = ~n376 & ~n379 ;
  assign n381 = n373 & n380 ;
  assign n383 = n169 & ~n382 ;
  assign n384 = n79 & n92 ;
  assign n385 = n384 ^ n79 ;
  assign n386 = n385 ^ n92 ;
  assign n387 = n383 & ~n386 ;
  assign n388 = n387 ^ n386 ;
  assign n389 = n56 ^ n54 ;
  assign n390 = n389 ^ n55 ;
  assign n240 = x19 & n96 ;
  assign n391 = n58 & n240 ;
  assign n392 = n391 ^ n58 ;
  assign n393 = n392 ^ n240 ;
  assign n394 = ~n390 & ~n393 ;
  assign n395 = ~n388 & n394 ;
  assign n396 = n381 & n395 ;
  assign n398 = n90 & ~n397 ;
  assign n402 = n75 & ~n401 ;
  assign n403 = n402 ^ n75 ;
  assign n404 = n177 ^ n176 ;
  assign n405 = n404 ^ n156 ;
  assign n406 = n403 & ~n405 ;
  assign n407 = n406 ^ n405 ;
  assign n408 = n398 & ~n407 ;
  assign n409 = n408 ^ n407 ;
  assign n410 = n135 & n139 ;
  assign n411 = n410 ^ n135 ;
  assign n412 = n411 ^ n139 ;
  assign n413 = n67 & n145 ;
  assign n414 = n413 ^ n67 ;
  assign n415 = n414 ^ n145 ;
  assign n416 = ~n412 & ~n415 ;
  assign n417 = n189 ^ n132 ;
  assign n418 = n417 ^ n160 ;
  assign n419 = n125 & n162 ;
  assign n420 = n419 ^ n125 ;
  assign n421 = n420 ^ n162 ;
  assign n422 = ~n418 & ~n421 ;
  assign n423 = n416 & n422 ;
  assign n424 = ~n409 & n423 ;
  assign n425 = n396 & n424 ;
  assign n481 = n480 ^ n425 ;
  assign n303 = n38 & n42 ;
  assign n304 = n161 & n171 ;
  assign n305 = n303 & n304 ;
  assign n306 = n305 ^ n303 ;
  assign n307 = n306 ^ n304 ;
  assign n308 = n62 & n65 ;
  assign n309 = n63 & n69 ;
  assign n310 = n308 & n309 ;
  assign n311 = n310 ^ n308 ;
  assign n312 = n311 ^ n309 ;
  assign n313 = ~n307 & ~n312 ;
  assign n314 = n155 & n157 ;
  assign n315 = n136 & n314 ;
  assign n316 = n315 ^ n314 ;
  assign n317 = n316 ^ n136 ;
  assign n318 = n34 & n41 ;
  assign n319 = n158 & n318 ;
  assign n320 = n319 ^ n158 ;
  assign n321 = n320 ^ n318 ;
  assign n322 = ~n317 & ~n321 ;
  assign n323 = n313 & n322 ;
  assign n324 = n63 & n76 ;
  assign n325 = n75 & n78 ;
  assign n326 = n180 & n325 ;
  assign n327 = n326 ^ n325 ;
  assign n328 = n327 ^ n180 ;
  assign n329 = n324 & ~n328 ;
  assign n330 = n329 ^ n328 ;
  assign n331 = n66 & n69 ;
  assign n332 = n127 & n331 ;
  assign n333 = n332 ^ n331 ;
  assign n334 = n333 ^ n127 ;
  assign n335 = n65 & n68 ;
  assign n336 = n39 & n41 ;
  assign n337 = n335 & n336 ;
  assign n338 = n337 ^ n335 ;
  assign n339 = n338 ^ n336 ;
  assign n340 = ~n334 & ~n339 ;
  assign n341 = ~n330 & n340 ;
  assign n342 = n323 & n341 ;
  assign n251 = n42 & n54 ;
  assign n252 = ~n52 & ~n251 ;
  assign n343 = n130 & n165 ;
  assign n344 = n343 ^ n130 ;
  assign n345 = n344 ^ n165 ;
  assign n346 = n168 & n170 ;
  assign n347 = n346 ^ n170 ;
  assign n348 = n347 ^ n168 ;
  assign n349 = ~n345 & ~n348 ;
  assign n350 = n252 & n349 ;
  assign n351 = n97 & n112 ;
  assign n352 = n351 ^ n97 ;
  assign n353 = n352 ^ n112 ;
  assign n250 = n36 & n49 ;
  assign n254 = n68 & n78 ;
  assign n354 = n250 & n254 ;
  assign n355 = n354 ^ n250 ;
  assign n356 = n355 ^ n254 ;
  assign n357 = ~n353 & ~n356 ;
  assign n358 = n35 & n192 ;
  assign n359 = n358 ^ n35 ;
  assign n360 = n359 ^ n192 ;
  assign n361 = n103 & n105 ;
  assign n362 = n361 ^ n103 ;
  assign n363 = n362 ^ n105 ;
  assign n364 = ~n360 & ~n363 ;
  assign n365 = n357 & n364 ;
  assign n366 = n350 & n365 ;
  assign n367 = n342 & n366 ;
  assign n482 = n481 ^ n367 ;
  assign n226 = n67 & n139 ;
  assign n266 = ~n119 & ~n226 ;
  assign n236 = n70 & n92 ;
  assign n241 = n118 & n240 ;
  assign n267 = ~n236 & ~n241 ;
  assign n268 = n266 & n267 ;
  assign n269 = ~n71 & ~n80 ;
  assign n270 = ~n86 & ~n93 ;
  assign n271 = n269 & n270 ;
  assign n272 = n268 & n271 ;
  assign n273 = n45 & n57 ;
  assign n274 = n272 & n273 ;
  assign n275 = ~n104 & ~n107 ;
  assign n276 = ~n113 & n275 ;
  assign n277 = n163 & n177 ;
  assign n278 = n277 ^ n177 ;
  assign n279 = n278 ^ n163 ;
  assign n280 = n166 & ~n279 ;
  assign n281 = n280 ^ n279 ;
  assign n282 = ~n133 & ~n172 ;
  assign n283 = ~n281 & n282 ;
  assign n284 = n140 & n146 ;
  assign n285 = n284 ^ n140 ;
  assign n286 = n285 ^ n146 ;
  assign n287 = n47 & n59 ;
  assign n288 = n287 ^ n47 ;
  assign n289 = n288 ^ n59 ;
  assign n290 = ~n286 & ~n289 ;
  assign n291 = n125 & n135 ;
  assign n292 = n183 & n291 ;
  assign n293 = n292 ^ n291 ;
  assign n294 = n293 ^ n183 ;
  assign n295 = n149 & n189 ;
  assign n296 = n295 ^ n149 ;
  assign n297 = n296 ^ n189 ;
  assign n298 = ~n294 & ~n297 ;
  assign n299 = n290 & n298 ;
  assign n300 = n283 & n299 ;
  assign n301 = n276 & n300 ;
  assign n302 = n274 & n301 ;
  assign n483 = n482 ^ n302 ;
  assign n206 = n160 & n183 ;
  assign n224 = ~n115 & ~n206 ;
  assign n225 = n44 & n54 ;
  assign n227 = n85 & n226 ;
  assign n228 = ~n225 & ~n227 ;
  assign n229 = n224 & n228 ;
  assign n230 = ~n137 & ~n147 ;
  assign n231 = ~n81 & ~n98 ;
  assign n232 = n230 & n231 ;
  assign n233 = n229 & n232 ;
  assign n235 = n119 & ~n234 ;
  assign n237 = ~x13 & ~x19 ;
  assign n238 = n236 & ~n237 ;
  assign n239 = ~n235 & ~n238 ;
  assign n242 = n40 & n241 ;
  assign n244 = n59 & n243 ;
  assign n245 = ~n242 & ~n244 ;
  assign n246 = n239 & n245 ;
  assign n247 = n174 & n246 ;
  assign n248 = n233 & n247 ;
  assign n249 = n103 & n107 ;
  assign n253 = n250 & ~n252 ;
  assign n255 = ~n140 & ~n254 ;
  assign n256 = n65 & ~n255 ;
  assign n257 = ~n253 & ~n256 ;
  assign n258 = ~n249 & n257 ;
  assign n259 = ~n159 & ~n178 ;
  assign n260 = ~n128 & ~n181 ;
  assign n261 = n259 & n260 ;
  assign n262 = ~n106 & ~n193 ;
  assign n263 = n261 & n262 ;
  assign n264 = n258 & n263 ;
  assign n265 = n248 & n264 ;
  assign n484 = n483 ^ n265 ;
  assign n199 = ~n48 & ~n60 ;
  assign n200 = ~n108 & n199 ;
  assign n201 = ~n187 & n190 ;
  assign n202 = n201 ^ n187 ;
  assign n203 = ~n144 & n194 ;
  assign n204 = n203 ^ n144 ;
  assign n205 = ~n202 & ~n204 ;
  assign n207 = n172 & n206 ;
  assign n208 = ~n99 & ~n114 ;
  assign n209 = ~n207 & n208 ;
  assign n210 = n88 & n95 ;
  assign n211 = n210 ^ n88 ;
  assign n212 = n211 ^ n95 ;
  assign n213 = n120 & ~n212 ;
  assign n214 = n213 ^ n212 ;
  assign n215 = n73 & n152 ;
  assign n216 = n215 ^ n73 ;
  assign n217 = n216 ^ n152 ;
  assign n218 = n164 & ~n217 ;
  assign n219 = n218 ^ n217 ;
  assign n220 = ~n214 & ~n219 ;
  assign n221 = n209 & n220 ;
  assign n222 = n205 & n221 ;
  assign n223 = n200 & n222 ;
  assign n485 = n484 ^ n223 ;
  assign n486 = ~n198 & ~n485 ;
  assign n497 = n454 & n479 ;
  assign n492 = n454 ^ n425 ;
  assign n493 = n492 ^ n479 ;
  assign n494 = n454 ^ n367 ;
  assign n495 = n494 ^ n479 ;
  assign n496 = n493 & n495 ;
  assign n498 = n497 ^ n496 ;
  assign n499 = n498 ^ n495 ;
  assign n500 = n499 ^ n493 ;
  assign n487 = n482 ^ n265 ;
  assign n488 = n483 & n487 ;
  assign n489 = n488 ^ n487 ;
  assign n490 = n489 ^ n483 ;
  assign n491 = n490 ^ n482 ;
  assign n501 = n500 ^ n491 ;
  assign n502 = n486 & ~n501 ;
  assign n503 = n223 & n484 ;
  assign n504 = n503 ^ n484 ;
  assign n505 = n501 & n504 ;
  assign n506 = n505 ^ n504 ;
  assign n511 = n301 ^ n274 ;
  assign n512 = n482 ^ n274 ;
  assign n513 = ~n482 & ~n512 ;
  assign n514 = n513 ^ n482 ;
  assign n515 = n514 ^ n301 ;
  assign n516 = n511 & ~n515 ;
  assign n517 = n516 ^ n513 ;
  assign n518 = n517 ^ n301 ;
  assign n519 = n500 & ~n518 ;
  assign n520 = n519 ^ n500 ;
  assign n507 = ~n454 & ~n479 ;
  assign n508 = n425 & n480 ;
  assign n509 = n508 ^ n480 ;
  assign n510 = ~n507 & ~n509 ;
  assign n522 = n520 ^ n510 ;
  assign n521 = n510 & n520 ;
  assign n523 = n522 ^ n521 ;
  assign n524 = n506 & n523 ;
  assign n525 = n524 ^ n523 ;
  assign n526 = n502 & ~n525 ;
  assign n527 = ~n265 & ~n483 ;
  assign n528 = n500 & n527 ;
  assign n529 = n528 ^ n502 ;
  assign n530 = n528 ^ n523 ;
  assign n531 = ~n528 & ~n530 ;
  assign n532 = n531 ^ n528 ;
  assign n533 = n532 ^ n506 ;
  assign n534 = n523 ^ n506 ;
  assign n535 = n533 & ~n534 ;
  assign n536 = n535 ^ n531 ;
  assign n537 = n536 ^ n506 ;
  assign n538 = n537 ^ n502 ;
  assign n539 = n529 & n538 ;
  assign n540 = n539 ^ n529 ;
  assign n541 = n540 ^ n538 ;
  assign n542 = n541 ^ n537 ;
  assign n543 = n542 ^ n525 ;
  assign n544 = ~n486 & ~n504 ;
  assign n545 = n544 ^ n501 ;
  assign n546 = n485 ^ n198 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = 1'b0 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = n526 ;
  assign y29 = ~n543 ;
  assign y30 = n545 ;
  assign y31 = n546 ;
endmodule
