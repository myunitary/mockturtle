module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 ;
  assign n8 = x3 & x4 ;
  assign n9 = ~x0 & ~x1 ;
  assign n10 = n8 & ~n9 ;
  assign n13 = ~x3 & ~x4 ;
  assign n14 = x1 & x2 ;
  assign n15 = n13 & n14 ;
  assign n11 = x2 & x3 ;
  assign n12 = x4 & n11 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = ~n10 & ~n16 ;
  assign n25 = x1 & n13 ;
  assign n26 = x2 & n25 ;
  assign n20 = ~x0 & x3 ;
  assign n21 = ~x1 & x4 ;
  assign n22 = n20 & n21 ;
  assign n18 = n8 ^ x4 ;
  assign n19 = x1 & n18 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = ~x2 & n23 ;
  assign n27 = n26 ^ n24 ;
  assign n34 = ~x2 & x4 ;
  assign n35 = n9 & n34 ;
  assign n31 = ~x0 & ~x2 ;
  assign n32 = n18 & n31 ;
  assign n28 = n8 ^ x3 ;
  assign n29 = x1 & ~x2 ;
  assign n30 = n28 & n29 ;
  assign n33 = n32 ^ n30 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = x0 & n8 ;
  assign n38 = n14 ^ x1 ;
  assign n39 = n38 ^ x2 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = x3 & ~n40 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = n37 & n43 ;
  assign n45 = n44 ^ n43 ;
  assign n54 = x0 & x2 ;
  assign n55 = n18 & n54 ;
  assign n48 = x5 & x6 ;
  assign n49 = n8 & n48 ;
  assign n50 = n49 ^ n28 ;
  assign n51 = x0 & n50 ;
  assign n46 = x4 & x5 ;
  assign n47 = n20 & n46 ;
  assign n52 = n51 ^ n47 ;
  assign n53 = n29 & n52 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = x4 & x6 ;
  assign n58 = n57 ^ x4 ;
  assign n59 = ~x2 & x3 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = n60 ^ x2 ;
  assign n62 = n14 & ~n18 ;
  assign n63 = n62 ^ x1 ;
  assign n64 = ~n61 & n63 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = x0 & x1 ;
  assign n67 = n8 & n66 ;
  assign n68 = n67 ^ n8 ;
  assign n69 = n68 ^ x2 ;
  assign n70 = x4 ^ x2 ;
  assign n71 = x4 ^ x3 ;
  assign n72 = n70 & n71 ;
  assign n73 = n72 ^ n71 ;
  assign n74 = n73 ^ x4 ;
  assign n75 = n74 ^ x2 ;
  assign n76 = ~n74 & n75 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = n77 ^ n68 ;
  assign n79 = ~n69 & ~n78 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = n80 ^ n68 ;
  assign n88 = x4 & n20 ;
  assign n89 = ~n39 & n88 ;
  assign n84 = x1 & ~x3 ;
  assign n85 = ~x4 & n84 ;
  assign n82 = x0 & x3 ;
  assign n83 = x4 & n82 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = x2 & n86 ;
  assign n90 = n89 ^ n87 ;
  assign n93 = x2 & ~x3 ;
  assign n92 = x2 & ~x4 ;
  assign n94 = n93 ^ n92 ;
  assign n97 = x1 & ~n94 ;
  assign n91 = ~x0 & n18 ;
  assign n95 = n29 & ~n94 ;
  assign n96 = ~n91 & n95 ;
  assign n98 = n97 ^ n96 ;
  assign n100 = n29 & n91 ;
  assign n99 = n8 & ~n39 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = n101 ^ n26 ;
  assign n109 = x2 & n18 ;
  assign n103 = ~x0 & x1 ;
  assign n104 = n18 & ~n103 ;
  assign n106 = ~n21 & n59 ;
  assign n107 = ~n104 & n106 ;
  assign n105 = ~x2 & n104 ;
  assign n108 = n107 ^ n105 ;
  assign n110 = n109 ^ n108 ;
  assign n111 = ~x0 & n13 ;
  assign n112 = ~n39 & n111 ;
  assign n115 = ~n9 & n18 ;
  assign n116 = n115 ^ x3 ;
  assign n117 = ~x2 & ~n116 ;
  assign n113 = ~x4 & ~n84 ;
  assign n114 = x2 & n113 ;
  assign n118 = n117 ^ n114 ;
  assign n119 = x2 & n13 ;
  assign n120 = x0 & n119 ;
  assign n121 = ~x0 & x2 ;
  assign n122 = n13 & n121 ;
  assign n123 = ~x1 & n28 ;
  assign n124 = n121 & n123 ;
  assign n125 = x0 & ~x1 ;
  assign n126 = n28 & n125 ;
  assign n127 = x2 & n126 ;
  assign n128 = x2 & n28 ;
  assign n129 = n66 & n128 ;
  assign n130 = n103 & n128 ;
  assign n131 = x2 & n68 ;
  assign n132 = n131 ^ x2 ;
  assign n136 = x2 & n66 ;
  assign n137 = n136 ^ n66 ;
  assign n138 = n46 ^ x4 ;
  assign n139 = x3 & n138 ;
  assign n140 = n139 ^ x3 ;
  assign n141 = n137 & n140 ;
  assign n133 = n128 ^ n28 ;
  assign n134 = n125 & n133 ;
  assign n135 = n134 ^ x2 ;
  assign n142 = n141 ^ n135 ;
  assign n143 = n132 & n142 ;
  assign n144 = n143 ^ n142 ;
  assign n149 = x1 & x5 ;
  assign n150 = ~x6 & n149 ;
  assign n146 = x0 & ~x2 ;
  assign n151 = n8 & n146 ;
  assign n152 = n150 & n151 ;
  assign n145 = ~x1 & x3 ;
  assign n147 = ~x4 & n146 ;
  assign n148 = n145 & n147 ;
  assign n153 = n152 ^ n148 ;
  assign n154 = n50 & n137 ;
  assign n155 = n154 ^ n131 ;
  assign n156 = x1 ^ x0 ;
  assign n157 = ~x2 & n18 ;
  assign n158 = ~n156 & n157 ;
  assign n159 = ~x1 & n18 ;
  assign n160 = n146 & n159 ;
  assign y0 = ~n17 ;
  assign y1 = n27 ;
  assign y2 = n36 ;
  assign y3 = n45 ;
  assign y4 = n56 ;
  assign y5 = n65 ;
  assign y6 = ~n81 ;
  assign y7 = n90 ;
  assign y8 = n98 ;
  assign y9 = n102 ;
  assign y10 = n110 ;
  assign y11 = n112 ;
  assign y12 = ~n118 ;
  assign y13 = n120 ;
  assign y14 = n122 ;
  assign y15 = n124 ;
  assign y16 = n127 ;
  assign y17 = n129 ;
  assign y18 = n130 ;
  assign y19 = n119 ;
  assign y20 = n144 ;
  assign y21 = n153 ;
  assign y22 = n155 ;
  assign y23 = ~1'b0 ;
  assign y24 = n158 ;
  assign y25 = n160 ;
endmodule
