module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 ;
  assign n33 = ~x0 & ~x1 ;
  assign n34 = x2 & x3 ;
  assign n35 = n34 ^ x2 ;
  assign n36 = n35 ^ x3 ;
  assign n37 = x4 & x5 ;
  assign n38 = n37 ^ x4 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = n36 & n39 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n33 & ~n42 ;
  assign n44 = x10 & x11 ;
  assign n45 = n44 ^ x10 ;
  assign n46 = n45 ^ x11 ;
  assign n47 = x13 & x14 ;
  assign n48 = n47 ^ x13 ;
  assign n49 = n48 ^ x14 ;
  assign n50 = n46 & n49 ;
  assign n51 = n50 ^ n46 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = x6 & x7 ;
  assign n54 = n53 ^ x6 ;
  assign n55 = n54 ^ x7 ;
  assign n56 = x8 & x9 ;
  assign n57 = n56 ^ x8 ;
  assign n58 = n57 ^ x9 ;
  assign n59 = n55 & n58 ;
  assign n60 = n59 ^ n55 ;
  assign n61 = n60 ^ n58 ;
  assign n62 = ~n52 & ~n61 ;
  assign n63 = n43 & n62 ;
  assign n64 = x21 & x22 ;
  assign n65 = n64 ^ x21 ;
  assign n66 = n65 ^ x22 ;
  assign n67 = x20 & x23 ;
  assign n68 = n67 ^ x20 ;
  assign n69 = n68 ^ x23 ;
  assign n70 = n66 & ~n69 ;
  assign n71 = n70 ^ n69 ;
  assign n72 = ~x24 & ~x25 ;
  assign n73 = ~n71 & n72 ;
  assign n74 = x16 & x17 ;
  assign n75 = n74 ^ x16 ;
  assign n76 = n75 ^ x17 ;
  assign n77 = x18 & n76 ;
  assign n78 = n77 ^ x18 ;
  assign n79 = n78 ^ n76 ;
  assign n80 = x12 & x15 ;
  assign n81 = n80 ^ x12 ;
  assign n82 = n81 ^ x15 ;
  assign n83 = x19 & ~n82 ;
  assign n84 = n83 ^ n82 ;
  assign n85 = n79 & ~n84 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = n86 ^ n73 ;
  assign n88 = n73 & ~n87 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = n89 ^ n86 ;
  assign n91 = n90 ^ n63 ;
  assign n92 = n63 & n91 ;
  assign n93 = n92 ^ n91 ;
  assign n94 = n93 ^ n89 ;
  assign n95 = n94 ^ n86 ;
  assign n96 = ~x28 & ~x29 ;
  assign n97 = ~x30 & ~x31 ;
  assign n98 = n96 & n97 ;
  assign n101 = ~x26 & ~x27 ;
  assign n102 = n98 & n101 ;
  assign n99 = x26 & ~x27 ;
  assign n100 = n98 & n99 ;
  assign n103 = n102 ^ n100 ;
  assign n104 = n95 & n103 ;
  assign n105 = n104 ^ n102 ;
  assign n106 = ~n79 & ~n82 ;
  assign n107 = n63 & n106 ;
  assign n108 = ~x19 & ~n71 ;
  assign n109 = x24 & ~x25 ;
  assign n110 = n109 ^ n72 ;
  assign n111 = n108 & n110 ;
  assign n112 = n107 & n111 ;
  assign n113 = n112 ^ n72 ;
  assign n114 = n105 & n113 ;
  assign n115 = n114 ^ n105 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = n116 ^ n105 ;
  assign n118 = n117 ^ n113 ;
  assign n119 = ~x16 & ~x17 ;
  assign n120 = x18 & ~n82 ;
  assign n121 = n119 & n120 ;
  assign n122 = n63 & n121 ;
  assign n123 = n122 ^ x18 ;
  assign n124 = n106 ^ n63 ;
  assign n125 = n108 ^ n106 ;
  assign n126 = ~n108 & ~n125 ;
  assign n127 = n126 ^ n108 ;
  assign n128 = n127 ^ n63 ;
  assign n129 = n124 & ~n128 ;
  assign n130 = n129 ^ n126 ;
  assign n131 = n130 ^ n63 ;
  assign n132 = n123 & ~n131 ;
  assign n133 = n132 ^ n131 ;
  assign n134 = ~n118 & ~n133 ;
  assign n135 = n134 ^ n133 ;
  assign n136 = n33 & ~n82 ;
  assign n137 = ~n42 & n136 ;
  assign n138 = n62 & n137 ;
  assign n139 = n138 ^ x16 ;
  assign n140 = ~x17 & ~n139 ;
  assign n141 = ~n135 & n140 ;
  assign n142 = n139 ^ n133 ;
  assign n143 = ~n139 & ~n142 ;
  assign n144 = n143 ^ n133 ;
  assign n145 = n144 ^ n118 ;
  assign n146 = ~n118 & ~n145 ;
  assign n147 = n146 ^ n143 ;
  assign n148 = n147 ^ n133 ;
  assign n149 = n148 ^ n135 ;
  assign n150 = x17 & n149 ;
  assign n151 = n95 & n102 ;
  assign n152 = n151 ^ n102 ;
  assign n153 = ~x24 & x25 ;
  assign n154 = ~n71 & n153 ;
  assign n155 = ~n86 & n154 ;
  assign n156 = n63 & n155 ;
  assign n157 = n156 ^ x25 ;
  assign n158 = n152 & ~n157 ;
  assign n159 = x19 & ~n107 ;
  assign n160 = n63 & ~n86 ;
  assign n161 = x24 & ~n71 ;
  assign n162 = n161 ^ n71 ;
  assign n163 = ~n160 & ~n162 ;
  assign n164 = ~n159 & n163 ;
  assign n165 = n158 & n164 ;
  assign n166 = x16 & n138 ;
  assign n167 = n166 ^ n138 ;
  assign n168 = x17 & ~n167 ;
  assign n169 = n119 & n138 ;
  assign n170 = ~x18 & ~n169 ;
  assign n171 = ~n168 & n170 ;
  assign n172 = n165 & n171 ;
  assign n173 = n150 & n172 ;
  assign n174 = n173 ^ n150 ;
  assign n175 = n174 ^ n149 ;
  assign n176 = n175 ^ n172 ;
  assign n177 = n172 ^ n135 ;
  assign n178 = ~n141 & ~n177 ;
  assign n179 = ~n135 & n165 ;
  assign n181 = n165 & ~n171 ;
  assign n180 = ~n135 & ~n165 ;
  assign n182 = n181 ^ n180 ;
  assign n183 = n179 & n182 ;
  assign n184 = n183 ^ n182 ;
  assign n185 = x23 & ~n66 ;
  assign n186 = n185 ^ n66 ;
  assign n188 = ~n86 & ~n186 ;
  assign n189 = n63 & n188 ;
  assign n187 = ~x20 & ~n186 ;
  assign n190 = n189 ^ n187 ;
  assign n192 = ~n123 & n190 ;
  assign n193 = ~n131 & n192 ;
  assign n194 = n118 & n193 ;
  assign n195 = ~n165 & n194 ;
  assign n196 = n195 ^ n165 ;
  assign n191 = n118 & n190 ;
  assign n197 = n196 ^ n191 ;
  assign n198 = n165 & ~n191 ;
  assign n199 = ~x20 & ~n86 ;
  assign n200 = n63 & n199 ;
  assign n201 = n200 ^ x21 ;
  assign n202 = ~x22 & ~x23 ;
  assign n203 = ~x24 & n202 ;
  assign n204 = ~n157 & n203 ;
  assign n205 = n152 & n204 ;
  assign n206 = ~n201 & n205 ;
  assign n207 = n198 & n206 ;
  assign n208 = n207 ^ n206 ;
  assign n209 = n208 ^ n191 ;
  assign n211 = ~n113 & ~n201 ;
  assign n212 = ~x24 & ~n157 ;
  assign n213 = n152 & n212 ;
  assign n214 = n211 & n213 ;
  assign n210 = ~x24 & ~n201 ;
  assign n215 = n214 ^ n210 ;
  assign n216 = ~n191 & ~n215 ;
  assign n217 = ~x20 & ~x21 ;
  assign n218 = ~n86 & n217 ;
  assign n219 = n63 & n218 ;
  assign n220 = ~x23 & n219 ;
  assign n221 = n220 ^ n202 ;
  assign n226 = ~x24 & n200 ;
  assign n227 = n221 & n226 ;
  assign n228 = ~n118 & n227 ;
  assign n223 = ~x21 & ~x24 ;
  assign n224 = n221 & n223 ;
  assign n225 = ~n118 & n224 ;
  assign n229 = n228 ^ n225 ;
  assign n222 = n118 & n221 ;
  assign n230 = n229 ^ n222 ;
  assign n231 = n216 & n230 ;
  assign n232 = ~x22 & n219 ;
  assign n233 = x23 & ~n232 ;
  assign n234 = n107 & n108 ;
  assign n235 = ~x24 & ~n234 ;
  assign n236 = n158 & n235 ;
  assign n237 = ~n233 & n236 ;
  assign n238 = ~n221 & n237 ;
  assign n239 = n118 & ~n237 ;
  assign n240 = ~n113 & n158 ;
  assign n241 = n105 & ~n113 ;
  assign n242 = ~n158 & n241 ;
  assign n243 = x26 & n95 ;
  assign n244 = n243 ^ n95 ;
  assign n245 = ~n99 & ~n244 ;
  assign n246 = ~x27 & n95 ;
  assign n247 = n98 & ~n246 ;
  assign n248 = ~n245 & n247 ;
  assign n249 = x27 & ~x28 ;
  assign n250 = ~n244 & n249 ;
  assign n251 = n95 & n101 ;
  assign n252 = x28 & n251 ;
  assign n253 = ~n250 & ~n252 ;
  assign n254 = ~x29 & n97 ;
  assign n255 = ~n253 & n254 ;
  assign n256 = x29 & ~n251 ;
  assign n257 = ~n96 & n97 ;
  assign n258 = ~n252 & n257 ;
  assign n259 = ~n256 & n258 ;
  assign n260 = n252 ^ n251 ;
  assign n262 = x30 & ~x31 ;
  assign n261 = x29 & n97 ;
  assign n263 = n262 ^ n261 ;
  assign n265 = n263 ^ n262 ;
  assign n264 = n263 ^ x29 ;
  assign n266 = n265 ^ n264 ;
  assign n267 = n265 ^ n263 ;
  assign n268 = n266 & n267 ;
  assign n269 = n268 ^ n265 ;
  assign n270 = n260 & n269 ;
  assign n271 = n270 ^ n263 ;
  assign n272 = n271 ^ n262 ;
  assign n273 = n96 & n101 ;
  assign n274 = n95 & n273 ;
  assign n275 = n274 ^ x31 ;
  assign n276 = n274 ^ x30 ;
  assign n277 = n275 & n276 ;
  assign n278 = n277 ^ n276 ;
  assign y0 = n141 ;
  assign y1 = n176 ;
  assign y2 = n178 ;
  assign y3 = n184 ;
  assign y4 = n197 ;
  assign y5 = n209 ;
  assign y6 = n231 ;
  assign y7 = n238 ;
  assign y8 = n239 ;
  assign y9 = n240 ;
  assign y10 = n242 ;
  assign y11 = n248 ;
  assign y12 = n255 ;
  assign y13 = n259 ;
  assign y14 = n272 ;
  assign y15 = n278 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
  assign y30 = 1'b0 ;
  assign y31 = 1'b0 ;
endmodule
