module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 ;
  assign n8 = x3 & x4 ;
  assign n9 = ~x0 & ~x1 ;
  assign n10 = n8 & ~n9 ;
  assign n13 = ~x3 & ~x4 ;
  assign n14 = x1 & x2 ;
  assign n15 = n13 & n14 ;
  assign n11 = x2 & x3 ;
  assign n12 = x4 & n11 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = ~n10 & ~n16 ;
  assign n25 = x1 & n13 ;
  assign n26 = x2 & n25 ;
  assign n20 = ~x0 & x3 ;
  assign n21 = ~x1 & x4 ;
  assign n22 = n20 & n21 ;
  assign n18 = ~x3 & x4 ;
  assign n19 = x1 & n18 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = ~x2 & n23 ;
  assign n27 = n26 ^ n24 ;
  assign n34 = ~x2 & x4 ;
  assign n35 = n9 & n34 ;
  assign n31 = ~x0 & ~x2 ;
  assign n32 = n18 & n31 ;
  assign n28 = x3 & ~x4 ;
  assign n29 = x1 & ~x2 ;
  assign n30 = n28 & n29 ;
  assign n33 = n32 ^ n30 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = x0 & n8 ;
  assign n38 = ~x1 & ~x2 ;
  assign n39 = x3 & n38 ;
  assign n40 = n39 ^ n18 ;
  assign n41 = ~n37 & n40 ;
  assign n51 = x0 & x2 ;
  assign n52 = n18 & n51 ;
  assign n47 = x4 & x5 ;
  assign n48 = n20 & n47 ;
  assign n49 = n29 & n48 ;
  assign n42 = x5 & x6 ;
  assign n43 = n8 & n42 ;
  assign n44 = n43 ^ n28 ;
  assign n45 = x0 & n29 ;
  assign n46 = n44 & n45 ;
  assign n50 = n49 ^ n46 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = x4 & ~x6 ;
  assign n55 = ~x2 & x3 ;
  assign n56 = ~n54 & n55 ;
  assign n57 = n56 ^ x2 ;
  assign n58 = n14 & ~n18 ;
  assign n59 = n58 ^ x1 ;
  assign n60 = n57 & n59 ;
  assign n61 = x0 & x1 ;
  assign n62 = n8 & ~n61 ;
  assign n63 = n34 ^ n11 ;
  assign n64 = n63 ^ n28 ;
  assign n65 = ~x2 & n64 ;
  assign n66 = n62 & n65 ;
  assign n67 = n66 ^ n64 ;
  assign n74 = x4 & n20 ;
  assign n75 = n38 & n74 ;
  assign n70 = x0 & x3 ;
  assign n71 = x4 & n70 ;
  assign n68 = x1 & ~x3 ;
  assign n69 = ~x4 & n68 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = x2 & n72 ;
  assign n76 = n75 ^ n73 ;
  assign n79 = x2 & ~x3 ;
  assign n78 = x2 & ~x4 ;
  assign n80 = n79 ^ n78 ;
  assign n83 = x1 & ~n80 ;
  assign n77 = ~x0 & n18 ;
  assign n81 = n29 & ~n80 ;
  assign n82 = ~n77 & n81 ;
  assign n84 = n83 ^ n82 ;
  assign n86 = n29 & n77 ;
  assign n85 = n8 & n38 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = n87 ^ n26 ;
  assign n95 = x2 & n18 ;
  assign n89 = ~x0 & x1 ;
  assign n90 = n18 & ~n89 ;
  assign n92 = ~n21 & n55 ;
  assign n93 = ~n90 & n92 ;
  assign n91 = ~x2 & n90 ;
  assign n94 = n93 ^ n91 ;
  assign n96 = n95 ^ n94 ;
  assign n97 = ~x0 & n13 ;
  assign n98 = n38 & n97 ;
  assign n101 = ~n9 & n18 ;
  assign n102 = n101 ^ x3 ;
  assign n103 = ~x2 & ~n102 ;
  assign n99 = ~x4 & ~n68 ;
  assign n100 = x2 & n99 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = x2 & n13 ;
  assign n106 = x0 & n105 ;
  assign n107 = ~x0 & x2 ;
  assign n108 = n13 & n107 ;
  assign n109 = ~x1 & n28 ;
  assign n110 = n107 & n109 ;
  assign n111 = x0 & ~x1 ;
  assign n112 = n28 & n111 ;
  assign n113 = x2 & n112 ;
  assign n114 = x2 & n28 ;
  assign n115 = n61 & n114 ;
  assign n116 = n89 & n114 ;
  assign n117 = x2 & ~n62 ;
  assign n121 = ~x2 & n61 ;
  assign n122 = x4 & ~x5 ;
  assign n123 = x3 & ~n122 ;
  assign n124 = n121 & n123 ;
  assign n118 = ~x2 & n28 ;
  assign n119 = n111 & n118 ;
  assign n120 = n119 ^ x2 ;
  assign n125 = n124 ^ n120 ;
  assign n126 = ~n117 & n125 ;
  assign n131 = x1 & x5 ;
  assign n132 = ~x6 & n131 ;
  assign n128 = x0 & ~x2 ;
  assign n133 = n8 & n128 ;
  assign n134 = n132 & n133 ;
  assign n127 = ~x1 & x3 ;
  assign n129 = ~x4 & n128 ;
  assign n130 = n127 & n129 ;
  assign n135 = n134 ^ n130 ;
  assign n137 = n44 & n121 ;
  assign n136 = x2 & n62 ;
  assign n138 = n137 ^ n136 ;
  assign n139 = ~x2 & n18 ;
  assign n140 = x1 ^ x0 ;
  assign n141 = n139 & ~n140 ;
  assign n142 = ~x1 & n18 ;
  assign n143 = n128 & n142 ;
  assign y0 = ~n17 ;
  assign y1 = n27 ;
  assign y2 = n36 ;
  assign y3 = n41 ;
  assign y4 = n53 ;
  assign y5 = n60 ;
  assign y6 = n67 ;
  assign y7 = n76 ;
  assign y8 = n84 ;
  assign y9 = n88 ;
  assign y10 = n96 ;
  assign y11 = n98 ;
  assign y12 = ~n104 ;
  assign y13 = n106 ;
  assign y14 = n108 ;
  assign y15 = n110 ;
  assign y16 = n113 ;
  assign y17 = n115 ;
  assign y18 = n116 ;
  assign y19 = n105 ;
  assign y20 = n126 ;
  assign y21 = n135 ;
  assign y22 = n138 ;
  assign y23 = ~1'b0 ;
  assign y24 = n141 ;
  assign y25 = n143 ;
endmodule
