// Benchmark "bitonic_sort_inc" written by ABC on Wed Jul  9 20:39:45 2025

module bitonic_sort_inc_2 ( 
    \in_array[0] , \in_array[1] , \in_array[2] , \in_array[3] ,
    \in_array[4] , \in_array[5] , \in_array[6] , \in_array[7] ,
    \in_array[8] , \in_array[9] , \in_array[10] , \in_array[11] ,
    \in_array[12] , \in_array[13] , \in_array[14] , \in_array[15] ,
    \out_array[0] , \out_array[1] , \out_array[2] , \out_array[3] ,
    \out_array[4] , \out_array[5] , \out_array[6] , \out_array[7] ,
    \out_array[8] , \out_array[9] , \out_array[10] , \out_array[11] ,
    \out_array[12] , \out_array[13] , \out_array[14] , \out_array[15]   );
  input  \in_array[0] , \in_array[1] , \in_array[2] , \in_array[3] ,
    \in_array[4] , \in_array[5] , \in_array[6] , \in_array[7] ,
    \in_array[8] , \in_array[9] , \in_array[10] , \in_array[11] ,
    \in_array[12] , \in_array[13] , \in_array[14] , \in_array[15] ;
  output \out_array[0] , \out_array[1] , \out_array[2] , \out_array[3] ,
    \out_array[4] , \out_array[5] , \out_array[6] , \out_array[7] ,
    \out_array[8] , \out_array[9] , \out_array[10] , \out_array[11] ,
    \out_array[12] , \out_array[13] , \out_array[14] , \out_array[15] ;
  wire new__347_, new__348_, new__349_, new__350_, new__351_, new__352_,
    new__353__neg, new__353_, new__354_, new__355_, new__356__neg,
    new__356_, new__357_, new__358_, new__359_, new__360__neg, new__360_,
    new__361_, new__362_, new__363_, new__364_, new__365_, new__366_,
    new__367_, new__000_, new__001_, new__002_, new__003_, new__004_,
    new__005_, new__006_, new__007_, new__008_, new__009_, new__010_,
    new__011_, new__012_, new__013_, new__014_, new__015_, new__016_,
    new__017_, new__018_, new__019_, new__020_, new__021_, new__022_,
    new__023__neg, new__023_, new__024_, new__025_, new__026_, new__027_,
    new__028_, new__029_, new__030_, new__031_, new__032_, new__033_,
    new__034_, new__035_, new__036_, new__037_, new__038_, new__039_,
    new__040__neg, new__040_, new__041_, new__042_, new__043_, new__044_,
    new__045_, new__046_, new__047_, new__048_, new__049_, new__050_,
    new__051_, new__052__neg, new__052_, new__053_, new__054__neg,
    new__054_, new__055_, new__056_, new__057_, new__058__neg, new__058_,
    new__059_, new__060_, new__061_, new__062_, new__063_, new__064_,
    new__065_, new__066__neg, new__066_, new__067_, new__068_, new__069_,
    new__070_, new__071_, new__072_, new__073_, new__074_, new__075_,
    new__076_, new__077_, new__078_, new__079__neg, new__079_, new__080_,
    new__081_, new__082_, new__083_, new__084_, new__085_, new__086_,
    new__087_, new__088__neg, new__088_, new__089_, new__090_, new__091_,
    new__092_, new__093_, new__094_, new__095_, new__096_, new__097_,
    new__098_, new__099_, new__100_, new__101_, new__102_, new__103_,
    new__104__neg, new__104_, new__105_, new__106_, new__107_, new__108_,
    new__109_, new__110_, new__111_, new__112_, new__113_, new__114_,
    new__115__neg, new__115_, new__116_, new__117_, new__118_, new__119_,
    new__120_, new__121_, new__122_, new__123_, new__124_, new__125_,
    new__126__neg, new__126_, new__127_, new__128_, new__129_, new__130_,
    new__131_, new__132__neg, new__132_, new__133_, new__134_,
    new__135__neg, new__135_, new__136_, new__137_, new__138_, new__139_,
    new__140__neg, new__140_, new__141_, new__142_, new__143_, new__144_,
    new__145_, new__146_, new__147_, new__148_, new__149_, new__150_,
    new__151_, new__152__neg, new__152_, new__153_, new__154_, new__155_,
    new__156_, new__157_, new__158_, new__159_, new__160_, new__161_,
    new__162_, new__163_, new__164_, new__165_, new__166_, new__167_,
    new__168__neg, new__168_, new__169_, new__170_, new__171_, new__172_,
    new__173_, new__174_, new__175_, new__176_, new__177_, new__178_,
    new__179_, new__180__neg, new__180_, new__181_, new__182_,
    new__183__neg, new__183_, new__184_, new__185_, new__186_, new__187_,
    new__188__neg, new__188_, new__189_, new__190_, new__191_, new__192_,
    new__193_, new__194_, new__195_, new__196__neg, new__196_, new__197_,
    new__198_, new__199_, new__200__neg, new__200_, new__201_, new__202_,
    new__203_, new__204__neg, new__204_, new__205_, new__206_, new__207_,
    new__208_, new__209_, new__210_, new__211_, new__212__neg, new__212_,
    new__213_, new__214_, new__215_, new__216_, new__217__neg, new__217_,
    new__218_, new__219_, new__220_, new__221_, new__222_, new__223_,
    new__224_, new__225_, new__226_, new__228_, new__229_, new__230__neg,
    new__230_, new__231_, new__232_, new__233_, new__235_, new__236_,
    new__237_, new__238__neg, new__238_, new__239_, new__240_, new__241_,
    new__242_, new__243_, new__245_, new__246_, new__247_, new__248_,
    new__249_, new__250_, new__251_, new__252_, new__253_, new__254_,
    new__256__neg, new__256_, new__257_, new__258_, new__259_, new__260_,
    new__261_, new__262_, new__263_, new__264_, new__265_, new__267_,
    new__268_, new__269__neg, new__269_, new__270_, new__271_, new__272_,
    new__273__neg, new__273_, new__274_, new__275_, new__276_,
    new__278__neg, new__278_, new__279_, new__280_, new__281_, new__282_,
    new__283_, new__284_, new__285_, new__287__neg, new__287_, new__288_,
    new__289_, new__290_, new__291_, new__292__neg, new__292_, new__293_,
    new__294_, new__295_, new__297_, new__298_, new__299_, new__300_,
    new__301_, new__302_, new__303_, new__304_, new__306__neg, new__306_,
    new__307_, new__308_, new__309_, new__227_, new__234_, new__244_,
    new__255_, new__266_, new__277_, new__286_, new__296_, new__305_,
    new__310_, new__311_, new__312_, new__313_, new__314_, new__315_,
    new__316_, new__317_, new__318_, new__319_, new__320_, new__321_,
    new__322_, new__323__neg, new__323_, new__324_, new__325_, new__326_,
    new__327_, new__328_, new__329_, new__330_, new__331_, new__332_,
    new__333_, new__334_, new__335_, new__336_, new__337_, new__338_,
    new__339_, new__340__neg, new__340_, new__341_, new__342_, new__343_,
    new__344_, new__345_, new__346_;
  assign new__347_ = ~new__346_;
  assign new__348_ = ~new__347_ ^ ~new__341_;
  assign new__349_ = new__348_ & new__345_;
  assign new__350_ = ~new__349_ ^ ~new__342_;
  assign new__351_ = new__350_ & new__340_;
  assign new__352_ = ~new__351_ ^ ~new__338_;
  assign new__353__neg = ~new__352_ ^ ~new__336_;
  assign new__353_ = ~new__353__neg;
  assign new__354_ = new__352_ & new__336_;
  assign new__355_ = ~new__354_;
  assign new__356__neg = ~new__331_ ^ ~new__328_;
  assign new__356_ = ~new__356__neg;
  assign new__357_ = new__356_ & new__334_;
  assign new__358_ = ~new__357_ ^ ~new__328_;
  assign new__359_ = ~new__358_ ^ ~new__354_;
  assign new__360__neg = ~new__346_ ^ ~new__343_;
  assign new__360_ = ~new__360__neg;
  assign new__361_ = new__360_ & new__350_;
  assign new__362_ = ~new__361_ ^ ~new__343_;
  assign new__363_ = ~new__362_ ^ ~new__354_;
  assign new__364_ = new__363_ & new__359_;
  assign new__365_ = ~new__364_ ^ ~new__355_;
  assign new__366_ = new__365_ & new__353_;
  assign new__367_ = ~new__366_ ^ ~new__336_;
  assign new__000_ = ~new__367_;
  assign new__001_ = ~\in_array[10] ;
  assign new__002_ = ~\in_array[10]  ^ ~\in_array[8] ;
  assign new__003_ = ~\in_array[8] ;
  assign new__004_ = \in_array[10]  & new__003_;
  assign new__005_ = ~new__004_;
  assign new__006_ = ~\in_array[9] ;
  assign new__007_ = ~new__004_ ^ ~new__006_;
  assign new__008_ = ~new__004_ ^ ~\in_array[11] ;
  assign new__009_ = new__008_ & new__007_;
  assign new__010_ = ~new__009_ ^ ~new__005_;
  assign new__011_ = new__010_ & new__002_;
  assign new__012_ = ~new__011_ ^ ~new__001_;
  assign new__013_ = ~\in_array[14]  ^ ~\in_array[12] ;
  assign new__014_ = ~\in_array[12] ;
  assign new__015_ = \in_array[14]  & new__014_;
  assign new__016_ = ~\in_array[13] ;
  assign new__017_ = ~new__015_ ^ ~new__016_;
  assign new__018_ = ~new__015_ ^ ~\in_array[15] ;
  assign new__019_ = new__018_ & new__017_;
  assign new__020_ = ~new__019_ ^ ~new__015_;
  assign new__021_ = new__020_ & new__013_;
  assign new__022_ = ~new__021_ ^ ~\in_array[14] ;
  assign new__023__neg = ~new__022_ ^ ~new__012_;
  assign new__023_ = ~new__023__neg;
  assign new__024_ = new__022_ & new__012_;
  assign new__025_ = ~\in_array[11] ;
  assign new__026_ = \in_array[9]  & new__025_;
  assign new__027_ = ~new__026_ ^ ~new__025_;
  assign new__028_ = ~new__027_ ^ ~new__024_;
  assign new__029_ = new__016_ & \in_array[15] ;
  assign new__030_ = ~new__029_ ^ ~\in_array[15] ;
  assign new__031_ = ~new__030_ ^ ~new__024_;
  assign new__032_ = new__031_ & new__028_;
  assign new__033_ = ~new__032_ ^ ~new__024_;
  assign new__034_ = new__033_ & new__023_;
  assign new__035_ = ~new__034_ ^ ~new__012_;
  assign new__036_ = ~new__035_;
  assign new__037_ = ~new__011_ ^ ~new__003_;
  assign new__038_ = ~new__037_;
  assign new__039_ = ~new__021_ ^ ~\in_array[12] ;
  assign new__040__neg = ~new__039_ ^ ~new__037_;
  assign new__040_ = ~new__040__neg;
  assign new__041_ = new__039_ & new__037_;
  assign new__042_ = ~new__026_ ^ ~\in_array[9] ;
  assign new__043_ = ~new__042_;
  assign new__044_ = ~new__043_ ^ ~new__041_;
  assign new__045_ = ~new__029_ ^ ~new__016_;
  assign new__046_ = ~new__045_;
  assign new__047_ = ~new__046_ ^ ~new__041_;
  assign new__048_ = new__047_ & new__044_;
  assign new__049_ = ~new__048_ ^ ~new__041_;
  assign new__050_ = new__049_ & new__040_;
  assign new__051_ = ~new__050_ ^ ~new__038_;
  assign new__052__neg = ~new__051_ ^ ~new__035_;
  assign new__052_ = ~new__052__neg;
  assign new__053_ = new__051_ & new__035_;
  assign new__054__neg = ~new__030_ ^ ~new__027_;
  assign new__054_ = ~new__054__neg;
  assign new__055_ = new__054_ & new__033_;
  assign new__056_ = ~new__055_ ^ ~new__027_;
  assign new__057_ = ~new__056_ ^ ~new__053_;
  assign new__058__neg = ~new__045_ ^ ~new__042_;
  assign new__058_ = ~new__058__neg;
  assign new__059_ = new__058_ & new__049_;
  assign new__060_ = ~new__059_ ^ ~new__042_;
  assign new__061_ = ~new__060_ ^ ~new__053_;
  assign new__062_ = new__061_ & new__057_;
  assign new__063_ = ~new__062_ ^ ~new__053_;
  assign new__064_ = new__063_ & new__052_;
  assign new__065_ = ~new__064_ ^ ~new__036_;
  assign new__066__neg = ~new__065_ ^ ~new__367_;
  assign new__066_ = ~new__066__neg;
  assign new__067_ = new__065_ & new__367_;
  assign new__068_ = ~new__067_;
  assign new__069_ = ~new__328_;
  assign new__070_ = ~new__357_ ^ ~new__069_;
  assign new__071_ = ~new__362_ ^ ~new__070_;
  assign new__072_ = new__071_ & new__365_;
  assign new__073_ = ~new__072_ ^ ~new__358_;
  assign new__074_ = ~new__073_ ^ ~new__067_;
  assign new__075_ = ~new__027_;
  assign new__076_ = ~new__055_ ^ ~new__075_;
  assign new__077_ = ~new__060_ ^ ~new__076_;
  assign new__078_ = new__077_ & new__063_;
  assign new__079__neg = ~new__078_ ^ ~new__056_;
  assign new__079_ = ~new__079__neg;
  assign new__080_ = ~new__079_ ^ ~new__067_;
  assign new__081_ = new__080_ & new__074_;
  assign new__082_ = ~new__081_ ^ ~new__068_;
  assign new__083_ = new__082_ & new__066_;
  assign new__084_ = ~new__083_ ^ ~new__000_;
  assign new__085_ = ~new__322_;
  assign new__086_ = ~new__335_ ^ ~new__085_;
  assign new__087_ = ~new__351_ ^ ~new__339_;
  assign new__088__neg = ~new__087_ ^ ~new__086_;
  assign new__088_ = ~new__088__neg;
  assign new__089_ = new__087_ & new__086_;
  assign new__090_ = ~new__089_;
  assign new__091_ = ~new__331_;
  assign new__092_ = ~new__357_ ^ ~new__091_;
  assign new__093_ = ~new__092_ ^ ~new__089_;
  assign new__094_ = ~new__361_ ^ ~new__347_;
  assign new__095_ = ~new__094_ ^ ~new__089_;
  assign new__096_ = new__095_ & new__093_;
  assign new__097_ = ~new__096_ ^ ~new__090_;
  assign new__098_ = new__097_ & new__088_;
  assign new__099_ = ~new__098_ ^ ~new__086_;
  assign new__100_ = ~new__022_;
  assign new__101_ = ~new__034_ ^ ~new__100_;
  assign new__102_ = ~new__101_;
  assign new__103_ = ~new__050_ ^ ~new__039_;
  assign new__104__neg = ~new__103_ ^ ~new__101_;
  assign new__104_ = ~new__104__neg;
  assign new__105_ = new__103_ & new__101_;
  assign new__106_ = ~new__030_;
  assign new__107_ = ~new__055_ ^ ~new__106_;
  assign new__108_ = ~new__107_ ^ ~new__105_;
  assign new__109_ = ~new__059_ ^ ~new__046_;
  assign new__110_ = ~new__109_ ^ ~new__105_;
  assign new__111_ = new__110_ & new__108_;
  assign new__112_ = ~new__111_ ^ ~new__105_;
  assign new__113_ = new__112_ & new__104_;
  assign new__114_ = ~new__113_ ^ ~new__102_;
  assign new__115__neg = ~new__114_ ^ ~new__099_;
  assign new__115_ = ~new__115__neg;
  assign new__116_ = new__114_ & new__099_;
  assign new__117_ = ~new__116_;
  assign new__118_ = ~new__357_ ^ ~new__331_;
  assign new__119_ = ~new__094_ ^ ~new__118_;
  assign new__120_ = new__119_ & new__097_;
  assign new__121_ = ~new__120_ ^ ~new__092_;
  assign new__122_ = ~new__121_ ^ ~new__116_;
  assign new__123_ = ~new__055_ ^ ~new__030_;
  assign new__124_ = ~new__109_ ^ ~new__123_;
  assign new__125_ = new__124_ & new__112_;
  assign new__126__neg = ~new__125_ ^ ~new__107_;
  assign new__126_ = ~new__126__neg;
  assign new__127_ = ~new__126_ ^ ~new__116_;
  assign new__128_ = new__127_ & new__122_;
  assign new__129_ = ~new__128_ ^ ~new__117_;
  assign new__130_ = new__129_ & new__115_;
  assign new__131_ = ~new__130_ ^ ~new__099_;
  assign new__132__neg = ~new__131_ ^ ~new__084_;
  assign new__132_ = ~new__132__neg;
  assign new__133_ = new__131_ & new__084_;
  assign new__134_ = ~new__133_;
  assign new__135__neg = ~new__126_ ^ ~new__121_;
  assign new__135_ = ~new__135__neg;
  assign new__136_ = new__135_ & new__129_;
  assign new__137_ = ~new__136_ ^ ~new__121_;
  assign new__138_ = ~new__137_ ^ ~new__133_;
  assign new__139_ = ~new__073_;
  assign new__140__neg = ~new__079_ ^ ~new__073_;
  assign new__140_ = ~new__140__neg;
  assign new__141_ = new__140_ & new__082_;
  assign new__142_ = ~new__141_ ^ ~new__139_;
  assign new__143_ = ~new__142_ ^ ~new__133_;
  assign new__144_ = new__143_ & new__138_;
  assign new__145_ = ~new__144_ ^ ~new__134_;
  assign new__146_ = new__145_ & new__132_;
  assign new__147_ = ~new__146_ ^ ~new__084_;
  assign new__148_ = ~new__352_;
  assign new__149_ = ~new__366_ ^ ~new__148_;
  assign new__150_ = ~new__149_;
  assign new__151_ = ~new__064_ ^ ~new__051_;
  assign new__152__neg = ~new__151_ ^ ~new__149_;
  assign new__152_ = ~new__152__neg;
  assign new__153_ = new__151_ & new__149_;
  assign new__154_ = ~new__153_;
  assign new__155_ = ~new__362_;
  assign new__156_ = ~new__072_ ^ ~new__155_;
  assign new__157_ = ~new__156_ ^ ~new__153_;
  assign new__158_ = ~new__078_ ^ ~new__060_;
  assign new__159_ = ~new__158_ ^ ~new__153_;
  assign new__160_ = new__159_ & new__157_;
  assign new__161_ = ~new__160_ ^ ~new__154_;
  assign new__162_ = new__161_ & new__152_;
  assign new__163_ = ~new__162_ ^ ~new__150_;
  assign new__164_ = ~new__163_;
  assign new__165_ = ~new__087_;
  assign new__166_ = ~new__098_ ^ ~new__165_;
  assign new__167_ = ~new__113_ ^ ~new__103_;
  assign new__168__neg = ~new__167_ ^ ~new__166_;
  assign new__168_ = ~new__168__neg;
  assign new__169_ = new__167_ & new__166_;
  assign new__170_ = ~new__169_;
  assign new__171_ = ~new__094_;
  assign new__172_ = ~new__120_ ^ ~new__171_;
  assign new__173_ = ~new__172_ ^ ~new__169_;
  assign new__174_ = ~new__125_ ^ ~new__109_;
  assign new__175_ = ~new__174_ ^ ~new__169_;
  assign new__176_ = new__175_ & new__173_;
  assign new__177_ = ~new__176_ ^ ~new__170_;
  assign new__178_ = new__177_ & new__168_;
  assign new__179_ = ~new__178_ ^ ~new__166_;
  assign new__180__neg = ~new__179_ ^ ~new__163_;
  assign new__180_ = ~new__180__neg;
  assign new__181_ = new__179_ & new__163_;
  assign new__182_ = ~new__181_;
  assign new__183__neg = ~new__174_ ^ ~new__172_;
  assign new__183_ = ~new__183__neg;
  assign new__184_ = new__183_ & new__177_;
  assign new__185_ = ~new__184_ ^ ~new__172_;
  assign new__186_ = ~new__185_ ^ ~new__181_;
  assign new__187_ = ~new__156_;
  assign new__188__neg = ~new__158_ ^ ~new__156_;
  assign new__188_ = ~new__188__neg;
  assign new__189_ = new__188_ & new__161_;
  assign new__190_ = ~new__189_ ^ ~new__187_;
  assign new__191_ = ~new__190_ ^ ~new__181_;
  assign new__192_ = new__191_ & new__186_;
  assign new__193_ = ~new__192_ ^ ~new__182_;
  assign new__194_ = new__193_ & new__180_;
  assign new__195_ = ~new__194_ ^ ~new__164_;
  assign new__196__neg = ~new__195_ ^ ~new__147_;
  assign new__196_ = ~new__196__neg;
  assign new__197_ = new__195_ & new__147_;
  assign new__198_ = ~new__197_;
  assign new__199_ = ~new__190_;
  assign new__200__neg = ~new__190_ ^ ~new__185_;
  assign new__200_ = ~new__200__neg;
  assign new__201_ = new__200_ & new__193_;
  assign new__202_ = ~new__201_ ^ ~new__199_;
  assign new__203_ = ~new__202_ ^ ~new__197_;
  assign new__204__neg = ~new__142_ ^ ~new__137_;
  assign new__204_ = ~new__204__neg;
  assign new__205_ = new__204_ & new__145_;
  assign new__206_ = ~new__205_ ^ ~new__142_;
  assign new__207_ = ~new__206_ ^ ~new__197_;
  assign new__208_ = new__207_ & new__203_;
  assign new__209_ = ~new__208_ ^ ~new__198_;
  assign new__210_ = new__209_ & new__196_;
  assign \out_array[8]  = ~new__210_ ^ ~new__147_;
  assign new__211_ = ~new__195_;
  assign \out_array[10]  = ~new__210_ ^ ~new__211_;
  assign new__212__neg = ~new__206_ ^ ~new__202_;
  assign new__212_ = ~new__212__neg;
  assign new__213_ = new__212_ & new__209_;
  assign \out_array[9]  = ~new__213_ ^ ~new__206_;
  assign new__214_ = ~new__131_;
  assign new__215_ = ~new__146_ ^ ~new__214_;
  assign new__216_ = ~new__194_ ^ ~new__179_;
  assign new__217__neg = ~new__216_ ^ ~new__215_;
  assign new__217_ = ~new__217__neg;
  assign new__218_ = new__216_ & new__215_;
  assign new__219_ = ~new__218_;
  assign new__220_ = ~new__201_ ^ ~new__185_;
  assign new__221_ = ~new__220_ ^ ~new__218_;
  assign new__222_ = ~new__137_;
  assign new__223_ = ~new__205_ ^ ~new__222_;
  assign new__224_ = ~new__223_ ^ ~new__218_;
  assign new__225_ = new__224_ & new__221_;
  assign new__226_ = ~new__225_ ^ ~new__219_;
  assign new__228_ = new__226_ & new__217_;
  assign \out_array[12]  = ~new__228_ ^ ~new__215_;
  assign new__229_ = ~new__216_;
  assign \out_array[14]  = ~new__228_ ^ ~new__229_;
  assign new__230__neg = ~new__223_ ^ ~new__220_;
  assign new__230_ = ~new__230__neg;
  assign new__231_ = new__230_ & new__226_;
  assign \out_array[13]  = ~new__231_ ^ ~new__223_;
  assign new__232_ = ~new__202_;
  assign \out_array[11]  = ~new__213_ ^ ~new__232_;
  assign new__233_ = ~new__220_;
  assign \out_array[15]  = ~new__231_ ^ ~new__233_;
  assign new__235_ = ~new__083_ ^ ~new__065_;
  assign new__236_ = ~new__114_;
  assign new__237_ = ~new__130_ ^ ~new__236_;
  assign new__238__neg = ~new__237_ ^ ~new__235_;
  assign new__238_ = ~new__238__neg;
  assign new__239_ = new__237_ & new__235_;
  assign new__240_ = ~new__239_;
  assign new__241_ = ~new__126_;
  assign new__242_ = ~new__136_ ^ ~new__241_;
  assign new__243_ = ~new__242_ ^ ~new__239_;
  assign new__245_ = ~new__141_ ^ ~new__079_;
  assign new__246_ = ~new__245_ ^ ~new__239_;
  assign new__247_ = new__246_ & new__243_;
  assign new__248_ = ~new__247_ ^ ~new__240_;
  assign new__249_ = new__248_ & new__238_;
  assign new__250_ = ~new__249_ ^ ~new__235_;
  assign new__251_ = ~new__162_ ^ ~new__151_;
  assign new__252_ = ~new__251_;
  assign new__253_ = ~new__167_;
  assign new__254_ = ~new__178_ ^ ~new__253_;
  assign new__256__neg = ~new__254_ ^ ~new__251_;
  assign new__256_ = ~new__256__neg;
  assign new__257_ = new__254_ & new__251_;
  assign new__258_ = ~new__257_;
  assign new__259_ = ~new__174_;
  assign new__260_ = ~new__184_ ^ ~new__259_;
  assign new__261_ = ~new__260_ ^ ~new__257_;
  assign new__262_ = ~new__189_ ^ ~new__158_;
  assign new__263_ = ~new__262_ ^ ~new__257_;
  assign new__264_ = new__263_ & new__261_;
  assign new__265_ = ~new__264_ ^ ~new__258_;
  assign new__267_ = new__265_ & new__256_;
  assign new__268_ = ~new__267_ ^ ~new__252_;
  assign new__269__neg = ~new__268_ ^ ~new__250_;
  assign new__269_ = ~new__269__neg;
  assign new__270_ = new__268_ & new__250_;
  assign new__271_ = ~new__270_;
  assign new__272_ = ~new__262_;
  assign new__273__neg = ~new__262_ ^ ~new__260_;
  assign new__273_ = ~new__273__neg;
  assign new__274_ = new__273_ & new__265_;
  assign new__275_ = ~new__274_ ^ ~new__272_;
  assign new__276_ = ~new__275_ ^ ~new__270_;
  assign new__278__neg = ~new__245_ ^ ~new__242_;
  assign new__278_ = ~new__278__neg;
  assign new__279_ = new__278_ & new__248_;
  assign new__280_ = ~new__279_ ^ ~new__245_;
  assign new__281_ = ~new__280_ ^ ~new__270_;
  assign new__282_ = new__281_ & new__276_;
  assign new__283_ = ~new__282_ ^ ~new__271_;
  assign new__284_ = new__283_ & new__269_;
  assign \out_array[0]  = ~new__284_ ^ ~new__250_;
  assign new__285_ = ~new__268_;
  assign \out_array[2]  = ~new__284_ ^ ~new__285_;
  assign new__287__neg = ~new__280_ ^ ~new__275_;
  assign new__287_ = ~new__287__neg;
  assign new__288_ = new__287_ & new__283_;
  assign \out_array[1]  = ~new__288_ ^ ~new__280_;
  assign new__289_ = ~new__237_;
  assign new__290_ = ~new__249_ ^ ~new__289_;
  assign new__291_ = ~new__267_ ^ ~new__254_;
  assign new__292__neg = ~new__291_ ^ ~new__290_;
  assign new__292_ = ~new__292__neg;
  assign new__293_ = new__291_ & new__290_;
  assign new__294_ = ~new__293_;
  assign new__295_ = ~new__274_ ^ ~new__260_;
  assign new__297_ = ~new__295_ ^ ~new__293_;
  assign new__298_ = ~new__242_;
  assign new__299_ = ~new__279_ ^ ~new__298_;
  assign new__300_ = ~new__299_ ^ ~new__293_;
  assign new__301_ = new__300_ & new__297_;
  assign new__302_ = ~new__301_ ^ ~new__294_;
  assign new__303_ = new__302_ & new__292_;
  assign \out_array[4]  = ~new__303_ ^ ~new__290_;
  assign new__304_ = ~new__291_;
  assign \out_array[6]  = ~new__303_ ^ ~new__304_;
  assign new__306__neg = ~new__299_ ^ ~new__295_;
  assign new__306_ = ~new__306__neg;
  assign new__307_ = new__306_ & new__302_;
  assign \out_array[5]  = ~new__307_ ^ ~new__299_;
  assign new__308_ = ~new__275_;
  assign \out_array[3]  = ~new__288_ ^ ~new__308_;
  assign new__309_ = ~new__295_;
  assign \out_array[7]  = ~new__307_ ^ ~new__309_;
  assign new__227_ = ~\in_array[2] ;
  assign new__234_ = ~\in_array[2]  ^ ~\in_array[0] ;
  assign new__244_ = ~\in_array[0] ;
  assign new__255_ = \in_array[2]  & new__244_;
  assign new__266_ = ~new__255_;
  assign new__277_ = ~\in_array[1] ;
  assign new__286_ = ~new__255_ ^ ~new__277_;
  assign new__296_ = ~new__255_ ^ ~\in_array[3] ;
  assign new__305_ = new__296_ & new__286_;
  assign new__310_ = ~new__305_ ^ ~new__266_;
  assign new__311_ = new__310_ & new__234_;
  assign new__312_ = ~new__311_ ^ ~new__227_;
  assign new__313_ = ~\in_array[6]  ^ ~\in_array[4] ;
  assign new__314_ = ~\in_array[4] ;
  assign new__315_ = \in_array[6]  & new__314_;
  assign new__316_ = ~\in_array[5] ;
  assign new__317_ = ~new__315_ ^ ~new__316_;
  assign new__318_ = ~new__315_ ^ ~\in_array[7] ;
  assign new__319_ = new__318_ & new__317_;
  assign new__320_ = ~new__319_ ^ ~new__315_;
  assign new__321_ = new__320_ & new__313_;
  assign new__322_ = ~new__321_ ^ ~\in_array[6] ;
  assign new__323__neg = ~new__322_ ^ ~new__312_;
  assign new__323_ = ~new__323__neg;
  assign new__324_ = new__322_ & new__312_;
  assign new__325_ = ~new__324_;
  assign new__326_ = ~\in_array[3] ;
  assign new__327_ = \in_array[1]  & new__326_;
  assign new__328_ = ~new__327_ ^ ~new__326_;
  assign new__329_ = ~new__328_ ^ ~new__324_;
  assign new__330_ = new__316_ & \in_array[7] ;
  assign new__331_ = ~new__330_ ^ ~\in_array[7] ;
  assign new__332_ = ~new__331_ ^ ~new__324_;
  assign new__333_ = new__332_ & new__329_;
  assign new__334_ = ~new__333_ ^ ~new__325_;
  assign new__335_ = new__334_ & new__323_;
  assign new__336_ = ~new__335_ ^ ~new__312_;
  assign new__337_ = ~new__311_ ^ ~new__244_;
  assign new__338_ = ~new__337_;
  assign new__339_ = ~new__321_ ^ ~\in_array[4] ;
  assign new__340__neg = ~new__339_ ^ ~new__337_;
  assign new__340_ = ~new__340__neg;
  assign new__341_ = new__339_ & new__337_;
  assign new__342_ = ~new__341_;
  assign new__343_ = ~new__327_ ^ ~\in_array[1] ;
  assign new__344_ = ~new__343_;
  assign new__345_ = ~new__344_ ^ ~new__341_;
  assign new__346_ = ~new__330_ ^ ~new__316_;
endmodule


