module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n9 = x6 & x7 ;
  assign n10 = x4 & x5 ;
  assign n11 = ~n9 & ~n10 ;
  assign n22 = ~x1 & x2 ;
  assign n23 = ~x3 & n22 ;
  assign n24 = n11 & n23 ;
  assign n19 = x0 & ~x1 ;
  assign n20 = ~x3 & n19 ;
  assign n21 = n11 & n20 ;
  assign n25 = n24 ^ n21 ;
  assign n16 = ~x0 & ~x2 ;
  assign n17 = n11 & n16 ;
  assign n12 = ~x0 & x1 ;
  assign n13 = ~x2 & x3 ;
  assign n14 = n12 & n13 ;
  assign n15 = n11 & n14 ;
  assign n18 = n17 ^ n15 ;
  assign n26 = n25 ^ n18 ;
  assign n33 = ~x4 & ~x5 ;
  assign n38 = n26 & n33 ;
  assign n28 = ~x0 & ~x1 ;
  assign n29 = ~x2 & ~x3 ;
  assign n30 = n28 & n29 ;
  assign n27 = ~x6 & ~x7 ;
  assign n34 = ~n27 & n33 ;
  assign n35 = ~n30 & n34 ;
  assign n36 = n26 & n35 ;
  assign n31 = n27 & n30 ;
  assign n32 = n26 & n31 ;
  assign n37 = n36 ^ n32 ;
  assign n39 = n38 ^ n37 ;
  assign y0 = n39 ;
endmodule
