module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 ;
  assign n33 = ~x0 & ~x1 ;
  assign n34 = x2 & x3 ;
  assign n35 = n34 ^ x2 ;
  assign n36 = n35 ^ x3 ;
  assign n37 = x4 & x5 ;
  assign n38 = n37 ^ x4 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = ~n36 & ~n39 ;
  assign n41 = n33 & n40 ;
  assign n42 = x10 & x11 ;
  assign n43 = n42 ^ x10 ;
  assign n44 = n43 ^ x11 ;
  assign n45 = x13 & x14 ;
  assign n46 = n45 ^ x13 ;
  assign n47 = n46 ^ x14 ;
  assign n48 = ~n44 & ~n47 ;
  assign n49 = x6 & x7 ;
  assign n50 = n49 ^ x6 ;
  assign n51 = n50 ^ x7 ;
  assign n52 = x8 & x9 ;
  assign n53 = n52 ^ x8 ;
  assign n54 = n53 ^ x9 ;
  assign n55 = ~n51 & ~n54 ;
  assign n56 = n48 & n55 ;
  assign n57 = n41 & n56 ;
  assign n58 = ~x16 & ~x17 ;
  assign n59 = ~x18 & n58 ;
  assign n60 = ~x12 & ~x15 ;
  assign n61 = ~x19 & n60 ;
  assign n62 = n59 & n61 ;
  assign n63 = ~x21 & ~x22 ;
  assign n64 = ~x20 & ~x23 ;
  assign n65 = n63 & n64 ;
  assign n66 = ~x24 & ~x25 ;
  assign n67 = n65 & n66 ;
  assign n68 = n62 & n67 ;
  assign n69 = n57 & n68 ;
  assign n70 = ~x28 & ~x29 ;
  assign n71 = ~x30 & ~x31 ;
  assign n72 = n70 & n71 ;
  assign n76 = x26 & ~x27 ;
  assign n77 = n72 & n76 ;
  assign n78 = n69 & ~n77 ;
  assign n73 = ~x26 & ~x27 ;
  assign n74 = n72 & n73 ;
  assign n75 = ~n69 & ~n74 ;
  assign n79 = n78 ^ n75 ;
  assign n80 = n59 & n60 ;
  assign n81 = x24 & ~x25 ;
  assign n82 = ~x19 & n81 ;
  assign n83 = n65 & n82 ;
  assign n84 = n80 & n83 ;
  assign n85 = n57 & n84 ;
  assign n86 = ~x19 & n66 ;
  assign n87 = n65 & n86 ;
  assign n88 = n80 & n87 ;
  assign n89 = n57 & n88 ;
  assign n90 = n89 ^ n66 ;
  assign n91 = ~n85 & ~n90 ;
  assign n92 = ~n79 & ~n91 ;
  assign n93 = n33 & n60 ;
  assign n94 = n40 & n93 ;
  assign n95 = n56 & n94 ;
  assign n96 = x18 & n58 ;
  assign n97 = n95 & n96 ;
  assign n98 = n97 ^ x18 ;
  assign n99 = ~x19 & n65 ;
  assign n101 = n80 & n99 ;
  assign n102 = n57 & n101 ;
  assign n103 = ~n98 & n102 ;
  assign n100 = ~n98 & n99 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = n95 ^ x16 ;
  assign n106 = ~x17 & ~n105 ;
  assign n107 = n104 & n106 ;
  assign n108 = n92 & n107 ;
  assign n112 = ~n69 & n74 ;
  assign n113 = ~x24 & n65 ;
  assign n114 = n113 ^ n62 ;
  assign n115 = ~n113 & n114 ;
  assign n116 = n115 ^ n62 ;
  assign n117 = n116 ^ n57 ;
  assign n118 = ~n57 & n117 ;
  assign n119 = n118 ^ n115 ;
  assign n120 = n119 ^ n62 ;
  assign n121 = x25 & n120 ;
  assign n122 = n121 ^ x25 ;
  assign n123 = n112 & n122 ;
  assign n124 = n123 ^ n112 ;
  assign n125 = n57 & n80 ;
  assign n126 = x19 & ~n125 ;
  assign n127 = n57 & n62 ;
  assign n128 = n113 & ~n127 ;
  assign n129 = ~n126 & n128 ;
  assign n130 = n124 & n129 ;
  assign n131 = ~x16 & n95 ;
  assign n136 = ~x17 & ~x18 ;
  assign n137 = ~n131 & n136 ;
  assign n138 = n130 & n137 ;
  assign n109 = n104 & ~n105 ;
  assign n110 = n92 & n109 ;
  assign n132 = x17 & ~x18 ;
  assign n133 = n131 & n132 ;
  assign n134 = ~n110 & n133 ;
  assign n135 = n130 & n134 ;
  assign n139 = n138 ^ n135 ;
  assign n111 = ~x17 & n110 ;
  assign n140 = n139 ^ n111 ;
  assign n142 = n58 & n95 ;
  assign n143 = ~x18 & ~n142 ;
  assign n144 = x17 & ~n131 ;
  assign n145 = n143 & ~n144 ;
  assign n146 = n130 & n145 ;
  assign n141 = n92 & n104 ;
  assign n147 = n146 ^ n141 ;
  assign n148 = ~n108 & n147 ;
  assign n149 = n130 & n141 ;
  assign n150 = n145 ^ n141 ;
  assign n151 = n130 & n150 ;
  assign n152 = n151 ^ n130 ;
  assign n153 = n152 ^ n141 ;
  assign n154 = n149 & n153 ;
  assign n155 = n154 ^ n153 ;
  assign n156 = ~n130 & n141 ;
  assign n157 = ~x23 & n63 ;
  assign n158 = n127 ^ x20 ;
  assign n159 = n157 & n158 ;
  assign n160 = n159 ^ n157 ;
  assign n161 = n92 & n160 ;
  assign n162 = n156 & n161 ;
  assign n163 = n162 ^ n130 ;
  assign n164 = n163 ^ n161 ;
  assign n165 = n130 & ~n161 ;
  assign n166 = ~x22 & ~x23 ;
  assign n167 = ~x24 & n166 ;
  assign n168 = n57 ^ x20 ;
  assign n169 = n62 ^ x20 ;
  assign n170 = ~n62 & ~n169 ;
  assign n171 = n170 ^ x20 ;
  assign n172 = ~n168 & n171 ;
  assign n173 = n172 ^ n170 ;
  assign n174 = n173 ^ n57 ;
  assign n175 = n174 ^ x21 ;
  assign n176 = n175 ^ n167 ;
  assign n177 = ~n167 & ~n176 ;
  assign n178 = n177 ^ n175 ;
  assign n179 = n178 ^ n124 ;
  assign n180 = ~n124 & ~n179 ;
  assign n181 = n180 ^ n177 ;
  assign n182 = n181 ^ n175 ;
  assign n183 = n165 & ~n182 ;
  assign n184 = n183 ^ n161 ;
  assign n185 = n184 ^ n182 ;
  assign n186 = x21 & n174 ;
  assign n187 = n186 ^ n174 ;
  assign n188 = n187 ^ x22 ;
  assign n189 = x23 & n188 ;
  assign n190 = n189 ^ n188 ;
  assign n191 = n190 ^ x23 ;
  assign n192 = ~n161 & ~n191 ;
  assign n194 = n91 & n124 ;
  assign n196 = n194 ^ n92 ;
  assign n197 = n196 ^ n194 ;
  assign n193 = ~x24 & ~n175 ;
  assign n195 = n194 ^ n193 ;
  assign n198 = n197 ^ n195 ;
  assign n199 = n197 ^ n194 ;
  assign n200 = ~n198 & n199 ;
  assign n201 = n200 ^ n197 ;
  assign n202 = n192 & n201 ;
  assign n203 = ~x22 & n187 ;
  assign n204 = x23 & ~n203 ;
  assign n205 = ~x24 & ~n102 ;
  assign n206 = n124 & n205 ;
  assign n207 = ~n204 & n206 ;
  assign n208 = n191 & n207 ;
  assign n209 = n92 & ~n207 ;
  assign n210 = ~n79 & n91 ;
  assign n211 = ~n124 & n210 ;
  assign n212 = ~x26 & n33 ;
  assign n213 = n40 & n212 ;
  assign n214 = n56 & n213 ;
  assign n215 = n68 & n214 ;
  assign n216 = ~n76 & ~n215 ;
  assign n217 = ~x27 & n69 ;
  assign n218 = n72 & ~n217 ;
  assign n219 = ~n216 & n218 ;
  assign n220 = x27 & ~x28 ;
  assign n221 = ~n215 & n220 ;
  assign n222 = ~x27 & n215 ;
  assign n223 = x28 & n222 ;
  assign n224 = ~n221 & ~n223 ;
  assign n225 = ~x29 & n71 ;
  assign n226 = ~n224 & n225 ;
  assign n227 = x29 & ~n222 ;
  assign n228 = ~n70 & n71 ;
  assign n229 = ~n223 & n228 ;
  assign n230 = ~n227 & n229 ;
  assign n231 = ~x27 & ~x28 ;
  assign n232 = n215 & n231 ;
  assign n235 = x30 & ~x31 ;
  assign n236 = ~x29 & n235 ;
  assign n237 = n232 & n236 ;
  assign n233 = x29 & n71 ;
  assign n234 = ~n232 & n233 ;
  assign n238 = n237 ^ n234 ;
  assign n239 = ~x29 & ~n235 ;
  assign n240 = n231 & n239 ;
  assign n241 = n215 & n240 ;
  assign n242 = n241 ^ n235 ;
  assign n243 = ~x30 & x31 ;
  assign n244 = ~x29 & ~n243 ;
  assign n245 = n231 & n244 ;
  assign n246 = n215 & n245 ;
  assign n247 = n242 & ~n246 ;
  assign y0 = n108 ;
  assign y1 = n140 ;
  assign y2 = n148 ;
  assign y3 = n155 ;
  assign y4 = n164 ;
  assign y5 = ~n185 ;
  assign y6 = n202 ;
  assign y7 = n208 ;
  assign y8 = n209 ;
  assign y9 = n194 ;
  assign y10 = n211 ;
  assign y11 = n219 ;
  assign y12 = n226 ;
  assign y13 = n230 ;
  assign y14 = n238 ;
  assign y15 = n247 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
  assign y30 = 1'b0 ;
  assign y31 = 1'b0 ;
endmodule
