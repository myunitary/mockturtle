module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 ;
  assign n485 = x8 ^ x0 ;
  assign n486 = x9 ^ x1 ;
  assign n487 = ~n485 & ~n486 ;
  assign n480 = x10 ^ x2 ;
  assign n496 = x11 ^ x3 ;
  assign n497 = ~n480 & ~n496 ;
  assign n498 = n487 & n497 ;
  assign n516 = x4 & ~x12 ;
  assign n499 = x12 ^ x4 ;
  assign n514 = x5 & ~x13 ;
  assign n515 = ~n499 & n514 ;
  assign n517 = n516 ^ n515 ;
  assign n500 = x13 ^ x5 ;
  assign n501 = ~n499 & ~n500 ;
  assign n511 = x6 & ~x14 ;
  assign n502 = x14 ^ x6 ;
  assign n509 = x7 & ~x15 ;
  assign n510 = ~n502 & n509 ;
  assign n512 = n511 ^ n510 ;
  assign n513 = n501 & n512 ;
  assign n518 = n517 ^ n513 ;
  assign n1100 = n498 & n518 ;
  assign n483 = x2 & ~x10 ;
  assign n481 = x3 & ~x11 ;
  assign n482 = ~n480 & n481 ;
  assign n484 = n483 ^ n482 ;
  assign n1098 = n484 & n487 ;
  assign n492 = x0 & ~x8 ;
  assign n490 = x1 & ~x9 ;
  assign n491 = ~n485 & n490 ;
  assign n493 = n492 ^ n491 ;
  assign n1099 = n1098 ^ n493 ;
  assign n1101 = n1100 ^ n1099 ;
  assign n503 = x15 ^ x7 ;
  assign n504 = ~n502 & ~n503 ;
  assign n505 = n501 & n504 ;
  assign n506 = n498 & n505 ;
  assign n1102 = n1101 ^ n506 ;
  assign n1104 = x0 & ~n1102 ;
  assign n1103 = x8 & n1102 ;
  assign n1105 = n1104 ^ n1103 ;
  assign n528 = x8 & n498 ;
  assign n529 = n518 & n528 ;
  assign n526 = x8 & ~n506 ;
  assign n524 = x8 & n493 ;
  assign n522 = x8 & n487 ;
  assign n523 = n484 & n522 ;
  assign n525 = n524 ^ n523 ;
  assign n527 = n526 ^ n525 ;
  assign n530 = n529 ^ n527 ;
  assign n519 = x0 & n498 ;
  assign n520 = n518 & n519 ;
  assign n507 = x0 & ~n506 ;
  assign n494 = x0 & ~n493 ;
  assign n488 = x0 & n487 ;
  assign n489 = n484 & n488 ;
  assign n495 = n494 ^ n489 ;
  assign n508 = n507 ^ n495 ;
  assign n521 = n520 ^ n508 ;
  assign n531 = n530 ^ n521 ;
  assign n52 = x16 & ~x24 ;
  assign n49 = x24 ^ x16 ;
  assign n50 = x17 & ~x25 ;
  assign n51 = ~n49 & n50 ;
  assign n53 = n52 ^ n51 ;
  assign n475 = x16 & n53 ;
  assign n58 = x18 & ~x26 ;
  assign n55 = x26 ^ x18 ;
  assign n56 = x19 & ~x27 ;
  assign n57 = ~n55 & n56 ;
  assign n59 = n58 ^ n57 ;
  assign n60 = x25 ^ x17 ;
  assign n61 = ~n49 & ~n60 ;
  assign n216 = x16 & n61 ;
  assign n217 = n59 & n216 ;
  assign n476 = n475 ^ n217 ;
  assign n65 = x27 ^ x19 ;
  assign n66 = ~n55 & ~n65 ;
  assign n67 = n61 & n66 ;
  assign n68 = x28 ^ x20 ;
  assign n69 = x29 ^ x21 ;
  assign n70 = ~n68 & ~n69 ;
  assign n71 = x30 ^ x22 ;
  assign n72 = x31 ^ x23 ;
  assign n73 = ~n71 & ~n72 ;
  assign n74 = n70 & n73 ;
  assign n75 = n67 & n74 ;
  assign n219 = x16 & ~n75 ;
  assign n477 = n476 ^ n219 ;
  assign n85 = x20 & ~x28 ;
  assign n83 = x21 & ~x29 ;
  assign n84 = ~n68 & n83 ;
  assign n86 = n85 ^ n84 ;
  assign n80 = x22 & ~x30 ;
  assign n78 = x23 & ~x31 ;
  assign n79 = ~n71 & n78 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = n70 & n81 ;
  assign n87 = n86 ^ n82 ;
  assign n221 = x16 & n67 ;
  assign n222 = n87 & n221 ;
  assign n478 = n477 ^ n222 ;
  assign n471 = x24 & ~n53 ;
  assign n225 = x24 & n61 ;
  assign n226 = n59 & n225 ;
  assign n472 = n471 ^ n226 ;
  assign n228 = x24 & ~n75 ;
  assign n473 = n472 ^ n228 ;
  assign n230 = x24 & n67 ;
  assign n231 = n87 & n230 ;
  assign n474 = n473 ^ n231 ;
  assign n479 = n478 ^ n474 ;
  assign n563 = ~n479 & n531 ;
  assign n532 = n531 ^ n479 ;
  assign n548 = x9 & n498 ;
  assign n549 = n518 & n548 ;
  assign n546 = x9 & ~n506 ;
  assign n544 = x9 & n493 ;
  assign n542 = x9 & n487 ;
  assign n543 = n484 & n542 ;
  assign n545 = n544 ^ n543 ;
  assign n547 = n546 ^ n545 ;
  assign n550 = n549 ^ n547 ;
  assign n539 = x1 & n498 ;
  assign n540 = n518 & n539 ;
  assign n537 = x1 & ~n506 ;
  assign n535 = x1 & ~n493 ;
  assign n533 = x1 & n487 ;
  assign n534 = n484 & n533 ;
  assign n536 = n535 ^ n534 ;
  assign n538 = n537 ^ n536 ;
  assign n541 = n540 ^ n538 ;
  assign n551 = n550 ^ n541 ;
  assign n556 = x17 & n53 ;
  assign n236 = x17 & n61 ;
  assign n237 = n59 & n236 ;
  assign n557 = n556 ^ n237 ;
  assign n239 = x17 & ~n75 ;
  assign n558 = n557 ^ n239 ;
  assign n241 = x17 & n67 ;
  assign n242 = n87 & n241 ;
  assign n559 = n558 ^ n242 ;
  assign n552 = x25 & ~n53 ;
  assign n245 = x25 & n61 ;
  assign n246 = n59 & n245 ;
  assign n553 = n552 ^ n246 ;
  assign n248 = x25 & ~n75 ;
  assign n554 = n553 ^ n248 ;
  assign n250 = x25 & n67 ;
  assign n251 = n87 & n250 ;
  assign n555 = n554 ^ n251 ;
  assign n560 = n559 ^ n555 ;
  assign n561 = n551 & ~n560 ;
  assign n562 = ~n532 & n561 ;
  assign n564 = n563 ^ n562 ;
  assign n1110 = n531 & n564 ;
  assign n580 = x10 & n498 ;
  assign n581 = n518 & n580 ;
  assign n578 = x10 & ~n506 ;
  assign n576 = x10 & n493 ;
  assign n574 = x10 & n487 ;
  assign n575 = n484 & n574 ;
  assign n577 = n576 ^ n575 ;
  assign n579 = n578 ^ n577 ;
  assign n582 = n581 ^ n579 ;
  assign n571 = x2 & n498 ;
  assign n572 = n518 & n571 ;
  assign n569 = x2 & ~n506 ;
  assign n567 = x2 & ~n493 ;
  assign n565 = x2 & n487 ;
  assign n566 = n484 & n565 ;
  assign n568 = n567 ^ n566 ;
  assign n570 = n569 ^ n568 ;
  assign n573 = n572 ^ n570 ;
  assign n583 = n582 ^ n573 ;
  assign n589 = x18 & n53 ;
  assign n62 = x18 & n61 ;
  assign n63 = n59 & n62 ;
  assign n590 = n589 ^ n63 ;
  assign n76 = x18 & ~n75 ;
  assign n591 = n590 ^ n76 ;
  assign n88 = x18 & n67 ;
  assign n89 = n87 & n88 ;
  assign n592 = n591 ^ n89 ;
  assign n585 = x26 & ~n53 ;
  assign n92 = x26 & n61 ;
  assign n93 = n59 & n92 ;
  assign n586 = n585 ^ n93 ;
  assign n95 = x26 & ~n75 ;
  assign n587 = n586 ^ n95 ;
  assign n97 = x26 & n67 ;
  assign n98 = n87 & n97 ;
  assign n588 = n587 ^ n98 ;
  assign n593 = n592 ^ n588 ;
  assign n625 = n583 & ~n593 ;
  assign n594 = n593 ^ n583 ;
  assign n599 = x19 & n53 ;
  assign n174 = x19 & n61 ;
  assign n175 = n59 & n174 ;
  assign n600 = n599 ^ n175 ;
  assign n177 = x19 & ~n75 ;
  assign n601 = n600 ^ n177 ;
  assign n179 = x19 & n67 ;
  assign n180 = n87 & n179 ;
  assign n602 = n601 ^ n180 ;
  assign n595 = x27 & ~n53 ;
  assign n183 = x27 & n61 ;
  assign n184 = n59 & n183 ;
  assign n596 = n595 ^ n184 ;
  assign n186 = x27 & ~n75 ;
  assign n597 = n596 ^ n186 ;
  assign n188 = x27 & n67 ;
  assign n189 = n87 & n188 ;
  assign n598 = n597 ^ n189 ;
  assign n603 = n602 ^ n598 ;
  assign n619 = x11 & n498 ;
  assign n620 = n518 & n619 ;
  assign n617 = x11 & ~n506 ;
  assign n615 = x11 & n493 ;
  assign n613 = x11 & n487 ;
  assign n614 = n484 & n613 ;
  assign n616 = n615 ^ n614 ;
  assign n618 = n617 ^ n616 ;
  assign n621 = n620 ^ n618 ;
  assign n610 = x3 & n498 ;
  assign n611 = n518 & n610 ;
  assign n608 = x3 & ~n506 ;
  assign n606 = x3 & ~n493 ;
  assign n604 = x3 & n487 ;
  assign n605 = n484 & n604 ;
  assign n607 = n606 ^ n605 ;
  assign n609 = n608 ^ n607 ;
  assign n612 = n611 ^ n609 ;
  assign n622 = n621 ^ n612 ;
  assign n623 = ~n603 & n622 ;
  assign n624 = ~n594 & n623 ;
  assign n626 = n625 ^ n624 ;
  assign n627 = n560 ^ n551 ;
  assign n628 = ~n532 & ~n627 ;
  assign n843 = n531 & n628 ;
  assign n844 = n626 & n843 ;
  assign n1111 = n1110 ^ n844 ;
  assign n632 = n622 ^ n603 ;
  assign n633 = ~n594 & ~n632 ;
  assign n634 = n628 & n633 ;
  assign n658 = x20 & n53 ;
  assign n287 = x20 & n61 ;
  assign n288 = n59 & n287 ;
  assign n659 = n658 ^ n288 ;
  assign n290 = x20 & ~n75 ;
  assign n660 = n659 ^ n290 ;
  assign n292 = x20 & n67 ;
  assign n293 = n87 & n292 ;
  assign n661 = n660 ^ n293 ;
  assign n654 = x28 & ~n53 ;
  assign n296 = x28 & n61 ;
  assign n297 = n59 & n296 ;
  assign n655 = n654 ^ n297 ;
  assign n299 = x28 & ~n75 ;
  assign n656 = n655 ^ n299 ;
  assign n301 = x28 & n67 ;
  assign n302 = n87 & n301 ;
  assign n657 = n656 ^ n302 ;
  assign n662 = n661 ^ n657 ;
  assign n650 = x12 & n498 ;
  assign n651 = n518 & n650 ;
  assign n648 = x12 & ~n506 ;
  assign n646 = x12 & n493 ;
  assign n644 = x12 & n487 ;
  assign n645 = n484 & n644 ;
  assign n647 = n646 ^ n645 ;
  assign n649 = n648 ^ n647 ;
  assign n652 = n651 ^ n649 ;
  assign n641 = x4 & n498 ;
  assign n642 = n518 & n641 ;
  assign n639 = x4 & ~n506 ;
  assign n637 = x4 & ~n493 ;
  assign n635 = x4 & n487 ;
  assign n636 = n484 & n635 ;
  assign n638 = n637 ^ n636 ;
  assign n640 = n639 ^ n638 ;
  assign n643 = n642 ^ n640 ;
  assign n653 = n652 ^ n643 ;
  assign n663 = n662 ^ n653 ;
  assign n687 = x21 & n53 ;
  assign n326 = x21 & n61 ;
  assign n327 = n59 & n326 ;
  assign n688 = n687 ^ n327 ;
  assign n329 = x21 & ~n75 ;
  assign n689 = n688 ^ n329 ;
  assign n331 = x21 & n67 ;
  assign n332 = n87 & n331 ;
  assign n690 = n689 ^ n332 ;
  assign n683 = x29 & ~n53 ;
  assign n335 = x29 & n61 ;
  assign n336 = n59 & n335 ;
  assign n684 = n683 ^ n336 ;
  assign n338 = x29 & ~n75 ;
  assign n685 = n684 ^ n338 ;
  assign n340 = x29 & n67 ;
  assign n341 = n87 & n340 ;
  assign n686 = n685 ^ n341 ;
  assign n691 = n690 ^ n686 ;
  assign n679 = x13 & n498 ;
  assign n680 = n518 & n679 ;
  assign n677 = x13 & ~n506 ;
  assign n675 = x13 & n493 ;
  assign n673 = x13 & n487 ;
  assign n674 = n484 & n673 ;
  assign n676 = n675 ^ n674 ;
  assign n678 = n677 ^ n676 ;
  assign n681 = n680 ^ n678 ;
  assign n670 = x5 & n498 ;
  assign n671 = n518 & n670 ;
  assign n668 = x5 & ~n506 ;
  assign n666 = x5 & ~n493 ;
  assign n664 = x5 & n487 ;
  assign n665 = n484 & n664 ;
  assign n667 = n666 ^ n665 ;
  assign n669 = n668 ^ n667 ;
  assign n672 = n671 ^ n669 ;
  assign n682 = n681 ^ n672 ;
  assign n692 = n691 ^ n682 ;
  assign n693 = ~n663 & ~n692 ;
  assign n717 = x22 & n53 ;
  assign n366 = x22 & n61 ;
  assign n367 = n59 & n366 ;
  assign n718 = n717 ^ n367 ;
  assign n369 = x22 & ~n75 ;
  assign n719 = n718 ^ n369 ;
  assign n371 = x22 & n67 ;
  assign n372 = n87 & n371 ;
  assign n720 = n719 ^ n372 ;
  assign n713 = x30 & ~n53 ;
  assign n375 = x30 & n61 ;
  assign n376 = n59 & n375 ;
  assign n714 = n713 ^ n376 ;
  assign n378 = x30 & ~n75 ;
  assign n715 = n714 ^ n378 ;
  assign n380 = x30 & n67 ;
  assign n381 = n87 & n380 ;
  assign n716 = n715 ^ n381 ;
  assign n721 = n720 ^ n716 ;
  assign n709 = x14 & n498 ;
  assign n710 = n518 & n709 ;
  assign n707 = x14 & ~n506 ;
  assign n705 = x14 & n493 ;
  assign n703 = x14 & n487 ;
  assign n704 = n484 & n703 ;
  assign n706 = n705 ^ n704 ;
  assign n708 = n707 ^ n706 ;
  assign n711 = n710 ^ n708 ;
  assign n700 = x6 & n498 ;
  assign n701 = n518 & n700 ;
  assign n698 = x6 & ~n506 ;
  assign n696 = x6 & ~n493 ;
  assign n694 = x6 & n487 ;
  assign n695 = n484 & n694 ;
  assign n697 = n696 ^ n695 ;
  assign n699 = n698 ^ n697 ;
  assign n702 = n701 ^ n699 ;
  assign n712 = n711 ^ n702 ;
  assign n722 = n721 ^ n712 ;
  assign n747 = x15 & n498 ;
  assign n748 = n518 & n747 ;
  assign n745 = x15 & ~n506 ;
  assign n743 = x15 & n493 ;
  assign n741 = x15 & n487 ;
  assign n742 = n484 & n741 ;
  assign n744 = n743 ^ n742 ;
  assign n746 = n745 ^ n744 ;
  assign n749 = n748 ^ n746 ;
  assign n738 = x7 & n498 ;
  assign n739 = n518 & n738 ;
  assign n736 = x7 & ~n506 ;
  assign n734 = x7 & ~n493 ;
  assign n732 = x7 & n487 ;
  assign n733 = n484 & n732 ;
  assign n735 = n734 ^ n733 ;
  assign n737 = n736 ^ n735 ;
  assign n740 = n739 ^ n737 ;
  assign n750 = n749 ^ n740 ;
  assign n727 = x23 & n53 ;
  assign n405 = x23 & n61 ;
  assign n406 = n59 & n405 ;
  assign n728 = n727 ^ n406 ;
  assign n408 = x23 & ~n75 ;
  assign n729 = n728 ^ n408 ;
  assign n410 = x23 & n67 ;
  assign n411 = n87 & n410 ;
  assign n730 = n729 ^ n411 ;
  assign n723 = x31 & ~n53 ;
  assign n414 = x31 & n61 ;
  assign n415 = n59 & n414 ;
  assign n724 = n723 ^ n415 ;
  assign n417 = x31 & ~n75 ;
  assign n725 = n724 ^ n417 ;
  assign n419 = x31 & n67 ;
  assign n420 = n87 & n419 ;
  assign n726 = n725 ^ n420 ;
  assign n731 = n730 ^ n726 ;
  assign n751 = n750 ^ n731 ;
  assign n752 = ~n722 & ~n751 ;
  assign n753 = n693 & n752 ;
  assign n754 = n634 & n753 ;
  assign n846 = n531 & ~n754 ;
  assign n1112 = n1111 ^ n846 ;
  assign n764 = n653 & ~n662 ;
  assign n762 = n682 & ~n691 ;
  assign n763 = ~n663 & n762 ;
  assign n765 = n764 ^ n763 ;
  assign n759 = n712 & ~n721 ;
  assign n757 = ~n731 & n750 ;
  assign n758 = ~n722 & n757 ;
  assign n760 = n759 ^ n758 ;
  assign n761 = n693 & n760 ;
  assign n766 = n765 ^ n761 ;
  assign n848 = n531 & n634 ;
  assign n849 = n766 & n848 ;
  assign n1113 = n1112 ^ n849 ;
  assign n1106 = n479 & ~n564 ;
  assign n852 = n479 & n628 ;
  assign n853 = n626 & n852 ;
  assign n1107 = n1106 ^ n853 ;
  assign n855 = n479 & ~n754 ;
  assign n1108 = n1107 ^ n855 ;
  assign n857 = n479 & n634 ;
  assign n858 = n766 & n857 ;
  assign n1109 = n1108 ^ n858 ;
  assign n1114 = n1113 ^ n1109 ;
  assign n1294 = n1105 & ~n1114 ;
  assign n1115 = n1114 ^ n1105 ;
  assign n1120 = n551 & n564 ;
  assign n882 = n551 & n628 ;
  assign n883 = n626 & n882 ;
  assign n1121 = n1120 ^ n883 ;
  assign n885 = n551 & ~n754 ;
  assign n1122 = n1121 ^ n885 ;
  assign n887 = n551 & n634 ;
  assign n888 = n766 & n887 ;
  assign n1123 = n1122 ^ n888 ;
  assign n1116 = n560 & ~n564 ;
  assign n891 = n560 & n628 ;
  assign n892 = n626 & n891 ;
  assign n1117 = n1116 ^ n892 ;
  assign n894 = n560 & ~n754 ;
  assign n1118 = n1117 ^ n894 ;
  assign n896 = n560 & n634 ;
  assign n897 = n766 & n896 ;
  assign n1119 = n1118 ^ n897 ;
  assign n1124 = n1123 ^ n1119 ;
  assign n1126 = x1 & ~n1102 ;
  assign n1125 = x9 & n1102 ;
  assign n1127 = n1126 ^ n1125 ;
  assign n1292 = ~n1124 & n1127 ;
  assign n1293 = ~n1115 & n1292 ;
  assign n1295 = n1294 ^ n1293 ;
  assign n1128 = n1127 ^ n1124 ;
  assign n1129 = ~n1115 & ~n1128 ;
  assign n1131 = x2 & ~n1102 ;
  assign n1130 = x10 & n1102 ;
  assign n1132 = n1131 ^ n1130 ;
  assign n1137 = n564 & n583 ;
  assign n629 = n583 & n628 ;
  assign n630 = n626 & n629 ;
  assign n1138 = n1137 ^ n630 ;
  assign n755 = n583 & ~n754 ;
  assign n1139 = n1138 ^ n755 ;
  assign n767 = n583 & n634 ;
  assign n768 = n766 & n767 ;
  assign n1140 = n1139 ^ n768 ;
  assign n1133 = ~n564 & n593 ;
  assign n771 = n593 & n628 ;
  assign n772 = n626 & n771 ;
  assign n1134 = n1133 ^ n772 ;
  assign n774 = n593 & ~n754 ;
  assign n1135 = n1134 ^ n774 ;
  assign n776 = n593 & n634 ;
  assign n777 = n766 & n776 ;
  assign n1136 = n1135 ^ n777 ;
  assign n1141 = n1140 ^ n1136 ;
  assign n1289 = n1132 & ~n1141 ;
  assign n1142 = n1141 ^ n1132 ;
  assign n1144 = x3 & ~n1102 ;
  assign n1143 = x11 & n1102 ;
  assign n1145 = n1144 ^ n1143 ;
  assign n1150 = n564 & n622 ;
  assign n801 = n622 & n628 ;
  assign n802 = n626 & n801 ;
  assign n1151 = n1150 ^ n802 ;
  assign n804 = n622 & ~n754 ;
  assign n1152 = n1151 ^ n804 ;
  assign n806 = n622 & n634 ;
  assign n807 = n766 & n806 ;
  assign n1153 = n1152 ^ n807 ;
  assign n1146 = ~n564 & n603 ;
  assign n810 = n603 & n628 ;
  assign n811 = n626 & n810 ;
  assign n1147 = n1146 ^ n811 ;
  assign n813 = n603 & ~n754 ;
  assign n1148 = n1147 ^ n813 ;
  assign n815 = n603 & n634 ;
  assign n816 = n766 & n815 ;
  assign n1149 = n1148 ^ n816 ;
  assign n1154 = n1153 ^ n1149 ;
  assign n1287 = n1145 & ~n1154 ;
  assign n1288 = ~n1142 & n1287 ;
  assign n1290 = n1289 ^ n1288 ;
  assign n1291 = n1129 & n1290 ;
  assign n1296 = n1295 ^ n1291 ;
  assign n1155 = n1154 ^ n1145 ;
  assign n1156 = ~n1142 & ~n1155 ;
  assign n1157 = n1129 & n1156 ;
  assign n1159 = x4 & ~n1102 ;
  assign n1158 = x12 & n1102 ;
  assign n1160 = n1159 ^ n1158 ;
  assign n1165 = n564 & n653 ;
  assign n914 = n628 & n653 ;
  assign n915 = n626 & n914 ;
  assign n1166 = n1165 ^ n915 ;
  assign n917 = n653 & ~n754 ;
  assign n1167 = n1166 ^ n917 ;
  assign n919 = n634 & n653 ;
  assign n920 = n766 & n919 ;
  assign n1168 = n1167 ^ n920 ;
  assign n1161 = ~n564 & n662 ;
  assign n923 = n628 & n662 ;
  assign n924 = n626 & n923 ;
  assign n1162 = n1161 ^ n924 ;
  assign n926 = n662 & ~n754 ;
  assign n1163 = n1162 ^ n926 ;
  assign n928 = n634 & n662 ;
  assign n929 = n766 & n928 ;
  assign n1164 = n1163 ^ n929 ;
  assign n1169 = n1168 ^ n1164 ;
  assign n1283 = n1160 & ~n1169 ;
  assign n1170 = n1169 ^ n1160 ;
  assign n1172 = x5 & ~n1102 ;
  assign n1171 = x13 & n1102 ;
  assign n1173 = n1172 ^ n1171 ;
  assign n1178 = n564 & n682 ;
  assign n953 = n628 & n682 ;
  assign n954 = n626 & n953 ;
  assign n1179 = n1178 ^ n954 ;
  assign n956 = n682 & ~n754 ;
  assign n1180 = n1179 ^ n956 ;
  assign n958 = n634 & n682 ;
  assign n959 = n766 & n958 ;
  assign n1181 = n1180 ^ n959 ;
  assign n1174 = ~n564 & n691 ;
  assign n962 = n628 & n691 ;
  assign n963 = n626 & n962 ;
  assign n1175 = n1174 ^ n963 ;
  assign n965 = n691 & ~n754 ;
  assign n1176 = n1175 ^ n965 ;
  assign n967 = n634 & n691 ;
  assign n968 = n766 & n967 ;
  assign n1177 = n1176 ^ n968 ;
  assign n1182 = n1181 ^ n1177 ;
  assign n1281 = n1173 & ~n1182 ;
  assign n1282 = ~n1170 & n1281 ;
  assign n1284 = n1283 ^ n1282 ;
  assign n1183 = n1182 ^ n1173 ;
  assign n1184 = ~n1170 & ~n1183 ;
  assign n1195 = x6 & ~n1102 ;
  assign n1194 = x14 & n1102 ;
  assign n1196 = n1195 ^ n1194 ;
  assign n1272 = ~n712 & n1196 ;
  assign n1276 = n634 & n1272 ;
  assign n1277 = n766 & n1276 ;
  assign n1218 = n626 & n628 ;
  assign n1219 = n1218 ^ n564 ;
  assign n1274 = ~n1219 & n1272 ;
  assign n1273 = n754 & n1272 ;
  assign n1275 = n1274 ^ n1273 ;
  assign n1278 = n1277 ^ n1275 ;
  assign n1210 = x7 & n1099 ;
  assign n1211 = n1210 ^ n736 ;
  assign n1212 = n1211 ^ n739 ;
  assign n1207 = x15 & ~n1099 ;
  assign n1208 = n1207 ^ n745 ;
  assign n1209 = n1208 ^ n748 ;
  assign n1213 = n1212 ^ n1209 ;
  assign n1237 = ~n731 & n1213 ;
  assign n1244 = n634 & n1237 ;
  assign n1245 = n766 & n1244 ;
  assign n1242 = ~n754 & n1237 ;
  assign n1240 = ~n564 & n1237 ;
  assign n1238 = n628 & n1237 ;
  assign n1239 = n626 & n1238 ;
  assign n1241 = n1240 ^ n1239 ;
  assign n1243 = n1242 ^ n1241 ;
  assign n1246 = n1245 ^ n1243 ;
  assign n1227 = ~n750 & n1213 ;
  assign n1234 = n634 & n1227 ;
  assign n1235 = n766 & n1234 ;
  assign n1232 = ~n754 & n1227 ;
  assign n1230 = n564 & n1227 ;
  assign n1228 = n628 & n1227 ;
  assign n1229 = n626 & n1228 ;
  assign n1231 = n1230 ^ n1229 ;
  assign n1233 = n1232 ^ n1231 ;
  assign n1236 = n1235 ^ n1233 ;
  assign n1247 = n1246 ^ n1236 ;
  assign n1269 = n1196 & n1247 ;
  assign n1264 = n634 & ~n712 ;
  assign n1265 = n766 & n1264 ;
  assign n1262 = ~n712 & ~n754 ;
  assign n1260 = n564 & ~n712 ;
  assign n1258 = n628 & ~n712 ;
  assign n1259 = n626 & n1258 ;
  assign n1261 = n1260 ^ n1259 ;
  assign n1263 = n1262 ^ n1261 ;
  assign n1266 = n1265 ^ n1263 ;
  assign n1267 = n1247 & n1266 ;
  assign n1254 = n634 & ~n721 ;
  assign n1255 = n766 & n1254 ;
  assign n1252 = ~n721 & ~n754 ;
  assign n1250 = ~n564 & ~n721 ;
  assign n1248 = n628 & ~n721 ;
  assign n1249 = n626 & n1248 ;
  assign n1251 = n1250 ^ n1249 ;
  assign n1253 = n1252 ^ n1251 ;
  assign n1256 = n1255 ^ n1253 ;
  assign n1257 = n1247 & n1256 ;
  assign n1268 = n1267 ^ n1257 ;
  assign n1270 = n1269 ^ n1268 ;
  assign n1220 = ~n721 & n1196 ;
  assign n1224 = n634 & n1220 ;
  assign n1225 = n766 & n1224 ;
  assign n1222 = ~n754 & n1220 ;
  assign n1221 = ~n1219 & n1220 ;
  assign n1223 = n1222 ^ n1221 ;
  assign n1226 = n1225 ^ n1223 ;
  assign n1271 = n1270 ^ n1226 ;
  assign n1279 = n1278 ^ n1271 ;
  assign n1280 = n1184 & n1279 ;
  assign n1285 = n1284 ^ n1280 ;
  assign n1286 = n1157 & n1285 ;
  assign n1297 = n1296 ^ n1286 ;
  assign n1189 = n564 & n712 ;
  assign n993 = n628 & n712 ;
  assign n994 = n626 & n993 ;
  assign n1190 = n1189 ^ n994 ;
  assign n996 = n712 & ~n754 ;
  assign n1191 = n1190 ^ n996 ;
  assign n998 = n634 & n712 ;
  assign n999 = n766 & n998 ;
  assign n1192 = n1191 ^ n999 ;
  assign n1185 = ~n564 & n721 ;
  assign n1002 = n628 & n721 ;
  assign n1003 = n626 & n1002 ;
  assign n1186 = n1185 ^ n1003 ;
  assign n1005 = n721 & ~n754 ;
  assign n1187 = n1186 ^ n1005 ;
  assign n1007 = n634 & n721 ;
  assign n1008 = n766 & n1007 ;
  assign n1188 = n1187 ^ n1008 ;
  assign n1193 = n1192 ^ n1188 ;
  assign n1197 = n1196 ^ n1193 ;
  assign n1202 = n564 & n750 ;
  assign n1032 = n628 & n750 ;
  assign n1033 = n626 & n1032 ;
  assign n1203 = n1202 ^ n1033 ;
  assign n1035 = n750 & ~n754 ;
  assign n1204 = n1203 ^ n1035 ;
  assign n1037 = n634 & n750 ;
  assign n1038 = n766 & n1037 ;
  assign n1205 = n1204 ^ n1038 ;
  assign n1198 = ~n564 & n731 ;
  assign n1041 = n628 & n731 ;
  assign n1042 = n626 & n1041 ;
  assign n1199 = n1198 ^ n1042 ;
  assign n1044 = n731 & ~n754 ;
  assign n1200 = n1199 ^ n1044 ;
  assign n1046 = n634 & n731 ;
  assign n1047 = n766 & n1046 ;
  assign n1201 = n1200 ^ n1047 ;
  assign n1206 = n1205 ^ n1201 ;
  assign n1214 = n1213 ^ n1206 ;
  assign n1215 = ~n1197 & ~n1214 ;
  assign n1216 = n1184 & n1215 ;
  assign n1217 = n1157 & n1216 ;
  assign n1298 = n1297 ^ n1217 ;
  assign n1505 = n1105 & ~n1298 ;
  assign n1504 = n1114 & n1298 ;
  assign n1506 = n1505 ^ n1504 ;
  assign n1387 = n1169 & ~n1298 ;
  assign n1386 = n1160 & n1298 ;
  assign n1388 = n1387 ^ n1386 ;
  assign n922 = n564 & n662 ;
  assign n925 = n924 ^ n922 ;
  assign n927 = n926 ^ n925 ;
  assign n930 = n929 ^ n927 ;
  assign n913 = ~n564 & n653 ;
  assign n916 = n915 ^ n913 ;
  assign n918 = n917 ^ n916 ;
  assign n921 = n920 ^ n918 ;
  assign n931 = n930 ^ n921 ;
  assign n295 = x28 & n53 ;
  assign n298 = n297 ^ n295 ;
  assign n300 = n299 ^ n298 ;
  assign n303 = n302 ^ n300 ;
  assign n286 = x20 & ~n53 ;
  assign n289 = n288 ^ n286 ;
  assign n291 = n290 ^ n289 ;
  assign n294 = n293 ^ n291 ;
  assign n304 = n303 ^ n294 ;
  assign n137 = x36 & ~x44 ;
  assign n120 = x44 ^ x36 ;
  assign n135 = x37 & ~x45 ;
  assign n136 = ~n120 & n135 ;
  assign n138 = n137 ^ n136 ;
  assign n121 = x45 ^ x37 ;
  assign n122 = ~n120 & ~n121 ;
  assign n132 = x38 & ~x46 ;
  assign n123 = x46 ^ x38 ;
  assign n130 = x39 & ~x47 ;
  assign n131 = ~n123 & n130 ;
  assign n133 = n132 ^ n131 ;
  assign n134 = n122 & n133 ;
  assign n139 = n138 ^ n134 ;
  assign n106 = x40 ^ x32 ;
  assign n107 = x41 ^ x33 ;
  assign n108 = ~n106 & ~n107 ;
  assign n101 = x42 ^ x34 ;
  assign n117 = x43 ^ x35 ;
  assign n118 = ~n101 & ~n117 ;
  assign n119 = n108 & n118 ;
  assign n320 = x36 & n119 ;
  assign n321 = n139 & n320 ;
  assign n124 = x47 ^ x39 ;
  assign n125 = ~n123 & ~n124 ;
  assign n126 = n122 & n125 ;
  assign n127 = n119 & n126 ;
  assign n318 = x36 & ~n127 ;
  assign n113 = x32 & ~x40 ;
  assign n111 = x33 & ~x41 ;
  assign n112 = ~n106 & n111 ;
  assign n114 = n113 ^ n112 ;
  assign n316 = x36 & n114 ;
  assign n104 = x34 & ~x42 ;
  assign n102 = x35 & ~x43 ;
  assign n103 = ~n101 & n102 ;
  assign n105 = n104 ^ n103 ;
  assign n314 = x36 & n108 ;
  assign n315 = n105 & n314 ;
  assign n317 = n316 ^ n315 ;
  assign n319 = n318 ^ n317 ;
  assign n322 = n321 ^ n319 ;
  assign n311 = x44 & n119 ;
  assign n312 = n139 & n311 ;
  assign n309 = x44 & ~n127 ;
  assign n307 = x44 & ~n114 ;
  assign n305 = x44 & n108 ;
  assign n306 = n105 & n305 ;
  assign n308 = n307 ^ n306 ;
  assign n310 = n309 ^ n308 ;
  assign n313 = n312 ^ n310 ;
  assign n323 = n322 ^ n313 ;
  assign n455 = n304 & ~n323 ;
  assign n324 = n323 ^ n304 ;
  assign n334 = x29 & n53 ;
  assign n337 = n336 ^ n334 ;
  assign n339 = n338 ^ n337 ;
  assign n342 = n341 ^ n339 ;
  assign n325 = x21 & ~n53 ;
  assign n328 = n327 ^ n325 ;
  assign n330 = n329 ^ n328 ;
  assign n333 = n332 ^ n330 ;
  assign n343 = n342 ^ n333 ;
  assign n359 = x37 & n119 ;
  assign n360 = n139 & n359 ;
  assign n357 = x37 & ~n127 ;
  assign n355 = x37 & n114 ;
  assign n353 = x37 & n108 ;
  assign n354 = n105 & n353 ;
  assign n356 = n355 ^ n354 ;
  assign n358 = n357 ^ n356 ;
  assign n361 = n360 ^ n358 ;
  assign n350 = x45 & n119 ;
  assign n351 = n139 & n350 ;
  assign n348 = x45 & ~n127 ;
  assign n346 = x45 & ~n114 ;
  assign n344 = x45 & n108 ;
  assign n345 = n105 & n344 ;
  assign n347 = n346 ^ n345 ;
  assign n349 = n348 ^ n347 ;
  assign n352 = n351 ^ n349 ;
  assign n362 = n361 ^ n352 ;
  assign n453 = n343 & ~n362 ;
  assign n454 = ~n324 & n453 ;
  assign n456 = n455 ^ n454 ;
  assign n363 = n362 ^ n343 ;
  assign n364 = ~n324 & ~n363 ;
  assign n374 = x30 & n53 ;
  assign n377 = n376 ^ n374 ;
  assign n379 = n378 ^ n377 ;
  assign n382 = n381 ^ n379 ;
  assign n365 = x22 & ~n53 ;
  assign n368 = n367 ^ n365 ;
  assign n370 = n369 ^ n368 ;
  assign n373 = n372 ^ n370 ;
  assign n383 = n382 ^ n373 ;
  assign n399 = x38 & n119 ;
  assign n400 = n139 & n399 ;
  assign n397 = x38 & ~n127 ;
  assign n395 = x38 & n114 ;
  assign n393 = x38 & n108 ;
  assign n394 = n105 & n393 ;
  assign n396 = n395 ^ n394 ;
  assign n398 = n397 ^ n396 ;
  assign n401 = n400 ^ n398 ;
  assign n390 = x46 & n119 ;
  assign n391 = n139 & n390 ;
  assign n388 = x46 & ~n127 ;
  assign n386 = x46 & ~n114 ;
  assign n384 = x46 & n108 ;
  assign n385 = n105 & n384 ;
  assign n387 = n386 ^ n385 ;
  assign n389 = n388 ^ n387 ;
  assign n392 = n391 ^ n389 ;
  assign n402 = n401 ^ n392 ;
  assign n450 = n383 & ~n402 ;
  assign n403 = n402 ^ n383 ;
  assign n413 = x31 & n53 ;
  assign n416 = n415 ^ n413 ;
  assign n418 = n417 ^ n416 ;
  assign n421 = n420 ^ n418 ;
  assign n404 = x23 & ~n53 ;
  assign n407 = n406 ^ n404 ;
  assign n409 = n408 ^ n407 ;
  assign n412 = n411 ^ n409 ;
  assign n422 = n421 ^ n412 ;
  assign n438 = x39 & n119 ;
  assign n439 = n139 & n438 ;
  assign n436 = x39 & ~n127 ;
  assign n434 = x39 & n114 ;
  assign n432 = x39 & n108 ;
  assign n433 = n105 & n432 ;
  assign n435 = n434 ^ n433 ;
  assign n437 = n436 ^ n435 ;
  assign n440 = n439 ^ n437 ;
  assign n429 = x47 & n119 ;
  assign n430 = n139 & n429 ;
  assign n427 = x47 & ~n127 ;
  assign n425 = x47 & ~n114 ;
  assign n423 = x47 & n108 ;
  assign n424 = n105 & n423 ;
  assign n426 = n425 ^ n424 ;
  assign n428 = n427 ^ n426 ;
  assign n431 = n430 ^ n428 ;
  assign n441 = n440 ^ n431 ;
  assign n448 = n422 & ~n441 ;
  assign n449 = ~n403 & n448 ;
  assign n451 = n450 ^ n449 ;
  assign n452 = n364 & n451 ;
  assign n457 = n456 ^ n452 ;
  assign n224 = x24 & n53 ;
  assign n227 = n226 ^ n224 ;
  assign n229 = n228 ^ n227 ;
  assign n232 = n231 ^ n229 ;
  assign n215 = x16 & ~n53 ;
  assign n218 = n217 ^ n215 ;
  assign n220 = n219 ^ n218 ;
  assign n223 = n222 ^ n220 ;
  assign n233 = n232 ^ n223 ;
  assign n211 = x32 & n119 ;
  assign n212 = n139 & n211 ;
  assign n209 = x32 & ~n127 ;
  assign n207 = x32 & n114 ;
  assign n205 = x32 & n108 ;
  assign n206 = n105 & n205 ;
  assign n208 = n207 ^ n206 ;
  assign n210 = n209 ^ n208 ;
  assign n213 = n212 ^ n210 ;
  assign n202 = x40 & n119 ;
  assign n203 = n139 & n202 ;
  assign n200 = x40 & ~n127 ;
  assign n198 = x40 & ~n114 ;
  assign n196 = x40 & n108 ;
  assign n197 = n105 & n196 ;
  assign n199 = n198 ^ n197 ;
  assign n201 = n200 ^ n199 ;
  assign n204 = n203 ^ n201 ;
  assign n214 = n213 ^ n204 ;
  assign n234 = n233 ^ n214 ;
  assign n269 = x33 & n119 ;
  assign n270 = n139 & n269 ;
  assign n267 = x33 & ~n127 ;
  assign n265 = x33 & n114 ;
  assign n263 = x33 & n108 ;
  assign n264 = n105 & n263 ;
  assign n266 = n265 ^ n264 ;
  assign n268 = n267 ^ n266 ;
  assign n271 = n270 ^ n268 ;
  assign n260 = x41 & n119 ;
  assign n261 = n139 & n260 ;
  assign n258 = x41 & ~n127 ;
  assign n256 = x41 & ~n114 ;
  assign n254 = x41 & n108 ;
  assign n255 = n105 & n254 ;
  assign n257 = n256 ^ n255 ;
  assign n259 = n258 ^ n257 ;
  assign n262 = n261 ^ n259 ;
  assign n272 = n271 ^ n262 ;
  assign n244 = x25 & n53 ;
  assign n247 = n246 ^ n244 ;
  assign n249 = n248 ^ n247 ;
  assign n252 = n251 ^ n249 ;
  assign n235 = x17 & ~n53 ;
  assign n238 = n237 ^ n235 ;
  assign n240 = n239 ^ n238 ;
  assign n243 = n242 ^ n240 ;
  assign n253 = n252 ^ n243 ;
  assign n273 = n272 ^ n253 ;
  assign n274 = ~n234 & ~n273 ;
  assign n149 = x34 & n119 ;
  assign n150 = n139 & n149 ;
  assign n147 = x34 & ~n127 ;
  assign n145 = x34 & n114 ;
  assign n143 = x34 & n108 ;
  assign n144 = n105 & n143 ;
  assign n146 = n145 ^ n144 ;
  assign n148 = n147 ^ n146 ;
  assign n151 = n150 ^ n148 ;
  assign n140 = x42 & n119 ;
  assign n141 = n139 & n140 ;
  assign n128 = x42 & ~n127 ;
  assign n115 = x42 & ~n114 ;
  assign n109 = x42 & n108 ;
  assign n110 = n105 & n109 ;
  assign n116 = n115 ^ n110 ;
  assign n129 = n128 ^ n116 ;
  assign n142 = n141 ^ n129 ;
  assign n152 = n151 ^ n142 ;
  assign n91 = x26 & n53 ;
  assign n94 = n93 ^ n91 ;
  assign n96 = n95 ^ n94 ;
  assign n99 = n98 ^ n96 ;
  assign n54 = x18 & ~n53 ;
  assign n64 = n63 ^ n54 ;
  assign n77 = n76 ^ n64 ;
  assign n90 = n89 ^ n77 ;
  assign n100 = n99 ^ n90 ;
  assign n153 = n152 ^ n100 ;
  assign n182 = x27 & n53 ;
  assign n185 = n184 ^ n182 ;
  assign n187 = n186 ^ n185 ;
  assign n190 = n189 ^ n187 ;
  assign n173 = x19 & ~n53 ;
  assign n176 = n175 ^ n173 ;
  assign n178 = n177 ^ n176 ;
  assign n181 = n180 ^ n178 ;
  assign n191 = n190 ^ n181 ;
  assign n169 = x35 & n119 ;
  assign n170 = n139 & n169 ;
  assign n167 = x35 & ~n127 ;
  assign n165 = x35 & n114 ;
  assign n163 = x35 & n108 ;
  assign n164 = n105 & n163 ;
  assign n166 = n165 ^ n164 ;
  assign n168 = n167 ^ n166 ;
  assign n171 = n170 ^ n168 ;
  assign n160 = x43 & n119 ;
  assign n161 = n139 & n160 ;
  assign n158 = x43 & ~n127 ;
  assign n156 = x43 & ~n114 ;
  assign n154 = x43 & n108 ;
  assign n155 = n105 & n154 ;
  assign n157 = n156 ^ n155 ;
  assign n159 = n158 ^ n157 ;
  assign n162 = n161 ^ n159 ;
  assign n172 = n171 ^ n162 ;
  assign n283 = n191 ^ n172 ;
  assign n284 = ~n153 & ~n283 ;
  assign n285 = n274 & n284 ;
  assign n947 = n285 & n304 ;
  assign n948 = n457 & n947 ;
  assign n442 = n441 ^ n422 ;
  assign n443 = ~n403 & ~n442 ;
  assign n444 = n364 & n443 ;
  assign n445 = n285 & n444 ;
  assign n945 = n304 & ~n445 ;
  assign n279 = ~n214 & n233 ;
  assign n277 = n253 & ~n272 ;
  assign n278 = ~n234 & n277 ;
  assign n280 = n279 ^ n278 ;
  assign n943 = n280 & n304 ;
  assign n194 = n100 & ~n152 ;
  assign n192 = ~n172 & n191 ;
  assign n193 = ~n153 & n192 ;
  assign n195 = n194 ^ n193 ;
  assign n941 = n274 & n304 ;
  assign n942 = n195 & n941 ;
  assign n944 = n943 ^ n942 ;
  assign n946 = n945 ^ n944 ;
  assign n949 = n948 ^ n946 ;
  assign n938 = n285 & n323 ;
  assign n939 = n457 & n938 ;
  assign n936 = n323 & ~n445 ;
  assign n934 = ~n280 & n323 ;
  assign n932 = n274 & n323 ;
  assign n933 = n195 & n932 ;
  assign n935 = n934 ^ n933 ;
  assign n937 = n936 ^ n935 ;
  assign n940 = n939 ^ n937 ;
  assign n950 = n949 ^ n940 ;
  assign n1082 = n931 & ~n950 ;
  assign n951 = n950 ^ n931 ;
  assign n961 = n564 & n691 ;
  assign n964 = n963 ^ n961 ;
  assign n966 = n965 ^ n964 ;
  assign n969 = n968 ^ n966 ;
  assign n952 = ~n564 & n682 ;
  assign n955 = n954 ^ n952 ;
  assign n957 = n956 ^ n955 ;
  assign n960 = n959 ^ n957 ;
  assign n970 = n969 ^ n960 ;
  assign n986 = n285 & n343 ;
  assign n987 = n457 & n986 ;
  assign n984 = n343 & ~n445 ;
  assign n982 = n280 & n343 ;
  assign n980 = n274 & n343 ;
  assign n981 = n195 & n980 ;
  assign n983 = n982 ^ n981 ;
  assign n985 = n984 ^ n983 ;
  assign n988 = n987 ^ n985 ;
  assign n977 = n285 & n362 ;
  assign n978 = n457 & n977 ;
  assign n975 = n362 & ~n445 ;
  assign n973 = ~n280 & n362 ;
  assign n971 = n274 & n362 ;
  assign n972 = n195 & n971 ;
  assign n974 = n973 ^ n972 ;
  assign n976 = n975 ^ n974 ;
  assign n979 = n978 ^ n976 ;
  assign n989 = n988 ^ n979 ;
  assign n1080 = n970 & ~n989 ;
  assign n1081 = ~n951 & n1080 ;
  assign n1083 = n1082 ^ n1081 ;
  assign n990 = n989 ^ n970 ;
  assign n991 = ~n951 & ~n990 ;
  assign n1001 = n564 & n721 ;
  assign n1004 = n1003 ^ n1001 ;
  assign n1006 = n1005 ^ n1004 ;
  assign n1009 = n1008 ^ n1006 ;
  assign n992 = ~n564 & n712 ;
  assign n995 = n994 ^ n992 ;
  assign n997 = n996 ^ n995 ;
  assign n1000 = n999 ^ n997 ;
  assign n1010 = n1009 ^ n1000 ;
  assign n1026 = n285 & n383 ;
  assign n1027 = n457 & n1026 ;
  assign n1024 = n383 & ~n445 ;
  assign n1022 = n280 & n383 ;
  assign n1020 = n274 & n383 ;
  assign n1021 = n195 & n1020 ;
  assign n1023 = n1022 ^ n1021 ;
  assign n1025 = n1024 ^ n1023 ;
  assign n1028 = n1027 ^ n1025 ;
  assign n1017 = n285 & n402 ;
  assign n1018 = n457 & n1017 ;
  assign n1015 = n402 & ~n445 ;
  assign n1013 = ~n280 & n402 ;
  assign n1011 = n274 & n402 ;
  assign n1012 = n195 & n1011 ;
  assign n1014 = n1013 ^ n1012 ;
  assign n1016 = n1015 ^ n1014 ;
  assign n1019 = n1018 ^ n1016 ;
  assign n1029 = n1028 ^ n1019 ;
  assign n1077 = n1010 & ~n1029 ;
  assign n1030 = n1029 ^ n1010 ;
  assign n1040 = n564 & n731 ;
  assign n1043 = n1042 ^ n1040 ;
  assign n1045 = n1044 ^ n1043 ;
  assign n1048 = n1047 ^ n1045 ;
  assign n1031 = ~n564 & n750 ;
  assign n1034 = n1033 ^ n1031 ;
  assign n1036 = n1035 ^ n1034 ;
  assign n1039 = n1038 ^ n1036 ;
  assign n1049 = n1048 ^ n1039 ;
  assign n1065 = n285 & n422 ;
  assign n1066 = n457 & n1065 ;
  assign n1063 = n422 & ~n445 ;
  assign n1061 = n280 & n422 ;
  assign n1059 = n274 & n422 ;
  assign n1060 = n195 & n1059 ;
  assign n1062 = n1061 ^ n1060 ;
  assign n1064 = n1063 ^ n1062 ;
  assign n1067 = n1066 ^ n1064 ;
  assign n1056 = n285 & n441 ;
  assign n1057 = n457 & n1056 ;
  assign n1054 = n441 & ~n445 ;
  assign n1052 = ~n280 & n441 ;
  assign n1050 = n274 & n441 ;
  assign n1051 = n195 & n1050 ;
  assign n1053 = n1052 ^ n1051 ;
  assign n1055 = n1054 ^ n1053 ;
  assign n1058 = n1057 ^ n1055 ;
  assign n1068 = n1067 ^ n1058 ;
  assign n1075 = n1049 & ~n1068 ;
  assign n1076 = ~n1030 & n1075 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1079 = n991 & n1078 ;
  assign n1084 = n1083 ^ n1079 ;
  assign n851 = n479 & n564 ;
  assign n854 = n853 ^ n851 ;
  assign n856 = n855 ^ n854 ;
  assign n859 = n858 ^ n856 ;
  assign n842 = n531 & ~n564 ;
  assign n845 = n844 ^ n842 ;
  assign n847 = n846 ^ n845 ;
  assign n850 = n849 ^ n847 ;
  assign n860 = n859 ^ n850 ;
  assign n838 = n233 & n285 ;
  assign n839 = n457 & n838 ;
  assign n836 = n233 & ~n445 ;
  assign n834 = n233 & n280 ;
  assign n832 = n233 & n274 ;
  assign n833 = n195 & n832 ;
  assign n835 = n834 ^ n833 ;
  assign n837 = n836 ^ n835 ;
  assign n840 = n839 ^ n837 ;
  assign n829 = n214 & n285 ;
  assign n830 = n457 & n829 ;
  assign n827 = n214 & ~n445 ;
  assign n825 = n214 & ~n280 ;
  assign n823 = n214 & n274 ;
  assign n824 = n195 & n823 ;
  assign n826 = n825 ^ n824 ;
  assign n828 = n827 ^ n826 ;
  assign n831 = n830 ^ n828 ;
  assign n841 = n840 ^ n831 ;
  assign n861 = n860 ^ n841 ;
  assign n890 = n560 & n564 ;
  assign n893 = n892 ^ n890 ;
  assign n895 = n894 ^ n893 ;
  assign n898 = n897 ^ n895 ;
  assign n881 = n551 & ~n564 ;
  assign n884 = n883 ^ n881 ;
  assign n886 = n885 ^ n884 ;
  assign n889 = n888 ^ n886 ;
  assign n899 = n898 ^ n889 ;
  assign n877 = n253 & n285 ;
  assign n878 = n457 & n877 ;
  assign n875 = n253 & ~n445 ;
  assign n873 = n253 & n280 ;
  assign n871 = n253 & n274 ;
  assign n872 = n195 & n871 ;
  assign n874 = n873 ^ n872 ;
  assign n876 = n875 ^ n874 ;
  assign n879 = n878 ^ n876 ;
  assign n868 = n272 & n285 ;
  assign n869 = n457 & n868 ;
  assign n866 = n272 & ~n445 ;
  assign n864 = n272 & ~n280 ;
  assign n862 = n272 & n274 ;
  assign n863 = n195 & n862 ;
  assign n865 = n864 ^ n863 ;
  assign n867 = n866 ^ n865 ;
  assign n870 = n869 ^ n867 ;
  assign n880 = n879 ^ n870 ;
  assign n900 = n899 ^ n880 ;
  assign n901 = ~n861 & ~n900 ;
  assign n770 = n564 & n593 ;
  assign n773 = n772 ^ n770 ;
  assign n775 = n774 ^ n773 ;
  assign n778 = n777 ^ n775 ;
  assign n584 = ~n564 & n583 ;
  assign n631 = n630 ^ n584 ;
  assign n756 = n755 ^ n631 ;
  assign n769 = n768 ^ n756 ;
  assign n779 = n778 ^ n769 ;
  assign n467 = n100 & n285 ;
  assign n468 = n457 & n467 ;
  assign n465 = n100 & ~n445 ;
  assign n463 = n100 & n280 ;
  assign n461 = n100 & n274 ;
  assign n462 = n195 & n461 ;
  assign n464 = n463 ^ n462 ;
  assign n466 = n465 ^ n464 ;
  assign n469 = n468 ^ n466 ;
  assign n458 = n152 & n285 ;
  assign n459 = n457 & n458 ;
  assign n446 = n152 & ~n445 ;
  assign n281 = n152 & ~n280 ;
  assign n275 = n152 & n274 ;
  assign n276 = n195 & n275 ;
  assign n282 = n281 ^ n276 ;
  assign n447 = n446 ^ n282 ;
  assign n460 = n459 ^ n447 ;
  assign n470 = n469 ^ n460 ;
  assign n780 = n779 ^ n470 ;
  assign n809 = n564 & n603 ;
  assign n812 = n811 ^ n809 ;
  assign n814 = n813 ^ n812 ;
  assign n817 = n816 ^ n814 ;
  assign n800 = ~n564 & n622 ;
  assign n803 = n802 ^ n800 ;
  assign n805 = n804 ^ n803 ;
  assign n808 = n807 ^ n805 ;
  assign n818 = n817 ^ n808 ;
  assign n796 = n191 & n285 ;
  assign n797 = n457 & n796 ;
  assign n794 = n191 & ~n445 ;
  assign n792 = n191 & n280 ;
  assign n790 = n191 & n274 ;
  assign n791 = n195 & n790 ;
  assign n793 = n792 ^ n791 ;
  assign n795 = n794 ^ n793 ;
  assign n798 = n797 ^ n795 ;
  assign n787 = n172 & n285 ;
  assign n788 = n457 & n787 ;
  assign n785 = n172 & ~n445 ;
  assign n783 = n172 & ~n280 ;
  assign n781 = n172 & n274 ;
  assign n782 = n195 & n781 ;
  assign n784 = n783 ^ n782 ;
  assign n786 = n785 ^ n784 ;
  assign n789 = n788 ^ n786 ;
  assign n799 = n798 ^ n789 ;
  assign n910 = n818 ^ n799 ;
  assign n911 = ~n780 & ~n910 ;
  assign n912 = n901 & n911 ;
  assign n1404 = n912 & n931 ;
  assign n1405 = n1084 & n1404 ;
  assign n1069 = n1068 ^ n1049 ;
  assign n1070 = ~n1030 & ~n1069 ;
  assign n1071 = n991 & n1070 ;
  assign n1072 = n912 & n1071 ;
  assign n1402 = n931 & ~n1072 ;
  assign n906 = ~n841 & n860 ;
  assign n904 = ~n880 & n899 ;
  assign n905 = ~n861 & n904 ;
  assign n907 = n906 ^ n905 ;
  assign n1400 = n907 & n931 ;
  assign n821 = ~n470 & n779 ;
  assign n819 = ~n799 & n818 ;
  assign n820 = ~n780 & n819 ;
  assign n822 = n821 ^ n820 ;
  assign n1398 = n901 & n931 ;
  assign n1399 = n822 & n1398 ;
  assign n1401 = n1400 ^ n1399 ;
  assign n1403 = n1402 ^ n1401 ;
  assign n1406 = n1405 ^ n1403 ;
  assign n1395 = n912 & n950 ;
  assign n1396 = n1084 & n1395 ;
  assign n1393 = n950 & ~n1072 ;
  assign n1391 = ~n907 & n950 ;
  assign n1389 = n901 & n950 ;
  assign n1390 = n822 & n1389 ;
  assign n1392 = n1391 ^ n1390 ;
  assign n1394 = n1393 ^ n1392 ;
  assign n1397 = n1396 ^ n1394 ;
  assign n1407 = n1406 ^ n1397 ;
  assign n1491 = n1388 & ~n1407 ;
  assign n1408 = n1407 ^ n1388 ;
  assign n1410 = n1182 & ~n1298 ;
  assign n1409 = n1173 & n1298 ;
  assign n1411 = n1410 ^ n1409 ;
  assign n1427 = n912 & n970 ;
  assign n1428 = n1084 & n1427 ;
  assign n1425 = n970 & ~n1072 ;
  assign n1423 = n907 & n970 ;
  assign n1421 = n901 & n970 ;
  assign n1422 = n822 & n1421 ;
  assign n1424 = n1423 ^ n1422 ;
  assign n1426 = n1425 ^ n1424 ;
  assign n1429 = n1428 ^ n1426 ;
  assign n1418 = n912 & n989 ;
  assign n1419 = n1084 & n1418 ;
  assign n1416 = n989 & ~n1072 ;
  assign n1414 = ~n907 & n989 ;
  assign n1412 = n901 & n989 ;
  assign n1413 = n822 & n1412 ;
  assign n1415 = n1414 ^ n1413 ;
  assign n1417 = n1416 ^ n1415 ;
  assign n1420 = n1419 ^ n1417 ;
  assign n1430 = n1429 ^ n1420 ;
  assign n1489 = n1411 & ~n1430 ;
  assign n1490 = ~n1408 & n1489 ;
  assign n1492 = n1491 ^ n1490 ;
  assign n1431 = n1430 ^ n1411 ;
  assign n1432 = ~n1408 & ~n1431 ;
  assign n1434 = n1193 & ~n1298 ;
  assign n1433 = n1196 & n1298 ;
  assign n1435 = n1434 ^ n1433 ;
  assign n1451 = n912 & n1010 ;
  assign n1452 = n1084 & n1451 ;
  assign n1449 = n1010 & ~n1072 ;
  assign n1447 = n907 & n1010 ;
  assign n1445 = n901 & n1010 ;
  assign n1446 = n822 & n1445 ;
  assign n1448 = n1447 ^ n1446 ;
  assign n1450 = n1449 ^ n1448 ;
  assign n1453 = n1452 ^ n1450 ;
  assign n1442 = n912 & n1029 ;
  assign n1443 = n1084 & n1442 ;
  assign n1440 = n1029 & ~n1072 ;
  assign n1438 = ~n907 & n1029 ;
  assign n1436 = n901 & n1029 ;
  assign n1437 = n822 & n1436 ;
  assign n1439 = n1438 ^ n1437 ;
  assign n1441 = n1440 ^ n1439 ;
  assign n1444 = n1443 ^ n1441 ;
  assign n1454 = n1453 ^ n1444 ;
  assign n1486 = n1435 & ~n1454 ;
  assign n1455 = n1454 ^ n1435 ;
  assign n1457 = n1206 & ~n1298 ;
  assign n1456 = n1213 & n1298 ;
  assign n1458 = n1457 ^ n1456 ;
  assign n1474 = n912 & n1049 ;
  assign n1475 = n1084 & n1474 ;
  assign n1472 = n1049 & ~n1072 ;
  assign n1470 = n907 & n1049 ;
  assign n1468 = n901 & n1049 ;
  assign n1469 = n822 & n1468 ;
  assign n1471 = n1470 ^ n1469 ;
  assign n1473 = n1472 ^ n1471 ;
  assign n1476 = n1475 ^ n1473 ;
  assign n1465 = n912 & n1068 ;
  assign n1466 = n1084 & n1465 ;
  assign n1463 = n1068 & ~n1072 ;
  assign n1461 = ~n907 & n1068 ;
  assign n1459 = n901 & n1068 ;
  assign n1460 = n822 & n1459 ;
  assign n1462 = n1461 ^ n1460 ;
  assign n1464 = n1463 ^ n1462 ;
  assign n1467 = n1466 ^ n1464 ;
  assign n1477 = n1476 ^ n1467 ;
  assign n1484 = n1458 & ~n1477 ;
  assign n1485 = ~n1455 & n1484 ;
  assign n1487 = n1486 ^ n1485 ;
  assign n1488 = n1432 & n1487 ;
  assign n1493 = n1492 ^ n1488 ;
  assign n1300 = n1114 & ~n1298 ;
  assign n1299 = n1105 & n1298 ;
  assign n1301 = n1300 ^ n1299 ;
  assign n1094 = n860 & n912 ;
  assign n1095 = n1084 & n1094 ;
  assign n1092 = n860 & ~n1072 ;
  assign n1090 = n860 & n907 ;
  assign n1088 = n860 & n901 ;
  assign n1089 = n822 & n1088 ;
  assign n1091 = n1090 ^ n1089 ;
  assign n1093 = n1092 ^ n1091 ;
  assign n1096 = n1095 ^ n1093 ;
  assign n1085 = n841 & n912 ;
  assign n1086 = n1084 & n1085 ;
  assign n1073 = n841 & ~n1072 ;
  assign n908 = n841 & ~n907 ;
  assign n902 = n841 & n901 ;
  assign n903 = n822 & n902 ;
  assign n909 = n908 ^ n903 ;
  assign n1074 = n1073 ^ n909 ;
  assign n1087 = n1086 ^ n1074 ;
  assign n1097 = n1096 ^ n1087 ;
  assign n1302 = n1301 ^ n1097 ;
  assign n1321 = n899 & n912 ;
  assign n1322 = n1084 & n1321 ;
  assign n1319 = n899 & ~n1072 ;
  assign n1317 = n899 & n907 ;
  assign n1315 = n899 & n901 ;
  assign n1316 = n822 & n1315 ;
  assign n1318 = n1317 ^ n1316 ;
  assign n1320 = n1319 ^ n1318 ;
  assign n1323 = n1322 ^ n1320 ;
  assign n1312 = n880 & n912 ;
  assign n1313 = n1084 & n1312 ;
  assign n1310 = n880 & ~n1072 ;
  assign n1308 = n880 & ~n907 ;
  assign n1306 = n880 & n901 ;
  assign n1307 = n822 & n1306 ;
  assign n1309 = n1308 ^ n1307 ;
  assign n1311 = n1310 ^ n1309 ;
  assign n1314 = n1313 ^ n1311 ;
  assign n1324 = n1323 ^ n1314 ;
  assign n1304 = n1124 & ~n1298 ;
  assign n1303 = n1127 & n1298 ;
  assign n1305 = n1304 ^ n1303 ;
  assign n1325 = n1324 ^ n1305 ;
  assign n1326 = ~n1302 & ~n1325 ;
  assign n1345 = n779 & n912 ;
  assign n1346 = n1084 & n1345 ;
  assign n1343 = n779 & ~n1072 ;
  assign n1341 = n779 & n907 ;
  assign n1339 = n779 & n901 ;
  assign n1340 = n822 & n1339 ;
  assign n1342 = n1341 ^ n1340 ;
  assign n1344 = n1343 ^ n1342 ;
  assign n1347 = n1346 ^ n1344 ;
  assign n1336 = n470 & n912 ;
  assign n1337 = n1084 & n1336 ;
  assign n1334 = n470 & ~n1072 ;
  assign n1332 = n470 & ~n907 ;
  assign n1330 = n470 & n901 ;
  assign n1331 = n822 & n1330 ;
  assign n1333 = n1332 ^ n1331 ;
  assign n1335 = n1334 ^ n1333 ;
  assign n1338 = n1337 ^ n1335 ;
  assign n1348 = n1347 ^ n1338 ;
  assign n1328 = n1141 & ~n1298 ;
  assign n1327 = n1132 & n1298 ;
  assign n1329 = n1328 ^ n1327 ;
  assign n1349 = n1348 ^ n1329 ;
  assign n1370 = n1154 & ~n1298 ;
  assign n1369 = n1145 & n1298 ;
  assign n1371 = n1370 ^ n1369 ;
  assign n1365 = n818 & n912 ;
  assign n1366 = n1084 & n1365 ;
  assign n1363 = n818 & ~n1072 ;
  assign n1361 = n818 & n907 ;
  assign n1359 = n818 & n901 ;
  assign n1360 = n822 & n1359 ;
  assign n1362 = n1361 ^ n1360 ;
  assign n1364 = n1363 ^ n1362 ;
  assign n1367 = n1366 ^ n1364 ;
  assign n1356 = n799 & n912 ;
  assign n1357 = n1084 & n1356 ;
  assign n1354 = n799 & ~n1072 ;
  assign n1352 = n799 & ~n907 ;
  assign n1350 = n799 & n901 ;
  assign n1351 = n822 & n1350 ;
  assign n1353 = n1352 ^ n1351 ;
  assign n1355 = n1354 ^ n1353 ;
  assign n1358 = n1357 ^ n1355 ;
  assign n1368 = n1367 ^ n1358 ;
  assign n1383 = n1371 ^ n1368 ;
  assign n1384 = ~n1349 & ~n1383 ;
  assign n1385 = n1326 & n1384 ;
  assign n1500 = n1301 & n1385 ;
  assign n1501 = n1493 & n1500 ;
  assign n1478 = n1477 ^ n1458 ;
  assign n1479 = ~n1455 & ~n1478 ;
  assign n1480 = n1432 & n1479 ;
  assign n1481 = n1385 & n1480 ;
  assign n1498 = n1301 & ~n1481 ;
  assign n1379 = ~n1097 & n1301 ;
  assign n1377 = n1305 & ~n1324 ;
  assign n1378 = ~n1302 & n1377 ;
  assign n1380 = n1379 ^ n1378 ;
  assign n1374 = n1329 & ~n1348 ;
  assign n1372 = ~n1368 & n1371 ;
  assign n1373 = ~n1349 & n1372 ;
  assign n1375 = n1374 ^ n1373 ;
  assign n1376 = n1326 & n1375 ;
  assign n1381 = n1380 ^ n1376 ;
  assign n1497 = n1301 & n1381 ;
  assign n1499 = n1498 ^ n1497 ;
  assign n1502 = n1501 ^ n1499 ;
  assign n1494 = n1097 & n1385 ;
  assign n1495 = n1493 & n1494 ;
  assign n1482 = n1097 & ~n1481 ;
  assign n1382 = n1097 & ~n1381 ;
  assign n1483 = n1482 ^ n1382 ;
  assign n1496 = n1495 ^ n1483 ;
  assign n1503 = n1502 ^ n1496 ;
  assign n1689 = ~n1503 & n1506 ;
  assign n1507 = n1506 ^ n1503 ;
  assign n1509 = n1127 & ~n1298 ;
  assign n1508 = n1124 & n1298 ;
  assign n1510 = n1509 ^ n1508 ;
  assign n1520 = n1305 & n1385 ;
  assign n1521 = n1493 & n1520 ;
  assign n1518 = n1305 & ~n1481 ;
  assign n1517 = n1305 & n1381 ;
  assign n1519 = n1518 ^ n1517 ;
  assign n1522 = n1521 ^ n1519 ;
  assign n1514 = n1324 & n1385 ;
  assign n1515 = n1493 & n1514 ;
  assign n1512 = n1324 & ~n1481 ;
  assign n1511 = n1324 & ~n1381 ;
  assign n1513 = n1512 ^ n1511 ;
  assign n1516 = n1515 ^ n1513 ;
  assign n1523 = n1522 ^ n1516 ;
  assign n1687 = n1510 & ~n1523 ;
  assign n1688 = ~n1507 & n1687 ;
  assign n1690 = n1689 ^ n1688 ;
  assign n1524 = n1523 ^ n1510 ;
  assign n1525 = ~n1507 & ~n1524 ;
  assign n1527 = n1132 & ~n1298 ;
  assign n1526 = n1141 & n1298 ;
  assign n1528 = n1527 ^ n1526 ;
  assign n1538 = n1329 & n1385 ;
  assign n1539 = n1493 & n1538 ;
  assign n1536 = n1329 & ~n1481 ;
  assign n1535 = n1329 & n1381 ;
  assign n1537 = n1536 ^ n1535 ;
  assign n1540 = n1539 ^ n1537 ;
  assign n1532 = n1348 & n1385 ;
  assign n1533 = n1493 & n1532 ;
  assign n1530 = n1348 & ~n1481 ;
  assign n1529 = n1348 & ~n1381 ;
  assign n1531 = n1530 ^ n1529 ;
  assign n1534 = n1533 ^ n1531 ;
  assign n1541 = n1540 ^ n1534 ;
  assign n1684 = n1528 & ~n1541 ;
  assign n1542 = n1541 ^ n1528 ;
  assign n1544 = n1145 & ~n1298 ;
  assign n1543 = n1154 & n1298 ;
  assign n1545 = n1544 ^ n1543 ;
  assign n1555 = n1371 & n1385 ;
  assign n1556 = n1493 & n1555 ;
  assign n1553 = n1371 & ~n1481 ;
  assign n1552 = n1371 & n1381 ;
  assign n1554 = n1553 ^ n1552 ;
  assign n1557 = n1556 ^ n1554 ;
  assign n1549 = n1368 & n1385 ;
  assign n1550 = n1493 & n1549 ;
  assign n1547 = n1368 & ~n1481 ;
  assign n1546 = n1368 & ~n1381 ;
  assign n1548 = n1547 ^ n1546 ;
  assign n1551 = n1550 ^ n1548 ;
  assign n1558 = n1557 ^ n1551 ;
  assign n1682 = n1545 & ~n1558 ;
  assign n1683 = ~n1542 & n1682 ;
  assign n1685 = n1684 ^ n1683 ;
  assign n1686 = n1525 & n1685 ;
  assign n1691 = n1690 ^ n1686 ;
  assign n1559 = n1558 ^ n1545 ;
  assign n1560 = ~n1542 & ~n1559 ;
  assign n1561 = n1525 & n1560 ;
  assign n1563 = n1160 & ~n1298 ;
  assign n1562 = n1169 & n1298 ;
  assign n1564 = n1563 ^ n1562 ;
  assign n1574 = n1385 & n1388 ;
  assign n1575 = n1493 & n1574 ;
  assign n1572 = n1388 & ~n1481 ;
  assign n1571 = n1381 & n1388 ;
  assign n1573 = n1572 ^ n1571 ;
  assign n1576 = n1575 ^ n1573 ;
  assign n1568 = n1385 & n1407 ;
  assign n1569 = n1493 & n1568 ;
  assign n1566 = n1407 & ~n1481 ;
  assign n1565 = ~n1381 & n1407 ;
  assign n1567 = n1566 ^ n1565 ;
  assign n1570 = n1569 ^ n1567 ;
  assign n1577 = n1576 ^ n1570 ;
  assign n1678 = n1564 & ~n1577 ;
  assign n1578 = n1577 ^ n1564 ;
  assign n1580 = n1173 & ~n1298 ;
  assign n1579 = n1182 & n1298 ;
  assign n1581 = n1580 ^ n1579 ;
  assign n1591 = n1385 & n1411 ;
  assign n1592 = n1493 & n1591 ;
  assign n1589 = n1411 & ~n1481 ;
  assign n1588 = n1381 & n1411 ;
  assign n1590 = n1589 ^ n1588 ;
  assign n1593 = n1592 ^ n1590 ;
  assign n1585 = n1385 & n1430 ;
  assign n1586 = n1493 & n1585 ;
  assign n1583 = n1430 & ~n1481 ;
  assign n1582 = ~n1381 & n1430 ;
  assign n1584 = n1583 ^ n1582 ;
  assign n1587 = n1586 ^ n1584 ;
  assign n1594 = n1593 ^ n1587 ;
  assign n1676 = n1581 & ~n1594 ;
  assign n1677 = ~n1578 & n1676 ;
  assign n1679 = n1678 ^ n1677 ;
  assign n1595 = n1594 ^ n1581 ;
  assign n1596 = ~n1578 & ~n1595 ;
  assign n1634 = n1385 & n1493 ;
  assign n1635 = n1634 ^ n1381 ;
  assign n1636 = n1635 ^ n1481 ;
  assign n1611 = n1196 & ~n1298 ;
  assign n1610 = n1193 & n1298 ;
  assign n1612 = n1611 ^ n1610 ;
  assign n1672 = ~n1435 & n1612 ;
  assign n1673 = ~n1636 & n1672 ;
  assign n1628 = n1213 & ~n1298 ;
  assign n1627 = n1206 & n1298 ;
  assign n1629 = n1628 ^ n1627 ;
  assign n1646 = ~n1458 & n1629 ;
  assign n1650 = n1385 & n1646 ;
  assign n1651 = n1493 & n1650 ;
  assign n1648 = ~n1481 & n1646 ;
  assign n1647 = n1381 & n1646 ;
  assign n1649 = n1648 ^ n1647 ;
  assign n1652 = n1651 ^ n1649 ;
  assign n1639 = ~n1477 & n1629 ;
  assign n1643 = n1385 & n1639 ;
  assign n1644 = n1493 & n1643 ;
  assign n1641 = ~n1481 & n1639 ;
  assign n1640 = ~n1381 & n1639 ;
  assign n1642 = n1641 ^ n1640 ;
  assign n1645 = n1644 ^ n1642 ;
  assign n1653 = n1652 ^ n1645 ;
  assign n1669 = n1612 & n1653 ;
  assign n1664 = n1385 & ~n1435 ;
  assign n1665 = n1493 & n1664 ;
  assign n1662 = ~n1435 & ~n1481 ;
  assign n1661 = n1381 & ~n1435 ;
  assign n1663 = n1662 ^ n1661 ;
  assign n1666 = n1665 ^ n1663 ;
  assign n1667 = n1653 & n1666 ;
  assign n1657 = n1385 & ~n1454 ;
  assign n1658 = n1493 & n1657 ;
  assign n1655 = ~n1454 & ~n1481 ;
  assign n1654 = ~n1381 & ~n1454 ;
  assign n1656 = n1655 ^ n1654 ;
  assign n1659 = n1658 ^ n1656 ;
  assign n1660 = n1653 & n1659 ;
  assign n1668 = n1667 ^ n1660 ;
  assign n1670 = n1669 ^ n1668 ;
  assign n1637 = ~n1454 & n1612 ;
  assign n1638 = n1636 & n1637 ;
  assign n1671 = n1670 ^ n1638 ;
  assign n1674 = n1673 ^ n1671 ;
  assign n1675 = n1596 & n1674 ;
  assign n1680 = n1679 ^ n1675 ;
  assign n1681 = n1561 & n1680 ;
  assign n1692 = n1691 ^ n1681 ;
  assign n1606 = n1385 & n1435 ;
  assign n1607 = n1493 & n1606 ;
  assign n1604 = n1435 & ~n1481 ;
  assign n1603 = n1381 & n1435 ;
  assign n1605 = n1604 ^ n1603 ;
  assign n1608 = n1607 ^ n1605 ;
  assign n1600 = n1385 & n1454 ;
  assign n1601 = n1493 & n1600 ;
  assign n1598 = n1454 & ~n1481 ;
  assign n1597 = ~n1381 & n1454 ;
  assign n1599 = n1598 ^ n1597 ;
  assign n1602 = n1601 ^ n1599 ;
  assign n1609 = n1608 ^ n1602 ;
  assign n1613 = n1612 ^ n1609 ;
  assign n1623 = n1385 & n1458 ;
  assign n1624 = n1493 & n1623 ;
  assign n1621 = n1458 & ~n1481 ;
  assign n1620 = n1381 & n1458 ;
  assign n1622 = n1621 ^ n1620 ;
  assign n1625 = n1624 ^ n1622 ;
  assign n1617 = n1385 & n1477 ;
  assign n1618 = n1493 & n1617 ;
  assign n1615 = n1477 & ~n1481 ;
  assign n1614 = ~n1381 & n1477 ;
  assign n1616 = n1615 ^ n1614 ;
  assign n1619 = n1618 ^ n1616 ;
  assign n1626 = n1625 ^ n1619 ;
  assign n1630 = n1629 ^ n1626 ;
  assign n1631 = ~n1613 & ~n1630 ;
  assign n1632 = n1596 & n1631 ;
  assign n1633 = n1561 & n1632 ;
  assign n1693 = n1692 ^ n1633 ;
  assign n1695 = n1506 & ~n1693 ;
  assign n1694 = n1503 & n1693 ;
  assign n1696 = n1695 ^ n1694 ;
  assign n1698 = n1510 & ~n1693 ;
  assign n1697 = n1523 & n1693 ;
  assign n1699 = n1698 ^ n1697 ;
  assign n1701 = n1528 & ~n1693 ;
  assign n1700 = n1541 & n1693 ;
  assign n1702 = n1701 ^ n1700 ;
  assign n1704 = n1545 & ~n1693 ;
  assign n1703 = n1558 & n1693 ;
  assign n1705 = n1704 ^ n1703 ;
  assign n1707 = n1564 & ~n1693 ;
  assign n1706 = n1577 & n1693 ;
  assign n1708 = n1707 ^ n1706 ;
  assign n1710 = n1581 & ~n1693 ;
  assign n1709 = n1594 & n1693 ;
  assign n1711 = n1710 ^ n1709 ;
  assign n1713 = n1612 & ~n1693 ;
  assign n1712 = n1609 & n1693 ;
  assign n1714 = n1713 ^ n1712 ;
  assign n1716 = n1629 & ~n1693 ;
  assign n1715 = n1626 & n1693 ;
  assign n1717 = n1716 ^ n1715 ;
  assign n1719 = n1503 & ~n1693 ;
  assign n1718 = n1506 & n1693 ;
  assign n1720 = n1719 ^ n1718 ;
  assign n1722 = n1523 & ~n1693 ;
  assign n1721 = n1510 & n1693 ;
  assign n1723 = n1722 ^ n1721 ;
  assign n1725 = n1541 & ~n1693 ;
  assign n1724 = n1528 & n1693 ;
  assign n1726 = n1725 ^ n1724 ;
  assign n1728 = n1558 & ~n1693 ;
  assign n1727 = n1545 & n1693 ;
  assign n1729 = n1728 ^ n1727 ;
  assign n1731 = n1577 & ~n1693 ;
  assign n1730 = n1564 & n1693 ;
  assign n1732 = n1731 ^ n1730 ;
  assign n1734 = n1594 & ~n1693 ;
  assign n1733 = n1581 & n1693 ;
  assign n1735 = n1734 ^ n1733 ;
  assign n1737 = n1609 & ~n1693 ;
  assign n1736 = n1612 & n1693 ;
  assign n1738 = n1737 ^ n1736 ;
  assign n1740 = n1626 & ~n1693 ;
  assign n1739 = n1629 & n1693 ;
  assign n1741 = n1740 ^ n1739 ;
  assign n2141 = n1381 & n1407 ;
  assign n2142 = n2141 ^ n1566 ;
  assign n2143 = n2142 ^ n1569 ;
  assign n2138 = ~n1381 & n1388 ;
  assign n2139 = n2138 ^ n1572 ;
  assign n2140 = n2139 ^ n1575 ;
  assign n2144 = n2143 ^ n2140 ;
  assign n1979 = n907 & n950 ;
  assign n1980 = n1979 ^ n1390 ;
  assign n1981 = n1980 ^ n1393 ;
  assign n1982 = n1981 ^ n1396 ;
  assign n1975 = ~n907 & n931 ;
  assign n1976 = n1975 ^ n1399 ;
  assign n1977 = n1976 ^ n1402 ;
  assign n1978 = n1977 ^ n1405 ;
  assign n1983 = n1982 ^ n1978 ;
  assign n1806 = n280 & n323 ;
  assign n1807 = n1806 ^ n933 ;
  assign n1808 = n1807 ^ n936 ;
  assign n1809 = n1808 ^ n939 ;
  assign n1802 = ~n280 & n304 ;
  assign n1803 = n1802 ^ n942 ;
  assign n1804 = n1803 ^ n945 ;
  assign n1805 = n1804 ^ n948 ;
  assign n1810 = n1809 ^ n1805 ;
  assign n1743 = n105 & n108 ;
  assign n1744 = n1743 ^ n114 ;
  assign n1742 = n119 & n139 ;
  assign n1745 = n1744 ^ n1742 ;
  assign n1746 = n1745 ^ n127 ;
  assign n1748 = x40 & ~n1746 ;
  assign n1747 = x32 & n1746 ;
  assign n1749 = n1748 ^ n1747 ;
  assign n1754 = n214 & n280 ;
  assign n1755 = n1754 ^ n824 ;
  assign n1756 = n1755 ^ n827 ;
  assign n1757 = n1756 ^ n830 ;
  assign n1750 = n233 & ~n280 ;
  assign n1751 = n1750 ^ n833 ;
  assign n1752 = n1751 ^ n836 ;
  assign n1753 = n1752 ^ n839 ;
  assign n1758 = n1757 ^ n1753 ;
  assign n1904 = ~n1749 & n1758 ;
  assign n1759 = n1758 ^ n1749 ;
  assign n1764 = n272 & n280 ;
  assign n1765 = n1764 ^ n863 ;
  assign n1766 = n1765 ^ n866 ;
  assign n1767 = n1766 ^ n869 ;
  assign n1760 = n253 & ~n280 ;
  assign n1761 = n1760 ^ n872 ;
  assign n1762 = n1761 ^ n875 ;
  assign n1763 = n1762 ^ n878 ;
  assign n1768 = n1767 ^ n1763 ;
  assign n1770 = x41 & ~n1746 ;
  assign n1769 = x33 & n1746 ;
  assign n1771 = n1770 ^ n1769 ;
  assign n1902 = n1768 & ~n1771 ;
  assign n1903 = ~n1759 & n1902 ;
  assign n1905 = n1904 ^ n1903 ;
  assign n1772 = n1771 ^ n1768 ;
  assign n1773 = ~n1759 & ~n1772 ;
  assign n1778 = n152 & n280 ;
  assign n1779 = n1778 ^ n276 ;
  assign n1780 = n1779 ^ n446 ;
  assign n1781 = n1780 ^ n459 ;
  assign n1774 = n100 & ~n280 ;
  assign n1775 = n1774 ^ n462 ;
  assign n1776 = n1775 ^ n465 ;
  assign n1777 = n1776 ^ n468 ;
  assign n1782 = n1781 ^ n1777 ;
  assign n1784 = x42 & ~n1746 ;
  assign n1783 = x34 & n1746 ;
  assign n1785 = n1784 ^ n1783 ;
  assign n1899 = n1782 & ~n1785 ;
  assign n1786 = n1785 ^ n1782 ;
  assign n1791 = n172 & n280 ;
  assign n1792 = n1791 ^ n782 ;
  assign n1793 = n1792 ^ n785 ;
  assign n1794 = n1793 ^ n788 ;
  assign n1787 = n191 & ~n280 ;
  assign n1788 = n1787 ^ n791 ;
  assign n1789 = n1788 ^ n794 ;
  assign n1790 = n1789 ^ n797 ;
  assign n1795 = n1794 ^ n1790 ;
  assign n1797 = x43 & ~n1746 ;
  assign n1796 = x35 & n1746 ;
  assign n1798 = n1797 ^ n1796 ;
  assign n1897 = n1795 & ~n1798 ;
  assign n1898 = ~n1786 & n1897 ;
  assign n1900 = n1899 ^ n1898 ;
  assign n1901 = n1773 & n1900 ;
  assign n1906 = n1905 ^ n1901 ;
  assign n1799 = n1798 ^ n1795 ;
  assign n1800 = ~n1786 & ~n1799 ;
  assign n1801 = n1773 & n1800 ;
  assign n1812 = x44 & ~n1746 ;
  assign n1811 = x36 & n1746 ;
  assign n1813 = n1812 ^ n1811 ;
  assign n1893 = n1810 & ~n1813 ;
  assign n1814 = n1813 ^ n1810 ;
  assign n1819 = n280 & n362 ;
  assign n1820 = n1819 ^ n972 ;
  assign n1821 = n1820 ^ n975 ;
  assign n1822 = n1821 ^ n978 ;
  assign n1815 = ~n280 & n343 ;
  assign n1816 = n1815 ^ n981 ;
  assign n1817 = n1816 ^ n984 ;
  assign n1818 = n1817 ^ n987 ;
  assign n1823 = n1822 ^ n1818 ;
  assign n1825 = x45 & ~n1746 ;
  assign n1824 = x37 & n1746 ;
  assign n1826 = n1825 ^ n1824 ;
  assign n1891 = n1823 & ~n1826 ;
  assign n1892 = ~n1814 & n1891 ;
  assign n1894 = n1893 ^ n1892 ;
  assign n1827 = n1826 ^ n1823 ;
  assign n1828 = ~n1814 & ~n1827 ;
  assign n1833 = n280 & n402 ;
  assign n1834 = n1833 ^ n1012 ;
  assign n1835 = n1834 ^ n1015 ;
  assign n1836 = n1835 ^ n1018 ;
  assign n1829 = ~n280 & n383 ;
  assign n1830 = n1829 ^ n1021 ;
  assign n1831 = n1830 ^ n1024 ;
  assign n1832 = n1831 ^ n1027 ;
  assign n1837 = n1836 ^ n1832 ;
  assign n1839 = x46 & ~n1746 ;
  assign n1838 = x38 & n1746 ;
  assign n1840 = n1839 ^ n1838 ;
  assign n1888 = n1837 & ~n1840 ;
  assign n1854 = x47 & n1744 ;
  assign n1855 = n1854 ^ n427 ;
  assign n1856 = n1855 ^ n430 ;
  assign n1851 = x39 & ~n1744 ;
  assign n1852 = n1851 ^ n436 ;
  assign n1853 = n1852 ^ n439 ;
  assign n1857 = n1856 ^ n1853 ;
  assign n1872 = n422 & ~n1857 ;
  assign n1879 = n285 & n1872 ;
  assign n1880 = n457 & n1879 ;
  assign n1877 = ~n445 & n1872 ;
  assign n1875 = ~n280 & n1872 ;
  assign n1873 = n274 & n1872 ;
  assign n1874 = n195 & n1873 ;
  assign n1876 = n1875 ^ n1874 ;
  assign n1878 = n1877 ^ n1876 ;
  assign n1881 = n1880 ^ n1878 ;
  assign n1862 = n441 & ~n1857 ;
  assign n1869 = n285 & n1862 ;
  assign n1870 = n457 & n1869 ;
  assign n1867 = ~n445 & n1862 ;
  assign n1865 = n280 & n1862 ;
  assign n1863 = n274 & n1862 ;
  assign n1864 = n195 & n1863 ;
  assign n1866 = n1865 ^ n1864 ;
  assign n1868 = n1867 ^ n1866 ;
  assign n1871 = n1870 ^ n1868 ;
  assign n1882 = n1881 ^ n1871 ;
  assign n1886 = ~n1840 & n1882 ;
  assign n1884 = n1836 & n1882 ;
  assign n1883 = n1832 & n1882 ;
  assign n1885 = n1884 ^ n1883 ;
  assign n1887 = n1886 ^ n1885 ;
  assign n1889 = n1888 ^ n1887 ;
  assign n1890 = n1828 & n1889 ;
  assign n1895 = n1894 ^ n1890 ;
  assign n1896 = n1801 & n1895 ;
  assign n1907 = n1906 ^ n1896 ;
  assign n1841 = n1840 ^ n1837 ;
  assign n1846 = n280 & n441 ;
  assign n1847 = n1846 ^ n1051 ;
  assign n1848 = n1847 ^ n1054 ;
  assign n1849 = n1848 ^ n1057 ;
  assign n1842 = ~n280 & n422 ;
  assign n1843 = n1842 ^ n1060 ;
  assign n1844 = n1843 ^ n1063 ;
  assign n1845 = n1844 ^ n1066 ;
  assign n1850 = n1849 ^ n1845 ;
  assign n1858 = n1857 ^ n1850 ;
  assign n1859 = ~n1841 & ~n1858 ;
  assign n1860 = n1828 & n1859 ;
  assign n1861 = n1801 & n1860 ;
  assign n1908 = n1907 ^ n1861 ;
  assign n1985 = n1810 & ~n1908 ;
  assign n1984 = n1813 & n1908 ;
  assign n1986 = n1985 ^ n1984 ;
  assign n2040 = n1983 & ~n1986 ;
  assign n1987 = n1986 ^ n1983 ;
  assign n1992 = n907 & n989 ;
  assign n1993 = n1992 ^ n1413 ;
  assign n1994 = n1993 ^ n1416 ;
  assign n1995 = n1994 ^ n1419 ;
  assign n1988 = ~n907 & n970 ;
  assign n1989 = n1988 ^ n1422 ;
  assign n1990 = n1989 ^ n1425 ;
  assign n1991 = n1990 ^ n1428 ;
  assign n1996 = n1995 ^ n1991 ;
  assign n1998 = n1823 & ~n1908 ;
  assign n1997 = n1826 & n1908 ;
  assign n1999 = n1998 ^ n1997 ;
  assign n2038 = n1996 & ~n1999 ;
  assign n2039 = ~n1987 & n2038 ;
  assign n2041 = n2040 ^ n2039 ;
  assign n2000 = n1999 ^ n1996 ;
  assign n2001 = ~n1987 & ~n2000 ;
  assign n2006 = n907 & n1029 ;
  assign n2007 = n2006 ^ n1437 ;
  assign n2008 = n2007 ^ n1440 ;
  assign n2009 = n2008 ^ n1443 ;
  assign n2002 = ~n907 & n1010 ;
  assign n2003 = n2002 ^ n1446 ;
  assign n2004 = n2003 ^ n1449 ;
  assign n2005 = n2004 ^ n1452 ;
  assign n2010 = n2009 ^ n2005 ;
  assign n2012 = n1837 & ~n1908 ;
  assign n2011 = n1840 & n1908 ;
  assign n2013 = n2012 ^ n2011 ;
  assign n2035 = n2010 & ~n2013 ;
  assign n2014 = n2013 ^ n2010 ;
  assign n2019 = n907 & n1068 ;
  assign n2020 = n2019 ^ n1460 ;
  assign n2021 = n2020 ^ n1463 ;
  assign n2022 = n2021 ^ n1466 ;
  assign n2015 = ~n907 & n1049 ;
  assign n2016 = n2015 ^ n1469 ;
  assign n2017 = n2016 ^ n1472 ;
  assign n2018 = n2017 ^ n1475 ;
  assign n2023 = n2022 ^ n2018 ;
  assign n2025 = n1850 & ~n1908 ;
  assign n2024 = n1857 & n1908 ;
  assign n2026 = n2025 ^ n2024 ;
  assign n2033 = n2023 & ~n2026 ;
  assign n2034 = ~n2014 & n2033 ;
  assign n2036 = n2035 ^ n2034 ;
  assign n2037 = n2001 & n2036 ;
  assign n2042 = n2041 ^ n2037 ;
  assign n1916 = n841 & n907 ;
  assign n1917 = n1916 ^ n903 ;
  assign n1918 = n1917 ^ n1073 ;
  assign n1919 = n1918 ^ n1086 ;
  assign n1912 = n860 & ~n907 ;
  assign n1913 = n1912 ^ n1089 ;
  assign n1914 = n1913 ^ n1092 ;
  assign n1915 = n1914 ^ n1095 ;
  assign n1920 = n1919 ^ n1915 ;
  assign n1910 = n1758 & ~n1908 ;
  assign n1909 = n1749 & n1908 ;
  assign n1911 = n1910 ^ n1909 ;
  assign n1921 = n1920 ^ n1911 ;
  assign n1932 = n1768 & ~n1908 ;
  assign n1931 = n1771 & n1908 ;
  assign n1933 = n1932 ^ n1931 ;
  assign n1926 = n880 & n907 ;
  assign n1927 = n1926 ^ n1307 ;
  assign n1928 = n1927 ^ n1310 ;
  assign n1929 = n1928 ^ n1313 ;
  assign n1922 = n899 & ~n907 ;
  assign n1923 = n1922 ^ n1316 ;
  assign n1924 = n1923 ^ n1319 ;
  assign n1925 = n1924 ^ n1322 ;
  assign n1930 = n1929 ^ n1925 ;
  assign n1934 = n1933 ^ n1930 ;
  assign n1935 = ~n1921 & ~n1934 ;
  assign n1946 = n1782 & ~n1908 ;
  assign n1945 = n1785 & n1908 ;
  assign n1947 = n1946 ^ n1945 ;
  assign n1940 = n470 & n907 ;
  assign n1941 = n1940 ^ n1331 ;
  assign n1942 = n1941 ^ n1334 ;
  assign n1943 = n1942 ^ n1337 ;
  assign n1936 = n779 & ~n907 ;
  assign n1937 = n1936 ^ n1340 ;
  assign n1938 = n1937 ^ n1343 ;
  assign n1939 = n1938 ^ n1346 ;
  assign n1944 = n1943 ^ n1939 ;
  assign n1948 = n1947 ^ n1944 ;
  assign n1956 = n799 & n907 ;
  assign n1957 = n1956 ^ n1351 ;
  assign n1958 = n1957 ^ n1354 ;
  assign n1959 = n1958 ^ n1357 ;
  assign n1952 = n818 & ~n907 ;
  assign n1953 = n1952 ^ n1360 ;
  assign n1954 = n1953 ^ n1363 ;
  assign n1955 = n1954 ^ n1366 ;
  assign n1960 = n1959 ^ n1955 ;
  assign n1950 = n1795 & ~n1908 ;
  assign n1949 = n1798 & n1908 ;
  assign n1951 = n1950 ^ n1949 ;
  assign n1972 = n1960 ^ n1951 ;
  assign n1973 = ~n1948 & ~n1972 ;
  assign n1974 = n1935 & n1973 ;
  assign n2154 = n1974 & n1983 ;
  assign n2155 = n2042 & n2154 ;
  assign n2027 = n2026 ^ n2023 ;
  assign n2028 = ~n2014 & ~n2027 ;
  assign n2029 = n2001 & n2028 ;
  assign n2030 = n1974 & n2029 ;
  assign n2152 = n1983 & ~n2030 ;
  assign n1968 = ~n1911 & n1920 ;
  assign n1966 = n1930 & ~n1933 ;
  assign n1967 = ~n1921 & n1966 ;
  assign n1969 = n1968 ^ n1967 ;
  assign n1963 = n1944 & ~n1947 ;
  assign n1961 = ~n1951 & n1960 ;
  assign n1962 = ~n1948 & n1961 ;
  assign n1964 = n1963 ^ n1962 ;
  assign n1965 = n1935 & n1964 ;
  assign n1970 = n1969 ^ n1965 ;
  assign n2151 = n1970 & n1983 ;
  assign n2153 = n2152 ^ n2151 ;
  assign n2156 = n2155 ^ n2153 ;
  assign n2148 = n1974 & n1986 ;
  assign n2149 = n2042 & n2148 ;
  assign n2146 = n1986 & ~n2030 ;
  assign n2145 = ~n1970 & n1986 ;
  assign n2147 = n2146 ^ n2145 ;
  assign n2150 = n2149 ^ n2147 ;
  assign n2157 = n2156 ^ n2150 ;
  assign n2247 = n2144 & ~n2157 ;
  assign n2158 = n2157 ^ n2144 ;
  assign n2162 = n1381 & n1430 ;
  assign n2163 = n2162 ^ n1583 ;
  assign n2164 = n2163 ^ n1586 ;
  assign n2159 = ~n1381 & n1411 ;
  assign n2160 = n2159 ^ n1589 ;
  assign n2161 = n2160 ^ n1592 ;
  assign n2165 = n2164 ^ n2161 ;
  assign n2175 = n1974 & n1996 ;
  assign n2176 = n2042 & n2175 ;
  assign n2173 = n1996 & ~n2030 ;
  assign n2172 = n1970 & n1996 ;
  assign n2174 = n2173 ^ n2172 ;
  assign n2177 = n2176 ^ n2174 ;
  assign n2169 = n1974 & n1999 ;
  assign n2170 = n2042 & n2169 ;
  assign n2167 = n1999 & ~n2030 ;
  assign n2166 = ~n1970 & n1999 ;
  assign n2168 = n2167 ^ n2166 ;
  assign n2171 = n2170 ^ n2168 ;
  assign n2178 = n2177 ^ n2171 ;
  assign n2245 = n2165 & ~n2178 ;
  assign n2246 = ~n2158 & n2245 ;
  assign n2248 = n2247 ^ n2246 ;
  assign n2179 = n2178 ^ n2165 ;
  assign n2180 = ~n2158 & ~n2179 ;
  assign n2184 = n1381 & n1454 ;
  assign n2185 = n2184 ^ n1598 ;
  assign n2186 = n2185 ^ n1601 ;
  assign n2181 = ~n1381 & n1435 ;
  assign n2182 = n2181 ^ n1604 ;
  assign n2183 = n2182 ^ n1607 ;
  assign n2187 = n2186 ^ n2183 ;
  assign n2197 = n1974 & n2010 ;
  assign n2198 = n2042 & n2197 ;
  assign n2195 = n2010 & ~n2030 ;
  assign n2194 = n1970 & n2010 ;
  assign n2196 = n2195 ^ n2194 ;
  assign n2199 = n2198 ^ n2196 ;
  assign n2191 = n1974 & n2013 ;
  assign n2192 = n2042 & n2191 ;
  assign n2189 = n2013 & ~n2030 ;
  assign n2188 = ~n1970 & n2013 ;
  assign n2190 = n2189 ^ n2188 ;
  assign n2193 = n2192 ^ n2190 ;
  assign n2200 = n2199 ^ n2193 ;
  assign n2242 = n2187 & ~n2200 ;
  assign n2201 = n2200 ^ n2187 ;
  assign n2210 = n1380 & n1477 ;
  assign n2208 = n1326 & n1477 ;
  assign n2209 = n1375 & n2208 ;
  assign n2211 = n2210 ^ n2209 ;
  assign n2212 = n2211 ^ n1615 ;
  assign n2213 = n2212 ^ n1618 ;
  assign n2204 = ~n1380 & n1458 ;
  assign n2202 = n1326 & n1458 ;
  assign n2203 = n1375 & n2202 ;
  assign n2205 = n2204 ^ n2203 ;
  assign n2206 = n2205 ^ n1621 ;
  assign n2207 = n2206 ^ n1624 ;
  assign n2214 = n2213 ^ n2207 ;
  assign n2230 = n1974 & n2023 ;
  assign n2231 = n2042 & n2230 ;
  assign n2228 = n2023 & ~n2030 ;
  assign n2226 = n1969 & n2023 ;
  assign n2224 = n1935 & n2023 ;
  assign n2225 = n1964 & n2224 ;
  assign n2227 = n2226 ^ n2225 ;
  assign n2229 = n2228 ^ n2227 ;
  assign n2232 = n2231 ^ n2229 ;
  assign n2221 = n1974 & n2026 ;
  assign n2222 = n2042 & n2221 ;
  assign n2219 = n2026 & ~n2030 ;
  assign n2217 = ~n1969 & n2026 ;
  assign n2215 = n1935 & n2026 ;
  assign n2216 = n1964 & n2215 ;
  assign n2218 = n2217 ^ n2216 ;
  assign n2220 = n2219 ^ n2218 ;
  assign n2223 = n2222 ^ n2220 ;
  assign n2233 = n2232 ^ n2223 ;
  assign n2240 = n2214 & ~n2233 ;
  assign n2241 = ~n2201 & n2240 ;
  assign n2243 = n2242 ^ n2241 ;
  assign n2244 = n2180 & n2243 ;
  assign n2249 = n2248 ^ n2244 ;
  assign n2056 = n1097 & n1381 ;
  assign n2057 = n2056 ^ n1482 ;
  assign n2058 = n2057 ^ n1495 ;
  assign n2053 = n1301 & ~n1381 ;
  assign n2054 = n2053 ^ n1498 ;
  assign n2055 = n2054 ^ n1501 ;
  assign n2059 = n2058 ^ n2055 ;
  assign n2049 = n1920 & n1974 ;
  assign n2050 = n2042 & n2049 ;
  assign n2047 = n1920 & ~n2030 ;
  assign n2046 = n1920 & n1970 ;
  assign n2048 = n2047 ^ n2046 ;
  assign n2051 = n2050 ^ n2048 ;
  assign n2043 = n1911 & n1974 ;
  assign n2044 = n2042 & n2043 ;
  assign n2031 = n1911 & ~n2030 ;
  assign n1971 = n1911 & ~n1970 ;
  assign n2032 = n2031 ^ n1971 ;
  assign n2045 = n2044 ^ n2032 ;
  assign n2052 = n2051 ^ n2045 ;
  assign n2060 = n2059 ^ n2052 ;
  assign n2077 = n1930 & n1974 ;
  assign n2078 = n2042 & n2077 ;
  assign n2075 = n1930 & ~n2030 ;
  assign n2074 = n1930 & n1970 ;
  assign n2076 = n2075 ^ n2074 ;
  assign n2079 = n2078 ^ n2076 ;
  assign n2071 = n1933 & n1974 ;
  assign n2072 = n2042 & n2071 ;
  assign n2069 = n1933 & ~n2030 ;
  assign n2068 = n1933 & ~n1970 ;
  assign n2070 = n2069 ^ n2068 ;
  assign n2073 = n2072 ^ n2070 ;
  assign n2080 = n2079 ^ n2073 ;
  assign n2064 = n1324 & n1381 ;
  assign n2065 = n2064 ^ n1512 ;
  assign n2066 = n2065 ^ n1515 ;
  assign n2061 = n1305 & ~n1381 ;
  assign n2062 = n2061 ^ n1518 ;
  assign n2063 = n2062 ^ n1521 ;
  assign n2067 = n2066 ^ n2063 ;
  assign n2081 = n2080 ^ n2067 ;
  assign n2082 = ~n2060 & ~n2081 ;
  assign n2099 = n1944 & n1974 ;
  assign n2100 = n2042 & n2099 ;
  assign n2097 = n1944 & ~n2030 ;
  assign n2096 = n1944 & n1970 ;
  assign n2098 = n2097 ^ n2096 ;
  assign n2101 = n2100 ^ n2098 ;
  assign n2093 = n1947 & n1974 ;
  assign n2094 = n2042 & n2093 ;
  assign n2091 = n1947 & ~n2030 ;
  assign n2090 = n1947 & ~n1970 ;
  assign n2092 = n2091 ^ n2090 ;
  assign n2095 = n2094 ^ n2092 ;
  assign n2102 = n2101 ^ n2095 ;
  assign n2086 = n1348 & n1381 ;
  assign n2087 = n2086 ^ n1530 ;
  assign n2088 = n2087 ^ n1533 ;
  assign n2083 = n1329 & ~n1381 ;
  assign n2084 = n2083 ^ n1536 ;
  assign n2085 = n2084 ^ n1539 ;
  assign n2089 = n2088 ^ n2085 ;
  assign n2103 = n2102 ^ n2089 ;
  assign n2120 = n1368 & n1381 ;
  assign n2121 = n2120 ^ n1547 ;
  assign n2122 = n2121 ^ n1550 ;
  assign n2117 = n1371 & ~n1381 ;
  assign n2118 = n2117 ^ n1553 ;
  assign n2119 = n2118 ^ n1556 ;
  assign n2123 = n2122 ^ n2119 ;
  assign n2113 = n1960 & n1974 ;
  assign n2114 = n2042 & n2113 ;
  assign n2111 = n1960 & ~n2030 ;
  assign n2110 = n1960 & n1970 ;
  assign n2112 = n2111 ^ n2110 ;
  assign n2115 = n2114 ^ n2112 ;
  assign n2107 = n1951 & n1974 ;
  assign n2108 = n2042 & n2107 ;
  assign n2105 = n1951 & ~n2030 ;
  assign n2104 = n1951 & ~n1970 ;
  assign n2106 = n2105 ^ n2104 ;
  assign n2109 = n2108 ^ n2106 ;
  assign n2116 = n2115 ^ n2109 ;
  assign n2135 = n2123 ^ n2116 ;
  assign n2136 = ~n2103 & ~n2135 ;
  assign n2137 = n2082 & n2136 ;
  assign n2256 = n2059 & n2137 ;
  assign n2257 = n2249 & n2256 ;
  assign n2234 = n2233 ^ n2214 ;
  assign n2235 = ~n2201 & ~n2234 ;
  assign n2236 = n2180 & n2235 ;
  assign n2237 = n2137 & n2236 ;
  assign n2254 = n2059 & ~n2237 ;
  assign n2131 = ~n2052 & n2059 ;
  assign n2129 = n2067 & ~n2080 ;
  assign n2130 = ~n2060 & n2129 ;
  assign n2132 = n2131 ^ n2130 ;
  assign n2126 = n2089 & ~n2102 ;
  assign n2124 = ~n2116 & n2123 ;
  assign n2125 = ~n2103 & n2124 ;
  assign n2127 = n2126 ^ n2125 ;
  assign n2128 = n2082 & n2127 ;
  assign n2133 = n2132 ^ n2128 ;
  assign n2253 = n2059 & n2133 ;
  assign n2255 = n2254 ^ n2253 ;
  assign n2258 = n2257 ^ n2255 ;
  assign n2250 = n2052 & n2137 ;
  assign n2251 = n2249 & n2250 ;
  assign n2238 = n2052 & ~n2237 ;
  assign n2134 = n2052 & ~n2133 ;
  assign n2239 = n2238 ^ n2134 ;
  assign n2252 = n2251 ^ n2239 ;
  assign n2259 = n2258 ^ n2252 ;
  assign n2269 = n2067 & n2137 ;
  assign n2270 = n2249 & n2269 ;
  assign n2267 = n2067 & ~n2237 ;
  assign n2266 = n2067 & n2133 ;
  assign n2268 = n2267 ^ n2266 ;
  assign n2271 = n2270 ^ n2268 ;
  assign n2263 = n2080 & n2137 ;
  assign n2264 = n2249 & n2263 ;
  assign n2261 = n2080 & ~n2237 ;
  assign n2260 = n2080 & ~n2133 ;
  assign n2262 = n2261 ^ n2260 ;
  assign n2265 = n2264 ^ n2262 ;
  assign n2272 = n2271 ^ n2265 ;
  assign n2282 = n2089 & n2137 ;
  assign n2283 = n2249 & n2282 ;
  assign n2280 = n2089 & ~n2237 ;
  assign n2279 = n2089 & n2133 ;
  assign n2281 = n2280 ^ n2279 ;
  assign n2284 = n2283 ^ n2281 ;
  assign n2276 = n2102 & n2137 ;
  assign n2277 = n2249 & n2276 ;
  assign n2274 = n2102 & ~n2237 ;
  assign n2273 = n2102 & ~n2133 ;
  assign n2275 = n2274 ^ n2273 ;
  assign n2278 = n2277 ^ n2275 ;
  assign n2285 = n2284 ^ n2278 ;
  assign n2295 = n2123 & n2137 ;
  assign n2296 = n2249 & n2295 ;
  assign n2293 = n2123 & ~n2237 ;
  assign n2292 = n2123 & n2133 ;
  assign n2294 = n2293 ^ n2292 ;
  assign n2297 = n2296 ^ n2294 ;
  assign n2289 = n2116 & n2137 ;
  assign n2290 = n2249 & n2289 ;
  assign n2287 = n2116 & ~n2237 ;
  assign n2286 = n2116 & ~n2133 ;
  assign n2288 = n2287 ^ n2286 ;
  assign n2291 = n2290 ^ n2288 ;
  assign n2298 = n2297 ^ n2291 ;
  assign n2308 = n2137 & n2144 ;
  assign n2309 = n2249 & n2308 ;
  assign n2306 = n2144 & ~n2237 ;
  assign n2305 = n2133 & n2144 ;
  assign n2307 = n2306 ^ n2305 ;
  assign n2310 = n2309 ^ n2307 ;
  assign n2302 = n2137 & n2157 ;
  assign n2303 = n2249 & n2302 ;
  assign n2300 = n2157 & ~n2237 ;
  assign n2299 = ~n2133 & n2157 ;
  assign n2301 = n2300 ^ n2299 ;
  assign n2304 = n2303 ^ n2301 ;
  assign n2311 = n2310 ^ n2304 ;
  assign n2321 = n2137 & n2165 ;
  assign n2322 = n2249 & n2321 ;
  assign n2319 = n2165 & ~n2237 ;
  assign n2318 = n2133 & n2165 ;
  assign n2320 = n2319 ^ n2318 ;
  assign n2323 = n2322 ^ n2320 ;
  assign n2315 = n2137 & n2178 ;
  assign n2316 = n2249 & n2315 ;
  assign n2313 = n2178 & ~n2237 ;
  assign n2312 = ~n2133 & n2178 ;
  assign n2314 = n2313 ^ n2312 ;
  assign n2317 = n2316 ^ n2314 ;
  assign n2324 = n2323 ^ n2317 ;
  assign n2334 = n2137 & n2187 ;
  assign n2335 = n2249 & n2334 ;
  assign n2332 = n2187 & ~n2237 ;
  assign n2331 = n2133 & n2187 ;
  assign n2333 = n2332 ^ n2331 ;
  assign n2336 = n2335 ^ n2333 ;
  assign n2328 = n2137 & n2200 ;
  assign n2329 = n2249 & n2328 ;
  assign n2326 = n2200 & ~n2237 ;
  assign n2325 = ~n2133 & n2200 ;
  assign n2327 = n2326 ^ n2325 ;
  assign n2330 = n2329 ^ n2327 ;
  assign n2337 = n2336 ^ n2330 ;
  assign n2347 = n2137 & n2214 ;
  assign n2348 = n2249 & n2347 ;
  assign n2345 = n2214 & ~n2237 ;
  assign n2344 = n2133 & n2214 ;
  assign n2346 = n2345 ^ n2344 ;
  assign n2349 = n2348 ^ n2346 ;
  assign n2341 = n2137 & n2233 ;
  assign n2342 = n2249 & n2341 ;
  assign n2339 = n2233 & ~n2237 ;
  assign n2338 = ~n2133 & n2233 ;
  assign n2340 = n2339 ^ n2338 ;
  assign n2343 = n2342 ^ n2340 ;
  assign n2350 = n2349 ^ n2343 ;
  assign n2354 = n2052 & n2133 ;
  assign n2355 = n2354 ^ n2238 ;
  assign n2356 = n2355 ^ n2251 ;
  assign n2351 = n2059 & ~n2133 ;
  assign n2352 = n2351 ^ n2254 ;
  assign n2353 = n2352 ^ n2257 ;
  assign n2357 = n2356 ^ n2353 ;
  assign n2361 = n2080 & n2133 ;
  assign n2362 = n2361 ^ n2261 ;
  assign n2363 = n2362 ^ n2264 ;
  assign n2358 = n2067 & ~n2133 ;
  assign n2359 = n2358 ^ n2267 ;
  assign n2360 = n2359 ^ n2270 ;
  assign n2364 = n2363 ^ n2360 ;
  assign n2368 = n2102 & n2133 ;
  assign n2369 = n2368 ^ n2274 ;
  assign n2370 = n2369 ^ n2277 ;
  assign n2365 = n2089 & ~n2133 ;
  assign n2366 = n2365 ^ n2280 ;
  assign n2367 = n2366 ^ n2283 ;
  assign n2371 = n2370 ^ n2367 ;
  assign n2375 = n2116 & n2133 ;
  assign n2376 = n2375 ^ n2287 ;
  assign n2377 = n2376 ^ n2290 ;
  assign n2372 = n2123 & ~n2133 ;
  assign n2373 = n2372 ^ n2293 ;
  assign n2374 = n2373 ^ n2296 ;
  assign n2378 = n2377 ^ n2374 ;
  assign n2382 = n2133 & n2157 ;
  assign n2383 = n2382 ^ n2300 ;
  assign n2384 = n2383 ^ n2303 ;
  assign n2379 = ~n2133 & n2144 ;
  assign n2380 = n2379 ^ n2306 ;
  assign n2381 = n2380 ^ n2309 ;
  assign n2385 = n2384 ^ n2381 ;
  assign n2389 = n2133 & n2178 ;
  assign n2390 = n2389 ^ n2313 ;
  assign n2391 = n2390 ^ n2316 ;
  assign n2386 = ~n2133 & n2165 ;
  assign n2387 = n2386 ^ n2319 ;
  assign n2388 = n2387 ^ n2322 ;
  assign n2392 = n2391 ^ n2388 ;
  assign n2396 = n2133 & n2200 ;
  assign n2397 = n2396 ^ n2326 ;
  assign n2398 = n2397 ^ n2329 ;
  assign n2393 = ~n2133 & n2187 ;
  assign n2394 = n2393 ^ n2332 ;
  assign n2395 = n2394 ^ n2335 ;
  assign n2399 = n2398 ^ n2395 ;
  assign n2403 = n2133 & n2233 ;
  assign n2404 = n2403 ^ n2339 ;
  assign n2405 = n2404 ^ n2342 ;
  assign n2400 = ~n2133 & n2214 ;
  assign n2401 = n2400 ^ n2345 ;
  assign n2402 = n2401 ^ n2348 ;
  assign n2406 = n2405 ^ n2402 ;
  assign n2413 = n1911 & n1970 ;
  assign n2414 = n2413 ^ n2031 ;
  assign n2415 = n2414 ^ n2044 ;
  assign n2410 = n1920 & ~n1970 ;
  assign n2411 = n2410 ^ n2047 ;
  assign n2412 = n2411 ^ n2050 ;
  assign n2416 = n2415 ^ n2412 ;
  assign n2408 = n1749 & ~n1908 ;
  assign n2407 = n1758 & n1908 ;
  assign n2409 = n2408 ^ n2407 ;
  assign n2538 = ~n2409 & n2416 ;
  assign n2417 = n2416 ^ n2409 ;
  assign n2421 = n1933 & n1970 ;
  assign n2422 = n2421 ^ n2069 ;
  assign n2423 = n2422 ^ n2072 ;
  assign n2418 = n1930 & ~n1970 ;
  assign n2419 = n2418 ^ n2075 ;
  assign n2420 = n2419 ^ n2078 ;
  assign n2424 = n2423 ^ n2420 ;
  assign n2426 = n1771 & ~n1908 ;
  assign n2425 = n1768 & n1908 ;
  assign n2427 = n2426 ^ n2425 ;
  assign n2536 = n2424 & ~n2427 ;
  assign n2537 = ~n2417 & n2536 ;
  assign n2539 = n2538 ^ n2537 ;
  assign n2428 = n2427 ^ n2424 ;
  assign n2429 = ~n2417 & ~n2428 ;
  assign n2433 = n1947 & n1970 ;
  assign n2434 = n2433 ^ n2091 ;
  assign n2435 = n2434 ^ n2094 ;
  assign n2430 = n1944 & ~n1970 ;
  assign n2431 = n2430 ^ n2097 ;
  assign n2432 = n2431 ^ n2100 ;
  assign n2436 = n2435 ^ n2432 ;
  assign n2438 = n1785 & ~n1908 ;
  assign n2437 = n1782 & n1908 ;
  assign n2439 = n2438 ^ n2437 ;
  assign n2533 = n2436 & ~n2439 ;
  assign n2440 = n2439 ^ n2436 ;
  assign n2444 = n1951 & n1970 ;
  assign n2445 = n2444 ^ n2105 ;
  assign n2446 = n2445 ^ n2108 ;
  assign n2441 = n1960 & ~n1970 ;
  assign n2442 = n2441 ^ n2111 ;
  assign n2443 = n2442 ^ n2114 ;
  assign n2447 = n2446 ^ n2443 ;
  assign n2449 = n1798 & ~n1908 ;
  assign n2448 = n1795 & n1908 ;
  assign n2450 = n2449 ^ n2448 ;
  assign n2531 = n2447 & ~n2450 ;
  assign n2532 = ~n2440 & n2531 ;
  assign n2534 = n2533 ^ n2532 ;
  assign n2535 = n2429 & n2534 ;
  assign n2540 = n2539 ^ n2535 ;
  assign n2451 = n2450 ^ n2447 ;
  assign n2452 = ~n2440 & ~n2451 ;
  assign n2453 = n2429 & n2452 ;
  assign n2457 = n1970 & n1986 ;
  assign n2458 = n2457 ^ n2146 ;
  assign n2459 = n2458 ^ n2149 ;
  assign n2454 = ~n1970 & n1983 ;
  assign n2455 = n2454 ^ n2152 ;
  assign n2456 = n2455 ^ n2155 ;
  assign n2460 = n2459 ^ n2456 ;
  assign n2462 = n1813 & ~n1908 ;
  assign n2461 = n1810 & n1908 ;
  assign n2463 = n2462 ^ n2461 ;
  assign n2527 = n2460 & ~n2463 ;
  assign n2464 = n2463 ^ n2460 ;
  assign n2468 = n1970 & n1999 ;
  assign n2469 = n2468 ^ n2167 ;
  assign n2470 = n2469 ^ n2170 ;
  assign n2465 = ~n1970 & n1996 ;
  assign n2466 = n2465 ^ n2173 ;
  assign n2467 = n2466 ^ n2176 ;
  assign n2471 = n2470 ^ n2467 ;
  assign n2473 = n1826 & ~n1908 ;
  assign n2472 = n1823 & n1908 ;
  assign n2474 = n2473 ^ n2472 ;
  assign n2525 = n2471 & ~n2474 ;
  assign n2526 = ~n2464 & n2525 ;
  assign n2528 = n2527 ^ n2526 ;
  assign n2475 = n2474 ^ n2471 ;
  assign n2476 = ~n2464 & ~n2475 ;
  assign n2480 = n1970 & n2013 ;
  assign n2481 = n2480 ^ n2189 ;
  assign n2482 = n2481 ^ n2192 ;
  assign n2477 = ~n1970 & n2010 ;
  assign n2478 = n2477 ^ n2195 ;
  assign n2479 = n2478 ^ n2198 ;
  assign n2483 = n2482 ^ n2479 ;
  assign n2485 = n1840 & ~n1908 ;
  assign n2484 = n1837 & n1908 ;
  assign n2486 = n2485 ^ n2484 ;
  assign n2522 = n2483 & ~n2486 ;
  assign n2496 = n1857 & ~n1908 ;
  assign n2495 = n1850 & n1908 ;
  assign n2497 = n2496 ^ n2495 ;
  assign n2509 = n2023 & ~n2497 ;
  assign n2513 = n1974 & n2509 ;
  assign n2514 = n2042 & n2513 ;
  assign n2511 = ~n2030 & n2509 ;
  assign n2510 = ~n1970 & n2509 ;
  assign n2512 = n2511 ^ n2510 ;
  assign n2515 = n2514 ^ n2512 ;
  assign n2502 = n2026 & ~n2497 ;
  assign n2506 = n1974 & n2502 ;
  assign n2507 = n2042 & n2506 ;
  assign n2504 = ~n2030 & n2502 ;
  assign n2503 = n1970 & n2502 ;
  assign n2505 = n2504 ^ n2503 ;
  assign n2508 = n2507 ^ n2505 ;
  assign n2516 = n2515 ^ n2508 ;
  assign n2520 = ~n2486 & n2516 ;
  assign n2518 = n2482 & n2516 ;
  assign n2517 = n2479 & n2516 ;
  assign n2519 = n2518 ^ n2517 ;
  assign n2521 = n2520 ^ n2519 ;
  assign n2523 = n2522 ^ n2521 ;
  assign n2524 = n2476 & n2523 ;
  assign n2529 = n2528 ^ n2524 ;
  assign n2530 = n2453 & n2529 ;
  assign n2541 = n2540 ^ n2530 ;
  assign n2487 = n2486 ^ n2483 ;
  assign n2491 = n1970 & n2026 ;
  assign n2492 = n2491 ^ n2219 ;
  assign n2493 = n2492 ^ n2222 ;
  assign n2488 = ~n1970 & n2023 ;
  assign n2489 = n2488 ^ n2228 ;
  assign n2490 = n2489 ^ n2231 ;
  assign n2494 = n2493 ^ n2490 ;
  assign n2498 = n2497 ^ n2494 ;
  assign n2499 = ~n2487 & ~n2498 ;
  assign n2500 = n2476 & n2499 ;
  assign n2501 = n2453 & n2500 ;
  assign n2542 = n2541 ^ n2501 ;
  assign n2544 = n2416 & ~n2542 ;
  assign n2543 = n2409 & n2542 ;
  assign n2545 = n2544 ^ n2543 ;
  assign n2547 = n2424 & ~n2542 ;
  assign n2546 = n2427 & n2542 ;
  assign n2548 = n2547 ^ n2546 ;
  assign n2550 = n2436 & ~n2542 ;
  assign n2549 = n2439 & n2542 ;
  assign n2551 = n2550 ^ n2549 ;
  assign n2553 = n2447 & ~n2542 ;
  assign n2552 = n2450 & n2542 ;
  assign n2554 = n2553 ^ n2552 ;
  assign n2556 = n2460 & ~n2542 ;
  assign n2555 = n2463 & n2542 ;
  assign n2557 = n2556 ^ n2555 ;
  assign n2559 = n2471 & ~n2542 ;
  assign n2558 = n2474 & n2542 ;
  assign n2560 = n2559 ^ n2558 ;
  assign n2562 = n2483 & ~n2542 ;
  assign n2561 = n2486 & n2542 ;
  assign n2563 = n2562 ^ n2561 ;
  assign n2565 = n2494 & ~n2542 ;
  assign n2564 = n2497 & n2542 ;
  assign n2566 = n2565 ^ n2564 ;
  assign n2568 = n2409 & ~n2542 ;
  assign n2567 = n2416 & n2542 ;
  assign n2569 = n2568 ^ n2567 ;
  assign n2571 = n2427 & ~n2542 ;
  assign n2570 = n2424 & n2542 ;
  assign n2572 = n2571 ^ n2570 ;
  assign n2574 = n2439 & ~n2542 ;
  assign n2573 = n2436 & n2542 ;
  assign n2575 = n2574 ^ n2573 ;
  assign n2577 = n2450 & ~n2542 ;
  assign n2576 = n2447 & n2542 ;
  assign n2578 = n2577 ^ n2576 ;
  assign n2580 = n2463 & ~n2542 ;
  assign n2579 = n2460 & n2542 ;
  assign n2581 = n2580 ^ n2579 ;
  assign n2583 = n2474 & ~n2542 ;
  assign n2582 = n2471 & n2542 ;
  assign n2584 = n2583 ^ n2582 ;
  assign n2586 = n2486 & ~n2542 ;
  assign n2585 = n2483 & n2542 ;
  assign n2587 = n2586 ^ n2585 ;
  assign n2589 = n2497 & ~n2542 ;
  assign n2588 = n2494 & n2542 ;
  assign n2590 = n2589 ^ n2588 ;
  assign y0 = n1696 ;
  assign y1 = n1699 ;
  assign y2 = n1702 ;
  assign y3 = n1705 ;
  assign y4 = n1708 ;
  assign y5 = n1711 ;
  assign y6 = n1714 ;
  assign y7 = n1717 ;
  assign y8 = n1720 ;
  assign y9 = n1723 ;
  assign y10 = n1726 ;
  assign y11 = n1729 ;
  assign y12 = n1732 ;
  assign y13 = n1735 ;
  assign y14 = n1738 ;
  assign y15 = n1741 ;
  assign y16 = n2259 ;
  assign y17 = n2272 ;
  assign y18 = n2285 ;
  assign y19 = n2298 ;
  assign y20 = n2311 ;
  assign y21 = n2324 ;
  assign y22 = n2337 ;
  assign y23 = n2350 ;
  assign y24 = n2357 ;
  assign y25 = n2364 ;
  assign y26 = n2371 ;
  assign y27 = n2378 ;
  assign y28 = n2385 ;
  assign y29 = n2392 ;
  assign y30 = n2399 ;
  assign y31 = n2406 ;
  assign y32 = n2545 ;
  assign y33 = n2548 ;
  assign y34 = n2551 ;
  assign y35 = n2554 ;
  assign y36 = n2557 ;
  assign y37 = n2560 ;
  assign y38 = n2563 ;
  assign y39 = n2566 ;
  assign y40 = n2569 ;
  assign y41 = n2572 ;
  assign y42 = n2575 ;
  assign y43 = n2578 ;
  assign y44 = n2581 ;
  assign y45 = n2584 ;
  assign y46 = n2587 ;
  assign y47 = n2590 ;
endmodule
