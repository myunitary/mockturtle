module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 ;
  assign n257 = ~x159 & ~x191 ;
  assign n258 = ~x223 & ~x255 ;
  assign n259 = n257 & n258 ;
  assign n260 = ~x31 & ~x63 ;
  assign n261 = ~x95 & ~x127 ;
  assign n262 = n260 & n261 ;
  assign n263 = n259 & ~n262 ;
  assign n264 = ~x31 & x63 ;
  assign n265 = x31 & ~x63 ;
  assign n266 = ~x30 & x62 ;
  assign n267 = x30 & ~x62 ;
  assign n268 = ~x29 & x61 ;
  assign n269 = x29 & ~x61 ;
  assign n270 = ~x28 & x60 ;
  assign n271 = x28 & ~x60 ;
  assign n272 = ~x27 & x59 ;
  assign n273 = x27 & ~x59 ;
  assign n274 = ~x26 & x58 ;
  assign n275 = x26 & ~x58 ;
  assign n276 = ~x25 & x57 ;
  assign n277 = x25 & ~x57 ;
  assign n278 = ~x24 & x56 ;
  assign n279 = x24 & ~x56 ;
  assign n280 = ~x23 & x55 ;
  assign n281 = x23 & ~x55 ;
  assign n282 = ~x22 & x54 ;
  assign n283 = x22 & ~x54 ;
  assign n284 = ~x21 & x53 ;
  assign n285 = x21 & ~x53 ;
  assign n286 = ~x20 & x52 ;
  assign n287 = x20 & ~x52 ;
  assign n288 = ~x19 & x51 ;
  assign n289 = x19 & ~x51 ;
  assign n290 = ~x18 & x50 ;
  assign n291 = x18 & ~x50 ;
  assign n292 = ~x17 & x49 ;
  assign n293 = x17 & ~x49 ;
  assign n294 = ~x16 & x48 ;
  assign n295 = x16 & ~x48 ;
  assign n296 = ~x15 & x47 ;
  assign n297 = x15 & ~x47 ;
  assign n298 = ~x14 & x46 ;
  assign n299 = x14 & ~x46 ;
  assign n300 = ~x13 & x45 ;
  assign n301 = x13 & ~x45 ;
  assign n302 = ~x12 & x44 ;
  assign n303 = x12 & ~x44 ;
  assign n304 = ~x11 & x43 ;
  assign n305 = x11 & ~x43 ;
  assign n306 = ~x10 & x42 ;
  assign n307 = x10 & ~x42 ;
  assign n308 = ~x9 & x41 ;
  assign n309 = x9 & ~x41 ;
  assign n310 = ~x8 & x40 ;
  assign n311 = x8 & ~x40 ;
  assign n312 = ~x7 & x39 ;
  assign n313 = x7 & ~x39 ;
  assign n314 = ~x6 & x38 ;
  assign n315 = x6 & ~x38 ;
  assign n316 = ~x5 & x37 ;
  assign n317 = x5 & ~x37 ;
  assign n318 = ~x4 & x36 ;
  assign n319 = x4 & ~x36 ;
  assign n320 = ~x3 & x35 ;
  assign n321 = x3 & ~x35 ;
  assign n322 = ~x2 & x34 ;
  assign n323 = x2 & ~x34 ;
  assign n324 = ~x1 & x33 ;
  assign n325 = x1 & ~x33 ;
  assign n326 = x0 & ~x32 ;
  assign n327 = ~n325 & ~n326 ;
  assign n328 = ~n324 & ~n327 ;
  assign n329 = ~n323 & ~n328 ;
  assign n330 = ~n322 & ~n329 ;
  assign n331 = ~n321 & ~n330 ;
  assign n332 = ~n320 & ~n331 ;
  assign n333 = ~n319 & ~n332 ;
  assign n334 = ~n318 & ~n333 ;
  assign n335 = ~n317 & ~n334 ;
  assign n336 = ~n316 & ~n335 ;
  assign n337 = ~n315 & ~n336 ;
  assign n338 = ~n314 & ~n337 ;
  assign n339 = ~n313 & ~n338 ;
  assign n340 = ~n312 & ~n339 ;
  assign n341 = ~n311 & ~n340 ;
  assign n342 = ~n310 & ~n341 ;
  assign n343 = ~n309 & ~n342 ;
  assign n344 = ~n308 & ~n343 ;
  assign n345 = ~n307 & ~n344 ;
  assign n346 = ~n306 & ~n345 ;
  assign n347 = ~n305 & ~n346 ;
  assign n348 = ~n304 & ~n347 ;
  assign n349 = ~n303 & ~n348 ;
  assign n350 = ~n302 & ~n349 ;
  assign n351 = ~n301 & ~n350 ;
  assign n352 = ~n300 & ~n351 ;
  assign n353 = ~n299 & ~n352 ;
  assign n354 = ~n298 & ~n353 ;
  assign n355 = ~n297 & ~n354 ;
  assign n356 = ~n296 & ~n355 ;
  assign n357 = ~n295 & ~n356 ;
  assign n358 = ~n294 & ~n357 ;
  assign n359 = ~n293 & ~n358 ;
  assign n360 = ~n292 & ~n359 ;
  assign n361 = ~n291 & ~n360 ;
  assign n362 = ~n290 & ~n361 ;
  assign n363 = ~n289 & ~n362 ;
  assign n364 = ~n288 & ~n363 ;
  assign n365 = ~n287 & ~n364 ;
  assign n366 = ~n286 & ~n365 ;
  assign n367 = ~n285 & ~n366 ;
  assign n368 = ~n284 & ~n367 ;
  assign n369 = ~n283 & ~n368 ;
  assign n370 = ~n282 & ~n369 ;
  assign n371 = ~n281 & ~n370 ;
  assign n372 = ~n280 & ~n371 ;
  assign n373 = ~n279 & ~n372 ;
  assign n374 = ~n278 & ~n373 ;
  assign n375 = ~n277 & ~n374 ;
  assign n376 = ~n276 & ~n375 ;
  assign n377 = ~n275 & ~n376 ;
  assign n378 = ~n274 & ~n377 ;
  assign n379 = ~n273 & ~n378 ;
  assign n380 = ~n272 & ~n379 ;
  assign n381 = ~n271 & ~n380 ;
  assign n382 = ~n270 & ~n381 ;
  assign n383 = ~n269 & ~n382 ;
  assign n384 = ~n268 & ~n383 ;
  assign n385 = ~n267 & ~n384 ;
  assign n386 = ~n266 & ~n385 ;
  assign n387 = ~n265 & ~n386 ;
  assign n388 = ~n264 & ~n387 ;
  assign n389 = x33 & ~n388 ;
  assign n390 = x1 & n388 ;
  assign n391 = ~n389 & ~n390 ;
  assign n392 = n260 & ~n261 ;
  assign n393 = ~n260 & n261 ;
  assign n394 = ~x95 & x127 ;
  assign n395 = x95 & ~x127 ;
  assign n396 = ~x94 & x126 ;
  assign n397 = x94 & ~x126 ;
  assign n398 = ~x93 & x125 ;
  assign n399 = x93 & ~x125 ;
  assign n400 = ~x92 & x124 ;
  assign n401 = x92 & ~x124 ;
  assign n402 = ~x91 & x123 ;
  assign n403 = x91 & ~x123 ;
  assign n404 = ~x90 & x122 ;
  assign n405 = x90 & ~x122 ;
  assign n406 = ~x89 & x121 ;
  assign n407 = x89 & ~x121 ;
  assign n408 = ~x88 & x120 ;
  assign n409 = x88 & ~x120 ;
  assign n410 = ~x87 & x119 ;
  assign n411 = x87 & ~x119 ;
  assign n412 = ~x86 & x118 ;
  assign n413 = x86 & ~x118 ;
  assign n414 = ~x85 & x117 ;
  assign n415 = x85 & ~x117 ;
  assign n416 = ~x84 & x116 ;
  assign n417 = x84 & ~x116 ;
  assign n418 = ~x83 & x115 ;
  assign n419 = x83 & ~x115 ;
  assign n420 = ~x82 & x114 ;
  assign n421 = x82 & ~x114 ;
  assign n422 = ~x81 & x113 ;
  assign n423 = x81 & ~x113 ;
  assign n424 = ~x80 & x112 ;
  assign n425 = x80 & ~x112 ;
  assign n426 = ~x79 & x111 ;
  assign n427 = x79 & ~x111 ;
  assign n428 = ~x78 & x110 ;
  assign n429 = x78 & ~x110 ;
  assign n430 = ~x77 & x109 ;
  assign n431 = x77 & ~x109 ;
  assign n432 = ~x76 & x108 ;
  assign n433 = x76 & ~x108 ;
  assign n434 = ~x75 & x107 ;
  assign n435 = x75 & ~x107 ;
  assign n436 = ~x74 & x106 ;
  assign n437 = x74 & ~x106 ;
  assign n438 = ~x73 & x105 ;
  assign n439 = x73 & ~x105 ;
  assign n440 = ~x72 & x104 ;
  assign n441 = x72 & ~x104 ;
  assign n442 = ~x71 & x103 ;
  assign n443 = x71 & ~x103 ;
  assign n444 = ~x70 & x102 ;
  assign n445 = x70 & ~x102 ;
  assign n446 = ~x69 & x101 ;
  assign n447 = x69 & ~x101 ;
  assign n448 = ~x68 & x100 ;
  assign n449 = x68 & ~x100 ;
  assign n450 = ~x67 & x99 ;
  assign n451 = x67 & ~x99 ;
  assign n452 = ~x66 & x98 ;
  assign n453 = x66 & ~x98 ;
  assign n454 = ~x65 & x97 ;
  assign n455 = x65 & ~x97 ;
  assign n456 = x64 & ~x96 ;
  assign n457 = ~n455 & ~n456 ;
  assign n458 = ~n454 & ~n457 ;
  assign n459 = ~n453 & ~n458 ;
  assign n460 = ~n452 & ~n459 ;
  assign n461 = ~n451 & ~n460 ;
  assign n462 = ~n450 & ~n461 ;
  assign n463 = ~n449 & ~n462 ;
  assign n464 = ~n448 & ~n463 ;
  assign n465 = ~n447 & ~n464 ;
  assign n466 = ~n446 & ~n465 ;
  assign n467 = ~n445 & ~n466 ;
  assign n468 = ~n444 & ~n467 ;
  assign n469 = ~n443 & ~n468 ;
  assign n470 = ~n442 & ~n469 ;
  assign n471 = ~n441 & ~n470 ;
  assign n472 = ~n440 & ~n471 ;
  assign n473 = ~n439 & ~n472 ;
  assign n474 = ~n438 & ~n473 ;
  assign n475 = ~n437 & ~n474 ;
  assign n476 = ~n436 & ~n475 ;
  assign n477 = ~n435 & ~n476 ;
  assign n478 = ~n434 & ~n477 ;
  assign n479 = ~n433 & ~n478 ;
  assign n480 = ~n432 & ~n479 ;
  assign n481 = ~n431 & ~n480 ;
  assign n482 = ~n430 & ~n481 ;
  assign n483 = ~n429 & ~n482 ;
  assign n484 = ~n428 & ~n483 ;
  assign n485 = ~n427 & ~n484 ;
  assign n486 = ~n426 & ~n485 ;
  assign n487 = ~n425 & ~n486 ;
  assign n488 = ~n424 & ~n487 ;
  assign n489 = ~n423 & ~n488 ;
  assign n490 = ~n422 & ~n489 ;
  assign n491 = ~n421 & ~n490 ;
  assign n492 = ~n420 & ~n491 ;
  assign n493 = ~n419 & ~n492 ;
  assign n494 = ~n418 & ~n493 ;
  assign n495 = ~n417 & ~n494 ;
  assign n496 = ~n416 & ~n495 ;
  assign n497 = ~n415 & ~n496 ;
  assign n498 = ~n414 & ~n497 ;
  assign n499 = ~n413 & ~n498 ;
  assign n500 = ~n412 & ~n499 ;
  assign n501 = ~n411 & ~n500 ;
  assign n502 = ~n410 & ~n501 ;
  assign n503 = ~n409 & ~n502 ;
  assign n504 = ~n408 & ~n503 ;
  assign n505 = ~n407 & ~n504 ;
  assign n506 = ~n406 & ~n505 ;
  assign n507 = ~n405 & ~n506 ;
  assign n508 = ~n404 & ~n507 ;
  assign n509 = ~n403 & ~n508 ;
  assign n510 = ~n402 & ~n509 ;
  assign n511 = ~n401 & ~n510 ;
  assign n512 = ~n400 & ~n511 ;
  assign n513 = ~n399 & ~n512 ;
  assign n514 = ~n398 & ~n513 ;
  assign n515 = ~n397 & ~n514 ;
  assign n516 = ~n396 & ~n515 ;
  assign n517 = ~n395 & ~n516 ;
  assign n518 = ~n394 & ~n517 ;
  assign n519 = x126 & ~n518 ;
  assign n520 = x94 & n518 ;
  assign n521 = ~n519 & ~n520 ;
  assign n522 = x62 & ~n388 ;
  assign n523 = x30 & n388 ;
  assign n524 = ~n522 & ~n523 ;
  assign n525 = ~n521 & n524 ;
  assign n526 = x97 & ~n518 ;
  assign n527 = x65 & n518 ;
  assign n528 = ~n526 & ~n527 ;
  assign n529 = n391 & ~n528 ;
  assign n530 = x96 & ~n518 ;
  assign n531 = x64 & n518 ;
  assign n532 = ~n530 & ~n531 ;
  assign n533 = x32 & ~n388 ;
  assign n534 = x0 & n388 ;
  assign n535 = ~n533 & ~n534 ;
  assign n536 = n532 & ~n535 ;
  assign n537 = ~n529 & n536 ;
  assign n538 = x98 & ~n518 ;
  assign n539 = x66 & n518 ;
  assign n540 = ~n538 & ~n539 ;
  assign n541 = x34 & ~n388 ;
  assign n542 = x2 & n388 ;
  assign n543 = ~n541 & ~n542 ;
  assign n544 = n540 & ~n543 ;
  assign n545 = ~n391 & n528 ;
  assign n546 = ~n544 & ~n545 ;
  assign n547 = ~n537 & n546 ;
  assign n548 = x35 & ~n388 ;
  assign n549 = x3 & n388 ;
  assign n550 = ~n548 & ~n549 ;
  assign n551 = x99 & ~n518 ;
  assign n552 = x67 & n518 ;
  assign n553 = ~n551 & ~n552 ;
  assign n554 = n550 & ~n553 ;
  assign n555 = ~n540 & n543 ;
  assign n556 = ~n554 & ~n555 ;
  assign n557 = ~n547 & n556 ;
  assign n558 = x100 & ~n518 ;
  assign n559 = x68 & n518 ;
  assign n560 = ~n558 & ~n559 ;
  assign n561 = x36 & ~n388 ;
  assign n562 = x4 & n388 ;
  assign n563 = ~n561 & ~n562 ;
  assign n564 = n560 & ~n563 ;
  assign n565 = ~n550 & n553 ;
  assign n566 = ~n564 & ~n565 ;
  assign n567 = ~n557 & n566 ;
  assign n568 = x101 & ~n518 ;
  assign n569 = x69 & n518 ;
  assign n570 = ~n568 & ~n569 ;
  assign n571 = x37 & ~n388 ;
  assign n572 = x5 & n388 ;
  assign n573 = ~n571 & ~n572 ;
  assign n574 = ~n570 & n573 ;
  assign n575 = ~n560 & n563 ;
  assign n576 = ~n574 & ~n575 ;
  assign n577 = ~n567 & n576 ;
  assign n578 = x38 & ~n388 ;
  assign n579 = x6 & n388 ;
  assign n580 = ~n578 & ~n579 ;
  assign n581 = x102 & ~n518 ;
  assign n582 = x70 & n518 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = ~n580 & n583 ;
  assign n585 = n570 & ~n573 ;
  assign n586 = ~n584 & ~n585 ;
  assign n587 = ~n577 & n586 ;
  assign n588 = x39 & ~n388 ;
  assign n589 = x7 & n388 ;
  assign n590 = ~n588 & ~n589 ;
  assign n591 = x103 & ~n518 ;
  assign n592 = x71 & n518 ;
  assign n593 = ~n591 & ~n592 ;
  assign n594 = n590 & ~n593 ;
  assign n595 = n580 & ~n583 ;
  assign n596 = ~n594 & ~n595 ;
  assign n597 = ~n587 & n596 ;
  assign n598 = ~n590 & n593 ;
  assign n599 = x104 & ~n518 ;
  assign n600 = x72 & n518 ;
  assign n601 = ~n599 & ~n600 ;
  assign n602 = x40 & ~n388 ;
  assign n603 = x8 & n388 ;
  assign n604 = ~n602 & ~n603 ;
  assign n605 = n601 & ~n604 ;
  assign n606 = ~n598 & ~n605 ;
  assign n607 = ~n597 & n606 ;
  assign n608 = ~n601 & n604 ;
  assign n609 = x105 & ~n518 ;
  assign n610 = x73 & n518 ;
  assign n611 = ~n609 & ~n610 ;
  assign n612 = x41 & ~n388 ;
  assign n613 = x9 & n388 ;
  assign n614 = ~n612 & ~n613 ;
  assign n615 = ~n611 & n614 ;
  assign n616 = ~n608 & ~n615 ;
  assign n617 = ~n607 & n616 ;
  assign n618 = n611 & ~n614 ;
  assign n619 = x42 & ~n388 ;
  assign n620 = x10 & n388 ;
  assign n621 = ~n619 & ~n620 ;
  assign n622 = x106 & ~n518 ;
  assign n623 = x74 & n518 ;
  assign n624 = ~n622 & ~n623 ;
  assign n625 = ~n621 & n624 ;
  assign n626 = ~n618 & ~n625 ;
  assign n627 = ~n617 & n626 ;
  assign n628 = x43 & ~n388 ;
  assign n629 = x11 & n388 ;
  assign n630 = ~n628 & ~n629 ;
  assign n631 = x107 & ~n518 ;
  assign n632 = x75 & n518 ;
  assign n633 = ~n631 & ~n632 ;
  assign n634 = n630 & ~n633 ;
  assign n635 = n621 & ~n624 ;
  assign n636 = ~n634 & ~n635 ;
  assign n637 = ~n627 & n636 ;
  assign n638 = x108 & ~n518 ;
  assign n639 = x76 & n518 ;
  assign n640 = ~n638 & ~n639 ;
  assign n641 = x44 & ~n388 ;
  assign n642 = x12 & n388 ;
  assign n643 = ~n641 & ~n642 ;
  assign n644 = n640 & ~n643 ;
  assign n645 = ~n630 & n633 ;
  assign n646 = ~n644 & ~n645 ;
  assign n647 = ~n637 & n646 ;
  assign n648 = ~n640 & n643 ;
  assign n649 = x109 & ~n518 ;
  assign n650 = x77 & n518 ;
  assign n651 = ~n649 & ~n650 ;
  assign n652 = x45 & ~n388 ;
  assign n653 = x13 & n388 ;
  assign n654 = ~n652 & ~n653 ;
  assign n655 = ~n651 & n654 ;
  assign n656 = ~n648 & ~n655 ;
  assign n657 = ~n647 & n656 ;
  assign n658 = n651 & ~n654 ;
  assign n659 = x46 & ~n388 ;
  assign n660 = x14 & n388 ;
  assign n661 = ~n659 & ~n660 ;
  assign n662 = x110 & ~n518 ;
  assign n663 = x78 & n518 ;
  assign n664 = ~n662 & ~n663 ;
  assign n665 = ~n661 & n664 ;
  assign n666 = ~n658 & ~n665 ;
  assign n667 = ~n657 & n666 ;
  assign n668 = x47 & ~n388 ;
  assign n669 = x15 & n388 ;
  assign n670 = ~n668 & ~n669 ;
  assign n671 = x111 & ~n518 ;
  assign n672 = x79 & n518 ;
  assign n673 = ~n671 & ~n672 ;
  assign n674 = n670 & ~n673 ;
  assign n675 = n661 & ~n664 ;
  assign n676 = ~n674 & ~n675 ;
  assign n677 = ~n667 & n676 ;
  assign n678 = x112 & ~n518 ;
  assign n679 = x80 & n518 ;
  assign n680 = ~n678 & ~n679 ;
  assign n681 = x48 & ~n388 ;
  assign n682 = x16 & n388 ;
  assign n683 = ~n681 & ~n682 ;
  assign n684 = n680 & ~n683 ;
  assign n685 = ~n670 & n673 ;
  assign n686 = ~n684 & ~n685 ;
  assign n687 = ~n677 & n686 ;
  assign n688 = ~n680 & n683 ;
  assign n689 = x113 & ~n518 ;
  assign n690 = x81 & n518 ;
  assign n691 = ~n689 & ~n690 ;
  assign n692 = x49 & ~n388 ;
  assign n693 = x17 & n388 ;
  assign n694 = ~n692 & ~n693 ;
  assign n695 = ~n691 & n694 ;
  assign n696 = ~n688 & ~n695 ;
  assign n697 = ~n687 & n696 ;
  assign n698 = n691 & ~n694 ;
  assign n699 = x50 & ~n388 ;
  assign n700 = x18 & n388 ;
  assign n701 = ~n699 & ~n700 ;
  assign n702 = x114 & ~n518 ;
  assign n703 = x82 & n518 ;
  assign n704 = ~n702 & ~n703 ;
  assign n705 = ~n701 & n704 ;
  assign n706 = ~n698 & ~n705 ;
  assign n707 = ~n697 & n706 ;
  assign n708 = x51 & ~n388 ;
  assign n709 = x19 & n388 ;
  assign n710 = ~n708 & ~n709 ;
  assign n711 = x115 & ~n518 ;
  assign n712 = x83 & n518 ;
  assign n713 = ~n711 & ~n712 ;
  assign n714 = n710 & ~n713 ;
  assign n715 = n701 & ~n704 ;
  assign n716 = ~n714 & ~n715 ;
  assign n717 = ~n707 & n716 ;
  assign n718 = x116 & ~n518 ;
  assign n719 = x84 & n518 ;
  assign n720 = ~n718 & ~n719 ;
  assign n721 = x52 & ~n388 ;
  assign n722 = x20 & n388 ;
  assign n723 = ~n721 & ~n722 ;
  assign n724 = n720 & ~n723 ;
  assign n725 = ~n710 & n713 ;
  assign n726 = ~n724 & ~n725 ;
  assign n727 = ~n717 & n726 ;
  assign n728 = ~n720 & n723 ;
  assign n729 = x117 & ~n518 ;
  assign n730 = x85 & n518 ;
  assign n731 = ~n729 & ~n730 ;
  assign n732 = x53 & ~n388 ;
  assign n733 = x21 & n388 ;
  assign n734 = ~n732 & ~n733 ;
  assign n735 = ~n731 & n734 ;
  assign n736 = ~n728 & ~n735 ;
  assign n737 = ~n727 & n736 ;
  assign n738 = n731 & ~n734 ;
  assign n739 = x54 & ~n388 ;
  assign n740 = x22 & n388 ;
  assign n741 = ~n739 & ~n740 ;
  assign n742 = x118 & ~n518 ;
  assign n743 = x86 & n518 ;
  assign n744 = ~n742 & ~n743 ;
  assign n745 = ~n741 & n744 ;
  assign n746 = ~n738 & ~n745 ;
  assign n747 = ~n737 & n746 ;
  assign n748 = x55 & ~n388 ;
  assign n749 = x23 & n388 ;
  assign n750 = ~n748 & ~n749 ;
  assign n751 = x119 & ~n518 ;
  assign n752 = x87 & n518 ;
  assign n753 = ~n751 & ~n752 ;
  assign n754 = n750 & ~n753 ;
  assign n755 = n741 & ~n744 ;
  assign n756 = ~n754 & ~n755 ;
  assign n757 = ~n747 & n756 ;
  assign n758 = x56 & ~n388 ;
  assign n759 = x24 & n388 ;
  assign n760 = ~n758 & ~n759 ;
  assign n761 = x120 & ~n518 ;
  assign n762 = x88 & n518 ;
  assign n763 = ~n761 & ~n762 ;
  assign n764 = ~n760 & n763 ;
  assign n765 = ~n750 & n753 ;
  assign n766 = ~n764 & ~n765 ;
  assign n767 = ~n757 & n766 ;
  assign n768 = n760 & ~n763 ;
  assign n769 = x121 & ~n518 ;
  assign n770 = x89 & n518 ;
  assign n771 = ~n769 & ~n770 ;
  assign n772 = x57 & ~n388 ;
  assign n773 = x25 & n388 ;
  assign n774 = ~n772 & ~n773 ;
  assign n775 = ~n771 & n774 ;
  assign n776 = ~n768 & ~n775 ;
  assign n777 = ~n767 & n776 ;
  assign n778 = n771 & ~n774 ;
  assign n779 = x58 & ~n388 ;
  assign n780 = x26 & n388 ;
  assign n781 = ~n779 & ~n780 ;
  assign n782 = x122 & ~n518 ;
  assign n783 = x90 & n518 ;
  assign n784 = ~n782 & ~n783 ;
  assign n785 = ~n781 & n784 ;
  assign n786 = ~n778 & ~n785 ;
  assign n787 = ~n777 & n786 ;
  assign n788 = x59 & ~n388 ;
  assign n789 = x27 & n388 ;
  assign n790 = ~n788 & ~n789 ;
  assign n791 = x123 & ~n518 ;
  assign n792 = x91 & n518 ;
  assign n793 = ~n791 & ~n792 ;
  assign n794 = n790 & ~n793 ;
  assign n795 = n781 & ~n784 ;
  assign n796 = ~n794 & ~n795 ;
  assign n797 = ~n787 & n796 ;
  assign n798 = x124 & ~n518 ;
  assign n799 = x92 & n518 ;
  assign n800 = ~n798 & ~n799 ;
  assign n801 = x60 & ~n388 ;
  assign n802 = x28 & n388 ;
  assign n803 = ~n801 & ~n802 ;
  assign n804 = n800 & ~n803 ;
  assign n805 = ~n790 & n793 ;
  assign n806 = ~n804 & ~n805 ;
  assign n807 = ~n797 & n806 ;
  assign n808 = ~n800 & n803 ;
  assign n809 = x61 & ~n388 ;
  assign n810 = x29 & n388 ;
  assign n811 = ~n809 & ~n810 ;
  assign n812 = x125 & ~n518 ;
  assign n813 = x93 & n518 ;
  assign n814 = ~n812 & ~n813 ;
  assign n815 = n811 & ~n814 ;
  assign n816 = ~n808 & ~n815 ;
  assign n817 = ~n807 & n816 ;
  assign n818 = n521 & ~n524 ;
  assign n819 = ~n811 & n814 ;
  assign n820 = ~n818 & ~n819 ;
  assign n821 = ~n817 & n820 ;
  assign n822 = ~n525 & ~n821 ;
  assign n823 = ~n393 & ~n822 ;
  assign n824 = ~n392 & ~n823 ;
  assign n825 = ~n391 & n824 ;
  assign n826 = ~n528 & ~n824 ;
  assign n827 = ~n825 & ~n826 ;
  assign n828 = ~x159 & x191 ;
  assign n829 = x159 & ~x191 ;
  assign n830 = ~x158 & x190 ;
  assign n831 = x158 & ~x190 ;
  assign n832 = ~x157 & x189 ;
  assign n833 = x157 & ~x189 ;
  assign n834 = ~x156 & x188 ;
  assign n835 = x156 & ~x188 ;
  assign n836 = ~x155 & x187 ;
  assign n837 = x155 & ~x187 ;
  assign n838 = ~x154 & x186 ;
  assign n839 = x154 & ~x186 ;
  assign n840 = ~x153 & x185 ;
  assign n841 = x153 & ~x185 ;
  assign n842 = ~x152 & x184 ;
  assign n843 = x152 & ~x184 ;
  assign n844 = ~x151 & x183 ;
  assign n845 = x151 & ~x183 ;
  assign n846 = ~x150 & x182 ;
  assign n847 = x150 & ~x182 ;
  assign n848 = ~x149 & x181 ;
  assign n849 = x149 & ~x181 ;
  assign n850 = ~x148 & x180 ;
  assign n851 = x148 & ~x180 ;
  assign n852 = ~x147 & x179 ;
  assign n853 = x147 & ~x179 ;
  assign n854 = ~x146 & x178 ;
  assign n855 = x146 & ~x178 ;
  assign n856 = ~x145 & x177 ;
  assign n857 = x145 & ~x177 ;
  assign n858 = ~x144 & x176 ;
  assign n859 = x144 & ~x176 ;
  assign n860 = ~x143 & x175 ;
  assign n861 = x143 & ~x175 ;
  assign n862 = ~x142 & x174 ;
  assign n863 = x142 & ~x174 ;
  assign n864 = ~x141 & x173 ;
  assign n865 = x141 & ~x173 ;
  assign n866 = ~x140 & x172 ;
  assign n867 = x140 & ~x172 ;
  assign n868 = ~x139 & x171 ;
  assign n869 = x139 & ~x171 ;
  assign n870 = ~x138 & x170 ;
  assign n871 = x138 & ~x170 ;
  assign n872 = ~x137 & x169 ;
  assign n873 = x137 & ~x169 ;
  assign n874 = ~x136 & x168 ;
  assign n875 = x136 & ~x168 ;
  assign n876 = ~x135 & x167 ;
  assign n877 = x135 & ~x167 ;
  assign n878 = ~x134 & x166 ;
  assign n879 = x134 & ~x166 ;
  assign n880 = ~x133 & x165 ;
  assign n881 = x133 & ~x165 ;
  assign n882 = ~x132 & x164 ;
  assign n883 = x132 & ~x164 ;
  assign n884 = ~x131 & x163 ;
  assign n885 = x131 & ~x163 ;
  assign n886 = ~x130 & x162 ;
  assign n887 = x130 & ~x162 ;
  assign n888 = ~x129 & x161 ;
  assign n889 = x129 & ~x161 ;
  assign n890 = x128 & ~x160 ;
  assign n891 = ~n889 & ~n890 ;
  assign n892 = ~n888 & ~n891 ;
  assign n893 = ~n887 & ~n892 ;
  assign n894 = ~n886 & ~n893 ;
  assign n895 = ~n885 & ~n894 ;
  assign n896 = ~n884 & ~n895 ;
  assign n897 = ~n883 & ~n896 ;
  assign n898 = ~n882 & ~n897 ;
  assign n899 = ~n881 & ~n898 ;
  assign n900 = ~n880 & ~n899 ;
  assign n901 = ~n879 & ~n900 ;
  assign n902 = ~n878 & ~n901 ;
  assign n903 = ~n877 & ~n902 ;
  assign n904 = ~n876 & ~n903 ;
  assign n905 = ~n875 & ~n904 ;
  assign n906 = ~n874 & ~n905 ;
  assign n907 = ~n873 & ~n906 ;
  assign n908 = ~n872 & ~n907 ;
  assign n909 = ~n871 & ~n908 ;
  assign n910 = ~n870 & ~n909 ;
  assign n911 = ~n869 & ~n910 ;
  assign n912 = ~n868 & ~n911 ;
  assign n913 = ~n867 & ~n912 ;
  assign n914 = ~n866 & ~n913 ;
  assign n915 = ~n865 & ~n914 ;
  assign n916 = ~n864 & ~n915 ;
  assign n917 = ~n863 & ~n916 ;
  assign n918 = ~n862 & ~n917 ;
  assign n919 = ~n861 & ~n918 ;
  assign n920 = ~n860 & ~n919 ;
  assign n921 = ~n859 & ~n920 ;
  assign n922 = ~n858 & ~n921 ;
  assign n923 = ~n857 & ~n922 ;
  assign n924 = ~n856 & ~n923 ;
  assign n925 = ~n855 & ~n924 ;
  assign n926 = ~n854 & ~n925 ;
  assign n927 = ~n853 & ~n926 ;
  assign n928 = ~n852 & ~n927 ;
  assign n929 = ~n851 & ~n928 ;
  assign n930 = ~n850 & ~n929 ;
  assign n931 = ~n849 & ~n930 ;
  assign n932 = ~n848 & ~n931 ;
  assign n933 = ~n847 & ~n932 ;
  assign n934 = ~n846 & ~n933 ;
  assign n935 = ~n845 & ~n934 ;
  assign n936 = ~n844 & ~n935 ;
  assign n937 = ~n843 & ~n936 ;
  assign n938 = ~n842 & ~n937 ;
  assign n939 = ~n841 & ~n938 ;
  assign n940 = ~n840 & ~n939 ;
  assign n941 = ~n839 & ~n940 ;
  assign n942 = ~n838 & ~n941 ;
  assign n943 = ~n837 & ~n942 ;
  assign n944 = ~n836 & ~n943 ;
  assign n945 = ~n835 & ~n944 ;
  assign n946 = ~n834 & ~n945 ;
  assign n947 = ~n833 & ~n946 ;
  assign n948 = ~n832 & ~n947 ;
  assign n949 = ~n831 & ~n948 ;
  assign n950 = ~n830 & ~n949 ;
  assign n951 = ~n829 & ~n950 ;
  assign n952 = ~n828 & ~n951 ;
  assign n953 = x161 & ~n952 ;
  assign n954 = x129 & n952 ;
  assign n955 = ~n953 & ~n954 ;
  assign n956 = n257 & ~n258 ;
  assign n957 = ~n257 & n258 ;
  assign n958 = ~x223 & x255 ;
  assign n959 = x223 & ~x255 ;
  assign n960 = ~x222 & x254 ;
  assign n961 = x222 & ~x254 ;
  assign n962 = ~x221 & x253 ;
  assign n963 = x221 & ~x253 ;
  assign n964 = ~x220 & x252 ;
  assign n965 = x220 & ~x252 ;
  assign n966 = ~x219 & x251 ;
  assign n967 = x219 & ~x251 ;
  assign n968 = ~x218 & x250 ;
  assign n969 = x218 & ~x250 ;
  assign n970 = ~x217 & x249 ;
  assign n971 = x217 & ~x249 ;
  assign n972 = ~x216 & x248 ;
  assign n973 = x216 & ~x248 ;
  assign n974 = ~x215 & x247 ;
  assign n975 = x215 & ~x247 ;
  assign n976 = ~x214 & x246 ;
  assign n977 = x214 & ~x246 ;
  assign n978 = ~x213 & x245 ;
  assign n979 = x213 & ~x245 ;
  assign n980 = ~x212 & x244 ;
  assign n981 = x212 & ~x244 ;
  assign n982 = ~x211 & x243 ;
  assign n983 = x211 & ~x243 ;
  assign n984 = ~x210 & x242 ;
  assign n985 = x210 & ~x242 ;
  assign n986 = ~x209 & x241 ;
  assign n987 = x209 & ~x241 ;
  assign n988 = ~x208 & x240 ;
  assign n989 = x208 & ~x240 ;
  assign n990 = ~x207 & x239 ;
  assign n991 = x207 & ~x239 ;
  assign n992 = ~x206 & x238 ;
  assign n993 = x206 & ~x238 ;
  assign n994 = ~x205 & x237 ;
  assign n995 = x205 & ~x237 ;
  assign n996 = ~x204 & x236 ;
  assign n997 = x204 & ~x236 ;
  assign n998 = ~x203 & x235 ;
  assign n999 = x203 & ~x235 ;
  assign n1000 = ~x202 & x234 ;
  assign n1001 = x202 & ~x234 ;
  assign n1002 = ~x201 & x233 ;
  assign n1003 = x201 & ~x233 ;
  assign n1004 = ~x200 & x232 ;
  assign n1005 = x200 & ~x232 ;
  assign n1006 = ~x199 & x231 ;
  assign n1007 = x199 & ~x231 ;
  assign n1008 = ~x198 & x230 ;
  assign n1009 = x198 & ~x230 ;
  assign n1010 = ~x197 & x229 ;
  assign n1011 = x197 & ~x229 ;
  assign n1012 = ~x196 & x228 ;
  assign n1013 = x196 & ~x228 ;
  assign n1014 = ~x195 & x227 ;
  assign n1015 = x195 & ~x227 ;
  assign n1016 = ~x194 & x226 ;
  assign n1017 = x194 & ~x226 ;
  assign n1018 = ~x193 & x225 ;
  assign n1019 = x193 & ~x225 ;
  assign n1020 = x192 & ~x224 ;
  assign n1021 = ~n1019 & ~n1020 ;
  assign n1022 = ~n1018 & ~n1021 ;
  assign n1023 = ~n1017 & ~n1022 ;
  assign n1024 = ~n1016 & ~n1023 ;
  assign n1025 = ~n1015 & ~n1024 ;
  assign n1026 = ~n1014 & ~n1025 ;
  assign n1027 = ~n1013 & ~n1026 ;
  assign n1028 = ~n1012 & ~n1027 ;
  assign n1029 = ~n1011 & ~n1028 ;
  assign n1030 = ~n1010 & ~n1029 ;
  assign n1031 = ~n1009 & ~n1030 ;
  assign n1032 = ~n1008 & ~n1031 ;
  assign n1033 = ~n1007 & ~n1032 ;
  assign n1034 = ~n1006 & ~n1033 ;
  assign n1035 = ~n1005 & ~n1034 ;
  assign n1036 = ~n1004 & ~n1035 ;
  assign n1037 = ~n1003 & ~n1036 ;
  assign n1038 = ~n1002 & ~n1037 ;
  assign n1039 = ~n1001 & ~n1038 ;
  assign n1040 = ~n1000 & ~n1039 ;
  assign n1041 = ~n999 & ~n1040 ;
  assign n1042 = ~n998 & ~n1041 ;
  assign n1043 = ~n997 & ~n1042 ;
  assign n1044 = ~n996 & ~n1043 ;
  assign n1045 = ~n995 & ~n1044 ;
  assign n1046 = ~n994 & ~n1045 ;
  assign n1047 = ~n993 & ~n1046 ;
  assign n1048 = ~n992 & ~n1047 ;
  assign n1049 = ~n991 & ~n1048 ;
  assign n1050 = ~n990 & ~n1049 ;
  assign n1051 = ~n989 & ~n1050 ;
  assign n1052 = ~n988 & ~n1051 ;
  assign n1053 = ~n987 & ~n1052 ;
  assign n1054 = ~n986 & ~n1053 ;
  assign n1055 = ~n985 & ~n1054 ;
  assign n1056 = ~n984 & ~n1055 ;
  assign n1057 = ~n983 & ~n1056 ;
  assign n1058 = ~n982 & ~n1057 ;
  assign n1059 = ~n981 & ~n1058 ;
  assign n1060 = ~n980 & ~n1059 ;
  assign n1061 = ~n979 & ~n1060 ;
  assign n1062 = ~n978 & ~n1061 ;
  assign n1063 = ~n977 & ~n1062 ;
  assign n1064 = ~n976 & ~n1063 ;
  assign n1065 = ~n975 & ~n1064 ;
  assign n1066 = ~n974 & ~n1065 ;
  assign n1067 = ~n973 & ~n1066 ;
  assign n1068 = ~n972 & ~n1067 ;
  assign n1069 = ~n971 & ~n1068 ;
  assign n1070 = ~n970 & ~n1069 ;
  assign n1071 = ~n969 & ~n1070 ;
  assign n1072 = ~n968 & ~n1071 ;
  assign n1073 = ~n967 & ~n1072 ;
  assign n1074 = ~n966 & ~n1073 ;
  assign n1075 = ~n965 & ~n1074 ;
  assign n1076 = ~n964 & ~n1075 ;
  assign n1077 = ~n963 & ~n1076 ;
  assign n1078 = ~n962 & ~n1077 ;
  assign n1079 = ~n961 & ~n1078 ;
  assign n1080 = ~n960 & ~n1079 ;
  assign n1081 = ~n959 & ~n1080 ;
  assign n1082 = ~n958 & ~n1081 ;
  assign n1083 = x225 & ~n1082 ;
  assign n1084 = x193 & n1082 ;
  assign n1085 = ~n1083 & ~n1084 ;
  assign n1086 = n955 & ~n1085 ;
  assign n1087 = x224 & ~n1082 ;
  assign n1088 = x192 & n1082 ;
  assign n1089 = ~n1087 & ~n1088 ;
  assign n1090 = x160 & ~n952 ;
  assign n1091 = x128 & n952 ;
  assign n1092 = ~n1090 & ~n1091 ;
  assign n1093 = n1089 & ~n1092 ;
  assign n1094 = ~n1086 & n1093 ;
  assign n1095 = x226 & ~n1082 ;
  assign n1096 = x194 & n1082 ;
  assign n1097 = ~n1095 & ~n1096 ;
  assign n1098 = x162 & ~n952 ;
  assign n1099 = x130 & n952 ;
  assign n1100 = ~n1098 & ~n1099 ;
  assign n1101 = n1097 & ~n1100 ;
  assign n1102 = ~n955 & n1085 ;
  assign n1103 = ~n1101 & ~n1102 ;
  assign n1104 = ~n1094 & n1103 ;
  assign n1105 = ~n1097 & n1100 ;
  assign n1106 = x227 & ~n1082 ;
  assign n1107 = x195 & n1082 ;
  assign n1108 = ~n1106 & ~n1107 ;
  assign n1109 = x163 & ~n952 ;
  assign n1110 = x131 & n952 ;
  assign n1111 = ~n1109 & ~n1110 ;
  assign n1112 = ~n1108 & n1111 ;
  assign n1113 = ~n1105 & ~n1112 ;
  assign n1114 = ~n1104 & n1113 ;
  assign n1115 = x164 & ~n952 ;
  assign n1116 = x132 & n952 ;
  assign n1117 = ~n1115 & ~n1116 ;
  assign n1118 = x228 & ~n1082 ;
  assign n1119 = x196 & n1082 ;
  assign n1120 = ~n1118 & ~n1119 ;
  assign n1121 = ~n1117 & n1120 ;
  assign n1122 = n1108 & ~n1111 ;
  assign n1123 = ~n1121 & ~n1122 ;
  assign n1124 = ~n1114 & n1123 ;
  assign n1125 = x229 & ~n1082 ;
  assign n1126 = x197 & n1082 ;
  assign n1127 = ~n1125 & ~n1126 ;
  assign n1128 = x165 & ~n952 ;
  assign n1129 = x133 & n952 ;
  assign n1130 = ~n1128 & ~n1129 ;
  assign n1131 = ~n1127 & n1130 ;
  assign n1132 = n1117 & ~n1120 ;
  assign n1133 = ~n1131 & ~n1132 ;
  assign n1134 = ~n1124 & n1133 ;
  assign n1135 = x230 & ~n1082 ;
  assign n1136 = x198 & n1082 ;
  assign n1137 = ~n1135 & ~n1136 ;
  assign n1138 = x166 & ~n952 ;
  assign n1139 = x134 & n952 ;
  assign n1140 = ~n1138 & ~n1139 ;
  assign n1141 = n1137 & ~n1140 ;
  assign n1142 = n1127 & ~n1130 ;
  assign n1143 = ~n1141 & ~n1142 ;
  assign n1144 = ~n1134 & n1143 ;
  assign n1145 = ~n1137 & n1140 ;
  assign n1146 = x167 & ~n952 ;
  assign n1147 = x135 & n952 ;
  assign n1148 = ~n1146 & ~n1147 ;
  assign n1149 = x231 & ~n1082 ;
  assign n1150 = x199 & n1082 ;
  assign n1151 = ~n1149 & ~n1150 ;
  assign n1152 = n1148 & ~n1151 ;
  assign n1153 = ~n1145 & ~n1152 ;
  assign n1154 = ~n1144 & n1153 ;
  assign n1155 = ~n1148 & n1151 ;
  assign n1156 = x232 & ~n1082 ;
  assign n1157 = x200 & n1082 ;
  assign n1158 = ~n1156 & ~n1157 ;
  assign n1159 = x168 & ~n952 ;
  assign n1160 = x136 & n952 ;
  assign n1161 = ~n1159 & ~n1160 ;
  assign n1162 = n1158 & ~n1161 ;
  assign n1163 = ~n1155 & ~n1162 ;
  assign n1164 = ~n1154 & n1163 ;
  assign n1165 = ~n1158 & n1161 ;
  assign n1166 = x233 & ~n1082 ;
  assign n1167 = x201 & n1082 ;
  assign n1168 = ~n1166 & ~n1167 ;
  assign n1169 = x169 & ~n952 ;
  assign n1170 = x137 & n952 ;
  assign n1171 = ~n1169 & ~n1170 ;
  assign n1172 = ~n1168 & n1171 ;
  assign n1173 = ~n1165 & ~n1172 ;
  assign n1174 = ~n1164 & n1173 ;
  assign n1175 = n1168 & ~n1171 ;
  assign n1176 = x170 & ~n952 ;
  assign n1177 = x138 & n952 ;
  assign n1178 = ~n1176 & ~n1177 ;
  assign n1179 = x234 & ~n1082 ;
  assign n1180 = x202 & n1082 ;
  assign n1181 = ~n1179 & ~n1180 ;
  assign n1182 = ~n1178 & n1181 ;
  assign n1183 = ~n1175 & ~n1182 ;
  assign n1184 = ~n1174 & n1183 ;
  assign n1185 = x171 & ~n952 ;
  assign n1186 = x139 & n952 ;
  assign n1187 = ~n1185 & ~n1186 ;
  assign n1188 = x235 & ~n1082 ;
  assign n1189 = x203 & n1082 ;
  assign n1190 = ~n1188 & ~n1189 ;
  assign n1191 = n1187 & ~n1190 ;
  assign n1192 = n1178 & ~n1181 ;
  assign n1193 = ~n1191 & ~n1192 ;
  assign n1194 = ~n1184 & n1193 ;
  assign n1195 = x236 & ~n1082 ;
  assign n1196 = x204 & n1082 ;
  assign n1197 = ~n1195 & ~n1196 ;
  assign n1198 = x172 & ~n952 ;
  assign n1199 = x140 & n952 ;
  assign n1200 = ~n1198 & ~n1199 ;
  assign n1201 = n1197 & ~n1200 ;
  assign n1202 = ~n1187 & n1190 ;
  assign n1203 = ~n1201 & ~n1202 ;
  assign n1204 = ~n1194 & n1203 ;
  assign n1205 = ~n1197 & n1200 ;
  assign n1206 = x237 & ~n1082 ;
  assign n1207 = x205 & n1082 ;
  assign n1208 = ~n1206 & ~n1207 ;
  assign n1209 = x173 & ~n952 ;
  assign n1210 = x141 & n952 ;
  assign n1211 = ~n1209 & ~n1210 ;
  assign n1212 = ~n1208 & n1211 ;
  assign n1213 = ~n1205 & ~n1212 ;
  assign n1214 = ~n1204 & n1213 ;
  assign n1215 = n1208 & ~n1211 ;
  assign n1216 = x174 & ~n952 ;
  assign n1217 = x142 & n952 ;
  assign n1218 = ~n1216 & ~n1217 ;
  assign n1219 = x238 & ~n1082 ;
  assign n1220 = x206 & n1082 ;
  assign n1221 = ~n1219 & ~n1220 ;
  assign n1222 = ~n1218 & n1221 ;
  assign n1223 = ~n1215 & ~n1222 ;
  assign n1224 = ~n1214 & n1223 ;
  assign n1225 = x175 & ~n952 ;
  assign n1226 = x143 & n952 ;
  assign n1227 = ~n1225 & ~n1226 ;
  assign n1228 = x239 & ~n1082 ;
  assign n1229 = x207 & n1082 ;
  assign n1230 = ~n1228 & ~n1229 ;
  assign n1231 = n1227 & ~n1230 ;
  assign n1232 = n1218 & ~n1221 ;
  assign n1233 = ~n1231 & ~n1232 ;
  assign n1234 = ~n1224 & n1233 ;
  assign n1235 = x240 & ~n1082 ;
  assign n1236 = x208 & n1082 ;
  assign n1237 = ~n1235 & ~n1236 ;
  assign n1238 = x176 & ~n952 ;
  assign n1239 = x144 & n952 ;
  assign n1240 = ~n1238 & ~n1239 ;
  assign n1241 = n1237 & ~n1240 ;
  assign n1242 = ~n1227 & n1230 ;
  assign n1243 = ~n1241 & ~n1242 ;
  assign n1244 = ~n1234 & n1243 ;
  assign n1245 = ~n1237 & n1240 ;
  assign n1246 = x241 & ~n1082 ;
  assign n1247 = x209 & n1082 ;
  assign n1248 = ~n1246 & ~n1247 ;
  assign n1249 = x177 & ~n952 ;
  assign n1250 = x145 & n952 ;
  assign n1251 = ~n1249 & ~n1250 ;
  assign n1252 = ~n1248 & n1251 ;
  assign n1253 = ~n1245 & ~n1252 ;
  assign n1254 = ~n1244 & n1253 ;
  assign n1255 = n1248 & ~n1251 ;
  assign n1256 = x178 & ~n952 ;
  assign n1257 = x146 & n952 ;
  assign n1258 = ~n1256 & ~n1257 ;
  assign n1259 = x242 & ~n1082 ;
  assign n1260 = x210 & n1082 ;
  assign n1261 = ~n1259 & ~n1260 ;
  assign n1262 = ~n1258 & n1261 ;
  assign n1263 = ~n1255 & ~n1262 ;
  assign n1264 = ~n1254 & n1263 ;
  assign n1265 = x179 & ~n952 ;
  assign n1266 = x147 & n952 ;
  assign n1267 = ~n1265 & ~n1266 ;
  assign n1268 = x243 & ~n1082 ;
  assign n1269 = x211 & n1082 ;
  assign n1270 = ~n1268 & ~n1269 ;
  assign n1271 = n1267 & ~n1270 ;
  assign n1272 = n1258 & ~n1261 ;
  assign n1273 = ~n1271 & ~n1272 ;
  assign n1274 = ~n1264 & n1273 ;
  assign n1275 = x244 & ~n1082 ;
  assign n1276 = x212 & n1082 ;
  assign n1277 = ~n1275 & ~n1276 ;
  assign n1278 = x180 & ~n952 ;
  assign n1279 = x148 & n952 ;
  assign n1280 = ~n1278 & ~n1279 ;
  assign n1281 = n1277 & ~n1280 ;
  assign n1282 = ~n1267 & n1270 ;
  assign n1283 = ~n1281 & ~n1282 ;
  assign n1284 = ~n1274 & n1283 ;
  assign n1285 = ~n1277 & n1280 ;
  assign n1286 = x245 & ~n1082 ;
  assign n1287 = x213 & n1082 ;
  assign n1288 = ~n1286 & ~n1287 ;
  assign n1289 = x181 & ~n952 ;
  assign n1290 = x149 & n952 ;
  assign n1291 = ~n1289 & ~n1290 ;
  assign n1292 = ~n1288 & n1291 ;
  assign n1293 = ~n1285 & ~n1292 ;
  assign n1294 = ~n1284 & n1293 ;
  assign n1295 = n1288 & ~n1291 ;
  assign n1296 = x182 & ~n952 ;
  assign n1297 = x150 & n952 ;
  assign n1298 = ~n1296 & ~n1297 ;
  assign n1299 = x246 & ~n1082 ;
  assign n1300 = x214 & n1082 ;
  assign n1301 = ~n1299 & ~n1300 ;
  assign n1302 = ~n1298 & n1301 ;
  assign n1303 = ~n1295 & ~n1302 ;
  assign n1304 = ~n1294 & n1303 ;
  assign n1305 = x183 & ~n952 ;
  assign n1306 = x151 & n952 ;
  assign n1307 = ~n1305 & ~n1306 ;
  assign n1308 = x247 & ~n1082 ;
  assign n1309 = x215 & n1082 ;
  assign n1310 = ~n1308 & ~n1309 ;
  assign n1311 = n1307 & ~n1310 ;
  assign n1312 = n1298 & ~n1301 ;
  assign n1313 = ~n1311 & ~n1312 ;
  assign n1314 = ~n1304 & n1313 ;
  assign n1315 = x248 & ~n1082 ;
  assign n1316 = x216 & n1082 ;
  assign n1317 = ~n1315 & ~n1316 ;
  assign n1318 = x184 & ~n952 ;
  assign n1319 = x152 & n952 ;
  assign n1320 = ~n1318 & ~n1319 ;
  assign n1321 = n1317 & ~n1320 ;
  assign n1322 = ~n1307 & n1310 ;
  assign n1323 = ~n1321 & ~n1322 ;
  assign n1324 = ~n1314 & n1323 ;
  assign n1325 = ~n1317 & n1320 ;
  assign n1326 = x249 & ~n1082 ;
  assign n1327 = x217 & n1082 ;
  assign n1328 = ~n1326 & ~n1327 ;
  assign n1329 = x185 & ~n952 ;
  assign n1330 = x153 & n952 ;
  assign n1331 = ~n1329 & ~n1330 ;
  assign n1332 = ~n1328 & n1331 ;
  assign n1333 = ~n1325 & ~n1332 ;
  assign n1334 = ~n1324 & n1333 ;
  assign n1335 = n1328 & ~n1331 ;
  assign n1336 = x186 & ~n952 ;
  assign n1337 = x154 & n952 ;
  assign n1338 = ~n1336 & ~n1337 ;
  assign n1339 = x250 & ~n1082 ;
  assign n1340 = x218 & n1082 ;
  assign n1341 = ~n1339 & ~n1340 ;
  assign n1342 = ~n1338 & n1341 ;
  assign n1343 = ~n1335 & ~n1342 ;
  assign n1344 = ~n1334 & n1343 ;
  assign n1345 = x251 & ~n1082 ;
  assign n1346 = x219 & n1082 ;
  assign n1347 = ~n1345 & ~n1346 ;
  assign n1348 = x187 & ~n952 ;
  assign n1349 = x155 & n952 ;
  assign n1350 = ~n1348 & ~n1349 ;
  assign n1351 = ~n1347 & n1350 ;
  assign n1352 = n1338 & ~n1341 ;
  assign n1353 = ~n1351 & ~n1352 ;
  assign n1354 = ~n1344 & n1353 ;
  assign n1355 = x188 & ~n952 ;
  assign n1356 = x156 & n952 ;
  assign n1357 = ~n1355 & ~n1356 ;
  assign n1358 = x252 & ~n1082 ;
  assign n1359 = x220 & n1082 ;
  assign n1360 = ~n1358 & ~n1359 ;
  assign n1361 = ~n1357 & n1360 ;
  assign n1362 = n1347 & ~n1350 ;
  assign n1363 = ~n1361 & ~n1362 ;
  assign n1364 = ~n1354 & n1363 ;
  assign n1365 = n1357 & ~n1360 ;
  assign n1366 = x189 & ~n952 ;
  assign n1367 = x157 & n952 ;
  assign n1368 = ~n1366 & ~n1367 ;
  assign n1369 = x253 & ~n1082 ;
  assign n1370 = x221 & n1082 ;
  assign n1371 = ~n1369 & ~n1370 ;
  assign n1372 = n1368 & ~n1371 ;
  assign n1373 = ~n1365 & ~n1372 ;
  assign n1374 = ~n1364 & n1373 ;
  assign n1375 = ~n1368 & n1371 ;
  assign n1376 = x190 & ~n952 ;
  assign n1377 = x158 & n952 ;
  assign n1378 = ~n1376 & ~n1377 ;
  assign n1379 = x254 & ~n1082 ;
  assign n1380 = x222 & n1082 ;
  assign n1381 = ~n1379 & ~n1380 ;
  assign n1382 = ~n1378 & n1381 ;
  assign n1383 = ~n1375 & ~n1382 ;
  assign n1384 = ~n1374 & n1383 ;
  assign n1385 = n1378 & ~n1381 ;
  assign n1386 = ~n1384 & ~n1385 ;
  assign n1387 = ~n957 & ~n1386 ;
  assign n1388 = ~n956 & ~n1387 ;
  assign n1389 = ~n955 & n1388 ;
  assign n1390 = ~n1085 & ~n1388 ;
  assign n1391 = ~n1389 & ~n1390 ;
  assign n1392 = n827 & ~n1391 ;
  assign n1393 = ~n1092 & n1388 ;
  assign n1394 = ~n1089 & ~n1388 ;
  assign n1395 = ~n1393 & ~n1394 ;
  assign n1396 = ~n535 & n824 ;
  assign n1397 = ~n532 & ~n824 ;
  assign n1398 = ~n1396 & ~n1397 ;
  assign n1399 = n1395 & ~n1398 ;
  assign n1400 = ~n1392 & n1399 ;
  assign n1401 = ~n1100 & n1388 ;
  assign n1402 = ~n1097 & ~n1388 ;
  assign n1403 = ~n1401 & ~n1402 ;
  assign n1404 = ~n543 & n824 ;
  assign n1405 = ~n540 & ~n824 ;
  assign n1406 = ~n1404 & ~n1405 ;
  assign n1407 = n1403 & ~n1406 ;
  assign n1408 = ~n827 & n1391 ;
  assign n1409 = ~n1407 & ~n1408 ;
  assign n1410 = ~n1400 & n1409 ;
  assign n1411 = ~n1403 & n1406 ;
  assign n1412 = ~n550 & n824 ;
  assign n1413 = ~n553 & ~n824 ;
  assign n1414 = ~n1412 & ~n1413 ;
  assign n1415 = ~n1111 & n1388 ;
  assign n1416 = ~n1108 & ~n1388 ;
  assign n1417 = ~n1415 & ~n1416 ;
  assign n1418 = n1414 & ~n1417 ;
  assign n1419 = ~n1411 & ~n1418 ;
  assign n1420 = ~n1410 & n1419 ;
  assign n1421 = ~n1117 & n1388 ;
  assign n1422 = ~n1120 & ~n1388 ;
  assign n1423 = ~n1421 & ~n1422 ;
  assign n1424 = ~n563 & n824 ;
  assign n1425 = ~n560 & ~n824 ;
  assign n1426 = ~n1424 & ~n1425 ;
  assign n1427 = n1423 & ~n1426 ;
  assign n1428 = ~n1414 & n1417 ;
  assign n1429 = ~n1427 & ~n1428 ;
  assign n1430 = ~n1420 & n1429 ;
  assign n1431 = ~n573 & n824 ;
  assign n1432 = ~n570 & ~n824 ;
  assign n1433 = ~n1431 & ~n1432 ;
  assign n1434 = ~n1130 & n1388 ;
  assign n1435 = ~n1127 & ~n1388 ;
  assign n1436 = ~n1434 & ~n1435 ;
  assign n1437 = n1433 & ~n1436 ;
  assign n1438 = ~n1423 & n1426 ;
  assign n1439 = ~n1437 & ~n1438 ;
  assign n1440 = ~n1430 & n1439 ;
  assign n1441 = ~n580 & n824 ;
  assign n1442 = ~n583 & ~n824 ;
  assign n1443 = ~n1441 & ~n1442 ;
  assign n1444 = ~n1140 & n1388 ;
  assign n1445 = ~n1137 & ~n1388 ;
  assign n1446 = ~n1444 & ~n1445 ;
  assign n1447 = ~n1443 & n1446 ;
  assign n1448 = ~n1433 & n1436 ;
  assign n1449 = ~n1447 & ~n1448 ;
  assign n1450 = ~n1440 & n1449 ;
  assign n1451 = ~n590 & n824 ;
  assign n1452 = ~n593 & ~n824 ;
  assign n1453 = ~n1451 & ~n1452 ;
  assign n1454 = ~n1148 & n1388 ;
  assign n1455 = ~n1151 & ~n1388 ;
  assign n1456 = ~n1454 & ~n1455 ;
  assign n1457 = n1453 & ~n1456 ;
  assign n1458 = n1443 & ~n1446 ;
  assign n1459 = ~n1457 & ~n1458 ;
  assign n1460 = ~n1450 & n1459 ;
  assign n1461 = ~n1161 & n1388 ;
  assign n1462 = ~n1158 & ~n1388 ;
  assign n1463 = ~n1461 & ~n1462 ;
  assign n1464 = ~n604 & n824 ;
  assign n1465 = ~n601 & ~n824 ;
  assign n1466 = ~n1464 & ~n1465 ;
  assign n1467 = n1463 & ~n1466 ;
  assign n1468 = ~n1453 & n1456 ;
  assign n1469 = ~n1467 & ~n1468 ;
  assign n1470 = ~n1460 & n1469 ;
  assign n1471 = ~n614 & n824 ;
  assign n1472 = ~n611 & ~n824 ;
  assign n1473 = ~n1471 & ~n1472 ;
  assign n1474 = ~n1171 & n1388 ;
  assign n1475 = ~n1168 & ~n1388 ;
  assign n1476 = ~n1474 & ~n1475 ;
  assign n1477 = n1473 & ~n1476 ;
  assign n1478 = ~n1463 & n1466 ;
  assign n1479 = ~n1477 & ~n1478 ;
  assign n1480 = ~n1470 & n1479 ;
  assign n1481 = ~n1178 & n1388 ;
  assign n1482 = ~n1181 & ~n1388 ;
  assign n1483 = ~n1481 & ~n1482 ;
  assign n1484 = ~n621 & n824 ;
  assign n1485 = ~n624 & ~n824 ;
  assign n1486 = ~n1484 & ~n1485 ;
  assign n1487 = n1483 & ~n1486 ;
  assign n1488 = ~n1473 & n1476 ;
  assign n1489 = ~n1487 & ~n1488 ;
  assign n1490 = ~n1480 & n1489 ;
  assign n1491 = ~n630 & n824 ;
  assign n1492 = ~n633 & ~n824 ;
  assign n1493 = ~n1491 & ~n1492 ;
  assign n1494 = ~n1187 & n1388 ;
  assign n1495 = ~n1190 & ~n1388 ;
  assign n1496 = ~n1494 & ~n1495 ;
  assign n1497 = n1493 & ~n1496 ;
  assign n1498 = ~n1483 & n1486 ;
  assign n1499 = ~n1497 & ~n1498 ;
  assign n1500 = ~n1490 & n1499 ;
  assign n1501 = ~n1200 & n1388 ;
  assign n1502 = ~n1197 & ~n1388 ;
  assign n1503 = ~n1501 & ~n1502 ;
  assign n1504 = ~n643 & n824 ;
  assign n1505 = ~n640 & ~n824 ;
  assign n1506 = ~n1504 & ~n1505 ;
  assign n1507 = n1503 & ~n1506 ;
  assign n1508 = ~n1493 & n1496 ;
  assign n1509 = ~n1507 & ~n1508 ;
  assign n1510 = ~n1500 & n1509 ;
  assign n1511 = ~n654 & n824 ;
  assign n1512 = ~n651 & ~n824 ;
  assign n1513 = ~n1511 & ~n1512 ;
  assign n1514 = ~n1211 & n1388 ;
  assign n1515 = ~n1208 & ~n1388 ;
  assign n1516 = ~n1514 & ~n1515 ;
  assign n1517 = n1513 & ~n1516 ;
  assign n1518 = ~n1503 & n1506 ;
  assign n1519 = ~n1517 & ~n1518 ;
  assign n1520 = ~n1510 & n1519 ;
  assign n1521 = ~n1218 & n1388 ;
  assign n1522 = ~n1221 & ~n1388 ;
  assign n1523 = ~n1521 & ~n1522 ;
  assign n1524 = ~n661 & n824 ;
  assign n1525 = ~n664 & ~n824 ;
  assign n1526 = ~n1524 & ~n1525 ;
  assign n1527 = n1523 & ~n1526 ;
  assign n1528 = ~n1513 & n1516 ;
  assign n1529 = ~n1527 & ~n1528 ;
  assign n1530 = ~n1520 & n1529 ;
  assign n1531 = ~n670 & n824 ;
  assign n1532 = ~n673 & ~n824 ;
  assign n1533 = ~n1531 & ~n1532 ;
  assign n1534 = ~n1227 & n1388 ;
  assign n1535 = ~n1230 & ~n1388 ;
  assign n1536 = ~n1534 & ~n1535 ;
  assign n1537 = n1533 & ~n1536 ;
  assign n1538 = ~n1523 & n1526 ;
  assign n1539 = ~n1537 & ~n1538 ;
  assign n1540 = ~n1530 & n1539 ;
  assign n1541 = ~n1240 & n1388 ;
  assign n1542 = ~n1237 & ~n1388 ;
  assign n1543 = ~n1541 & ~n1542 ;
  assign n1544 = ~n683 & n824 ;
  assign n1545 = ~n680 & ~n824 ;
  assign n1546 = ~n1544 & ~n1545 ;
  assign n1547 = n1543 & ~n1546 ;
  assign n1548 = ~n1533 & n1536 ;
  assign n1549 = ~n1547 & ~n1548 ;
  assign n1550 = ~n1540 & n1549 ;
  assign n1551 = ~n694 & n824 ;
  assign n1552 = ~n691 & ~n824 ;
  assign n1553 = ~n1551 & ~n1552 ;
  assign n1554 = ~n1251 & n1388 ;
  assign n1555 = ~n1248 & ~n1388 ;
  assign n1556 = ~n1554 & ~n1555 ;
  assign n1557 = n1553 & ~n1556 ;
  assign n1558 = ~n1543 & n1546 ;
  assign n1559 = ~n1557 & ~n1558 ;
  assign n1560 = ~n1550 & n1559 ;
  assign n1561 = ~n1258 & n1388 ;
  assign n1562 = ~n1261 & ~n1388 ;
  assign n1563 = ~n1561 & ~n1562 ;
  assign n1564 = ~n701 & n824 ;
  assign n1565 = ~n704 & ~n824 ;
  assign n1566 = ~n1564 & ~n1565 ;
  assign n1567 = n1563 & ~n1566 ;
  assign n1568 = ~n1553 & n1556 ;
  assign n1569 = ~n1567 & ~n1568 ;
  assign n1570 = ~n1560 & n1569 ;
  assign n1571 = ~n710 & n824 ;
  assign n1572 = ~n713 & ~n824 ;
  assign n1573 = ~n1571 & ~n1572 ;
  assign n1574 = ~n1267 & n1388 ;
  assign n1575 = ~n1270 & ~n1388 ;
  assign n1576 = ~n1574 & ~n1575 ;
  assign n1577 = n1573 & ~n1576 ;
  assign n1578 = ~n1563 & n1566 ;
  assign n1579 = ~n1577 & ~n1578 ;
  assign n1580 = ~n1570 & n1579 ;
  assign n1581 = ~n1280 & n1388 ;
  assign n1582 = ~n1277 & ~n1388 ;
  assign n1583 = ~n1581 & ~n1582 ;
  assign n1584 = ~n723 & n824 ;
  assign n1585 = ~n720 & ~n824 ;
  assign n1586 = ~n1584 & ~n1585 ;
  assign n1587 = n1583 & ~n1586 ;
  assign n1588 = ~n1573 & n1576 ;
  assign n1589 = ~n1587 & ~n1588 ;
  assign n1590 = ~n1580 & n1589 ;
  assign n1591 = ~n734 & n824 ;
  assign n1592 = ~n731 & ~n824 ;
  assign n1593 = ~n1591 & ~n1592 ;
  assign n1594 = ~n1291 & n1388 ;
  assign n1595 = ~n1288 & ~n1388 ;
  assign n1596 = ~n1594 & ~n1595 ;
  assign n1597 = n1593 & ~n1596 ;
  assign n1598 = ~n1583 & n1586 ;
  assign n1599 = ~n1597 & ~n1598 ;
  assign n1600 = ~n1590 & n1599 ;
  assign n1601 = ~n1298 & n1388 ;
  assign n1602 = ~n1301 & ~n1388 ;
  assign n1603 = ~n1601 & ~n1602 ;
  assign n1604 = ~n741 & n824 ;
  assign n1605 = ~n744 & ~n824 ;
  assign n1606 = ~n1604 & ~n1605 ;
  assign n1607 = n1603 & ~n1606 ;
  assign n1608 = ~n1593 & n1596 ;
  assign n1609 = ~n1607 & ~n1608 ;
  assign n1610 = ~n1600 & n1609 ;
  assign n1611 = ~n750 & n824 ;
  assign n1612 = ~n753 & ~n824 ;
  assign n1613 = ~n1611 & ~n1612 ;
  assign n1614 = ~n1307 & n1388 ;
  assign n1615 = ~n1310 & ~n1388 ;
  assign n1616 = ~n1614 & ~n1615 ;
  assign n1617 = n1613 & ~n1616 ;
  assign n1618 = ~n1603 & n1606 ;
  assign n1619 = ~n1617 & ~n1618 ;
  assign n1620 = ~n1610 & n1619 ;
  assign n1621 = ~n760 & n824 ;
  assign n1622 = ~n763 & ~n824 ;
  assign n1623 = ~n1621 & ~n1622 ;
  assign n1624 = ~n1320 & n1388 ;
  assign n1625 = ~n1317 & ~n1388 ;
  assign n1626 = ~n1624 & ~n1625 ;
  assign n1627 = ~n1623 & n1626 ;
  assign n1628 = ~n1613 & n1616 ;
  assign n1629 = ~n1627 & ~n1628 ;
  assign n1630 = ~n1620 & n1629 ;
  assign n1631 = ~n774 & n824 ;
  assign n1632 = ~n771 & ~n824 ;
  assign n1633 = ~n1631 & ~n1632 ;
  assign n1634 = ~n1331 & n1388 ;
  assign n1635 = ~n1328 & ~n1388 ;
  assign n1636 = ~n1634 & ~n1635 ;
  assign n1637 = n1633 & ~n1636 ;
  assign n1638 = n1623 & ~n1626 ;
  assign n1639 = ~n1637 & ~n1638 ;
  assign n1640 = ~n1630 & n1639 ;
  assign n1641 = ~n1338 & n1388 ;
  assign n1642 = ~n1341 & ~n1388 ;
  assign n1643 = ~n1641 & ~n1642 ;
  assign n1644 = ~n781 & n824 ;
  assign n1645 = ~n784 & ~n824 ;
  assign n1646 = ~n1644 & ~n1645 ;
  assign n1647 = n1643 & ~n1646 ;
  assign n1648 = ~n1633 & n1636 ;
  assign n1649 = ~n1647 & ~n1648 ;
  assign n1650 = ~n1640 & n1649 ;
  assign n1651 = ~n1643 & n1646 ;
  assign n1652 = ~n790 & n824 ;
  assign n1653 = ~n793 & ~n824 ;
  assign n1654 = ~n1652 & ~n1653 ;
  assign n1655 = ~n1350 & n1388 ;
  assign n1656 = ~n1347 & ~n1388 ;
  assign n1657 = ~n1655 & ~n1656 ;
  assign n1658 = n1654 & ~n1657 ;
  assign n1659 = ~n1651 & ~n1658 ;
  assign n1660 = ~n1650 & n1659 ;
  assign n1661 = ~n1654 & n1657 ;
  assign n1662 = ~n1357 & n1388 ;
  assign n1663 = ~n1360 & ~n1388 ;
  assign n1664 = ~n1662 & ~n1663 ;
  assign n1665 = ~n803 & n824 ;
  assign n1666 = ~n800 & ~n824 ;
  assign n1667 = ~n1665 & ~n1666 ;
  assign n1668 = n1664 & ~n1667 ;
  assign n1669 = ~n1661 & ~n1668 ;
  assign n1670 = ~n1660 & n1669 ;
  assign n1671 = ~n1664 & n1667 ;
  assign n1672 = ~n1368 & n1388 ;
  assign n1673 = ~n1371 & ~n1388 ;
  assign n1674 = ~n1672 & ~n1673 ;
  assign n1675 = ~n811 & n824 ;
  assign n1676 = ~n814 & ~n824 ;
  assign n1677 = ~n1675 & ~n1676 ;
  assign n1678 = ~n1674 & n1677 ;
  assign n1679 = ~n1671 & ~n1678 ;
  assign n1680 = ~n1670 & n1679 ;
  assign n1681 = n1674 & ~n1677 ;
  assign n1682 = ~n1378 & n1388 ;
  assign n1683 = ~n1381 & ~n1388 ;
  assign n1684 = ~n1682 & ~n1683 ;
  assign n1685 = ~n524 & n824 ;
  assign n1686 = ~n521 & ~n824 ;
  assign n1687 = ~n1685 & ~n1686 ;
  assign n1688 = n1684 & ~n1687 ;
  assign n1689 = ~n1681 & ~n1688 ;
  assign n1690 = ~n1680 & n1689 ;
  assign n1691 = ~n259 & n262 ;
  assign n1692 = ~n1684 & n1687 ;
  assign n1693 = ~n1691 & ~n1692 ;
  assign n1694 = ~n1690 & n1693 ;
  assign n1695 = ~n263 & ~n1694 ;
  assign n1696 = ~n1388 & n1695 ;
  assign n1697 = ~n824 & ~n1695 ;
  assign n1698 = ~n1696 & ~n1697 ;
  assign n1699 = n952 & n1698 ;
  assign n1700 = n1082 & ~n1388 ;
  assign n1701 = ~n1699 & ~n1700 ;
  assign n1702 = n1695 & ~n1701 ;
  assign n1703 = n388 & n1698 ;
  assign n1704 = n518 & ~n824 ;
  assign n1705 = ~n1703 & ~n1704 ;
  assign n1706 = ~n1695 & ~n1705 ;
  assign n1707 = ~n1702 & ~n1706 ;
  assign n1708 = ~n1398 & ~n1695 ;
  assign n1709 = ~n1395 & n1695 ;
  assign n1710 = ~n1708 & ~n1709 ;
  assign n1711 = ~n827 & ~n1695 ;
  assign n1712 = ~n1391 & n1695 ;
  assign n1713 = ~n1711 & ~n1712 ;
  assign n1714 = ~n1406 & ~n1695 ;
  assign n1715 = ~n1403 & n1695 ;
  assign n1716 = ~n1714 & ~n1715 ;
  assign n1717 = ~n1417 & n1695 ;
  assign n1718 = ~n1414 & ~n1695 ;
  assign n1719 = ~n1717 & ~n1718 ;
  assign n1720 = ~n1426 & ~n1695 ;
  assign n1721 = ~n1423 & n1695 ;
  assign n1722 = ~n1720 & ~n1721 ;
  assign n1723 = ~n1433 & ~n1695 ;
  assign n1724 = ~n1436 & n1695 ;
  assign n1725 = ~n1723 & ~n1724 ;
  assign n1726 = ~n1446 & n1695 ;
  assign n1727 = ~n1443 & ~n1695 ;
  assign n1728 = ~n1726 & ~n1727 ;
  assign n1729 = ~n1453 & ~n1695 ;
  assign n1730 = ~n1456 & n1695 ;
  assign n1731 = ~n1729 & ~n1730 ;
  assign n1732 = ~n1466 & ~n1695 ;
  assign n1733 = ~n1463 & n1695 ;
  assign n1734 = ~n1732 & ~n1733 ;
  assign n1735 = ~n1473 & ~n1695 ;
  assign n1736 = ~n1476 & n1695 ;
  assign n1737 = ~n1735 & ~n1736 ;
  assign n1738 = n1486 & ~n1695 ;
  assign n1739 = n1483 & n1695 ;
  assign n1740 = ~n1738 & ~n1739 ;
  assign n1741 = ~n1493 & ~n1695 ;
  assign n1742 = ~n1496 & n1695 ;
  assign n1743 = ~n1741 & ~n1742 ;
  assign n1744 = ~n1506 & ~n1695 ;
  assign n1745 = ~n1503 & n1695 ;
  assign n1746 = ~n1744 & ~n1745 ;
  assign n1747 = ~n1513 & ~n1695 ;
  assign n1748 = ~n1516 & n1695 ;
  assign n1749 = ~n1747 & ~n1748 ;
  assign n1750 = n1526 & ~n1695 ;
  assign n1751 = n1523 & n1695 ;
  assign n1752 = ~n1750 & ~n1751 ;
  assign n1753 = ~n1533 & ~n1695 ;
  assign n1754 = ~n1536 & n1695 ;
  assign n1755 = ~n1753 & ~n1754 ;
  assign n1756 = ~n1546 & ~n1695 ;
  assign n1757 = ~n1543 & n1695 ;
  assign n1758 = ~n1756 & ~n1757 ;
  assign n1759 = ~n1553 & ~n1695 ;
  assign n1760 = ~n1556 & n1695 ;
  assign n1761 = ~n1759 & ~n1760 ;
  assign n1762 = n1566 & ~n1695 ;
  assign n1763 = n1563 & n1695 ;
  assign n1764 = ~n1762 & ~n1763 ;
  assign n1765 = ~n1573 & ~n1695 ;
  assign n1766 = ~n1576 & n1695 ;
  assign n1767 = ~n1765 & ~n1766 ;
  assign n1768 = ~n1586 & ~n1695 ;
  assign n1769 = ~n1583 & n1695 ;
  assign n1770 = ~n1768 & ~n1769 ;
  assign n1771 = ~n1593 & ~n1695 ;
  assign n1772 = ~n1596 & n1695 ;
  assign n1773 = ~n1771 & ~n1772 ;
  assign n1774 = n1606 & ~n1695 ;
  assign n1775 = n1603 & n1695 ;
  assign n1776 = ~n1774 & ~n1775 ;
  assign n1777 = ~n1613 & ~n1695 ;
  assign n1778 = ~n1616 & n1695 ;
  assign n1779 = ~n1777 & ~n1778 ;
  assign n1780 = ~n1626 & n1695 ;
  assign n1781 = ~n1623 & ~n1695 ;
  assign n1782 = ~n1780 & ~n1781 ;
  assign n1783 = ~n1633 & ~n1695 ;
  assign n1784 = ~n1636 & n1695 ;
  assign n1785 = ~n1783 & ~n1784 ;
  assign n1786 = n1646 & ~n1695 ;
  assign n1787 = n1643 & n1695 ;
  assign n1788 = ~n1786 & ~n1787 ;
  assign n1789 = ~n1657 & n1695 ;
  assign n1790 = ~n1654 & ~n1695 ;
  assign n1791 = ~n1789 & ~n1790 ;
  assign n1792 = ~n1667 & ~n1695 ;
  assign n1793 = ~n1664 & n1695 ;
  assign n1794 = ~n1792 & ~n1793 ;
  assign n1795 = n1677 & ~n1695 ;
  assign n1796 = n1674 & n1695 ;
  assign n1797 = ~n1795 & ~n1796 ;
  assign n1798 = ~n1687 & ~n1695 ;
  assign n1799 = ~n1684 & n1695 ;
  assign n1800 = ~n1798 & ~n1799 ;
  assign n1801 = n259 & n262 ;
  assign y0 = n1707 ;
  assign y1 = ~n1698 ;
  assign y2 = n1695 ;
  assign y3 = ~n1710 ;
  assign y4 = ~n1713 ;
  assign y5 = ~n1716 ;
  assign y6 = ~n1719 ;
  assign y7 = ~n1722 ;
  assign y8 = ~n1725 ;
  assign y9 = ~n1728 ;
  assign y10 = ~n1731 ;
  assign y11 = ~n1734 ;
  assign y12 = ~n1737 ;
  assign y13 = n1740 ;
  assign y14 = ~n1743 ;
  assign y15 = ~n1746 ;
  assign y16 = ~n1749 ;
  assign y17 = n1752 ;
  assign y18 = ~n1755 ;
  assign y19 = ~n1758 ;
  assign y20 = ~n1761 ;
  assign y21 = n1764 ;
  assign y22 = ~n1767 ;
  assign y23 = ~n1770 ;
  assign y24 = ~n1773 ;
  assign y25 = n1776 ;
  assign y26 = ~n1779 ;
  assign y27 = ~n1782 ;
  assign y28 = ~n1785 ;
  assign y29 = n1788 ;
  assign y30 = ~n1791 ;
  assign y31 = ~n1794 ;
  assign y32 = n1797 ;
  assign y33 = ~n1800 ;
  assign y34 = ~n1801 ;
endmodule
