module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 ;
  assign n31 = ~x4 & x7 ;
  assign n57 = x1 & ~x2 ;
  assign n58 = ~n31 & n57 ;
  assign n47 = x4 & x8 ;
  assign n59 = x3 & x4 ;
  assign n60 = ~n47 & ~n59 ;
  assign n61 = n58 & n60 ;
  assign n62 = ~x7 & ~x8 ;
  assign n63 = ~x1 & x2 ;
  assign n64 = n62 & n63 ;
  assign n65 = ~x9 & ~n64 ;
  assign n66 = ~n61 & n65 ;
  assign n54 = ~x5 & x6 ;
  assign n55 = x9 & ~n54 ;
  assign n67 = x5 & ~x6 ;
  assign n71 = n55 & n67 ;
  assign n72 = ~n66 & n71 ;
  assign n40 = x1 & x4 ;
  assign n41 = ~x4 & x8 ;
  assign n42 = ~n40 & ~n41 ;
  assign n43 = x0 & ~n42 ;
  assign n12 = ~x6 & ~x7 ;
  assign n44 = ~x0 & ~n40 ;
  assign n45 = n12 & ~n44 ;
  assign n46 = ~n43 & n45 ;
  assign n28 = ~x2 & ~x7 ;
  assign n29 = x1 & x5 ;
  assign n30 = n28 & n29 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = x3 & ~x8 ;
  assign n34 = n32 & n33 ;
  assign n25 = ~x3 & x4 ;
  assign n26 = x7 & ~x8 ;
  assign n27 = n25 & n26 ;
  assign n35 = n34 ^ n27 ;
  assign n36 = ~x4 & x5 ;
  assign n37 = x8 & n36 ;
  assign n48 = ~x5 & ~n47 ;
  assign n49 = ~n37 & n48 ;
  assign n50 = ~n35 & n49 ;
  assign n51 = ~n46 & n50 ;
  assign n38 = x5 & ~n37 ;
  assign n39 = ~n35 & n38 ;
  assign n52 = n51 ^ n39 ;
  assign n68 = ~x9 & n67 ;
  assign n69 = ~n66 & n68 ;
  assign n70 = n52 & n69 ;
  assign n73 = n72 ^ n70 ;
  assign n53 = ~x9 & n52 ;
  assign n56 = n55 ^ n53 ;
  assign n74 = n73 ^ n56 ;
  assign n78 = ~x10 & n74 ;
  assign n14 = ~x8 & ~x9 ;
  assign n15 = x3 ^ x2 ;
  assign n16 = n14 & n15 ;
  assign n17 = ~x10 & ~n16 ;
  assign n18 = ~x7 & ~n17 ;
  assign n19 = x8 & x10 ;
  assign n20 = x9 & n19 ;
  assign n21 = ~n18 & ~n20 ;
  assign n75 = x6 & ~x10 ;
  assign n76 = ~n21 & n75 ;
  assign n77 = n74 & n76 ;
  assign n79 = n78 ^ n77 ;
  assign n22 = x6 & x10 ;
  assign n23 = n21 & n22 ;
  assign n13 = x10 & n12 ;
  assign n24 = n23 ^ n13 ;
  assign n80 = n79 ^ n24 ;
  assign n93 = ~x4 & ~x9 ;
  assign n110 = ~n28 & ~n93 ;
  assign n111 = x8 & ~x9 ;
  assign n112 = ~x1 & ~n111 ;
  assign n113 = ~n110 & n112 ;
  assign n114 = n113 ^ n111 ;
  assign n115 = ~x0 & x2 ;
  assign n116 = x4 & ~x7 ;
  assign n117 = ~n115 & n116 ;
  assign n85 = x1 & x2 ;
  assign n121 = x0 & ~x6 ;
  assign n122 = ~n85 & n121 ;
  assign n123 = n117 & n122 ;
  assign n124 = ~n114 & n123 ;
  assign n118 = ~x6 & ~n117 ;
  assign n119 = ~n114 & n118 ;
  assign n120 = n119 ^ x6 ;
  assign n125 = n124 ^ n120 ;
  assign n81 = ~x7 & x9 ;
  assign n126 = x7 & n14 ;
  assign n127 = ~n59 & n126 ;
  assign n128 = ~n81 & ~n127 ;
  assign n129 = n125 & n128 ;
  assign n82 = ~x9 & n41 ;
  assign n83 = ~n81 & ~n82 ;
  assign n84 = ~x6 & ~n83 ;
  assign n130 = ~x5 & ~x10 ;
  assign n131 = ~n84 & n130 ;
  assign n132 = n129 & n131 ;
  assign n94 = ~n81 & ~n93 ;
  assign n101 = ~x3 & x6 ;
  assign n102 = ~n14 & n101 ;
  assign n103 = n94 & n102 ;
  assign n104 = n103 ^ x3 ;
  assign n89 = ~x4 & ~x6 ;
  assign n90 = ~x7 & n85 ;
  assign n91 = n89 & n90 ;
  assign n86 = ~x7 & ~n85 ;
  assign n87 = x4 & n14 ;
  assign n88 = ~n86 & n87 ;
  assign n92 = n91 ^ n88 ;
  assign n99 = x3 & ~n92 ;
  assign n95 = x3 & x6 ;
  assign n96 = ~n14 & n95 ;
  assign n97 = n94 & n96 ;
  assign n98 = ~n92 & n97 ;
  assign n100 = n99 ^ n98 ;
  assign n105 = n104 ^ n100 ;
  assign n106 = x5 & ~x10 ;
  assign n107 = ~n105 & n106 ;
  assign n108 = ~n84 & n107 ;
  assign n109 = n108 ^ x10 ;
  assign n133 = n132 ^ n109 ;
  assign n146 = ~x4 & x6 ;
  assign n147 = ~x9 & n146 ;
  assign n144 = ~x3 & x5 ;
  assign n145 = ~x6 & n144 ;
  assign n148 = n147 ^ n145 ;
  assign n149 = ~x2 & n148 ;
  assign n141 = x6 & ~x9 ;
  assign n142 = x2 & n59 ;
  assign n143 = n141 & n142 ;
  assign n150 = n149 ^ n143 ;
  assign n151 = ~x4 & n141 ;
  assign n155 = ~x1 & ~x3 ;
  assign n156 = n67 & n155 ;
  assign n157 = ~n151 & n156 ;
  assign n158 = ~n150 & n157 ;
  assign n152 = ~x3 & n151 ;
  assign n153 = ~n150 & n152 ;
  assign n154 = n153 ^ n150 ;
  assign n159 = n158 ^ n154 ;
  assign n134 = x6 & x7 ;
  assign n135 = ~x9 & n134 ;
  assign n136 = n19 & n135 ;
  assign n137 = ~x8 & ~n134 ;
  assign n160 = ~x7 & ~x10 ;
  assign n161 = n137 & n160 ;
  assign n162 = ~n136 & n161 ;
  assign n163 = n159 & n162 ;
  assign n138 = x10 & n137 ;
  assign n139 = ~n136 & n138 ;
  assign n140 = n139 ^ n136 ;
  assign n164 = n163 ^ n140 ;
  assign n165 = n133 & ~n164 ;
  assign n197 = x5 & x6 ;
  assign n198 = ~x8 & ~n59 ;
  assign n199 = ~n197 & n198 ;
  assign n192 = ~x1 & x5 ;
  assign n193 = ~x6 & n192 ;
  assign n178 = x2 & ~x5 ;
  assign n191 = x6 & n178 ;
  assign n194 = n193 ^ n191 ;
  assign n195 = ~x8 & n59 ;
  assign n196 = ~n194 & n195 ;
  assign n200 = n199 ^ n196 ;
  assign n175 = x0 & x1 ;
  assign n176 = n59 & ~n175 ;
  assign n177 = n176 ^ n89 ;
  assign n179 = n177 & n178 ;
  assign n205 = ~x7 & n179 ;
  assign n180 = ~x5 & n177 ;
  assign n182 = n25 & n121 ;
  assign n181 = x3 & n36 ;
  assign n183 = n182 ^ n181 ;
  assign n203 = n90 & n183 ;
  assign n204 = ~n180 & n203 ;
  assign n206 = n205 ^ n204 ;
  assign n207 = n200 & ~n206 ;
  assign n184 = n85 & n183 ;
  assign n185 = ~n180 & n184 ;
  assign n186 = n185 ^ n179 ;
  assign n187 = ~x2 & x3 ;
  assign n188 = ~x6 & n187 ;
  assign n189 = n188 ^ n144 ;
  assign n190 = n116 & n189 ;
  assign n201 = n190 & n200 ;
  assign n202 = ~n186 & n201 ;
  assign n208 = n207 ^ n202 ;
  assign n209 = n208 ^ x8 ;
  assign n166 = x4 & x5 ;
  assign n213 = x3 & ~x6 ;
  assign n214 = x7 & n213 ;
  assign n211 = ~x2 & x6 ;
  assign n212 = ~x7 & n211 ;
  assign n215 = n214 ^ n212 ;
  assign n216 = n166 & ~n215 ;
  assign n210 = ~n134 & ~n166 ;
  assign n217 = n216 ^ n210 ;
  assign n167 = x6 & ~x7 ;
  assign n168 = ~n166 & n167 ;
  assign n169 = n168 ^ x6 ;
  assign n170 = n169 ^ x7 ;
  assign n218 = ~x9 & ~x10 ;
  assign n219 = x8 & n218 ;
  assign n220 = n170 & n219 ;
  assign n221 = n220 ^ n218 ;
  assign n222 = n217 & n221 ;
  assign n223 = n209 & n222 ;
  assign n171 = x8 & n170 ;
  assign n172 = x9 & ~x10 ;
  assign n173 = ~n171 & n172 ;
  assign n174 = n173 ^ x10 ;
  assign n224 = n223 ^ n174 ;
  assign n225 = x5 & ~x8 ;
  assign n226 = x9 & n225 ;
  assign n227 = ~n19 & ~n226 ;
  assign n228 = n134 & ~n227 ;
  assign n229 = x5 & x7 ;
  assign n230 = x8 & ~n229 ;
  assign n231 = ~x10 & ~n230 ;
  assign n232 = x9 & ~n231 ;
  assign n233 = ~n228 & ~n232 ;
  assign n234 = n224 & n233 ;
  assign n235 = x7 & n197 ;
  assign n236 = ~x2 & n47 ;
  assign n237 = n235 & n236 ;
  assign n238 = ~x5 & ~x6 ;
  assign n239 = ~x4 & ~x7 ;
  assign n240 = ~x8 & n239 ;
  assign n241 = n238 & n240 ;
  assign n242 = ~n237 & ~n241 ;
  assign n243 = ~x3 & n218 ;
  assign n244 = ~n242 & n243 ;
  assign n249 = x3 & ~x7 ;
  assign n250 = n85 & n249 ;
  assign n245 = ~x5 & ~x7 ;
  assign n251 = ~n197 & ~n245 ;
  assign n252 = n250 & n251 ;
  assign n246 = x3 & n197 ;
  assign n247 = ~n245 & n246 ;
  assign n248 = n247 ^ n245 ;
  assign n253 = n252 ^ n248 ;
  assign n255 = ~x4 & ~n167 ;
  assign n256 = n253 & n255 ;
  assign n254 = ~n167 & ~n253 ;
  assign n257 = n256 ^ n254 ;
  assign n259 = n166 & n167 ;
  assign n260 = n175 & n238 ;
  assign n261 = ~n259 & ~n260 ;
  assign n262 = x2 & x3 ;
  assign n263 = ~x8 & n262 ;
  assign n264 = ~n261 & n263 ;
  assign n265 = ~n257 & n264 ;
  assign n258 = ~x8 & n257 ;
  assign n266 = n265 ^ n258 ;
  assign n267 = x7 & x8 ;
  assign n268 = n197 & n267 ;
  assign n269 = x9 & ~n268 ;
  assign n278 = ~x10 & ~n269 ;
  assign n279 = ~n266 & n278 ;
  assign n270 = n135 & n166 ;
  assign n271 = x2 & ~x3 ;
  assign n272 = x3 & x8 ;
  assign n273 = ~n271 & ~n272 ;
  assign n274 = ~x10 & ~n273 ;
  assign n275 = n270 & n274 ;
  assign n276 = ~n269 & n275 ;
  assign n277 = ~n266 & n276 ;
  assign n280 = n279 ^ n277 ;
  assign n281 = n280 ^ x10 ;
  assign n291 = x4 & n272 ;
  assign n292 = n235 & n291 ;
  assign n282 = n33 & n175 ;
  assign n283 = n245 & n282 ;
  assign n284 = n283 ^ n268 ;
  assign n285 = x2 & x4 ;
  assign n289 = n284 & n285 ;
  assign n286 = n272 & n285 ;
  assign n287 = n235 & n286 ;
  assign n288 = n284 & n287 ;
  assign n290 = n289 ^ n288 ;
  assign n293 = n292 ^ n290 ;
  assign n299 = n218 & ~n293 ;
  assign n294 = n142 & n197 ;
  assign n295 = n62 & ~n238 ;
  assign n296 = n218 & n295 ;
  assign n297 = ~n294 & n296 ;
  assign n298 = ~n293 & n297 ;
  assign n300 = n299 ^ n298 ;
  assign n301 = n62 & n218 ;
  assign n302 = ~n294 & n301 ;
  assign y0 = ~n80 ;
  assign y1 = n165 ;
  assign y2 = ~n234 ;
  assign y3 = ~n244 ;
  assign y4 = n281 ;
  assign y5 = ~n300 ;
  assign y6 = ~n302 ;
endmodule
