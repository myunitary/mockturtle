module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 ;
  assign n338 = x0 & ~x8 ;
  assign n293 = x8 ^ x0 ;
  assign n336 = x1 & ~x9 ;
  assign n337 = ~n293 & n336 ;
  assign n339 = n338 ^ n337 ;
  assign n294 = x9 ^ x1 ;
  assign n295 = n293 & n294 ;
  assign n296 = n295 ^ n293 ;
  assign n297 = n296 ^ n294 ;
  assign n333 = x2 & ~x10 ;
  assign n298 = x10 ^ x2 ;
  assign n329 = x3 & x11 ;
  assign n330 = n329 ^ x3 ;
  assign n331 = n298 & n330 ;
  assign n332 = n331 ^ n330 ;
  assign n334 = n333 ^ n332 ;
  assign n335 = ~n297 & n334 ;
  assign n340 = n339 ^ n335 ;
  assign n299 = x11 ^ x3 ;
  assign n300 = n298 & n299 ;
  assign n301 = n300 ^ n298 ;
  assign n302 = n301 ^ n299 ;
  assign n303 = ~n297 & ~n302 ;
  assign n325 = x4 & ~x12 ;
  assign n304 = x12 ^ x4 ;
  assign n323 = x5 & ~x13 ;
  assign n324 = ~n304 & n323 ;
  assign n326 = n325 ^ n324 ;
  assign n305 = x13 ^ x5 ;
  assign n306 = n304 & n305 ;
  assign n307 = n306 ^ n304 ;
  assign n308 = n307 ^ n305 ;
  assign n320 = x6 & ~x14 ;
  assign n309 = x14 ^ x6 ;
  assign n316 = x7 & x15 ;
  assign n317 = n316 ^ x7 ;
  assign n318 = n309 & n317 ;
  assign n319 = n318 ^ n317 ;
  assign n321 = n320 ^ n319 ;
  assign n322 = ~n308 & n321 ;
  assign n327 = n326 ^ n322 ;
  assign n328 = n303 & n327 ;
  assign n341 = n340 ^ n328 ;
  assign n310 = x15 ^ x7 ;
  assign n311 = n309 & n310 ;
  assign n312 = n311 ^ n309 ;
  assign n313 = n312 ^ n310 ;
  assign n314 = ~n308 & ~n313 ;
  assign n315 = n303 & n314 ;
  assign n342 = n341 ^ n315 ;
  assign n550 = x0 & ~n342 ;
  assign n344 = x8 & n342 ;
  assign n551 = n550 ^ n344 ;
  assign n345 = n344 ^ x8 ;
  assign n343 = x0 & n342 ;
  assign n346 = n345 ^ n343 ;
  assign n148 = x16 & ~x24 ;
  assign n103 = x24 ^ x16 ;
  assign n146 = x17 & ~x25 ;
  assign n147 = ~n103 & n146 ;
  assign n149 = n148 ^ n147 ;
  assign n104 = x25 ^ x17 ;
  assign n105 = n103 & n104 ;
  assign n106 = n105 ^ n103 ;
  assign n107 = n106 ^ n104 ;
  assign n143 = x18 & ~x26 ;
  assign n108 = x26 ^ x18 ;
  assign n139 = x19 & x27 ;
  assign n140 = n139 ^ x19 ;
  assign n141 = n108 & n140 ;
  assign n142 = n141 ^ n140 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = ~n107 & n144 ;
  assign n150 = n149 ^ n145 ;
  assign n109 = x27 ^ x19 ;
  assign n110 = n108 & n109 ;
  assign n111 = n110 ^ n108 ;
  assign n112 = n111 ^ n109 ;
  assign n113 = ~n107 & ~n112 ;
  assign n135 = x20 & ~x28 ;
  assign n114 = x28 ^ x20 ;
  assign n133 = x21 & ~x29 ;
  assign n134 = ~n114 & n133 ;
  assign n136 = n135 ^ n134 ;
  assign n115 = x29 ^ x21 ;
  assign n116 = n114 & n115 ;
  assign n117 = n116 ^ n114 ;
  assign n118 = n117 ^ n115 ;
  assign n130 = x22 & ~x30 ;
  assign n119 = x30 ^ x22 ;
  assign n126 = x23 & x31 ;
  assign n127 = n126 ^ x23 ;
  assign n128 = n119 & n127 ;
  assign n129 = n128 ^ n127 ;
  assign n131 = n130 ^ n129 ;
  assign n132 = ~n118 & n131 ;
  assign n137 = n136 ^ n132 ;
  assign n138 = n113 & n137 ;
  assign n151 = n150 ^ n138 ;
  assign n120 = x31 ^ x23 ;
  assign n121 = n119 & n120 ;
  assign n122 = n121 ^ n119 ;
  assign n123 = n122 ^ n120 ;
  assign n124 = ~n118 & ~n123 ;
  assign n125 = n113 & n124 ;
  assign n152 = n151 ^ n125 ;
  assign n155 = x16 & n152 ;
  assign n347 = n155 ^ x16 ;
  assign n153 = x24 & n152 ;
  assign n348 = n347 ^ n153 ;
  assign n455 = n346 & ~n348 ;
  assign n349 = n348 ^ n346 ;
  assign n351 = x9 & n342 ;
  assign n352 = n351 ^ x9 ;
  assign n350 = x1 & n342 ;
  assign n353 = n352 ^ n350 ;
  assign n164 = x17 & n152 ;
  assign n354 = n164 ^ x17 ;
  assign n162 = x25 & n152 ;
  assign n355 = n354 ^ n162 ;
  assign n453 = n353 & ~n355 ;
  assign n454 = ~n349 & n453 ;
  assign n456 = n455 ^ n454 ;
  assign n356 = n355 ^ n353 ;
  assign n357 = n349 & n356 ;
  assign n358 = n357 ^ n349 ;
  assign n359 = n358 ^ n356 ;
  assign n176 = x18 & n152 ;
  assign n360 = n176 ^ x18 ;
  assign n174 = x26 & n152 ;
  assign n361 = n360 ^ n174 ;
  assign n363 = x10 & n342 ;
  assign n364 = n363 ^ x10 ;
  assign n362 = x2 & n342 ;
  assign n365 = n364 ^ n362 ;
  assign n450 = ~n361 & n365 ;
  assign n366 = n365 ^ n361 ;
  assign n185 = x19 & n152 ;
  assign n367 = n185 ^ x19 ;
  assign n183 = x27 & n152 ;
  assign n368 = n367 ^ n183 ;
  assign n370 = x11 & n342 ;
  assign n371 = n370 ^ x11 ;
  assign n369 = x3 & n342 ;
  assign n372 = n371 ^ n369 ;
  assign n446 = n368 & n372 ;
  assign n447 = n446 ^ n372 ;
  assign n448 = n366 & n447 ;
  assign n449 = n448 ^ n447 ;
  assign n451 = n450 ^ n449 ;
  assign n452 = ~n359 & n451 ;
  assign n457 = n456 ^ n452 ;
  assign n373 = n372 ^ n368 ;
  assign n374 = n366 & n373 ;
  assign n375 = n374 ^ n366 ;
  assign n376 = n375 ^ n373 ;
  assign n377 = ~n359 & ~n376 ;
  assign n198 = x20 & n152 ;
  assign n378 = n198 ^ x20 ;
  assign n196 = x28 & n152 ;
  assign n379 = n378 ^ n196 ;
  assign n381 = x12 & n342 ;
  assign n382 = n381 ^ x12 ;
  assign n380 = x4 & n342 ;
  assign n383 = n382 ^ n380 ;
  assign n442 = ~n379 & n383 ;
  assign n384 = n383 ^ n379 ;
  assign n207 = x21 & n152 ;
  assign n385 = n207 ^ x21 ;
  assign n205 = x29 & n152 ;
  assign n386 = n385 ^ n205 ;
  assign n388 = x13 & n342 ;
  assign n389 = n388 ^ x13 ;
  assign n387 = x5 & n342 ;
  assign n390 = n389 ^ n387 ;
  assign n438 = n386 & n390 ;
  assign n439 = n438 ^ n390 ;
  assign n440 = n384 & n439 ;
  assign n441 = n440 ^ n439 ;
  assign n443 = n442 ^ n441 ;
  assign n391 = n390 ^ n386 ;
  assign n392 = n384 & n391 ;
  assign n393 = n392 ^ n384 ;
  assign n394 = n393 ^ n391 ;
  assign n219 = x22 & n152 ;
  assign n395 = n219 ^ x22 ;
  assign n217 = x30 & n152 ;
  assign n396 = n395 ^ n217 ;
  assign n398 = x14 & n342 ;
  assign n399 = n398 ^ x14 ;
  assign n397 = x6 & n342 ;
  assign n400 = n399 ^ n397 ;
  assign n434 = n396 & n400 ;
  assign n435 = n434 ^ n400 ;
  assign n401 = n400 ^ n396 ;
  assign n414 = x15 & n303 ;
  assign n415 = n327 & n414 ;
  assign n411 = x15 & n315 ;
  assign n412 = n411 ^ x15 ;
  assign n410 = x15 & n340 ;
  assign n413 = n412 ^ n410 ;
  assign n416 = n415 ^ n413 ;
  assign n407 = x7 & n303 ;
  assign n408 = n327 & n407 ;
  assign n404 = x7 & n315 ;
  assign n405 = n404 ^ x7 ;
  assign n402 = x7 & n340 ;
  assign n403 = n402 ^ x7 ;
  assign n406 = n405 ^ n403 ;
  assign n409 = n408 ^ n406 ;
  assign n417 = n416 ^ n409 ;
  assign n240 = x23 & n125 ;
  assign n241 = n240 ^ x23 ;
  assign n238 = x23 & n150 ;
  assign n421 = n241 ^ n238 ;
  assign n243 = x23 & n113 ;
  assign n244 = n137 & n243 ;
  assign n422 = n421 ^ n244 ;
  assign n248 = x31 & n150 ;
  assign n418 = n248 ^ x31 ;
  assign n246 = x31 & n125 ;
  assign n247 = n246 ^ x31 ;
  assign n419 = n418 ^ n247 ;
  assign n250 = x31 & n113 ;
  assign n251 = n137 & n250 ;
  assign n420 = n419 ^ n251 ;
  assign n423 = n422 ^ n420 ;
  assign n430 = n417 & n423 ;
  assign n431 = n430 ^ n417 ;
  assign n432 = n401 & n431 ;
  assign n433 = n432 ^ n431 ;
  assign n436 = n435 ^ n433 ;
  assign n437 = ~n394 & n436 ;
  assign n444 = n443 ^ n437 ;
  assign n445 = n377 & n444 ;
  assign n458 = n457 ^ n445 ;
  assign n424 = n423 ^ n417 ;
  assign n425 = n401 & n424 ;
  assign n426 = n425 ^ n401 ;
  assign n427 = n426 ^ n424 ;
  assign n428 = ~n394 & ~n427 ;
  assign n429 = n377 & n428 ;
  assign n459 = n458 ^ n429 ;
  assign n553 = n346 & ~n459 ;
  assign n552 = n348 & n459 ;
  assign n554 = n553 ^ n552 ;
  assign n637 = n551 & ~n554 ;
  assign n555 = n554 ^ n551 ;
  assign n556 = x1 & ~n342 ;
  assign n557 = n556 ^ n351 ;
  assign n559 = n353 & ~n459 ;
  assign n558 = n355 & n459 ;
  assign n560 = n559 ^ n558 ;
  assign n635 = n557 & ~n560 ;
  assign n636 = ~n555 & n635 ;
  assign n638 = n637 ^ n636 ;
  assign n561 = n560 ^ n557 ;
  assign n562 = ~n555 & ~n561 ;
  assign n564 = n365 & ~n459 ;
  assign n563 = n361 & n459 ;
  assign n565 = n564 ^ n563 ;
  assign n566 = x2 & ~n342 ;
  assign n567 = n566 ^ n363 ;
  assign n632 = ~n565 & n567 ;
  assign n568 = n567 ^ n565 ;
  assign n570 = n372 & ~n459 ;
  assign n569 = n368 & n459 ;
  assign n571 = n570 ^ n569 ;
  assign n572 = x3 & ~n342 ;
  assign n573 = n572 ^ n370 ;
  assign n630 = ~n571 & n573 ;
  assign n631 = ~n568 & n630 ;
  assign n633 = n632 ^ n631 ;
  assign n634 = n562 & n633 ;
  assign n639 = n638 ^ n634 ;
  assign n574 = n573 ^ n571 ;
  assign n575 = ~n568 & ~n574 ;
  assign n576 = n562 & n575 ;
  assign n578 = n383 & ~n459 ;
  assign n577 = n379 & n459 ;
  assign n579 = n578 ^ n577 ;
  assign n580 = x4 & ~n342 ;
  assign n581 = n580 ^ n381 ;
  assign n626 = ~n579 & n581 ;
  assign n582 = n581 ^ n579 ;
  assign n584 = n390 & ~n459 ;
  assign n583 = n386 & n459 ;
  assign n585 = n584 ^ n583 ;
  assign n586 = x5 & ~n342 ;
  assign n587 = n586 ^ n388 ;
  assign n624 = ~n585 & n587 ;
  assign n625 = ~n582 & n624 ;
  assign n627 = n626 ^ n625 ;
  assign n588 = n587 ^ n585 ;
  assign n589 = ~n582 & ~n588 ;
  assign n593 = x6 & ~n342 ;
  assign n594 = n593 ^ n398 ;
  assign n620 = ~n400 & n594 ;
  assign n621 = ~n459 & n620 ;
  assign n599 = x7 & ~n342 ;
  assign n598 = x15 & n342 ;
  assign n600 = n599 ^ n598 ;
  assign n609 = ~n423 & n600 ;
  assign n610 = n459 & n609 ;
  assign n607 = ~n417 & n600 ;
  assign n608 = ~n459 & n607 ;
  assign n611 = n610 ^ n608 ;
  assign n617 = n594 & n611 ;
  assign n614 = ~n400 & ~n459 ;
  assign n615 = n611 & n614 ;
  assign n612 = ~n396 & n459 ;
  assign n613 = n611 & n612 ;
  assign n616 = n615 ^ n613 ;
  assign n618 = n617 ^ n616 ;
  assign n605 = ~n396 & n594 ;
  assign n606 = n459 & n605 ;
  assign n619 = n618 ^ n606 ;
  assign n622 = n621 ^ n619 ;
  assign n623 = n589 & n622 ;
  assign n628 = n627 ^ n623 ;
  assign n629 = n576 & n628 ;
  assign n640 = n639 ^ n629 ;
  assign n591 = n400 & ~n459 ;
  assign n590 = n396 & n459 ;
  assign n592 = n591 ^ n590 ;
  assign n595 = n594 ^ n592 ;
  assign n596 = n417 & ~n459 ;
  assign n515 = n423 & n459 ;
  assign n597 = n596 ^ n515 ;
  assign n601 = n600 ^ n597 ;
  assign n602 = ~n595 & ~n601 ;
  assign n603 = n589 & n602 ;
  assign n604 = n576 & n603 ;
  assign n641 = n640 ^ n604 ;
  assign n732 = n551 & ~n641 ;
  assign n731 = n554 & n641 ;
  assign n733 = n732 ^ n731 ;
  assign n643 = n554 & ~n641 ;
  assign n642 = n551 & n641 ;
  assign n644 = n643 ^ n642 ;
  assign n461 = n348 & ~n459 ;
  assign n460 = n346 & n459 ;
  assign n462 = n461 ^ n460 ;
  assign n154 = n153 ^ x24 ;
  assign n156 = n155 ^ n154 ;
  assign n94 = x32 & ~x40 ;
  assign n49 = x40 ^ x32 ;
  assign n92 = x33 & ~x41 ;
  assign n93 = ~n49 & n92 ;
  assign n95 = n94 ^ n93 ;
  assign n50 = x41 ^ x33 ;
  assign n51 = n49 & n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n52 ^ n50 ;
  assign n89 = x34 & ~x42 ;
  assign n54 = x42 ^ x34 ;
  assign n85 = x35 & x43 ;
  assign n86 = n85 ^ x35 ;
  assign n87 = n54 & n86 ;
  assign n88 = n87 ^ n86 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = ~n53 & n90 ;
  assign n96 = n95 ^ n91 ;
  assign n55 = x43 ^ x35 ;
  assign n56 = n54 & n55 ;
  assign n57 = n56 ^ n54 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = ~n53 & ~n58 ;
  assign n81 = x36 & ~x44 ;
  assign n60 = x44 ^ x36 ;
  assign n79 = x37 & ~x45 ;
  assign n80 = ~n60 & n79 ;
  assign n82 = n81 ^ n80 ;
  assign n61 = x45 ^ x37 ;
  assign n62 = n60 & n61 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = n63 ^ n61 ;
  assign n76 = x38 & ~x46 ;
  assign n65 = x46 ^ x38 ;
  assign n72 = x39 & x47 ;
  assign n73 = n72 ^ x39 ;
  assign n74 = n65 & n73 ;
  assign n75 = n74 ^ n73 ;
  assign n77 = n76 ^ n75 ;
  assign n78 = ~n64 & n77 ;
  assign n83 = n82 ^ n78 ;
  assign n84 = n59 & n83 ;
  assign n97 = n96 ^ n84 ;
  assign n66 = x47 ^ x39 ;
  assign n67 = n65 & n66 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = n68 ^ n66 ;
  assign n70 = ~n64 & ~n69 ;
  assign n71 = n59 & n70 ;
  assign n98 = n97 ^ n71 ;
  assign n100 = x32 & n98 ;
  assign n101 = n100 ^ x32 ;
  assign n99 = x40 & n98 ;
  assign n102 = n101 ^ n99 ;
  assign n285 = ~n102 & n156 ;
  assign n157 = n156 ^ n102 ;
  assign n159 = x33 & n98 ;
  assign n160 = n159 ^ x33 ;
  assign n158 = x41 & n98 ;
  assign n161 = n160 ^ n158 ;
  assign n163 = n162 ^ x25 ;
  assign n165 = n164 ^ n163 ;
  assign n283 = ~n161 & n165 ;
  assign n284 = ~n157 & n283 ;
  assign n286 = n285 ^ n284 ;
  assign n166 = n165 ^ n161 ;
  assign n167 = n157 & n166 ;
  assign n168 = n167 ^ n157 ;
  assign n169 = n168 ^ n166 ;
  assign n171 = x34 & n98 ;
  assign n172 = n171 ^ x34 ;
  assign n170 = x42 & n98 ;
  assign n173 = n172 ^ n170 ;
  assign n175 = n174 ^ x26 ;
  assign n177 = n176 ^ n175 ;
  assign n280 = ~n173 & n177 ;
  assign n178 = n177 ^ n173 ;
  assign n180 = x35 & n98 ;
  assign n181 = n180 ^ x35 ;
  assign n179 = x43 & n98 ;
  assign n182 = n181 ^ n179 ;
  assign n184 = n183 ^ x27 ;
  assign n186 = n185 ^ n184 ;
  assign n276 = n182 & n186 ;
  assign n277 = n276 ^ n186 ;
  assign n278 = n178 & n277 ;
  assign n279 = n278 ^ n277 ;
  assign n281 = n280 ^ n279 ;
  assign n282 = ~n169 & n281 ;
  assign n287 = n286 ^ n282 ;
  assign n187 = n186 ^ n182 ;
  assign n188 = n178 & n187 ;
  assign n189 = n188 ^ n178 ;
  assign n190 = n189 ^ n187 ;
  assign n191 = ~n169 & ~n190 ;
  assign n193 = x36 & n98 ;
  assign n194 = n193 ^ x36 ;
  assign n192 = x44 & n98 ;
  assign n195 = n194 ^ n192 ;
  assign n197 = n196 ^ x28 ;
  assign n199 = n198 ^ n197 ;
  assign n272 = ~n195 & n199 ;
  assign n200 = n199 ^ n195 ;
  assign n202 = x37 & n98 ;
  assign n203 = n202 ^ x37 ;
  assign n201 = x45 & n98 ;
  assign n204 = n203 ^ n201 ;
  assign n206 = n205 ^ x29 ;
  assign n208 = n207 ^ n206 ;
  assign n268 = n204 & n208 ;
  assign n269 = n268 ^ n208 ;
  assign n270 = n200 & n269 ;
  assign n271 = n270 ^ n269 ;
  assign n273 = n272 ^ n271 ;
  assign n209 = n208 ^ n204 ;
  assign n210 = n200 & n209 ;
  assign n211 = n210 ^ n200 ;
  assign n212 = n211 ^ n209 ;
  assign n214 = x38 & n98 ;
  assign n215 = n214 ^ x38 ;
  assign n213 = x46 & n98 ;
  assign n216 = n215 ^ n213 ;
  assign n218 = n217 ^ x30 ;
  assign n220 = n219 ^ n218 ;
  assign n264 = n216 & n220 ;
  assign n265 = n264 ^ n220 ;
  assign n221 = n220 ^ n216 ;
  assign n234 = x39 & n59 ;
  assign n235 = n83 & n234 ;
  assign n231 = x39 & n71 ;
  assign n232 = n231 ^ x39 ;
  assign n230 = x39 & n96 ;
  assign n233 = n232 ^ n230 ;
  assign n236 = n235 ^ n233 ;
  assign n227 = x47 & n59 ;
  assign n228 = n83 & n227 ;
  assign n224 = x47 & n71 ;
  assign n225 = n224 ^ x47 ;
  assign n222 = x47 & n96 ;
  assign n223 = n222 ^ x47 ;
  assign n226 = n225 ^ n223 ;
  assign n229 = n228 ^ n226 ;
  assign n237 = n236 ^ n229 ;
  assign n249 = n248 ^ n247 ;
  assign n252 = n251 ^ n249 ;
  assign n239 = n238 ^ x23 ;
  assign n242 = n241 ^ n239 ;
  assign n245 = n244 ^ n242 ;
  assign n253 = n252 ^ n245 ;
  assign n260 = n237 & n253 ;
  assign n261 = n260 ^ n253 ;
  assign n262 = n221 & n261 ;
  assign n263 = n262 ^ n261 ;
  assign n266 = n265 ^ n263 ;
  assign n267 = ~n212 & n266 ;
  assign n274 = n273 ^ n267 ;
  assign n275 = n191 & n274 ;
  assign n288 = n287 ^ n275 ;
  assign n254 = n253 ^ n237 ;
  assign n255 = n221 & n254 ;
  assign n256 = n255 ^ n221 ;
  assign n257 = n256 ^ n254 ;
  assign n258 = ~n212 & ~n257 ;
  assign n259 = n191 & n258 ;
  assign n289 = n288 ^ n259 ;
  assign n291 = n156 & ~n289 ;
  assign n290 = n102 & n289 ;
  assign n292 = n291 ^ n290 ;
  assign n542 = ~n292 & n462 ;
  assign n463 = n462 ^ n292 ;
  assign n465 = n165 & ~n289 ;
  assign n464 = n161 & n289 ;
  assign n466 = n465 ^ n464 ;
  assign n468 = n355 & ~n459 ;
  assign n467 = n353 & n459 ;
  assign n469 = n468 ^ n467 ;
  assign n540 = ~n466 & n469 ;
  assign n541 = ~n463 & n540 ;
  assign n543 = n542 ^ n541 ;
  assign n470 = n469 ^ n466 ;
  assign n471 = ~n463 & ~n470 ;
  assign n473 = n177 & ~n289 ;
  assign n472 = n173 & n289 ;
  assign n474 = n473 ^ n472 ;
  assign n476 = n361 & ~n459 ;
  assign n475 = n365 & n459 ;
  assign n477 = n476 ^ n475 ;
  assign n537 = ~n474 & n477 ;
  assign n478 = n477 ^ n474 ;
  assign n480 = n186 & ~n289 ;
  assign n479 = n182 & n289 ;
  assign n481 = n480 ^ n479 ;
  assign n483 = n368 & ~n459 ;
  assign n482 = n372 & n459 ;
  assign n484 = n483 ^ n482 ;
  assign n535 = ~n481 & n484 ;
  assign n536 = ~n478 & n535 ;
  assign n538 = n537 ^ n536 ;
  assign n539 = n471 & n538 ;
  assign n544 = n543 ^ n539 ;
  assign n485 = n484 ^ n481 ;
  assign n486 = ~n478 & ~n485 ;
  assign n487 = n471 & n486 ;
  assign n489 = n199 & ~n289 ;
  assign n488 = n195 & n289 ;
  assign n490 = n489 ^ n488 ;
  assign n492 = n379 & ~n459 ;
  assign n491 = n383 & n459 ;
  assign n493 = n492 ^ n491 ;
  assign n531 = ~n490 & n493 ;
  assign n494 = n493 ^ n490 ;
  assign n496 = n208 & ~n289 ;
  assign n495 = n204 & n289 ;
  assign n497 = n496 ^ n495 ;
  assign n499 = n386 & ~n459 ;
  assign n498 = n390 & n459 ;
  assign n500 = n499 ^ n498 ;
  assign n529 = ~n497 & n500 ;
  assign n530 = ~n494 & n529 ;
  assign n532 = n531 ^ n530 ;
  assign n501 = n500 ^ n497 ;
  assign n502 = ~n494 & ~n501 ;
  assign n504 = n220 & ~n289 ;
  assign n503 = n216 & n289 ;
  assign n505 = n504 ^ n503 ;
  assign n507 = n396 & ~n459 ;
  assign n506 = n400 & n459 ;
  assign n508 = n507 ^ n506 ;
  assign n526 = ~n505 & n508 ;
  assign n509 = n508 ^ n505 ;
  assign n511 = n253 & n289 ;
  assign n512 = n511 ^ n253 ;
  assign n510 = n237 & n289 ;
  assign n513 = n512 ^ n510 ;
  assign n516 = n515 ^ n423 ;
  assign n514 = n417 & n459 ;
  assign n517 = n516 ^ n514 ;
  assign n522 = n513 & n517 ;
  assign n523 = n522 ^ n517 ;
  assign n524 = n509 & n523 ;
  assign n525 = n524 ^ n523 ;
  assign n527 = n526 ^ n525 ;
  assign n528 = n502 & n527 ;
  assign n533 = n532 ^ n528 ;
  assign n534 = n487 & n533 ;
  assign n545 = n544 ^ n534 ;
  assign n518 = n517 ^ n513 ;
  assign n519 = ~n509 & ~n518 ;
  assign n520 = n502 & n519 ;
  assign n521 = n487 & n520 ;
  assign n546 = n545 ^ n521 ;
  assign n548 = n462 & ~n546 ;
  assign n547 = n292 & n546 ;
  assign n549 = n548 ^ n547 ;
  assign n723 = ~n549 & n644 ;
  assign n645 = n644 ^ n549 ;
  assign n647 = n469 & ~n546 ;
  assign n646 = n466 & n546 ;
  assign n648 = n647 ^ n646 ;
  assign n650 = n560 & ~n641 ;
  assign n649 = n557 & n641 ;
  assign n651 = n650 ^ n649 ;
  assign n721 = ~n648 & n651 ;
  assign n722 = ~n645 & n721 ;
  assign n724 = n723 ^ n722 ;
  assign n652 = n651 ^ n648 ;
  assign n653 = ~n645 & ~n652 ;
  assign n655 = n477 & ~n546 ;
  assign n654 = n474 & n546 ;
  assign n656 = n655 ^ n654 ;
  assign n658 = n565 & ~n641 ;
  assign n657 = n567 & n641 ;
  assign n659 = n658 ^ n657 ;
  assign n718 = ~n656 & n659 ;
  assign n660 = n659 ^ n656 ;
  assign n662 = n484 & ~n546 ;
  assign n661 = n481 & n546 ;
  assign n663 = n662 ^ n661 ;
  assign n665 = n571 & ~n641 ;
  assign n664 = n573 & n641 ;
  assign n666 = n665 ^ n664 ;
  assign n716 = ~n663 & n666 ;
  assign n717 = ~n660 & n716 ;
  assign n719 = n718 ^ n717 ;
  assign n720 = n653 & n719 ;
  assign n725 = n724 ^ n720 ;
  assign n667 = n666 ^ n663 ;
  assign n668 = ~n660 & ~n667 ;
  assign n669 = n653 & n668 ;
  assign n671 = n493 & ~n546 ;
  assign n670 = n490 & n546 ;
  assign n672 = n671 ^ n670 ;
  assign n674 = n579 & ~n641 ;
  assign n673 = n581 & n641 ;
  assign n675 = n674 ^ n673 ;
  assign n712 = ~n672 & n675 ;
  assign n676 = n675 ^ n672 ;
  assign n678 = n500 & ~n546 ;
  assign n677 = n497 & n546 ;
  assign n679 = n678 ^ n677 ;
  assign n681 = n585 & ~n641 ;
  assign n680 = n587 & n641 ;
  assign n682 = n681 ^ n680 ;
  assign n710 = ~n679 & n682 ;
  assign n711 = ~n676 & n710 ;
  assign n713 = n712 ^ n711 ;
  assign n683 = n682 ^ n679 ;
  assign n684 = ~n676 & ~n683 ;
  assign n686 = n508 & ~n546 ;
  assign n685 = n505 & n546 ;
  assign n687 = n686 ^ n685 ;
  assign n689 = n592 & ~n641 ;
  assign n688 = n594 & n641 ;
  assign n690 = n689 ^ n688 ;
  assign n707 = ~n687 & n690 ;
  assign n691 = n690 ^ n687 ;
  assign n693 = n517 & n546 ;
  assign n694 = n693 ^ n517 ;
  assign n692 = n513 & n546 ;
  assign n695 = n694 ^ n692 ;
  assign n697 = n597 & ~n641 ;
  assign n696 = n600 & n641 ;
  assign n698 = n697 ^ n696 ;
  assign n703 = n695 & n698 ;
  assign n704 = n703 ^ n698 ;
  assign n705 = n691 & n704 ;
  assign n706 = n705 ^ n704 ;
  assign n708 = n707 ^ n706 ;
  assign n709 = n684 & n708 ;
  assign n714 = n713 ^ n709 ;
  assign n715 = n669 & n714 ;
  assign n726 = n725 ^ n715 ;
  assign n699 = n698 ^ n695 ;
  assign n700 = ~n691 & ~n699 ;
  assign n701 = n684 & n700 ;
  assign n702 = n669 & n701 ;
  assign n727 = n726 ^ n702 ;
  assign n729 = n644 & ~n727 ;
  assign n728 = n549 & n727 ;
  assign n730 = n729 ^ n728 ;
  assign n823 = ~n730 & n733 ;
  assign n734 = n733 ^ n730 ;
  assign n736 = n651 & ~n727 ;
  assign n735 = n648 & n727 ;
  assign n737 = n736 ^ n735 ;
  assign n739 = n557 & ~n641 ;
  assign n738 = n560 & n641 ;
  assign n740 = n739 ^ n738 ;
  assign n821 = ~n737 & n740 ;
  assign n822 = ~n734 & n821 ;
  assign n824 = n823 ^ n822 ;
  assign n741 = n740 ^ n737 ;
  assign n742 = ~n734 & ~n741 ;
  assign n744 = n659 & ~n727 ;
  assign n743 = n656 & n727 ;
  assign n745 = n744 ^ n743 ;
  assign n747 = n567 & ~n641 ;
  assign n746 = n565 & n641 ;
  assign n748 = n747 ^ n746 ;
  assign n818 = ~n745 & n748 ;
  assign n749 = n748 ^ n745 ;
  assign n751 = n666 & ~n727 ;
  assign n750 = n663 & n727 ;
  assign n752 = n751 ^ n750 ;
  assign n754 = n573 & ~n641 ;
  assign n753 = n571 & n641 ;
  assign n755 = n754 ^ n753 ;
  assign n816 = ~n752 & n755 ;
  assign n817 = ~n749 & n816 ;
  assign n819 = n818 ^ n817 ;
  assign n820 = n742 & n819 ;
  assign n825 = n824 ^ n820 ;
  assign n756 = n755 ^ n752 ;
  assign n757 = ~n749 & ~n756 ;
  assign n758 = n742 & n757 ;
  assign n760 = n675 & ~n727 ;
  assign n759 = n672 & n727 ;
  assign n761 = n760 ^ n759 ;
  assign n763 = n581 & ~n641 ;
  assign n762 = n579 & n641 ;
  assign n764 = n763 ^ n762 ;
  assign n812 = ~n761 & n764 ;
  assign n765 = n764 ^ n761 ;
  assign n767 = n682 & ~n727 ;
  assign n766 = n679 & n727 ;
  assign n768 = n767 ^ n766 ;
  assign n770 = n587 & ~n641 ;
  assign n769 = n585 & n641 ;
  assign n771 = n770 ^ n769 ;
  assign n810 = ~n768 & n771 ;
  assign n811 = ~n765 & n810 ;
  assign n813 = n812 ^ n811 ;
  assign n772 = n771 ^ n768 ;
  assign n773 = ~n765 & ~n772 ;
  assign n778 = n594 & ~n641 ;
  assign n777 = n592 & n641 ;
  assign n779 = n778 ^ n777 ;
  assign n806 = ~n690 & n779 ;
  assign n807 = ~n727 & n806 ;
  assign n785 = n600 & ~n641 ;
  assign n784 = n597 & n641 ;
  assign n786 = n785 ^ n784 ;
  assign n795 = ~n698 & n786 ;
  assign n796 = ~n727 & n795 ;
  assign n793 = ~n695 & n786 ;
  assign n794 = n727 & n793 ;
  assign n797 = n796 ^ n794 ;
  assign n803 = n779 & n797 ;
  assign n800 = ~n690 & ~n727 ;
  assign n801 = n797 & n800 ;
  assign n798 = ~n687 & n727 ;
  assign n799 = n797 & n798 ;
  assign n802 = n801 ^ n799 ;
  assign n804 = n803 ^ n802 ;
  assign n791 = ~n687 & n779 ;
  assign n792 = n727 & n791 ;
  assign n805 = n804 ^ n792 ;
  assign n808 = n807 ^ n805 ;
  assign n809 = n773 & n808 ;
  assign n814 = n813 ^ n809 ;
  assign n815 = n758 & n814 ;
  assign n826 = n825 ^ n815 ;
  assign n775 = n690 & ~n727 ;
  assign n774 = n687 & n727 ;
  assign n776 = n775 ^ n774 ;
  assign n780 = n779 ^ n776 ;
  assign n782 = n698 & ~n727 ;
  assign n781 = n695 & n727 ;
  assign n783 = n782 ^ n781 ;
  assign n787 = n786 ^ n783 ;
  assign n788 = ~n780 & ~n787 ;
  assign n789 = n773 & n788 ;
  assign n790 = n758 & n789 ;
  assign n827 = n826 ^ n790 ;
  assign n829 = n733 & ~n827 ;
  assign n828 = n730 & n827 ;
  assign n830 = n829 ^ n828 ;
  assign n832 = n740 & ~n827 ;
  assign n831 = n737 & n827 ;
  assign n833 = n832 ^ n831 ;
  assign n835 = n748 & ~n827 ;
  assign n834 = n745 & n827 ;
  assign n836 = n835 ^ n834 ;
  assign n838 = n755 & ~n827 ;
  assign n837 = n752 & n827 ;
  assign n839 = n838 ^ n837 ;
  assign n841 = n764 & ~n827 ;
  assign n840 = n761 & n827 ;
  assign n842 = n841 ^ n840 ;
  assign n844 = n771 & ~n827 ;
  assign n843 = n768 & n827 ;
  assign n845 = n844 ^ n843 ;
  assign n847 = n779 & ~n827 ;
  assign n846 = n776 & n827 ;
  assign n848 = n847 ^ n846 ;
  assign n850 = n786 & ~n827 ;
  assign n849 = n783 & n827 ;
  assign n851 = n850 ^ n849 ;
  assign n853 = n730 & ~n827 ;
  assign n852 = n733 & n827 ;
  assign n854 = n853 ^ n852 ;
  assign n856 = n737 & ~n827 ;
  assign n855 = n740 & n827 ;
  assign n857 = n856 ^ n855 ;
  assign n859 = n745 & ~n827 ;
  assign n858 = n748 & n827 ;
  assign n860 = n859 ^ n858 ;
  assign n862 = n752 & ~n827 ;
  assign n861 = n755 & n827 ;
  assign n863 = n862 ^ n861 ;
  assign n865 = n761 & ~n827 ;
  assign n864 = n764 & n827 ;
  assign n866 = n865 ^ n864 ;
  assign n868 = n768 & ~n827 ;
  assign n867 = n771 & n827 ;
  assign n869 = n868 ^ n867 ;
  assign n871 = n776 & ~n827 ;
  assign n870 = n779 & n827 ;
  assign n872 = n871 ^ n870 ;
  assign n874 = n783 & ~n827 ;
  assign n873 = n786 & n827 ;
  assign n875 = n874 ^ n873 ;
  assign n1053 = n549 & ~n727 ;
  assign n1052 = n644 & n727 ;
  assign n1054 = n1053 ^ n1052 ;
  assign n966 = n292 & ~n546 ;
  assign n965 = n462 & n546 ;
  assign n967 = n966 ^ n965 ;
  assign n879 = n102 & ~n289 ;
  assign n878 = n156 & n289 ;
  assign n880 = n879 ^ n878 ;
  assign n876 = x40 & ~n98 ;
  assign n877 = n876 ^ n100 ;
  assign n957 = ~n877 & n880 ;
  assign n881 = n880 ^ n877 ;
  assign n882 = x41 & ~n98 ;
  assign n883 = n882 ^ n159 ;
  assign n885 = n161 & ~n289 ;
  assign n884 = n165 & n289 ;
  assign n886 = n885 ^ n884 ;
  assign n955 = ~n883 & n886 ;
  assign n956 = ~n881 & n955 ;
  assign n958 = n957 ^ n956 ;
  assign n887 = n886 ^ n883 ;
  assign n888 = ~n881 & ~n887 ;
  assign n889 = x42 & ~n98 ;
  assign n890 = n889 ^ n171 ;
  assign n892 = n173 & ~n289 ;
  assign n891 = n177 & n289 ;
  assign n893 = n892 ^ n891 ;
  assign n952 = ~n890 & n893 ;
  assign n894 = n893 ^ n890 ;
  assign n895 = x43 & ~n98 ;
  assign n896 = n895 ^ n180 ;
  assign n898 = n182 & ~n289 ;
  assign n897 = n186 & n289 ;
  assign n899 = n898 ^ n897 ;
  assign n950 = ~n896 & n899 ;
  assign n951 = ~n894 & n950 ;
  assign n953 = n952 ^ n951 ;
  assign n954 = n888 & n953 ;
  assign n959 = n958 ^ n954 ;
  assign n900 = n899 ^ n896 ;
  assign n901 = ~n894 & ~n900 ;
  assign n902 = n888 & n901 ;
  assign n903 = x44 & ~n98 ;
  assign n904 = n903 ^ n193 ;
  assign n906 = n195 & ~n289 ;
  assign n905 = n199 & n289 ;
  assign n907 = n906 ^ n905 ;
  assign n946 = ~n904 & n907 ;
  assign n908 = n907 ^ n904 ;
  assign n909 = x45 & ~n98 ;
  assign n910 = n909 ^ n202 ;
  assign n912 = n204 & ~n289 ;
  assign n911 = n208 & n289 ;
  assign n913 = n912 ^ n911 ;
  assign n944 = ~n910 & n913 ;
  assign n945 = ~n908 & n944 ;
  assign n947 = n946 ^ n945 ;
  assign n914 = n913 ^ n910 ;
  assign n915 = ~n908 & ~n914 ;
  assign n916 = x46 & ~n98 ;
  assign n917 = n916 ^ n214 ;
  assign n919 = n216 & ~n289 ;
  assign n918 = n220 & n289 ;
  assign n920 = n919 ^ n918 ;
  assign n941 = ~n917 & n920 ;
  assign n925 = x47 & ~n98 ;
  assign n924 = x39 & n98 ;
  assign n926 = n925 ^ n924 ;
  assign n933 = n253 & ~n926 ;
  assign n934 = n289 & n933 ;
  assign n931 = n237 & ~n926 ;
  assign n932 = ~n289 & n931 ;
  assign n935 = n934 ^ n932 ;
  assign n939 = ~n917 & n935 ;
  assign n937 = n919 & n935 ;
  assign n936 = n918 & n935 ;
  assign n938 = n937 ^ n936 ;
  assign n940 = n939 ^ n938 ;
  assign n942 = n941 ^ n940 ;
  assign n943 = n915 & n942 ;
  assign n948 = n947 ^ n943 ;
  assign n949 = n902 & n948 ;
  assign n960 = n959 ^ n949 ;
  assign n921 = n920 ^ n917 ;
  assign n922 = n237 & ~n289 ;
  assign n923 = n922 ^ n511 ;
  assign n927 = n926 ^ n923 ;
  assign n928 = ~n921 & ~n927 ;
  assign n929 = n915 & n928 ;
  assign n930 = n902 & n929 ;
  assign n961 = n960 ^ n930 ;
  assign n963 = n880 & ~n961 ;
  assign n962 = n877 & n961 ;
  assign n964 = n963 ^ n962 ;
  assign n1044 = ~n964 & n967 ;
  assign n968 = n967 ^ n964 ;
  assign n970 = n886 & ~n961 ;
  assign n969 = n883 & n961 ;
  assign n971 = n970 ^ n969 ;
  assign n973 = n466 & ~n546 ;
  assign n972 = n469 & n546 ;
  assign n974 = n973 ^ n972 ;
  assign n1042 = ~n971 & n974 ;
  assign n1043 = ~n968 & n1042 ;
  assign n1045 = n1044 ^ n1043 ;
  assign n975 = n974 ^ n971 ;
  assign n976 = ~n968 & ~n975 ;
  assign n978 = n893 & ~n961 ;
  assign n977 = n890 & n961 ;
  assign n979 = n978 ^ n977 ;
  assign n981 = n474 & ~n546 ;
  assign n980 = n477 & n546 ;
  assign n982 = n981 ^ n980 ;
  assign n1039 = ~n979 & n982 ;
  assign n983 = n982 ^ n979 ;
  assign n985 = n899 & ~n961 ;
  assign n984 = n896 & n961 ;
  assign n986 = n985 ^ n984 ;
  assign n988 = n481 & ~n546 ;
  assign n987 = n484 & n546 ;
  assign n989 = n988 ^ n987 ;
  assign n1037 = ~n986 & n989 ;
  assign n1038 = ~n983 & n1037 ;
  assign n1040 = n1039 ^ n1038 ;
  assign n1041 = n976 & n1040 ;
  assign n1046 = n1045 ^ n1041 ;
  assign n990 = n989 ^ n986 ;
  assign n991 = ~n983 & ~n990 ;
  assign n992 = n976 & n991 ;
  assign n994 = n907 & ~n961 ;
  assign n993 = n904 & n961 ;
  assign n995 = n994 ^ n993 ;
  assign n997 = n490 & ~n546 ;
  assign n996 = n493 & n546 ;
  assign n998 = n997 ^ n996 ;
  assign n1033 = ~n995 & n998 ;
  assign n999 = n998 ^ n995 ;
  assign n1001 = n913 & ~n961 ;
  assign n1000 = n910 & n961 ;
  assign n1002 = n1001 ^ n1000 ;
  assign n1004 = n497 & ~n546 ;
  assign n1003 = n500 & n546 ;
  assign n1005 = n1004 ^ n1003 ;
  assign n1031 = ~n1002 & n1005 ;
  assign n1032 = ~n999 & n1031 ;
  assign n1034 = n1033 ^ n1032 ;
  assign n1006 = n1005 ^ n1002 ;
  assign n1007 = ~n999 & ~n1006 ;
  assign n1009 = n920 & ~n961 ;
  assign n1008 = n917 & n961 ;
  assign n1010 = n1009 ^ n1008 ;
  assign n1012 = n505 & ~n546 ;
  assign n1011 = n508 & n546 ;
  assign n1013 = n1012 ^ n1011 ;
  assign n1028 = ~n1010 & n1013 ;
  assign n1014 = n1013 ^ n1010 ;
  assign n1016 = n923 & ~n961 ;
  assign n1015 = n926 & n961 ;
  assign n1017 = n1016 ^ n1015 ;
  assign n1018 = n692 ^ n513 ;
  assign n1019 = n1018 ^ n693 ;
  assign n1024 = n1017 & n1019 ;
  assign n1025 = n1024 ^ n1019 ;
  assign n1026 = n1014 & n1025 ;
  assign n1027 = n1026 ^ n1025 ;
  assign n1029 = n1028 ^ n1027 ;
  assign n1030 = n1007 & n1029 ;
  assign n1035 = n1034 ^ n1030 ;
  assign n1036 = n992 & n1035 ;
  assign n1047 = n1046 ^ n1036 ;
  assign n1020 = n1019 ^ n1017 ;
  assign n1021 = ~n1014 & ~n1020 ;
  assign n1022 = n1007 & n1021 ;
  assign n1023 = n992 & n1022 ;
  assign n1048 = n1047 ^ n1023 ;
  assign n1050 = n967 & ~n1048 ;
  assign n1049 = n964 & n1048 ;
  assign n1051 = n1050 ^ n1049 ;
  assign n1133 = ~n1051 & n1054 ;
  assign n1055 = n1054 ^ n1051 ;
  assign n1057 = n974 & ~n1048 ;
  assign n1056 = n971 & n1048 ;
  assign n1058 = n1057 ^ n1056 ;
  assign n1060 = n648 & ~n727 ;
  assign n1059 = n651 & n727 ;
  assign n1061 = n1060 ^ n1059 ;
  assign n1131 = ~n1058 & n1061 ;
  assign n1132 = ~n1055 & n1131 ;
  assign n1134 = n1133 ^ n1132 ;
  assign n1062 = n1061 ^ n1058 ;
  assign n1063 = ~n1055 & ~n1062 ;
  assign n1065 = n982 & ~n1048 ;
  assign n1064 = n979 & n1048 ;
  assign n1066 = n1065 ^ n1064 ;
  assign n1068 = n656 & ~n727 ;
  assign n1067 = n659 & n727 ;
  assign n1069 = n1068 ^ n1067 ;
  assign n1128 = ~n1066 & n1069 ;
  assign n1070 = n1069 ^ n1066 ;
  assign n1072 = n989 & ~n1048 ;
  assign n1071 = n986 & n1048 ;
  assign n1073 = n1072 ^ n1071 ;
  assign n1075 = n663 & ~n727 ;
  assign n1074 = n666 & n727 ;
  assign n1076 = n1075 ^ n1074 ;
  assign n1126 = ~n1073 & n1076 ;
  assign n1127 = ~n1070 & n1126 ;
  assign n1129 = n1128 ^ n1127 ;
  assign n1130 = n1063 & n1129 ;
  assign n1135 = n1134 ^ n1130 ;
  assign n1077 = n1076 ^ n1073 ;
  assign n1078 = ~n1070 & ~n1077 ;
  assign n1079 = n1063 & n1078 ;
  assign n1081 = n998 & ~n1048 ;
  assign n1080 = n995 & n1048 ;
  assign n1082 = n1081 ^ n1080 ;
  assign n1084 = n672 & ~n727 ;
  assign n1083 = n675 & n727 ;
  assign n1085 = n1084 ^ n1083 ;
  assign n1122 = ~n1082 & n1085 ;
  assign n1086 = n1085 ^ n1082 ;
  assign n1088 = n1005 & ~n1048 ;
  assign n1087 = n1002 & n1048 ;
  assign n1089 = n1088 ^ n1087 ;
  assign n1091 = n679 & ~n727 ;
  assign n1090 = n682 & n727 ;
  assign n1092 = n1091 ^ n1090 ;
  assign n1120 = ~n1089 & n1092 ;
  assign n1121 = ~n1086 & n1120 ;
  assign n1123 = n1122 ^ n1121 ;
  assign n1093 = n1092 ^ n1089 ;
  assign n1094 = ~n1086 & ~n1093 ;
  assign n1096 = n1013 & ~n1048 ;
  assign n1095 = n1010 & n1048 ;
  assign n1097 = n1096 ^ n1095 ;
  assign n1099 = n687 & ~n727 ;
  assign n1098 = n690 & n727 ;
  assign n1100 = n1099 ^ n1098 ;
  assign n1117 = ~n1097 & n1100 ;
  assign n1101 = n1100 ^ n1097 ;
  assign n1103 = n1019 & n1048 ;
  assign n1104 = n1103 ^ n1019 ;
  assign n1102 = n1017 & n1048 ;
  assign n1105 = n1104 ^ n1102 ;
  assign n1107 = n781 ^ n695 ;
  assign n1106 = n698 & n727 ;
  assign n1108 = n1107 ^ n1106 ;
  assign n1113 = n1105 & n1108 ;
  assign n1114 = n1113 ^ n1108 ;
  assign n1115 = n1101 & n1114 ;
  assign n1116 = n1115 ^ n1114 ;
  assign n1118 = n1117 ^ n1116 ;
  assign n1119 = n1094 & n1118 ;
  assign n1124 = n1123 ^ n1119 ;
  assign n1125 = n1079 & n1124 ;
  assign n1136 = n1135 ^ n1125 ;
  assign n1109 = n1108 ^ n1105 ;
  assign n1110 = ~n1101 & ~n1109 ;
  assign n1111 = n1094 & n1110 ;
  assign n1112 = n1079 & n1111 ;
  assign n1137 = n1136 ^ n1112 ;
  assign n1139 = n1054 & n1137 ;
  assign n1140 = n1139 ^ n1054 ;
  assign n1138 = n1051 & n1137 ;
  assign n1141 = n1140 ^ n1138 ;
  assign n1143 = n1061 & n1137 ;
  assign n1144 = n1143 ^ n1061 ;
  assign n1142 = n1058 & n1137 ;
  assign n1145 = n1144 ^ n1142 ;
  assign n1147 = n1069 & n1137 ;
  assign n1148 = n1147 ^ n1069 ;
  assign n1146 = n1066 & n1137 ;
  assign n1149 = n1148 ^ n1146 ;
  assign n1151 = n1076 & n1137 ;
  assign n1152 = n1151 ^ n1076 ;
  assign n1150 = n1073 & n1137 ;
  assign n1153 = n1152 ^ n1150 ;
  assign n1155 = n1085 & n1137 ;
  assign n1156 = n1155 ^ n1085 ;
  assign n1154 = n1082 & n1137 ;
  assign n1157 = n1156 ^ n1154 ;
  assign n1159 = n1092 & n1137 ;
  assign n1160 = n1159 ^ n1092 ;
  assign n1158 = n1089 & n1137 ;
  assign n1161 = n1160 ^ n1158 ;
  assign n1163 = n1100 & n1137 ;
  assign n1164 = n1163 ^ n1100 ;
  assign n1162 = n1097 & n1137 ;
  assign n1165 = n1164 ^ n1162 ;
  assign n1167 = n1108 & n1137 ;
  assign n1168 = n1167 ^ n1108 ;
  assign n1166 = n1105 & n1137 ;
  assign n1169 = n1168 ^ n1166 ;
  assign n1170 = n1138 ^ n1051 ;
  assign n1171 = n1170 ^ n1139 ;
  assign n1172 = n1142 ^ n1058 ;
  assign n1173 = n1172 ^ n1143 ;
  assign n1174 = n1146 ^ n1066 ;
  assign n1175 = n1174 ^ n1147 ;
  assign n1176 = n1150 ^ n1073 ;
  assign n1177 = n1176 ^ n1151 ;
  assign n1178 = n1154 ^ n1082 ;
  assign n1179 = n1178 ^ n1155 ;
  assign n1180 = n1158 ^ n1089 ;
  assign n1181 = n1180 ^ n1159 ;
  assign n1182 = n1162 ^ n1097 ;
  assign n1183 = n1182 ^ n1163 ;
  assign n1184 = n1166 ^ n1105 ;
  assign n1185 = n1184 ^ n1167 ;
  assign n1190 = n964 & ~n1048 ;
  assign n1189 = n967 & n1048 ;
  assign n1191 = n1190 ^ n1189 ;
  assign n1187 = n877 & ~n961 ;
  assign n1186 = n880 & n961 ;
  assign n1188 = n1187 ^ n1186 ;
  assign n1274 = ~n1188 & n1191 ;
  assign n1192 = n1191 ^ n1188 ;
  assign n1194 = n883 & ~n961 ;
  assign n1193 = n886 & n961 ;
  assign n1195 = n1194 ^ n1193 ;
  assign n1197 = n971 & ~n1048 ;
  assign n1196 = n974 & n1048 ;
  assign n1198 = n1197 ^ n1196 ;
  assign n1272 = ~n1195 & n1198 ;
  assign n1273 = ~n1192 & n1272 ;
  assign n1275 = n1274 ^ n1273 ;
  assign n1199 = n1198 ^ n1195 ;
  assign n1200 = ~n1192 & ~n1199 ;
  assign n1202 = n890 & ~n961 ;
  assign n1201 = n893 & n961 ;
  assign n1203 = n1202 ^ n1201 ;
  assign n1205 = n979 & ~n1048 ;
  assign n1204 = n982 & n1048 ;
  assign n1206 = n1205 ^ n1204 ;
  assign n1269 = ~n1203 & n1206 ;
  assign n1207 = n1206 ^ n1203 ;
  assign n1209 = n896 & ~n961 ;
  assign n1208 = n899 & n961 ;
  assign n1210 = n1209 ^ n1208 ;
  assign n1212 = n986 & ~n1048 ;
  assign n1211 = n989 & n1048 ;
  assign n1213 = n1212 ^ n1211 ;
  assign n1267 = ~n1210 & n1213 ;
  assign n1268 = ~n1207 & n1267 ;
  assign n1270 = n1269 ^ n1268 ;
  assign n1271 = n1200 & n1270 ;
  assign n1276 = n1275 ^ n1271 ;
  assign n1214 = n1213 ^ n1210 ;
  assign n1215 = ~n1207 & ~n1214 ;
  assign n1216 = n1200 & n1215 ;
  assign n1218 = n904 & ~n961 ;
  assign n1217 = n907 & n961 ;
  assign n1219 = n1218 ^ n1217 ;
  assign n1221 = n995 & ~n1048 ;
  assign n1220 = n998 & n1048 ;
  assign n1222 = n1221 ^ n1220 ;
  assign n1263 = ~n1219 & n1222 ;
  assign n1223 = n1222 ^ n1219 ;
  assign n1225 = n910 & ~n961 ;
  assign n1224 = n913 & n961 ;
  assign n1226 = n1225 ^ n1224 ;
  assign n1228 = n1002 & ~n1048 ;
  assign n1227 = n1005 & n1048 ;
  assign n1229 = n1228 ^ n1227 ;
  assign n1261 = ~n1226 & n1229 ;
  assign n1262 = ~n1223 & n1261 ;
  assign n1264 = n1263 ^ n1262 ;
  assign n1230 = n1229 ^ n1226 ;
  assign n1231 = ~n1223 & ~n1230 ;
  assign n1233 = n917 & ~n961 ;
  assign n1232 = n920 & n961 ;
  assign n1234 = n1233 ^ n1232 ;
  assign n1236 = n1010 & ~n1048 ;
  assign n1235 = n1013 & n1048 ;
  assign n1237 = n1236 ^ n1235 ;
  assign n1258 = ~n1234 & n1237 ;
  assign n1242 = n926 & ~n961 ;
  assign n1241 = n923 & n961 ;
  assign n1243 = n1242 ^ n1241 ;
  assign n1250 = n1019 & ~n1243 ;
  assign n1251 = n1048 & n1250 ;
  assign n1248 = n1017 & ~n1243 ;
  assign n1249 = ~n1048 & n1248 ;
  assign n1252 = n1251 ^ n1249 ;
  assign n1256 = ~n1234 & n1252 ;
  assign n1254 = n1236 & n1252 ;
  assign n1253 = n1235 & n1252 ;
  assign n1255 = n1254 ^ n1253 ;
  assign n1257 = n1256 ^ n1255 ;
  assign n1259 = n1258 ^ n1257 ;
  assign n1260 = n1231 & n1259 ;
  assign n1265 = n1264 ^ n1260 ;
  assign n1266 = n1216 & n1265 ;
  assign n1277 = n1276 ^ n1266 ;
  assign n1238 = n1237 ^ n1234 ;
  assign n1239 = n1017 & ~n1048 ;
  assign n1240 = n1239 ^ n1103 ;
  assign n1244 = n1243 ^ n1240 ;
  assign n1245 = ~n1238 & ~n1244 ;
  assign n1246 = n1231 & n1245 ;
  assign n1247 = n1216 & n1246 ;
  assign n1278 = n1277 ^ n1247 ;
  assign n1280 = n1191 & ~n1278 ;
  assign n1279 = n1188 & n1278 ;
  assign n1281 = n1280 ^ n1279 ;
  assign n1283 = n1198 & ~n1278 ;
  assign n1282 = n1195 & n1278 ;
  assign n1284 = n1283 ^ n1282 ;
  assign n1286 = n1206 & ~n1278 ;
  assign n1285 = n1203 & n1278 ;
  assign n1287 = n1286 ^ n1285 ;
  assign n1289 = n1213 & ~n1278 ;
  assign n1288 = n1210 & n1278 ;
  assign n1290 = n1289 ^ n1288 ;
  assign n1292 = n1222 & ~n1278 ;
  assign n1291 = n1219 & n1278 ;
  assign n1293 = n1292 ^ n1291 ;
  assign n1295 = n1229 & ~n1278 ;
  assign n1294 = n1226 & n1278 ;
  assign n1296 = n1295 ^ n1294 ;
  assign n1298 = n1237 & ~n1278 ;
  assign n1297 = n1234 & n1278 ;
  assign n1299 = n1298 ^ n1297 ;
  assign n1301 = n1240 & ~n1278 ;
  assign n1300 = n1243 & n1278 ;
  assign n1302 = n1301 ^ n1300 ;
  assign n1304 = n1188 & ~n1278 ;
  assign n1303 = n1191 & n1278 ;
  assign n1305 = n1304 ^ n1303 ;
  assign n1307 = n1195 & ~n1278 ;
  assign n1306 = n1198 & n1278 ;
  assign n1308 = n1307 ^ n1306 ;
  assign n1310 = n1203 & ~n1278 ;
  assign n1309 = n1206 & n1278 ;
  assign n1311 = n1310 ^ n1309 ;
  assign n1313 = n1210 & ~n1278 ;
  assign n1312 = n1213 & n1278 ;
  assign n1314 = n1313 ^ n1312 ;
  assign n1316 = n1219 & ~n1278 ;
  assign n1315 = n1222 & n1278 ;
  assign n1317 = n1316 ^ n1315 ;
  assign n1319 = n1226 & ~n1278 ;
  assign n1318 = n1229 & n1278 ;
  assign n1320 = n1319 ^ n1318 ;
  assign n1322 = n1234 & ~n1278 ;
  assign n1321 = n1237 & n1278 ;
  assign n1323 = n1322 ^ n1321 ;
  assign n1325 = n1243 & ~n1278 ;
  assign n1324 = n1240 & n1278 ;
  assign n1326 = n1325 ^ n1324 ;
  assign y0 = n830 ;
  assign y1 = n833 ;
  assign y2 = n836 ;
  assign y3 = n839 ;
  assign y4 = n842 ;
  assign y5 = n845 ;
  assign y6 = n848 ;
  assign y7 = n851 ;
  assign y8 = n854 ;
  assign y9 = n857 ;
  assign y10 = n860 ;
  assign y11 = n863 ;
  assign y12 = n866 ;
  assign y13 = n869 ;
  assign y14 = n872 ;
  assign y15 = n875 ;
  assign y16 = n1141 ;
  assign y17 = n1145 ;
  assign y18 = n1149 ;
  assign y19 = n1153 ;
  assign y20 = n1157 ;
  assign y21 = n1161 ;
  assign y22 = n1165 ;
  assign y23 = n1169 ;
  assign y24 = n1171 ;
  assign y25 = n1173 ;
  assign y26 = n1175 ;
  assign y27 = n1177 ;
  assign y28 = n1179 ;
  assign y29 = n1181 ;
  assign y30 = n1183 ;
  assign y31 = n1185 ;
  assign y32 = n1281 ;
  assign y33 = n1284 ;
  assign y34 = n1287 ;
  assign y35 = n1290 ;
  assign y36 = n1293 ;
  assign y37 = n1296 ;
  assign y38 = n1299 ;
  assign y39 = n1302 ;
  assign y40 = n1305 ;
  assign y41 = n1308 ;
  assign y42 = n1311 ;
  assign y43 = n1314 ;
  assign y44 = n1317 ;
  assign y45 = n1320 ;
  assign y46 = n1323 ;
  assign y47 = n1326 ;
endmodule
