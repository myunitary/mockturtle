// nine parties (one provide the reference data), each holding a 32-bit data, finding the two closest to the reference
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 ;
  assign n378 = x285 ^ x29 ;
  assign n377 = x286 ^ x30 ;
  assign n379 = n378 ^ n377 ;
  assign n376 = x287 ^ x31 ;
  assign n411 = n377 ^ n376 ;
  assign n412 = n379 & ~n411 ;
  assign n413 = n412 ^ n378 ;
  assign n381 = x281 ^ x25 ;
  assign n380 = n379 ^ n376 ;
  assign n382 = n381 ^ n380 ;
  assign n373 = x283 ^ x27 ;
  assign n372 = x282 ^ x26 ;
  assign n374 = n373 ^ n372 ;
  assign n371 = x284 ^ x28 ;
  assign n375 = n374 ^ n371 ;
  assign n408 = n380 ^ n375 ;
  assign n409 = n382 & ~n408 ;
  assign n410 = n409 ^ n381 ;
  assign n414 = n413 ^ n410 ;
  assign n405 = n372 ^ n371 ;
  assign n406 = n374 & ~n405 ;
  assign n407 = n406 ^ n373 ;
  assign n429 = n410 ^ n407 ;
  assign n430 = n414 & ~n429 ;
  assign n431 = n430 ^ n413 ;
  assign n415 = n414 ^ n407 ;
  assign n383 = n382 ^ n375 ;
  assign n370 = x273 ^ x17 ;
  assign n384 = n383 ^ n370 ;
  assign n365 = x279 ^ x23 ;
  assign n364 = x278 ^ x22 ;
  assign n366 = n365 ^ n364 ;
  assign n363 = x280 ^ x24 ;
  assign n367 = n366 ^ n363 ;
  assign n362 = x274 ^ x18 ;
  assign n368 = n367 ^ n362 ;
  assign n359 = x276 ^ x20 ;
  assign n358 = x275 ^ x19 ;
  assign n360 = n359 ^ n358 ;
  assign n357 = x277 ^ x21 ;
  assign n361 = n360 ^ n357 ;
  assign n369 = n368 ^ n361 ;
  assign n402 = n370 ^ n369 ;
  assign n403 = n384 & ~n402 ;
  assign n404 = n403 ^ n383 ;
  assign n416 = n415 ^ n404 ;
  assign n397 = n362 ^ n361 ;
  assign n398 = n368 & ~n397 ;
  assign n399 = n398 ^ n367 ;
  assign n394 = n364 ^ n363 ;
  assign n395 = n366 & ~n394 ;
  assign n396 = n395 ^ n365 ;
  assign n400 = n399 ^ n396 ;
  assign n391 = n358 ^ n357 ;
  assign n392 = n360 & ~n391 ;
  assign n393 = n392 ^ n359 ;
  assign n401 = n400 ^ n393 ;
  assign n426 = n415 ^ n401 ;
  assign n427 = n416 & ~n426 ;
  assign n428 = n427 ^ n404 ;
  assign n432 = n431 ^ n428 ;
  assign n423 = n396 ^ n393 ;
  assign n424 = n400 & ~n423 ;
  assign n425 = n424 ^ n399 ;
  assign n439 = n428 ^ n425 ;
  assign n440 = n432 & ~n439 ;
  assign n441 = n440 ^ n431 ;
  assign n433 = n432 ^ n425 ;
  assign n417 = n416 ^ n401 ;
  assign n385 = n384 ^ n369 ;
  assign n356 = x257 ^ x1 ;
  assign n386 = n385 ^ n356 ;
  assign n326 = x261 ^ x5 ;
  assign n325 = x260 ^ x4 ;
  assign n327 = n326 ^ n325 ;
  assign n324 = x262 ^ x6 ;
  assign n328 = n327 ^ n324 ;
  assign n320 = x264 ^ x8 ;
  assign n319 = x263 ^ x7 ;
  assign n321 = n320 ^ n319 ;
  assign n318 = x265 ^ x9 ;
  assign n322 = n321 ^ n318 ;
  assign n317 = x259 ^ x3 ;
  assign n323 = n322 ^ n317 ;
  assign n329 = n328 ^ n323 ;
  assign n315 = x258 ^ x2 ;
  assign n301 = x268 ^ x12 ;
  assign n300 = x267 ^ x11 ;
  assign n302 = n301 ^ n300 ;
  assign n299 = x269 ^ x13 ;
  assign n303 = n302 ^ n299 ;
  assign n292 = x272 ^ x16 ;
  assign n290 = x271 ^ x15 ;
  assign n289 = x270 ^ x14 ;
  assign n291 = n290 ^ n289 ;
  assign n297 = n292 ^ n291 ;
  assign n296 = x266 ^ x10 ;
  assign n298 = n297 ^ n296 ;
  assign n314 = n303 ^ n298 ;
  assign n316 = n315 ^ n314 ;
  assign n387 = n329 ^ n316 ;
  assign n388 = n387 ^ n356 ;
  assign n389 = n386 & ~n388 ;
  assign n390 = n389 ^ n385 ;
  assign n418 = n417 ^ n390 ;
  assign n341 = n319 ^ n318 ;
  assign n342 = n321 & ~n341 ;
  assign n343 = n342 ^ n320 ;
  assign n338 = n328 ^ n322 ;
  assign n339 = ~n323 & n338 ;
  assign n340 = n339 ^ n328 ;
  assign n344 = n343 ^ n340 ;
  assign n335 = n325 ^ n324 ;
  assign n336 = n327 & ~n335 ;
  assign n337 = n336 ^ n326 ;
  assign n345 = n344 ^ n337 ;
  assign n308 = n300 ^ n299 ;
  assign n309 = n302 & ~n308 ;
  assign n310 = n309 ^ n301 ;
  assign n304 = n303 ^ n296 ;
  assign n305 = n298 & ~n304 ;
  assign n306 = n305 ^ n297 ;
  assign n293 = n292 ^ n289 ;
  assign n294 = n291 & ~n293 ;
  assign n295 = n294 ^ n290 ;
  assign n307 = n306 ^ n295 ;
  assign n333 = n310 ^ n307 ;
  assign n330 = n329 ^ n314 ;
  assign n331 = n316 & ~n330 ;
  assign n332 = n331 ^ n315 ;
  assign n334 = n333 ^ n332 ;
  assign n419 = n345 ^ n334 ;
  assign n420 = n419 ^ n417 ;
  assign n421 = n418 & ~n420 ;
  assign n422 = n421 ^ n390 ;
  assign n434 = n433 ^ n422 ;
  assign n350 = n340 ^ n337 ;
  assign n351 = n344 & ~n350 ;
  assign n352 = n351 ^ n343 ;
  assign n346 = n345 ^ n333 ;
  assign n347 = n334 & ~n346 ;
  assign n348 = n347 ^ n332 ;
  assign n311 = n310 ^ n295 ;
  assign n312 = n307 & ~n311 ;
  assign n313 = n312 ^ n306 ;
  assign n349 = n348 ^ n313 ;
  assign n435 = n352 ^ n349 ;
  assign n436 = n435 ^ n422 ;
  assign n437 = n434 & ~n436 ;
  assign n438 = n437 ^ n433 ;
  assign n442 = n441 ^ n438 ;
  assign n353 = n352 ^ n313 ;
  assign n354 = n349 & ~n353 ;
  assign n355 = n354 ^ n348 ;
  assign n443 = n442 ^ n355 ;
  assign n444 = n419 ^ n418 ;
  assign n445 = n387 ^ n386 ;
  assign n446 = x256 ^ x0 ;
  assign n447 = n445 & n446 ;
  assign n448 = n444 & n447 ;
  assign n449 = n435 ^ n434 ;
  assign n450 = n448 & n449 ;
  assign n451 = n443 & n450 ;
  assign n452 = n441 ^ n355 ;
  assign n453 = ~n442 & n452 ;
  assign n454 = n453 ^ n355 ;
  assign n455 = n451 & n454 ;
  assign n545 = x285 ^ x61 ;
  assign n544 = x286 ^ x62 ;
  assign n546 = n545 ^ n544 ;
  assign n543 = x287 ^ x63 ;
  assign n578 = n544 ^ n543 ;
  assign n579 = n546 & ~n578 ;
  assign n580 = n579 ^ n545 ;
  assign n548 = x281 ^ x57 ;
  assign n547 = n546 ^ n543 ;
  assign n549 = n548 ^ n547 ;
  assign n540 = x283 ^ x59 ;
  assign n539 = x282 ^ x58 ;
  assign n541 = n540 ^ n539 ;
  assign n538 = x284 ^ x60 ;
  assign n542 = n541 ^ n538 ;
  assign n575 = n547 ^ n542 ;
  assign n576 = n549 & ~n575 ;
  assign n577 = n576 ^ n548 ;
  assign n581 = n580 ^ n577 ;
  assign n572 = n539 ^ n538 ;
  assign n573 = n541 & ~n572 ;
  assign n574 = n573 ^ n540 ;
  assign n596 = n577 ^ n574 ;
  assign n597 = n581 & ~n596 ;
  assign n598 = n597 ^ n580 ;
  assign n582 = n581 ^ n574 ;
  assign n550 = n549 ^ n542 ;
  assign n537 = x273 ^ x49 ;
  assign n551 = n550 ^ n537 ;
  assign n532 = x279 ^ x55 ;
  assign n531 = x278 ^ x54 ;
  assign n533 = n532 ^ n531 ;
  assign n530 = x280 ^ x56 ;
  assign n534 = n533 ^ n530 ;
  assign n529 = x274 ^ x50 ;
  assign n535 = n534 ^ n529 ;
  assign n526 = x276 ^ x52 ;
  assign n525 = x275 ^ x51 ;
  assign n527 = n526 ^ n525 ;
  assign n524 = x277 ^ x53 ;
  assign n528 = n527 ^ n524 ;
  assign n536 = n535 ^ n528 ;
  assign n569 = n537 ^ n536 ;
  assign n570 = n551 & ~n569 ;
  assign n571 = n570 ^ n550 ;
  assign n583 = n582 ^ n571 ;
  assign n564 = n529 ^ n528 ;
  assign n565 = n535 & ~n564 ;
  assign n566 = n565 ^ n534 ;
  assign n561 = n531 ^ n530 ;
  assign n562 = n533 & ~n561 ;
  assign n563 = n562 ^ n532 ;
  assign n567 = n566 ^ n563 ;
  assign n558 = n525 ^ n524 ;
  assign n559 = n527 & ~n558 ;
  assign n560 = n559 ^ n526 ;
  assign n568 = n567 ^ n560 ;
  assign n593 = n582 ^ n568 ;
  assign n594 = n583 & ~n593 ;
  assign n595 = n594 ^ n571 ;
  assign n599 = n598 ^ n595 ;
  assign n590 = n563 ^ n560 ;
  assign n591 = n567 & ~n590 ;
  assign n592 = n591 ^ n566 ;
  assign n606 = n595 ^ n592 ;
  assign n607 = n599 & ~n606 ;
  assign n608 = n607 ^ n598 ;
  assign n600 = n599 ^ n592 ;
  assign n584 = n583 ^ n568 ;
  assign n552 = n551 ^ n536 ;
  assign n523 = x257 ^ x33 ;
  assign n553 = n552 ^ n523 ;
  assign n493 = x261 ^ x37 ;
  assign n492 = x260 ^ x36 ;
  assign n494 = n493 ^ n492 ;
  assign n491 = x262 ^ x38 ;
  assign n495 = n494 ^ n491 ;
  assign n487 = x264 ^ x40 ;
  assign n486 = x263 ^ x39 ;
  assign n488 = n487 ^ n486 ;
  assign n485 = x265 ^ x41 ;
  assign n489 = n488 ^ n485 ;
  assign n484 = x259 ^ x35 ;
  assign n490 = n489 ^ n484 ;
  assign n496 = n495 ^ n490 ;
  assign n482 = x258 ^ x34 ;
  assign n468 = x268 ^ x44 ;
  assign n467 = x267 ^ x43 ;
  assign n469 = n468 ^ n467 ;
  assign n466 = x269 ^ x45 ;
  assign n470 = n469 ^ n466 ;
  assign n459 = x272 ^ x48 ;
  assign n457 = x271 ^ x47 ;
  assign n456 = x270 ^ x46 ;
  assign n458 = n457 ^ n456 ;
  assign n464 = n459 ^ n458 ;
  assign n463 = x266 ^ x42 ;
  assign n465 = n464 ^ n463 ;
  assign n481 = n470 ^ n465 ;
  assign n483 = n482 ^ n481 ;
  assign n554 = n496 ^ n483 ;
  assign n555 = n554 ^ n523 ;
  assign n556 = n553 & ~n555 ;
  assign n557 = n556 ^ n552 ;
  assign n585 = n584 ^ n557 ;
  assign n508 = n486 ^ n485 ;
  assign n509 = n488 & ~n508 ;
  assign n510 = n509 ^ n487 ;
  assign n505 = n495 ^ n489 ;
  assign n506 = ~n490 & n505 ;
  assign n507 = n506 ^ n495 ;
  assign n511 = n510 ^ n507 ;
  assign n502 = n492 ^ n491 ;
  assign n503 = n494 & ~n502 ;
  assign n504 = n503 ^ n493 ;
  assign n512 = n511 ^ n504 ;
  assign n475 = n467 ^ n466 ;
  assign n476 = n469 & ~n475 ;
  assign n477 = n476 ^ n468 ;
  assign n471 = n470 ^ n463 ;
  assign n472 = n465 & ~n471 ;
  assign n473 = n472 ^ n464 ;
  assign n460 = n459 ^ n456 ;
  assign n461 = n458 & ~n460 ;
  assign n462 = n461 ^ n457 ;
  assign n474 = n473 ^ n462 ;
  assign n500 = n477 ^ n474 ;
  assign n497 = n496 ^ n481 ;
  assign n498 = n483 & ~n497 ;
  assign n499 = n498 ^ n482 ;
  assign n501 = n500 ^ n499 ;
  assign n586 = n512 ^ n501 ;
  assign n587 = n586 ^ n584 ;
  assign n588 = n585 & ~n587 ;
  assign n589 = n588 ^ n557 ;
  assign n601 = n600 ^ n589 ;
  assign n517 = n507 ^ n504 ;
  assign n518 = n511 & ~n517 ;
  assign n519 = n518 ^ n510 ;
  assign n513 = n512 ^ n500 ;
  assign n514 = n501 & ~n513 ;
  assign n515 = n514 ^ n499 ;
  assign n478 = n477 ^ n462 ;
  assign n479 = n474 & ~n478 ;
  assign n480 = n479 ^ n473 ;
  assign n516 = n515 ^ n480 ;
  assign n602 = n519 ^ n516 ;
  assign n603 = n602 ^ n589 ;
  assign n604 = n601 & ~n603 ;
  assign n605 = n604 ^ n600 ;
  assign n609 = n608 ^ n605 ;
  assign n520 = n519 ^ n480 ;
  assign n521 = n516 & ~n520 ;
  assign n522 = n521 ^ n515 ;
  assign n610 = n609 ^ n522 ;
  assign n611 = n586 ^ n585 ;
  assign n612 = n554 ^ n553 ;
  assign n613 = x256 ^ x32 ;
  assign n614 = n612 & n613 ;
  assign n615 = n611 & n614 ;
  assign n616 = n602 ^ n601 ;
  assign n617 = n615 & n616 ;
  assign n618 = n610 & n617 ;
  assign n619 = n608 ^ n522 ;
  assign n620 = ~n609 & n619 ;
  assign n621 = n620 ^ n522 ;
  assign n622 = n618 & n621 ;
  assign n1564 = x285 ^ x125 ;
  assign n1563 = x286 ^ x126 ;
  assign n1565 = n1564 ^ n1563 ;
  assign n1562 = x287 ^ x127 ;
  assign n1597 = n1563 ^ n1562 ;
  assign n1598 = n1565 & ~n1597 ;
  assign n1599 = n1598 ^ n1564 ;
  assign n1567 = x281 ^ x121 ;
  assign n1566 = n1565 ^ n1562 ;
  assign n1568 = n1567 ^ n1566 ;
  assign n1559 = x283 ^ x123 ;
  assign n1558 = x282 ^ x122 ;
  assign n1560 = n1559 ^ n1558 ;
  assign n1557 = x284 ^ x124 ;
  assign n1561 = n1560 ^ n1557 ;
  assign n1594 = n1566 ^ n1561 ;
  assign n1595 = n1568 & ~n1594 ;
  assign n1596 = n1595 ^ n1567 ;
  assign n1600 = n1599 ^ n1596 ;
  assign n1591 = n1558 ^ n1557 ;
  assign n1592 = n1560 & ~n1591 ;
  assign n1593 = n1592 ^ n1559 ;
  assign n1615 = n1596 ^ n1593 ;
  assign n1616 = n1600 & ~n1615 ;
  assign n1617 = n1616 ^ n1599 ;
  assign n1601 = n1600 ^ n1593 ;
  assign n1569 = n1568 ^ n1561 ;
  assign n1556 = x273 ^ x113 ;
  assign n1570 = n1569 ^ n1556 ;
  assign n1551 = x279 ^ x119 ;
  assign n1550 = x278 ^ x118 ;
  assign n1552 = n1551 ^ n1550 ;
  assign n1549 = x280 ^ x120 ;
  assign n1553 = n1552 ^ n1549 ;
  assign n1548 = x274 ^ x114 ;
  assign n1554 = n1553 ^ n1548 ;
  assign n1545 = x276 ^ x116 ;
  assign n1544 = x275 ^ x115 ;
  assign n1546 = n1545 ^ n1544 ;
  assign n1543 = x277 ^ x117 ;
  assign n1547 = n1546 ^ n1543 ;
  assign n1555 = n1554 ^ n1547 ;
  assign n1588 = n1556 ^ n1555 ;
  assign n1589 = n1570 & ~n1588 ;
  assign n1590 = n1589 ^ n1569 ;
  assign n1602 = n1601 ^ n1590 ;
  assign n1583 = n1548 ^ n1547 ;
  assign n1584 = n1554 & ~n1583 ;
  assign n1585 = n1584 ^ n1553 ;
  assign n1580 = n1550 ^ n1549 ;
  assign n1581 = n1552 & ~n1580 ;
  assign n1582 = n1581 ^ n1551 ;
  assign n1586 = n1585 ^ n1582 ;
  assign n1577 = n1544 ^ n1543 ;
  assign n1578 = n1546 & ~n1577 ;
  assign n1579 = n1578 ^ n1545 ;
  assign n1587 = n1586 ^ n1579 ;
  assign n1612 = n1601 ^ n1587 ;
  assign n1613 = n1602 & ~n1612 ;
  assign n1614 = n1613 ^ n1590 ;
  assign n1618 = n1617 ^ n1614 ;
  assign n1609 = n1582 ^ n1579 ;
  assign n1610 = n1586 & ~n1609 ;
  assign n1611 = n1610 ^ n1585 ;
  assign n1625 = n1614 ^ n1611 ;
  assign n1626 = n1618 & ~n1625 ;
  assign n1627 = n1626 ^ n1617 ;
  assign n1619 = n1618 ^ n1611 ;
  assign n1603 = n1602 ^ n1587 ;
  assign n1571 = n1570 ^ n1555 ;
  assign n1542 = x257 ^ x97 ;
  assign n1572 = n1571 ^ n1542 ;
  assign n1512 = x261 ^ x101 ;
  assign n1511 = x260 ^ x100 ;
  assign n1513 = n1512 ^ n1511 ;
  assign n1510 = x262 ^ x102 ;
  assign n1514 = n1513 ^ n1510 ;
  assign n1506 = x264 ^ x104 ;
  assign n1505 = x263 ^ x103 ;
  assign n1507 = n1506 ^ n1505 ;
  assign n1504 = x265 ^ x105 ;
  assign n1508 = n1507 ^ n1504 ;
  assign n1503 = x259 ^ x99 ;
  assign n1509 = n1508 ^ n1503 ;
  assign n1515 = n1514 ^ n1509 ;
  assign n1501 = x258 ^ x98 ;
  assign n1487 = x268 ^ x108 ;
  assign n1486 = x267 ^ x107 ;
  assign n1488 = n1487 ^ n1486 ;
  assign n1485 = x269 ^ x109 ;
  assign n1489 = n1488 ^ n1485 ;
  assign n1478 = x272 ^ x112 ;
  assign n1476 = x271 ^ x111 ;
  assign n1475 = x270 ^ x110 ;
  assign n1477 = n1476 ^ n1475 ;
  assign n1483 = n1478 ^ n1477 ;
  assign n1482 = x266 ^ x106 ;
  assign n1484 = n1483 ^ n1482 ;
  assign n1500 = n1489 ^ n1484 ;
  assign n1502 = n1501 ^ n1500 ;
  assign n1573 = n1515 ^ n1502 ;
  assign n1574 = n1573 ^ n1542 ;
  assign n1575 = n1572 & ~n1574 ;
  assign n1576 = n1575 ^ n1571 ;
  assign n1604 = n1603 ^ n1576 ;
  assign n1527 = n1505 ^ n1504 ;
  assign n1528 = n1507 & ~n1527 ;
  assign n1529 = n1528 ^ n1506 ;
  assign n1524 = n1514 ^ n1508 ;
  assign n1525 = ~n1509 & n1524 ;
  assign n1526 = n1525 ^ n1514 ;
  assign n1530 = n1529 ^ n1526 ;
  assign n1521 = n1511 ^ n1510 ;
  assign n1522 = n1513 & ~n1521 ;
  assign n1523 = n1522 ^ n1512 ;
  assign n1531 = n1530 ^ n1523 ;
  assign n1494 = n1486 ^ n1485 ;
  assign n1495 = n1488 & ~n1494 ;
  assign n1496 = n1495 ^ n1487 ;
  assign n1490 = n1489 ^ n1482 ;
  assign n1491 = n1484 & ~n1490 ;
  assign n1492 = n1491 ^ n1483 ;
  assign n1479 = n1478 ^ n1475 ;
  assign n1480 = n1477 & ~n1479 ;
  assign n1481 = n1480 ^ n1476 ;
  assign n1493 = n1492 ^ n1481 ;
  assign n1519 = n1496 ^ n1493 ;
  assign n1516 = n1515 ^ n1500 ;
  assign n1517 = n1502 & ~n1516 ;
  assign n1518 = n1517 ^ n1501 ;
  assign n1520 = n1519 ^ n1518 ;
  assign n1605 = n1531 ^ n1520 ;
  assign n1606 = n1605 ^ n1603 ;
  assign n1607 = n1604 & ~n1606 ;
  assign n1608 = n1607 ^ n1576 ;
  assign n1620 = n1619 ^ n1608 ;
  assign n1536 = n1526 ^ n1523 ;
  assign n1537 = n1530 & ~n1536 ;
  assign n1538 = n1537 ^ n1529 ;
  assign n1532 = n1531 ^ n1519 ;
  assign n1533 = n1520 & ~n1532 ;
  assign n1534 = n1533 ^ n1518 ;
  assign n1497 = n1496 ^ n1481 ;
  assign n1498 = n1493 & ~n1497 ;
  assign n1499 = n1498 ^ n1492 ;
  assign n1535 = n1534 ^ n1499 ;
  assign n1621 = n1538 ^ n1535 ;
  assign n1622 = n1621 ^ n1608 ;
  assign n1623 = n1620 & ~n1622 ;
  assign n1624 = n1623 ^ n1619 ;
  assign n1628 = n1627 ^ n1624 ;
  assign n1539 = n1538 ^ n1499 ;
  assign n1540 = n1535 & ~n1539 ;
  assign n1541 = n1540 ^ n1534 ;
  assign n1629 = n1628 ^ n1541 ;
  assign n1630 = n1605 ^ n1604 ;
  assign n1631 = n1573 ^ n1572 ;
  assign n1632 = x256 ^ x96 ;
  assign n1633 = n1631 & n1632 ;
  assign n1634 = n1630 & n1633 ;
  assign n1635 = n1621 ^ n1620 ;
  assign n1636 = n1634 & n1635 ;
  assign n1637 = n1629 & n1636 ;
  assign n1638 = n1627 ^ n1541 ;
  assign n1639 = ~n1628 & n1638 ;
  assign n1640 = n1639 ^ n1541 ;
  assign n1641 = n1637 & n1640 ;
  assign n879 = x285 ^ x157 ;
  assign n878 = x286 ^ x158 ;
  assign n880 = n879 ^ n878 ;
  assign n877 = x287 ^ x159 ;
  assign n912 = n878 ^ n877 ;
  assign n913 = n880 & ~n912 ;
  assign n914 = n913 ^ n879 ;
  assign n882 = x281 ^ x153 ;
  assign n881 = n880 ^ n877 ;
  assign n883 = n882 ^ n881 ;
  assign n874 = x283 ^ x155 ;
  assign n873 = x282 ^ x154 ;
  assign n875 = n874 ^ n873 ;
  assign n872 = x284 ^ x156 ;
  assign n876 = n875 ^ n872 ;
  assign n909 = n881 ^ n876 ;
  assign n910 = n883 & ~n909 ;
  assign n911 = n910 ^ n882 ;
  assign n915 = n914 ^ n911 ;
  assign n906 = n873 ^ n872 ;
  assign n907 = n875 & ~n906 ;
  assign n908 = n907 ^ n874 ;
  assign n930 = n911 ^ n908 ;
  assign n931 = n915 & ~n930 ;
  assign n932 = n931 ^ n914 ;
  assign n916 = n915 ^ n908 ;
  assign n884 = n883 ^ n876 ;
  assign n871 = x273 ^ x145 ;
  assign n885 = n884 ^ n871 ;
  assign n866 = x279 ^ x151 ;
  assign n865 = x278 ^ x150 ;
  assign n867 = n866 ^ n865 ;
  assign n864 = x280 ^ x152 ;
  assign n868 = n867 ^ n864 ;
  assign n863 = x274 ^ x146 ;
  assign n869 = n868 ^ n863 ;
  assign n860 = x276 ^ x148 ;
  assign n859 = x275 ^ x147 ;
  assign n861 = n860 ^ n859 ;
  assign n858 = x277 ^ x149 ;
  assign n862 = n861 ^ n858 ;
  assign n870 = n869 ^ n862 ;
  assign n903 = n871 ^ n870 ;
  assign n904 = n885 & ~n903 ;
  assign n905 = n904 ^ n884 ;
  assign n917 = n916 ^ n905 ;
  assign n898 = n863 ^ n862 ;
  assign n899 = n869 & ~n898 ;
  assign n900 = n899 ^ n868 ;
  assign n895 = n865 ^ n864 ;
  assign n896 = n867 & ~n895 ;
  assign n897 = n896 ^ n866 ;
  assign n901 = n900 ^ n897 ;
  assign n892 = n859 ^ n858 ;
  assign n893 = n861 & ~n892 ;
  assign n894 = n893 ^ n860 ;
  assign n902 = n901 ^ n894 ;
  assign n927 = n916 ^ n902 ;
  assign n928 = n917 & ~n927 ;
  assign n929 = n928 ^ n905 ;
  assign n933 = n932 ^ n929 ;
  assign n924 = n897 ^ n894 ;
  assign n925 = n901 & ~n924 ;
  assign n926 = n925 ^ n900 ;
  assign n940 = n929 ^ n926 ;
  assign n941 = n933 & ~n940 ;
  assign n942 = n941 ^ n932 ;
  assign n934 = n933 ^ n926 ;
  assign n918 = n917 ^ n902 ;
  assign n886 = n885 ^ n870 ;
  assign n857 = x257 ^ x129 ;
  assign n887 = n886 ^ n857 ;
  assign n827 = x261 ^ x133 ;
  assign n826 = x260 ^ x132 ;
  assign n828 = n827 ^ n826 ;
  assign n825 = x262 ^ x134 ;
  assign n829 = n828 ^ n825 ;
  assign n821 = x264 ^ x136 ;
  assign n820 = x263 ^ x135 ;
  assign n822 = n821 ^ n820 ;
  assign n819 = x265 ^ x137 ;
  assign n823 = n822 ^ n819 ;
  assign n818 = x259 ^ x131 ;
  assign n824 = n823 ^ n818 ;
  assign n830 = n829 ^ n824 ;
  assign n816 = x258 ^ x130 ;
  assign n802 = x268 ^ x140 ;
  assign n801 = x267 ^ x139 ;
  assign n803 = n802 ^ n801 ;
  assign n800 = x269 ^ x141 ;
  assign n804 = n803 ^ n800 ;
  assign n793 = x272 ^ x144 ;
  assign n791 = x271 ^ x143 ;
  assign n790 = x270 ^ x142 ;
  assign n792 = n791 ^ n790 ;
  assign n798 = n793 ^ n792 ;
  assign n797 = x266 ^ x138 ;
  assign n799 = n798 ^ n797 ;
  assign n815 = n804 ^ n799 ;
  assign n817 = n816 ^ n815 ;
  assign n888 = n830 ^ n817 ;
  assign n889 = n888 ^ n857 ;
  assign n890 = n887 & ~n889 ;
  assign n891 = n890 ^ n886 ;
  assign n919 = n918 ^ n891 ;
  assign n842 = n820 ^ n819 ;
  assign n843 = n822 & ~n842 ;
  assign n844 = n843 ^ n821 ;
  assign n839 = n829 ^ n823 ;
  assign n840 = ~n824 & n839 ;
  assign n841 = n840 ^ n829 ;
  assign n845 = n844 ^ n841 ;
  assign n836 = n826 ^ n825 ;
  assign n837 = n828 & ~n836 ;
  assign n838 = n837 ^ n827 ;
  assign n846 = n845 ^ n838 ;
  assign n809 = n801 ^ n800 ;
  assign n810 = n803 & ~n809 ;
  assign n811 = n810 ^ n802 ;
  assign n805 = n804 ^ n797 ;
  assign n806 = n799 & ~n805 ;
  assign n807 = n806 ^ n798 ;
  assign n794 = n793 ^ n790 ;
  assign n795 = n792 & ~n794 ;
  assign n796 = n795 ^ n791 ;
  assign n808 = n807 ^ n796 ;
  assign n834 = n811 ^ n808 ;
  assign n831 = n830 ^ n815 ;
  assign n832 = n817 & ~n831 ;
  assign n833 = n832 ^ n816 ;
  assign n835 = n834 ^ n833 ;
  assign n920 = n846 ^ n835 ;
  assign n921 = n920 ^ n918 ;
  assign n922 = n919 & ~n921 ;
  assign n923 = n922 ^ n891 ;
  assign n935 = n934 ^ n923 ;
  assign n851 = n841 ^ n838 ;
  assign n852 = n845 & ~n851 ;
  assign n853 = n852 ^ n844 ;
  assign n847 = n846 ^ n834 ;
  assign n848 = n835 & ~n847 ;
  assign n849 = n848 ^ n833 ;
  assign n812 = n811 ^ n796 ;
  assign n813 = n808 & ~n812 ;
  assign n814 = n813 ^ n807 ;
  assign n850 = n849 ^ n814 ;
  assign n936 = n853 ^ n850 ;
  assign n937 = n936 ^ n923 ;
  assign n938 = n935 & ~n937 ;
  assign n939 = n938 ^ n934 ;
  assign n943 = n942 ^ n939 ;
  assign n854 = n853 ^ n814 ;
  assign n855 = n850 & ~n854 ;
  assign n856 = n855 ^ n849 ;
  assign n944 = n943 ^ n856 ;
  assign n945 = n920 ^ n919 ;
  assign n946 = n888 ^ n887 ;
  assign n947 = x256 ^ x128 ;
  assign n948 = n946 & n947 ;
  assign n949 = n945 & n948 ;
  assign n950 = n936 ^ n935 ;
  assign n951 = n949 & n950 ;
  assign n952 = n944 & n951 ;
  assign n953 = n942 ^ n856 ;
  assign n954 = ~n943 & n953 ;
  assign n955 = n954 ^ n856 ;
  assign n956 = n952 & n955 ;
  assign n1031 = x276 ^ x244 ;
  assign n1030 = x275 ^ x243 ;
  assign n1032 = n1031 ^ n1030 ;
  assign n1029 = x277 ^ x245 ;
  assign n1041 = n1030 ^ n1029 ;
  assign n1042 = n1032 & ~n1041 ;
  assign n1043 = n1042 ^ n1031 ;
  assign n1025 = x279 ^ x247 ;
  assign n1024 = x278 ^ x246 ;
  assign n1026 = n1025 ^ n1024 ;
  assign n1023 = x280 ^ x248 ;
  assign n1037 = n1024 ^ n1023 ;
  assign n1038 = n1026 & ~n1037 ;
  assign n1039 = n1038 ^ n1025 ;
  assign n1027 = n1026 ^ n1023 ;
  assign n1022 = x274 ^ x242 ;
  assign n1028 = n1027 ^ n1022 ;
  assign n1033 = n1032 ^ n1029 ;
  assign n1034 = n1033 ^ n1022 ;
  assign n1035 = n1028 & ~n1034 ;
  assign n1036 = n1035 ^ n1027 ;
  assign n1040 = n1039 ^ n1036 ;
  assign n1081 = n1043 ^ n1040 ;
  assign n1059 = x283 ^ x251 ;
  assign n1058 = x282 ^ x250 ;
  assign n1060 = n1059 ^ n1058 ;
  assign n1057 = x284 ^ x252 ;
  assign n1066 = n1058 ^ n1057 ;
  assign n1067 = n1060 & ~n1066 ;
  assign n1068 = n1067 ^ n1059 ;
  assign n1055 = x281 ^ x249 ;
  assign n1050 = x287 ^ x255 ;
  assign n1048 = x286 ^ x254 ;
  assign n1047 = x285 ^ x253 ;
  assign n1049 = n1048 ^ n1047 ;
  assign n1054 = n1050 ^ n1049 ;
  assign n1056 = n1055 ^ n1054 ;
  assign n1061 = n1060 ^ n1057 ;
  assign n1062 = n1061 ^ n1054 ;
  assign n1063 = n1056 & ~n1062 ;
  assign n1064 = n1063 ^ n1055 ;
  assign n1051 = n1050 ^ n1048 ;
  assign n1052 = ~n1049 & n1051 ;
  assign n1053 = n1052 ^ n1050 ;
  assign n1065 = n1064 ^ n1053 ;
  assign n1079 = n1068 ^ n1065 ;
  assign n1073 = n1061 ^ n1056 ;
  assign n1072 = x273 ^ x241 ;
  assign n1074 = n1073 ^ n1072 ;
  assign n1075 = n1033 ^ n1028 ;
  assign n1076 = n1075 ^ n1072 ;
  assign n1077 = n1074 & ~n1076 ;
  assign n1078 = n1077 ^ n1073 ;
  assign n1080 = n1079 ^ n1078 ;
  assign n1094 = n1081 ^ n1080 ;
  assign n1088 = x257 ^ x225 ;
  assign n1087 = n1075 ^ n1074 ;
  assign n1089 = n1088 ^ n1087 ;
  assign n966 = x261 ^ x229 ;
  assign n965 = x260 ^ x228 ;
  assign n967 = n966 ^ n965 ;
  assign n964 = x262 ^ x230 ;
  assign n968 = n967 ^ n964 ;
  assign n960 = x264 ^ x232 ;
  assign n959 = x263 ^ x231 ;
  assign n961 = n960 ^ n959 ;
  assign n958 = x265 ^ x233 ;
  assign n962 = n961 ^ n958 ;
  assign n957 = x259 ^ x227 ;
  assign n963 = n962 ^ n957 ;
  assign n1013 = n968 ^ n963 ;
  assign n1011 = x258 ^ x226 ;
  assign n994 = x268 ^ x236 ;
  assign n993 = x267 ^ x235 ;
  assign n995 = n994 ^ n993 ;
  assign n992 = x269 ^ x237 ;
  assign n996 = n995 ^ n992 ;
  assign n990 = x266 ^ x234 ;
  assign n985 = x272 ^ x240 ;
  assign n983 = x271 ^ x239 ;
  assign n982 = x270 ^ x238 ;
  assign n984 = n983 ^ n982 ;
  assign n989 = n985 ^ n984 ;
  assign n991 = n990 ^ n989 ;
  assign n1010 = n996 ^ n991 ;
  assign n1012 = n1011 ^ n1010 ;
  assign n1090 = n1013 ^ n1012 ;
  assign n1091 = n1090 ^ n1087 ;
  assign n1092 = n1089 & ~n1091 ;
  assign n1093 = n1092 ^ n1088 ;
  assign n1095 = n1094 ^ n1093 ;
  assign n1014 = n1013 ^ n1011 ;
  assign n1015 = ~n1012 & n1014 ;
  assign n1016 = n1015 ^ n1013 ;
  assign n1001 = n993 ^ n992 ;
  assign n1002 = n995 & ~n1001 ;
  assign n1003 = n1002 ^ n994 ;
  assign n997 = n996 ^ n989 ;
  assign n998 = n991 & ~n997 ;
  assign n999 = n998 ^ n990 ;
  assign n986 = n985 ^ n983 ;
  assign n987 = ~n984 & n986 ;
  assign n988 = n987 ^ n985 ;
  assign n1000 = n999 ^ n988 ;
  assign n1008 = n1003 ^ n1000 ;
  assign n976 = n965 ^ n964 ;
  assign n977 = n967 & ~n976 ;
  assign n978 = n977 ^ n966 ;
  assign n972 = n959 ^ n958 ;
  assign n973 = n961 & ~n972 ;
  assign n974 = n973 ^ n960 ;
  assign n969 = n968 ^ n957 ;
  assign n970 = n963 & ~n969 ;
  assign n971 = n970 ^ n962 ;
  assign n975 = n974 ^ n971 ;
  assign n1007 = n978 ^ n975 ;
  assign n1009 = n1008 ^ n1007 ;
  assign n1096 = n1016 ^ n1009 ;
  assign n1097 = n1096 ^ n1094 ;
  assign n1098 = n1095 & ~n1097 ;
  assign n1099 = n1098 ^ n1093 ;
  assign n1082 = n1081 ^ n1079 ;
  assign n1083 = n1080 & ~n1082 ;
  assign n1084 = n1083 ^ n1078 ;
  assign n1069 = n1068 ^ n1064 ;
  assign n1070 = ~n1065 & n1069 ;
  assign n1071 = n1070 ^ n1068 ;
  assign n1085 = n1084 ^ n1071 ;
  assign n1044 = n1043 ^ n1036 ;
  assign n1045 = ~n1040 & n1044 ;
  assign n1046 = n1045 ^ n1043 ;
  assign n1086 = n1085 ^ n1046 ;
  assign n1100 = n1099 ^ n1086 ;
  assign n1017 = n1016 ^ n1007 ;
  assign n1018 = n1009 & ~n1017 ;
  assign n1019 = n1018 ^ n1008 ;
  assign n1004 = n1003 ^ n999 ;
  assign n1005 = ~n1000 & n1004 ;
  assign n1006 = n1005 ^ n1003 ;
  assign n1020 = n1019 ^ n1006 ;
  assign n979 = n978 ^ n971 ;
  assign n980 = ~n975 & n979 ;
  assign n981 = n980 ^ n978 ;
  assign n1021 = n1020 ^ n981 ;
  assign n1101 = n1100 ^ n1021 ;
  assign n1102 = n1096 ^ n1095 ;
  assign n1103 = x256 ^ x224 ;
  assign n1104 = n1090 ^ n1089 ;
  assign n1105 = n1103 & n1104 ;
  assign n1106 = n1102 & n1105 ;
  assign n1107 = n1101 & n1106 ;
  assign n1114 = n1086 ^ n1021 ;
  assign n1115 = n1100 & ~n1114 ;
  assign n1116 = n1115 ^ n1099 ;
  assign n1111 = n1071 ^ n1046 ;
  assign n1112 = n1085 & ~n1111 ;
  assign n1113 = n1112 ^ n1084 ;
  assign n1117 = n1116 ^ n1113 ;
  assign n1108 = n1006 ^ n981 ;
  assign n1109 = n1020 & ~n1108 ;
  assign n1110 = n1109 ^ n1019 ;
  assign n1118 = n1117 ^ n1110 ;
  assign n1119 = n1107 & n1118 ;
  assign n1120 = n1113 ^ n1110 ;
  assign n1121 = n1117 & ~n1120 ;
  assign n1122 = n1121 ^ n1116 ;
  assign n1123 = n1119 & n1122 ;
  assign n1179 = x266 ^ x202 ;
  assign n1177 = x272 ^ x208 ;
  assign n1175 = x271 ^ x207 ;
  assign n1174 = x270 ^ x206 ;
  assign n1176 = n1175 ^ n1174 ;
  assign n1178 = n1177 ^ n1176 ;
  assign n1180 = n1179 ^ n1178 ;
  assign n1171 = x268 ^ x204 ;
  assign n1170 = x267 ^ x203 ;
  assign n1172 = n1171 ^ n1170 ;
  assign n1169 = x269 ^ x205 ;
  assign n1173 = n1172 ^ n1169 ;
  assign n1235 = n1178 ^ n1173 ;
  assign n1236 = n1180 & ~n1235 ;
  assign n1237 = n1236 ^ n1179 ;
  assign n1232 = n1177 ^ n1175 ;
  assign n1233 = ~n1176 & n1232 ;
  assign n1234 = n1233 ^ n1177 ;
  assign n1238 = n1237 ^ n1234 ;
  assign n1229 = n1170 ^ n1169 ;
  assign n1230 = n1172 & ~n1229 ;
  assign n1231 = n1230 ^ n1171 ;
  assign n1239 = n1238 ^ n1231 ;
  assign n1163 = x264 ^ x200 ;
  assign n1162 = x263 ^ x199 ;
  assign n1164 = n1163 ^ n1162 ;
  assign n1161 = x265 ^ x201 ;
  assign n1224 = n1162 ^ n1161 ;
  assign n1225 = n1164 & ~n1224 ;
  assign n1226 = n1225 ^ n1163 ;
  assign n1165 = n1164 ^ n1161 ;
  assign n1160 = x259 ^ x195 ;
  assign n1166 = n1165 ^ n1160 ;
  assign n1157 = x261 ^ x197 ;
  assign n1156 = x260 ^ x196 ;
  assign n1158 = n1157 ^ n1156 ;
  assign n1155 = x262 ^ x198 ;
  assign n1159 = n1158 ^ n1155 ;
  assign n1221 = n1160 ^ n1159 ;
  assign n1222 = n1166 & ~n1221 ;
  assign n1223 = n1222 ^ n1165 ;
  assign n1227 = n1226 ^ n1223 ;
  assign n1218 = n1156 ^ n1155 ;
  assign n1219 = n1158 & ~n1218 ;
  assign n1220 = n1219 ^ n1157 ;
  assign n1228 = n1227 ^ n1220 ;
  assign n1240 = n1239 ^ n1228 ;
  assign n1181 = n1180 ^ n1173 ;
  assign n1168 = x258 ^ x194 ;
  assign n1182 = n1181 ^ n1168 ;
  assign n1167 = n1166 ^ n1159 ;
  assign n1215 = n1168 ^ n1167 ;
  assign n1216 = n1182 & ~n1215 ;
  assign n1217 = n1216 ^ n1181 ;
  assign n1263 = n1239 ^ n1217 ;
  assign n1264 = ~n1240 & n1263 ;
  assign n1265 = n1264 ^ n1217 ;
  assign n1260 = n1237 ^ n1231 ;
  assign n1261 = ~n1238 & n1260 ;
  assign n1262 = n1261 ^ n1231 ;
  assign n1266 = n1265 ^ n1262 ;
  assign n1257 = n1223 ^ n1220 ;
  assign n1258 = ~n1227 & n1257 ;
  assign n1259 = n1258 ^ n1220 ;
  assign n1267 = n1266 ^ n1259 ;
  assign n1146 = x285 ^ x221 ;
  assign n1145 = x286 ^ x222 ;
  assign n1147 = n1146 ^ n1145 ;
  assign n1144 = x287 ^ x223 ;
  assign n1207 = n1145 ^ n1144 ;
  assign n1208 = n1147 & ~n1207 ;
  assign n1209 = n1208 ^ n1146 ;
  assign n1148 = n1147 ^ n1144 ;
  assign n1143 = x281 ^ x217 ;
  assign n1149 = n1148 ^ n1143 ;
  assign n1140 = x283 ^ x219 ;
  assign n1139 = x282 ^ x218 ;
  assign n1141 = n1140 ^ n1139 ;
  assign n1138 = x284 ^ x220 ;
  assign n1142 = n1141 ^ n1138 ;
  assign n1204 = n1143 ^ n1142 ;
  assign n1205 = n1149 & ~n1204 ;
  assign n1206 = n1205 ^ n1148 ;
  assign n1210 = n1209 ^ n1206 ;
  assign n1201 = n1139 ^ n1138 ;
  assign n1202 = n1141 & ~n1201 ;
  assign n1203 = n1202 ^ n1140 ;
  assign n1251 = n1206 ^ n1203 ;
  assign n1252 = n1210 & ~n1251 ;
  assign n1253 = n1252 ^ n1209 ;
  assign n1211 = n1210 ^ n1203 ;
  assign n1150 = n1149 ^ n1142 ;
  assign n1137 = x273 ^ x209 ;
  assign n1151 = n1150 ^ n1137 ;
  assign n1134 = x277 ^ x213 ;
  assign n1132 = x275 ^ x211 ;
  assign n1131 = x276 ^ x212 ;
  assign n1133 = n1132 ^ n1131 ;
  assign n1135 = n1134 ^ n1133 ;
  assign n1129 = x274 ^ x210 ;
  assign n1127 = x280 ^ x216 ;
  assign n1125 = x278 ^ x214 ;
  assign n1124 = x279 ^ x215 ;
  assign n1126 = n1125 ^ n1124 ;
  assign n1128 = n1127 ^ n1126 ;
  assign n1130 = n1129 ^ n1128 ;
  assign n1136 = n1135 ^ n1130 ;
  assign n1198 = n1137 ^ n1136 ;
  assign n1199 = n1151 & ~n1198 ;
  assign n1200 = n1199 ^ n1150 ;
  assign n1212 = n1211 ^ n1200 ;
  assign n1193 = n1127 ^ n1124 ;
  assign n1194 = n1126 & ~n1193 ;
  assign n1195 = n1194 ^ n1125 ;
  assign n1190 = n1135 ^ n1128 ;
  assign n1191 = n1130 & ~n1190 ;
  assign n1192 = n1191 ^ n1129 ;
  assign n1196 = n1195 ^ n1192 ;
  assign n1187 = n1134 ^ n1131 ;
  assign n1188 = n1133 & ~n1187 ;
  assign n1189 = n1188 ^ n1132 ;
  assign n1197 = n1196 ^ n1189 ;
  assign n1248 = n1211 ^ n1197 ;
  assign n1249 = ~n1212 & n1248 ;
  assign n1250 = n1249 ^ n1197 ;
  assign n1254 = n1253 ^ n1250 ;
  assign n1245 = n1192 ^ n1189 ;
  assign n1246 = ~n1196 & n1245 ;
  assign n1247 = n1246 ^ n1189 ;
  assign n1255 = n1254 ^ n1247 ;
  assign n1213 = n1212 ^ n1197 ;
  assign n1153 = x257 ^ x193 ;
  assign n1152 = n1151 ^ n1136 ;
  assign n1154 = n1153 ^ n1152 ;
  assign n1183 = n1182 ^ n1167 ;
  assign n1184 = n1183 ^ n1152 ;
  assign n1185 = n1154 & ~n1184 ;
  assign n1186 = n1185 ^ n1153 ;
  assign n1214 = n1213 ^ n1186 ;
  assign n1241 = n1240 ^ n1217 ;
  assign n1242 = n1241 ^ n1213 ;
  assign n1243 = n1214 & ~n1242 ;
  assign n1244 = n1243 ^ n1186 ;
  assign n1256 = n1255 ^ n1244 ;
  assign n1281 = n1267 ^ n1256 ;
  assign n1282 = n1241 ^ n1214 ;
  assign n1283 = x256 ^ x192 ;
  assign n1284 = n1183 ^ n1154 ;
  assign n1285 = n1283 & n1284 ;
  assign n1286 = n1282 & n1285 ;
  assign n1287 = n1281 & n1286 ;
  assign n1275 = n1262 ^ n1259 ;
  assign n1276 = n1266 & ~n1275 ;
  assign n1277 = n1276 ^ n1265 ;
  assign n1271 = n1250 ^ n1247 ;
  assign n1272 = n1254 & ~n1271 ;
  assign n1273 = n1272 ^ n1253 ;
  assign n1268 = n1267 ^ n1255 ;
  assign n1269 = ~n1256 & n1268 ;
  assign n1270 = n1269 ^ n1267 ;
  assign n1274 = n1273 ^ n1270 ;
  assign n1288 = n1277 ^ n1274 ;
  assign n1289 = n1287 & n1288 ;
  assign n1278 = n1277 ^ n1270 ;
  assign n1279 = n1274 & ~n1278 ;
  assign n1280 = n1279 ^ n1273 ;
  assign n1291 = n1289 ^ n1280 ;
  assign n1290 = ~n1280 & ~n1289 ;
  assign n1292 = n1291 ^ n1290 ;
  assign n1293 = ~n1123 & ~n1292 ;
  assign n1294 = n1293 ^ n1123 ;
  assign n1386 = x285 ^ x189 ;
  assign n1385 = x286 ^ x190 ;
  assign n1387 = n1386 ^ n1385 ;
  assign n1384 = x287 ^ x191 ;
  assign n1419 = n1385 ^ n1384 ;
  assign n1420 = n1387 & ~n1419 ;
  assign n1421 = n1420 ^ n1386 ;
  assign n1389 = x281 ^ x185 ;
  assign n1388 = n1387 ^ n1384 ;
  assign n1390 = n1389 ^ n1388 ;
  assign n1381 = x283 ^ x187 ;
  assign n1380 = x282 ^ x186 ;
  assign n1382 = n1381 ^ n1380 ;
  assign n1379 = x284 ^ x188 ;
  assign n1383 = n1382 ^ n1379 ;
  assign n1416 = n1388 ^ n1383 ;
  assign n1417 = n1390 & ~n1416 ;
  assign n1418 = n1417 ^ n1389 ;
  assign n1422 = n1421 ^ n1418 ;
  assign n1413 = n1380 ^ n1379 ;
  assign n1414 = n1382 & ~n1413 ;
  assign n1415 = n1414 ^ n1381 ;
  assign n1437 = n1418 ^ n1415 ;
  assign n1438 = n1422 & ~n1437 ;
  assign n1439 = n1438 ^ n1421 ;
  assign n1423 = n1422 ^ n1415 ;
  assign n1391 = n1390 ^ n1383 ;
  assign n1378 = x273 ^ x177 ;
  assign n1392 = n1391 ^ n1378 ;
  assign n1373 = x279 ^ x183 ;
  assign n1372 = x278 ^ x182 ;
  assign n1374 = n1373 ^ n1372 ;
  assign n1371 = x280 ^ x184 ;
  assign n1375 = n1374 ^ n1371 ;
  assign n1370 = x274 ^ x178 ;
  assign n1376 = n1375 ^ n1370 ;
  assign n1367 = x276 ^ x180 ;
  assign n1366 = x275 ^ x179 ;
  assign n1368 = n1367 ^ n1366 ;
  assign n1365 = x277 ^ x181 ;
  assign n1369 = n1368 ^ n1365 ;
  assign n1377 = n1376 ^ n1369 ;
  assign n1410 = n1378 ^ n1377 ;
  assign n1411 = n1392 & ~n1410 ;
  assign n1412 = n1411 ^ n1391 ;
  assign n1424 = n1423 ^ n1412 ;
  assign n1405 = n1370 ^ n1369 ;
  assign n1406 = n1376 & ~n1405 ;
  assign n1407 = n1406 ^ n1375 ;
  assign n1402 = n1372 ^ n1371 ;
  assign n1403 = n1374 & ~n1402 ;
  assign n1404 = n1403 ^ n1373 ;
  assign n1408 = n1407 ^ n1404 ;
  assign n1399 = n1366 ^ n1365 ;
  assign n1400 = n1368 & ~n1399 ;
  assign n1401 = n1400 ^ n1367 ;
  assign n1409 = n1408 ^ n1401 ;
  assign n1434 = n1423 ^ n1409 ;
  assign n1435 = n1424 & ~n1434 ;
  assign n1436 = n1435 ^ n1412 ;
  assign n1440 = n1439 ^ n1436 ;
  assign n1431 = n1404 ^ n1401 ;
  assign n1432 = n1408 & ~n1431 ;
  assign n1433 = n1432 ^ n1407 ;
  assign n1447 = n1436 ^ n1433 ;
  assign n1448 = n1440 & ~n1447 ;
  assign n1449 = n1448 ^ n1439 ;
  assign n1441 = n1440 ^ n1433 ;
  assign n1425 = n1424 ^ n1409 ;
  assign n1393 = n1392 ^ n1377 ;
  assign n1364 = x257 ^ x161 ;
  assign n1394 = n1393 ^ n1364 ;
  assign n1334 = x261 ^ x165 ;
  assign n1333 = x260 ^ x164 ;
  assign n1335 = n1334 ^ n1333 ;
  assign n1332 = x262 ^ x166 ;
  assign n1336 = n1335 ^ n1332 ;
  assign n1328 = x264 ^ x168 ;
  assign n1327 = x263 ^ x167 ;
  assign n1329 = n1328 ^ n1327 ;
  assign n1326 = x265 ^ x169 ;
  assign n1330 = n1329 ^ n1326 ;
  assign n1325 = x259 ^ x163 ;
  assign n1331 = n1330 ^ n1325 ;
  assign n1337 = n1336 ^ n1331 ;
  assign n1323 = x258 ^ x162 ;
  assign n1309 = x268 ^ x172 ;
  assign n1308 = x267 ^ x171 ;
  assign n1310 = n1309 ^ n1308 ;
  assign n1307 = x269 ^ x173 ;
  assign n1311 = n1310 ^ n1307 ;
  assign n1300 = x272 ^ x176 ;
  assign n1298 = x271 ^ x175 ;
  assign n1297 = x270 ^ x174 ;
  assign n1299 = n1298 ^ n1297 ;
  assign n1305 = n1300 ^ n1299 ;
  assign n1304 = x266 ^ x170 ;
  assign n1306 = n1305 ^ n1304 ;
  assign n1322 = n1311 ^ n1306 ;
  assign n1324 = n1323 ^ n1322 ;
  assign n1395 = n1337 ^ n1324 ;
  assign n1396 = n1395 ^ n1364 ;
  assign n1397 = n1394 & ~n1396 ;
  assign n1398 = n1397 ^ n1393 ;
  assign n1426 = n1425 ^ n1398 ;
  assign n1349 = n1327 ^ n1326 ;
  assign n1350 = n1329 & ~n1349 ;
  assign n1351 = n1350 ^ n1328 ;
  assign n1346 = n1336 ^ n1330 ;
  assign n1347 = ~n1331 & n1346 ;
  assign n1348 = n1347 ^ n1336 ;
  assign n1352 = n1351 ^ n1348 ;
  assign n1343 = n1333 ^ n1332 ;
  assign n1344 = n1335 & ~n1343 ;
  assign n1345 = n1344 ^ n1334 ;
  assign n1353 = n1352 ^ n1345 ;
  assign n1316 = n1308 ^ n1307 ;
  assign n1317 = n1310 & ~n1316 ;
  assign n1318 = n1317 ^ n1309 ;
  assign n1312 = n1311 ^ n1304 ;
  assign n1313 = n1306 & ~n1312 ;
  assign n1314 = n1313 ^ n1305 ;
  assign n1301 = n1300 ^ n1297 ;
  assign n1302 = n1299 & ~n1301 ;
  assign n1303 = n1302 ^ n1298 ;
  assign n1315 = n1314 ^ n1303 ;
  assign n1341 = n1318 ^ n1315 ;
  assign n1338 = n1337 ^ n1322 ;
  assign n1339 = n1324 & ~n1338 ;
  assign n1340 = n1339 ^ n1323 ;
  assign n1342 = n1341 ^ n1340 ;
  assign n1427 = n1353 ^ n1342 ;
  assign n1428 = n1427 ^ n1425 ;
  assign n1429 = n1426 & ~n1428 ;
  assign n1430 = n1429 ^ n1398 ;
  assign n1442 = n1441 ^ n1430 ;
  assign n1358 = n1348 ^ n1345 ;
  assign n1359 = n1352 & ~n1358 ;
  assign n1360 = n1359 ^ n1351 ;
  assign n1354 = n1353 ^ n1341 ;
  assign n1355 = n1342 & ~n1354 ;
  assign n1356 = n1355 ^ n1340 ;
  assign n1319 = n1318 ^ n1303 ;
  assign n1320 = n1315 & ~n1319 ;
  assign n1321 = n1320 ^ n1314 ;
  assign n1357 = n1356 ^ n1321 ;
  assign n1443 = n1360 ^ n1357 ;
  assign n1444 = n1443 ^ n1430 ;
  assign n1445 = n1442 & ~n1444 ;
  assign n1446 = n1445 ^ n1441 ;
  assign n1450 = n1449 ^ n1446 ;
  assign n1361 = n1360 ^ n1321 ;
  assign n1362 = n1357 & ~n1361 ;
  assign n1363 = n1362 ^ n1356 ;
  assign n1451 = n1450 ^ n1363 ;
  assign n1452 = n1427 ^ n1426 ;
  assign n1453 = n1395 ^ n1394 ;
  assign n1454 = x256 ^ x160 ;
  assign n1455 = n1453 & n1454 ;
  assign n1456 = n1452 & n1455 ;
  assign n1457 = n1443 ^ n1442 ;
  assign n1458 = n1456 & n1457 ;
  assign n1459 = n1451 & n1458 ;
  assign n1460 = n1449 ^ n1363 ;
  assign n1461 = ~n1450 & n1460 ;
  assign n1462 = n1461 ^ n1363 ;
  assign n1463 = n1459 & n1462 ;
  assign n1464 = n1294 & ~n1463 ;
  assign n1465 = n1464 ^ n1294 ;
  assign n1295 = n1294 ^ n1292 ;
  assign n1296 = n1295 ^ n1123 ;
  assign n1467 = n1465 ^ n1296 ;
  assign n1466 = n1296 & n1465 ;
  assign n1468 = n1467 ^ n1466 ;
  assign n1469 = n1468 ^ n1465 ;
  assign n1470 = ~n956 & ~n1469 ;
  assign n1471 = n1470 ^ n1469 ;
  assign n1472 = n1468 ^ n1296 ;
  assign n1473 = ~n1471 & ~n1472 ;
  assign n1474 = n1473 ^ n1471 ;
  assign n1642 = n1474 ^ n1472 ;
  assign n1643 = n1642 ^ n1471 ;
  assign n1644 = ~n1641 & n1643 ;
  assign n1645 = n1644 ^ n1643 ;
  assign n1649 = n1645 ^ n1474 ;
  assign n712 = x285 ^ x93 ;
  assign n711 = x286 ^ x94 ;
  assign n713 = n712 ^ n711 ;
  assign n710 = x287 ^ x95 ;
  assign n745 = n711 ^ n710 ;
  assign n746 = n713 & ~n745 ;
  assign n747 = n746 ^ n712 ;
  assign n715 = x281 ^ x89 ;
  assign n714 = n713 ^ n710 ;
  assign n716 = n715 ^ n714 ;
  assign n707 = x283 ^ x91 ;
  assign n706 = x282 ^ x90 ;
  assign n708 = n707 ^ n706 ;
  assign n705 = x284 ^ x92 ;
  assign n709 = n708 ^ n705 ;
  assign n742 = n714 ^ n709 ;
  assign n743 = n716 & ~n742 ;
  assign n744 = n743 ^ n715 ;
  assign n748 = n747 ^ n744 ;
  assign n739 = n706 ^ n705 ;
  assign n740 = n708 & ~n739 ;
  assign n741 = n740 ^ n707 ;
  assign n763 = n744 ^ n741 ;
  assign n764 = n748 & ~n763 ;
  assign n765 = n764 ^ n747 ;
  assign n749 = n748 ^ n741 ;
  assign n717 = n716 ^ n709 ;
  assign n704 = x273 ^ x81 ;
  assign n718 = n717 ^ n704 ;
  assign n699 = x279 ^ x87 ;
  assign n698 = x278 ^ x86 ;
  assign n700 = n699 ^ n698 ;
  assign n697 = x280 ^ x88 ;
  assign n701 = n700 ^ n697 ;
  assign n696 = x274 ^ x82 ;
  assign n702 = n701 ^ n696 ;
  assign n693 = x276 ^ x84 ;
  assign n692 = x275 ^ x83 ;
  assign n694 = n693 ^ n692 ;
  assign n691 = x277 ^ x85 ;
  assign n695 = n694 ^ n691 ;
  assign n703 = n702 ^ n695 ;
  assign n736 = n704 ^ n703 ;
  assign n737 = n718 & ~n736 ;
  assign n738 = n737 ^ n717 ;
  assign n750 = n749 ^ n738 ;
  assign n731 = n696 ^ n695 ;
  assign n732 = n702 & ~n731 ;
  assign n733 = n732 ^ n701 ;
  assign n728 = n698 ^ n697 ;
  assign n729 = n700 & ~n728 ;
  assign n730 = n729 ^ n699 ;
  assign n734 = n733 ^ n730 ;
  assign n725 = n692 ^ n691 ;
  assign n726 = n694 & ~n725 ;
  assign n727 = n726 ^ n693 ;
  assign n735 = n734 ^ n727 ;
  assign n760 = n749 ^ n735 ;
  assign n761 = n750 & ~n760 ;
  assign n762 = n761 ^ n738 ;
  assign n766 = n765 ^ n762 ;
  assign n757 = n730 ^ n727 ;
  assign n758 = n734 & ~n757 ;
  assign n759 = n758 ^ n733 ;
  assign n773 = n762 ^ n759 ;
  assign n774 = n766 & ~n773 ;
  assign n775 = n774 ^ n765 ;
  assign n767 = n766 ^ n759 ;
  assign n751 = n750 ^ n735 ;
  assign n719 = n718 ^ n703 ;
  assign n690 = x257 ^ x65 ;
  assign n720 = n719 ^ n690 ;
  assign n660 = x261 ^ x69 ;
  assign n659 = x260 ^ x68 ;
  assign n661 = n660 ^ n659 ;
  assign n658 = x262 ^ x70 ;
  assign n662 = n661 ^ n658 ;
  assign n654 = x264 ^ x72 ;
  assign n653 = x263 ^ x71 ;
  assign n655 = n654 ^ n653 ;
  assign n652 = x265 ^ x73 ;
  assign n656 = n655 ^ n652 ;
  assign n651 = x259 ^ x67 ;
  assign n657 = n656 ^ n651 ;
  assign n663 = n662 ^ n657 ;
  assign n649 = x258 ^ x66 ;
  assign n635 = x268 ^ x76 ;
  assign n634 = x267 ^ x75 ;
  assign n636 = n635 ^ n634 ;
  assign n633 = x269 ^ x77 ;
  assign n637 = n636 ^ n633 ;
  assign n626 = x272 ^ x80 ;
  assign n624 = x271 ^ x79 ;
  assign n623 = x270 ^ x78 ;
  assign n625 = n624 ^ n623 ;
  assign n631 = n626 ^ n625 ;
  assign n630 = x266 ^ x74 ;
  assign n632 = n631 ^ n630 ;
  assign n648 = n637 ^ n632 ;
  assign n650 = n649 ^ n648 ;
  assign n721 = n663 ^ n650 ;
  assign n722 = n721 ^ n690 ;
  assign n723 = n720 & ~n722 ;
  assign n724 = n723 ^ n719 ;
  assign n752 = n751 ^ n724 ;
  assign n675 = n653 ^ n652 ;
  assign n676 = n655 & ~n675 ;
  assign n677 = n676 ^ n654 ;
  assign n672 = n662 ^ n656 ;
  assign n673 = ~n657 & n672 ;
  assign n674 = n673 ^ n662 ;
  assign n678 = n677 ^ n674 ;
  assign n669 = n659 ^ n658 ;
  assign n670 = n661 & ~n669 ;
  assign n671 = n670 ^ n660 ;
  assign n679 = n678 ^ n671 ;
  assign n642 = n634 ^ n633 ;
  assign n643 = n636 & ~n642 ;
  assign n644 = n643 ^ n635 ;
  assign n638 = n637 ^ n630 ;
  assign n639 = n632 & ~n638 ;
  assign n640 = n639 ^ n631 ;
  assign n627 = n626 ^ n623 ;
  assign n628 = n625 & ~n627 ;
  assign n629 = n628 ^ n624 ;
  assign n641 = n640 ^ n629 ;
  assign n667 = n644 ^ n641 ;
  assign n664 = n663 ^ n648 ;
  assign n665 = n650 & ~n664 ;
  assign n666 = n665 ^ n649 ;
  assign n668 = n667 ^ n666 ;
  assign n753 = n679 ^ n668 ;
  assign n754 = n753 ^ n751 ;
  assign n755 = n752 & ~n754 ;
  assign n756 = n755 ^ n724 ;
  assign n768 = n767 ^ n756 ;
  assign n684 = n674 ^ n671 ;
  assign n685 = n678 & ~n684 ;
  assign n686 = n685 ^ n677 ;
  assign n680 = n679 ^ n667 ;
  assign n681 = n668 & ~n680 ;
  assign n682 = n681 ^ n666 ;
  assign n645 = n644 ^ n629 ;
  assign n646 = n641 & ~n645 ;
  assign n647 = n646 ^ n640 ;
  assign n683 = n682 ^ n647 ;
  assign n769 = n686 ^ n683 ;
  assign n770 = n769 ^ n756 ;
  assign n771 = n768 & ~n770 ;
  assign n772 = n771 ^ n767 ;
  assign n776 = n775 ^ n772 ;
  assign n687 = n686 ^ n647 ;
  assign n688 = n683 & ~n687 ;
  assign n689 = n688 ^ n682 ;
  assign n777 = n776 ^ n689 ;
  assign n778 = n753 ^ n752 ;
  assign n779 = n721 ^ n720 ;
  assign n780 = x256 ^ x64 ;
  assign n781 = n779 & n780 ;
  assign n782 = n778 & n781 ;
  assign n783 = n769 ^ n768 ;
  assign n784 = n782 & n783 ;
  assign n785 = n777 & n784 ;
  assign n786 = n775 ^ n689 ;
  assign n787 = ~n776 & n786 ;
  assign n788 = n787 ^ n689 ;
  assign n789 = n785 & n788 ;
  assign n1646 = n1474 & ~n1645 ;
  assign n1647 = ~n789 & ~n1646 ;
  assign n1652 = n1649 ^ n1647 ;
  assign n1648 = n1647 ^ n1646 ;
  assign n1650 = n1649 ^ n1646 ;
  assign n1651 = ~n1648 & ~n1650 ;
  assign n1653 = n1652 ^ n1651 ;
  assign n1654 = n1653 ^ n1648 ;
  assign n1655 = ~n622 & n1654 ;
  assign n1656 = n1655 ^ n1654 ;
  assign n1657 = n1653 ^ n1650 ;
  assign n1658 = n1656 & n1657 ;
  assign n1659 = n1658 ^ n1656 ;
  assign n1660 = n1659 ^ n1657 ;
  assign n1661 = n1660 ^ n1656 ;
  assign n1662 = ~n455 & ~n1661 ;
  assign n1663 = n1662 ^ n1661 ;
  assign n1664 = n1663 ^ n1659 ;
  assign n1667 = n1122 ^ n1119 ;
  assign n1668 = n1667 ^ n1291 ;
  assign n1669 = n1291 & ~n1667 ;
  assign n1670 = n1669 ^ n1293 ;
  assign n1671 = n1669 ^ n1668 ;
  assign n1673 = n1118 ^ n1107 ;
  assign n1672 = n1288 ^ n1287 ;
  assign n1674 = n1673 ^ n1672 ;
  assign n1676 = n1286 ^ n1281 ;
  assign n1675 = n1106 ^ n1101 ;
  assign n1677 = n1676 ^ n1675 ;
  assign n1681 = n1105 ^ n1102 ;
  assign n1678 = n1284 ^ n1283 ;
  assign n1679 = n1104 ^ n1103 ;
  assign n1680 = n1678 & ~n1679 ;
  assign n1682 = n1681 ^ n1680 ;
  assign n1683 = n1285 ^ n1282 ;
  assign n1684 = n1683 ^ n1680 ;
  assign n1685 = ~n1682 & ~n1684 ;
  assign n1686 = n1685 ^ n1681 ;
  assign n1687 = n1686 ^ n1676 ;
  assign n1688 = ~n1677 & n1687 ;
  assign n1689 = n1688 ^ n1675 ;
  assign n1690 = n1689 ^ n1673 ;
  assign n1691 = ~n1674 & n1690 ;
  assign n1692 = n1691 ^ n1673 ;
  assign n1693 = ~n1671 & ~n1692 ;
  assign n1694 = ~n1670 & ~n1693 ;
  assign n1695 = n1295 & ~n1694 ;
  assign n1696 = n1668 & ~n1695 ;
  assign n1741 = n1696 ^ n1667 ;
  assign n1666 = n1291 ^ n1123 ;
  assign n1697 = n1696 ^ n1666 ;
  assign n1698 = n1697 ^ n1123 ;
  assign n1665 = n1462 ^ n1459 ;
  assign n1699 = n1698 ^ n1665 ;
  assign n1700 = n1455 ^ n1452 ;
  assign n1701 = n1683 ^ n1681 ;
  assign n1702 = n1695 & n1701 ;
  assign n1703 = n1702 ^ n1701 ;
  assign n1704 = n1703 ^ n1683 ;
  assign n1705 = n1700 & ~n1704 ;
  assign n1706 = n1454 ^ n1453 ;
  assign n1707 = n1679 ^ n1678 ;
  assign n1708 = n1695 & n1707 ;
  assign n1709 = n1708 ^ n1707 ;
  assign n1710 = n1709 ^ n1678 ;
  assign n1711 = n1706 & ~n1710 ;
  assign n1712 = ~n1705 & ~n1711 ;
  assign n1713 = ~n1452 & n1704 ;
  assign n1715 = n1677 & ~n1695 ;
  assign n1716 = n1715 ^ n1677 ;
  assign n1717 = n1716 ^ n1675 ;
  assign n1714 = n1457 ^ n1456 ;
  assign n1719 = n1717 ^ n1714 ;
  assign n1718 = n1714 & ~n1717 ;
  assign n1720 = n1719 ^ n1718 ;
  assign n1721 = ~n1713 & ~n1720 ;
  assign n1722 = ~n1712 & n1721 ;
  assign n1724 = n1674 & ~n1695 ;
  assign n1725 = n1724 ^ n1672 ;
  assign n1723 = n1458 ^ n1451 ;
  assign n1727 = n1725 ^ n1723 ;
  assign n1726 = ~n1723 & n1725 ;
  assign n1728 = n1727 ^ n1726 ;
  assign n1729 = ~n1718 & ~n1728 ;
  assign n1730 = ~n1722 & n1729 ;
  assign n1731 = ~n1665 & n1698 ;
  assign n1732 = n1731 ^ n1464 ;
  assign n1733 = ~n1726 & ~n1732 ;
  assign n1734 = ~n1730 & n1733 ;
  assign n1735 = n1699 ^ n1463 ;
  assign n1736 = n1735 ^ n1731 ;
  assign n1737 = ~n1294 & n1736 ;
  assign n1738 = ~n1734 & ~n1737 ;
  assign n1739 = n1699 & ~n1738 ;
  assign n1740 = n1739 ^ n1665 ;
  assign n1742 = n1741 ^ n1740 ;
  assign n1743 = ~n1740 & n1741 ;
  assign n1744 = n1743 ^ n1468 ;
  assign n1745 = n1743 ^ n1742 ;
  assign n1747 = n1727 & ~n1738 ;
  assign n1748 = n1747 ^ n1723 ;
  assign n1746 = n1724 ^ n1673 ;
  assign n1749 = n1748 ^ n1746 ;
  assign n1751 = n1719 & ~n1738 ;
  assign n1752 = n1751 ^ n1714 ;
  assign n1750 = n1715 ^ n1675 ;
  assign n1753 = n1752 ^ n1750 ;
  assign n1757 = n1702 ^ n1683 ;
  assign n1754 = n1704 ^ n1700 ;
  assign n1755 = ~n1738 & n1754 ;
  assign n1756 = n1755 ^ n1700 ;
  assign n1758 = n1757 ^ n1756 ;
  assign n1759 = n1710 ^ n1706 ;
  assign n1760 = ~n1738 & n1759 ;
  assign n1761 = n1760 ^ n1706 ;
  assign n1762 = n1708 ^ n1678 ;
  assign n1763 = n1761 & ~n1762 ;
  assign n1764 = n1763 ^ n1757 ;
  assign n1765 = ~n1758 & ~n1764 ;
  assign n1766 = n1765 ^ n1757 ;
  assign n1767 = n1766 ^ n1752 ;
  assign n1768 = ~n1753 & ~n1767 ;
  assign n1769 = n1768 ^ n1752 ;
  assign n1770 = n1769 ^ n1748 ;
  assign n1771 = ~n1749 & n1770 ;
  assign n1772 = n1771 ^ n1748 ;
  assign n1773 = ~n1745 & ~n1772 ;
  assign n1774 = n1744 & ~n1773 ;
  assign n1775 = ~n1466 & ~n1774 ;
  assign n1776 = n1742 & n1775 ;
  assign n1819 = n1776 ^ n1741 ;
  assign n1778 = n955 ^ n952 ;
  assign n1777 = n1776 ^ n1740 ;
  assign n1779 = n1778 ^ n1777 ;
  assign n1780 = n947 ^ n946 ;
  assign n1781 = n1762 ^ n1761 ;
  assign n1782 = ~n1775 & n1781 ;
  assign n1783 = n1782 ^ n1781 ;
  assign n1784 = n1783 ^ n1761 ;
  assign n1785 = n1780 & ~n1784 ;
  assign n1786 = n945 & n1785 ;
  assign n1787 = n1758 & n1775 ;
  assign n1788 = n1787 ^ n1756 ;
  assign n1789 = ~n1786 & n1788 ;
  assign n1790 = n948 ^ n945 ;
  assign n1791 = ~n1785 & ~n1790 ;
  assign n1793 = n1753 & n1775 ;
  assign n1794 = n1793 ^ n1753 ;
  assign n1795 = n1794 ^ n1750 ;
  assign n1792 = n950 ^ n949 ;
  assign n1797 = n1795 ^ n1792 ;
  assign n1796 = n1792 & ~n1795 ;
  assign n1798 = n1797 ^ n1796 ;
  assign n1799 = ~n1791 & ~n1798 ;
  assign n1800 = ~n1789 & n1799 ;
  assign n1802 = n1749 & n1775 ;
  assign n1803 = n1802 ^ n1748 ;
  assign n1801 = n951 ^ n944 ;
  assign n1805 = n1803 ^ n1801 ;
  assign n1804 = ~n1801 & n1803 ;
  assign n1806 = n1805 ^ n1804 ;
  assign n1807 = ~n1796 & ~n1806 ;
  assign n1808 = ~n1800 & n1807 ;
  assign n1809 = n1777 & ~n1778 ;
  assign n1810 = ~n1470 & ~n1804 ;
  assign n1811 = ~n1809 & n1810 ;
  assign n1812 = ~n1808 & n1811 ;
  assign n1813 = n1779 ^ n956 ;
  assign n1814 = n1813 ^ n1809 ;
  assign n1815 = n1469 & n1814 ;
  assign n1816 = ~n1812 & ~n1815 ;
  assign n1817 = n1779 & ~n1816 ;
  assign n1818 = n1817 ^ n1778 ;
  assign n1820 = n1819 ^ n1818 ;
  assign n1821 = n1472 ^ n1471 ;
  assign n1823 = n1805 & ~n1816 ;
  assign n1824 = n1823 ^ n1801 ;
  assign n1822 = n1802 ^ n1746 ;
  assign n1825 = n1824 ^ n1822 ;
  assign n1827 = n1797 & ~n1816 ;
  assign n1828 = n1827 ^ n1792 ;
  assign n1826 = n1793 ^ n1750 ;
  assign n1829 = n1828 ^ n1826 ;
  assign n1832 = n1790 ^ n1788 ;
  assign n1833 = n1816 & n1832 ;
  assign n1834 = n1833 ^ n1788 ;
  assign n1830 = n1788 ^ n1757 ;
  assign n1831 = n1830 ^ n1756 ;
  assign n1835 = n1834 ^ n1831 ;
  assign n1836 = n1782 ^ n1761 ;
  assign n1837 = n1784 ^ n1780 ;
  assign n1838 = ~n1816 & n1837 ;
  assign n1839 = n1838 ^ n1780 ;
  assign n1840 = ~n1836 & n1839 ;
  assign n1841 = n1840 ^ n1834 ;
  assign n1842 = ~n1835 & n1841 ;
  assign n1843 = n1842 ^ n1834 ;
  assign n1844 = n1843 ^ n1828 ;
  assign n1845 = ~n1829 & n1844 ;
  assign n1846 = n1845 ^ n1828 ;
  assign n1847 = n1846 ^ n1824 ;
  assign n1848 = ~n1825 & n1847 ;
  assign n1849 = n1848 ^ n1824 ;
  assign n1850 = n1849 ^ n1819 ;
  assign n1851 = ~n1820 & ~n1850 ;
  assign n1852 = n1851 ^ n1819 ;
  assign n1853 = n1852 ^ n1472 ;
  assign n1854 = n1821 & ~n1853 ;
  assign n1855 = n1854 ^ n1471 ;
  assign n1856 = n1820 & n1855 ;
  assign n1901 = n1856 ^ n1819 ;
  assign n1858 = n1640 ^ n1637 ;
  assign n1857 = n1856 ^ n1818 ;
  assign n1859 = n1858 ^ n1857 ;
  assign n1860 = n1633 ^ n1630 ;
  assign n1861 = n1835 & n1855 ;
  assign n1862 = n1861 ^ n1831 ;
  assign n1863 = n1862 ^ n1834 ;
  assign n1864 = n1863 ^ n1831 ;
  assign n1865 = n1860 & ~n1864 ;
  assign n1866 = n1632 ^ n1631 ;
  assign n1867 = n1839 ^ n1836 ;
  assign n1868 = n1855 & n1867 ;
  assign n1869 = n1868 ^ n1867 ;
  assign n1870 = n1869 ^ n1836 ;
  assign n1871 = n1866 & ~n1870 ;
  assign n1872 = ~n1865 & ~n1871 ;
  assign n1873 = ~n1630 & n1864 ;
  assign n1875 = n1829 & n1855 ;
  assign n1876 = n1875 ^ n1829 ;
  assign n1877 = n1876 ^ n1826 ;
  assign n1874 = n1635 ^ n1634 ;
  assign n1879 = n1877 ^ n1874 ;
  assign n1878 = n1874 & ~n1877 ;
  assign n1880 = n1879 ^ n1878 ;
  assign n1881 = ~n1873 & ~n1880 ;
  assign n1882 = ~n1872 & n1881 ;
  assign n1884 = n1825 & n1855 ;
  assign n1885 = n1884 ^ n1824 ;
  assign n1883 = n1636 ^ n1629 ;
  assign n1887 = n1885 ^ n1883 ;
  assign n1886 = ~n1883 & n1885 ;
  assign n1888 = n1887 ^ n1886 ;
  assign n1889 = ~n1878 & ~n1888 ;
  assign n1890 = ~n1882 & n1889 ;
  assign n1891 = n1857 & ~n1858 ;
  assign n1892 = ~n1644 & ~n1891 ;
  assign n1893 = ~n1886 & n1892 ;
  assign n1894 = ~n1890 & n1893 ;
  assign n1895 = n1859 ^ n1641 ;
  assign n1896 = n1895 ^ n1891 ;
  assign n1897 = ~n1643 & n1896 ;
  assign n1898 = ~n1894 & ~n1897 ;
  assign n1899 = n1859 & ~n1898 ;
  assign n1900 = n1899 ^ n1858 ;
  assign n1902 = n1901 ^ n1900 ;
  assign n1903 = n1900 & ~n1901 ;
  assign n1904 = n1903 ^ n1902 ;
  assign n1905 = n1904 ^ n1474 ;
  assign n1906 = n1905 ^ n1474 ;
  assign n1908 = n1887 & ~n1898 ;
  assign n1909 = n1908 ^ n1883 ;
  assign n1907 = n1884 ^ n1822 ;
  assign n1910 = n1909 ^ n1907 ;
  assign n1912 = n1879 & ~n1898 ;
  assign n1913 = n1912 ^ n1874 ;
  assign n1911 = n1875 ^ n1826 ;
  assign n1914 = n1913 ^ n1911 ;
  assign n1915 = n1864 ^ n1860 ;
  assign n1916 = ~n1898 & n1915 ;
  assign n1917 = n1916 ^ n1860 ;
  assign n1918 = n1917 ^ n1862 ;
  assign n1919 = n1868 ^ n1836 ;
  assign n1920 = n1870 ^ n1866 ;
  assign n1921 = ~n1898 & n1920 ;
  assign n1922 = n1921 ^ n1866 ;
  assign n1923 = ~n1919 & n1922 ;
  assign n1924 = n1923 ^ n1862 ;
  assign n1925 = ~n1918 & ~n1924 ;
  assign n1926 = n1925 ^ n1862 ;
  assign n1927 = n1926 ^ n1913 ;
  assign n1928 = ~n1914 & ~n1927 ;
  assign n1929 = n1928 ^ n1913 ;
  assign n1930 = n1929 ^ n1907 ;
  assign n1931 = ~n1910 & ~n1930 ;
  assign n1932 = n1931 ^ n1907 ;
  assign n1933 = ~n1903 & n1932 ;
  assign n1934 = n1933 ^ n1474 ;
  assign n1935 = n1934 ^ n1474 ;
  assign n1936 = ~n1906 & ~n1935 ;
  assign n1937 = n1936 ^ n1474 ;
  assign n1938 = n1649 & ~n1937 ;
  assign n1939 = n1938 ^ n1645 ;
  assign n1940 = n1902 & ~n1939 ;
  assign n1984 = n1940 ^ n1901 ;
  assign n1942 = n788 ^ n785 ;
  assign n1941 = n1940 ^ n1900 ;
  assign n1943 = n1942 ^ n1941 ;
  assign n1944 = n781 ^ n778 ;
  assign n1945 = n1918 & n1939 ;
  assign n1946 = n1945 ^ n1918 ;
  assign n1947 = n1946 ^ n1917 ;
  assign n1948 = n1944 & ~n1947 ;
  assign n1949 = n780 ^ n779 ;
  assign n1950 = n1922 ^ n1919 ;
  assign n1951 = ~n1939 & n1950 ;
  assign n1952 = n1951 ^ n1950 ;
  assign n1953 = n1952 ^ n1919 ;
  assign n1954 = n1949 & ~n1953 ;
  assign n1955 = ~n1948 & ~n1954 ;
  assign n1956 = ~n778 & n1947 ;
  assign n1958 = n1914 & ~n1939 ;
  assign n1959 = n1958 ^ n1914 ;
  assign n1960 = n1959 ^ n1911 ;
  assign n1957 = n783 ^ n782 ;
  assign n1962 = n1960 ^ n1957 ;
  assign n1961 = n1957 & ~n1960 ;
  assign n1963 = n1962 ^ n1961 ;
  assign n1964 = ~n1956 & ~n1963 ;
  assign n1965 = ~n1955 & n1964 ;
  assign n1967 = n1910 & ~n1939 ;
  assign n1968 = n1967 ^ n1909 ;
  assign n1966 = n784 ^ n777 ;
  assign n1970 = n1968 ^ n1966 ;
  assign n1969 = ~n1966 & n1968 ;
  assign n1971 = n1970 ^ n1969 ;
  assign n1972 = ~n1961 & ~n1971 ;
  assign n1973 = ~n1965 & n1972 ;
  assign n1974 = n1941 & ~n1942 ;
  assign n1975 = ~n1647 & ~n1974 ;
  assign n1976 = ~n1969 & n1975 ;
  assign n1977 = ~n1973 & n1976 ;
  assign n1978 = n1943 ^ n789 ;
  assign n1979 = n1978 ^ n1974 ;
  assign n1980 = n1646 & n1979 ;
  assign n1981 = ~n1977 & ~n1980 ;
  assign n1982 = n1943 & ~n1981 ;
  assign n1983 = n1982 ^ n1942 ;
  assign n1985 = n1984 ^ n1983 ;
  assign n1987 = n1970 & ~n1981 ;
  assign n1988 = n1987 ^ n1966 ;
  assign n1986 = n1967 ^ n1907 ;
  assign n1989 = n1988 ^ n1986 ;
  assign n1991 = n1962 & ~n1981 ;
  assign n1992 = n1991 ^ n1957 ;
  assign n1990 = n1958 ^ n1911 ;
  assign n1993 = n1992 ^ n1990 ;
  assign n1997 = n1945 ^ n1917 ;
  assign n1994 = n1947 ^ n1944 ;
  assign n1995 = ~n1981 & n1994 ;
  assign n1996 = n1995 ^ n1944 ;
  assign n1998 = n1997 ^ n1996 ;
  assign n1999 = n1951 ^ n1919 ;
  assign n2000 = n1953 ^ n1949 ;
  assign n2001 = ~n1981 & n2000 ;
  assign n2002 = n2001 ^ n1949 ;
  assign n2003 = ~n1999 & n2002 ;
  assign n2004 = n2003 ^ n1997 ;
  assign n2005 = ~n1998 & ~n2004 ;
  assign n2006 = n2005 ^ n1997 ;
  assign n2007 = n2006 ^ n1992 ;
  assign n2008 = ~n1993 & ~n2007 ;
  assign n2009 = n2008 ^ n1992 ;
  assign n2010 = n2009 ^ n1988 ;
  assign n2011 = ~n1989 & n2010 ;
  assign n2012 = n2011 ^ n1988 ;
  assign n2013 = n2012 ^ n1984 ;
  assign n2014 = ~n1985 & ~n2013 ;
  assign n2015 = n2014 ^ n1984 ;
  assign n2016 = n2015 ^ n1650 ;
  assign n2017 = ~n1652 & n2016 ;
  assign n2018 = n2017 ^ n2015 ;
  assign n2019 = n1985 & n2018 ;
  assign n2064 = n2019 ^ n1984 ;
  assign n2021 = n621 ^ n618 ;
  assign n2020 = n2019 ^ n1983 ;
  assign n2022 = n2021 ^ n2020 ;
  assign n2023 = n614 ^ n611 ;
  assign n2024 = n1998 & ~n2018 ;
  assign n2025 = n2024 ^ n1996 ;
  assign n2026 = n2025 ^ n1997 ;
  assign n2027 = n2026 ^ n1996 ;
  assign n2028 = n2023 & ~n2027 ;
  assign n2029 = n613 ^ n612 ;
  assign n2030 = n2002 ^ n1999 ;
  assign n2031 = n2018 & n2030 ;
  assign n2032 = n2031 ^ n2030 ;
  assign n2033 = n2032 ^ n1999 ;
  assign n2034 = n2029 & ~n2033 ;
  assign n2035 = ~n2028 & ~n2034 ;
  assign n2036 = ~n611 & n2027 ;
  assign n2038 = n1993 & n2018 ;
  assign n2039 = n2038 ^ n1993 ;
  assign n2040 = n2039 ^ n1990 ;
  assign n2037 = n616 ^ n615 ;
  assign n2042 = n2040 ^ n2037 ;
  assign n2041 = n2037 & ~n2040 ;
  assign n2043 = n2042 ^ n2041 ;
  assign n2044 = ~n2036 & ~n2043 ;
  assign n2045 = ~n2035 & n2044 ;
  assign n2047 = n1989 & n2018 ;
  assign n2048 = n2047 ^ n1988 ;
  assign n2046 = n617 ^ n610 ;
  assign n2050 = n2048 ^ n2046 ;
  assign n2049 = ~n2046 & n2048 ;
  assign n2051 = n2050 ^ n2049 ;
  assign n2052 = ~n2041 & ~n2051 ;
  assign n2053 = ~n2045 & n2052 ;
  assign n2054 = n2020 & ~n2021 ;
  assign n2055 = ~n1655 & ~n2054 ;
  assign n2056 = ~n2049 & n2055 ;
  assign n2057 = ~n2053 & n2056 ;
  assign n2058 = n2022 ^ n622 ;
  assign n2059 = n2058 ^ n2054 ;
  assign n2060 = ~n1654 & n2059 ;
  assign n2061 = ~n2057 & ~n2060 ;
  assign n2062 = n2022 & ~n2061 ;
  assign n2063 = n2062 ^ n2021 ;
  assign n2065 = n2064 ^ n2063 ;
  assign n2066 = n1657 ^ n1656 ;
  assign n2067 = ~n2063 & n2064 ;
  assign n2068 = n2067 ^ n2065 ;
  assign n2070 = n2050 & ~n2061 ;
  assign n2071 = n2070 ^ n2046 ;
  assign n2069 = n2047 ^ n1986 ;
  assign n2072 = n2071 ^ n2069 ;
  assign n2074 = n2042 & ~n2061 ;
  assign n2075 = n2074 ^ n2037 ;
  assign n2073 = n2038 ^ n1990 ;
  assign n2076 = n2075 ^ n2073 ;
  assign n2077 = n2027 ^ n2023 ;
  assign n2078 = ~n2061 & n2077 ;
  assign n2079 = n2078 ^ n2023 ;
  assign n2080 = n2079 ^ n2025 ;
  assign n2081 = n2033 ^ n2029 ;
  assign n2082 = ~n2061 & n2081 ;
  assign n2083 = n2082 ^ n2029 ;
  assign n2084 = n2031 ^ n1999 ;
  assign n2085 = n2083 & ~n2084 ;
  assign n2086 = n2085 ^ n2025 ;
  assign n2087 = ~n2080 & ~n2086 ;
  assign n2088 = n2087 ^ n2025 ;
  assign n2089 = n2088 ^ n2075 ;
  assign n2090 = ~n2076 & ~n2089 ;
  assign n2091 = n2090 ^ n2075 ;
  assign n2092 = n2091 ^ n2071 ;
  assign n2093 = ~n2072 & n2092 ;
  assign n2094 = n2093 ^ n2071 ;
  assign n2095 = ~n2068 & ~n2094 ;
  assign n2096 = n2095 ^ n1657 ;
  assign n2097 = n2096 ^ n1657 ;
  assign n2098 = ~n2067 & ~n2097 ;
  assign n2099 = n2098 ^ n1657 ;
  assign n2100 = n2066 & ~n2099 ;
  assign n2101 = n2100 ^ n1656 ;
  assign n2102 = n2065 & ~n2101 ;
  assign n2105 = n2102 ^ n2063 ;
  assign n2104 = n454 ^ n451 ;
  assign n2106 = n2105 ^ n2104 ;
  assign n2107 = n447 ^ n444 ;
  assign n2108 = n2080 & n2101 ;
  assign n2109 = n2108 ^ n2079 ;
  assign n2110 = n2109 ^ n2025 ;
  assign n2111 = n2110 ^ n2079 ;
  assign n2112 = n2107 & ~n2111 ;
  assign n2113 = n446 ^ n445 ;
  assign n2114 = n2084 ^ n2083 ;
  assign n2115 = n2101 & n2114 ;
  assign n2116 = n2115 ^ n2114 ;
  assign n2117 = n2116 ^ n2083 ;
  assign n2118 = n2113 & ~n2117 ;
  assign n2119 = ~n2112 & ~n2118 ;
  assign n2120 = ~n444 & n2111 ;
  assign n2122 = n2076 & ~n2101 ;
  assign n2123 = n2122 ^ n2076 ;
  assign n2124 = n2123 ^ n2073 ;
  assign n2121 = n449 ^ n448 ;
  assign n2126 = n2124 ^ n2121 ;
  assign n2125 = n2121 & ~n2124 ;
  assign n2127 = n2126 ^ n2125 ;
  assign n2128 = ~n2120 & ~n2127 ;
  assign n2129 = ~n2119 & n2128 ;
  assign n2131 = n2072 & ~n2101 ;
  assign n2132 = n2131 ^ n2071 ;
  assign n2130 = n450 ^ n443 ;
  assign n2134 = n2132 ^ n2130 ;
  assign n2133 = ~n2130 & n2132 ;
  assign n2135 = n2134 ^ n2133 ;
  assign n2136 = ~n2125 & ~n2135 ;
  assign n2137 = ~n2129 & n2136 ;
  assign n2138 = ~n2104 & n2105 ;
  assign n2139 = ~n1662 & ~n2138 ;
  assign n2140 = ~n2133 & n2139 ;
  assign n2141 = ~n2137 & n2140 ;
  assign n2142 = n2106 ^ n455 ;
  assign n2143 = n2142 ^ n2138 ;
  assign n2144 = n1661 & n2143 ;
  assign n2145 = ~n2141 & ~n2144 ;
  assign n2146 = n2106 & n2145 ;
  assign n2147 = n2146 ^ n2105 ;
  assign n2103 = n2102 ^ n2064 ;
  assign n2148 = n2147 ^ n2103 ;
  assign n2150 = n2134 & n2145 ;
  assign n2151 = n2150 ^ n2132 ;
  assign n2149 = n2131 ^ n2069 ;
  assign n2152 = n2151 ^ n2149 ;
  assign n2154 = n2126 & ~n2145 ;
  assign n2155 = n2154 ^ n2121 ;
  assign n2153 = n2122 ^ n2073 ;
  assign n2156 = n2155 ^ n2153 ;
  assign n2162 = n2111 ^ n2107 ;
  assign n2163 = ~n2145 & n2162 ;
  assign n2164 = n2163 ^ n2107 ;
  assign n2157 = n2115 ^ n2083 ;
  assign n2158 = n2117 ^ n2113 ;
  assign n2159 = n2145 & n2158 ;
  assign n2160 = n2159 ^ n2117 ;
  assign n2161 = ~n2157 & n2160 ;
  assign n2165 = n2164 ^ n2161 ;
  assign n2166 = n2161 ^ n2109 ;
  assign n2167 = n2165 & ~n2166 ;
  assign n2168 = n2167 ^ n2161 ;
  assign n2169 = n2168 ^ n2155 ;
  assign n2170 = ~n2156 & n2169 ;
  assign n2171 = n2170 ^ n2155 ;
  assign n2172 = n2171 ^ n2149 ;
  assign n2173 = ~n2152 & ~n2172 ;
  assign n2174 = n2173 ^ n2149 ;
  assign n2175 = n2174 ^ n2103 ;
  assign n2176 = ~n2148 & ~n2175 ;
  assign n2177 = n2176 ^ n2147 ;
  assign n2178 = n2177 ^ n1659 ;
  assign n2179 = n1664 & n2178 ;
  assign n2180 = n2179 ^ n1663 ;
  assign n2181 = x224 ^ x192 ;
  assign n2182 = ~n1695 & n2181 ;
  assign n2185 = n2182 ^ x192 ;
  assign n2186 = n2185 ^ x160 ;
  assign n2187 = ~n1738 & n2186 ;
  assign n2188 = n2187 ^ x160 ;
  assign n2183 = n2182 ^ n2181 ;
  assign n2184 = n2183 ^ x192 ;
  assign n2189 = n2188 ^ n2184 ;
  assign n2190 = ~n1775 & n2189 ;
  assign n2193 = n2190 ^ n2184 ;
  assign n2194 = n2193 ^ x128 ;
  assign n2195 = ~n1816 & n2194 ;
  assign n2196 = n2195 ^ x128 ;
  assign n2191 = n2190 ^ n2189 ;
  assign n2192 = n2191 ^ n2184 ;
  assign n2197 = n2196 ^ n2192 ;
  assign n2198 = ~n1855 & n2197 ;
  assign n2201 = n2198 ^ n2192 ;
  assign n2202 = n2201 ^ x96 ;
  assign n2203 = ~n1898 & n2202 ;
  assign n2204 = n2203 ^ x96 ;
  assign n2199 = n2198 ^ n2197 ;
  assign n2200 = n2199 ^ n2192 ;
  assign n2205 = n2204 ^ n2200 ;
  assign n2206 = n1939 & n2205 ;
  assign n2209 = n2206 ^ n2200 ;
  assign n2210 = n2209 ^ x64 ;
  assign n2211 = ~n1981 & n2210 ;
  assign n2212 = n2211 ^ x64 ;
  assign n2207 = n2206 ^ n2205 ;
  assign n2208 = n2207 ^ n2200 ;
  assign n2213 = n2212 ^ n2208 ;
  assign n2214 = ~n2018 & n2213 ;
  assign n2217 = n2214 ^ n2208 ;
  assign n2218 = n2217 ^ x32 ;
  assign n2219 = ~n2061 & n2218 ;
  assign n2220 = n2219 ^ x32 ;
  assign n2215 = n2214 ^ n2213 ;
  assign n2216 = n2215 ^ n2208 ;
  assign n2221 = n2220 ^ n2216 ;
  assign n2222 = n2101 & n2221 ;
  assign n2225 = n2222 ^ n2216 ;
  assign n2226 = n2225 ^ x0 ;
  assign n2227 = ~n2145 & n2226 ;
  assign n2228 = n2227 ^ x0 ;
  assign n2223 = n2222 ^ n2221 ;
  assign n2224 = n2223 ^ n2216 ;
  assign n2229 = n2228 ^ n2224 ;
  assign n2230 = ~n2180 & n2229 ;
  assign n2231 = n2230 ^ n2229 ;
  assign n2232 = n2231 ^ n2224 ;
  assign n2233 = x225 ^ x193 ;
  assign n2234 = ~n1695 & n2233 ;
  assign n2237 = n2234 ^ x193 ;
  assign n2238 = n2237 ^ x161 ;
  assign n2239 = ~n1738 & n2238 ;
  assign n2240 = n2239 ^ x161 ;
  assign n2235 = n2234 ^ n2233 ;
  assign n2236 = n2235 ^ x193 ;
  assign n2241 = n2240 ^ n2236 ;
  assign n2242 = ~n1775 & n2241 ;
  assign n2245 = n2242 ^ n2236 ;
  assign n2246 = n2245 ^ x129 ;
  assign n2247 = ~n1816 & n2246 ;
  assign n2248 = n2247 ^ x129 ;
  assign n2243 = n2242 ^ n2241 ;
  assign n2244 = n2243 ^ n2236 ;
  assign n2249 = n2248 ^ n2244 ;
  assign n2250 = ~n1855 & n2249 ;
  assign n2253 = n2250 ^ n2244 ;
  assign n2254 = n2253 ^ x97 ;
  assign n2255 = ~n1898 & n2254 ;
  assign n2256 = n2255 ^ x97 ;
  assign n2251 = n2250 ^ n2249 ;
  assign n2252 = n2251 ^ n2244 ;
  assign n2257 = n2256 ^ n2252 ;
  assign n2258 = n1939 & n2257 ;
  assign n2261 = n2258 ^ n2252 ;
  assign n2262 = n2261 ^ x65 ;
  assign n2263 = ~n1981 & n2262 ;
  assign n2264 = n2263 ^ x65 ;
  assign n2259 = n2258 ^ n2257 ;
  assign n2260 = n2259 ^ n2252 ;
  assign n2265 = n2264 ^ n2260 ;
  assign n2266 = ~n2018 & n2265 ;
  assign n2269 = n2266 ^ n2260 ;
  assign n2270 = n2269 ^ x33 ;
  assign n2271 = ~n2061 & n2270 ;
  assign n2272 = n2271 ^ x33 ;
  assign n2267 = n2266 ^ n2265 ;
  assign n2268 = n2267 ^ n2260 ;
  assign n2273 = n2272 ^ n2268 ;
  assign n2274 = n2101 & n2273 ;
  assign n2277 = n2274 ^ n2268 ;
  assign n2278 = n2277 ^ x1 ;
  assign n2279 = ~n2145 & n2278 ;
  assign n2280 = n2279 ^ x1 ;
  assign n2275 = n2274 ^ n2273 ;
  assign n2276 = n2275 ^ n2268 ;
  assign n2281 = n2280 ^ n2276 ;
  assign n2282 = ~n2180 & n2281 ;
  assign n2283 = n2282 ^ n2281 ;
  assign n2284 = n2283 ^ n2276 ;
  assign n2285 = x226 ^ x194 ;
  assign n2286 = ~n1695 & n2285 ;
  assign n2289 = n2286 ^ x194 ;
  assign n2290 = n2289 ^ x162 ;
  assign n2291 = ~n1738 & n2290 ;
  assign n2292 = n2291 ^ x162 ;
  assign n2287 = n2286 ^ n2285 ;
  assign n2288 = n2287 ^ x194 ;
  assign n2293 = n2292 ^ n2288 ;
  assign n2294 = ~n1775 & n2293 ;
  assign n2297 = n2294 ^ n2288 ;
  assign n2298 = n2297 ^ x130 ;
  assign n2299 = ~n1816 & n2298 ;
  assign n2300 = n2299 ^ x130 ;
  assign n2295 = n2294 ^ n2293 ;
  assign n2296 = n2295 ^ n2288 ;
  assign n2301 = n2300 ^ n2296 ;
  assign n2302 = ~n1855 & n2301 ;
  assign n2305 = n2302 ^ n2296 ;
  assign n2306 = n2305 ^ x98 ;
  assign n2307 = ~n1898 & n2306 ;
  assign n2308 = n2307 ^ x98 ;
  assign n2303 = n2302 ^ n2301 ;
  assign n2304 = n2303 ^ n2296 ;
  assign n2309 = n2308 ^ n2304 ;
  assign n2310 = n1939 & n2309 ;
  assign n2313 = n2310 ^ n2304 ;
  assign n2314 = n2313 ^ x66 ;
  assign n2315 = ~n1981 & n2314 ;
  assign n2316 = n2315 ^ x66 ;
  assign n2311 = n2310 ^ n2309 ;
  assign n2312 = n2311 ^ n2304 ;
  assign n2317 = n2316 ^ n2312 ;
  assign n2318 = ~n2018 & n2317 ;
  assign n2321 = n2318 ^ n2312 ;
  assign n2322 = n2321 ^ x34 ;
  assign n2323 = ~n2061 & n2322 ;
  assign n2324 = n2323 ^ x34 ;
  assign n2319 = n2318 ^ n2317 ;
  assign n2320 = n2319 ^ n2312 ;
  assign n2325 = n2324 ^ n2320 ;
  assign n2326 = n2101 & n2325 ;
  assign n2329 = n2326 ^ n2320 ;
  assign n2330 = n2329 ^ x2 ;
  assign n2331 = ~n2145 & n2330 ;
  assign n2332 = n2331 ^ x2 ;
  assign n2327 = n2326 ^ n2325 ;
  assign n2328 = n2327 ^ n2320 ;
  assign n2333 = n2332 ^ n2328 ;
  assign n2334 = ~n2180 & n2333 ;
  assign n2335 = n2334 ^ n2333 ;
  assign n2336 = n2335 ^ n2328 ;
  assign n2337 = x227 ^ x195 ;
  assign n2338 = ~n1695 & n2337 ;
  assign n2341 = n2338 ^ x195 ;
  assign n2342 = n2341 ^ x163 ;
  assign n2343 = ~n1738 & n2342 ;
  assign n2344 = n2343 ^ x163 ;
  assign n2339 = n2338 ^ n2337 ;
  assign n2340 = n2339 ^ x195 ;
  assign n2345 = n2344 ^ n2340 ;
  assign n2346 = ~n1775 & n2345 ;
  assign n2349 = n2346 ^ n2340 ;
  assign n2350 = n2349 ^ x131 ;
  assign n2351 = ~n1816 & n2350 ;
  assign n2352 = n2351 ^ x131 ;
  assign n2347 = n2346 ^ n2345 ;
  assign n2348 = n2347 ^ n2340 ;
  assign n2353 = n2352 ^ n2348 ;
  assign n2354 = ~n1855 & n2353 ;
  assign n2357 = n2354 ^ n2348 ;
  assign n2358 = n2357 ^ x99 ;
  assign n2359 = ~n1898 & n2358 ;
  assign n2360 = n2359 ^ x99 ;
  assign n2355 = n2354 ^ n2353 ;
  assign n2356 = n2355 ^ n2348 ;
  assign n2361 = n2360 ^ n2356 ;
  assign n2362 = n1939 & n2361 ;
  assign n2365 = n2362 ^ n2356 ;
  assign n2366 = n2365 ^ x67 ;
  assign n2367 = ~n1981 & n2366 ;
  assign n2368 = n2367 ^ x67 ;
  assign n2363 = n2362 ^ n2361 ;
  assign n2364 = n2363 ^ n2356 ;
  assign n2369 = n2368 ^ n2364 ;
  assign n2370 = ~n2018 & n2369 ;
  assign n2373 = n2370 ^ n2364 ;
  assign n2374 = n2373 ^ x35 ;
  assign n2375 = ~n2061 & n2374 ;
  assign n2376 = n2375 ^ x35 ;
  assign n2371 = n2370 ^ n2369 ;
  assign n2372 = n2371 ^ n2364 ;
  assign n2377 = n2376 ^ n2372 ;
  assign n2378 = n2101 & n2377 ;
  assign n2381 = n2378 ^ n2372 ;
  assign n2382 = n2381 ^ x3 ;
  assign n2383 = ~n2145 & n2382 ;
  assign n2384 = n2383 ^ x3 ;
  assign n2379 = n2378 ^ n2377 ;
  assign n2380 = n2379 ^ n2372 ;
  assign n2385 = n2384 ^ n2380 ;
  assign n2386 = ~n2180 & n2385 ;
  assign n2387 = n2386 ^ n2385 ;
  assign n2388 = n2387 ^ n2380 ;
  assign n2389 = x228 ^ x196 ;
  assign n2390 = ~n1695 & n2389 ;
  assign n2393 = n2390 ^ x196 ;
  assign n2394 = n2393 ^ x164 ;
  assign n2395 = ~n1738 & n2394 ;
  assign n2396 = n2395 ^ x164 ;
  assign n2391 = n2390 ^ n2389 ;
  assign n2392 = n2391 ^ x196 ;
  assign n2397 = n2396 ^ n2392 ;
  assign n2398 = ~n1775 & n2397 ;
  assign n2401 = n2398 ^ n2392 ;
  assign n2402 = n2401 ^ x132 ;
  assign n2403 = ~n1816 & n2402 ;
  assign n2404 = n2403 ^ x132 ;
  assign n2399 = n2398 ^ n2397 ;
  assign n2400 = n2399 ^ n2392 ;
  assign n2405 = n2404 ^ n2400 ;
  assign n2406 = ~n1855 & n2405 ;
  assign n2409 = n2406 ^ n2400 ;
  assign n2410 = n2409 ^ x100 ;
  assign n2411 = ~n1898 & n2410 ;
  assign n2412 = n2411 ^ x100 ;
  assign n2407 = n2406 ^ n2405 ;
  assign n2408 = n2407 ^ n2400 ;
  assign n2413 = n2412 ^ n2408 ;
  assign n2414 = n1939 & n2413 ;
  assign n2417 = n2414 ^ n2408 ;
  assign n2418 = n2417 ^ x68 ;
  assign n2419 = ~n1981 & n2418 ;
  assign n2420 = n2419 ^ x68 ;
  assign n2415 = n2414 ^ n2413 ;
  assign n2416 = n2415 ^ n2408 ;
  assign n2421 = n2420 ^ n2416 ;
  assign n2422 = ~n2018 & n2421 ;
  assign n2425 = n2422 ^ n2416 ;
  assign n2426 = n2425 ^ x36 ;
  assign n2427 = ~n2061 & n2426 ;
  assign n2428 = n2427 ^ x36 ;
  assign n2423 = n2422 ^ n2421 ;
  assign n2424 = n2423 ^ n2416 ;
  assign n2429 = n2428 ^ n2424 ;
  assign n2430 = n2101 & n2429 ;
  assign n2433 = n2430 ^ n2424 ;
  assign n2434 = n2433 ^ x4 ;
  assign n2435 = ~n2145 & n2434 ;
  assign n2436 = n2435 ^ x4 ;
  assign n2431 = n2430 ^ n2429 ;
  assign n2432 = n2431 ^ n2424 ;
  assign n2437 = n2436 ^ n2432 ;
  assign n2438 = ~n2180 & n2437 ;
  assign n2439 = n2438 ^ n2437 ;
  assign n2440 = n2439 ^ n2432 ;
  assign n2441 = x229 ^ x197 ;
  assign n2442 = ~n1695 & n2441 ;
  assign n2445 = n2442 ^ x197 ;
  assign n2446 = n2445 ^ x165 ;
  assign n2447 = ~n1738 & n2446 ;
  assign n2448 = n2447 ^ x165 ;
  assign n2443 = n2442 ^ n2441 ;
  assign n2444 = n2443 ^ x197 ;
  assign n2449 = n2448 ^ n2444 ;
  assign n2450 = ~n1775 & n2449 ;
  assign n2453 = n2450 ^ n2444 ;
  assign n2454 = n2453 ^ x133 ;
  assign n2455 = ~n1816 & n2454 ;
  assign n2456 = n2455 ^ x133 ;
  assign n2451 = n2450 ^ n2449 ;
  assign n2452 = n2451 ^ n2444 ;
  assign n2457 = n2456 ^ n2452 ;
  assign n2458 = ~n1855 & n2457 ;
  assign n2461 = n2458 ^ n2452 ;
  assign n2462 = n2461 ^ x101 ;
  assign n2463 = ~n1898 & n2462 ;
  assign n2464 = n2463 ^ x101 ;
  assign n2459 = n2458 ^ n2457 ;
  assign n2460 = n2459 ^ n2452 ;
  assign n2465 = n2464 ^ n2460 ;
  assign n2466 = n1939 & n2465 ;
  assign n2469 = n2466 ^ n2460 ;
  assign n2470 = n2469 ^ x69 ;
  assign n2471 = ~n1981 & n2470 ;
  assign n2472 = n2471 ^ x69 ;
  assign n2467 = n2466 ^ n2465 ;
  assign n2468 = n2467 ^ n2460 ;
  assign n2473 = n2472 ^ n2468 ;
  assign n2474 = ~n2018 & n2473 ;
  assign n2477 = n2474 ^ n2468 ;
  assign n2478 = n2477 ^ x37 ;
  assign n2479 = ~n2061 & n2478 ;
  assign n2480 = n2479 ^ x37 ;
  assign n2475 = n2474 ^ n2473 ;
  assign n2476 = n2475 ^ n2468 ;
  assign n2481 = n2480 ^ n2476 ;
  assign n2482 = n2101 & n2481 ;
  assign n2485 = n2482 ^ n2476 ;
  assign n2486 = n2485 ^ x5 ;
  assign n2487 = ~n2145 & n2486 ;
  assign n2488 = n2487 ^ x5 ;
  assign n2483 = n2482 ^ n2481 ;
  assign n2484 = n2483 ^ n2476 ;
  assign n2489 = n2488 ^ n2484 ;
  assign n2490 = ~n2180 & n2489 ;
  assign n2491 = n2490 ^ n2489 ;
  assign n2492 = n2491 ^ n2484 ;
  assign n2493 = x230 ^ x198 ;
  assign n2494 = ~n1695 & n2493 ;
  assign n2497 = n2494 ^ x198 ;
  assign n2498 = n2497 ^ x166 ;
  assign n2499 = ~n1738 & n2498 ;
  assign n2500 = n2499 ^ x166 ;
  assign n2495 = n2494 ^ n2493 ;
  assign n2496 = n2495 ^ x198 ;
  assign n2501 = n2500 ^ n2496 ;
  assign n2502 = ~n1775 & n2501 ;
  assign n2505 = n2502 ^ n2496 ;
  assign n2506 = n2505 ^ x134 ;
  assign n2507 = ~n1816 & n2506 ;
  assign n2508 = n2507 ^ x134 ;
  assign n2503 = n2502 ^ n2501 ;
  assign n2504 = n2503 ^ n2496 ;
  assign n2509 = n2508 ^ n2504 ;
  assign n2510 = ~n1855 & n2509 ;
  assign n2513 = n2510 ^ n2504 ;
  assign n2514 = n2513 ^ x102 ;
  assign n2515 = ~n1898 & n2514 ;
  assign n2516 = n2515 ^ x102 ;
  assign n2511 = n2510 ^ n2509 ;
  assign n2512 = n2511 ^ n2504 ;
  assign n2517 = n2516 ^ n2512 ;
  assign n2518 = n1939 & n2517 ;
  assign n2521 = n2518 ^ n2512 ;
  assign n2522 = n2521 ^ x70 ;
  assign n2523 = ~n1981 & n2522 ;
  assign n2524 = n2523 ^ x70 ;
  assign n2519 = n2518 ^ n2517 ;
  assign n2520 = n2519 ^ n2512 ;
  assign n2525 = n2524 ^ n2520 ;
  assign n2526 = ~n2018 & n2525 ;
  assign n2529 = n2526 ^ n2520 ;
  assign n2530 = n2529 ^ x38 ;
  assign n2531 = ~n2061 & n2530 ;
  assign n2532 = n2531 ^ x38 ;
  assign n2527 = n2526 ^ n2525 ;
  assign n2528 = n2527 ^ n2520 ;
  assign n2533 = n2532 ^ n2528 ;
  assign n2534 = n2101 & n2533 ;
  assign n2537 = n2534 ^ n2528 ;
  assign n2538 = n2537 ^ x6 ;
  assign n2539 = ~n2145 & n2538 ;
  assign n2540 = n2539 ^ x6 ;
  assign n2535 = n2534 ^ n2533 ;
  assign n2536 = n2535 ^ n2528 ;
  assign n2541 = n2540 ^ n2536 ;
  assign n2542 = ~n2180 & n2541 ;
  assign n2543 = n2542 ^ n2541 ;
  assign n2544 = n2543 ^ n2536 ;
  assign n2545 = x231 ^ x199 ;
  assign n2546 = ~n1695 & n2545 ;
  assign n2549 = n2546 ^ x199 ;
  assign n2550 = n2549 ^ x167 ;
  assign n2551 = ~n1738 & n2550 ;
  assign n2552 = n2551 ^ x167 ;
  assign n2547 = n2546 ^ n2545 ;
  assign n2548 = n2547 ^ x199 ;
  assign n2553 = n2552 ^ n2548 ;
  assign n2554 = ~n1775 & n2553 ;
  assign n2557 = n2554 ^ n2548 ;
  assign n2558 = n2557 ^ x135 ;
  assign n2559 = ~n1816 & n2558 ;
  assign n2560 = n2559 ^ x135 ;
  assign n2555 = n2554 ^ n2553 ;
  assign n2556 = n2555 ^ n2548 ;
  assign n2561 = n2560 ^ n2556 ;
  assign n2562 = ~n1855 & n2561 ;
  assign n2565 = n2562 ^ n2556 ;
  assign n2566 = n2565 ^ x103 ;
  assign n2567 = ~n1898 & n2566 ;
  assign n2568 = n2567 ^ x103 ;
  assign n2563 = n2562 ^ n2561 ;
  assign n2564 = n2563 ^ n2556 ;
  assign n2569 = n2568 ^ n2564 ;
  assign n2570 = n1939 & n2569 ;
  assign n2573 = n2570 ^ n2564 ;
  assign n2574 = n2573 ^ x71 ;
  assign n2575 = ~n1981 & n2574 ;
  assign n2576 = n2575 ^ x71 ;
  assign n2571 = n2570 ^ n2569 ;
  assign n2572 = n2571 ^ n2564 ;
  assign n2577 = n2576 ^ n2572 ;
  assign n2578 = ~n2018 & n2577 ;
  assign n2581 = n2578 ^ n2572 ;
  assign n2582 = n2581 ^ x39 ;
  assign n2583 = ~n2061 & n2582 ;
  assign n2584 = n2583 ^ x39 ;
  assign n2579 = n2578 ^ n2577 ;
  assign n2580 = n2579 ^ n2572 ;
  assign n2585 = n2584 ^ n2580 ;
  assign n2586 = n2101 & n2585 ;
  assign n2589 = n2586 ^ n2580 ;
  assign n2590 = n2589 ^ x7 ;
  assign n2591 = ~n2145 & n2590 ;
  assign n2592 = n2591 ^ x7 ;
  assign n2587 = n2586 ^ n2585 ;
  assign n2588 = n2587 ^ n2580 ;
  assign n2593 = n2592 ^ n2588 ;
  assign n2594 = ~n2180 & n2593 ;
  assign n2595 = n2594 ^ n2593 ;
  assign n2596 = n2595 ^ n2588 ;
  assign n2597 = x232 ^ x200 ;
  assign n2598 = ~n1695 & n2597 ;
  assign n2601 = n2598 ^ x200 ;
  assign n2602 = n2601 ^ x168 ;
  assign n2603 = ~n1738 & n2602 ;
  assign n2604 = n2603 ^ x168 ;
  assign n2599 = n2598 ^ n2597 ;
  assign n2600 = n2599 ^ x200 ;
  assign n2605 = n2604 ^ n2600 ;
  assign n2606 = ~n1775 & n2605 ;
  assign n2609 = n2606 ^ n2600 ;
  assign n2610 = n2609 ^ x136 ;
  assign n2611 = ~n1816 & n2610 ;
  assign n2612 = n2611 ^ x136 ;
  assign n2607 = n2606 ^ n2605 ;
  assign n2608 = n2607 ^ n2600 ;
  assign n2613 = n2612 ^ n2608 ;
  assign n2614 = ~n1855 & n2613 ;
  assign n2617 = n2614 ^ n2608 ;
  assign n2618 = n2617 ^ x104 ;
  assign n2619 = ~n1898 & n2618 ;
  assign n2620 = n2619 ^ x104 ;
  assign n2615 = n2614 ^ n2613 ;
  assign n2616 = n2615 ^ n2608 ;
  assign n2621 = n2620 ^ n2616 ;
  assign n2622 = n1939 & n2621 ;
  assign n2625 = n2622 ^ n2616 ;
  assign n2626 = n2625 ^ x72 ;
  assign n2627 = ~n1981 & n2626 ;
  assign n2628 = n2627 ^ x72 ;
  assign n2623 = n2622 ^ n2621 ;
  assign n2624 = n2623 ^ n2616 ;
  assign n2629 = n2628 ^ n2624 ;
  assign n2630 = ~n2018 & n2629 ;
  assign n2633 = n2630 ^ n2624 ;
  assign n2634 = n2633 ^ x40 ;
  assign n2635 = ~n2061 & n2634 ;
  assign n2636 = n2635 ^ x40 ;
  assign n2631 = n2630 ^ n2629 ;
  assign n2632 = n2631 ^ n2624 ;
  assign n2637 = n2636 ^ n2632 ;
  assign n2638 = n2101 & n2637 ;
  assign n2641 = n2638 ^ n2632 ;
  assign n2642 = n2641 ^ x8 ;
  assign n2643 = ~n2145 & n2642 ;
  assign n2644 = n2643 ^ x8 ;
  assign n2639 = n2638 ^ n2637 ;
  assign n2640 = n2639 ^ n2632 ;
  assign n2645 = n2644 ^ n2640 ;
  assign n2646 = ~n2180 & n2645 ;
  assign n2647 = n2646 ^ n2645 ;
  assign n2648 = n2647 ^ n2640 ;
  assign n2649 = x233 ^ x201 ;
  assign n2650 = ~n1695 & n2649 ;
  assign n2653 = n2650 ^ x201 ;
  assign n2654 = n2653 ^ x169 ;
  assign n2655 = ~n1738 & n2654 ;
  assign n2656 = n2655 ^ x169 ;
  assign n2651 = n2650 ^ n2649 ;
  assign n2652 = n2651 ^ x201 ;
  assign n2657 = n2656 ^ n2652 ;
  assign n2658 = ~n1775 & n2657 ;
  assign n2661 = n2658 ^ n2652 ;
  assign n2662 = n2661 ^ x137 ;
  assign n2663 = ~n1816 & n2662 ;
  assign n2664 = n2663 ^ x137 ;
  assign n2659 = n2658 ^ n2657 ;
  assign n2660 = n2659 ^ n2652 ;
  assign n2665 = n2664 ^ n2660 ;
  assign n2666 = ~n1855 & n2665 ;
  assign n2669 = n2666 ^ n2660 ;
  assign n2670 = n2669 ^ x105 ;
  assign n2671 = ~n1898 & n2670 ;
  assign n2672 = n2671 ^ x105 ;
  assign n2667 = n2666 ^ n2665 ;
  assign n2668 = n2667 ^ n2660 ;
  assign n2673 = n2672 ^ n2668 ;
  assign n2674 = n1939 & n2673 ;
  assign n2677 = n2674 ^ n2668 ;
  assign n2678 = n2677 ^ x73 ;
  assign n2679 = ~n1981 & n2678 ;
  assign n2680 = n2679 ^ x73 ;
  assign n2675 = n2674 ^ n2673 ;
  assign n2676 = n2675 ^ n2668 ;
  assign n2681 = n2680 ^ n2676 ;
  assign n2682 = ~n2018 & n2681 ;
  assign n2685 = n2682 ^ n2676 ;
  assign n2686 = n2685 ^ x41 ;
  assign n2687 = ~n2061 & n2686 ;
  assign n2688 = n2687 ^ x41 ;
  assign n2683 = n2682 ^ n2681 ;
  assign n2684 = n2683 ^ n2676 ;
  assign n2689 = n2688 ^ n2684 ;
  assign n2690 = n2101 & n2689 ;
  assign n2693 = n2690 ^ n2684 ;
  assign n2694 = n2693 ^ x9 ;
  assign n2695 = ~n2145 & n2694 ;
  assign n2696 = n2695 ^ x9 ;
  assign n2691 = n2690 ^ n2689 ;
  assign n2692 = n2691 ^ n2684 ;
  assign n2697 = n2696 ^ n2692 ;
  assign n2698 = ~n2180 & n2697 ;
  assign n2699 = n2698 ^ n2697 ;
  assign n2700 = n2699 ^ n2692 ;
  assign n2701 = x234 ^ x202 ;
  assign n2702 = ~n1695 & n2701 ;
  assign n2705 = n2702 ^ x202 ;
  assign n2706 = n2705 ^ x170 ;
  assign n2707 = ~n1738 & n2706 ;
  assign n2708 = n2707 ^ x170 ;
  assign n2703 = n2702 ^ n2701 ;
  assign n2704 = n2703 ^ x202 ;
  assign n2709 = n2708 ^ n2704 ;
  assign n2710 = ~n1775 & n2709 ;
  assign n2713 = n2710 ^ n2704 ;
  assign n2714 = n2713 ^ x138 ;
  assign n2715 = ~n1816 & n2714 ;
  assign n2716 = n2715 ^ x138 ;
  assign n2711 = n2710 ^ n2709 ;
  assign n2712 = n2711 ^ n2704 ;
  assign n2717 = n2716 ^ n2712 ;
  assign n2718 = ~n1855 & n2717 ;
  assign n2721 = n2718 ^ n2712 ;
  assign n2722 = n2721 ^ x106 ;
  assign n2723 = ~n1898 & n2722 ;
  assign n2724 = n2723 ^ x106 ;
  assign n2719 = n2718 ^ n2717 ;
  assign n2720 = n2719 ^ n2712 ;
  assign n2725 = n2724 ^ n2720 ;
  assign n2726 = n1939 & n2725 ;
  assign n2729 = n2726 ^ n2720 ;
  assign n2730 = n2729 ^ x74 ;
  assign n2731 = ~n1981 & n2730 ;
  assign n2732 = n2731 ^ x74 ;
  assign n2727 = n2726 ^ n2725 ;
  assign n2728 = n2727 ^ n2720 ;
  assign n2733 = n2732 ^ n2728 ;
  assign n2734 = ~n2018 & n2733 ;
  assign n2737 = n2734 ^ n2728 ;
  assign n2738 = n2737 ^ x42 ;
  assign n2739 = ~n2061 & n2738 ;
  assign n2740 = n2739 ^ x42 ;
  assign n2735 = n2734 ^ n2733 ;
  assign n2736 = n2735 ^ n2728 ;
  assign n2741 = n2740 ^ n2736 ;
  assign n2742 = n2101 & n2741 ;
  assign n2745 = n2742 ^ n2736 ;
  assign n2746 = n2745 ^ x10 ;
  assign n2747 = ~n2145 & n2746 ;
  assign n2748 = n2747 ^ x10 ;
  assign n2743 = n2742 ^ n2741 ;
  assign n2744 = n2743 ^ n2736 ;
  assign n2749 = n2748 ^ n2744 ;
  assign n2750 = ~n2180 & n2749 ;
  assign n2751 = n2750 ^ n2749 ;
  assign n2752 = n2751 ^ n2744 ;
  assign n2753 = x235 ^ x203 ;
  assign n2754 = ~n1695 & n2753 ;
  assign n2757 = n2754 ^ x203 ;
  assign n2758 = n2757 ^ x171 ;
  assign n2759 = ~n1738 & n2758 ;
  assign n2760 = n2759 ^ x171 ;
  assign n2755 = n2754 ^ n2753 ;
  assign n2756 = n2755 ^ x203 ;
  assign n2761 = n2760 ^ n2756 ;
  assign n2762 = ~n1775 & n2761 ;
  assign n2765 = n2762 ^ n2756 ;
  assign n2766 = n2765 ^ x139 ;
  assign n2767 = ~n1816 & n2766 ;
  assign n2768 = n2767 ^ x139 ;
  assign n2763 = n2762 ^ n2761 ;
  assign n2764 = n2763 ^ n2756 ;
  assign n2769 = n2768 ^ n2764 ;
  assign n2770 = ~n1855 & n2769 ;
  assign n2773 = n2770 ^ n2764 ;
  assign n2774 = n2773 ^ x107 ;
  assign n2775 = ~n1898 & n2774 ;
  assign n2776 = n2775 ^ x107 ;
  assign n2771 = n2770 ^ n2769 ;
  assign n2772 = n2771 ^ n2764 ;
  assign n2777 = n2776 ^ n2772 ;
  assign n2778 = n1939 & n2777 ;
  assign n2781 = n2778 ^ n2772 ;
  assign n2782 = n2781 ^ x75 ;
  assign n2783 = ~n1981 & n2782 ;
  assign n2784 = n2783 ^ x75 ;
  assign n2779 = n2778 ^ n2777 ;
  assign n2780 = n2779 ^ n2772 ;
  assign n2785 = n2784 ^ n2780 ;
  assign n2786 = ~n2018 & n2785 ;
  assign n2789 = n2786 ^ n2780 ;
  assign n2790 = n2789 ^ x43 ;
  assign n2791 = ~n2061 & n2790 ;
  assign n2792 = n2791 ^ x43 ;
  assign n2787 = n2786 ^ n2785 ;
  assign n2788 = n2787 ^ n2780 ;
  assign n2793 = n2792 ^ n2788 ;
  assign n2794 = n2101 & n2793 ;
  assign n2797 = n2794 ^ n2788 ;
  assign n2798 = n2797 ^ x11 ;
  assign n2799 = ~n2145 & n2798 ;
  assign n2800 = n2799 ^ x11 ;
  assign n2795 = n2794 ^ n2793 ;
  assign n2796 = n2795 ^ n2788 ;
  assign n2801 = n2800 ^ n2796 ;
  assign n2802 = ~n2180 & n2801 ;
  assign n2803 = n2802 ^ n2801 ;
  assign n2804 = n2803 ^ n2796 ;
  assign n2805 = x236 ^ x204 ;
  assign n2806 = ~n1695 & n2805 ;
  assign n2809 = n2806 ^ x204 ;
  assign n2810 = n2809 ^ x172 ;
  assign n2811 = ~n1738 & n2810 ;
  assign n2812 = n2811 ^ x172 ;
  assign n2807 = n2806 ^ n2805 ;
  assign n2808 = n2807 ^ x204 ;
  assign n2813 = n2812 ^ n2808 ;
  assign n2814 = ~n1775 & n2813 ;
  assign n2817 = n2814 ^ n2808 ;
  assign n2818 = n2817 ^ x140 ;
  assign n2819 = ~n1816 & n2818 ;
  assign n2820 = n2819 ^ x140 ;
  assign n2815 = n2814 ^ n2813 ;
  assign n2816 = n2815 ^ n2808 ;
  assign n2821 = n2820 ^ n2816 ;
  assign n2822 = ~n1855 & n2821 ;
  assign n2825 = n2822 ^ n2816 ;
  assign n2826 = n2825 ^ x108 ;
  assign n2827 = ~n1898 & n2826 ;
  assign n2828 = n2827 ^ x108 ;
  assign n2823 = n2822 ^ n2821 ;
  assign n2824 = n2823 ^ n2816 ;
  assign n2829 = n2828 ^ n2824 ;
  assign n2830 = n1939 & n2829 ;
  assign n2833 = n2830 ^ n2824 ;
  assign n2834 = n2833 ^ x76 ;
  assign n2835 = ~n1981 & n2834 ;
  assign n2836 = n2835 ^ x76 ;
  assign n2831 = n2830 ^ n2829 ;
  assign n2832 = n2831 ^ n2824 ;
  assign n2837 = n2836 ^ n2832 ;
  assign n2838 = ~n2018 & n2837 ;
  assign n2841 = n2838 ^ n2832 ;
  assign n2842 = n2841 ^ x44 ;
  assign n2843 = ~n2061 & n2842 ;
  assign n2844 = n2843 ^ x44 ;
  assign n2839 = n2838 ^ n2837 ;
  assign n2840 = n2839 ^ n2832 ;
  assign n2845 = n2844 ^ n2840 ;
  assign n2846 = n2101 & n2845 ;
  assign n2849 = n2846 ^ n2840 ;
  assign n2850 = n2849 ^ x12 ;
  assign n2851 = ~n2145 & n2850 ;
  assign n2852 = n2851 ^ x12 ;
  assign n2847 = n2846 ^ n2845 ;
  assign n2848 = n2847 ^ n2840 ;
  assign n2853 = n2852 ^ n2848 ;
  assign n2854 = ~n2180 & n2853 ;
  assign n2855 = n2854 ^ n2853 ;
  assign n2856 = n2855 ^ n2848 ;
  assign n2857 = x237 ^ x205 ;
  assign n2858 = ~n1695 & n2857 ;
  assign n2861 = n2858 ^ x205 ;
  assign n2862 = n2861 ^ x173 ;
  assign n2863 = ~n1738 & n2862 ;
  assign n2864 = n2863 ^ x173 ;
  assign n2859 = n2858 ^ n2857 ;
  assign n2860 = n2859 ^ x205 ;
  assign n2865 = n2864 ^ n2860 ;
  assign n2866 = ~n1775 & n2865 ;
  assign n2869 = n2866 ^ n2860 ;
  assign n2870 = n2869 ^ x141 ;
  assign n2871 = ~n1816 & n2870 ;
  assign n2872 = n2871 ^ x141 ;
  assign n2867 = n2866 ^ n2865 ;
  assign n2868 = n2867 ^ n2860 ;
  assign n2873 = n2872 ^ n2868 ;
  assign n2874 = ~n1855 & n2873 ;
  assign n2877 = n2874 ^ n2868 ;
  assign n2878 = n2877 ^ x109 ;
  assign n2879 = ~n1898 & n2878 ;
  assign n2880 = n2879 ^ x109 ;
  assign n2875 = n2874 ^ n2873 ;
  assign n2876 = n2875 ^ n2868 ;
  assign n2881 = n2880 ^ n2876 ;
  assign n2882 = n1939 & n2881 ;
  assign n2885 = n2882 ^ n2876 ;
  assign n2886 = n2885 ^ x77 ;
  assign n2887 = ~n1981 & n2886 ;
  assign n2888 = n2887 ^ x77 ;
  assign n2883 = n2882 ^ n2881 ;
  assign n2884 = n2883 ^ n2876 ;
  assign n2889 = n2888 ^ n2884 ;
  assign n2890 = ~n2018 & n2889 ;
  assign n2893 = n2890 ^ n2884 ;
  assign n2894 = n2893 ^ x45 ;
  assign n2895 = ~n2061 & n2894 ;
  assign n2896 = n2895 ^ x45 ;
  assign n2891 = n2890 ^ n2889 ;
  assign n2892 = n2891 ^ n2884 ;
  assign n2897 = n2896 ^ n2892 ;
  assign n2898 = n2101 & n2897 ;
  assign n2901 = n2898 ^ n2892 ;
  assign n2902 = n2901 ^ x13 ;
  assign n2903 = ~n2145 & n2902 ;
  assign n2904 = n2903 ^ x13 ;
  assign n2899 = n2898 ^ n2897 ;
  assign n2900 = n2899 ^ n2892 ;
  assign n2905 = n2904 ^ n2900 ;
  assign n2906 = ~n2180 & n2905 ;
  assign n2907 = n2906 ^ n2905 ;
  assign n2908 = n2907 ^ n2900 ;
  assign n2909 = x238 ^ x206 ;
  assign n2910 = ~n1695 & n2909 ;
  assign n2913 = n2910 ^ x206 ;
  assign n2914 = n2913 ^ x174 ;
  assign n2915 = ~n1738 & n2914 ;
  assign n2916 = n2915 ^ x174 ;
  assign n2911 = n2910 ^ n2909 ;
  assign n2912 = n2911 ^ x206 ;
  assign n2917 = n2916 ^ n2912 ;
  assign n2918 = ~n1775 & n2917 ;
  assign n2921 = n2918 ^ n2912 ;
  assign n2922 = n2921 ^ x142 ;
  assign n2923 = ~n1816 & n2922 ;
  assign n2924 = n2923 ^ x142 ;
  assign n2919 = n2918 ^ n2917 ;
  assign n2920 = n2919 ^ n2912 ;
  assign n2925 = n2924 ^ n2920 ;
  assign n2926 = ~n1855 & n2925 ;
  assign n2929 = n2926 ^ n2920 ;
  assign n2930 = n2929 ^ x110 ;
  assign n2931 = ~n1898 & n2930 ;
  assign n2932 = n2931 ^ x110 ;
  assign n2927 = n2926 ^ n2925 ;
  assign n2928 = n2927 ^ n2920 ;
  assign n2933 = n2932 ^ n2928 ;
  assign n2934 = n1939 & n2933 ;
  assign n2937 = n2934 ^ n2928 ;
  assign n2938 = n2937 ^ x78 ;
  assign n2939 = ~n1981 & n2938 ;
  assign n2940 = n2939 ^ x78 ;
  assign n2935 = n2934 ^ n2933 ;
  assign n2936 = n2935 ^ n2928 ;
  assign n2941 = n2940 ^ n2936 ;
  assign n2942 = ~n2018 & n2941 ;
  assign n2945 = n2942 ^ n2936 ;
  assign n2946 = n2945 ^ x46 ;
  assign n2947 = ~n2061 & n2946 ;
  assign n2948 = n2947 ^ x46 ;
  assign n2943 = n2942 ^ n2941 ;
  assign n2944 = n2943 ^ n2936 ;
  assign n2949 = n2948 ^ n2944 ;
  assign n2950 = n2101 & n2949 ;
  assign n2953 = n2950 ^ n2944 ;
  assign n2954 = n2953 ^ x14 ;
  assign n2955 = ~n2145 & n2954 ;
  assign n2956 = n2955 ^ x14 ;
  assign n2951 = n2950 ^ n2949 ;
  assign n2952 = n2951 ^ n2944 ;
  assign n2957 = n2956 ^ n2952 ;
  assign n2958 = ~n2180 & n2957 ;
  assign n2959 = n2958 ^ n2957 ;
  assign n2960 = n2959 ^ n2952 ;
  assign n2961 = x239 ^ x207 ;
  assign n2962 = ~n1695 & n2961 ;
  assign n2965 = n2962 ^ x207 ;
  assign n2966 = n2965 ^ x175 ;
  assign n2967 = ~n1738 & n2966 ;
  assign n2968 = n2967 ^ x175 ;
  assign n2963 = n2962 ^ n2961 ;
  assign n2964 = n2963 ^ x207 ;
  assign n2969 = n2968 ^ n2964 ;
  assign n2970 = ~n1775 & n2969 ;
  assign n2973 = n2970 ^ n2964 ;
  assign n2974 = n2973 ^ x143 ;
  assign n2975 = ~n1816 & n2974 ;
  assign n2976 = n2975 ^ x143 ;
  assign n2971 = n2970 ^ n2969 ;
  assign n2972 = n2971 ^ n2964 ;
  assign n2977 = n2976 ^ n2972 ;
  assign n2978 = ~n1855 & n2977 ;
  assign n2981 = n2978 ^ n2972 ;
  assign n2982 = n2981 ^ x111 ;
  assign n2983 = ~n1898 & n2982 ;
  assign n2984 = n2983 ^ x111 ;
  assign n2979 = n2978 ^ n2977 ;
  assign n2980 = n2979 ^ n2972 ;
  assign n2985 = n2984 ^ n2980 ;
  assign n2986 = n1939 & n2985 ;
  assign n2989 = n2986 ^ n2980 ;
  assign n2990 = n2989 ^ x79 ;
  assign n2991 = ~n1981 & n2990 ;
  assign n2992 = n2991 ^ x79 ;
  assign n2987 = n2986 ^ n2985 ;
  assign n2988 = n2987 ^ n2980 ;
  assign n2993 = n2992 ^ n2988 ;
  assign n2994 = ~n2018 & n2993 ;
  assign n2997 = n2994 ^ n2988 ;
  assign n2998 = n2997 ^ x47 ;
  assign n2999 = ~n2061 & n2998 ;
  assign n3000 = n2999 ^ x47 ;
  assign n2995 = n2994 ^ n2993 ;
  assign n2996 = n2995 ^ n2988 ;
  assign n3001 = n3000 ^ n2996 ;
  assign n3002 = n2101 & n3001 ;
  assign n3005 = n3002 ^ n2996 ;
  assign n3006 = n3005 ^ x15 ;
  assign n3007 = ~n2145 & n3006 ;
  assign n3008 = n3007 ^ x15 ;
  assign n3003 = n3002 ^ n3001 ;
  assign n3004 = n3003 ^ n2996 ;
  assign n3009 = n3008 ^ n3004 ;
  assign n3010 = ~n2180 & n3009 ;
  assign n3011 = n3010 ^ n3009 ;
  assign n3012 = n3011 ^ n3004 ;
  assign n3013 = x240 ^ x208 ;
  assign n3014 = ~n1695 & n3013 ;
  assign n3017 = n3014 ^ x208 ;
  assign n3018 = n3017 ^ x176 ;
  assign n3019 = ~n1738 & n3018 ;
  assign n3020 = n3019 ^ x176 ;
  assign n3015 = n3014 ^ n3013 ;
  assign n3016 = n3015 ^ x208 ;
  assign n3021 = n3020 ^ n3016 ;
  assign n3022 = ~n1775 & n3021 ;
  assign n3025 = n3022 ^ n3016 ;
  assign n3026 = n3025 ^ x144 ;
  assign n3027 = ~n1816 & n3026 ;
  assign n3028 = n3027 ^ x144 ;
  assign n3023 = n3022 ^ n3021 ;
  assign n3024 = n3023 ^ n3016 ;
  assign n3029 = n3028 ^ n3024 ;
  assign n3030 = ~n1855 & n3029 ;
  assign n3033 = n3030 ^ n3024 ;
  assign n3034 = n3033 ^ x112 ;
  assign n3035 = ~n1898 & n3034 ;
  assign n3036 = n3035 ^ x112 ;
  assign n3031 = n3030 ^ n3029 ;
  assign n3032 = n3031 ^ n3024 ;
  assign n3037 = n3036 ^ n3032 ;
  assign n3038 = n1939 & n3037 ;
  assign n3041 = n3038 ^ n3032 ;
  assign n3042 = n3041 ^ x80 ;
  assign n3043 = ~n1981 & n3042 ;
  assign n3044 = n3043 ^ x80 ;
  assign n3039 = n3038 ^ n3037 ;
  assign n3040 = n3039 ^ n3032 ;
  assign n3045 = n3044 ^ n3040 ;
  assign n3046 = ~n2018 & n3045 ;
  assign n3049 = n3046 ^ n3040 ;
  assign n3050 = n3049 ^ x48 ;
  assign n3051 = ~n2061 & n3050 ;
  assign n3052 = n3051 ^ x48 ;
  assign n3047 = n3046 ^ n3045 ;
  assign n3048 = n3047 ^ n3040 ;
  assign n3053 = n3052 ^ n3048 ;
  assign n3054 = n2101 & n3053 ;
  assign n3057 = n3054 ^ n3048 ;
  assign n3058 = n3057 ^ x16 ;
  assign n3059 = ~n2145 & n3058 ;
  assign n3060 = n3059 ^ x16 ;
  assign n3055 = n3054 ^ n3053 ;
  assign n3056 = n3055 ^ n3048 ;
  assign n3061 = n3060 ^ n3056 ;
  assign n3062 = ~n2180 & n3061 ;
  assign n3063 = n3062 ^ n3061 ;
  assign n3064 = n3063 ^ n3056 ;
  assign n3065 = x241 ^ x209 ;
  assign n3066 = ~n1695 & n3065 ;
  assign n3069 = n3066 ^ x209 ;
  assign n3070 = n3069 ^ x177 ;
  assign n3071 = ~n1738 & n3070 ;
  assign n3072 = n3071 ^ x177 ;
  assign n3067 = n3066 ^ n3065 ;
  assign n3068 = n3067 ^ x209 ;
  assign n3073 = n3072 ^ n3068 ;
  assign n3074 = ~n1775 & n3073 ;
  assign n3077 = n3074 ^ n3068 ;
  assign n3078 = n3077 ^ x145 ;
  assign n3079 = ~n1816 & n3078 ;
  assign n3080 = n3079 ^ x145 ;
  assign n3075 = n3074 ^ n3073 ;
  assign n3076 = n3075 ^ n3068 ;
  assign n3081 = n3080 ^ n3076 ;
  assign n3082 = ~n1855 & n3081 ;
  assign n3085 = n3082 ^ n3076 ;
  assign n3086 = n3085 ^ x113 ;
  assign n3087 = ~n1898 & n3086 ;
  assign n3088 = n3087 ^ x113 ;
  assign n3083 = n3082 ^ n3081 ;
  assign n3084 = n3083 ^ n3076 ;
  assign n3089 = n3088 ^ n3084 ;
  assign n3090 = n1939 & n3089 ;
  assign n3093 = n3090 ^ n3084 ;
  assign n3094 = n3093 ^ x81 ;
  assign n3095 = ~n1981 & n3094 ;
  assign n3096 = n3095 ^ x81 ;
  assign n3091 = n3090 ^ n3089 ;
  assign n3092 = n3091 ^ n3084 ;
  assign n3097 = n3096 ^ n3092 ;
  assign n3098 = ~n2018 & n3097 ;
  assign n3101 = n3098 ^ n3092 ;
  assign n3102 = n3101 ^ x49 ;
  assign n3103 = ~n2061 & n3102 ;
  assign n3104 = n3103 ^ x49 ;
  assign n3099 = n3098 ^ n3097 ;
  assign n3100 = n3099 ^ n3092 ;
  assign n3105 = n3104 ^ n3100 ;
  assign n3106 = n2101 & n3105 ;
  assign n3109 = n3106 ^ n3100 ;
  assign n3110 = n3109 ^ x17 ;
  assign n3111 = ~n2145 & n3110 ;
  assign n3112 = n3111 ^ x17 ;
  assign n3107 = n3106 ^ n3105 ;
  assign n3108 = n3107 ^ n3100 ;
  assign n3113 = n3112 ^ n3108 ;
  assign n3114 = ~n2180 & n3113 ;
  assign n3115 = n3114 ^ n3113 ;
  assign n3116 = n3115 ^ n3108 ;
  assign n3117 = x242 ^ x210 ;
  assign n3118 = ~n1695 & n3117 ;
  assign n3121 = n3118 ^ x210 ;
  assign n3122 = n3121 ^ x178 ;
  assign n3123 = ~n1738 & n3122 ;
  assign n3124 = n3123 ^ x178 ;
  assign n3119 = n3118 ^ n3117 ;
  assign n3120 = n3119 ^ x210 ;
  assign n3125 = n3124 ^ n3120 ;
  assign n3126 = ~n1775 & n3125 ;
  assign n3129 = n3126 ^ n3120 ;
  assign n3130 = n3129 ^ x146 ;
  assign n3131 = ~n1816 & n3130 ;
  assign n3132 = n3131 ^ x146 ;
  assign n3127 = n3126 ^ n3125 ;
  assign n3128 = n3127 ^ n3120 ;
  assign n3133 = n3132 ^ n3128 ;
  assign n3134 = ~n1855 & n3133 ;
  assign n3137 = n3134 ^ n3128 ;
  assign n3138 = n3137 ^ x114 ;
  assign n3139 = ~n1898 & n3138 ;
  assign n3140 = n3139 ^ x114 ;
  assign n3135 = n3134 ^ n3133 ;
  assign n3136 = n3135 ^ n3128 ;
  assign n3141 = n3140 ^ n3136 ;
  assign n3142 = n1939 & n3141 ;
  assign n3145 = n3142 ^ n3136 ;
  assign n3146 = n3145 ^ x82 ;
  assign n3147 = ~n1981 & n3146 ;
  assign n3148 = n3147 ^ x82 ;
  assign n3143 = n3142 ^ n3141 ;
  assign n3144 = n3143 ^ n3136 ;
  assign n3149 = n3148 ^ n3144 ;
  assign n3150 = ~n2018 & n3149 ;
  assign n3153 = n3150 ^ n3144 ;
  assign n3154 = n3153 ^ x50 ;
  assign n3155 = ~n2061 & n3154 ;
  assign n3156 = n3155 ^ x50 ;
  assign n3151 = n3150 ^ n3149 ;
  assign n3152 = n3151 ^ n3144 ;
  assign n3157 = n3156 ^ n3152 ;
  assign n3158 = n2101 & n3157 ;
  assign n3161 = n3158 ^ n3152 ;
  assign n3162 = n3161 ^ x18 ;
  assign n3163 = ~n2145 & n3162 ;
  assign n3164 = n3163 ^ x18 ;
  assign n3159 = n3158 ^ n3157 ;
  assign n3160 = n3159 ^ n3152 ;
  assign n3165 = n3164 ^ n3160 ;
  assign n3166 = ~n2180 & n3165 ;
  assign n3167 = n3166 ^ n3165 ;
  assign n3168 = n3167 ^ n3160 ;
  assign n3169 = x243 ^ x211 ;
  assign n3170 = ~n1695 & n3169 ;
  assign n3173 = n3170 ^ x211 ;
  assign n3174 = n3173 ^ x179 ;
  assign n3175 = ~n1738 & n3174 ;
  assign n3176 = n3175 ^ x179 ;
  assign n3171 = n3170 ^ n3169 ;
  assign n3172 = n3171 ^ x211 ;
  assign n3177 = n3176 ^ n3172 ;
  assign n3178 = ~n1775 & n3177 ;
  assign n3181 = n3178 ^ n3172 ;
  assign n3182 = n3181 ^ x147 ;
  assign n3183 = ~n1816 & n3182 ;
  assign n3184 = n3183 ^ x147 ;
  assign n3179 = n3178 ^ n3177 ;
  assign n3180 = n3179 ^ n3172 ;
  assign n3185 = n3184 ^ n3180 ;
  assign n3186 = ~n1855 & n3185 ;
  assign n3189 = n3186 ^ n3180 ;
  assign n3190 = n3189 ^ x115 ;
  assign n3191 = ~n1898 & n3190 ;
  assign n3192 = n3191 ^ x115 ;
  assign n3187 = n3186 ^ n3185 ;
  assign n3188 = n3187 ^ n3180 ;
  assign n3193 = n3192 ^ n3188 ;
  assign n3194 = n1939 & n3193 ;
  assign n3197 = n3194 ^ n3188 ;
  assign n3198 = n3197 ^ x83 ;
  assign n3199 = ~n1981 & n3198 ;
  assign n3200 = n3199 ^ x83 ;
  assign n3195 = n3194 ^ n3193 ;
  assign n3196 = n3195 ^ n3188 ;
  assign n3201 = n3200 ^ n3196 ;
  assign n3202 = ~n2018 & n3201 ;
  assign n3205 = n3202 ^ n3196 ;
  assign n3206 = n3205 ^ x51 ;
  assign n3207 = ~n2061 & n3206 ;
  assign n3208 = n3207 ^ x51 ;
  assign n3203 = n3202 ^ n3201 ;
  assign n3204 = n3203 ^ n3196 ;
  assign n3209 = n3208 ^ n3204 ;
  assign n3210 = n2101 & n3209 ;
  assign n3213 = n3210 ^ n3204 ;
  assign n3214 = n3213 ^ x19 ;
  assign n3215 = ~n2145 & n3214 ;
  assign n3216 = n3215 ^ x19 ;
  assign n3211 = n3210 ^ n3209 ;
  assign n3212 = n3211 ^ n3204 ;
  assign n3217 = n3216 ^ n3212 ;
  assign n3218 = ~n2180 & n3217 ;
  assign n3219 = n3218 ^ n3217 ;
  assign n3220 = n3219 ^ n3212 ;
  assign n3221 = x244 ^ x212 ;
  assign n3222 = ~n1695 & n3221 ;
  assign n3225 = n3222 ^ x212 ;
  assign n3226 = n3225 ^ x180 ;
  assign n3227 = ~n1738 & n3226 ;
  assign n3228 = n3227 ^ x180 ;
  assign n3223 = n3222 ^ n3221 ;
  assign n3224 = n3223 ^ x212 ;
  assign n3229 = n3228 ^ n3224 ;
  assign n3230 = ~n1775 & n3229 ;
  assign n3233 = n3230 ^ n3224 ;
  assign n3234 = n3233 ^ x148 ;
  assign n3235 = ~n1816 & n3234 ;
  assign n3236 = n3235 ^ x148 ;
  assign n3231 = n3230 ^ n3229 ;
  assign n3232 = n3231 ^ n3224 ;
  assign n3237 = n3236 ^ n3232 ;
  assign n3238 = ~n1855 & n3237 ;
  assign n3241 = n3238 ^ n3232 ;
  assign n3242 = n3241 ^ x116 ;
  assign n3243 = ~n1898 & n3242 ;
  assign n3244 = n3243 ^ x116 ;
  assign n3239 = n3238 ^ n3237 ;
  assign n3240 = n3239 ^ n3232 ;
  assign n3245 = n3244 ^ n3240 ;
  assign n3246 = n1939 & n3245 ;
  assign n3249 = n3246 ^ n3240 ;
  assign n3250 = n3249 ^ x84 ;
  assign n3251 = ~n1981 & n3250 ;
  assign n3252 = n3251 ^ x84 ;
  assign n3247 = n3246 ^ n3245 ;
  assign n3248 = n3247 ^ n3240 ;
  assign n3253 = n3252 ^ n3248 ;
  assign n3254 = ~n2018 & n3253 ;
  assign n3257 = n3254 ^ n3248 ;
  assign n3258 = n3257 ^ x52 ;
  assign n3259 = ~n2061 & n3258 ;
  assign n3260 = n3259 ^ x52 ;
  assign n3255 = n3254 ^ n3253 ;
  assign n3256 = n3255 ^ n3248 ;
  assign n3261 = n3260 ^ n3256 ;
  assign n3262 = n2101 & n3261 ;
  assign n3265 = n3262 ^ n3256 ;
  assign n3266 = n3265 ^ x20 ;
  assign n3267 = ~n2145 & n3266 ;
  assign n3268 = n3267 ^ x20 ;
  assign n3263 = n3262 ^ n3261 ;
  assign n3264 = n3263 ^ n3256 ;
  assign n3269 = n3268 ^ n3264 ;
  assign n3270 = ~n2180 & n3269 ;
  assign n3271 = n3270 ^ n3269 ;
  assign n3272 = n3271 ^ n3264 ;
  assign n3273 = x245 ^ x213 ;
  assign n3274 = ~n1695 & n3273 ;
  assign n3277 = n3274 ^ x213 ;
  assign n3278 = n3277 ^ x181 ;
  assign n3279 = ~n1738 & n3278 ;
  assign n3280 = n3279 ^ x181 ;
  assign n3275 = n3274 ^ n3273 ;
  assign n3276 = n3275 ^ x213 ;
  assign n3281 = n3280 ^ n3276 ;
  assign n3282 = ~n1775 & n3281 ;
  assign n3285 = n3282 ^ n3276 ;
  assign n3286 = n3285 ^ x149 ;
  assign n3287 = ~n1816 & n3286 ;
  assign n3288 = n3287 ^ x149 ;
  assign n3283 = n3282 ^ n3281 ;
  assign n3284 = n3283 ^ n3276 ;
  assign n3289 = n3288 ^ n3284 ;
  assign n3290 = ~n1855 & n3289 ;
  assign n3293 = n3290 ^ n3284 ;
  assign n3294 = n3293 ^ x117 ;
  assign n3295 = ~n1898 & n3294 ;
  assign n3296 = n3295 ^ x117 ;
  assign n3291 = n3290 ^ n3289 ;
  assign n3292 = n3291 ^ n3284 ;
  assign n3297 = n3296 ^ n3292 ;
  assign n3298 = n1939 & n3297 ;
  assign n3301 = n3298 ^ n3292 ;
  assign n3302 = n3301 ^ x85 ;
  assign n3303 = ~n1981 & n3302 ;
  assign n3304 = n3303 ^ x85 ;
  assign n3299 = n3298 ^ n3297 ;
  assign n3300 = n3299 ^ n3292 ;
  assign n3305 = n3304 ^ n3300 ;
  assign n3306 = ~n2018 & n3305 ;
  assign n3309 = n3306 ^ n3300 ;
  assign n3310 = n3309 ^ x53 ;
  assign n3311 = ~n2061 & n3310 ;
  assign n3312 = n3311 ^ x53 ;
  assign n3307 = n3306 ^ n3305 ;
  assign n3308 = n3307 ^ n3300 ;
  assign n3313 = n3312 ^ n3308 ;
  assign n3314 = n2101 & n3313 ;
  assign n3317 = n3314 ^ n3308 ;
  assign n3318 = n3317 ^ x21 ;
  assign n3319 = ~n2145 & n3318 ;
  assign n3320 = n3319 ^ x21 ;
  assign n3315 = n3314 ^ n3313 ;
  assign n3316 = n3315 ^ n3308 ;
  assign n3321 = n3320 ^ n3316 ;
  assign n3322 = ~n2180 & n3321 ;
  assign n3323 = n3322 ^ n3321 ;
  assign n3324 = n3323 ^ n3316 ;
  assign n3325 = x246 ^ x214 ;
  assign n3326 = ~n1695 & n3325 ;
  assign n3329 = n3326 ^ x214 ;
  assign n3330 = n3329 ^ x182 ;
  assign n3331 = ~n1738 & n3330 ;
  assign n3332 = n3331 ^ x182 ;
  assign n3327 = n3326 ^ n3325 ;
  assign n3328 = n3327 ^ x214 ;
  assign n3333 = n3332 ^ n3328 ;
  assign n3334 = ~n1775 & n3333 ;
  assign n3337 = n3334 ^ n3328 ;
  assign n3338 = n3337 ^ x150 ;
  assign n3339 = ~n1816 & n3338 ;
  assign n3340 = n3339 ^ x150 ;
  assign n3335 = n3334 ^ n3333 ;
  assign n3336 = n3335 ^ n3328 ;
  assign n3341 = n3340 ^ n3336 ;
  assign n3342 = ~n1855 & n3341 ;
  assign n3345 = n3342 ^ n3336 ;
  assign n3346 = n3345 ^ x118 ;
  assign n3347 = ~n1898 & n3346 ;
  assign n3348 = n3347 ^ x118 ;
  assign n3343 = n3342 ^ n3341 ;
  assign n3344 = n3343 ^ n3336 ;
  assign n3349 = n3348 ^ n3344 ;
  assign n3350 = n1939 & n3349 ;
  assign n3353 = n3350 ^ n3344 ;
  assign n3354 = n3353 ^ x86 ;
  assign n3355 = ~n1981 & n3354 ;
  assign n3356 = n3355 ^ x86 ;
  assign n3351 = n3350 ^ n3349 ;
  assign n3352 = n3351 ^ n3344 ;
  assign n3357 = n3356 ^ n3352 ;
  assign n3358 = ~n2018 & n3357 ;
  assign n3361 = n3358 ^ n3352 ;
  assign n3362 = n3361 ^ x54 ;
  assign n3363 = ~n2061 & n3362 ;
  assign n3364 = n3363 ^ x54 ;
  assign n3359 = n3358 ^ n3357 ;
  assign n3360 = n3359 ^ n3352 ;
  assign n3365 = n3364 ^ n3360 ;
  assign n3366 = n2101 & n3365 ;
  assign n3369 = n3366 ^ n3360 ;
  assign n3370 = n3369 ^ x22 ;
  assign n3371 = ~n2145 & n3370 ;
  assign n3372 = n3371 ^ x22 ;
  assign n3367 = n3366 ^ n3365 ;
  assign n3368 = n3367 ^ n3360 ;
  assign n3373 = n3372 ^ n3368 ;
  assign n3374 = ~n2180 & n3373 ;
  assign n3375 = n3374 ^ n3373 ;
  assign n3376 = n3375 ^ n3368 ;
  assign n3377 = x247 ^ x215 ;
  assign n3378 = ~n1695 & n3377 ;
  assign n3381 = n3378 ^ x215 ;
  assign n3382 = n3381 ^ x183 ;
  assign n3383 = ~n1738 & n3382 ;
  assign n3384 = n3383 ^ x183 ;
  assign n3379 = n3378 ^ n3377 ;
  assign n3380 = n3379 ^ x215 ;
  assign n3385 = n3384 ^ n3380 ;
  assign n3386 = ~n1775 & n3385 ;
  assign n3389 = n3386 ^ n3380 ;
  assign n3390 = n3389 ^ x151 ;
  assign n3391 = ~n1816 & n3390 ;
  assign n3392 = n3391 ^ x151 ;
  assign n3387 = n3386 ^ n3385 ;
  assign n3388 = n3387 ^ n3380 ;
  assign n3393 = n3392 ^ n3388 ;
  assign n3394 = ~n1855 & n3393 ;
  assign n3397 = n3394 ^ n3388 ;
  assign n3398 = n3397 ^ x119 ;
  assign n3399 = ~n1898 & n3398 ;
  assign n3400 = n3399 ^ x119 ;
  assign n3395 = n3394 ^ n3393 ;
  assign n3396 = n3395 ^ n3388 ;
  assign n3401 = n3400 ^ n3396 ;
  assign n3402 = n1939 & n3401 ;
  assign n3405 = n3402 ^ n3396 ;
  assign n3406 = n3405 ^ x87 ;
  assign n3407 = ~n1981 & n3406 ;
  assign n3408 = n3407 ^ x87 ;
  assign n3403 = n3402 ^ n3401 ;
  assign n3404 = n3403 ^ n3396 ;
  assign n3409 = n3408 ^ n3404 ;
  assign n3410 = ~n2018 & n3409 ;
  assign n3413 = n3410 ^ n3404 ;
  assign n3414 = n3413 ^ x55 ;
  assign n3415 = ~n2061 & n3414 ;
  assign n3416 = n3415 ^ x55 ;
  assign n3411 = n3410 ^ n3409 ;
  assign n3412 = n3411 ^ n3404 ;
  assign n3417 = n3416 ^ n3412 ;
  assign n3418 = n2101 & n3417 ;
  assign n3421 = n3418 ^ n3412 ;
  assign n3422 = n3421 ^ x23 ;
  assign n3423 = ~n2145 & n3422 ;
  assign n3424 = n3423 ^ x23 ;
  assign n3419 = n3418 ^ n3417 ;
  assign n3420 = n3419 ^ n3412 ;
  assign n3425 = n3424 ^ n3420 ;
  assign n3426 = ~n2180 & n3425 ;
  assign n3427 = n3426 ^ n3425 ;
  assign n3428 = n3427 ^ n3420 ;
  assign n3429 = x248 ^ x216 ;
  assign n3430 = ~n1695 & n3429 ;
  assign n3433 = n3430 ^ x216 ;
  assign n3434 = n3433 ^ x184 ;
  assign n3435 = ~n1738 & n3434 ;
  assign n3436 = n3435 ^ x184 ;
  assign n3431 = n3430 ^ n3429 ;
  assign n3432 = n3431 ^ x216 ;
  assign n3437 = n3436 ^ n3432 ;
  assign n3438 = ~n1775 & n3437 ;
  assign n3441 = n3438 ^ n3432 ;
  assign n3442 = n3441 ^ x152 ;
  assign n3443 = ~n1816 & n3442 ;
  assign n3444 = n3443 ^ x152 ;
  assign n3439 = n3438 ^ n3437 ;
  assign n3440 = n3439 ^ n3432 ;
  assign n3445 = n3444 ^ n3440 ;
  assign n3446 = ~n1855 & n3445 ;
  assign n3449 = n3446 ^ n3440 ;
  assign n3450 = n3449 ^ x120 ;
  assign n3451 = ~n1898 & n3450 ;
  assign n3452 = n3451 ^ x120 ;
  assign n3447 = n3446 ^ n3445 ;
  assign n3448 = n3447 ^ n3440 ;
  assign n3453 = n3452 ^ n3448 ;
  assign n3454 = n1939 & n3453 ;
  assign n3457 = n3454 ^ n3448 ;
  assign n3458 = n3457 ^ x88 ;
  assign n3459 = ~n1981 & n3458 ;
  assign n3460 = n3459 ^ x88 ;
  assign n3455 = n3454 ^ n3453 ;
  assign n3456 = n3455 ^ n3448 ;
  assign n3461 = n3460 ^ n3456 ;
  assign n3462 = ~n2018 & n3461 ;
  assign n3465 = n3462 ^ n3456 ;
  assign n3466 = n3465 ^ x56 ;
  assign n3467 = ~n2061 & n3466 ;
  assign n3468 = n3467 ^ x56 ;
  assign n3463 = n3462 ^ n3461 ;
  assign n3464 = n3463 ^ n3456 ;
  assign n3469 = n3468 ^ n3464 ;
  assign n3470 = n2101 & n3469 ;
  assign n3473 = n3470 ^ n3464 ;
  assign n3474 = n3473 ^ x24 ;
  assign n3475 = ~n2145 & n3474 ;
  assign n3476 = n3475 ^ x24 ;
  assign n3471 = n3470 ^ n3469 ;
  assign n3472 = n3471 ^ n3464 ;
  assign n3477 = n3476 ^ n3472 ;
  assign n3478 = ~n2180 & n3477 ;
  assign n3479 = n3478 ^ n3477 ;
  assign n3480 = n3479 ^ n3472 ;
  assign n3481 = x249 ^ x217 ;
  assign n3482 = ~n1695 & n3481 ;
  assign n3485 = n3482 ^ x217 ;
  assign n3486 = n3485 ^ x185 ;
  assign n3487 = ~n1738 & n3486 ;
  assign n3488 = n3487 ^ x185 ;
  assign n3483 = n3482 ^ n3481 ;
  assign n3484 = n3483 ^ x217 ;
  assign n3489 = n3488 ^ n3484 ;
  assign n3490 = ~n1775 & n3489 ;
  assign n3493 = n3490 ^ n3484 ;
  assign n3494 = n3493 ^ x153 ;
  assign n3495 = ~n1816 & n3494 ;
  assign n3496 = n3495 ^ x153 ;
  assign n3491 = n3490 ^ n3489 ;
  assign n3492 = n3491 ^ n3484 ;
  assign n3497 = n3496 ^ n3492 ;
  assign n3498 = ~n1855 & n3497 ;
  assign n3501 = n3498 ^ n3492 ;
  assign n3502 = n3501 ^ x121 ;
  assign n3503 = ~n1898 & n3502 ;
  assign n3504 = n3503 ^ x121 ;
  assign n3499 = n3498 ^ n3497 ;
  assign n3500 = n3499 ^ n3492 ;
  assign n3505 = n3504 ^ n3500 ;
  assign n3506 = n1939 & n3505 ;
  assign n3509 = n3506 ^ n3500 ;
  assign n3510 = n3509 ^ x89 ;
  assign n3511 = ~n1981 & n3510 ;
  assign n3512 = n3511 ^ x89 ;
  assign n3507 = n3506 ^ n3505 ;
  assign n3508 = n3507 ^ n3500 ;
  assign n3513 = n3512 ^ n3508 ;
  assign n3514 = ~n2018 & n3513 ;
  assign n3517 = n3514 ^ n3508 ;
  assign n3518 = n3517 ^ x57 ;
  assign n3519 = ~n2061 & n3518 ;
  assign n3520 = n3519 ^ x57 ;
  assign n3515 = n3514 ^ n3513 ;
  assign n3516 = n3515 ^ n3508 ;
  assign n3521 = n3520 ^ n3516 ;
  assign n3522 = n2101 & n3521 ;
  assign n3525 = n3522 ^ n3516 ;
  assign n3526 = n3525 ^ x25 ;
  assign n3527 = ~n2145 & n3526 ;
  assign n3528 = n3527 ^ x25 ;
  assign n3523 = n3522 ^ n3521 ;
  assign n3524 = n3523 ^ n3516 ;
  assign n3529 = n3528 ^ n3524 ;
  assign n3530 = ~n2180 & n3529 ;
  assign n3531 = n3530 ^ n3529 ;
  assign n3532 = n3531 ^ n3524 ;
  assign n3533 = x250 ^ x218 ;
  assign n3534 = ~n1695 & n3533 ;
  assign n3537 = n3534 ^ x218 ;
  assign n3538 = n3537 ^ x186 ;
  assign n3539 = ~n1738 & n3538 ;
  assign n3540 = n3539 ^ x186 ;
  assign n3535 = n3534 ^ n3533 ;
  assign n3536 = n3535 ^ x218 ;
  assign n3541 = n3540 ^ n3536 ;
  assign n3542 = ~n1775 & n3541 ;
  assign n3545 = n3542 ^ n3536 ;
  assign n3546 = n3545 ^ x154 ;
  assign n3547 = ~n1816 & n3546 ;
  assign n3548 = n3547 ^ x154 ;
  assign n3543 = n3542 ^ n3541 ;
  assign n3544 = n3543 ^ n3536 ;
  assign n3549 = n3548 ^ n3544 ;
  assign n3550 = ~n1855 & n3549 ;
  assign n3553 = n3550 ^ n3544 ;
  assign n3554 = n3553 ^ x122 ;
  assign n3555 = ~n1898 & n3554 ;
  assign n3556 = n3555 ^ x122 ;
  assign n3551 = n3550 ^ n3549 ;
  assign n3552 = n3551 ^ n3544 ;
  assign n3557 = n3556 ^ n3552 ;
  assign n3558 = n1939 & n3557 ;
  assign n3561 = n3558 ^ n3552 ;
  assign n3562 = n3561 ^ x90 ;
  assign n3563 = ~n1981 & n3562 ;
  assign n3564 = n3563 ^ x90 ;
  assign n3559 = n3558 ^ n3557 ;
  assign n3560 = n3559 ^ n3552 ;
  assign n3565 = n3564 ^ n3560 ;
  assign n3566 = ~n2018 & n3565 ;
  assign n3569 = n3566 ^ n3560 ;
  assign n3570 = n3569 ^ x58 ;
  assign n3571 = ~n2061 & n3570 ;
  assign n3572 = n3571 ^ x58 ;
  assign n3567 = n3566 ^ n3565 ;
  assign n3568 = n3567 ^ n3560 ;
  assign n3573 = n3572 ^ n3568 ;
  assign n3574 = n2101 & n3573 ;
  assign n3577 = n3574 ^ n3568 ;
  assign n3578 = n3577 ^ x26 ;
  assign n3579 = ~n2145 & n3578 ;
  assign n3580 = n3579 ^ x26 ;
  assign n3575 = n3574 ^ n3573 ;
  assign n3576 = n3575 ^ n3568 ;
  assign n3581 = n3580 ^ n3576 ;
  assign n3582 = ~n2180 & n3581 ;
  assign n3583 = n3582 ^ n3581 ;
  assign n3584 = n3583 ^ n3576 ;
  assign n3585 = x251 ^ x219 ;
  assign n3586 = ~n1695 & n3585 ;
  assign n3589 = n3586 ^ x219 ;
  assign n3590 = n3589 ^ x187 ;
  assign n3591 = ~n1738 & n3590 ;
  assign n3592 = n3591 ^ x187 ;
  assign n3587 = n3586 ^ n3585 ;
  assign n3588 = n3587 ^ x219 ;
  assign n3593 = n3592 ^ n3588 ;
  assign n3594 = ~n1775 & n3593 ;
  assign n3597 = n3594 ^ n3588 ;
  assign n3598 = n3597 ^ x155 ;
  assign n3599 = ~n1816 & n3598 ;
  assign n3600 = n3599 ^ x155 ;
  assign n3595 = n3594 ^ n3593 ;
  assign n3596 = n3595 ^ n3588 ;
  assign n3601 = n3600 ^ n3596 ;
  assign n3602 = ~n1855 & n3601 ;
  assign n3605 = n3602 ^ n3596 ;
  assign n3606 = n3605 ^ x123 ;
  assign n3607 = ~n1898 & n3606 ;
  assign n3608 = n3607 ^ x123 ;
  assign n3603 = n3602 ^ n3601 ;
  assign n3604 = n3603 ^ n3596 ;
  assign n3609 = n3608 ^ n3604 ;
  assign n3610 = n1939 & n3609 ;
  assign n3613 = n3610 ^ n3604 ;
  assign n3614 = n3613 ^ x91 ;
  assign n3615 = ~n1981 & n3614 ;
  assign n3616 = n3615 ^ x91 ;
  assign n3611 = n3610 ^ n3609 ;
  assign n3612 = n3611 ^ n3604 ;
  assign n3617 = n3616 ^ n3612 ;
  assign n3618 = ~n2018 & n3617 ;
  assign n3621 = n3618 ^ n3612 ;
  assign n3622 = n3621 ^ x59 ;
  assign n3623 = ~n2061 & n3622 ;
  assign n3624 = n3623 ^ x59 ;
  assign n3619 = n3618 ^ n3617 ;
  assign n3620 = n3619 ^ n3612 ;
  assign n3625 = n3624 ^ n3620 ;
  assign n3626 = n2101 & n3625 ;
  assign n3629 = n3626 ^ n3620 ;
  assign n3630 = n3629 ^ x27 ;
  assign n3631 = ~n2145 & n3630 ;
  assign n3632 = n3631 ^ x27 ;
  assign n3627 = n3626 ^ n3625 ;
  assign n3628 = n3627 ^ n3620 ;
  assign n3633 = n3632 ^ n3628 ;
  assign n3634 = ~n2180 & n3633 ;
  assign n3635 = n3634 ^ n3633 ;
  assign n3636 = n3635 ^ n3628 ;
  assign n3637 = x252 ^ x220 ;
  assign n3638 = ~n1695 & n3637 ;
  assign n3641 = n3638 ^ x220 ;
  assign n3642 = n3641 ^ x188 ;
  assign n3643 = ~n1738 & n3642 ;
  assign n3644 = n3643 ^ x188 ;
  assign n3639 = n3638 ^ n3637 ;
  assign n3640 = n3639 ^ x220 ;
  assign n3645 = n3644 ^ n3640 ;
  assign n3646 = ~n1775 & n3645 ;
  assign n3649 = n3646 ^ n3640 ;
  assign n3650 = n3649 ^ x156 ;
  assign n3651 = ~n1816 & n3650 ;
  assign n3652 = n3651 ^ x156 ;
  assign n3647 = n3646 ^ n3645 ;
  assign n3648 = n3647 ^ n3640 ;
  assign n3653 = n3652 ^ n3648 ;
  assign n3654 = ~n1855 & n3653 ;
  assign n3657 = n3654 ^ n3648 ;
  assign n3658 = n3657 ^ x124 ;
  assign n3659 = ~n1898 & n3658 ;
  assign n3660 = n3659 ^ x124 ;
  assign n3655 = n3654 ^ n3653 ;
  assign n3656 = n3655 ^ n3648 ;
  assign n3661 = n3660 ^ n3656 ;
  assign n3662 = n1939 & n3661 ;
  assign n3665 = n3662 ^ n3656 ;
  assign n3666 = n3665 ^ x92 ;
  assign n3667 = ~n1981 & n3666 ;
  assign n3668 = n3667 ^ x92 ;
  assign n3663 = n3662 ^ n3661 ;
  assign n3664 = n3663 ^ n3656 ;
  assign n3669 = n3668 ^ n3664 ;
  assign n3670 = ~n2018 & n3669 ;
  assign n3673 = n3670 ^ n3664 ;
  assign n3674 = n3673 ^ x60 ;
  assign n3675 = ~n2061 & n3674 ;
  assign n3676 = n3675 ^ x60 ;
  assign n3671 = n3670 ^ n3669 ;
  assign n3672 = n3671 ^ n3664 ;
  assign n3677 = n3676 ^ n3672 ;
  assign n3678 = n2101 & n3677 ;
  assign n3681 = n3678 ^ n3672 ;
  assign n3682 = n3681 ^ x28 ;
  assign n3683 = ~n2145 & n3682 ;
  assign n3684 = n3683 ^ x28 ;
  assign n3679 = n3678 ^ n3677 ;
  assign n3680 = n3679 ^ n3672 ;
  assign n3685 = n3684 ^ n3680 ;
  assign n3686 = ~n2180 & n3685 ;
  assign n3687 = n3686 ^ n3685 ;
  assign n3688 = n3687 ^ n3680 ;
  assign n3689 = x253 ^ x221 ;
  assign n3690 = ~n1695 & n3689 ;
  assign n3693 = n3690 ^ x221 ;
  assign n3694 = n3693 ^ x189 ;
  assign n3695 = ~n1738 & n3694 ;
  assign n3696 = n3695 ^ x189 ;
  assign n3691 = n3690 ^ n3689 ;
  assign n3692 = n3691 ^ x221 ;
  assign n3697 = n3696 ^ n3692 ;
  assign n3698 = ~n1775 & n3697 ;
  assign n3701 = n3698 ^ n3692 ;
  assign n3702 = n3701 ^ x157 ;
  assign n3703 = ~n1816 & n3702 ;
  assign n3704 = n3703 ^ x157 ;
  assign n3699 = n3698 ^ n3697 ;
  assign n3700 = n3699 ^ n3692 ;
  assign n3705 = n3704 ^ n3700 ;
  assign n3706 = ~n1855 & n3705 ;
  assign n3709 = n3706 ^ n3700 ;
  assign n3710 = n3709 ^ x125 ;
  assign n3711 = ~n1898 & n3710 ;
  assign n3712 = n3711 ^ x125 ;
  assign n3707 = n3706 ^ n3705 ;
  assign n3708 = n3707 ^ n3700 ;
  assign n3713 = n3712 ^ n3708 ;
  assign n3714 = n1939 & n3713 ;
  assign n3717 = n3714 ^ n3708 ;
  assign n3718 = n3717 ^ x93 ;
  assign n3719 = ~n1981 & n3718 ;
  assign n3720 = n3719 ^ x93 ;
  assign n3715 = n3714 ^ n3713 ;
  assign n3716 = n3715 ^ n3708 ;
  assign n3721 = n3720 ^ n3716 ;
  assign n3722 = ~n2018 & n3721 ;
  assign n3725 = n3722 ^ n3716 ;
  assign n3726 = n3725 ^ x61 ;
  assign n3727 = ~n2061 & n3726 ;
  assign n3728 = n3727 ^ x61 ;
  assign n3723 = n3722 ^ n3721 ;
  assign n3724 = n3723 ^ n3716 ;
  assign n3729 = n3728 ^ n3724 ;
  assign n3730 = n2101 & n3729 ;
  assign n3733 = n3730 ^ n3724 ;
  assign n3734 = n3733 ^ x29 ;
  assign n3735 = ~n2145 & n3734 ;
  assign n3736 = n3735 ^ x29 ;
  assign n3731 = n3730 ^ n3729 ;
  assign n3732 = n3731 ^ n3724 ;
  assign n3737 = n3736 ^ n3732 ;
  assign n3738 = ~n2180 & n3737 ;
  assign n3739 = n3738 ^ n3737 ;
  assign n3740 = n3739 ^ n3732 ;
  assign n3741 = x254 ^ x222 ;
  assign n3742 = ~n1695 & n3741 ;
  assign n3745 = n3742 ^ x222 ;
  assign n3746 = n3745 ^ x190 ;
  assign n3747 = ~n1738 & n3746 ;
  assign n3748 = n3747 ^ x190 ;
  assign n3743 = n3742 ^ n3741 ;
  assign n3744 = n3743 ^ x222 ;
  assign n3749 = n3748 ^ n3744 ;
  assign n3750 = ~n1775 & n3749 ;
  assign n3753 = n3750 ^ n3744 ;
  assign n3754 = n3753 ^ x158 ;
  assign n3755 = ~n1816 & n3754 ;
  assign n3756 = n3755 ^ x158 ;
  assign n3751 = n3750 ^ n3749 ;
  assign n3752 = n3751 ^ n3744 ;
  assign n3757 = n3756 ^ n3752 ;
  assign n3758 = ~n1855 & n3757 ;
  assign n3761 = n3758 ^ n3752 ;
  assign n3762 = n3761 ^ x126 ;
  assign n3763 = ~n1898 & n3762 ;
  assign n3764 = n3763 ^ x126 ;
  assign n3759 = n3758 ^ n3757 ;
  assign n3760 = n3759 ^ n3752 ;
  assign n3765 = n3764 ^ n3760 ;
  assign n3766 = n1939 & n3765 ;
  assign n3769 = n3766 ^ n3760 ;
  assign n3770 = n3769 ^ x94 ;
  assign n3771 = ~n1981 & n3770 ;
  assign n3772 = n3771 ^ x94 ;
  assign n3767 = n3766 ^ n3765 ;
  assign n3768 = n3767 ^ n3760 ;
  assign n3773 = n3772 ^ n3768 ;
  assign n3774 = ~n2018 & n3773 ;
  assign n3777 = n3774 ^ n3768 ;
  assign n3778 = n3777 ^ x62 ;
  assign n3779 = ~n2061 & n3778 ;
  assign n3780 = n3779 ^ x62 ;
  assign n3775 = n3774 ^ n3773 ;
  assign n3776 = n3775 ^ n3768 ;
  assign n3781 = n3780 ^ n3776 ;
  assign n3782 = n2101 & n3781 ;
  assign n3785 = n3782 ^ n3776 ;
  assign n3786 = n3785 ^ x30 ;
  assign n3787 = ~n2145 & n3786 ;
  assign n3788 = n3787 ^ x30 ;
  assign n3783 = n3782 ^ n3781 ;
  assign n3784 = n3783 ^ n3776 ;
  assign n3789 = n3788 ^ n3784 ;
  assign n3790 = ~n2180 & n3789 ;
  assign n3791 = n3790 ^ n3789 ;
  assign n3792 = n3791 ^ n3784 ;
  assign n3793 = x255 ^ x223 ;
  assign n3794 = ~n1695 & n3793 ;
  assign n3797 = n3794 ^ x223 ;
  assign n3798 = n3797 ^ x191 ;
  assign n3799 = ~n1738 & n3798 ;
  assign n3800 = n3799 ^ x191 ;
  assign n3795 = n3794 ^ n3793 ;
  assign n3796 = n3795 ^ x223 ;
  assign n3801 = n3800 ^ n3796 ;
  assign n3802 = ~n1775 & n3801 ;
  assign n3805 = n3802 ^ n3796 ;
  assign n3806 = n3805 ^ x159 ;
  assign n3807 = ~n1816 & n3806 ;
  assign n3808 = n3807 ^ x159 ;
  assign n3803 = n3802 ^ n3801 ;
  assign n3804 = n3803 ^ n3796 ;
  assign n3809 = n3808 ^ n3804 ;
  assign n3810 = ~n1855 & n3809 ;
  assign n3813 = n3810 ^ n3804 ;
  assign n3814 = n3813 ^ x127 ;
  assign n3815 = ~n1898 & n3814 ;
  assign n3816 = n3815 ^ x127 ;
  assign n3811 = n3810 ^ n3809 ;
  assign n3812 = n3811 ^ n3804 ;
  assign n3817 = n3816 ^ n3812 ;
  assign n3818 = n1939 & n3817 ;
  assign n3821 = n3818 ^ n3812 ;
  assign n3822 = n3821 ^ x95 ;
  assign n3823 = ~n1981 & n3822 ;
  assign n3824 = n3823 ^ x95 ;
  assign n3819 = n3818 ^ n3817 ;
  assign n3820 = n3819 ^ n3812 ;
  assign n3825 = n3824 ^ n3820 ;
  assign n3826 = ~n2018 & n3825 ;
  assign n3829 = n3826 ^ n3820 ;
  assign n3830 = n3829 ^ x63 ;
  assign n3831 = ~n2061 & n3830 ;
  assign n3832 = n3831 ^ x63 ;
  assign n3827 = n3826 ^ n3825 ;
  assign n3828 = n3827 ^ n3820 ;
  assign n3833 = n3832 ^ n3828 ;
  assign n3834 = n2101 & n3833 ;
  assign n3837 = n3834 ^ n3828 ;
  assign n3838 = n3837 ^ x31 ;
  assign n3839 = ~n2145 & n3838 ;
  assign n3840 = n3839 ^ x31 ;
  assign n3835 = n3834 ^ n3833 ;
  assign n3836 = n3835 ^ n3828 ;
  assign n3841 = n3840 ^ n3836 ;
  assign n3842 = ~n2180 & n3841 ;
  assign n3843 = n3842 ^ n3841 ;
  assign n3844 = n3843 ^ n3836 ;
  assign n3845 = n2230 ^ n2224 ;
  assign n3846 = n2282 ^ n2276 ;
  assign n3847 = n2334 ^ n2328 ;
  assign n3848 = n2386 ^ n2380 ;
  assign n3849 = n2438 ^ n2432 ;
  assign n3850 = n2490 ^ n2484 ;
  assign n3851 = n2542 ^ n2536 ;
  assign n3852 = n2594 ^ n2588 ;
  assign n3853 = n2646 ^ n2640 ;
  assign n3854 = n2698 ^ n2692 ;
  assign n3855 = n2750 ^ n2744 ;
  assign n3856 = n2802 ^ n2796 ;
  assign n3857 = n2854 ^ n2848 ;
  assign n3858 = n2906 ^ n2900 ;
  assign n3859 = n2958 ^ n2952 ;
  assign n3860 = n3010 ^ n3004 ;
  assign n3861 = n3062 ^ n3056 ;
  assign n3862 = n3114 ^ n3108 ;
  assign n3863 = n3166 ^ n3160 ;
  assign n3864 = n3218 ^ n3212 ;
  assign n3865 = n3270 ^ n3264 ;
  assign n3866 = n3322 ^ n3316 ;
  assign n3867 = n3374 ^ n3368 ;
  assign n3868 = n3426 ^ n3420 ;
  assign n3869 = n3478 ^ n3472 ;
  assign n3870 = n3530 ^ n3524 ;
  assign n3871 = n3582 ^ n3576 ;
  assign n3872 = n3634 ^ n3628 ;
  assign n3873 = n3686 ^ n3680 ;
  assign n3874 = n3738 ^ n3732 ;
  assign n3875 = n3790 ^ n3784 ;
  assign n3876 = n3842 ^ n3836 ;
  assign y0 = n2232 ;
  assign y1 = n2284 ;
  assign y2 = n2336 ;
  assign y3 = n2388 ;
  assign y4 = n2440 ;
  assign y5 = n2492 ;
  assign y6 = n2544 ;
  assign y7 = n2596 ;
  assign y8 = n2648 ;
  assign y9 = n2700 ;
  assign y10 = n2752 ;
  assign y11 = n2804 ;
  assign y12 = n2856 ;
  assign y13 = n2908 ;
  assign y14 = n2960 ;
  assign y15 = n3012 ;
  assign y16 = n3064 ;
  assign y17 = n3116 ;
  assign y18 = n3168 ;
  assign y19 = n3220 ;
  assign y20 = n3272 ;
  assign y21 = n3324 ;
  assign y22 = n3376 ;
  assign y23 = n3428 ;
  assign y24 = n3480 ;
  assign y25 = n3532 ;
  assign y26 = n3584 ;
  assign y27 = n3636 ;
  assign y28 = n3688 ;
  assign y29 = n3740 ;
  assign y30 = n3792 ;
  assign y31 = n3844 ;
  assign y32 = n3845 ;
  assign y33 = n3846 ;
  assign y34 = n3847 ;
  assign y35 = n3848 ;
  assign y36 = n3849 ;
  assign y37 = n3850 ;
  assign y38 = n3851 ;
  assign y39 = n3852 ;
  assign y40 = n3853 ;
  assign y41 = n3854 ;
  assign y42 = n3855 ;
  assign y43 = n3856 ;
  assign y44 = n3857 ;
  assign y45 = n3858 ;
  assign y46 = n3859 ;
  assign y47 = n3860 ;
  assign y48 = n3861 ;
  assign y49 = n3862 ;
  assign y50 = n3863 ;
  assign y51 = n3864 ;
  assign y52 = n3865 ;
  assign y53 = n3866 ;
  assign y54 = n3867 ;
  assign y55 = n3868 ;
  assign y56 = n3869 ;
  assign y57 = n3870 ;
  assign y58 = n3871 ;
  assign y59 = n3872 ;
  assign y60 = n3873 ;
  assign y61 = n3874 ;
  assign y62 = n3875 ;
  assign y63 = n3876 ;
endmodule
