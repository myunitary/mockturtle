module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 ;
  assign n33 = x31 ^ x0 ;
  assign n34 = n33 ^ x31 ;
  assign n36 = ~x0 & x31 ;
  assign n35 = x31 ^ x1 ;
  assign n37 = n36 ^ n35 ;
  assign n39 = n35 & n36 ;
  assign n38 = x31 ^ x2 ;
  assign n40 = n39 ^ n38 ;
  assign n42 = n38 & n39 ;
  assign n41 = x31 ^ x3 ;
  assign n43 = n42 ^ n41 ;
  assign n45 = n38 & n41 ;
  assign n46 = n39 & n45 ;
  assign n44 = x31 ^ x4 ;
  assign n47 = n46 ^ n44 ;
  assign n49 = n44 & n46 ;
  assign n48 = x31 ^ x5 ;
  assign n50 = n49 ^ n48 ;
  assign n52 = n44 & n48 ;
  assign n53 = n46 & n52 ;
  assign n51 = x31 ^ x6 ;
  assign n54 = n53 ^ n51 ;
  assign n56 = n51 & n52 ;
  assign n57 = n46 & n56 ;
  assign n55 = x31 ^ x7 ;
  assign n58 = n57 ^ n55 ;
  assign n60 = n51 & n55 ;
  assign n61 = n52 & n60 ;
  assign n62 = n46 & n61 ;
  assign n59 = x31 ^ x8 ;
  assign n63 = n62 ^ n59 ;
  assign n65 = n59 & n62 ;
  assign n64 = x31 ^ x9 ;
  assign n66 = n65 ^ n64 ;
  assign n68 = n59 & n64 ;
  assign n69 = n62 & n68 ;
  assign n67 = x31 ^ x10 ;
  assign n70 = n69 ^ n67 ;
  assign n72 = n67 & n68 ;
  assign n73 = n62 & n72 ;
  assign n71 = x31 ^ x11 ;
  assign n74 = n73 ^ n71 ;
  assign n76 = n67 & n71 ;
  assign n77 = n68 & n76 ;
  assign n78 = n62 & n77 ;
  assign n75 = x31 ^ x12 ;
  assign n79 = n78 ^ n75 ;
  assign n81 = n75 & n77 ;
  assign n82 = n62 & n81 ;
  assign n80 = x31 ^ x13 ;
  assign n83 = n82 ^ n80 ;
  assign n85 = n75 & n80 ;
  assign n86 = n77 & n85 ;
  assign n87 = n62 & n86 ;
  assign n84 = x31 ^ x14 ;
  assign n88 = n87 ^ n84 ;
  assign n90 = n84 & n85 ;
  assign n91 = n77 & n90 ;
  assign n92 = n62 & n91 ;
  assign n89 = x31 ^ x15 ;
  assign n93 = n92 ^ n89 ;
  assign n95 = n84 & n89 ;
  assign n96 = n85 & n95 ;
  assign n97 = n77 & n96 ;
  assign n98 = n62 & n97 ;
  assign n94 = x31 ^ x16 ;
  assign n99 = n98 ^ n94 ;
  assign n101 = n94 & n98 ;
  assign n100 = x31 ^ x17 ;
  assign n102 = n101 ^ n100 ;
  assign n104 = n94 & n100 ;
  assign n105 = n98 & n104 ;
  assign n103 = x31 ^ x18 ;
  assign n106 = n105 ^ n103 ;
  assign n108 = n103 & n104 ;
  assign n109 = n98 & n108 ;
  assign n107 = x31 ^ x19 ;
  assign n110 = n109 ^ n107 ;
  assign n112 = n103 & n107 ;
  assign n113 = n104 & n112 ;
  assign n114 = n98 & n113 ;
  assign n111 = x31 ^ x20 ;
  assign n115 = n114 ^ n111 ;
  assign n117 = n111 & n113 ;
  assign n118 = n98 & n117 ;
  assign n116 = x31 ^ x21 ;
  assign n119 = n118 ^ n116 ;
  assign n121 = n111 & n116 ;
  assign n122 = n113 & n121 ;
  assign n123 = n98 & n122 ;
  assign n120 = x31 ^ x22 ;
  assign n124 = n123 ^ n120 ;
  assign n126 = n120 & n121 ;
  assign n127 = n113 & n126 ;
  assign n128 = n98 & n127 ;
  assign n125 = x31 ^ x23 ;
  assign n129 = n128 ^ n125 ;
  assign n131 = n120 & n125 ;
  assign n132 = n121 & n131 ;
  assign n133 = n113 & n132 ;
  assign n134 = n98 & n133 ;
  assign n130 = x31 ^ x24 ;
  assign n135 = n134 ^ n130 ;
  assign n137 = n130 & n133 ;
  assign n138 = n98 & n137 ;
  assign n136 = x31 ^ x25 ;
  assign n139 = n138 ^ n136 ;
  assign n141 = n130 & n136 ;
  assign n142 = n133 & n141 ;
  assign n143 = n98 & n142 ;
  assign n140 = x31 ^ x26 ;
  assign n144 = n143 ^ n140 ;
  assign n146 = n140 & n141 ;
  assign n147 = n133 & n146 ;
  assign n148 = n98 & n147 ;
  assign n145 = x31 ^ x27 ;
  assign n149 = n148 ^ n145 ;
  assign n151 = n140 & n145 ;
  assign n152 = n141 & n151 ;
  assign n153 = n133 & n152 ;
  assign n154 = n98 & n153 ;
  assign n150 = x31 ^ x28 ;
  assign n155 = n154 ^ n150 ;
  assign n157 = n150 & n152 ;
  assign n158 = n133 & n157 ;
  assign n159 = n98 & n158 ;
  assign n156 = x31 ^ x29 ;
  assign n160 = n159 ^ n156 ;
  assign n162 = n150 & n156 ;
  assign n163 = n152 & n162 ;
  assign n164 = n133 & n163 ;
  assign n165 = n98 & n164 ;
  assign n161 = x31 ^ x30 ;
  assign n166 = n165 ^ n161 ;
  assign n167 = n161 & n162 ;
  assign n168 = n152 & n167 ;
  assign n169 = n133 & n168 ;
  assign n170 = n98 & n169 ;
  assign y0 = n34 ;
  assign y1 = n37 ;
  assign y2 = n40 ;
  assign y3 = n43 ;
  assign y4 = n47 ;
  assign y5 = n50 ;
  assign y6 = n54 ;
  assign y7 = n58 ;
  assign y8 = n63 ;
  assign y9 = n66 ;
  assign y10 = n70 ;
  assign y11 = n74 ;
  assign y12 = n79 ;
  assign y13 = n83 ;
  assign y14 = n88 ;
  assign y15 = n93 ;
  assign y16 = n99 ;
  assign y17 = n102 ;
  assign y18 = n106 ;
  assign y19 = n110 ;
  assign y20 = n115 ;
  assign y21 = n119 ;
  assign y22 = n124 ;
  assign y23 = n129 ;
  assign y24 = n135 ;
  assign y25 = n139 ;
  assign y26 = n144 ;
  assign y27 = n149 ;
  assign y28 = n155 ;
  assign y29 = n160 ;
  assign y30 = n166 ;
  assign y31 = n170 ;
endmodule
