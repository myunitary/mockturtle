module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 ;
  assign n190 = x33 ^ x1 ;
  assign n191 = x0 & ~x32 ;
  assign n192 = ~n190 & n191 ;
  assign n189 = x1 & ~x33 ;
  assign n193 = n192 ^ n189 ;
  assign n185 = x35 ^ x3 ;
  assign n194 = x34 ^ x2 ;
  assign n195 = ~n185 & ~n194 ;
  assign n196 = n193 & n195 ;
  assign n186 = x2 & ~x34 ;
  assign n187 = ~n185 & n186 ;
  assign n184 = x3 & ~x35 ;
  assign n188 = n187 ^ n184 ;
  assign n197 = n196 ^ n188 ;
  assign n171 = x39 ^ x7 ;
  assign n175 = x38 ^ x6 ;
  assign n176 = ~n171 & ~n175 ;
  assign n178 = x37 ^ x5 ;
  assign n198 = x36 ^ x4 ;
  assign n199 = ~n178 & ~n198 ;
  assign n200 = n176 & n199 ;
  assign n201 = n197 & n200 ;
  assign n179 = x4 & ~x36 ;
  assign n180 = ~n178 & n179 ;
  assign n177 = x5 & ~x37 ;
  assign n181 = n180 ^ n177 ;
  assign n182 = n176 & n181 ;
  assign n172 = x6 & ~x38 ;
  assign n173 = ~n171 & n172 ;
  assign n170 = x7 & ~x39 ;
  assign n174 = n173 ^ n170 ;
  assign n183 = n182 ^ n174 ;
  assign n202 = n201 ^ n183 ;
  assign n138 = x47 ^ x15 ;
  assign n142 = x46 ^ x14 ;
  assign n143 = ~n138 & ~n142 ;
  assign n145 = x45 ^ x13 ;
  assign n151 = x44 ^ x12 ;
  assign n152 = ~n145 & ~n151 ;
  assign n153 = n143 & n152 ;
  assign n155 = x43 ^ x11 ;
  assign n159 = x42 ^ x10 ;
  assign n160 = ~n155 & ~n159 ;
  assign n162 = x41 ^ x9 ;
  assign n203 = x40 ^ x8 ;
  assign n204 = ~n162 & ~n203 ;
  assign n205 = n160 & n204 ;
  assign n206 = n153 & n205 ;
  assign n207 = n202 & n206 ;
  assign n163 = x8 & ~x40 ;
  assign n164 = ~n162 & n163 ;
  assign n161 = x9 & ~x41 ;
  assign n165 = n164 ^ n161 ;
  assign n166 = n160 & n165 ;
  assign n156 = x10 & ~x42 ;
  assign n157 = ~n155 & n156 ;
  assign n154 = x11 & ~x43 ;
  assign n158 = n157 ^ n154 ;
  assign n167 = n166 ^ n158 ;
  assign n168 = n153 & n167 ;
  assign n146 = x12 & ~x44 ;
  assign n147 = ~n145 & n146 ;
  assign n144 = x13 & ~x45 ;
  assign n148 = n147 ^ n144 ;
  assign n149 = n143 & n148 ;
  assign n139 = x14 & ~x46 ;
  assign n140 = ~n138 & n139 ;
  assign n137 = x15 & ~x47 ;
  assign n141 = n140 ^ n137 ;
  assign n150 = n149 ^ n141 ;
  assign n169 = n168 ^ n150 ;
  assign n208 = n207 ^ n169 ;
  assign n66 = x63 ^ x31 ;
  assign n70 = x62 ^ x30 ;
  assign n71 = ~n66 & ~n70 ;
  assign n73 = x61 ^ x29 ;
  assign n79 = x60 ^ x28 ;
  assign n80 = ~n73 & ~n79 ;
  assign n81 = n71 & n80 ;
  assign n83 = x59 ^ x27 ;
  assign n87 = x58 ^ x26 ;
  assign n88 = ~n83 & ~n87 ;
  assign n90 = x57 ^ x25 ;
  assign n98 = x56 ^ x24 ;
  assign n99 = ~n90 & ~n98 ;
  assign n100 = n88 & n99 ;
  assign n101 = n81 & n100 ;
  assign n103 = x55 ^ x23 ;
  assign n107 = x54 ^ x22 ;
  assign n108 = ~n103 & ~n107 ;
  assign n110 = x53 ^ x21 ;
  assign n116 = x52 ^ x20 ;
  assign n117 = ~n110 & ~n116 ;
  assign n118 = n108 & n117 ;
  assign n120 = x51 ^ x19 ;
  assign n124 = x50 ^ x18 ;
  assign n125 = ~n120 & ~n124 ;
  assign n127 = x49 ^ x17 ;
  assign n209 = x48 ^ x16 ;
  assign n210 = ~n127 & ~n209 ;
  assign n211 = n125 & n210 ;
  assign n212 = n118 & n211 ;
  assign n213 = n101 & n212 ;
  assign n214 = n208 & n213 ;
  assign n128 = x16 & ~x48 ;
  assign n129 = ~n127 & n128 ;
  assign n126 = x17 & ~x49 ;
  assign n130 = n129 ^ n126 ;
  assign n131 = n125 & n130 ;
  assign n121 = x18 & ~x50 ;
  assign n122 = ~n120 & n121 ;
  assign n119 = x19 & ~x51 ;
  assign n123 = n122 ^ n119 ;
  assign n132 = n131 ^ n123 ;
  assign n133 = n118 & n132 ;
  assign n111 = x20 & ~x52 ;
  assign n112 = ~n110 & n111 ;
  assign n109 = x21 & ~x53 ;
  assign n113 = n112 ^ n109 ;
  assign n114 = n108 & n113 ;
  assign n104 = x22 & ~x54 ;
  assign n105 = ~n103 & n104 ;
  assign n102 = x23 & ~x55 ;
  assign n106 = n105 ^ n102 ;
  assign n115 = n114 ^ n106 ;
  assign n134 = n133 ^ n115 ;
  assign n135 = n101 & n134 ;
  assign n91 = x24 & ~x56 ;
  assign n92 = ~n90 & n91 ;
  assign n89 = x25 & ~x57 ;
  assign n93 = n92 ^ n89 ;
  assign n94 = n88 & n93 ;
  assign n84 = x26 & ~x58 ;
  assign n85 = ~n83 & n84 ;
  assign n82 = x27 & ~x59 ;
  assign n86 = n85 ^ n82 ;
  assign n95 = n94 ^ n86 ;
  assign n96 = n81 & n95 ;
  assign n74 = x28 & ~x60 ;
  assign n75 = ~n73 & n74 ;
  assign n72 = x29 & ~x61 ;
  assign n76 = n75 ^ n72 ;
  assign n77 = n71 & n76 ;
  assign n67 = x30 & ~x62 ;
  assign n68 = ~n66 & n67 ;
  assign n65 = x31 & ~x63 ;
  assign n69 = n68 ^ n65 ;
  assign n78 = n77 ^ n69 ;
  assign n97 = n96 ^ n78 ;
  assign n136 = n135 ^ n97 ;
  assign n215 = n214 ^ n136 ;
  assign n216 = x32 ^ x0 ;
  assign n217 = n215 & n216 ;
  assign n218 = n217 ^ x32 ;
  assign n219 = n190 & n215 ;
  assign n220 = n219 ^ x33 ;
  assign n221 = n194 & n215 ;
  assign n222 = n221 ^ x34 ;
  assign n223 = n185 & n215 ;
  assign n224 = n223 ^ x35 ;
  assign n225 = n198 & n215 ;
  assign n226 = n225 ^ x36 ;
  assign n227 = n178 & n215 ;
  assign n228 = n227 ^ x37 ;
  assign n229 = n175 & n215 ;
  assign n230 = n229 ^ x38 ;
  assign n231 = n171 & n215 ;
  assign n232 = n231 ^ x39 ;
  assign n233 = n203 & n215 ;
  assign n234 = n233 ^ x40 ;
  assign n235 = n162 & n215 ;
  assign n236 = n235 ^ x41 ;
  assign n237 = n159 & n215 ;
  assign n238 = n237 ^ x42 ;
  assign n239 = n155 & n215 ;
  assign n240 = n239 ^ x43 ;
  assign n241 = n151 & n215 ;
  assign n242 = n241 ^ x44 ;
  assign n243 = n145 & n215 ;
  assign n244 = n243 ^ x45 ;
  assign n245 = n142 & n215 ;
  assign n246 = n245 ^ x46 ;
  assign n247 = n138 & n215 ;
  assign n248 = n247 ^ x47 ;
  assign n249 = n209 & n215 ;
  assign n250 = n249 ^ x48 ;
  assign n251 = n127 & n215 ;
  assign n252 = n251 ^ x49 ;
  assign n253 = n124 & n215 ;
  assign n254 = n253 ^ x50 ;
  assign n255 = n120 & n215 ;
  assign n256 = n255 ^ x51 ;
  assign n257 = n116 & n215 ;
  assign n258 = n257 ^ x52 ;
  assign n259 = n110 & n215 ;
  assign n260 = n259 ^ x53 ;
  assign n261 = n107 & n215 ;
  assign n262 = n261 ^ x54 ;
  assign n263 = n103 & n215 ;
  assign n264 = n263 ^ x55 ;
  assign n265 = n98 & n215 ;
  assign n266 = n265 ^ x56 ;
  assign n267 = n90 & n215 ;
  assign n268 = n267 ^ x57 ;
  assign n269 = n87 & n215 ;
  assign n270 = n269 ^ x58 ;
  assign n271 = n83 & n215 ;
  assign n272 = n271 ^ x59 ;
  assign n273 = n79 & n215 ;
  assign n274 = n273 ^ x60 ;
  assign n275 = n73 & n215 ;
  assign n276 = n275 ^ x61 ;
  assign n277 = n70 & n215 ;
  assign n278 = n277 ^ x62 ;
  assign n279 = n66 & n215 ;
  assign n280 = n279 ^ x63 ;
  assign y0 = n218 ;
  assign y1 = n220 ;
  assign y2 = n222 ;
  assign y3 = n224 ;
  assign y4 = n226 ;
  assign y5 = n228 ;
  assign y6 = n230 ;
  assign y7 = n232 ;
  assign y8 = n234 ;
  assign y9 = n236 ;
  assign y10 = n238 ;
  assign y11 = n240 ;
  assign y12 = n242 ;
  assign y13 = n244 ;
  assign y14 = n246 ;
  assign y15 = n248 ;
  assign y16 = n250 ;
  assign y17 = n252 ;
  assign y18 = n254 ;
  assign y19 = n256 ;
  assign y20 = n258 ;
  assign y21 = n260 ;
  assign y22 = n262 ;
  assign y23 = n264 ;
  assign y24 = n266 ;
  assign y25 = n268 ;
  assign y26 = n270 ;
  assign y27 = n272 ;
  assign y28 = n274 ;
  assign y29 = n276 ;
  assign y30 = n278 ;
  assign y31 = n280 ;
endmodule
