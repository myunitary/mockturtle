module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 ;
  assign n136 = ~x132 & ~x133 ;
  assign n148 = x130 & ~x131 ;
  assign n152 = x60 ^ x59 ;
  assign n153 = x128 & n152 ;
  assign n154 = n153 ^ x60 ;
  assign n149 = x58 ^ x57 ;
  assign n150 = x128 & n149 ;
  assign n151 = n150 ^ x58 ;
  assign n155 = n154 ^ n151 ;
  assign n156 = x129 & n155 ;
  assign n157 = n156 ^ n154 ;
  assign n158 = n148 & n157 ;
  assign n137 = ~x130 & ~x131 ;
  assign n141 = x64 ^ x63 ;
  assign n142 = x128 & n141 ;
  assign n143 = n142 ^ x64 ;
  assign n138 = x62 ^ x61 ;
  assign n139 = x128 & n138 ;
  assign n140 = n139 ^ x62 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = x129 & n144 ;
  assign n146 = n145 ^ n143 ;
  assign n147 = n137 & n146 ;
  assign n159 = n158 ^ n147 ;
  assign n171 = ~x130 & x131 ;
  assign n175 = x56 ^ x55 ;
  assign n176 = x128 & n175 ;
  assign n177 = n176 ^ x56 ;
  assign n172 = x54 ^ x53 ;
  assign n173 = x128 & n172 ;
  assign n174 = n173 ^ x54 ;
  assign n178 = n177 ^ n174 ;
  assign n179 = x129 & n178 ;
  assign n180 = n179 ^ n177 ;
  assign n181 = n171 & n180 ;
  assign n160 = x130 & x131 ;
  assign n164 = x52 ^ x51 ;
  assign n165 = x128 & n164 ;
  assign n166 = n165 ^ x52 ;
  assign n161 = x50 ^ x49 ;
  assign n162 = x128 & n161 ;
  assign n163 = n162 ^ x50 ;
  assign n167 = n166 ^ n163 ;
  assign n168 = x129 & n167 ;
  assign n169 = n168 ^ n166 ;
  assign n170 = n160 & n169 ;
  assign n182 = n181 ^ n170 ;
  assign n183 = ~n159 & ~n182 ;
  assign n184 = n136 & n183 ;
  assign n185 = n184 ^ n136 ;
  assign n197 = x38 & x128 ;
  assign n198 = n197 ^ x38 ;
  assign n196 = x39 & x128 ;
  assign n199 = n198 ^ n196 ;
  assign n200 = x129 & n199 ;
  assign n201 = n200 ^ n199 ;
  assign n202 = n201 ^ n198 ;
  assign n204 = x40 & x128 ;
  assign n205 = n204 ^ x40 ;
  assign n203 = x37 & x128 ;
  assign n206 = n205 ^ n203 ;
  assign n207 = x129 & n206 ;
  assign n208 = n207 ^ n205 ;
  assign n209 = n202 & ~n208 ;
  assign n210 = n209 ^ n208 ;
  assign n211 = n171 & ~n210 ;
  assign n212 = n211 ^ n171 ;
  assign n189 = x36 ^ x35 ;
  assign n190 = x128 & n189 ;
  assign n191 = n190 ^ x36 ;
  assign n186 = x34 ^ x33 ;
  assign n187 = x128 & n186 ;
  assign n188 = n187 ^ x34 ;
  assign n192 = n191 ^ n188 ;
  assign n193 = x129 & n192 ;
  assign n194 = n193 ^ n191 ;
  assign n195 = n160 & n194 ;
  assign n213 = n212 ^ n195 ;
  assign n214 = x132 & ~x133 ;
  assign n226 = n137 & n214 ;
  assign n230 = x48 ^ x47 ;
  assign n231 = x128 & n230 ;
  assign n232 = n231 ^ x48 ;
  assign n227 = x46 ^ x45 ;
  assign n228 = x128 & n227 ;
  assign n229 = n228 ^ x46 ;
  assign n233 = n232 ^ n229 ;
  assign n234 = x129 & n233 ;
  assign n235 = n234 ^ n232 ;
  assign n236 = n226 & n235 ;
  assign n237 = n236 ^ n214 ;
  assign n215 = n148 & n214 ;
  assign n219 = x44 ^ x43 ;
  assign n220 = x128 & n219 ;
  assign n221 = n220 ^ x44 ;
  assign n216 = x42 ^ x41 ;
  assign n217 = x128 & n216 ;
  assign n218 = n217 ^ x42 ;
  assign n222 = n221 ^ n218 ;
  assign n223 = x129 & n222 ;
  assign n224 = n223 ^ n221 ;
  assign n225 = n215 & n224 ;
  assign n238 = n237 ^ n225 ;
  assign n239 = ~n213 & n238 ;
  assign n240 = n239 ^ n214 ;
  assign n241 = n185 & n240 ;
  assign n242 = n241 ^ n185 ;
  assign n243 = n242 ^ n240 ;
  assign n289 = ~x132 & x133 ;
  assign n303 = x28 ^ x27 ;
  assign n304 = x128 & n303 ;
  assign n305 = n304 ^ x28 ;
  assign n300 = x26 ^ x25 ;
  assign n301 = x128 & n300 ;
  assign n302 = n301 ^ x26 ;
  assign n306 = n305 ^ n302 ;
  assign n307 = x129 & n306 ;
  assign n308 = n307 ^ n305 ;
  assign n309 = n148 & n308 ;
  assign n293 = x32 ^ x31 ;
  assign n294 = x128 & n293 ;
  assign n295 = n294 ^ x32 ;
  assign n290 = x30 ^ x29 ;
  assign n291 = x128 & n290 ;
  assign n292 = n291 ^ x30 ;
  assign n296 = n295 ^ n292 ;
  assign n297 = x129 & n296 ;
  assign n298 = n297 ^ n295 ;
  assign n299 = n137 & n298 ;
  assign n310 = n309 ^ n299 ;
  assign n324 = x24 ^ x23 ;
  assign n325 = x128 & n324 ;
  assign n326 = n325 ^ x24 ;
  assign n321 = x22 ^ x21 ;
  assign n322 = x128 & n321 ;
  assign n323 = n322 ^ x22 ;
  assign n327 = n326 ^ n323 ;
  assign n328 = x129 & n327 ;
  assign n329 = n328 ^ n326 ;
  assign n330 = n171 & n329 ;
  assign n314 = x20 ^ x19 ;
  assign n315 = x128 & n314 ;
  assign n316 = n315 ^ x20 ;
  assign n311 = x18 ^ x17 ;
  assign n312 = x128 & n311 ;
  assign n313 = n312 ^ x18 ;
  assign n317 = n316 ^ n313 ;
  assign n318 = x129 & n317 ;
  assign n319 = n318 ^ n316 ;
  assign n320 = n160 & n319 ;
  assign n331 = n330 ^ n320 ;
  assign n332 = ~n310 & ~n331 ;
  assign n333 = n289 & n332 ;
  assign n334 = n333 ^ n289 ;
  assign n244 = x132 & x133 ;
  assign n258 = x12 ^ x11 ;
  assign n259 = x128 & n258 ;
  assign n260 = n259 ^ x12 ;
  assign n255 = x10 ^ x9 ;
  assign n256 = x128 & n255 ;
  assign n257 = n256 ^ x10 ;
  assign n261 = n260 ^ n257 ;
  assign n262 = x129 & n261 ;
  assign n263 = n262 ^ n260 ;
  assign n264 = n148 & n263 ;
  assign n248 = x16 ^ x15 ;
  assign n249 = x128 & n248 ;
  assign n250 = n249 ^ x16 ;
  assign n245 = x14 ^ x13 ;
  assign n246 = x128 & n245 ;
  assign n247 = n246 ^ x14 ;
  assign n251 = n250 ^ n247 ;
  assign n252 = x129 & n251 ;
  assign n253 = n252 ^ n250 ;
  assign n254 = n137 & n253 ;
  assign n265 = n264 ^ n254 ;
  assign n279 = x8 ^ x7 ;
  assign n280 = x128 & n279 ;
  assign n281 = n280 ^ x8 ;
  assign n276 = x6 ^ x5 ;
  assign n277 = x128 & n276 ;
  assign n278 = n277 ^ x6 ;
  assign n282 = n281 ^ n278 ;
  assign n283 = x129 & n282 ;
  assign n284 = n283 ^ n281 ;
  assign n285 = n171 & n284 ;
  assign n269 = x4 ^ x3 ;
  assign n270 = x128 & n269 ;
  assign n271 = n270 ^ x4 ;
  assign n266 = x2 ^ x1 ;
  assign n267 = x128 & n266 ;
  assign n268 = n267 ^ x2 ;
  assign n272 = n271 ^ n268 ;
  assign n273 = x129 & n272 ;
  assign n274 = n273 ^ n271 ;
  assign n275 = n160 & n274 ;
  assign n286 = n285 ^ n275 ;
  assign n287 = ~n265 & ~n286 ;
  assign n288 = n244 & ~n287 ;
  assign n335 = n334 ^ n288 ;
  assign n521 = x134 & ~n335 ;
  assign n522 = ~n243 & n521 ;
  assign n394 = x92 ^ x91 ;
  assign n395 = x128 & n394 ;
  assign n396 = n395 ^ x92 ;
  assign n391 = x90 ^ x89 ;
  assign n392 = x128 & n391 ;
  assign n393 = n392 ^ x90 ;
  assign n397 = n396 ^ n393 ;
  assign n398 = x129 & n397 ;
  assign n399 = n398 ^ n396 ;
  assign n400 = n148 & n399 ;
  assign n384 = x96 ^ x95 ;
  assign n385 = x128 & n384 ;
  assign n386 = n385 ^ x96 ;
  assign n381 = x94 ^ x93 ;
  assign n382 = x128 & n381 ;
  assign n383 = n382 ^ x94 ;
  assign n387 = n386 ^ n383 ;
  assign n388 = x129 & n387 ;
  assign n389 = n388 ^ n386 ;
  assign n390 = n137 & n389 ;
  assign n401 = n400 ^ n390 ;
  assign n415 = x88 ^ x87 ;
  assign n416 = x128 & n415 ;
  assign n417 = n416 ^ x88 ;
  assign n412 = x86 ^ x85 ;
  assign n413 = x128 & n412 ;
  assign n414 = n413 ^ x86 ;
  assign n418 = n417 ^ n414 ;
  assign n419 = x129 & n418 ;
  assign n420 = n419 ^ n417 ;
  assign n421 = n171 & n420 ;
  assign n405 = x84 ^ x83 ;
  assign n406 = x128 & n405 ;
  assign n407 = n406 ^ x84 ;
  assign n402 = x82 ^ x81 ;
  assign n403 = x128 & n402 ;
  assign n404 = n403 ^ x82 ;
  assign n408 = n407 ^ n404 ;
  assign n409 = x129 & n408 ;
  assign n410 = n409 ^ n407 ;
  assign n411 = n160 & n410 ;
  assign n422 = n421 ^ n411 ;
  assign n423 = ~n401 & ~n422 ;
  assign n424 = n289 & n423 ;
  assign n425 = n424 ^ n289 ;
  assign n350 = x76 ^ x75 ;
  assign n351 = x128 & n350 ;
  assign n352 = n351 ^ x76 ;
  assign n347 = x74 ^ x73 ;
  assign n348 = x128 & n347 ;
  assign n349 = n348 ^ x74 ;
  assign n353 = n352 ^ n349 ;
  assign n354 = x129 & n353 ;
  assign n355 = n354 ^ n352 ;
  assign n356 = n148 & n355 ;
  assign n340 = x80 ^ x79 ;
  assign n341 = x128 & n340 ;
  assign n342 = n341 ^ x80 ;
  assign n337 = x78 ^ x77 ;
  assign n338 = x128 & n337 ;
  assign n339 = n338 ^ x78 ;
  assign n343 = n342 ^ n339 ;
  assign n344 = x129 & n343 ;
  assign n345 = n344 ^ n342 ;
  assign n346 = n137 & n345 ;
  assign n357 = n356 ^ n346 ;
  assign n371 = x72 ^ x71 ;
  assign n372 = x128 & n371 ;
  assign n373 = n372 ^ x72 ;
  assign n368 = x70 ^ x69 ;
  assign n369 = x128 & n368 ;
  assign n370 = n369 ^ x70 ;
  assign n374 = n373 ^ n370 ;
  assign n375 = x129 & n374 ;
  assign n376 = n375 ^ n373 ;
  assign n377 = n171 & n376 ;
  assign n361 = x68 ^ x67 ;
  assign n362 = x128 & n361 ;
  assign n363 = n362 ^ x68 ;
  assign n358 = x66 ^ x65 ;
  assign n359 = x128 & n358 ;
  assign n360 = n359 ^ x66 ;
  assign n364 = n363 ^ n360 ;
  assign n365 = x129 & n364 ;
  assign n366 = n365 ^ n363 ;
  assign n367 = n160 & n366 ;
  assign n378 = n377 ^ n367 ;
  assign n379 = ~n357 & ~n378 ;
  assign n380 = n244 & ~n379 ;
  assign n426 = n425 ^ n380 ;
  assign n485 = x108 ^ x107 ;
  assign n486 = x128 & n485 ;
  assign n487 = n486 ^ x108 ;
  assign n482 = x106 ^ x105 ;
  assign n483 = x128 & n482 ;
  assign n484 = n483 ^ x106 ;
  assign n488 = n487 ^ n484 ;
  assign n489 = x129 & n488 ;
  assign n490 = n489 ^ n487 ;
  assign n491 = n148 & n490 ;
  assign n475 = x112 ^ x111 ;
  assign n476 = x128 & n475 ;
  assign n477 = n476 ^ x112 ;
  assign n472 = x110 ^ x109 ;
  assign n473 = x128 & n472 ;
  assign n474 = n473 ^ x110 ;
  assign n478 = n477 ^ n474 ;
  assign n479 = x129 & n478 ;
  assign n480 = n479 ^ n477 ;
  assign n481 = n137 & n480 ;
  assign n492 = n491 ^ n481 ;
  assign n506 = x104 ^ x103 ;
  assign n507 = x128 & n506 ;
  assign n508 = n507 ^ x104 ;
  assign n503 = x102 ^ x101 ;
  assign n504 = x128 & n503 ;
  assign n505 = n504 ^ x102 ;
  assign n509 = n508 ^ n505 ;
  assign n510 = x129 & n509 ;
  assign n511 = n510 ^ n508 ;
  assign n512 = n171 & n511 ;
  assign n496 = x100 ^ x99 ;
  assign n497 = x128 & n496 ;
  assign n498 = n497 ^ x100 ;
  assign n493 = x98 ^ x97 ;
  assign n494 = x128 & n493 ;
  assign n495 = n494 ^ x98 ;
  assign n499 = n498 ^ n495 ;
  assign n500 = x129 & n499 ;
  assign n501 = n500 ^ n498 ;
  assign n502 = n160 & n501 ;
  assign n513 = n512 ^ n502 ;
  assign n514 = ~n492 & ~n513 ;
  assign n515 = n214 & n514 ;
  assign n516 = n515 ^ n214 ;
  assign n441 = x124 ^ x123 ;
  assign n442 = x128 & n441 ;
  assign n443 = n442 ^ x124 ;
  assign n438 = x122 ^ x121 ;
  assign n439 = x128 & n438 ;
  assign n440 = n439 ^ x122 ;
  assign n444 = n443 ^ n440 ;
  assign n445 = x129 & n444 ;
  assign n446 = n445 ^ n443 ;
  assign n447 = n148 & n446 ;
  assign n430 = x127 ^ x0 ;
  assign n431 = x128 & n430 ;
  assign n432 = n431 ^ n430 ;
  assign n433 = n432 ^ x127 ;
  assign n427 = x126 ^ x125 ;
  assign n428 = x128 & n427 ;
  assign n429 = n428 ^ x126 ;
  assign n434 = n433 ^ n429 ;
  assign n435 = x129 & n434 ;
  assign n436 = n435 ^ n433 ;
  assign n437 = n137 & n436 ;
  assign n448 = n447 ^ n437 ;
  assign n462 = x120 ^ x119 ;
  assign n463 = x128 & n462 ;
  assign n464 = n463 ^ x120 ;
  assign n459 = x118 ^ x117 ;
  assign n460 = x128 & n459 ;
  assign n461 = n460 ^ x118 ;
  assign n465 = n464 ^ n461 ;
  assign n466 = x129 & n465 ;
  assign n467 = n466 ^ n464 ;
  assign n468 = n171 & n467 ;
  assign n452 = x116 ^ x115 ;
  assign n453 = x128 & n452 ;
  assign n454 = n453 ^ x116 ;
  assign n449 = x114 ^ x113 ;
  assign n450 = x128 & n449 ;
  assign n451 = n450 ^ x114 ;
  assign n455 = n454 ^ n451 ;
  assign n456 = x129 & n455 ;
  assign n457 = n456 ^ n454 ;
  assign n458 = n160 & n457 ;
  assign n469 = n468 ^ n458 ;
  assign n470 = ~n448 & ~n469 ;
  assign n471 = n136 & ~n470 ;
  assign n517 = n516 ^ n471 ;
  assign n518 = ~n426 & ~n517 ;
  assign n520 = x134 & n518 ;
  assign n523 = n522 ^ n520 ;
  assign n336 = ~n243 & ~n335 ;
  assign n519 = n518 ^ n336 ;
  assign n524 = n523 ^ n519 ;
  assign n525 = n524 ^ n336 ;
  assign n898 = x11 & x128 ;
  assign n899 = n898 ^ x11 ;
  assign n897 = x12 & x128 ;
  assign n900 = n899 ^ n897 ;
  assign n901 = x129 & n900 ;
  assign n902 = n901 ^ n900 ;
  assign n903 = n902 ^ n899 ;
  assign n905 = x13 & x128 ;
  assign n906 = n905 ^ x13 ;
  assign n904 = x10 & x128 ;
  assign n907 = n906 ^ n904 ;
  assign n908 = x129 & n907 ;
  assign n909 = n908 ^ n906 ;
  assign n910 = n903 & ~n909 ;
  assign n911 = n910 ^ n909 ;
  assign n912 = n148 & ~n911 ;
  assign n913 = n912 ^ n148 ;
  assign n882 = x15 & x128 ;
  assign n883 = n882 ^ x15 ;
  assign n881 = x16 & x128 ;
  assign n884 = n883 ^ n881 ;
  assign n885 = x129 & n884 ;
  assign n886 = n885 ^ n884 ;
  assign n887 = n886 ^ n883 ;
  assign n889 = x17 & x128 ;
  assign n890 = n889 ^ x17 ;
  assign n888 = x14 & x128 ;
  assign n891 = n890 ^ n888 ;
  assign n892 = x129 & n891 ;
  assign n893 = n892 ^ n890 ;
  assign n894 = n887 & ~n893 ;
  assign n895 = n894 ^ n893 ;
  assign n896 = n137 & n895 ;
  assign n914 = n913 ^ n896 ;
  assign n932 = x7 & x128 ;
  assign n933 = n932 ^ x7 ;
  assign n931 = x8 & x128 ;
  assign n934 = n933 ^ n931 ;
  assign n935 = x129 & n934 ;
  assign n936 = n935 ^ n934 ;
  assign n937 = n936 ^ n933 ;
  assign n939 = x9 & x128 ;
  assign n940 = n939 ^ x9 ;
  assign n938 = x6 & x128 ;
  assign n941 = n940 ^ n938 ;
  assign n942 = x129 & n941 ;
  assign n943 = n942 ^ n940 ;
  assign n944 = n937 & ~n943 ;
  assign n945 = n944 ^ n943 ;
  assign n946 = n171 & ~n945 ;
  assign n947 = n946 ^ n171 ;
  assign n916 = x3 & x128 ;
  assign n917 = n916 ^ x3 ;
  assign n915 = x4 & x128 ;
  assign n918 = n917 ^ n915 ;
  assign n919 = x129 & n918 ;
  assign n920 = n919 ^ n918 ;
  assign n921 = n920 ^ n917 ;
  assign n923 = x5 & x128 ;
  assign n924 = n923 ^ x5 ;
  assign n922 = x2 & x128 ;
  assign n925 = n924 ^ n922 ;
  assign n926 = x129 & n925 ;
  assign n927 = n926 ^ n924 ;
  assign n928 = n921 & ~n927 ;
  assign n929 = n928 ^ n927 ;
  assign n930 = n160 & n929 ;
  assign n948 = n947 ^ n930 ;
  assign n949 = ~n914 & ~n948 ;
  assign n950 = n244 & n949 ;
  assign n951 = n950 ^ n244 ;
  assign n828 = x59 & x128 ;
  assign n829 = n828 ^ x59 ;
  assign n827 = x60 & x128 ;
  assign n830 = n829 ^ n827 ;
  assign n831 = x129 & n830 ;
  assign n832 = n831 ^ n830 ;
  assign n833 = n832 ^ n829 ;
  assign n835 = x61 & x128 ;
  assign n836 = n835 ^ x61 ;
  assign n834 = x58 & x128 ;
  assign n837 = n836 ^ n834 ;
  assign n838 = x129 & n837 ;
  assign n839 = n838 ^ n836 ;
  assign n840 = n833 & ~n839 ;
  assign n841 = n840 ^ n839 ;
  assign n842 = n148 & ~n841 ;
  assign n843 = n842 ^ n148 ;
  assign n812 = x63 & x128 ;
  assign n813 = n812 ^ x63 ;
  assign n811 = x64 & x128 ;
  assign n814 = n813 ^ n811 ;
  assign n815 = x129 & n814 ;
  assign n816 = n815 ^ n814 ;
  assign n817 = n816 ^ n813 ;
  assign n819 = x65 & x128 ;
  assign n820 = n819 ^ x65 ;
  assign n818 = x62 & x128 ;
  assign n821 = n820 ^ n818 ;
  assign n822 = x129 & n821 ;
  assign n823 = n822 ^ n820 ;
  assign n824 = n817 & ~n823 ;
  assign n825 = n824 ^ n823 ;
  assign n826 = n137 & n825 ;
  assign n844 = n843 ^ n826 ;
  assign n862 = x55 & x128 ;
  assign n863 = n862 ^ x55 ;
  assign n861 = x56 & x128 ;
  assign n864 = n863 ^ n861 ;
  assign n865 = x129 & n864 ;
  assign n866 = n865 ^ n864 ;
  assign n867 = n866 ^ n863 ;
  assign n869 = x57 & x128 ;
  assign n870 = n869 ^ x57 ;
  assign n868 = x54 & x128 ;
  assign n871 = n870 ^ n868 ;
  assign n872 = x129 & n871 ;
  assign n873 = n872 ^ n870 ;
  assign n874 = n867 & ~n873 ;
  assign n875 = n874 ^ n873 ;
  assign n876 = n171 & ~n875 ;
  assign n877 = n876 ^ n171 ;
  assign n846 = x51 & x128 ;
  assign n847 = n846 ^ x51 ;
  assign n845 = x52 & x128 ;
  assign n848 = n847 ^ n845 ;
  assign n849 = x129 & n848 ;
  assign n850 = n849 ^ n848 ;
  assign n851 = n850 ^ n847 ;
  assign n853 = x53 & x128 ;
  assign n854 = n853 ^ x53 ;
  assign n852 = x50 & x128 ;
  assign n855 = n854 ^ n852 ;
  assign n856 = x129 & n855 ;
  assign n857 = n856 ^ n854 ;
  assign n858 = n851 & ~n857 ;
  assign n859 = n858 ^ n857 ;
  assign n860 = n160 & n859 ;
  assign n878 = n877 ^ n860 ;
  assign n879 = ~n844 & ~n878 ;
  assign n880 = n136 & ~n879 ;
  assign n952 = n951 ^ n880 ;
  assign n1039 = x27 & x128 ;
  assign n1040 = n1039 ^ x27 ;
  assign n1038 = x28 & x128 ;
  assign n1041 = n1040 ^ n1038 ;
  assign n1042 = x129 & n1041 ;
  assign n1043 = n1042 ^ n1041 ;
  assign n1044 = n1043 ^ n1040 ;
  assign n1046 = x29 & x128 ;
  assign n1047 = n1046 ^ x29 ;
  assign n1045 = x26 & x128 ;
  assign n1048 = n1047 ^ n1045 ;
  assign n1049 = x129 & n1048 ;
  assign n1050 = n1049 ^ n1047 ;
  assign n1051 = n1044 & ~n1050 ;
  assign n1052 = n1051 ^ n1050 ;
  assign n1053 = n148 & ~n1052 ;
  assign n1054 = n1053 ^ n148 ;
  assign n1023 = x31 & x128 ;
  assign n1024 = n1023 ^ x31 ;
  assign n1022 = x32 & x128 ;
  assign n1025 = n1024 ^ n1022 ;
  assign n1026 = x129 & n1025 ;
  assign n1027 = n1026 ^ n1025 ;
  assign n1028 = n1027 ^ n1024 ;
  assign n1030 = x33 & x128 ;
  assign n1031 = n1030 ^ x33 ;
  assign n1029 = x30 & x128 ;
  assign n1032 = n1031 ^ n1029 ;
  assign n1033 = x129 & n1032 ;
  assign n1034 = n1033 ^ n1031 ;
  assign n1035 = n1028 & ~n1034 ;
  assign n1036 = n1035 ^ n1034 ;
  assign n1037 = n137 & n1036 ;
  assign n1055 = n1054 ^ n1037 ;
  assign n1073 = x23 & x128 ;
  assign n1074 = n1073 ^ x23 ;
  assign n1072 = x24 & x128 ;
  assign n1075 = n1074 ^ n1072 ;
  assign n1076 = x129 & n1075 ;
  assign n1077 = n1076 ^ n1075 ;
  assign n1078 = n1077 ^ n1074 ;
  assign n1080 = x25 & x128 ;
  assign n1081 = n1080 ^ x25 ;
  assign n1079 = x22 & x128 ;
  assign n1082 = n1081 ^ n1079 ;
  assign n1083 = x129 & n1082 ;
  assign n1084 = n1083 ^ n1081 ;
  assign n1085 = n1078 & ~n1084 ;
  assign n1086 = n1085 ^ n1084 ;
  assign n1087 = n171 & ~n1086 ;
  assign n1088 = n1087 ^ n171 ;
  assign n1057 = x19 & x128 ;
  assign n1058 = n1057 ^ x19 ;
  assign n1056 = x20 & x128 ;
  assign n1059 = n1058 ^ n1056 ;
  assign n1060 = x129 & n1059 ;
  assign n1061 = n1060 ^ n1059 ;
  assign n1062 = n1061 ^ n1058 ;
  assign n1064 = x21 & x128 ;
  assign n1065 = n1064 ^ x21 ;
  assign n1063 = x18 & x128 ;
  assign n1066 = n1065 ^ n1063 ;
  assign n1067 = x129 & n1066 ;
  assign n1068 = n1067 ^ n1065 ;
  assign n1069 = n1062 & ~n1068 ;
  assign n1070 = n1069 ^ n1068 ;
  assign n1071 = n160 & n1070 ;
  assign n1089 = n1088 ^ n1071 ;
  assign n1090 = ~n1055 & ~n1089 ;
  assign n1091 = n289 & n1090 ;
  assign n1092 = n1091 ^ n289 ;
  assign n966 = x47 & x128 ;
  assign n967 = n966 ^ x47 ;
  assign n965 = x48 & x128 ;
  assign n968 = n967 ^ n965 ;
  assign n969 = x129 & n968 ;
  assign n970 = n969 ^ n968 ;
  assign n971 = n970 ^ n967 ;
  assign n973 = x49 & x128 ;
  assign n974 = n973 ^ x49 ;
  assign n972 = x46 & x128 ;
  assign n975 = n974 ^ n972 ;
  assign n976 = x129 & n975 ;
  assign n977 = n976 ^ n974 ;
  assign n978 = n971 & ~n977 ;
  assign n979 = n978 ^ n977 ;
  assign n956 = x45 ^ x44 ;
  assign n957 = x128 & n956 ;
  assign n958 = n957 ^ x45 ;
  assign n953 = x43 ^ x42 ;
  assign n954 = x128 & n953 ;
  assign n955 = n954 ^ x43 ;
  assign n959 = n958 ^ n955 ;
  assign n960 = x129 & ~n959 ;
  assign n961 = n960 ^ x129 ;
  assign n962 = n961 ^ n958 ;
  assign n982 = n137 & n148 ;
  assign n983 = n962 & n982 ;
  assign n984 = n979 & n983 ;
  assign n980 = n137 & ~n979 ;
  assign n981 = n980 ^ n137 ;
  assign n985 = n984 ^ n981 ;
  assign n963 = n148 & ~n962 ;
  assign n964 = n963 ^ n148 ;
  assign n986 = n985 ^ n964 ;
  assign n1000 = x35 & x128 ;
  assign n1001 = n1000 ^ x35 ;
  assign n999 = x36 & x128 ;
  assign n1002 = n1001 ^ n999 ;
  assign n1003 = x129 & n1002 ;
  assign n1004 = n1003 ^ n1002 ;
  assign n1005 = n1004 ^ n1001 ;
  assign n1007 = n203 ^ x37 ;
  assign n1006 = x34 & x128 ;
  assign n1008 = n1007 ^ n1006 ;
  assign n1009 = x129 & n1008 ;
  assign n1010 = n1009 ^ n1007 ;
  assign n1011 = n1005 & ~n1010 ;
  assign n1012 = n1011 ^ n1010 ;
  assign n990 = x39 ^ x38 ;
  assign n991 = x128 & n990 ;
  assign n992 = n991 ^ x39 ;
  assign n987 = x41 ^ x40 ;
  assign n988 = x128 & n987 ;
  assign n989 = n988 ^ x41 ;
  assign n993 = n992 ^ n989 ;
  assign n994 = x129 & n993 ;
  assign n995 = n994 ^ n993 ;
  assign n996 = n995 ^ n992 ;
  assign n1015 = n160 & n171 ;
  assign n1016 = n996 & n1015 ;
  assign n1017 = n1012 & n1016 ;
  assign n1013 = n160 & ~n1012 ;
  assign n1014 = n1013 ^ n160 ;
  assign n1018 = n1017 ^ n1014 ;
  assign n997 = n171 & ~n996 ;
  assign n998 = n997 ^ n171 ;
  assign n1019 = n1018 ^ n998 ;
  assign n1020 = ~n986 & ~n1019 ;
  assign n1021 = n214 & ~n1020 ;
  assign n1093 = n1092 ^ n1021 ;
  assign n1094 = ~n952 & ~n1093 ;
  assign n613 = x91 & x128 ;
  assign n614 = n613 ^ x91 ;
  assign n612 = x92 & x128 ;
  assign n615 = n614 ^ n612 ;
  assign n616 = x129 & n615 ;
  assign n617 = n616 ^ n615 ;
  assign n618 = n617 ^ n614 ;
  assign n620 = x93 & x128 ;
  assign n621 = n620 ^ x93 ;
  assign n619 = x90 & x128 ;
  assign n622 = n621 ^ n619 ;
  assign n623 = x129 & n622 ;
  assign n624 = n623 ^ n621 ;
  assign n625 = n618 & ~n624 ;
  assign n626 = n625 ^ n624 ;
  assign n627 = n148 & ~n626 ;
  assign n628 = n627 ^ n148 ;
  assign n597 = x95 & x128 ;
  assign n598 = n597 ^ x95 ;
  assign n596 = x96 & x128 ;
  assign n599 = n598 ^ n596 ;
  assign n600 = x129 & n599 ;
  assign n601 = n600 ^ n599 ;
  assign n602 = n601 ^ n598 ;
  assign n604 = x97 & x128 ;
  assign n605 = n604 ^ x97 ;
  assign n603 = x94 & x128 ;
  assign n606 = n605 ^ n603 ;
  assign n607 = x129 & n606 ;
  assign n608 = n607 ^ n605 ;
  assign n609 = n602 & ~n608 ;
  assign n610 = n609 ^ n608 ;
  assign n611 = n137 & n610 ;
  assign n629 = n628 ^ n611 ;
  assign n647 = x87 & x128 ;
  assign n648 = n647 ^ x87 ;
  assign n646 = x88 & x128 ;
  assign n649 = n648 ^ n646 ;
  assign n650 = x129 & n649 ;
  assign n651 = n650 ^ n649 ;
  assign n652 = n651 ^ n648 ;
  assign n654 = x89 & x128 ;
  assign n655 = n654 ^ x89 ;
  assign n653 = x86 & x128 ;
  assign n656 = n655 ^ n653 ;
  assign n657 = x129 & n656 ;
  assign n658 = n657 ^ n655 ;
  assign n659 = n652 & ~n658 ;
  assign n660 = n659 ^ n658 ;
  assign n661 = n171 & ~n660 ;
  assign n662 = n661 ^ n171 ;
  assign n631 = x83 & x128 ;
  assign n632 = n631 ^ x83 ;
  assign n630 = x84 & x128 ;
  assign n633 = n632 ^ n630 ;
  assign n634 = x129 & n633 ;
  assign n635 = n634 ^ n633 ;
  assign n636 = n635 ^ n632 ;
  assign n638 = x85 & x128 ;
  assign n639 = n638 ^ x85 ;
  assign n637 = x82 & x128 ;
  assign n640 = n639 ^ n637 ;
  assign n641 = x129 & n640 ;
  assign n642 = n641 ^ n639 ;
  assign n643 = n636 & ~n642 ;
  assign n644 = n643 ^ n642 ;
  assign n645 = n160 & n644 ;
  assign n663 = n662 ^ n645 ;
  assign n664 = ~n629 & ~n663 ;
  assign n665 = n289 & n664 ;
  assign n666 = n665 ^ n289 ;
  assign n543 = x75 & x128 ;
  assign n544 = n543 ^ x75 ;
  assign n542 = x76 & x128 ;
  assign n545 = n544 ^ n542 ;
  assign n546 = x129 & n545 ;
  assign n547 = n546 ^ n545 ;
  assign n548 = n547 ^ n544 ;
  assign n550 = x77 & x128 ;
  assign n551 = n550 ^ x77 ;
  assign n549 = x74 & x128 ;
  assign n552 = n551 ^ n549 ;
  assign n553 = x129 & n552 ;
  assign n554 = n553 ^ n551 ;
  assign n555 = n548 & ~n554 ;
  assign n556 = n555 ^ n554 ;
  assign n557 = n148 & ~n556 ;
  assign n558 = n557 ^ n148 ;
  assign n527 = x79 & x128 ;
  assign n528 = n527 ^ x79 ;
  assign n526 = x80 & x128 ;
  assign n529 = n528 ^ n526 ;
  assign n530 = x129 & n529 ;
  assign n531 = n530 ^ n529 ;
  assign n532 = n531 ^ n528 ;
  assign n534 = x81 & x128 ;
  assign n535 = n534 ^ x81 ;
  assign n533 = x78 & x128 ;
  assign n536 = n535 ^ n533 ;
  assign n537 = x129 & n536 ;
  assign n538 = n537 ^ n535 ;
  assign n539 = n532 & ~n538 ;
  assign n540 = n539 ^ n538 ;
  assign n541 = n137 & n540 ;
  assign n559 = n558 ^ n541 ;
  assign n577 = x71 & x128 ;
  assign n578 = n577 ^ x71 ;
  assign n576 = x72 & x128 ;
  assign n579 = n578 ^ n576 ;
  assign n580 = x129 & n579 ;
  assign n581 = n580 ^ n579 ;
  assign n582 = n581 ^ n578 ;
  assign n584 = x73 & x128 ;
  assign n585 = n584 ^ x73 ;
  assign n583 = x70 & x128 ;
  assign n586 = n585 ^ n583 ;
  assign n587 = x129 & n586 ;
  assign n588 = n587 ^ n585 ;
  assign n589 = n582 & ~n588 ;
  assign n590 = n589 ^ n588 ;
  assign n591 = n171 & ~n590 ;
  assign n592 = n591 ^ n171 ;
  assign n561 = x67 & x128 ;
  assign n562 = n561 ^ x67 ;
  assign n560 = x68 & x128 ;
  assign n563 = n562 ^ n560 ;
  assign n564 = x129 & n563 ;
  assign n565 = n564 ^ n563 ;
  assign n566 = n565 ^ n562 ;
  assign n568 = x69 & x128 ;
  assign n569 = n568 ^ x69 ;
  assign n567 = x66 & x128 ;
  assign n570 = n569 ^ n567 ;
  assign n571 = x129 & n570 ;
  assign n572 = n571 ^ n569 ;
  assign n573 = n566 & ~n572 ;
  assign n574 = n573 ^ n572 ;
  assign n575 = n160 & n574 ;
  assign n593 = n592 ^ n575 ;
  assign n594 = ~n559 & ~n593 ;
  assign n595 = n244 & ~n594 ;
  assign n667 = n666 ^ n595 ;
  assign n755 = x107 & x128 ;
  assign n756 = n755 ^ x107 ;
  assign n754 = x108 & x128 ;
  assign n757 = n756 ^ n754 ;
  assign n758 = x129 & n757 ;
  assign n759 = n758 ^ n757 ;
  assign n760 = n759 ^ n756 ;
  assign n762 = x109 & x128 ;
  assign n763 = n762 ^ x109 ;
  assign n761 = x106 & x128 ;
  assign n764 = n763 ^ n761 ;
  assign n765 = x129 & n764 ;
  assign n766 = n765 ^ n763 ;
  assign n767 = n760 & ~n766 ;
  assign n768 = n767 ^ n766 ;
  assign n769 = n148 & ~n768 ;
  assign n770 = n769 ^ n148 ;
  assign n739 = x111 & x128 ;
  assign n740 = n739 ^ x111 ;
  assign n738 = x112 & x128 ;
  assign n741 = n740 ^ n738 ;
  assign n742 = x129 & n741 ;
  assign n743 = n742 ^ n741 ;
  assign n744 = n743 ^ n740 ;
  assign n746 = x113 & x128 ;
  assign n747 = n746 ^ x113 ;
  assign n745 = x110 & x128 ;
  assign n748 = n747 ^ n745 ;
  assign n749 = x129 & n748 ;
  assign n750 = n749 ^ n747 ;
  assign n751 = n744 & ~n750 ;
  assign n752 = n751 ^ n750 ;
  assign n753 = n137 & n752 ;
  assign n771 = n770 ^ n753 ;
  assign n789 = x103 & x128 ;
  assign n790 = n789 ^ x103 ;
  assign n788 = x104 & x128 ;
  assign n791 = n790 ^ n788 ;
  assign n792 = x129 & n791 ;
  assign n793 = n792 ^ n791 ;
  assign n794 = n793 ^ n790 ;
  assign n796 = x105 & x128 ;
  assign n797 = n796 ^ x105 ;
  assign n795 = x102 & x128 ;
  assign n798 = n797 ^ n795 ;
  assign n799 = x129 & n798 ;
  assign n800 = n799 ^ n797 ;
  assign n801 = n794 & ~n800 ;
  assign n802 = n801 ^ n800 ;
  assign n803 = n171 & ~n802 ;
  assign n804 = n803 ^ n171 ;
  assign n773 = x99 & x128 ;
  assign n774 = n773 ^ x99 ;
  assign n772 = x100 & x128 ;
  assign n775 = n774 ^ n772 ;
  assign n776 = x129 & n775 ;
  assign n777 = n776 ^ n775 ;
  assign n778 = n777 ^ n774 ;
  assign n780 = x101 & x128 ;
  assign n781 = n780 ^ x101 ;
  assign n779 = x98 & x128 ;
  assign n782 = n781 ^ n779 ;
  assign n783 = x129 & n782 ;
  assign n784 = n783 ^ n781 ;
  assign n785 = n778 & ~n784 ;
  assign n786 = n785 ^ n784 ;
  assign n787 = n160 & n786 ;
  assign n805 = n804 ^ n787 ;
  assign n806 = ~n771 & ~n805 ;
  assign n807 = n214 & n806 ;
  assign n808 = n807 ^ n214 ;
  assign n685 = x123 & x128 ;
  assign n686 = n685 ^ x123 ;
  assign n684 = x124 & x128 ;
  assign n687 = n686 ^ n684 ;
  assign n688 = x129 & n687 ;
  assign n689 = n688 ^ n687 ;
  assign n690 = n689 ^ n686 ;
  assign n692 = x125 & x128 ;
  assign n693 = n692 ^ x125 ;
  assign n691 = x122 & x128 ;
  assign n694 = n693 ^ n691 ;
  assign n695 = x129 & n694 ;
  assign n696 = n695 ^ n693 ;
  assign n697 = n690 & ~n696 ;
  assign n698 = n697 ^ n696 ;
  assign n699 = n148 & ~n698 ;
  assign n700 = n699 ^ n148 ;
  assign n669 = x127 & x128 ;
  assign n670 = n669 ^ x127 ;
  assign n668 = x0 & x128 ;
  assign n671 = n670 ^ n668 ;
  assign n672 = x129 & n671 ;
  assign n673 = n672 ^ n671 ;
  assign n674 = n673 ^ n670 ;
  assign n676 = x1 & x128 ;
  assign n677 = n676 ^ x1 ;
  assign n675 = x126 & x128 ;
  assign n678 = n677 ^ n675 ;
  assign n679 = x129 & n678 ;
  assign n680 = n679 ^ n677 ;
  assign n681 = n674 & ~n680 ;
  assign n682 = n681 ^ n680 ;
  assign n683 = n137 & n682 ;
  assign n701 = n700 ^ n683 ;
  assign n719 = x119 & x128 ;
  assign n720 = n719 ^ x119 ;
  assign n718 = x120 & x128 ;
  assign n721 = n720 ^ n718 ;
  assign n722 = x129 & n721 ;
  assign n723 = n722 ^ n721 ;
  assign n724 = n723 ^ n720 ;
  assign n726 = x121 & x128 ;
  assign n727 = n726 ^ x121 ;
  assign n725 = x118 & x128 ;
  assign n728 = n727 ^ n725 ;
  assign n729 = x129 & n728 ;
  assign n730 = n729 ^ n727 ;
  assign n731 = n724 & ~n730 ;
  assign n732 = n731 ^ n730 ;
  assign n733 = n171 & ~n732 ;
  assign n734 = n733 ^ n171 ;
  assign n703 = x115 & x128 ;
  assign n704 = n703 ^ x115 ;
  assign n702 = x116 & x128 ;
  assign n705 = n704 ^ n702 ;
  assign n706 = x129 & n705 ;
  assign n707 = n706 ^ n705 ;
  assign n708 = n707 ^ n704 ;
  assign n710 = x117 & x128 ;
  assign n711 = n710 ^ x117 ;
  assign n709 = x114 & x128 ;
  assign n712 = n711 ^ n709 ;
  assign n713 = x129 & n712 ;
  assign n714 = n713 ^ n711 ;
  assign n715 = n708 & ~n714 ;
  assign n716 = n715 ^ n714 ;
  assign n717 = n160 & n716 ;
  assign n735 = n734 ^ n717 ;
  assign n736 = ~n701 & ~n735 ;
  assign n737 = n136 & ~n736 ;
  assign n809 = n808 ^ n737 ;
  assign n810 = ~n667 & ~n809 ;
  assign n1095 = n1094 ^ n810 ;
  assign n1096 = x134 & n1095 ;
  assign n1097 = n1096 ^ n1095 ;
  assign n1098 = n1097 ^ n1094 ;
  assign n1220 = n260 ^ n247 ;
  assign n1221 = x129 & n1220 ;
  assign n1222 = n1221 ^ n1220 ;
  assign n1223 = n1222 ^ n260 ;
  assign n1224 = n148 & n1223 ;
  assign n1216 = n313 ^ n250 ;
  assign n1217 = x129 & n1216 ;
  assign n1218 = n1217 ^ n313 ;
  assign n1219 = n137 & n1218 ;
  assign n1225 = n1224 ^ n1219 ;
  assign n1230 = n281 ^ n257 ;
  assign n1231 = x129 & n1230 ;
  assign n1232 = n1231 ^ n1230 ;
  assign n1233 = n1232 ^ n281 ;
  assign n1234 = n171 & n1233 ;
  assign n1226 = n278 ^ n271 ;
  assign n1227 = x129 & n1226 ;
  assign n1228 = n1227 ^ n278 ;
  assign n1229 = n160 & n1228 ;
  assign n1235 = n1234 ^ n1229 ;
  assign n1236 = ~n1225 & ~n1235 ;
  assign n1237 = n244 & n1236 ;
  assign n1238 = n1237 ^ n244 ;
  assign n1198 = n154 ^ n140 ;
  assign n1199 = x129 & n1198 ;
  assign n1200 = n1199 ^ n1198 ;
  assign n1201 = n1200 ^ n154 ;
  assign n1202 = n148 & n1201 ;
  assign n1193 = n360 ^ n143 ;
  assign n1194 = x129 & n1193 ;
  assign n1195 = n1194 ^ n1193 ;
  assign n1196 = n1195 ^ n143 ;
  assign n1197 = n137 & n1196 ;
  assign n1203 = n1202 ^ n1197 ;
  assign n1208 = n177 ^ n151 ;
  assign n1209 = x129 & n1208 ;
  assign n1210 = n1209 ^ n1208 ;
  assign n1211 = n1210 ^ n177 ;
  assign n1212 = n171 & n1211 ;
  assign n1204 = n174 ^ n166 ;
  assign n1205 = x129 & n1204 ;
  assign n1206 = n1205 ^ n174 ;
  assign n1207 = n160 & n1206 ;
  assign n1213 = n1212 ^ n1207 ;
  assign n1214 = ~n1203 & ~n1213 ;
  assign n1215 = n136 & ~n1214 ;
  assign n1239 = n1238 ^ n1215 ;
  assign n1276 = n305 ^ n292 ;
  assign n1277 = x129 & n1276 ;
  assign n1278 = n1277 ^ n1276 ;
  assign n1279 = n1278 ^ n305 ;
  assign n1280 = n148 & n1279 ;
  assign n1272 = n295 ^ n188 ;
  assign n1273 = x129 & n1272 ;
  assign n1274 = n1273 ^ n188 ;
  assign n1275 = n137 & n1274 ;
  assign n1281 = n1280 ^ n1275 ;
  assign n1286 = n326 ^ n302 ;
  assign n1287 = x129 & n1286 ;
  assign n1288 = n1287 ^ n1286 ;
  assign n1289 = n1288 ^ n326 ;
  assign n1290 = n171 & n1289 ;
  assign n1282 = n323 ^ n316 ;
  assign n1283 = x129 & n1282 ;
  assign n1284 = n1283 ^ n323 ;
  assign n1285 = n160 & n1284 ;
  assign n1291 = n1290 ^ n1285 ;
  assign n1292 = ~n1281 & ~n1291 ;
  assign n1293 = n289 & n1292 ;
  assign n1294 = n1293 ^ n289 ;
  assign n1245 = n229 ^ n221 ;
  assign n1246 = x129 & n1245 ;
  assign n1247 = n1246 ^ n1245 ;
  assign n1248 = n1247 ^ n221 ;
  assign n1249 = n148 & n1248 ;
  assign n1240 = n232 ^ n163 ;
  assign n1241 = x129 & n1240 ;
  assign n1242 = n1241 ^ n1240 ;
  assign n1243 = n1242 ^ n232 ;
  assign n1244 = n137 & n1243 ;
  assign n1250 = n1249 ^ n1244 ;
  assign n1259 = x40 ^ x39 ;
  assign n1260 = x128 & n1259 ;
  assign n1261 = n1260 ^ x40 ;
  assign n1262 = n1261 ^ n218 ;
  assign n1263 = x129 & ~n1262 ;
  assign n1264 = n1263 ^ x129 ;
  assign n1265 = n1264 ^ n1262 ;
  assign n1266 = n1265 ^ n1261 ;
  assign n1267 = n171 & ~n1266 ;
  assign n1268 = n1267 ^ n171 ;
  assign n1251 = x38 ^ x37 ;
  assign n1252 = x128 & n1251 ;
  assign n1253 = n1252 ^ x38 ;
  assign n1254 = n1253 ^ n191 ;
  assign n1255 = x129 & ~n1254 ;
  assign n1256 = n1255 ^ x129 ;
  assign n1257 = n1256 ^ n1253 ;
  assign n1258 = n160 & n1257 ;
  assign n1269 = n1268 ^ n1258 ;
  assign n1270 = ~n1250 & ~n1269 ;
  assign n1271 = n214 & ~n1270 ;
  assign n1295 = n1294 ^ n1271 ;
  assign n1296 = ~n1239 & ~n1295 ;
  assign n1125 = n396 ^ n383 ;
  assign n1126 = x129 & n1125 ;
  assign n1127 = n1126 ^ n1125 ;
  assign n1128 = n1127 ^ n396 ;
  assign n1129 = n148 & n1128 ;
  assign n1121 = n495 ^ n386 ;
  assign n1122 = x129 & n1121 ;
  assign n1123 = n1122 ^ n495 ;
  assign n1124 = n137 & n1123 ;
  assign n1130 = n1129 ^ n1124 ;
  assign n1135 = n417 ^ n393 ;
  assign n1136 = x129 & n1135 ;
  assign n1137 = n1136 ^ n1135 ;
  assign n1138 = n1137 ^ n417 ;
  assign n1139 = n171 & n1138 ;
  assign n1131 = n414 ^ n407 ;
  assign n1132 = x129 & n1131 ;
  assign n1133 = n1132 ^ n414 ;
  assign n1134 = n160 & n1133 ;
  assign n1140 = n1139 ^ n1134 ;
  assign n1141 = ~n1130 & ~n1140 ;
  assign n1142 = n289 & n1141 ;
  assign n1143 = n1142 ^ n289 ;
  assign n1103 = n352 ^ n339 ;
  assign n1104 = x129 & n1103 ;
  assign n1105 = n1104 ^ n1103 ;
  assign n1106 = n1105 ^ n352 ;
  assign n1107 = n148 & n1106 ;
  assign n1099 = n404 ^ n342 ;
  assign n1100 = x129 & n1099 ;
  assign n1101 = n1100 ^ n404 ;
  assign n1102 = n137 & n1101 ;
  assign n1108 = n1107 ^ n1102 ;
  assign n1113 = n373 ^ n349 ;
  assign n1114 = x129 & n1113 ;
  assign n1115 = n1114 ^ n1113 ;
  assign n1116 = n1115 ^ n373 ;
  assign n1117 = n171 & n1116 ;
  assign n1109 = n370 ^ n363 ;
  assign n1110 = x129 & n1109 ;
  assign n1111 = n1110 ^ n370 ;
  assign n1112 = n160 & n1111 ;
  assign n1118 = n1117 ^ n1112 ;
  assign n1119 = ~n1108 & ~n1118 ;
  assign n1120 = n244 & ~n1119 ;
  assign n1144 = n1143 ^ n1120 ;
  assign n1172 = n487 ^ n474 ;
  assign n1173 = x129 & n1172 ;
  assign n1174 = n1173 ^ n1172 ;
  assign n1175 = n1174 ^ n487 ;
  assign n1176 = n148 & n1175 ;
  assign n1167 = n477 ^ n451 ;
  assign n1168 = x129 & n1167 ;
  assign n1169 = n1168 ^ n1167 ;
  assign n1170 = n1169 ^ n477 ;
  assign n1171 = n137 & n1170 ;
  assign n1177 = n1176 ^ n1171 ;
  assign n1182 = n508 ^ n484 ;
  assign n1183 = x129 & n1182 ;
  assign n1184 = n1183 ^ n1182 ;
  assign n1185 = n1184 ^ n508 ;
  assign n1186 = n171 & n1185 ;
  assign n1178 = n505 ^ n498 ;
  assign n1179 = x129 & n1178 ;
  assign n1180 = n1179 ^ n505 ;
  assign n1181 = n160 & n1180 ;
  assign n1187 = n1186 ^ n1181 ;
  assign n1188 = ~n1177 & ~n1187 ;
  assign n1189 = n214 & n1188 ;
  assign n1190 = n1189 ^ n214 ;
  assign n1149 = n443 ^ n429 ;
  assign n1150 = x129 & n1149 ;
  assign n1151 = n1150 ^ n1149 ;
  assign n1152 = n1151 ^ n443 ;
  assign n1153 = n148 & n1152 ;
  assign n1145 = n433 ^ n268 ;
  assign n1146 = x129 & n1145 ;
  assign n1147 = n1146 ^ n268 ;
  assign n1148 = n137 & n1147 ;
  assign n1154 = n1153 ^ n1148 ;
  assign n1159 = n464 ^ n440 ;
  assign n1160 = x129 & n1159 ;
  assign n1161 = n1160 ^ n1159 ;
  assign n1162 = n1161 ^ n464 ;
  assign n1163 = n171 & n1162 ;
  assign n1155 = n461 ^ n454 ;
  assign n1156 = x129 & n1155 ;
  assign n1157 = n1156 ^ n461 ;
  assign n1158 = n160 & n1157 ;
  assign n1164 = n1163 ^ n1158 ;
  assign n1165 = ~n1154 & ~n1164 ;
  assign n1166 = n136 & ~n1165 ;
  assign n1191 = n1190 ^ n1166 ;
  assign n1192 = ~n1144 & ~n1191 ;
  assign n1297 = n1296 ^ n1192 ;
  assign n1298 = x134 & n1297 ;
  assign n1299 = n1298 ^ n1297 ;
  assign n1300 = n1299 ^ n1296 ;
  assign n1549 = n965 ^ n847 ;
  assign n1550 = x129 & n1549 ;
  assign n1551 = n1550 ^ n1549 ;
  assign n1552 = n1551 ^ n965 ;
  assign n1553 = n974 ^ n852 ;
  assign n1554 = x129 & n1553 ;
  assign n1555 = n1554 ^ n1553 ;
  assign n1556 = n1555 ^ n974 ;
  assign n1557 = n1552 & ~n1556 ;
  assign n1558 = n1557 ^ n1556 ;
  assign n1540 = x47 ^ x46 ;
  assign n1541 = x128 & n1540 ;
  assign n1542 = n1541 ^ x47 ;
  assign n1543 = n1542 ^ n958 ;
  assign n1544 = x129 & ~n1543 ;
  assign n1545 = n1544 ^ x129 ;
  assign n1546 = n1545 ^ n1542 ;
  assign n1561 = n982 & n1546 ;
  assign n1562 = n1558 & n1561 ;
  assign n1559 = n137 & ~n1558 ;
  assign n1560 = n1559 ^ n137 ;
  assign n1563 = n1562 ^ n1560 ;
  assign n1547 = n148 & ~n1546 ;
  assign n1548 = n1547 ^ n148 ;
  assign n1564 = n1563 ^ n1548 ;
  assign n1575 = x43 & x128 ;
  assign n1576 = n1575 ^ x43 ;
  assign n1577 = n1576 ^ n204 ;
  assign n1578 = x129 & n1577 ;
  assign n1579 = n1578 ^ n1577 ;
  assign n1580 = n1579 ^ n204 ;
  assign n1582 = x41 & x128 ;
  assign n1583 = n1582 ^ x41 ;
  assign n1581 = x42 & x128 ;
  assign n1584 = n1583 ^ n1581 ;
  assign n1585 = x129 & n1584 ;
  assign n1586 = n1585 ^ n1584 ;
  assign n1587 = n1586 ^ n1583 ;
  assign n1588 = n1580 & ~n1587 ;
  assign n1589 = n1588 ^ n1587 ;
  assign n1590 = n171 & ~n1589 ;
  assign n1591 = n1590 ^ n171 ;
  assign n1565 = n196 ^ x39 ;
  assign n1566 = n1565 ^ n999 ;
  assign n1567 = x129 & n1566 ;
  assign n1568 = n1567 ^ n1565 ;
  assign n1569 = n1007 ^ n197 ;
  assign n1570 = x129 & n1569 ;
  assign n1571 = n1570 ^ n197 ;
  assign n1572 = n1568 & ~n1571 ;
  assign n1573 = n1572 ^ n1571 ;
  assign n1574 = n160 & n1573 ;
  assign n1592 = n1591 ^ n1574 ;
  assign n1593 = ~n1564 & ~n1592 ;
  assign n1594 = n214 & n1593 ;
  assign n1595 = n1594 ^ n214 ;
  assign n1503 = n827 ^ n813 ;
  assign n1504 = x129 & n1503 ;
  assign n1505 = n1504 ^ n1503 ;
  assign n1506 = n1505 ^ n827 ;
  assign n1507 = n836 ^ n818 ;
  assign n1508 = x129 & n1507 ;
  assign n1509 = n1508 ^ n1507 ;
  assign n1510 = n1509 ^ n836 ;
  assign n1511 = n1506 & ~n1510 ;
  assign n1512 = n1511 ^ n1510 ;
  assign n1513 = n148 & ~n1512 ;
  assign n1514 = n1513 ^ n148 ;
  assign n1492 = n811 ^ n562 ;
  assign n1493 = x129 & n1492 ;
  assign n1494 = n1493 ^ n1492 ;
  assign n1495 = n1494 ^ n811 ;
  assign n1496 = n820 ^ n567 ;
  assign n1497 = x129 & n1496 ;
  assign n1498 = n1497 ^ n1496 ;
  assign n1499 = n1498 ^ n820 ;
  assign n1500 = n1495 & ~n1499 ;
  assign n1501 = n1500 ^ n1499 ;
  assign n1502 = n137 & n1501 ;
  assign n1515 = n1514 ^ n1502 ;
  assign n1525 = n861 ^ n829 ;
  assign n1526 = x129 & n1525 ;
  assign n1527 = n1526 ^ n1525 ;
  assign n1528 = n1527 ^ n861 ;
  assign n1529 = n870 ^ n834 ;
  assign n1530 = x129 & n1529 ;
  assign n1531 = n1530 ^ n1529 ;
  assign n1532 = n1531 ^ n870 ;
  assign n1533 = n1528 & ~n1532 ;
  assign n1534 = n1533 ^ n1532 ;
  assign n1535 = n171 & ~n1534 ;
  assign n1536 = n1535 ^ n171 ;
  assign n1516 = n863 ^ n845 ;
  assign n1517 = x129 & n1516 ;
  assign n1518 = n1517 ^ n863 ;
  assign n1519 = n868 ^ n854 ;
  assign n1520 = x129 & n1519 ;
  assign n1521 = n1520 ^ n868 ;
  assign n1522 = n1518 & ~n1521 ;
  assign n1523 = n1522 ^ n1521 ;
  assign n1524 = n160 & n1523 ;
  assign n1537 = n1536 ^ n1524 ;
  assign n1538 = ~n1515 & ~n1537 ;
  assign n1539 = n136 & ~n1538 ;
  assign n1596 = n1595 ^ n1539 ;
  assign n1654 = n1038 ^ n1024 ;
  assign n1655 = x129 & n1654 ;
  assign n1656 = n1655 ^ n1654 ;
  assign n1657 = n1656 ^ n1038 ;
  assign n1658 = n1047 ^ n1029 ;
  assign n1659 = x129 & n1658 ;
  assign n1660 = n1659 ^ n1658 ;
  assign n1661 = n1660 ^ n1047 ;
  assign n1662 = n1657 & ~n1661 ;
  assign n1663 = n1662 ^ n1661 ;
  assign n1664 = n148 & ~n1663 ;
  assign n1665 = n1664 ^ n148 ;
  assign n1643 = n1022 ^ n1001 ;
  assign n1644 = x129 & n1643 ;
  assign n1645 = n1644 ^ n1643 ;
  assign n1646 = n1645 ^ n1022 ;
  assign n1647 = n1031 ^ n1006 ;
  assign n1648 = x129 & n1647 ;
  assign n1649 = n1648 ^ n1647 ;
  assign n1650 = n1649 ^ n1031 ;
  assign n1651 = n1646 & ~n1650 ;
  assign n1652 = n1651 ^ n1650 ;
  assign n1653 = n137 & n1652 ;
  assign n1666 = n1665 ^ n1653 ;
  assign n1676 = n1072 ^ n1040 ;
  assign n1677 = x129 & n1676 ;
  assign n1678 = n1677 ^ n1676 ;
  assign n1679 = n1678 ^ n1072 ;
  assign n1680 = n1081 ^ n1045 ;
  assign n1681 = x129 & n1680 ;
  assign n1682 = n1681 ^ n1680 ;
  assign n1683 = n1682 ^ n1081 ;
  assign n1684 = n1679 & ~n1683 ;
  assign n1685 = n1684 ^ n1683 ;
  assign n1686 = n171 & ~n1685 ;
  assign n1687 = n1686 ^ n171 ;
  assign n1667 = n1074 ^ n1056 ;
  assign n1668 = x129 & n1667 ;
  assign n1669 = n1668 ^ n1074 ;
  assign n1670 = n1079 ^ n1065 ;
  assign n1671 = x129 & n1670 ;
  assign n1672 = n1671 ^ n1079 ;
  assign n1673 = n1669 & ~n1672 ;
  assign n1674 = n1673 ^ n1672 ;
  assign n1675 = n160 & n1674 ;
  assign n1688 = n1687 ^ n1675 ;
  assign n1689 = ~n1666 & ~n1688 ;
  assign n1690 = n289 & n1689 ;
  assign n1691 = n1690 ^ n289 ;
  assign n1606 = n897 ^ n883 ;
  assign n1607 = x129 & n1606 ;
  assign n1608 = n1607 ^ n1606 ;
  assign n1609 = n1608 ^ n897 ;
  assign n1610 = n906 ^ n888 ;
  assign n1611 = x129 & n1610 ;
  assign n1612 = n1611 ^ n1610 ;
  assign n1613 = n1612 ^ n906 ;
  assign n1614 = n1609 & ~n1613 ;
  assign n1615 = n1614 ^ n1613 ;
  assign n1616 = n148 & ~n1615 ;
  assign n1617 = n1616 ^ n148 ;
  assign n1597 = n1058 ^ n881 ;
  assign n1598 = x129 & n1597 ;
  assign n1599 = n1598 ^ n1058 ;
  assign n1600 = n1063 ^ n890 ;
  assign n1601 = x129 & n1600 ;
  assign n1602 = n1601 ^ n1063 ;
  assign n1603 = n1599 & ~n1602 ;
  assign n1604 = n1603 ^ n1602 ;
  assign n1605 = n137 & n1604 ;
  assign n1618 = n1617 ^ n1605 ;
  assign n1628 = n931 ^ n899 ;
  assign n1629 = x129 & n1628 ;
  assign n1630 = n1629 ^ n1628 ;
  assign n1631 = n1630 ^ n931 ;
  assign n1632 = n940 ^ n904 ;
  assign n1633 = x129 & n1632 ;
  assign n1634 = n1633 ^ n1632 ;
  assign n1635 = n1634 ^ n940 ;
  assign n1636 = n1631 & ~n1635 ;
  assign n1637 = n1636 ^ n1635 ;
  assign n1638 = n171 & ~n1637 ;
  assign n1639 = n1638 ^ n171 ;
  assign n1619 = n933 ^ n915 ;
  assign n1620 = x129 & n1619 ;
  assign n1621 = n1620 ^ n933 ;
  assign n1622 = n938 ^ n924 ;
  assign n1623 = x129 & n1622 ;
  assign n1624 = n1623 ^ n938 ;
  assign n1625 = n1621 & ~n1624 ;
  assign n1626 = n1625 ^ n1624 ;
  assign n1627 = n160 & n1626 ;
  assign n1640 = n1639 ^ n1627 ;
  assign n1641 = ~n1618 & ~n1640 ;
  assign n1642 = n244 & ~n1641 ;
  assign n1692 = n1691 ^ n1642 ;
  assign n1693 = ~n1596 & ~n1692 ;
  assign n1358 = n612 ^ n598 ;
  assign n1359 = x129 & n1358 ;
  assign n1360 = n1359 ^ n1358 ;
  assign n1361 = n1360 ^ n612 ;
  assign n1362 = n621 ^ n603 ;
  assign n1363 = x129 & n1362 ;
  assign n1364 = n1363 ^ n1362 ;
  assign n1365 = n1364 ^ n621 ;
  assign n1366 = n1361 & ~n1365 ;
  assign n1367 = n1366 ^ n1365 ;
  assign n1368 = n148 & ~n1367 ;
  assign n1369 = n1368 ^ n148 ;
  assign n1349 = n774 ^ n596 ;
  assign n1350 = x129 & n1349 ;
  assign n1351 = n1350 ^ n774 ;
  assign n1352 = n779 ^ n605 ;
  assign n1353 = x129 & n1352 ;
  assign n1354 = n1353 ^ n779 ;
  assign n1355 = n1351 & ~n1354 ;
  assign n1356 = n1355 ^ n1354 ;
  assign n1357 = n137 & n1356 ;
  assign n1370 = n1369 ^ n1357 ;
  assign n1380 = n646 ^ n614 ;
  assign n1381 = x129 & n1380 ;
  assign n1382 = n1381 ^ n1380 ;
  assign n1383 = n1382 ^ n646 ;
  assign n1384 = n655 ^ n619 ;
  assign n1385 = x129 & n1384 ;
  assign n1386 = n1385 ^ n1384 ;
  assign n1387 = n1386 ^ n655 ;
  assign n1388 = n1383 & ~n1387 ;
  assign n1389 = n1388 ^ n1387 ;
  assign n1390 = n171 & ~n1389 ;
  assign n1391 = n1390 ^ n171 ;
  assign n1371 = n648 ^ n630 ;
  assign n1372 = x129 & n1371 ;
  assign n1373 = n1372 ^ n648 ;
  assign n1374 = n653 ^ n639 ;
  assign n1375 = x129 & n1374 ;
  assign n1376 = n1375 ^ n653 ;
  assign n1377 = n1373 & ~n1376 ;
  assign n1378 = n1377 ^ n1376 ;
  assign n1379 = n160 & n1378 ;
  assign n1392 = n1391 ^ n1379 ;
  assign n1393 = ~n1370 & ~n1392 ;
  assign n1394 = n289 & n1393 ;
  assign n1395 = n1394 ^ n289 ;
  assign n1312 = n754 ^ n740 ;
  assign n1313 = x129 & n1312 ;
  assign n1314 = n1313 ^ n1312 ;
  assign n1315 = n1314 ^ n754 ;
  assign n1316 = n763 ^ n745 ;
  assign n1317 = x129 & n1316 ;
  assign n1318 = n1317 ^ n1316 ;
  assign n1319 = n1318 ^ n763 ;
  assign n1320 = n1315 & ~n1319 ;
  assign n1321 = n1320 ^ n1319 ;
  assign n1322 = n148 & ~n1321 ;
  assign n1323 = n1322 ^ n148 ;
  assign n1301 = n738 ^ n704 ;
  assign n1302 = x129 & n1301 ;
  assign n1303 = n1302 ^ n1301 ;
  assign n1304 = n1303 ^ n738 ;
  assign n1305 = n747 ^ n709 ;
  assign n1306 = x129 & n1305 ;
  assign n1307 = n1306 ^ n1305 ;
  assign n1308 = n1307 ^ n747 ;
  assign n1309 = n1304 & ~n1308 ;
  assign n1310 = n1309 ^ n1308 ;
  assign n1311 = n137 & n1310 ;
  assign n1324 = n1323 ^ n1311 ;
  assign n1334 = n788 ^ n756 ;
  assign n1335 = x129 & n1334 ;
  assign n1336 = n1335 ^ n1334 ;
  assign n1337 = n1336 ^ n788 ;
  assign n1338 = n797 ^ n761 ;
  assign n1339 = x129 & n1338 ;
  assign n1340 = n1339 ^ n1338 ;
  assign n1341 = n1340 ^ n797 ;
  assign n1342 = n1337 & ~n1341 ;
  assign n1343 = n1342 ^ n1341 ;
  assign n1344 = n171 & ~n1343 ;
  assign n1345 = n1344 ^ n171 ;
  assign n1325 = n790 ^ n772 ;
  assign n1326 = x129 & n1325 ;
  assign n1327 = n1326 ^ n790 ;
  assign n1328 = n795 ^ n781 ;
  assign n1329 = x129 & n1328 ;
  assign n1330 = n1329 ^ n795 ;
  assign n1331 = n1327 & ~n1330 ;
  assign n1332 = n1331 ^ n1330 ;
  assign n1333 = n160 & n1332 ;
  assign n1346 = n1345 ^ n1333 ;
  assign n1347 = ~n1324 & ~n1346 ;
  assign n1348 = n214 & ~n1347 ;
  assign n1396 = n1395 ^ n1348 ;
  assign n1452 = n542 ^ n528 ;
  assign n1453 = x129 & n1452 ;
  assign n1454 = n1453 ^ n1452 ;
  assign n1455 = n1454 ^ n542 ;
  assign n1456 = n551 ^ n533 ;
  assign n1457 = x129 & n1456 ;
  assign n1458 = n1457 ^ n1456 ;
  assign n1459 = n1458 ^ n551 ;
  assign n1460 = n1455 & ~n1459 ;
  assign n1461 = n1460 ^ n1459 ;
  assign n1462 = n148 & ~n1461 ;
  assign n1463 = n1462 ^ n148 ;
  assign n1443 = n632 ^ n526 ;
  assign n1444 = x129 & n1443 ;
  assign n1445 = n1444 ^ n632 ;
  assign n1446 = n637 ^ n535 ;
  assign n1447 = x129 & n1446 ;
  assign n1448 = n1447 ^ n637 ;
  assign n1449 = n1445 & ~n1448 ;
  assign n1450 = n1449 ^ n1448 ;
  assign n1451 = n137 & n1450 ;
  assign n1464 = n1463 ^ n1451 ;
  assign n1474 = n576 ^ n544 ;
  assign n1475 = x129 & n1474 ;
  assign n1476 = n1475 ^ n1474 ;
  assign n1477 = n1476 ^ n576 ;
  assign n1478 = n585 ^ n549 ;
  assign n1479 = x129 & n1478 ;
  assign n1480 = n1479 ^ n1478 ;
  assign n1481 = n1480 ^ n585 ;
  assign n1482 = n1477 & ~n1481 ;
  assign n1483 = n1482 ^ n1481 ;
  assign n1484 = n171 & ~n1483 ;
  assign n1485 = n1484 ^ n171 ;
  assign n1465 = n578 ^ n560 ;
  assign n1466 = x129 & n1465 ;
  assign n1467 = n1466 ^ n578 ;
  assign n1468 = n583 ^ n569 ;
  assign n1469 = x129 & n1468 ;
  assign n1470 = n1469 ^ n583 ;
  assign n1471 = n1467 & ~n1470 ;
  assign n1472 = n1471 ^ n1470 ;
  assign n1473 = n160 & n1472 ;
  assign n1486 = n1485 ^ n1473 ;
  assign n1487 = ~n1464 & ~n1486 ;
  assign n1488 = n244 & n1487 ;
  assign n1489 = n1488 ^ n244 ;
  assign n1406 = n684 ^ n670 ;
  assign n1407 = x129 & n1406 ;
  assign n1408 = n1407 ^ n1406 ;
  assign n1409 = n1408 ^ n684 ;
  assign n1410 = n693 ^ n675 ;
  assign n1411 = x129 & n1410 ;
  assign n1412 = n1411 ^ n1410 ;
  assign n1413 = n1412 ^ n693 ;
  assign n1414 = n1409 & ~n1413 ;
  assign n1415 = n1414 ^ n1413 ;
  assign n1416 = n148 & ~n1415 ;
  assign n1417 = n1416 ^ n148 ;
  assign n1397 = n917 ^ n668 ;
  assign n1398 = x129 & n1397 ;
  assign n1399 = n1398 ^ n917 ;
  assign n1400 = n922 ^ n677 ;
  assign n1401 = x129 & n1400 ;
  assign n1402 = n1401 ^ n922 ;
  assign n1403 = n1399 & ~n1402 ;
  assign n1404 = n1403 ^ n1402 ;
  assign n1405 = n137 & n1404 ;
  assign n1418 = n1417 ^ n1405 ;
  assign n1428 = n718 ^ n686 ;
  assign n1429 = x129 & n1428 ;
  assign n1430 = n1429 ^ n1428 ;
  assign n1431 = n1430 ^ n718 ;
  assign n1432 = n727 ^ n691 ;
  assign n1433 = x129 & n1432 ;
  assign n1434 = n1433 ^ n1432 ;
  assign n1435 = n1434 ^ n727 ;
  assign n1436 = n1431 & ~n1435 ;
  assign n1437 = n1436 ^ n1435 ;
  assign n1438 = n171 & ~n1437 ;
  assign n1439 = n1438 ^ n171 ;
  assign n1419 = n720 ^ n702 ;
  assign n1420 = x129 & n1419 ;
  assign n1421 = n1420 ^ n720 ;
  assign n1422 = n725 ^ n711 ;
  assign n1423 = x129 & n1422 ;
  assign n1424 = n1423 ^ n725 ;
  assign n1425 = n1421 & ~n1424 ;
  assign n1426 = n1425 ^ n1424 ;
  assign n1427 = n160 & n1426 ;
  assign n1440 = n1439 ^ n1427 ;
  assign n1441 = ~n1418 & ~n1440 ;
  assign n1442 = n136 & ~n1441 ;
  assign n1490 = n1489 ^ n1442 ;
  assign n1491 = ~n1396 & ~n1490 ;
  assign n1694 = n1693 ^ n1491 ;
  assign n1695 = x134 & n1694 ;
  assign n1696 = n1695 ^ n1694 ;
  assign n1697 = n1696 ^ n1693 ;
  assign n1701 = n224 & n1015 ;
  assign n1702 = n210 & n1701 ;
  assign n1699 = n160 & ~n210 ;
  assign n1700 = n1699 ^ n160 ;
  assign n1703 = n1702 ^ n1700 ;
  assign n1698 = n171 & n224 ;
  assign n1704 = n1703 ^ n1698 ;
  assign n1706 = n169 & n226 ;
  assign n1707 = n1706 ^ n214 ;
  assign n1705 = n215 & n235 ;
  assign n1708 = n1707 ^ n1705 ;
  assign n1709 = ~n1704 & n1708 ;
  assign n1710 = n1709 ^ n214 ;
  assign n1712 = n146 & n148 ;
  assign n1711 = n137 & n366 ;
  assign n1713 = n1712 ^ n1711 ;
  assign n1715 = n157 & n171 ;
  assign n1714 = n160 & n180 ;
  assign n1716 = n1715 ^ n1714 ;
  assign n1717 = ~n1713 & ~n1716 ;
  assign n1718 = n136 & n1717 ;
  assign n1719 = n1718 ^ n136 ;
  assign n1720 = n1710 & n1719 ;
  assign n1721 = n1720 ^ n1710 ;
  assign n1722 = n1721 ^ n1719 ;
  assign n1732 = n137 & n319 ;
  assign n1731 = n148 & n253 ;
  assign n1733 = n1732 ^ n1731 ;
  assign n1735 = n171 & n263 ;
  assign n1734 = n160 & n284 ;
  assign n1736 = n1735 ^ n1734 ;
  assign n1737 = ~n1733 & ~n1736 ;
  assign n1738 = n244 & n1737 ;
  assign n1739 = n1738 ^ n244 ;
  assign n1724 = n148 & n298 ;
  assign n1723 = n137 & n194 ;
  assign n1725 = n1724 ^ n1723 ;
  assign n1727 = n171 & n308 ;
  assign n1726 = n160 & n329 ;
  assign n1728 = n1727 ^ n1726 ;
  assign n1729 = ~n1725 & ~n1728 ;
  assign n1730 = n289 & ~n1729 ;
  assign n1740 = n1739 ^ n1730 ;
  assign n1781 = x134 & ~n1740 ;
  assign n1782 = ~n1722 & n1781 ;
  assign n1751 = n148 & n389 ;
  assign n1750 = n137 & n501 ;
  assign n1752 = n1751 ^ n1750 ;
  assign n1754 = n171 & n399 ;
  assign n1753 = n160 & n420 ;
  assign n1755 = n1754 ^ n1753 ;
  assign n1756 = ~n1752 & ~n1755 ;
  assign n1757 = n289 & n1756 ;
  assign n1758 = n1757 ^ n289 ;
  assign n1743 = n148 & n345 ;
  assign n1742 = n137 & n410 ;
  assign n1744 = n1743 ^ n1742 ;
  assign n1746 = n171 & n355 ;
  assign n1745 = n160 & n376 ;
  assign n1747 = n1746 ^ n1745 ;
  assign n1748 = ~n1744 & ~n1747 ;
  assign n1749 = n244 & ~n1748 ;
  assign n1759 = n1758 ^ n1749 ;
  assign n1769 = n148 & n480 ;
  assign n1768 = n137 & n457 ;
  assign n1770 = n1769 ^ n1768 ;
  assign n1772 = n171 & n490 ;
  assign n1771 = n160 & n511 ;
  assign n1773 = n1772 ^ n1771 ;
  assign n1774 = ~n1770 & ~n1773 ;
  assign n1775 = n214 & n1774 ;
  assign n1776 = n1775 ^ n214 ;
  assign n1761 = n148 & n436 ;
  assign n1760 = n137 & n274 ;
  assign n1762 = n1761 ^ n1760 ;
  assign n1764 = n171 & n446 ;
  assign n1763 = n160 & n467 ;
  assign n1765 = n1764 ^ n1763 ;
  assign n1766 = ~n1762 & ~n1765 ;
  assign n1767 = n136 & ~n1766 ;
  assign n1777 = n1776 ^ n1767 ;
  assign n1778 = ~n1759 & ~n1777 ;
  assign n1780 = x134 & n1778 ;
  assign n1783 = n1782 ^ n1780 ;
  assign n1741 = ~n1722 & ~n1740 ;
  assign n1779 = n1778 ^ n1741 ;
  assign n1784 = n1783 ^ n1779 ;
  assign n1785 = n1784 ^ n1741 ;
  assign n1793 = n160 & ~n996 ;
  assign n1794 = n1793 ^ n160 ;
  assign n1795 = n171 & ~n962 ;
  assign n1796 = n1795 ^ n171 ;
  assign n1797 = n1794 & n1796 ;
  assign n1798 = n1797 ^ n1794 ;
  assign n1799 = n1798 ^ n1796 ;
  assign n1786 = n137 & ~n859 ;
  assign n1787 = n1786 ^ n137 ;
  assign n1788 = n148 & ~n979 ;
  assign n1789 = n1788 ^ n148 ;
  assign n1790 = n1787 & n1789 ;
  assign n1791 = n1790 ^ n1787 ;
  assign n1792 = n1791 ^ n1789 ;
  assign n1800 = n1799 ^ n1792 ;
  assign n1801 = n1799 ^ n214 ;
  assign n1802 = ~n214 & n1801 ;
  assign n1803 = n1802 ^ n214 ;
  assign n1804 = n1803 ^ n1792 ;
  assign n1805 = n1800 & n1804 ;
  assign n1806 = n1805 ^ n1802 ;
  assign n1807 = n1806 ^ n1792 ;
  assign n1809 = n148 & ~n825 ;
  assign n1810 = n1809 ^ n148 ;
  assign n1808 = n137 & n574 ;
  assign n1811 = n1810 ^ n1808 ;
  assign n1813 = n171 & ~n841 ;
  assign n1814 = n1813 ^ n171 ;
  assign n1812 = n160 & n875 ;
  assign n1815 = n1814 ^ n1812 ;
  assign n1816 = ~n1811 & ~n1815 ;
  assign n1817 = n136 & n1816 ;
  assign n1818 = n1817 ^ n136 ;
  assign n1819 = n1807 & n1818 ;
  assign n1820 = n1819 ^ n1807 ;
  assign n1821 = n1820 ^ n1818 ;
  assign n1833 = n148 & ~n895 ;
  assign n1834 = n1833 ^ n148 ;
  assign n1832 = n137 & n1070 ;
  assign n1835 = n1834 ^ n1832 ;
  assign n1837 = n171 & ~n911 ;
  assign n1838 = n1837 ^ n171 ;
  assign n1836 = n160 & n945 ;
  assign n1839 = n1838 ^ n1836 ;
  assign n1840 = ~n1835 & ~n1839 ;
  assign n1841 = n244 & n1840 ;
  assign n1842 = n1841 ^ n244 ;
  assign n1823 = n148 & ~n1036 ;
  assign n1824 = n1823 ^ n148 ;
  assign n1822 = n137 & n1012 ;
  assign n1825 = n1824 ^ n1822 ;
  assign n1827 = n171 & ~n1052 ;
  assign n1828 = n1827 ^ n171 ;
  assign n1826 = n160 & n1086 ;
  assign n1829 = n1828 ^ n1826 ;
  assign n1830 = ~n1825 & ~n1829 ;
  assign n1831 = n289 & ~n1830 ;
  assign n1843 = n1842 ^ n1831 ;
  assign n1892 = x134 & ~n1843 ;
  assign n1893 = ~n1821 & n1892 ;
  assign n1856 = n148 & ~n610 ;
  assign n1857 = n1856 ^ n148 ;
  assign n1855 = n137 & n786 ;
  assign n1858 = n1857 ^ n1855 ;
  assign n1860 = n171 & ~n626 ;
  assign n1861 = n1860 ^ n171 ;
  assign n1859 = n160 & n660 ;
  assign n1862 = n1861 ^ n1859 ;
  assign n1863 = ~n1858 & ~n1862 ;
  assign n1864 = n289 & n1863 ;
  assign n1865 = n1864 ^ n289 ;
  assign n1846 = n148 & ~n540 ;
  assign n1847 = n1846 ^ n148 ;
  assign n1845 = n137 & n644 ;
  assign n1848 = n1847 ^ n1845 ;
  assign n1850 = n171 & ~n556 ;
  assign n1851 = n1850 ^ n171 ;
  assign n1849 = n160 & n590 ;
  assign n1852 = n1851 ^ n1849 ;
  assign n1853 = ~n1848 & ~n1852 ;
  assign n1854 = n244 & ~n1853 ;
  assign n1866 = n1865 ^ n1854 ;
  assign n1878 = n148 & ~n752 ;
  assign n1879 = n1878 ^ n148 ;
  assign n1877 = n137 & n716 ;
  assign n1880 = n1879 ^ n1877 ;
  assign n1882 = n171 & ~n768 ;
  assign n1883 = n1882 ^ n171 ;
  assign n1881 = n160 & n802 ;
  assign n1884 = n1883 ^ n1881 ;
  assign n1885 = ~n1880 & ~n1884 ;
  assign n1886 = n214 & n1885 ;
  assign n1887 = n1886 ^ n214 ;
  assign n1868 = n148 & ~n682 ;
  assign n1869 = n1868 ^ n148 ;
  assign n1867 = n137 & n929 ;
  assign n1870 = n1869 ^ n1867 ;
  assign n1872 = n171 & ~n698 ;
  assign n1873 = n1872 ^ n171 ;
  assign n1871 = n160 & n732 ;
  assign n1874 = n1873 ^ n1871 ;
  assign n1875 = ~n1870 & ~n1874 ;
  assign n1876 = n136 & ~n1875 ;
  assign n1888 = n1887 ^ n1876 ;
  assign n1889 = ~n1866 & ~n1888 ;
  assign n1891 = x134 & n1889 ;
  assign n1894 = n1893 ^ n1891 ;
  assign n1844 = ~n1821 & ~n1843 ;
  assign n1890 = n1889 ^ n1844 ;
  assign n1895 = n1894 ^ n1890 ;
  assign n1896 = n1895 ^ n1844 ;
  assign n1943 = n148 & n1196 ;
  assign n1942 = n137 & n1111 ;
  assign n1944 = n1943 ^ n1942 ;
  assign n1946 = n171 & n1201 ;
  assign n1945 = n160 & n1211 ;
  assign n1947 = n1946 ^ n1945 ;
  assign n1948 = ~n1944 & ~n1947 ;
  assign n1949 = n136 & n1948 ;
  assign n1950 = n1949 ^ n136 ;
  assign n1935 = n148 & n1243 ;
  assign n1934 = n137 & n1206 ;
  assign n1936 = n1935 ^ n1934 ;
  assign n1938 = n171 & n1248 ;
  assign n1937 = n160 & n1266 ;
  assign n1939 = n1938 ^ n1937 ;
  assign n1940 = ~n1936 & ~n1939 ;
  assign n1941 = n214 & ~n1940 ;
  assign n1951 = n1950 ^ n1941 ;
  assign n1961 = n148 & n1218 ;
  assign n1960 = n137 & n1284 ;
  assign n1962 = n1961 ^ n1960 ;
  assign n1964 = n171 & n1223 ;
  assign n1963 = n160 & n1233 ;
  assign n1965 = n1964 ^ n1963 ;
  assign n1966 = ~n1962 & ~n1965 ;
  assign n1967 = n244 & n1966 ;
  assign n1968 = n1967 ^ n244 ;
  assign n1953 = n148 & n1274 ;
  assign n1952 = n137 & n1257 ;
  assign n1954 = n1953 ^ n1952 ;
  assign n1956 = n171 & n1279 ;
  assign n1955 = n160 & n1289 ;
  assign n1957 = n1956 ^ n1955 ;
  assign n1958 = ~n1954 & ~n1957 ;
  assign n1959 = n289 & ~n1958 ;
  assign n1969 = n1968 ^ n1959 ;
  assign n1970 = ~n1951 & ~n1969 ;
  assign n1906 = n148 & n1123 ;
  assign n1905 = n137 & n1180 ;
  assign n1907 = n1906 ^ n1905 ;
  assign n1909 = n171 & n1128 ;
  assign n1908 = n160 & n1138 ;
  assign n1910 = n1909 ^ n1908 ;
  assign n1911 = ~n1907 & ~n1910 ;
  assign n1912 = n289 & n1911 ;
  assign n1913 = n1912 ^ n289 ;
  assign n1898 = n148 & n1101 ;
  assign n1897 = n137 & n1133 ;
  assign n1899 = n1898 ^ n1897 ;
  assign n1901 = n171 & n1106 ;
  assign n1900 = n160 & n1116 ;
  assign n1902 = n1901 ^ n1900 ;
  assign n1903 = ~n1899 & ~n1902 ;
  assign n1904 = n244 & ~n1903 ;
  assign n1914 = n1913 ^ n1904 ;
  assign n1924 = n148 & n1170 ;
  assign n1923 = n137 & n1157 ;
  assign n1925 = n1924 ^ n1923 ;
  assign n1927 = n171 & n1175 ;
  assign n1926 = n160 & n1185 ;
  assign n1928 = n1927 ^ n1926 ;
  assign n1929 = ~n1925 & ~n1928 ;
  assign n1930 = n214 & n1929 ;
  assign n1931 = n1930 ^ n214 ;
  assign n1916 = n148 & n1147 ;
  assign n1915 = n137 & n1228 ;
  assign n1917 = n1916 ^ n1915 ;
  assign n1919 = n171 & n1152 ;
  assign n1918 = n160 & n1162 ;
  assign n1920 = n1919 ^ n1918 ;
  assign n1921 = ~n1917 & ~n1920 ;
  assign n1922 = n136 & ~n1921 ;
  assign n1932 = n1931 ^ n1922 ;
  assign n1933 = ~n1914 & ~n1932 ;
  assign n1971 = n1970 ^ n1933 ;
  assign n1972 = x134 & n1971 ;
  assign n1973 = n1972 ^ n1971 ;
  assign n1974 = n1973 ^ n1970 ;
  assign n2036 = n148 & ~n1501 ;
  assign n2037 = n2036 ^ n148 ;
  assign n2035 = n137 & n1472 ;
  assign n2038 = n2037 ^ n2035 ;
  assign n2040 = n171 & ~n1512 ;
  assign n2041 = n2040 ^ n171 ;
  assign n2039 = n160 & n1534 ;
  assign n2042 = n2041 ^ n2039 ;
  assign n2043 = ~n2038 & ~n2042 ;
  assign n2044 = n136 & n2043 ;
  assign n2045 = n2044 ^ n136 ;
  assign n2024 = n148 & n171 ;
  assign n2025 = n1546 & n2024 ;
  assign n2026 = n1558 & n2025 ;
  assign n2022 = n148 & ~n1558 ;
  assign n2023 = n2022 ^ n148 ;
  assign n2027 = n2026 ^ n2023 ;
  assign n2020 = n171 & ~n1546 ;
  assign n2021 = n2020 ^ n171 ;
  assign n2028 = n2027 ^ n2021 ;
  assign n2030 = n137 & ~n1523 ;
  assign n2031 = n2030 ^ n137 ;
  assign n2029 = n160 & n1589 ;
  assign n2032 = n2031 ^ n2029 ;
  assign n2033 = ~n2028 & ~n2032 ;
  assign n2034 = n214 & ~n2033 ;
  assign n2046 = n2045 ^ n2034 ;
  assign n2058 = n148 & ~n1604 ;
  assign n2059 = n2058 ^ n148 ;
  assign n2057 = n137 & n1674 ;
  assign n2060 = n2059 ^ n2057 ;
  assign n2062 = n171 & ~n1615 ;
  assign n2063 = n2062 ^ n171 ;
  assign n2061 = n160 & n1637 ;
  assign n2064 = n2063 ^ n2061 ;
  assign n2065 = ~n2060 & ~n2064 ;
  assign n2066 = n244 & n2065 ;
  assign n2067 = n2066 ^ n244 ;
  assign n2048 = n148 & ~n1652 ;
  assign n2049 = n2048 ^ n148 ;
  assign n2047 = n137 & n1573 ;
  assign n2050 = n2049 ^ n2047 ;
  assign n2052 = n171 & ~n1663 ;
  assign n2053 = n2052 ^ n171 ;
  assign n2051 = n160 & n1685 ;
  assign n2054 = n2053 ^ n2051 ;
  assign n2055 = ~n2050 & ~n2054 ;
  assign n2056 = n289 & ~n2055 ;
  assign n2068 = n2067 ^ n2056 ;
  assign n2069 = ~n2046 & ~n2068 ;
  assign n1986 = n148 & ~n1356 ;
  assign n1987 = n1986 ^ n148 ;
  assign n1985 = n137 & n1332 ;
  assign n1988 = n1987 ^ n1985 ;
  assign n1990 = n171 & ~n1367 ;
  assign n1991 = n1990 ^ n171 ;
  assign n1989 = n160 & n1389 ;
  assign n1992 = n1991 ^ n1989 ;
  assign n1993 = ~n1988 & ~n1992 ;
  assign n1994 = n289 & n1993 ;
  assign n1995 = n1994 ^ n289 ;
  assign n1976 = n148 & ~n1450 ;
  assign n1977 = n1976 ^ n148 ;
  assign n1975 = n137 & n1378 ;
  assign n1978 = n1977 ^ n1975 ;
  assign n1980 = n171 & ~n1461 ;
  assign n1981 = n1980 ^ n171 ;
  assign n1979 = n160 & n1483 ;
  assign n1982 = n1981 ^ n1979 ;
  assign n1983 = ~n1978 & ~n1982 ;
  assign n1984 = n244 & ~n1983 ;
  assign n1996 = n1995 ^ n1984 ;
  assign n2008 = n148 & ~n1310 ;
  assign n2009 = n2008 ^ n148 ;
  assign n2007 = n137 & n1426 ;
  assign n2010 = n2009 ^ n2007 ;
  assign n2012 = n171 & ~n1321 ;
  assign n2013 = n2012 ^ n171 ;
  assign n2011 = n160 & n1343 ;
  assign n2014 = n2013 ^ n2011 ;
  assign n2015 = ~n2010 & ~n2014 ;
  assign n2016 = n214 & n2015 ;
  assign n2017 = n2016 ^ n214 ;
  assign n1998 = n148 & ~n1404 ;
  assign n1999 = n1998 ^ n148 ;
  assign n1997 = n137 & n1626 ;
  assign n2000 = n1999 ^ n1997 ;
  assign n2002 = n171 & ~n1415 ;
  assign n2003 = n2002 ^ n171 ;
  assign n2001 = n160 & n1437 ;
  assign n2004 = n2003 ^ n2001 ;
  assign n2005 = ~n2000 & ~n2004 ;
  assign n2006 = n136 & ~n2005 ;
  assign n2018 = n2017 ^ n2006 ;
  assign n2019 = ~n1996 & ~n2018 ;
  assign n2070 = n2069 ^ n2019 ;
  assign n2071 = x134 & n2070 ;
  assign n2072 = n2071 ^ n2070 ;
  assign n2073 = n2072 ^ n2069 ;
  assign n2082 = n171 & n298 ;
  assign n2081 = n160 & n308 ;
  assign n2083 = n2082 ^ n2081 ;
  assign n2077 = n194 & n982 ;
  assign n2078 = n210 & n2077 ;
  assign n2075 = n137 & ~n210 ;
  assign n2076 = n2075 ^ n137 ;
  assign n2079 = n2078 ^ n2076 ;
  assign n2074 = n148 & n194 ;
  assign n2080 = n2079 ^ n2074 ;
  assign n2084 = n2083 ^ n2080 ;
  assign n2087 = n160 & ~n289 ;
  assign n2088 = n308 & n2087 ;
  assign n2085 = n171 & ~n289 ;
  assign n2086 = n298 & n2085 ;
  assign n2089 = n2088 ^ n2086 ;
  assign n2090 = n2089 ^ n289 ;
  assign n2091 = n2090 ^ n2080 ;
  assign n2092 = n2084 & n2091 ;
  assign n2093 = n2092 ^ n2089 ;
  assign n2094 = n2093 ^ n2080 ;
  assign n2096 = n137 & n329 ;
  assign n2095 = n148 & n319 ;
  assign n2097 = n2096 ^ n2095 ;
  assign n2099 = n171 & n253 ;
  assign n2098 = n160 & n263 ;
  assign n2100 = n2099 ^ n2098 ;
  assign n2101 = ~n2097 & ~n2100 ;
  assign n2102 = n244 & n2101 ;
  assign n2103 = n2102 ^ n244 ;
  assign n2104 = n2094 & n2103 ;
  assign n2105 = n2104 ^ n2094 ;
  assign n2106 = n2105 ^ n2103 ;
  assign n2116 = n148 & n366 ;
  assign n2115 = n137 & n376 ;
  assign n2117 = n2116 ^ n2115 ;
  assign n2119 = n146 & n171 ;
  assign n2118 = n157 & n160 ;
  assign n2120 = n2119 ^ n2118 ;
  assign n2121 = ~n2117 & ~n2120 ;
  assign n2122 = n136 & n2121 ;
  assign n2123 = n2122 ^ n136 ;
  assign n2108 = n148 & n169 ;
  assign n2107 = n137 & n180 ;
  assign n2109 = n2108 ^ n2107 ;
  assign n2111 = n171 & n235 ;
  assign n2110 = n160 & n224 ;
  assign n2112 = n2111 ^ n2110 ;
  assign n2113 = ~n2109 & ~n2112 ;
  assign n2114 = n214 & ~n2113 ;
  assign n2124 = n2123 ^ n2114 ;
  assign n2165 = x134 & ~n2124 ;
  assign n2166 = ~n2106 & n2165 ;
  assign n2135 = n148 & n501 ;
  assign n2134 = n137 & n511 ;
  assign n2136 = n2135 ^ n2134 ;
  assign n2138 = n171 & n389 ;
  assign n2137 = n160 & n399 ;
  assign n2139 = n2138 ^ n2137 ;
  assign n2140 = ~n2136 & ~n2139 ;
  assign n2141 = n289 & n2140 ;
  assign n2142 = n2141 ^ n289 ;
  assign n2127 = n148 & n410 ;
  assign n2126 = n137 & n420 ;
  assign n2128 = n2127 ^ n2126 ;
  assign n2130 = n171 & n345 ;
  assign n2129 = n160 & n355 ;
  assign n2131 = n2130 ^ n2129 ;
  assign n2132 = ~n2128 & ~n2131 ;
  assign n2133 = n244 & ~n2132 ;
  assign n2143 = n2142 ^ n2133 ;
  assign n2153 = n148 & n457 ;
  assign n2152 = n137 & n467 ;
  assign n2154 = n2153 ^ n2152 ;
  assign n2156 = n171 & n480 ;
  assign n2155 = n160 & n490 ;
  assign n2157 = n2156 ^ n2155 ;
  assign n2158 = ~n2154 & ~n2157 ;
  assign n2159 = n214 & n2158 ;
  assign n2160 = n2159 ^ n214 ;
  assign n2145 = n148 & n274 ;
  assign n2144 = n137 & n284 ;
  assign n2146 = n2145 ^ n2144 ;
  assign n2148 = n171 & n436 ;
  assign n2147 = n160 & n446 ;
  assign n2149 = n2148 ^ n2147 ;
  assign n2150 = ~n2146 & ~n2149 ;
  assign n2151 = n136 & ~n2150 ;
  assign n2161 = n2160 ^ n2151 ;
  assign n2162 = ~n2143 & ~n2161 ;
  assign n2164 = x134 & n2162 ;
  assign n2167 = n2166 ^ n2164 ;
  assign n2125 = ~n2106 & ~n2124 ;
  assign n2163 = n2162 ^ n2125 ;
  assign n2168 = n2167 ^ n2163 ;
  assign n2169 = n2168 ^ n2125 ;
  assign n2226 = n148 & ~n574 ;
  assign n2227 = n2226 ^ n148 ;
  assign n2225 = n137 & n590 ;
  assign n2228 = n2227 ^ n2225 ;
  assign n2230 = n171 & ~n825 ;
  assign n2231 = n2230 ^ n171 ;
  assign n2229 = n160 & n841 ;
  assign n2232 = n2231 ^ n2229 ;
  assign n2233 = ~n2228 & ~n2232 ;
  assign n2234 = n136 & n2233 ;
  assign n2235 = n2234 ^ n136 ;
  assign n2216 = n148 & ~n859 ;
  assign n2217 = n2216 ^ n148 ;
  assign n2215 = n137 & n875 ;
  assign n2218 = n2217 ^ n2215 ;
  assign n2221 = n160 & n962 ;
  assign n2219 = n171 & ~n979 ;
  assign n2220 = n2219 ^ n171 ;
  assign n2222 = n2221 ^ n2220 ;
  assign n2223 = ~n2218 & ~n2222 ;
  assign n2224 = n214 & ~n2223 ;
  assign n2236 = n2235 ^ n2224 ;
  assign n2248 = n148 & ~n1070 ;
  assign n2249 = n2248 ^ n148 ;
  assign n2247 = n137 & n1086 ;
  assign n2250 = n2249 ^ n2247 ;
  assign n2252 = n171 & ~n895 ;
  assign n2253 = n2252 ^ n171 ;
  assign n2251 = n160 & n911 ;
  assign n2254 = n2253 ^ n2251 ;
  assign n2255 = ~n2250 & ~n2254 ;
  assign n2256 = n244 & n2255 ;
  assign n2257 = n2256 ^ n244 ;
  assign n2239 = n137 & n996 ;
  assign n2237 = n148 & ~n1012 ;
  assign n2238 = n2237 ^ n148 ;
  assign n2240 = n2239 ^ n2238 ;
  assign n2242 = n171 & ~n1036 ;
  assign n2243 = n2242 ^ n171 ;
  assign n2241 = n160 & n1052 ;
  assign n2244 = n2243 ^ n2241 ;
  assign n2245 = ~n2240 & ~n2244 ;
  assign n2246 = n289 & ~n2245 ;
  assign n2258 = n2257 ^ n2246 ;
  assign n2259 = ~n2236 & ~n2258 ;
  assign n2181 = n148 & ~n786 ;
  assign n2182 = n2181 ^ n148 ;
  assign n2180 = n137 & n802 ;
  assign n2183 = n2182 ^ n2180 ;
  assign n2185 = n171 & ~n610 ;
  assign n2186 = n2185 ^ n171 ;
  assign n2184 = n160 & n626 ;
  assign n2187 = n2186 ^ n2184 ;
  assign n2188 = ~n2183 & ~n2187 ;
  assign n2189 = n289 & n2188 ;
  assign n2190 = n2189 ^ n289 ;
  assign n2171 = n148 & ~n644 ;
  assign n2172 = n2171 ^ n148 ;
  assign n2170 = n137 & n660 ;
  assign n2173 = n2172 ^ n2170 ;
  assign n2175 = n171 & ~n540 ;
  assign n2176 = n2175 ^ n171 ;
  assign n2174 = n160 & n556 ;
  assign n2177 = n2176 ^ n2174 ;
  assign n2178 = ~n2173 & ~n2177 ;
  assign n2179 = n244 & ~n2178 ;
  assign n2191 = n2190 ^ n2179 ;
  assign n2203 = n148 & ~n716 ;
  assign n2204 = n2203 ^ n148 ;
  assign n2202 = n137 & n732 ;
  assign n2205 = n2204 ^ n2202 ;
  assign n2207 = n171 & ~n752 ;
  assign n2208 = n2207 ^ n171 ;
  assign n2206 = n160 & n768 ;
  assign n2209 = n2208 ^ n2206 ;
  assign n2210 = ~n2205 & ~n2209 ;
  assign n2211 = n214 & n2210 ;
  assign n2212 = n2211 ^ n214 ;
  assign n2193 = n148 & ~n929 ;
  assign n2194 = n2193 ^ n148 ;
  assign n2192 = n137 & n945 ;
  assign n2195 = n2194 ^ n2192 ;
  assign n2197 = n171 & ~n682 ;
  assign n2198 = n2197 ^ n171 ;
  assign n2196 = n160 & n698 ;
  assign n2199 = n2198 ^ n2196 ;
  assign n2200 = ~n2195 & ~n2199 ;
  assign n2201 = n136 & ~n2200 ;
  assign n2213 = n2212 ^ n2201 ;
  assign n2214 = ~n2191 & ~n2213 ;
  assign n2260 = n2259 ^ n2214 ;
  assign n2261 = x134 & n2260 ;
  assign n2262 = n2261 ^ n2260 ;
  assign n2263 = n2262 ^ n2259 ;
  assign n2310 = n148 & n1111 ;
  assign n2309 = n137 & n1116 ;
  assign n2311 = n2310 ^ n2309 ;
  assign n2313 = n171 & n1196 ;
  assign n2312 = n160 & n1201 ;
  assign n2314 = n2313 ^ n2312 ;
  assign n2315 = ~n2311 & ~n2314 ;
  assign n2316 = n136 & n2315 ;
  assign n2317 = n2316 ^ n136 ;
  assign n2302 = n148 & n1206 ;
  assign n2301 = n137 & n1211 ;
  assign n2303 = n2302 ^ n2301 ;
  assign n2305 = n171 & n1243 ;
  assign n2304 = n160 & n1248 ;
  assign n2306 = n2305 ^ n2304 ;
  assign n2307 = ~n2303 & ~n2306 ;
  assign n2308 = n214 & ~n2307 ;
  assign n2318 = n2317 ^ n2308 ;
  assign n2329 = n148 & n1284 ;
  assign n2328 = n137 & n1289 ;
  assign n2330 = n2329 ^ n2328 ;
  assign n2332 = n171 & n1218 ;
  assign n2331 = n160 & n1223 ;
  assign n2333 = n2332 ^ n2331 ;
  assign n2334 = ~n2330 & ~n2333 ;
  assign n2335 = n244 & n2334 ;
  assign n2336 = n2335 ^ n244 ;
  assign n2320 = n148 & ~n1257 ;
  assign n2321 = n2320 ^ n148 ;
  assign n2319 = n137 & n1266 ;
  assign n2322 = n2321 ^ n2319 ;
  assign n2324 = n171 & n1274 ;
  assign n2323 = n160 & n1279 ;
  assign n2325 = n2324 ^ n2323 ;
  assign n2326 = ~n2322 & ~n2325 ;
  assign n2327 = n289 & ~n2326 ;
  assign n2337 = n2336 ^ n2327 ;
  assign n2338 = ~n2318 & ~n2337 ;
  assign n2273 = n148 & n1180 ;
  assign n2272 = n137 & n1185 ;
  assign n2274 = n2273 ^ n2272 ;
  assign n2276 = n171 & n1123 ;
  assign n2275 = n160 & n1128 ;
  assign n2277 = n2276 ^ n2275 ;
  assign n2278 = ~n2274 & ~n2277 ;
  assign n2279 = n289 & n2278 ;
  assign n2280 = n2279 ^ n289 ;
  assign n2265 = n148 & n1133 ;
  assign n2264 = n137 & n1138 ;
  assign n2266 = n2265 ^ n2264 ;
  assign n2268 = n171 & n1101 ;
  assign n2267 = n160 & n1106 ;
  assign n2269 = n2268 ^ n2267 ;
  assign n2270 = ~n2266 & ~n2269 ;
  assign n2271 = n244 & ~n2270 ;
  assign n2281 = n2280 ^ n2271 ;
  assign n2291 = n148 & n1157 ;
  assign n2290 = n137 & n1162 ;
  assign n2292 = n2291 ^ n2290 ;
  assign n2294 = n171 & n1170 ;
  assign n2293 = n160 & n1175 ;
  assign n2295 = n2294 ^ n2293 ;
  assign n2296 = ~n2292 & ~n2295 ;
  assign n2297 = n214 & n2296 ;
  assign n2298 = n2297 ^ n214 ;
  assign n2283 = n148 & n1228 ;
  assign n2282 = n137 & n1233 ;
  assign n2284 = n2283 ^ n2282 ;
  assign n2286 = n171 & n1147 ;
  assign n2285 = n160 & n1152 ;
  assign n2287 = n2286 ^ n2285 ;
  assign n2288 = ~n2284 & ~n2287 ;
  assign n2289 = n136 & ~n2288 ;
  assign n2299 = n2298 ^ n2289 ;
  assign n2300 = ~n2281 & ~n2299 ;
  assign n2339 = n2338 ^ n2300 ;
  assign n2340 = x134 & n2339 ;
  assign n2341 = n2340 ^ n2339 ;
  assign n2342 = n2341 ^ n2338 ;
  assign n2399 = n148 & ~n1472 ;
  assign n2400 = n2399 ^ n148 ;
  assign n2398 = n137 & n1483 ;
  assign n2401 = n2400 ^ n2398 ;
  assign n2403 = n171 & ~n1501 ;
  assign n2404 = n2403 ^ n171 ;
  assign n2402 = n160 & n1512 ;
  assign n2405 = n2404 ^ n2402 ;
  assign n2406 = ~n2401 & ~n2405 ;
  assign n2407 = n136 & n2406 ;
  assign n2408 = n2407 ^ n136 ;
  assign n2389 = n171 & ~n1558 ;
  assign n2390 = n2389 ^ n171 ;
  assign n2388 = n137 & n1534 ;
  assign n2391 = n2390 ^ n2388 ;
  assign n2394 = n160 & n1546 ;
  assign n2392 = n148 & ~n1523 ;
  assign n2393 = n2392 ^ n148 ;
  assign n2395 = n2394 ^ n2393 ;
  assign n2396 = ~n2391 & ~n2395 ;
  assign n2397 = n214 & ~n2396 ;
  assign n2409 = n2408 ^ n2397 ;
  assign n2421 = n148 & ~n1674 ;
  assign n2422 = n2421 ^ n148 ;
  assign n2420 = n137 & n1685 ;
  assign n2423 = n2422 ^ n2420 ;
  assign n2425 = n171 & ~n1604 ;
  assign n2426 = n2425 ^ n171 ;
  assign n2424 = n160 & n1615 ;
  assign n2427 = n2426 ^ n2424 ;
  assign n2428 = ~n2423 & ~n2427 ;
  assign n2429 = n244 & n2428 ;
  assign n2430 = n2429 ^ n244 ;
  assign n2411 = n148 & ~n1573 ;
  assign n2412 = n2411 ^ n148 ;
  assign n2410 = n137 & n1589 ;
  assign n2413 = n2412 ^ n2410 ;
  assign n2415 = n171 & ~n1652 ;
  assign n2416 = n2415 ^ n171 ;
  assign n2414 = n160 & n1663 ;
  assign n2417 = n2416 ^ n2414 ;
  assign n2418 = ~n2413 & ~n2417 ;
  assign n2419 = n289 & ~n2418 ;
  assign n2431 = n2430 ^ n2419 ;
  assign n2432 = ~n2409 & ~n2431 ;
  assign n2354 = n148 & ~n1332 ;
  assign n2355 = n2354 ^ n148 ;
  assign n2353 = n137 & n1343 ;
  assign n2356 = n2355 ^ n2353 ;
  assign n2358 = n171 & ~n1356 ;
  assign n2359 = n2358 ^ n171 ;
  assign n2357 = n160 & n1367 ;
  assign n2360 = n2359 ^ n2357 ;
  assign n2361 = ~n2356 & ~n2360 ;
  assign n2362 = n289 & n2361 ;
  assign n2363 = n2362 ^ n289 ;
  assign n2344 = n148 & ~n1378 ;
  assign n2345 = n2344 ^ n148 ;
  assign n2343 = n137 & n1389 ;
  assign n2346 = n2345 ^ n2343 ;
  assign n2348 = n171 & ~n1450 ;
  assign n2349 = n2348 ^ n171 ;
  assign n2347 = n160 & n1461 ;
  assign n2350 = n2349 ^ n2347 ;
  assign n2351 = ~n2346 & ~n2350 ;
  assign n2352 = n244 & ~n2351 ;
  assign n2364 = n2363 ^ n2352 ;
  assign n2376 = n148 & ~n1426 ;
  assign n2377 = n2376 ^ n148 ;
  assign n2375 = n137 & n1437 ;
  assign n2378 = n2377 ^ n2375 ;
  assign n2380 = n171 & ~n1310 ;
  assign n2381 = n2380 ^ n171 ;
  assign n2379 = n160 & n1321 ;
  assign n2382 = n2381 ^ n2379 ;
  assign n2383 = ~n2378 & ~n2382 ;
  assign n2384 = n214 & n2383 ;
  assign n2385 = n2384 ^ n214 ;
  assign n2366 = n148 & ~n1626 ;
  assign n2367 = n2366 ^ n148 ;
  assign n2365 = n137 & n1637 ;
  assign n2368 = n2367 ^ n2365 ;
  assign n2370 = n171 & ~n1404 ;
  assign n2371 = n2370 ^ n171 ;
  assign n2369 = n160 & n1415 ;
  assign n2372 = n2371 ^ n2369 ;
  assign n2373 = ~n2368 & ~n2372 ;
  assign n2374 = n136 & ~n2373 ;
  assign n2386 = n2385 ^ n2374 ;
  assign n2387 = ~n2364 & ~n2386 ;
  assign n2433 = n2432 ^ n2387 ;
  assign n2434 = x134 & n2433 ;
  assign n2435 = n2434 ^ n2433 ;
  assign n2436 = n2435 ^ n2432 ;
  assign n2442 = n171 & n194 ;
  assign n2441 = n160 & n298 ;
  assign n2443 = n2442 ^ n2441 ;
  assign n2438 = n148 & ~n210 ;
  assign n2439 = n2438 ^ n148 ;
  assign n2437 = n137 & n224 ;
  assign n2440 = n2439 ^ n2437 ;
  assign n2444 = n2443 ^ n2440 ;
  assign n2446 = n298 & n2087 ;
  assign n2445 = n194 & n2085 ;
  assign n2447 = n2446 ^ n2445 ;
  assign n2448 = n2447 ^ n289 ;
  assign n2449 = n2448 ^ n2440 ;
  assign n2450 = n2444 & n2449 ;
  assign n2451 = n2450 ^ n2447 ;
  assign n2452 = n2451 ^ n2440 ;
  assign n2454 = n148 & n329 ;
  assign n2453 = n137 & n308 ;
  assign n2455 = n2454 ^ n2453 ;
  assign n2457 = n171 & n319 ;
  assign n2456 = n160 & n253 ;
  assign n2458 = n2457 ^ n2456 ;
  assign n2459 = ~n2455 & ~n2458 ;
  assign n2460 = n244 & n2459 ;
  assign n2461 = n2460 ^ n244 ;
  assign n2462 = n2452 & n2461 ;
  assign n2463 = n2462 ^ n2452 ;
  assign n2464 = n2463 ^ n2461 ;
  assign n2474 = n148 & n376 ;
  assign n2473 = n137 & n355 ;
  assign n2475 = n2474 ^ n2473 ;
  assign n2477 = n171 & n366 ;
  assign n2476 = n146 & n160 ;
  assign n2478 = n2477 ^ n2476 ;
  assign n2479 = ~n2475 & ~n2478 ;
  assign n2480 = n136 & n2479 ;
  assign n2481 = n2480 ^ n136 ;
  assign n2466 = n148 & n180 ;
  assign n2465 = n137 & n157 ;
  assign n2467 = n2466 ^ n2465 ;
  assign n2469 = n169 & n171 ;
  assign n2468 = n160 & n235 ;
  assign n2470 = n2469 ^ n2468 ;
  assign n2471 = ~n2467 & ~n2470 ;
  assign n2472 = n214 & ~n2471 ;
  assign n2482 = n2481 ^ n2472 ;
  assign n2523 = x134 & ~n2482 ;
  assign n2524 = ~n2464 & n2523 ;
  assign n2493 = n148 & n511 ;
  assign n2492 = n137 & n490 ;
  assign n2494 = n2493 ^ n2492 ;
  assign n2496 = n171 & n501 ;
  assign n2495 = n160 & n389 ;
  assign n2497 = n2496 ^ n2495 ;
  assign n2498 = ~n2494 & ~n2497 ;
  assign n2499 = n289 & n2498 ;
  assign n2500 = n2499 ^ n289 ;
  assign n2485 = n148 & n420 ;
  assign n2484 = n137 & n399 ;
  assign n2486 = n2485 ^ n2484 ;
  assign n2488 = n171 & n410 ;
  assign n2487 = n160 & n345 ;
  assign n2489 = n2488 ^ n2487 ;
  assign n2490 = ~n2486 & ~n2489 ;
  assign n2491 = n244 & ~n2490 ;
  assign n2501 = n2500 ^ n2491 ;
  assign n2511 = n148 & n467 ;
  assign n2510 = n137 & n446 ;
  assign n2512 = n2511 ^ n2510 ;
  assign n2514 = n171 & n457 ;
  assign n2513 = n160 & n480 ;
  assign n2515 = n2514 ^ n2513 ;
  assign n2516 = ~n2512 & ~n2515 ;
  assign n2517 = n214 & n2516 ;
  assign n2518 = n2517 ^ n214 ;
  assign n2503 = n148 & n284 ;
  assign n2502 = n137 & n263 ;
  assign n2504 = n2503 ^ n2502 ;
  assign n2506 = n160 & n436 ;
  assign n2505 = n171 & n274 ;
  assign n2507 = n2506 ^ n2505 ;
  assign n2508 = ~n2504 & ~n2507 ;
  assign n2509 = n136 & ~n2508 ;
  assign n2519 = n2518 ^ n2509 ;
  assign n2520 = ~n2501 & ~n2519 ;
  assign n2522 = x134 & n2520 ;
  assign n2525 = n2524 ^ n2522 ;
  assign n2483 = ~n2464 & ~n2482 ;
  assign n2521 = n2520 ^ n2483 ;
  assign n2526 = n2525 ^ n2521 ;
  assign n2527 = n2526 ^ n2483 ;
  assign n2528 = n160 & ~n1036 ;
  assign n2529 = n2528 ^ n160 ;
  assign n2530 = n171 & ~n1012 ;
  assign n2531 = n2530 ^ n171 ;
  assign n2532 = n2529 & n2531 ;
  assign n2533 = n2532 ^ n2529 ;
  assign n2534 = n2533 ^ n2531 ;
  assign n2535 = n137 & ~n962 ;
  assign n2536 = n2535 ^ n137 ;
  assign n2537 = n148 & ~n996 ;
  assign n2538 = n2537 ^ n148 ;
  assign n2539 = n2536 & n2538 ;
  assign n2540 = n2539 ^ n2536 ;
  assign n2541 = n2540 ^ n2538 ;
  assign n2542 = n289 & ~n2541 ;
  assign n2543 = ~n2534 & n2542 ;
  assign n2544 = n2543 ^ n289 ;
  assign n2546 = n148 & ~n1086 ;
  assign n2547 = n2546 ^ n148 ;
  assign n2545 = n137 & n1052 ;
  assign n2548 = n2547 ^ n2545 ;
  assign n2550 = n171 & ~n1070 ;
  assign n2551 = n2550 ^ n171 ;
  assign n2549 = n160 & n895 ;
  assign n2552 = n2551 ^ n2549 ;
  assign n2553 = ~n2548 & ~n2552 ;
  assign n2554 = n244 & n2553 ;
  assign n2555 = n2554 ^ n244 ;
  assign n2556 = n2544 & n2555 ;
  assign n2557 = n2556 ^ n2544 ;
  assign n2558 = n2557 ^ n2555 ;
  assign n2570 = n148 & ~n590 ;
  assign n2571 = n2570 ^ n148 ;
  assign n2569 = n137 & n556 ;
  assign n2572 = n2571 ^ n2569 ;
  assign n2574 = n171 & ~n574 ;
  assign n2575 = n2574 ^ n171 ;
  assign n2573 = n160 & n825 ;
  assign n2576 = n2575 ^ n2573 ;
  assign n2577 = ~n2572 & ~n2576 ;
  assign n2578 = n136 & n2577 ;
  assign n2579 = n2578 ^ n136 ;
  assign n2560 = n148 & ~n875 ;
  assign n2561 = n2560 ^ n148 ;
  assign n2559 = n137 & n841 ;
  assign n2562 = n2561 ^ n2559 ;
  assign n2564 = n171 & ~n859 ;
  assign n2565 = n2564 ^ n171 ;
  assign n2563 = n160 & n979 ;
  assign n2566 = n2565 ^ n2563 ;
  assign n2567 = ~n2562 & ~n2566 ;
  assign n2568 = n214 & ~n2567 ;
  assign n2580 = n2579 ^ n2568 ;
  assign n2629 = x134 & ~n2580 ;
  assign n2630 = ~n2558 & n2629 ;
  assign n2593 = n148 & ~n802 ;
  assign n2594 = n2593 ^ n148 ;
  assign n2592 = n137 & n768 ;
  assign n2595 = n2594 ^ n2592 ;
  assign n2597 = n171 & ~n786 ;
  assign n2598 = n2597 ^ n171 ;
  assign n2596 = n160 & n610 ;
  assign n2599 = n2598 ^ n2596 ;
  assign n2600 = ~n2595 & ~n2599 ;
  assign n2601 = n289 & n2600 ;
  assign n2602 = n2601 ^ n289 ;
  assign n2583 = n148 & ~n660 ;
  assign n2584 = n2583 ^ n148 ;
  assign n2582 = n137 & n626 ;
  assign n2585 = n2584 ^ n2582 ;
  assign n2587 = n171 & ~n644 ;
  assign n2588 = n2587 ^ n171 ;
  assign n2586 = n160 & n540 ;
  assign n2589 = n2588 ^ n2586 ;
  assign n2590 = ~n2585 & ~n2589 ;
  assign n2591 = n244 & ~n2590 ;
  assign n2603 = n2602 ^ n2591 ;
  assign n2615 = n148 & ~n732 ;
  assign n2616 = n2615 ^ n148 ;
  assign n2614 = n137 & n698 ;
  assign n2617 = n2616 ^ n2614 ;
  assign n2619 = n171 & ~n716 ;
  assign n2620 = n2619 ^ n171 ;
  assign n2618 = n160 & n752 ;
  assign n2621 = n2620 ^ n2618 ;
  assign n2622 = ~n2617 & ~n2621 ;
  assign n2623 = n214 & n2622 ;
  assign n2624 = n2623 ^ n214 ;
  assign n2605 = n148 & ~n945 ;
  assign n2606 = n2605 ^ n148 ;
  assign n2604 = n137 & n911 ;
  assign n2607 = n2606 ^ n2604 ;
  assign n2609 = n171 & ~n929 ;
  assign n2610 = n2609 ^ n171 ;
  assign n2608 = n160 & n682 ;
  assign n2611 = n2610 ^ n2608 ;
  assign n2612 = ~n2607 & ~n2611 ;
  assign n2613 = n136 & ~n2612 ;
  assign n2625 = n2624 ^ n2613 ;
  assign n2626 = ~n2603 & ~n2625 ;
  assign n2628 = x134 & n2626 ;
  assign n2631 = n2630 ^ n2628 ;
  assign n2581 = ~n2558 & ~n2580 ;
  assign n2627 = n2626 ^ n2581 ;
  assign n2632 = n2631 ^ n2627 ;
  assign n2633 = n2632 ^ n2581 ;
  assign n2680 = n148 & n1116 ;
  assign n2679 = n137 & n1106 ;
  assign n2681 = n2680 ^ n2679 ;
  assign n2683 = n171 & n1111 ;
  assign n2682 = n160 & n1196 ;
  assign n2684 = n2683 ^ n2682 ;
  assign n2685 = ~n2681 & ~n2684 ;
  assign n2686 = n136 & n2685 ;
  assign n2687 = n2686 ^ n136 ;
  assign n2672 = n148 & n1211 ;
  assign n2671 = n137 & n1201 ;
  assign n2673 = n2672 ^ n2671 ;
  assign n2675 = n171 & n1206 ;
  assign n2674 = n160 & n1243 ;
  assign n2676 = n2675 ^ n2674 ;
  assign n2677 = ~n2673 & ~n2676 ;
  assign n2678 = n214 & ~n2677 ;
  assign n2688 = n2687 ^ n2678 ;
  assign n2700 = n148 & n1289 ;
  assign n2699 = n137 & n1279 ;
  assign n2701 = n2700 ^ n2699 ;
  assign n2703 = n171 & n1284 ;
  assign n2702 = n160 & n1218 ;
  assign n2704 = n2703 ^ n2702 ;
  assign n2705 = ~n2701 & ~n2704 ;
  assign n2706 = n244 & n2705 ;
  assign n2707 = n2706 ^ n244 ;
  assign n2690 = n148 & ~n1266 ;
  assign n2691 = n2690 ^ n148 ;
  assign n2689 = n137 & n1248 ;
  assign n2692 = n2691 ^ n2689 ;
  assign n2694 = n171 & ~n1257 ;
  assign n2695 = n2694 ^ n171 ;
  assign n2693 = n160 & n1274 ;
  assign n2696 = n2695 ^ n2693 ;
  assign n2697 = ~n2692 & ~n2696 ;
  assign n2698 = n289 & ~n2697 ;
  assign n2708 = n2707 ^ n2698 ;
  assign n2709 = ~n2688 & ~n2708 ;
  assign n2643 = n148 & n1185 ;
  assign n2642 = n137 & n1175 ;
  assign n2644 = n2643 ^ n2642 ;
  assign n2646 = n171 & n1180 ;
  assign n2645 = n160 & n1123 ;
  assign n2647 = n2646 ^ n2645 ;
  assign n2648 = ~n2644 & ~n2647 ;
  assign n2649 = n289 & n2648 ;
  assign n2650 = n2649 ^ n289 ;
  assign n2635 = n148 & n1138 ;
  assign n2634 = n137 & n1128 ;
  assign n2636 = n2635 ^ n2634 ;
  assign n2638 = n171 & n1133 ;
  assign n2637 = n160 & n1101 ;
  assign n2639 = n2638 ^ n2637 ;
  assign n2640 = ~n2636 & ~n2639 ;
  assign n2641 = n244 & ~n2640 ;
  assign n2651 = n2650 ^ n2641 ;
  assign n2661 = n148 & n1162 ;
  assign n2660 = n137 & n1152 ;
  assign n2662 = n2661 ^ n2660 ;
  assign n2664 = n171 & n1157 ;
  assign n2663 = n160 & n1170 ;
  assign n2665 = n2664 ^ n2663 ;
  assign n2666 = ~n2662 & ~n2665 ;
  assign n2667 = n214 & n2666 ;
  assign n2668 = n2667 ^ n214 ;
  assign n2653 = n148 & n1233 ;
  assign n2652 = n137 & n1223 ;
  assign n2654 = n2653 ^ n2652 ;
  assign n2656 = n171 & n1228 ;
  assign n2655 = n160 & n1147 ;
  assign n2657 = n2656 ^ n2655 ;
  assign n2658 = ~n2654 & ~n2657 ;
  assign n2659 = n136 & ~n2658 ;
  assign n2669 = n2668 ^ n2659 ;
  assign n2670 = ~n2651 & ~n2669 ;
  assign n2710 = n2709 ^ n2670 ;
  assign n2711 = x134 & n2710 ;
  assign n2712 = n2711 ^ n2710 ;
  assign n2713 = n2712 ^ n2709 ;
  assign n2770 = n148 & ~n1483 ;
  assign n2771 = n2770 ^ n148 ;
  assign n2769 = n137 & n1461 ;
  assign n2772 = n2771 ^ n2769 ;
  assign n2774 = n171 & ~n1472 ;
  assign n2775 = n2774 ^ n171 ;
  assign n2773 = n160 & n1501 ;
  assign n2776 = n2775 ^ n2773 ;
  assign n2777 = ~n2772 & ~n2776 ;
  assign n2778 = n136 & n2777 ;
  assign n2779 = n2778 ^ n136 ;
  assign n2760 = n148 & ~n1534 ;
  assign n2761 = n2760 ^ n148 ;
  assign n2759 = n137 & n1512 ;
  assign n2762 = n2761 ^ n2759 ;
  assign n2764 = n171 & ~n1523 ;
  assign n2765 = n2764 ^ n171 ;
  assign n2763 = n160 & n1558 ;
  assign n2766 = n2765 ^ n2763 ;
  assign n2767 = ~n2762 & ~n2766 ;
  assign n2768 = n214 & ~n2767 ;
  assign n2780 = n2779 ^ n2768 ;
  assign n2792 = n148 & ~n1685 ;
  assign n2793 = n2792 ^ n148 ;
  assign n2791 = n137 & n1663 ;
  assign n2794 = n2793 ^ n2791 ;
  assign n2796 = n171 & ~n1674 ;
  assign n2797 = n2796 ^ n171 ;
  assign n2795 = n160 & n1604 ;
  assign n2798 = n2797 ^ n2795 ;
  assign n2799 = ~n2794 & ~n2798 ;
  assign n2800 = n244 & n2799 ;
  assign n2801 = n2800 ^ n244 ;
  assign n2783 = n137 & n1546 ;
  assign n2781 = n148 & ~n1589 ;
  assign n2782 = n2781 ^ n148 ;
  assign n2784 = n2783 ^ n2782 ;
  assign n2786 = n171 & ~n1573 ;
  assign n2787 = n2786 ^ n171 ;
  assign n2785 = n160 & n1652 ;
  assign n2788 = n2787 ^ n2785 ;
  assign n2789 = ~n2784 & ~n2788 ;
  assign n2790 = n289 & ~n2789 ;
  assign n2802 = n2801 ^ n2790 ;
  assign n2803 = ~n2780 & ~n2802 ;
  assign n2725 = n148 & ~n1343 ;
  assign n2726 = n2725 ^ n148 ;
  assign n2724 = n137 & n1321 ;
  assign n2727 = n2726 ^ n2724 ;
  assign n2729 = n171 & ~n1332 ;
  assign n2730 = n2729 ^ n171 ;
  assign n2728 = n160 & n1356 ;
  assign n2731 = n2730 ^ n2728 ;
  assign n2732 = ~n2727 & ~n2731 ;
  assign n2733 = n289 & n2732 ;
  assign n2734 = n2733 ^ n289 ;
  assign n2715 = n148 & ~n1389 ;
  assign n2716 = n2715 ^ n148 ;
  assign n2714 = n137 & n1367 ;
  assign n2717 = n2716 ^ n2714 ;
  assign n2719 = n171 & ~n1378 ;
  assign n2720 = n2719 ^ n171 ;
  assign n2718 = n160 & n1450 ;
  assign n2721 = n2720 ^ n2718 ;
  assign n2722 = ~n2717 & ~n2721 ;
  assign n2723 = n244 & ~n2722 ;
  assign n2735 = n2734 ^ n2723 ;
  assign n2747 = n148 & ~n1437 ;
  assign n2748 = n2747 ^ n148 ;
  assign n2746 = n137 & n1415 ;
  assign n2749 = n2748 ^ n2746 ;
  assign n2751 = n171 & ~n1426 ;
  assign n2752 = n2751 ^ n171 ;
  assign n2750 = n160 & n1310 ;
  assign n2753 = n2752 ^ n2750 ;
  assign n2754 = ~n2749 & ~n2753 ;
  assign n2755 = n214 & n2754 ;
  assign n2756 = n2755 ^ n214 ;
  assign n2737 = n148 & ~n1637 ;
  assign n2738 = n2737 ^ n148 ;
  assign n2736 = n137 & n1615 ;
  assign n2739 = n2738 ^ n2736 ;
  assign n2741 = n171 & ~n1626 ;
  assign n2742 = n2741 ^ n171 ;
  assign n2740 = n160 & n1404 ;
  assign n2743 = n2742 ^ n2740 ;
  assign n2744 = ~n2739 & ~n2743 ;
  assign n2745 = n136 & ~n2744 ;
  assign n2757 = n2756 ^ n2745 ;
  assign n2758 = ~n2735 & ~n2757 ;
  assign n2804 = n2803 ^ n2758 ;
  assign n2805 = x134 & n2804 ;
  assign n2806 = n2805 ^ n2804 ;
  assign n2807 = n2806 ^ n2803 ;
  assign n2808 = n183 & n214 ;
  assign n2809 = n2808 ^ n214 ;
  assign n2812 = n137 & n289 ;
  assign n2813 = n235 & n2812 ;
  assign n2814 = n2813 ^ n289 ;
  assign n2810 = n148 & n289 ;
  assign n2811 = n224 & n2810 ;
  assign n2815 = n2814 ^ n2811 ;
  assign n2816 = ~n213 & n2815 ;
  assign n2817 = n2816 ^ n289 ;
  assign n2818 = n2809 & n2817 ;
  assign n2819 = n2818 ^ n2809 ;
  assign n2820 = n2819 ^ n2817 ;
  assign n2822 = n244 & n332 ;
  assign n2823 = n2822 ^ n244 ;
  assign n2821 = n136 & ~n379 ;
  assign n2824 = n2823 ^ n2821 ;
  assign n2837 = x134 & ~n2824 ;
  assign n2838 = ~n2820 & n2837 ;
  assign n2827 = n289 & n514 ;
  assign n2828 = n2827 ^ n289 ;
  assign n2826 = n244 & ~n423 ;
  assign n2829 = n2828 ^ n2826 ;
  assign n2831 = n214 & n470 ;
  assign n2832 = n2831 ^ n214 ;
  assign n2830 = n136 & ~n287 ;
  assign n2833 = n2832 ^ n2830 ;
  assign n2834 = ~n2829 & ~n2833 ;
  assign n2836 = x134 & n2834 ;
  assign n2839 = n2838 ^ n2836 ;
  assign n2825 = ~n2820 & ~n2824 ;
  assign n2835 = n2834 ^ n2825 ;
  assign n2840 = n2839 ^ n2835 ;
  assign n2841 = n2840 ^ n2825 ;
  assign n2852 = n136 & n594 ;
  assign n2853 = n2852 ^ n136 ;
  assign n2851 = n214 & ~n879 ;
  assign n2854 = n2853 ^ n2851 ;
  assign n2856 = n244 & n1090 ;
  assign n2857 = n2856 ^ n244 ;
  assign n2855 = n289 & ~n1020 ;
  assign n2858 = n2857 ^ n2855 ;
  assign n2859 = ~n2854 & ~n2858 ;
  assign n2843 = n289 & n806 ;
  assign n2844 = n2843 ^ n289 ;
  assign n2842 = n244 & ~n664 ;
  assign n2845 = n2844 ^ n2842 ;
  assign n2847 = n214 & n736 ;
  assign n2848 = n2847 ^ n214 ;
  assign n2846 = n136 & ~n949 ;
  assign n2849 = n2848 ^ n2846 ;
  assign n2850 = ~n2845 & ~n2849 ;
  assign n2860 = n2859 ^ n2850 ;
  assign n2861 = x134 & n2860 ;
  assign n2862 = n2861 ^ n2860 ;
  assign n2863 = n2862 ^ n2859 ;
  assign n2874 = n136 & n1119 ;
  assign n2875 = n2874 ^ n136 ;
  assign n2873 = n214 & ~n1214 ;
  assign n2876 = n2875 ^ n2873 ;
  assign n2878 = n244 & n1292 ;
  assign n2879 = n2878 ^ n244 ;
  assign n2877 = n289 & ~n1270 ;
  assign n2880 = n2879 ^ n2877 ;
  assign n2881 = ~n2876 & ~n2880 ;
  assign n2865 = n289 & n1188 ;
  assign n2866 = n2865 ^ n289 ;
  assign n2864 = n244 & ~n1141 ;
  assign n2867 = n2866 ^ n2864 ;
  assign n2869 = n214 & n1165 ;
  assign n2870 = n2869 ^ n214 ;
  assign n2868 = n136 & ~n1236 ;
  assign n2871 = n2870 ^ n2868 ;
  assign n2872 = ~n2867 & ~n2871 ;
  assign n2882 = n2881 ^ n2872 ;
  assign n2883 = x134 & n2882 ;
  assign n2884 = n2883 ^ n2882 ;
  assign n2885 = n2884 ^ n2881 ;
  assign n2896 = n136 & n1487 ;
  assign n2897 = n2896 ^ n136 ;
  assign n2895 = n214 & ~n1538 ;
  assign n2898 = n2897 ^ n2895 ;
  assign n2900 = n289 & n1593 ;
  assign n2901 = n2900 ^ n289 ;
  assign n2899 = n244 & ~n1689 ;
  assign n2902 = n2901 ^ n2899 ;
  assign n2903 = ~n2898 & ~n2902 ;
  assign n2887 = n244 & n1393 ;
  assign n2888 = n2887 ^ n244 ;
  assign n2886 = n289 & ~n1347 ;
  assign n2889 = n2888 ^ n2886 ;
  assign n2891 = n136 & n1641 ;
  assign n2892 = n2891 ^ n136 ;
  assign n2890 = n214 & ~n1441 ;
  assign n2893 = n2892 ^ n2890 ;
  assign n2894 = ~n2889 & ~n2893 ;
  assign n2904 = n2903 ^ n2894 ;
  assign n2905 = x134 & n2904 ;
  assign n2906 = n2905 ^ n2904 ;
  assign n2907 = n2906 ^ n2903 ;
  assign n2908 = n136 & n1748 ;
  assign n2909 = n2908 ^ n136 ;
  assign n2911 = n169 & n2812 ;
  assign n2912 = n2911 ^ n289 ;
  assign n2910 = n235 & n2810 ;
  assign n2913 = n2912 ^ n2910 ;
  assign n2914 = ~n1704 & n2913 ;
  assign n2915 = n2914 ^ n289 ;
  assign n2916 = n2909 & n2915 ;
  assign n2917 = n2916 ^ n2909 ;
  assign n2918 = n2917 ^ n2915 ;
  assign n2920 = n214 & n1717 ;
  assign n2921 = n2920 ^ n214 ;
  assign n2919 = n244 & ~n1729 ;
  assign n2922 = n2921 ^ n2919 ;
  assign n2935 = x134 & ~n2922 ;
  assign n2936 = ~n2918 & n2935 ;
  assign n2925 = n289 & n1774 ;
  assign n2926 = n2925 ^ n289 ;
  assign n2924 = n244 & ~n1756 ;
  assign n2927 = n2926 ^ n2924 ;
  assign n2929 = n214 & n1766 ;
  assign n2930 = n2929 ^ n214 ;
  assign n2928 = n136 & ~n1737 ;
  assign n2931 = n2930 ^ n2928 ;
  assign n2932 = ~n2927 & ~n2931 ;
  assign n2934 = x134 & n2932 ;
  assign n2937 = n2936 ^ n2934 ;
  assign n2923 = ~n2918 & ~n2922 ;
  assign n2933 = n2932 ^ n2923 ;
  assign n2938 = n2937 ^ n2933 ;
  assign n2939 = n2938 ^ n2923 ;
  assign n2940 = n136 & n1853 ;
  assign n2941 = n2940 ^ n136 ;
  assign n2942 = n1799 ^ n289 ;
  assign n2943 = ~n289 & n2942 ;
  assign n2944 = n2943 ^ n289 ;
  assign n2945 = n2944 ^ n1792 ;
  assign n2946 = n1800 & n2945 ;
  assign n2947 = n2946 ^ n2943 ;
  assign n2948 = n2947 ^ n1792 ;
  assign n2949 = n2941 & n2948 ;
  assign n2950 = n2949 ^ n2941 ;
  assign n2951 = n2950 ^ n2948 ;
  assign n2953 = n214 & n1816 ;
  assign n2954 = n2953 ^ n214 ;
  assign n2952 = n244 & ~n1830 ;
  assign n2955 = n2954 ^ n2952 ;
  assign n2968 = x134 & ~n2955 ;
  assign n2969 = ~n2951 & n2968 ;
  assign n2958 = n289 & n1885 ;
  assign n2959 = n2958 ^ n289 ;
  assign n2957 = n244 & ~n1863 ;
  assign n2960 = n2959 ^ n2957 ;
  assign n2962 = n214 & n1875 ;
  assign n2963 = n2962 ^ n214 ;
  assign n2961 = n136 & ~n1840 ;
  assign n2964 = n2963 ^ n2961 ;
  assign n2965 = ~n2960 & ~n2964 ;
  assign n2967 = x134 & n2965 ;
  assign n2970 = n2969 ^ n2967 ;
  assign n2956 = ~n2951 & ~n2955 ;
  assign n2966 = n2965 ^ n2956 ;
  assign n2971 = n2970 ^ n2966 ;
  assign n2972 = n2971 ^ n2956 ;
  assign n2983 = n289 & n1940 ;
  assign n2984 = n2983 ^ n289 ;
  assign n2982 = n136 & ~n1903 ;
  assign n2985 = n2984 ^ n2982 ;
  assign n2987 = n214 & n1948 ;
  assign n2988 = n2987 ^ n214 ;
  assign n2986 = n244 & ~n1958 ;
  assign n2989 = n2988 ^ n2986 ;
  assign n2990 = ~n2985 & ~n2989 ;
  assign n2974 = n289 & n1929 ;
  assign n2975 = n2974 ^ n289 ;
  assign n2973 = n244 & ~n1911 ;
  assign n2976 = n2975 ^ n2973 ;
  assign n2978 = n214 & n1921 ;
  assign n2979 = n2978 ^ n214 ;
  assign n2977 = n136 & ~n1966 ;
  assign n2980 = n2979 ^ n2977 ;
  assign n2981 = ~n2976 & ~n2980 ;
  assign n2991 = n2990 ^ n2981 ;
  assign n2992 = x134 & n2991 ;
  assign n2993 = n2992 ^ n2991 ;
  assign n2994 = n2993 ^ n2990 ;
  assign n3005 = n214 & n2043 ;
  assign n3006 = n3005 ^ n214 ;
  assign n3004 = n289 & ~n2033 ;
  assign n3007 = n3006 ^ n3004 ;
  assign n3009 = n136 & n1983 ;
  assign n3010 = n3009 ^ n136 ;
  assign n3008 = n244 & ~n2055 ;
  assign n3011 = n3010 ^ n3008 ;
  assign n3012 = ~n3007 & ~n3011 ;
  assign n2996 = n136 & n2065 ;
  assign n2997 = n2996 ^ n136 ;
  assign n2995 = n244 & ~n1993 ;
  assign n2998 = n2997 ^ n2995 ;
  assign n3000 = n289 & n2015 ;
  assign n3001 = n3000 ^ n289 ;
  assign n2999 = n214 & ~n2005 ;
  assign n3002 = n3001 ^ n2999 ;
  assign n3003 = ~n2998 & ~n3002 ;
  assign n3013 = n3012 ^ n3003 ;
  assign n3014 = x134 & n3013 ;
  assign n3015 = n3014 ^ n3013 ;
  assign n3016 = n3015 ^ n3012 ;
  assign n3019 = n160 & ~n244 ;
  assign n3020 = n308 & n3019 ;
  assign n3017 = n171 & ~n244 ;
  assign n3018 = n298 & n3017 ;
  assign n3021 = n3020 ^ n3018 ;
  assign n3022 = n3021 ^ n244 ;
  assign n3023 = n3022 ^ n2080 ;
  assign n3024 = n2084 & n3023 ;
  assign n3025 = n3024 ^ n3021 ;
  assign n3026 = n3025 ^ n2080 ;
  assign n3027 = n136 & n2132 ;
  assign n3028 = n3027 ^ n136 ;
  assign n3029 = n3026 & n3028 ;
  assign n3030 = n3029 ^ n3026 ;
  assign n3031 = n3030 ^ n3028 ;
  assign n3033 = n214 & n2121 ;
  assign n3034 = n3033 ^ n214 ;
  assign n3032 = n289 & ~n2113 ;
  assign n3035 = n3034 ^ n3032 ;
  assign n3048 = x134 & ~n3035 ;
  assign n3049 = ~n3031 & n3048 ;
  assign n3038 = n136 & n2101 ;
  assign n3039 = n3038 ^ n136 ;
  assign n3037 = n244 & ~n2140 ;
  assign n3040 = n3039 ^ n3037 ;
  assign n3042 = n289 & n2158 ;
  assign n3043 = n3042 ^ n289 ;
  assign n3041 = n214 & ~n2150 ;
  assign n3044 = n3043 ^ n3041 ;
  assign n3045 = ~n3040 & ~n3044 ;
  assign n3047 = x134 & n3045 ;
  assign n3050 = n3049 ^ n3047 ;
  assign n3036 = ~n3031 & ~n3035 ;
  assign n3046 = n3045 ^ n3036 ;
  assign n3051 = n3050 ^ n3046 ;
  assign n3052 = n3051 ^ n3036 ;
  assign n3063 = n214 & n2233 ;
  assign n3064 = n3063 ^ n214 ;
  assign n3062 = n289 & ~n2223 ;
  assign n3065 = n3064 ^ n3062 ;
  assign n3067 = n136 & n2178 ;
  assign n3068 = n3067 ^ n136 ;
  assign n3066 = n244 & ~n2245 ;
  assign n3069 = n3068 ^ n3066 ;
  assign n3070 = ~n3065 & ~n3069 ;
  assign n3054 = n136 & n2255 ;
  assign n3055 = n3054 ^ n136 ;
  assign n3053 = n244 & ~n2188 ;
  assign n3056 = n3055 ^ n3053 ;
  assign n3058 = n289 & n2210 ;
  assign n3059 = n3058 ^ n289 ;
  assign n3057 = n214 & ~n2200 ;
  assign n3060 = n3059 ^ n3057 ;
  assign n3061 = ~n3056 & ~n3060 ;
  assign n3071 = n3070 ^ n3061 ;
  assign n3072 = x134 & n3071 ;
  assign n3073 = n3072 ^ n3071 ;
  assign n3074 = n3073 ^ n3070 ;
  assign n3085 = n214 & n2315 ;
  assign n3086 = n3085 ^ n214 ;
  assign n3084 = n289 & ~n2307 ;
  assign n3087 = n3086 ^ n3084 ;
  assign n3089 = n136 & n2270 ;
  assign n3090 = n3089 ^ n136 ;
  assign n3088 = n244 & ~n2326 ;
  assign n3091 = n3090 ^ n3088 ;
  assign n3092 = ~n3087 & ~n3091 ;
  assign n3076 = n289 & n2296 ;
  assign n3077 = n3076 ^ n289 ;
  assign n3075 = n244 & ~n2278 ;
  assign n3078 = n3077 ^ n3075 ;
  assign n3080 = n214 & n2288 ;
  assign n3081 = n3080 ^ n214 ;
  assign n3079 = n136 & ~n2334 ;
  assign n3082 = n3081 ^ n3079 ;
  assign n3083 = ~n3078 & ~n3082 ;
  assign n3093 = n3092 ^ n3083 ;
  assign n3094 = x134 & n3093 ;
  assign n3095 = n3094 ^ n3093 ;
  assign n3096 = n3095 ^ n3092 ;
  assign n3107 = n214 & n2406 ;
  assign n3108 = n3107 ^ n214 ;
  assign n3106 = n289 & ~n2396 ;
  assign n3109 = n3108 ^ n3106 ;
  assign n3111 = n136 & n2351 ;
  assign n3112 = n3111 ^ n136 ;
  assign n3110 = n244 & ~n2418 ;
  assign n3113 = n3112 ^ n3110 ;
  assign n3114 = ~n3109 & ~n3113 ;
  assign n3098 = n289 & n2383 ;
  assign n3099 = n3098 ^ n289 ;
  assign n3097 = n244 & ~n2361 ;
  assign n3100 = n3099 ^ n3097 ;
  assign n3102 = n214 & n2373 ;
  assign n3103 = n3102 ^ n214 ;
  assign n3101 = n136 & ~n2428 ;
  assign n3104 = n3103 ^ n3101 ;
  assign n3105 = ~n3100 & ~n3104 ;
  assign n3115 = n3114 ^ n3105 ;
  assign n3116 = x134 & n3115 ;
  assign n3117 = n3116 ^ n3115 ;
  assign n3118 = n3117 ^ n3114 ;
  assign n3120 = n298 & n3019 ;
  assign n3119 = n194 & n3017 ;
  assign n3121 = n3120 ^ n3119 ;
  assign n3122 = n3121 ^ n244 ;
  assign n3123 = n3122 ^ n2440 ;
  assign n3124 = n2444 & n3123 ;
  assign n3125 = n3124 ^ n3121 ;
  assign n3126 = n3125 ^ n2440 ;
  assign n3127 = n136 & n2490 ;
  assign n3128 = n3127 ^ n136 ;
  assign n3129 = n3126 & n3128 ;
  assign n3130 = n3129 ^ n3126 ;
  assign n3131 = n3130 ^ n3128 ;
  assign n3133 = n214 & n2479 ;
  assign n3134 = n3133 ^ n214 ;
  assign n3132 = n289 & ~n2471 ;
  assign n3135 = n3134 ^ n3132 ;
  assign n3148 = x134 & ~n3135 ;
  assign n3149 = ~n3131 & n3148 ;
  assign n3138 = n289 & n2516 ;
  assign n3139 = n3138 ^ n289 ;
  assign n3137 = n244 & ~n2498 ;
  assign n3140 = n3139 ^ n3137 ;
  assign n3142 = n214 & n2508 ;
  assign n3143 = n3142 ^ n214 ;
  assign n3141 = n136 & ~n2459 ;
  assign n3144 = n3143 ^ n3141 ;
  assign n3145 = ~n3140 & ~n3144 ;
  assign n3147 = x134 & n3145 ;
  assign n3150 = n3149 ^ n3147 ;
  assign n3136 = ~n3131 & ~n3135 ;
  assign n3146 = n3145 ^ n3136 ;
  assign n3151 = n3150 ^ n3146 ;
  assign n3152 = n3151 ^ n3136 ;
  assign n3153 = n244 & ~n2541 ;
  assign n3154 = ~n2534 & n3153 ;
  assign n3155 = n3154 ^ n244 ;
  assign n3156 = n136 & n2590 ;
  assign n3157 = n3156 ^ n136 ;
  assign n3158 = n3155 & n3157 ;
  assign n3159 = n3158 ^ n3155 ;
  assign n3160 = n3159 ^ n3157 ;
  assign n3162 = n214 & n2577 ;
  assign n3163 = n3162 ^ n214 ;
  assign n3161 = n289 & ~n2567 ;
  assign n3164 = n3163 ^ n3161 ;
  assign n3177 = x134 & ~n3164 ;
  assign n3178 = ~n3160 & n3177 ;
  assign n3167 = n289 & n2622 ;
  assign n3168 = n3167 ^ n289 ;
  assign n3166 = n244 & ~n2600 ;
  assign n3169 = n3168 ^ n3166 ;
  assign n3171 = n214 & n2612 ;
  assign n3172 = n3171 ^ n214 ;
  assign n3170 = n136 & ~n2553 ;
  assign n3173 = n3172 ^ n3170 ;
  assign n3174 = ~n3169 & ~n3173 ;
  assign n3176 = x134 & n3174 ;
  assign n3179 = n3178 ^ n3176 ;
  assign n3165 = ~n3160 & ~n3164 ;
  assign n3175 = n3174 ^ n3165 ;
  assign n3180 = n3179 ^ n3175 ;
  assign n3181 = n3180 ^ n3165 ;
  assign n3192 = n214 & n2685 ;
  assign n3193 = n3192 ^ n214 ;
  assign n3191 = n289 & ~n2677 ;
  assign n3194 = n3193 ^ n3191 ;
  assign n3196 = n136 & n2640 ;
  assign n3197 = n3196 ^ n136 ;
  assign n3195 = n244 & ~n2697 ;
  assign n3198 = n3197 ^ n3195 ;
  assign n3199 = ~n3194 & ~n3198 ;
  assign n3183 = n289 & n2666 ;
  assign n3184 = n3183 ^ n289 ;
  assign n3182 = n244 & ~n2648 ;
  assign n3185 = n3184 ^ n3182 ;
  assign n3187 = n214 & n2658 ;
  assign n3188 = n3187 ^ n214 ;
  assign n3186 = n136 & ~n2705 ;
  assign n3189 = n3188 ^ n3186 ;
  assign n3190 = ~n3185 & ~n3189 ;
  assign n3200 = n3199 ^ n3190 ;
  assign n3201 = x134 & n3200 ;
  assign n3202 = n3201 ^ n3200 ;
  assign n3203 = n3202 ^ n3199 ;
  assign n3214 = n214 & n2777 ;
  assign n3215 = n3214 ^ n214 ;
  assign n3213 = n289 & ~n2767 ;
  assign n3216 = n3215 ^ n3213 ;
  assign n3218 = n136 & n2722 ;
  assign n3219 = n3218 ^ n136 ;
  assign n3217 = n244 & ~n2789 ;
  assign n3220 = n3219 ^ n3217 ;
  assign n3221 = ~n3216 & ~n3220 ;
  assign n3205 = n289 & n2754 ;
  assign n3206 = n3205 ^ n289 ;
  assign n3204 = n244 & ~n2732 ;
  assign n3207 = n3206 ^ n3204 ;
  assign n3209 = n214 & n2744 ;
  assign n3210 = n3209 ^ n214 ;
  assign n3208 = n136 & ~n2799 ;
  assign n3211 = n3210 ^ n3208 ;
  assign n3212 = ~n3207 & ~n3211 ;
  assign n3222 = n3221 ^ n3212 ;
  assign n3223 = x134 & n3222 ;
  assign n3224 = n3223 ^ n3222 ;
  assign n3225 = n3224 ^ n3221 ;
  assign n3226 = n183 & n289 ;
  assign n3227 = n3226 ^ n289 ;
  assign n3230 = n137 & n244 ;
  assign n3231 = n235 & n3230 ;
  assign n3232 = n3231 ^ n244 ;
  assign n3228 = n148 & n244 ;
  assign n3229 = n224 & n3228 ;
  assign n3233 = n3232 ^ n3229 ;
  assign n3234 = ~n213 & n3233 ;
  assign n3235 = n3234 ^ n244 ;
  assign n3236 = n3227 & n3235 ;
  assign n3237 = n3236 ^ n3227 ;
  assign n3238 = n3237 ^ n3235 ;
  assign n3240 = n136 & n423 ;
  assign n3241 = n3240 ^ n136 ;
  assign n3239 = n214 & ~n379 ;
  assign n3242 = n3241 ^ n3239 ;
  assign n3255 = x134 & ~n3242 ;
  assign n3256 = ~n3238 & n3255 ;
  assign n3245 = n289 & n470 ;
  assign n3246 = n3245 ^ n289 ;
  assign n3244 = n244 & ~n514 ;
  assign n3247 = n3246 ^ n3244 ;
  assign n3249 = n214 & n287 ;
  assign n3250 = n3249 ^ n214 ;
  assign n3248 = n136 & ~n332 ;
  assign n3251 = n3250 ^ n3248 ;
  assign n3252 = ~n3247 & ~n3251 ;
  assign n3254 = x134 & n3252 ;
  assign n3257 = n3256 ^ n3254 ;
  assign n3243 = ~n3238 & ~n3242 ;
  assign n3253 = n3252 ^ n3243 ;
  assign n3258 = n3257 ^ n3253 ;
  assign n3259 = n3258 ^ n3243 ;
  assign n3270 = n214 & n594 ;
  assign n3271 = n3270 ^ n214 ;
  assign n3269 = n289 & ~n879 ;
  assign n3272 = n3271 ^ n3269 ;
  assign n3274 = n136 & n664 ;
  assign n3275 = n3274 ^ n136 ;
  assign n3273 = n244 & ~n1020 ;
  assign n3276 = n3275 ^ n3273 ;
  assign n3277 = ~n3272 & ~n3276 ;
  assign n3261 = n289 & n736 ;
  assign n3262 = n3261 ^ n289 ;
  assign n3260 = n244 & ~n806 ;
  assign n3263 = n3262 ^ n3260 ;
  assign n3265 = n214 & n949 ;
  assign n3266 = n3265 ^ n214 ;
  assign n3264 = n136 & ~n1090 ;
  assign n3267 = n3266 ^ n3264 ;
  assign n3268 = ~n3263 & ~n3267 ;
  assign n3278 = n3277 ^ n3268 ;
  assign n3279 = x134 & n3278 ;
  assign n3280 = n3279 ^ n3278 ;
  assign n3281 = n3280 ^ n3277 ;
  assign n3292 = n214 & n1119 ;
  assign n3293 = n3292 ^ n214 ;
  assign n3291 = n289 & ~n1214 ;
  assign n3294 = n3293 ^ n3291 ;
  assign n3296 = n136 & n1141 ;
  assign n3297 = n3296 ^ n136 ;
  assign n3295 = n244 & ~n1270 ;
  assign n3298 = n3297 ^ n3295 ;
  assign n3299 = ~n3294 & ~n3298 ;
  assign n3283 = n289 & n1165 ;
  assign n3284 = n3283 ^ n289 ;
  assign n3282 = n244 & ~n1188 ;
  assign n3285 = n3284 ^ n3282 ;
  assign n3287 = n214 & n1236 ;
  assign n3288 = n3287 ^ n214 ;
  assign n3286 = n136 & ~n1292 ;
  assign n3289 = n3288 ^ n3286 ;
  assign n3290 = ~n3285 & ~n3289 ;
  assign n3300 = n3299 ^ n3290 ;
  assign n3301 = x134 & n3300 ;
  assign n3302 = n3301 ^ n3300 ;
  assign n3303 = n3302 ^ n3299 ;
  assign n3314 = n136 & n1393 ;
  assign n3315 = n3314 ^ n136 ;
  assign n3313 = n289 & ~n1538 ;
  assign n3316 = n3315 ^ n3313 ;
  assign n3318 = n214 & n1487 ;
  assign n3319 = n3318 ^ n214 ;
  assign n3317 = n244 & ~n1593 ;
  assign n3320 = n3319 ^ n3317 ;
  assign n3321 = ~n3316 & ~n3320 ;
  assign n3305 = n136 & n1689 ;
  assign n3306 = n3305 ^ n136 ;
  assign n3304 = n244 & ~n1347 ;
  assign n3307 = n3306 ^ n3304 ;
  assign n3309 = n214 & n1641 ;
  assign n3310 = n3309 ^ n214 ;
  assign n3308 = n289 & ~n1441 ;
  assign n3311 = n3310 ^ n3308 ;
  assign n3312 = ~n3307 & ~n3311 ;
  assign n3322 = n3321 ^ n3312 ;
  assign n3323 = x134 & n3322 ;
  assign n3324 = n3323 ^ n3322 ;
  assign n3325 = n3324 ^ n3321 ;
  assign n3326 = n289 & n1717 ;
  assign n3327 = n3326 ^ n289 ;
  assign n3329 = n169 & n3230 ;
  assign n3330 = n3329 ^ n244 ;
  assign n3328 = n235 & n3228 ;
  assign n3331 = n3330 ^ n3328 ;
  assign n3332 = ~n1704 & n3331 ;
  assign n3333 = n3332 ^ n244 ;
  assign n3334 = n3327 & n3333 ;
  assign n3335 = n3334 ^ n3327 ;
  assign n3336 = n3335 ^ n3333 ;
  assign n3338 = n136 & n1756 ;
  assign n3339 = n3338 ^ n136 ;
  assign n3337 = n214 & ~n1748 ;
  assign n3340 = n3339 ^ n3337 ;
  assign n3353 = x134 & ~n3340 ;
  assign n3354 = ~n3336 & n3353 ;
  assign n3343 = n289 & n1766 ;
  assign n3344 = n3343 ^ n289 ;
  assign n3342 = n244 & ~n1774 ;
  assign n3345 = n3344 ^ n3342 ;
  assign n3347 = n214 & n1737 ;
  assign n3348 = n3347 ^ n214 ;
  assign n3346 = n136 & ~n1729 ;
  assign n3349 = n3348 ^ n3346 ;
  assign n3350 = ~n3345 & ~n3349 ;
  assign n3352 = x134 & n3350 ;
  assign n3355 = n3354 ^ n3352 ;
  assign n3341 = ~n3336 & ~n3340 ;
  assign n3351 = n3350 ^ n3341 ;
  assign n3356 = n3355 ^ n3351 ;
  assign n3357 = n3356 ^ n3341 ;
  assign n3358 = n289 & n1816 ;
  assign n3359 = n3358 ^ n289 ;
  assign n3360 = n1799 ^ n244 ;
  assign n3361 = ~n244 & n3360 ;
  assign n3362 = n3361 ^ n244 ;
  assign n3363 = n3362 ^ n1792 ;
  assign n3364 = n1800 & n3363 ;
  assign n3365 = n3364 ^ n3361 ;
  assign n3366 = n3365 ^ n1792 ;
  assign n3367 = n3359 & n3366 ;
  assign n3368 = n3367 ^ n3359 ;
  assign n3369 = n3368 ^ n3366 ;
  assign n3371 = n136 & n1863 ;
  assign n3372 = n3371 ^ n136 ;
  assign n3370 = n214 & ~n1853 ;
  assign n3373 = n3372 ^ n3370 ;
  assign n3386 = x134 & ~n3373 ;
  assign n3387 = ~n3369 & n3386 ;
  assign n3376 = n289 & n1875 ;
  assign n3377 = n3376 ^ n289 ;
  assign n3375 = n244 & ~n1885 ;
  assign n3378 = n3377 ^ n3375 ;
  assign n3380 = n214 & n1840 ;
  assign n3381 = n3380 ^ n214 ;
  assign n3379 = n136 & ~n1830 ;
  assign n3382 = n3381 ^ n3379 ;
  assign n3383 = ~n3378 & ~n3382 ;
  assign n3385 = x134 & n3383 ;
  assign n3388 = n3387 ^ n3385 ;
  assign n3374 = ~n3369 & ~n3373 ;
  assign n3384 = n3383 ^ n3374 ;
  assign n3389 = n3388 ^ n3384 ;
  assign n3390 = n3389 ^ n3374 ;
  assign n3401 = n136 & n1911 ;
  assign n3402 = n3401 ^ n136 ;
  assign n3400 = n214 & ~n1903 ;
  assign n3403 = n3402 ^ n3400 ;
  assign n3405 = n244 & n1940 ;
  assign n3406 = n3405 ^ n244 ;
  assign n3404 = n289 & ~n1948 ;
  assign n3407 = n3406 ^ n3404 ;
  assign n3408 = ~n3403 & ~n3407 ;
  assign n3392 = n289 & n1921 ;
  assign n3393 = n3392 ^ n289 ;
  assign n3391 = n244 & ~n1929 ;
  assign n3394 = n3393 ^ n3391 ;
  assign n3396 = n214 & n1966 ;
  assign n3397 = n3396 ^ n214 ;
  assign n3395 = n136 & ~n1958 ;
  assign n3398 = n3397 ^ n3395 ;
  assign n3399 = ~n3394 & ~n3398 ;
  assign n3409 = n3408 ^ n3399 ;
  assign n3410 = x134 & n3409 ;
  assign n3411 = n3410 ^ n3409 ;
  assign n3412 = n3411 ^ n3408 ;
  assign n3423 = n289 & n2043 ;
  assign n3424 = n3423 ^ n289 ;
  assign n3422 = n244 & ~n2033 ;
  assign n3425 = n3424 ^ n3422 ;
  assign n3427 = n214 & n1983 ;
  assign n3428 = n3427 ^ n214 ;
  assign n3426 = n136 & ~n1993 ;
  assign n3429 = n3428 ^ n3426 ;
  assign n3430 = ~n3425 & ~n3429 ;
  assign n3414 = n136 & n2055 ;
  assign n3415 = n3414 ^ n136 ;
  assign n3413 = n214 & ~n2065 ;
  assign n3416 = n3415 ^ n3413 ;
  assign n3418 = n244 & n2015 ;
  assign n3419 = n3418 ^ n244 ;
  assign n3417 = n289 & ~n2005 ;
  assign n3420 = n3419 ^ n3417 ;
  assign n3421 = ~n3416 & ~n3420 ;
  assign n3431 = n3430 ^ n3421 ;
  assign n3432 = x134 & n3431 ;
  assign n3433 = n3432 ^ n3431 ;
  assign n3434 = n3433 ^ n3430 ;
  assign n3435 = n214 & n2101 ;
  assign n3436 = n3435 ^ n214 ;
  assign n3439 = ~n136 & n160 ;
  assign n3440 = n308 & n3439 ;
  assign n3437 = ~n136 & n171 ;
  assign n3438 = n298 & n3437 ;
  assign n3441 = n3440 ^ n3438 ;
  assign n3442 = n3441 ^ n136 ;
  assign n3443 = n3442 ^ n2080 ;
  assign n3444 = n2084 & n3443 ;
  assign n3445 = n3444 ^ n3441 ;
  assign n3446 = n3445 ^ n2080 ;
  assign n3447 = n3436 & n3446 ;
  assign n3448 = n3447 ^ n3436 ;
  assign n3449 = n3448 ^ n3446 ;
  assign n3451 = n244 & n2158 ;
  assign n3452 = n3451 ^ n244 ;
  assign n3450 = n289 & ~n2150 ;
  assign n3453 = n3452 ^ n3450 ;
  assign n3466 = x134 & ~n3453 ;
  assign n3467 = ~n3449 & n3466 ;
  assign n3456 = n289 & n2121 ;
  assign n3457 = n3456 ^ n289 ;
  assign n3455 = n244 & ~n2113 ;
  assign n3458 = n3457 ^ n3455 ;
  assign n3460 = n214 & n2132 ;
  assign n3461 = n3460 ^ n214 ;
  assign n3459 = n136 & ~n2140 ;
  assign n3462 = n3461 ^ n3459 ;
  assign n3463 = ~n3458 & ~n3462 ;
  assign n3465 = x134 & n3463 ;
  assign n3468 = n3467 ^ n3465 ;
  assign n3454 = ~n3449 & ~n3453 ;
  assign n3464 = n3463 ^ n3454 ;
  assign n3469 = n3468 ^ n3464 ;
  assign n3470 = n3469 ^ n3463 ;
  assign n3486 = n289 & n2233 ;
  assign n3487 = n3486 ^ n289 ;
  assign n3485 = n244 & ~n2223 ;
  assign n3488 = n3487 ^ n3485 ;
  assign n3490 = n214 & n2178 ;
  assign n3491 = n3490 ^ n214 ;
  assign n3489 = n136 & ~n2188 ;
  assign n3492 = n3491 ^ n3489 ;
  assign n3493 = ~n3488 & ~n3492 ;
  assign n3474 = n136 & n148 ;
  assign n3475 = n1012 & n3474 ;
  assign n3476 = ~n2244 & n3475 ;
  assign n3472 = n136 & ~n2239 ;
  assign n3473 = ~n2244 & n3472 ;
  assign n3477 = n3476 ^ n3473 ;
  assign n3478 = n3477 ^ n136 ;
  assign n3471 = n214 & ~n2255 ;
  assign n3479 = n3478 ^ n3471 ;
  assign n3481 = n244 & n2210 ;
  assign n3482 = n3481 ^ n244 ;
  assign n3480 = n289 & ~n2200 ;
  assign n3483 = n3482 ^ n3480 ;
  assign n3484 = ~n3479 & ~n3483 ;
  assign n3494 = n3493 ^ n3484 ;
  assign n3495 = x134 & n3494 ;
  assign n3496 = n3495 ^ n3494 ;
  assign n3497 = n3496 ^ n3493 ;
  assign n3508 = n289 & n2315 ;
  assign n3509 = n3508 ^ n289 ;
  assign n3507 = n244 & ~n2307 ;
  assign n3510 = n3509 ^ n3507 ;
  assign n3512 = n214 & n2270 ;
  assign n3513 = n3512 ^ n214 ;
  assign n3511 = n136 & ~n2278 ;
  assign n3514 = n3513 ^ n3511 ;
  assign n3515 = ~n3510 & ~n3514 ;
  assign n3499 = n289 & n2288 ;
  assign n3500 = n3499 ^ n289 ;
  assign n3498 = n244 & ~n2296 ;
  assign n3501 = n3500 ^ n3498 ;
  assign n3503 = n214 & n2334 ;
  assign n3504 = n3503 ^ n214 ;
  assign n3502 = n136 & ~n2326 ;
  assign n3505 = n3504 ^ n3502 ;
  assign n3506 = ~n3501 & ~n3505 ;
  assign n3516 = n3515 ^ n3506 ;
  assign n3517 = x134 & n3516 ;
  assign n3518 = n3517 ^ n3516 ;
  assign n3519 = n3518 ^ n3515 ;
  assign n3530 = n289 & n2406 ;
  assign n3531 = n3530 ^ n289 ;
  assign n3529 = n244 & ~n2396 ;
  assign n3532 = n3531 ^ n3529 ;
  assign n3534 = n214 & n2351 ;
  assign n3535 = n3534 ^ n214 ;
  assign n3533 = n136 & ~n2361 ;
  assign n3536 = n3535 ^ n3533 ;
  assign n3537 = ~n3532 & ~n3536 ;
  assign n3521 = n289 & n2373 ;
  assign n3522 = n3521 ^ n289 ;
  assign n3520 = n244 & ~n2383 ;
  assign n3523 = n3522 ^ n3520 ;
  assign n3525 = n214 & n2428 ;
  assign n3526 = n3525 ^ n214 ;
  assign n3524 = n136 & ~n2418 ;
  assign n3527 = n3526 ^ n3524 ;
  assign n3528 = ~n3523 & ~n3527 ;
  assign n3538 = n3537 ^ n3528 ;
  assign n3539 = x134 & n3538 ;
  assign n3540 = n3539 ^ n3538 ;
  assign n3541 = n3540 ^ n3537 ;
  assign n3543 = n298 & n3439 ;
  assign n3542 = n194 & n3437 ;
  assign n3544 = n3543 ^ n3542 ;
  assign n3545 = n3544 ^ n136 ;
  assign n3546 = n3545 ^ n2440 ;
  assign n3547 = n2444 & n3546 ;
  assign n3548 = n3547 ^ n3544 ;
  assign n3549 = n3548 ^ n2440 ;
  assign n3550 = n214 & n2459 ;
  assign n3551 = n3550 ^ n214 ;
  assign n3552 = n3549 & n3551 ;
  assign n3553 = n3552 ^ n3549 ;
  assign n3554 = n3553 ^ n3551 ;
  assign n3556 = n289 & n2508 ;
  assign n3557 = n3556 ^ n289 ;
  assign n3555 = n244 & ~n2516 ;
  assign n3558 = n3557 ^ n3555 ;
  assign n3571 = x134 & ~n3558 ;
  assign n3572 = ~n3554 & n3571 ;
  assign n3561 = n289 & n2479 ;
  assign n3562 = n3561 ^ n289 ;
  assign n3560 = n244 & ~n2471 ;
  assign n3563 = n3562 ^ n3560 ;
  assign n3565 = n214 & n2490 ;
  assign n3566 = n3565 ^ n214 ;
  assign n3564 = n136 & ~n2498 ;
  assign n3567 = n3566 ^ n3564 ;
  assign n3568 = ~n3563 & ~n3567 ;
  assign n3570 = x134 & n3568 ;
  assign n3573 = n3572 ^ n3570 ;
  assign n3559 = ~n3554 & ~n3558 ;
  assign n3569 = n3568 ^ n3559 ;
  assign n3574 = n3573 ^ n3569 ;
  assign n3575 = n3574 ^ n3568 ;
  assign n3576 = n136 & ~n2541 ;
  assign n3577 = ~n2534 & n3576 ;
  assign n3578 = n3577 ^ n136 ;
  assign n3579 = n214 & n2553 ;
  assign n3580 = n3579 ^ n214 ;
  assign n3581 = n3578 & n3580 ;
  assign n3582 = n3581 ^ n3578 ;
  assign n3583 = n3582 ^ n3580 ;
  assign n3585 = n289 & n2612 ;
  assign n3586 = n3585 ^ n289 ;
  assign n3584 = n244 & ~n2622 ;
  assign n3587 = n3586 ^ n3584 ;
  assign n3600 = x134 & ~n3587 ;
  assign n3601 = ~n3583 & n3600 ;
  assign n3590 = n289 & n2577 ;
  assign n3591 = n3590 ^ n289 ;
  assign n3589 = n244 & ~n2567 ;
  assign n3592 = n3591 ^ n3589 ;
  assign n3594 = n214 & n2590 ;
  assign n3595 = n3594 ^ n214 ;
  assign n3593 = n136 & ~n2600 ;
  assign n3596 = n3595 ^ n3593 ;
  assign n3597 = ~n3592 & ~n3596 ;
  assign n3599 = x134 & n3597 ;
  assign n3602 = n3601 ^ n3599 ;
  assign n3588 = ~n3583 & ~n3587 ;
  assign n3598 = n3597 ^ n3588 ;
  assign n3603 = n3602 ^ n3598 ;
  assign n3604 = n3603 ^ n3597 ;
  assign n3615 = n289 & n2685 ;
  assign n3616 = n3615 ^ n289 ;
  assign n3614 = n244 & ~n2677 ;
  assign n3617 = n3616 ^ n3614 ;
  assign n3619 = n214 & n2640 ;
  assign n3620 = n3619 ^ n214 ;
  assign n3618 = n136 & ~n2648 ;
  assign n3621 = n3620 ^ n3618 ;
  assign n3622 = ~n3617 & ~n3621 ;
  assign n3606 = n289 & n2658 ;
  assign n3607 = n3606 ^ n289 ;
  assign n3605 = n244 & ~n2666 ;
  assign n3608 = n3607 ^ n3605 ;
  assign n3610 = n214 & n2705 ;
  assign n3611 = n3610 ^ n214 ;
  assign n3609 = n136 & ~n2697 ;
  assign n3612 = n3611 ^ n3609 ;
  assign n3613 = ~n3608 & ~n3612 ;
  assign n3623 = n3622 ^ n3613 ;
  assign n3624 = x134 & n3623 ;
  assign n3625 = n3624 ^ n3623 ;
  assign n3626 = n3625 ^ n3622 ;
  assign n3637 = n289 & n2777 ;
  assign n3638 = n3637 ^ n289 ;
  assign n3636 = n244 & ~n2767 ;
  assign n3639 = n3638 ^ n3636 ;
  assign n3641 = n214 & n2722 ;
  assign n3642 = n3641 ^ n214 ;
  assign n3640 = n136 & ~n2732 ;
  assign n3643 = n3642 ^ n3640 ;
  assign n3644 = ~n3639 & ~n3643 ;
  assign n3628 = n289 & n2744 ;
  assign n3629 = n3628 ^ n289 ;
  assign n3627 = n244 & ~n2754 ;
  assign n3630 = n3629 ^ n3627 ;
  assign n3632 = n214 & n2799 ;
  assign n3633 = n3632 ^ n214 ;
  assign n3631 = n136 & ~n2789 ;
  assign n3634 = n3633 ^ n3631 ;
  assign n3635 = ~n3630 & ~n3634 ;
  assign n3645 = n3644 ^ n3635 ;
  assign n3646 = x134 & n3645 ;
  assign n3647 = n3646 ^ n3645 ;
  assign n3648 = n3647 ^ n3644 ;
  assign n3650 = n136 & n137 ;
  assign n3651 = n235 & n3650 ;
  assign n3652 = n3651 ^ n136 ;
  assign n3649 = n224 & n3474 ;
  assign n3653 = n3652 ^ n3649 ;
  assign n3654 = ~n213 & n3653 ;
  assign n3655 = n3654 ^ n136 ;
  assign n3656 = n214 & n332 ;
  assign n3657 = n3656 ^ n214 ;
  assign n3658 = n3655 & n3657 ;
  assign n3659 = n3658 ^ n3655 ;
  assign n3660 = n3659 ^ n3657 ;
  assign n3662 = n287 & n289 ;
  assign n3663 = n3662 ^ n289 ;
  assign n3661 = n244 & ~n470 ;
  assign n3664 = n3663 ^ n3661 ;
  assign n3677 = x134 & ~n3664 ;
  assign n3678 = ~n3660 & n3677 ;
  assign n3667 = n214 & n423 ;
  assign n3668 = n3667 ^ n214 ;
  assign n3666 = n289 & ~n379 ;
  assign n3669 = n3668 ^ n3666 ;
  assign n3671 = n136 & n514 ;
  assign n3672 = n3671 ^ n136 ;
  assign n3670 = ~n183 & n244 ;
  assign n3673 = n3672 ^ n3670 ;
  assign n3674 = ~n3669 & ~n3673 ;
  assign n3676 = x134 & n3674 ;
  assign n3679 = n3678 ^ n3676 ;
  assign n3665 = ~n3660 & ~n3664 ;
  assign n3675 = n3674 ^ n3665 ;
  assign n3680 = n3679 ^ n3675 ;
  assign n3681 = n3680 ^ n3674 ;
  assign n3692 = n289 & n594 ;
  assign n3693 = n3692 ^ n289 ;
  assign n3691 = n244 & ~n879 ;
  assign n3694 = n3693 ^ n3691 ;
  assign n3696 = n214 & n664 ;
  assign n3697 = n3696 ^ n214 ;
  assign n3695 = n136 & ~n806 ;
  assign n3698 = n3697 ^ n3695 ;
  assign n3699 = ~n3694 & ~n3698 ;
  assign n3683 = n289 & n949 ;
  assign n3684 = n3683 ^ n289 ;
  assign n3682 = n244 & ~n736 ;
  assign n3685 = n3684 ^ n3682 ;
  assign n3687 = n214 & n1090 ;
  assign n3688 = n3687 ^ n214 ;
  assign n3686 = n136 & ~n1020 ;
  assign n3689 = n3688 ^ n3686 ;
  assign n3690 = ~n3685 & ~n3689 ;
  assign n3700 = n3699 ^ n3690 ;
  assign n3701 = x134 & n3700 ;
  assign n3702 = n3701 ^ n3700 ;
  assign n3703 = n3702 ^ n3699 ;
  assign n3714 = n289 & n1119 ;
  assign n3715 = n3714 ^ n289 ;
  assign n3713 = n244 & ~n1214 ;
  assign n3716 = n3715 ^ n3713 ;
  assign n3718 = n214 & n1141 ;
  assign n3719 = n3718 ^ n214 ;
  assign n3717 = n136 & ~n1188 ;
  assign n3720 = n3719 ^ n3717 ;
  assign n3721 = ~n3716 & ~n3720 ;
  assign n3705 = n289 & n1236 ;
  assign n3706 = n3705 ^ n289 ;
  assign n3704 = n244 & ~n1165 ;
  assign n3707 = n3706 ^ n3704 ;
  assign n3709 = n214 & n1292 ;
  assign n3710 = n3709 ^ n214 ;
  assign n3708 = n136 & ~n1270 ;
  assign n3711 = n3710 ^ n3708 ;
  assign n3712 = ~n3707 & ~n3711 ;
  assign n3722 = n3721 ^ n3712 ;
  assign n3723 = x134 & n3722 ;
  assign n3724 = n3723 ^ n3722 ;
  assign n3725 = n3724 ^ n3721 ;
  assign n3736 = n136 & n1347 ;
  assign n3737 = n3736 ^ n136 ;
  assign n3735 = n244 & ~n1538 ;
  assign n3738 = n3737 ^ n3735 ;
  assign n3740 = n214 & n1393 ;
  assign n3741 = n3740 ^ n214 ;
  assign n3739 = n289 & ~n1487 ;
  assign n3742 = n3741 ^ n3739 ;
  assign n3743 = ~n3738 & ~n3742 ;
  assign n3727 = n214 & n1689 ;
  assign n3728 = n3727 ^ n214 ;
  assign n3726 = n136 & ~n1593 ;
  assign n3729 = n3728 ^ n3726 ;
  assign n3731 = n289 & n1641 ;
  assign n3732 = n3731 ^ n289 ;
  assign n3730 = n244 & ~n1441 ;
  assign n3733 = n3732 ^ n3730 ;
  assign n3734 = ~n3729 & ~n3733 ;
  assign n3744 = n3743 ^ n3734 ;
  assign n3745 = x134 & n3744 ;
  assign n3746 = n3745 ^ n3744 ;
  assign n3747 = n3746 ^ n3743 ;
  assign n3749 = n169 & n3650 ;
  assign n3750 = n3749 ^ n136 ;
  assign n3748 = n235 & n3474 ;
  assign n3751 = n3750 ^ n3748 ;
  assign n3752 = ~n1704 & n3751 ;
  assign n3753 = n3752 ^ n136 ;
  assign n3754 = n244 & n1766 ;
  assign n3755 = n3754 ^ n244 ;
  assign n3756 = n3753 & n3755 ;
  assign n3757 = n3756 ^ n3753 ;
  assign n3758 = n3757 ^ n3755 ;
  assign n3760 = n289 & n1737 ;
  assign n3761 = n3760 ^ n289 ;
  assign n3759 = n214 & ~n1729 ;
  assign n3762 = n3761 ^ n3759 ;
  assign n3775 = x134 & ~n3762 ;
  assign n3776 = ~n3758 & n3775 ;
  assign n3765 = n214 & n1756 ;
  assign n3766 = n3765 ^ n214 ;
  assign n3764 = n289 & ~n1748 ;
  assign n3767 = n3766 ^ n3764 ;
  assign n3769 = n244 & n1717 ;
  assign n3770 = n3769 ^ n244 ;
  assign n3768 = n136 & ~n1774 ;
  assign n3771 = n3770 ^ n3768 ;
  assign n3772 = ~n3767 & ~n3771 ;
  assign n3774 = x134 & n3772 ;
  assign n3777 = n3776 ^ n3774 ;
  assign n3763 = ~n3758 & ~n3762 ;
  assign n3773 = n3772 ^ n3763 ;
  assign n3778 = n3777 ^ n3773 ;
  assign n3779 = n3778 ^ n3772 ;
  assign n3780 = n1799 ^ n136 ;
  assign n3781 = ~n136 & n3780 ;
  assign n3782 = n3781 ^ n136 ;
  assign n3783 = n3782 ^ n1792 ;
  assign n3784 = n1800 & n3783 ;
  assign n3785 = n3784 ^ n3781 ;
  assign n3786 = n3785 ^ n1792 ;
  assign n3787 = n244 & n1875 ;
  assign n3788 = n3787 ^ n244 ;
  assign n3789 = n3786 & n3788 ;
  assign n3790 = n3789 ^ n3786 ;
  assign n3791 = n3790 ^ n3788 ;
  assign n3793 = n289 & n1840 ;
  assign n3794 = n3793 ^ n289 ;
  assign n3792 = n214 & ~n1830 ;
  assign n3795 = n3794 ^ n3792 ;
  assign n3808 = x134 & ~n3795 ;
  assign n3809 = ~n3791 & n3808 ;
  assign n3798 = n214 & n1863 ;
  assign n3799 = n3798 ^ n214 ;
  assign n3797 = n289 & ~n1853 ;
  assign n3800 = n3799 ^ n3797 ;
  assign n3802 = n244 & n1816 ;
  assign n3803 = n3802 ^ n244 ;
  assign n3801 = n136 & ~n1885 ;
  assign n3804 = n3803 ^ n3801 ;
  assign n3805 = ~n3800 & ~n3804 ;
  assign n3807 = x134 & n3805 ;
  assign n3810 = n3809 ^ n3807 ;
  assign n3796 = ~n3791 & ~n3795 ;
  assign n3806 = n3805 ^ n3796 ;
  assign n3811 = n3810 ^ n3806 ;
  assign n3812 = n3811 ^ n3805 ;
  assign n3823 = n214 & n1911 ;
  assign n3824 = n3823 ^ n214 ;
  assign n3822 = n289 & ~n1903 ;
  assign n3825 = n3824 ^ n3822 ;
  assign n3827 = n244 & n1948 ;
  assign n3828 = n3827 ^ n244 ;
  assign n3826 = n136 & ~n1929 ;
  assign n3829 = n3828 ^ n3826 ;
  assign n3830 = ~n3825 & ~n3829 ;
  assign n3814 = n244 & n1921 ;
  assign n3815 = n3814 ^ n244 ;
  assign n3813 = n136 & ~n1940 ;
  assign n3816 = n3815 ^ n3813 ;
  assign n3818 = n289 & n1966 ;
  assign n3819 = n3818 ^ n289 ;
  assign n3817 = n214 & ~n1958 ;
  assign n3820 = n3819 ^ n3817 ;
  assign n3821 = ~n3816 & ~n3820 ;
  assign n3831 = n3830 ^ n3821 ;
  assign n3832 = x134 & n3831 ;
  assign n3833 = n3832 ^ n3831 ;
  assign n3834 = n3833 ^ n3830 ;
  assign n3845 = n289 & n1983 ;
  assign n3846 = n3845 ^ n289 ;
  assign n3844 = n244 & ~n2043 ;
  assign n3847 = n3846 ^ n3844 ;
  assign n3849 = n214 & n1993 ;
  assign n3850 = n3849 ^ n214 ;
  assign n3848 = n136 & ~n2015 ;
  assign n3851 = n3850 ^ n3848 ;
  assign n3852 = ~n3847 & ~n3851 ;
  assign n3836 = n289 & n2065 ;
  assign n3837 = n3836 ^ n289 ;
  assign n3835 = n136 & ~n2033 ;
  assign n3838 = n3837 ^ n3835 ;
  assign n3840 = n214 & n2055 ;
  assign n3841 = n3840 ^ n214 ;
  assign n3839 = n244 & ~n2005 ;
  assign n3842 = n3841 ^ n3839 ;
  assign n3843 = ~n3838 & ~n3842 ;
  assign n3853 = n3852 ^ n3843 ;
  assign n3854 = x134 & n3853 ;
  assign n3855 = n3854 ^ n3853 ;
  assign n3856 = n3855 ^ n3852 ;
  assign n3857 = n244 & n2150 ;
  assign n3858 = n3857 ^ n244 ;
  assign n3861 = n160 & ~n214 ;
  assign n3862 = n308 & n3861 ;
  assign n3859 = n171 & ~n214 ;
  assign n3860 = n298 & n3859 ;
  assign n3863 = n3862 ^ n3860 ;
  assign n3864 = n3863 ^ n214 ;
  assign n3865 = n3864 ^ n2080 ;
  assign n3866 = n2084 & n3865 ;
  assign n3867 = n3866 ^ n3863 ;
  assign n3868 = n3867 ^ n2080 ;
  assign n3869 = n3858 & n3868 ;
  assign n3870 = n3869 ^ n3858 ;
  assign n3871 = n3870 ^ n3868 ;
  assign n3873 = n289 & n2101 ;
  assign n3874 = n3873 ^ n289 ;
  assign n3872 = n136 & ~n2113 ;
  assign n3875 = n3874 ^ n3872 ;
  assign n3888 = x134 & ~n3875 ;
  assign n3889 = ~n3871 & n3888 ;
  assign n3878 = n289 & n2132 ;
  assign n3879 = n3878 ^ n289 ;
  assign n3877 = n244 & ~n2121 ;
  assign n3880 = n3879 ^ n3877 ;
  assign n3882 = n214 & n2140 ;
  assign n3883 = n3882 ^ n214 ;
  assign n3881 = n136 & ~n2158 ;
  assign n3884 = n3883 ^ n3881 ;
  assign n3885 = ~n3880 & ~n3884 ;
  assign n3887 = x134 & n3885 ;
  assign n3890 = n3889 ^ n3887 ;
  assign n3876 = ~n3871 & ~n3875 ;
  assign n3886 = n3885 ^ n3876 ;
  assign n3891 = n3890 ^ n3886 ;
  assign n3892 = n3891 ^ n3885 ;
  assign n3907 = n289 & n2178 ;
  assign n3908 = n3907 ^ n289 ;
  assign n3906 = n244 & ~n2233 ;
  assign n3909 = n3908 ^ n3906 ;
  assign n3911 = n214 & n2188 ;
  assign n3912 = n3911 ^ n214 ;
  assign n3910 = n136 & ~n2210 ;
  assign n3913 = n3912 ^ n3910 ;
  assign n3914 = ~n3909 & ~n3913 ;
  assign n3894 = n289 & n2255 ;
  assign n3895 = n3894 ^ n289 ;
  assign n3893 = n136 & ~n2223 ;
  assign n3896 = n3895 ^ n3893 ;
  assign n3900 = n215 & n1012 ;
  assign n3901 = ~n2244 & n3900 ;
  assign n3898 = n214 & ~n2239 ;
  assign n3899 = ~n2244 & n3898 ;
  assign n3902 = n3901 ^ n3899 ;
  assign n3903 = n3902 ^ n214 ;
  assign n3897 = n244 & ~n2200 ;
  assign n3904 = n3903 ^ n3897 ;
  assign n3905 = ~n3896 & ~n3904 ;
  assign n3915 = n3914 ^ n3905 ;
  assign n3916 = x134 & n3915 ;
  assign n3917 = n3916 ^ n3915 ;
  assign n3918 = n3917 ^ n3914 ;
  assign n3929 = n289 & n2270 ;
  assign n3930 = n3929 ^ n289 ;
  assign n3928 = n244 & ~n2315 ;
  assign n3931 = n3930 ^ n3928 ;
  assign n3933 = n214 & n2278 ;
  assign n3934 = n3933 ^ n214 ;
  assign n3932 = n136 & ~n2296 ;
  assign n3935 = n3934 ^ n3932 ;
  assign n3936 = ~n3931 & ~n3935 ;
  assign n3920 = n244 & n2288 ;
  assign n3921 = n3920 ^ n244 ;
  assign n3919 = n136 & ~n2307 ;
  assign n3922 = n3921 ^ n3919 ;
  assign n3924 = n289 & n2334 ;
  assign n3925 = n3924 ^ n289 ;
  assign n3923 = n214 & ~n2326 ;
  assign n3926 = n3925 ^ n3923 ;
  assign n3927 = ~n3922 & ~n3926 ;
  assign n3937 = n3936 ^ n3927 ;
  assign n3938 = x134 & n3937 ;
  assign n3939 = n3938 ^ n3937 ;
  assign n3940 = n3939 ^ n3936 ;
  assign n3951 = n289 & n2351 ;
  assign n3952 = n3951 ^ n289 ;
  assign n3950 = n244 & ~n2406 ;
  assign n3953 = n3952 ^ n3950 ;
  assign n3955 = n214 & n2361 ;
  assign n3956 = n3955 ^ n214 ;
  assign n3954 = n136 & ~n2383 ;
  assign n3957 = n3956 ^ n3954 ;
  assign n3958 = ~n3953 & ~n3957 ;
  assign n3942 = n244 & n2373 ;
  assign n3943 = n3942 ^ n244 ;
  assign n3941 = n136 & ~n2396 ;
  assign n3944 = n3943 ^ n3941 ;
  assign n3946 = n289 & n2428 ;
  assign n3947 = n3946 ^ n289 ;
  assign n3945 = n214 & ~n2418 ;
  assign n3948 = n3947 ^ n3945 ;
  assign n3949 = ~n3944 & ~n3948 ;
  assign n3959 = n3958 ^ n3949 ;
  assign n3960 = x134 & n3959 ;
  assign n3961 = n3960 ^ n3959 ;
  assign n3962 = n3961 ^ n3958 ;
  assign n3964 = n298 & n3861 ;
  assign n3963 = n194 & n3859 ;
  assign n3965 = n3964 ^ n3963 ;
  assign n3966 = n3965 ^ n214 ;
  assign n3967 = n3966 ^ n2440 ;
  assign n3968 = n2444 & n3967 ;
  assign n3969 = n3968 ^ n3965 ;
  assign n3970 = n3969 ^ n2440 ;
  assign n3971 = n289 & n2459 ;
  assign n3972 = n3971 ^ n289 ;
  assign n3973 = n3970 & n3972 ;
  assign n3974 = n3973 ^ n3970 ;
  assign n3975 = n3974 ^ n3972 ;
  assign n3977 = n244 & n2508 ;
  assign n3978 = n3977 ^ n244 ;
  assign n3976 = n136 & ~n2471 ;
  assign n3979 = n3978 ^ n3976 ;
  assign n3992 = x134 & ~n3979 ;
  assign n3993 = ~n3975 & n3992 ;
  assign n3982 = n289 & n2490 ;
  assign n3983 = n3982 ^ n289 ;
  assign n3981 = n244 & ~n2479 ;
  assign n3984 = n3983 ^ n3981 ;
  assign n3986 = n214 & n2498 ;
  assign n3987 = n3986 ^ n214 ;
  assign n3985 = n136 & ~n2516 ;
  assign n3988 = n3987 ^ n3985 ;
  assign n3989 = ~n3984 & ~n3988 ;
  assign n3991 = x134 & n3989 ;
  assign n3994 = n3993 ^ n3991 ;
  assign n3980 = ~n3975 & ~n3979 ;
  assign n3990 = n3989 ^ n3980 ;
  assign n3995 = n3994 ^ n3990 ;
  assign n3996 = n3995 ^ n3989 ;
  assign n3997 = n214 & ~n2541 ;
  assign n3998 = ~n2534 & n3997 ;
  assign n3999 = n3998 ^ n214 ;
  assign n4000 = n289 & n2553 ;
  assign n4001 = n4000 ^ n289 ;
  assign n4002 = n3999 & n4001 ;
  assign n4003 = n4002 ^ n3999 ;
  assign n4004 = n4003 ^ n4001 ;
  assign n4006 = n244 & n2612 ;
  assign n4007 = n4006 ^ n244 ;
  assign n4005 = n136 & ~n2567 ;
  assign n4008 = n4007 ^ n4005 ;
  assign n4021 = x134 & ~n4008 ;
  assign n4022 = ~n4004 & n4021 ;
  assign n4011 = n289 & n2590 ;
  assign n4012 = n4011 ^ n289 ;
  assign n4010 = n244 & ~n2577 ;
  assign n4013 = n4012 ^ n4010 ;
  assign n4015 = n214 & n2600 ;
  assign n4016 = n4015 ^ n214 ;
  assign n4014 = n136 & ~n2622 ;
  assign n4017 = n4016 ^ n4014 ;
  assign n4018 = ~n4013 & ~n4017 ;
  assign n4020 = x134 & n4018 ;
  assign n4023 = n4022 ^ n4020 ;
  assign n4009 = ~n4004 & ~n4008 ;
  assign n4019 = n4018 ^ n4009 ;
  assign n4024 = n4023 ^ n4019 ;
  assign n4025 = n4024 ^ n4018 ;
  assign n4036 = n289 & n2640 ;
  assign n4037 = n4036 ^ n289 ;
  assign n4035 = n244 & ~n2685 ;
  assign n4038 = n4037 ^ n4035 ;
  assign n4040 = n214 & n2648 ;
  assign n4041 = n4040 ^ n214 ;
  assign n4039 = n136 & ~n2666 ;
  assign n4042 = n4041 ^ n4039 ;
  assign n4043 = ~n4038 & ~n4042 ;
  assign n4027 = n244 & n2658 ;
  assign n4028 = n4027 ^ n244 ;
  assign n4026 = n136 & ~n2677 ;
  assign n4029 = n4028 ^ n4026 ;
  assign n4031 = n289 & n2705 ;
  assign n4032 = n4031 ^ n289 ;
  assign n4030 = n214 & ~n2697 ;
  assign n4033 = n4032 ^ n4030 ;
  assign n4034 = ~n4029 & ~n4033 ;
  assign n4044 = n4043 ^ n4034 ;
  assign n4045 = x134 & n4044 ;
  assign n4046 = n4045 ^ n4044 ;
  assign n4047 = n4046 ^ n4043 ;
  assign n4058 = n289 & n2722 ;
  assign n4059 = n4058 ^ n289 ;
  assign n4057 = n244 & ~n2777 ;
  assign n4060 = n4059 ^ n4057 ;
  assign n4062 = n214 & n2732 ;
  assign n4063 = n4062 ^ n214 ;
  assign n4061 = n136 & ~n2754 ;
  assign n4064 = n4063 ^ n4061 ;
  assign n4065 = ~n4060 & ~n4064 ;
  assign n4049 = n244 & n2744 ;
  assign n4050 = n4049 ^ n244 ;
  assign n4048 = n136 & ~n2767 ;
  assign n4051 = n4050 ^ n4048 ;
  assign n4053 = n289 & n2799 ;
  assign n4054 = n4053 ^ n289 ;
  assign n4052 = n214 & ~n2789 ;
  assign n4055 = n4054 ^ n4052 ;
  assign n4056 = ~n4051 & ~n4055 ;
  assign n4066 = n4065 ^ n4056 ;
  assign n4067 = x134 & n4066 ;
  assign n4068 = n4067 ^ n4066 ;
  assign n4069 = n4068 ^ n4065 ;
  assign n4070 = n523 ^ n336 ;
  assign n4071 = n1096 ^ n1094 ;
  assign n4072 = n1298 ^ n1296 ;
  assign n4073 = n1695 ^ n1693 ;
  assign n4074 = n1783 ^ n1741 ;
  assign n4075 = n1894 ^ n1844 ;
  assign n4076 = n1972 ^ n1970 ;
  assign n4077 = n2071 ^ n2069 ;
  assign n4078 = n2167 ^ n2125 ;
  assign n4079 = n2261 ^ n2259 ;
  assign n4080 = n2340 ^ n2338 ;
  assign n4081 = n2434 ^ n2432 ;
  assign n4082 = n2525 ^ n2483 ;
  assign n4083 = n2631 ^ n2581 ;
  assign n4084 = n2711 ^ n2709 ;
  assign n4085 = n2805 ^ n2803 ;
  assign n4086 = n2839 ^ n2825 ;
  assign n4087 = n2861 ^ n2859 ;
  assign n4088 = n2883 ^ n2881 ;
  assign n4089 = n2905 ^ n2903 ;
  assign n4090 = n2937 ^ n2923 ;
  assign n4091 = n2970 ^ n2956 ;
  assign n4092 = n2992 ^ n2990 ;
  assign n4093 = n3014 ^ n3012 ;
  assign n4094 = n3050 ^ n3036 ;
  assign n4095 = n3072 ^ n3070 ;
  assign n4096 = n3094 ^ n3092 ;
  assign n4097 = n3116 ^ n3114 ;
  assign n4098 = n3150 ^ n3136 ;
  assign n4099 = n3179 ^ n3165 ;
  assign n4100 = n3201 ^ n3199 ;
  assign n4101 = n3223 ^ n3221 ;
  assign n4102 = n3257 ^ n3243 ;
  assign n4103 = n3279 ^ n3277 ;
  assign n4104 = n3301 ^ n3299 ;
  assign n4105 = n3323 ^ n3321 ;
  assign n4106 = n3355 ^ n3341 ;
  assign n4107 = n3388 ^ n3374 ;
  assign n4108 = n3410 ^ n3408 ;
  assign n4109 = n3432 ^ n3430 ;
  assign n4110 = n3468 ^ n3463 ;
  assign n4111 = n3495 ^ n3493 ;
  assign n4112 = n3517 ^ n3515 ;
  assign n4113 = n3539 ^ n3537 ;
  assign n4114 = n3573 ^ n3568 ;
  assign n4115 = n3602 ^ n3597 ;
  assign n4116 = n3624 ^ n3622 ;
  assign n4117 = n3646 ^ n3644 ;
  assign n4118 = n3679 ^ n3674 ;
  assign n4119 = n3701 ^ n3699 ;
  assign n4120 = n3723 ^ n3721 ;
  assign n4121 = n3745 ^ n3743 ;
  assign n4122 = n3777 ^ n3772 ;
  assign n4123 = n3810 ^ n3805 ;
  assign n4124 = n3832 ^ n3830 ;
  assign n4125 = n3854 ^ n3852 ;
  assign n4126 = n3890 ^ n3885 ;
  assign n4127 = n3916 ^ n3914 ;
  assign n4128 = n3938 ^ n3936 ;
  assign n4129 = n3960 ^ n3958 ;
  assign n4130 = n3994 ^ n3989 ;
  assign n4131 = n4023 ^ n4018 ;
  assign n4132 = n4045 ^ n4043 ;
  assign n4133 = n4067 ^ n4065 ;
  assign y0 = ~n525 ;
  assign y1 = ~n1098 ;
  assign y2 = ~n1300 ;
  assign y3 = ~n1697 ;
  assign y4 = ~n1785 ;
  assign y5 = ~n1896 ;
  assign y6 = ~n1974 ;
  assign y7 = ~n2073 ;
  assign y8 = ~n2169 ;
  assign y9 = ~n2263 ;
  assign y10 = ~n2342 ;
  assign y11 = ~n2436 ;
  assign y12 = ~n2527 ;
  assign y13 = ~n2633 ;
  assign y14 = ~n2713 ;
  assign y15 = ~n2807 ;
  assign y16 = ~n2841 ;
  assign y17 = ~n2863 ;
  assign y18 = ~n2885 ;
  assign y19 = ~n2907 ;
  assign y20 = ~n2939 ;
  assign y21 = ~n2972 ;
  assign y22 = ~n2994 ;
  assign y23 = ~n3016 ;
  assign y24 = ~n3052 ;
  assign y25 = ~n3074 ;
  assign y26 = ~n3096 ;
  assign y27 = ~n3118 ;
  assign y28 = ~n3152 ;
  assign y29 = ~n3181 ;
  assign y30 = ~n3203 ;
  assign y31 = ~n3225 ;
  assign y32 = ~n3259 ;
  assign y33 = ~n3281 ;
  assign y34 = ~n3303 ;
  assign y35 = ~n3325 ;
  assign y36 = ~n3357 ;
  assign y37 = ~n3390 ;
  assign y38 = ~n3412 ;
  assign y39 = ~n3434 ;
  assign y40 = ~n3470 ;
  assign y41 = ~n3497 ;
  assign y42 = ~n3519 ;
  assign y43 = ~n3541 ;
  assign y44 = ~n3575 ;
  assign y45 = ~n3604 ;
  assign y46 = ~n3626 ;
  assign y47 = ~n3648 ;
  assign y48 = ~n3681 ;
  assign y49 = ~n3703 ;
  assign y50 = ~n3725 ;
  assign y51 = ~n3747 ;
  assign y52 = ~n3779 ;
  assign y53 = ~n3812 ;
  assign y54 = ~n3834 ;
  assign y55 = ~n3856 ;
  assign y56 = ~n3892 ;
  assign y57 = ~n3918 ;
  assign y58 = ~n3940 ;
  assign y59 = ~n3962 ;
  assign y60 = ~n3996 ;
  assign y61 = ~n4025 ;
  assign y62 = ~n4047 ;
  assign y63 = ~n4069 ;
  assign y64 = ~n4070 ;
  assign y65 = ~n4071 ;
  assign y66 = ~n4072 ;
  assign y67 = ~n4073 ;
  assign y68 = ~n4074 ;
  assign y69 = ~n4075 ;
  assign y70 = ~n4076 ;
  assign y71 = ~n4077 ;
  assign y72 = ~n4078 ;
  assign y73 = ~n4079 ;
  assign y74 = ~n4080 ;
  assign y75 = ~n4081 ;
  assign y76 = ~n4082 ;
  assign y77 = ~n4083 ;
  assign y78 = ~n4084 ;
  assign y79 = ~n4085 ;
  assign y80 = ~n4086 ;
  assign y81 = ~n4087 ;
  assign y82 = ~n4088 ;
  assign y83 = ~n4089 ;
  assign y84 = ~n4090 ;
  assign y85 = ~n4091 ;
  assign y86 = ~n4092 ;
  assign y87 = ~n4093 ;
  assign y88 = ~n4094 ;
  assign y89 = ~n4095 ;
  assign y90 = ~n4096 ;
  assign y91 = ~n4097 ;
  assign y92 = ~n4098 ;
  assign y93 = ~n4099 ;
  assign y94 = ~n4100 ;
  assign y95 = ~n4101 ;
  assign y96 = ~n4102 ;
  assign y97 = ~n4103 ;
  assign y98 = ~n4104 ;
  assign y99 = ~n4105 ;
  assign y100 = ~n4106 ;
  assign y101 = ~n4107 ;
  assign y102 = ~n4108 ;
  assign y103 = ~n4109 ;
  assign y104 = ~n4110 ;
  assign y105 = ~n4111 ;
  assign y106 = ~n4112 ;
  assign y107 = ~n4113 ;
  assign y108 = ~n4114 ;
  assign y109 = ~n4115 ;
  assign y110 = ~n4116 ;
  assign y111 = ~n4117 ;
  assign y112 = ~n4118 ;
  assign y113 = ~n4119 ;
  assign y114 = ~n4120 ;
  assign y115 = ~n4121 ;
  assign y116 = ~n4122 ;
  assign y117 = ~n4123 ;
  assign y118 = ~n4124 ;
  assign y119 = ~n4125 ;
  assign y120 = ~n4126 ;
  assign y121 = ~n4127 ;
  assign y122 = ~n4128 ;
  assign y123 = ~n4129 ;
  assign y124 = ~n4130 ;
  assign y125 = ~n4131 ;
  assign y126 = ~n4132 ;
  assign y127 = ~n4133 ;
endmodule
