module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 ;
  assign n257 = ~x143 & ~x159 ;
  assign n258 = ~x175 & ~x191 ;
  assign n259 = n257 & n258 ;
  assign n260 = ~x207 & ~x223 ;
  assign n261 = ~x239 & ~x255 ;
  assign n262 = n260 & n261 ;
  assign n263 = n259 & n262 ;
  assign n264 = ~x15 & ~x31 ;
  assign n265 = ~x47 & ~x63 ;
  assign n266 = n264 & n265 ;
  assign n267 = ~x79 & ~x95 ;
  assign n268 = ~x111 & ~x127 ;
  assign n269 = n267 & n268 ;
  assign n270 = n266 & n269 ;
  assign n271 = n263 & ~n270 ;
  assign n272 = ~x143 & x159 ;
  assign n273 = x143 & ~x159 ;
  assign n274 = ~x142 & x158 ;
  assign n275 = x142 & ~x158 ;
  assign n276 = ~x141 & x157 ;
  assign n277 = x141 & ~x157 ;
  assign n278 = ~x140 & x156 ;
  assign n279 = x140 & ~x156 ;
  assign n280 = ~x139 & x155 ;
  assign n281 = x139 & ~x155 ;
  assign n282 = ~x138 & x154 ;
  assign n283 = x138 & ~x154 ;
  assign n284 = ~x137 & x153 ;
  assign n285 = x137 & ~x153 ;
  assign n286 = ~x136 & x152 ;
  assign n287 = x136 & ~x152 ;
  assign n288 = ~x135 & x151 ;
  assign n289 = x135 & ~x151 ;
  assign n290 = ~x134 & x150 ;
  assign n291 = x134 & ~x150 ;
  assign n292 = ~x133 & x149 ;
  assign n293 = x133 & ~x149 ;
  assign n294 = ~x132 & x148 ;
  assign n295 = x132 & ~x148 ;
  assign n296 = ~x131 & x147 ;
  assign n297 = x131 & ~x147 ;
  assign n298 = ~x130 & x146 ;
  assign n299 = x130 & ~x146 ;
  assign n300 = ~x129 & x145 ;
  assign n301 = x129 & ~x145 ;
  assign n302 = x128 & ~x144 ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = ~n300 & ~n303 ;
  assign n305 = ~n299 & ~n304 ;
  assign n306 = ~n298 & ~n305 ;
  assign n307 = ~n297 & ~n306 ;
  assign n308 = ~n296 & ~n307 ;
  assign n309 = ~n295 & ~n308 ;
  assign n310 = ~n294 & ~n309 ;
  assign n311 = ~n293 & ~n310 ;
  assign n312 = ~n292 & ~n311 ;
  assign n313 = ~n291 & ~n312 ;
  assign n314 = ~n290 & ~n313 ;
  assign n315 = ~n289 & ~n314 ;
  assign n316 = ~n288 & ~n315 ;
  assign n317 = ~n287 & ~n316 ;
  assign n318 = ~n286 & ~n317 ;
  assign n319 = ~n285 & ~n318 ;
  assign n320 = ~n284 & ~n319 ;
  assign n321 = ~n283 & ~n320 ;
  assign n322 = ~n282 & ~n321 ;
  assign n323 = ~n281 & ~n322 ;
  assign n324 = ~n280 & ~n323 ;
  assign n325 = ~n279 & ~n324 ;
  assign n326 = ~n278 & ~n325 ;
  assign n327 = ~n277 & ~n326 ;
  assign n328 = ~n276 & ~n327 ;
  assign n329 = ~n275 & ~n328 ;
  assign n330 = ~n274 & ~n329 ;
  assign n331 = ~n273 & ~n330 ;
  assign n332 = ~n272 & ~n331 ;
  assign n333 = x152 & ~n332 ;
  assign n334 = x136 & n332 ;
  assign n335 = ~n333 & ~n334 ;
  assign n336 = n257 & ~n258 ;
  assign n337 = ~n257 & n258 ;
  assign n338 = x145 & ~n332 ;
  assign n339 = x129 & n332 ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = ~x175 & x191 ;
  assign n342 = x175 & ~x191 ;
  assign n343 = ~x174 & x190 ;
  assign n344 = x174 & ~x190 ;
  assign n345 = ~x173 & x189 ;
  assign n346 = x173 & ~x189 ;
  assign n347 = ~x172 & x188 ;
  assign n348 = x172 & ~x188 ;
  assign n349 = ~x171 & x187 ;
  assign n350 = x171 & ~x187 ;
  assign n351 = ~x170 & x186 ;
  assign n352 = x170 & ~x186 ;
  assign n353 = ~x169 & x185 ;
  assign n354 = x169 & ~x185 ;
  assign n355 = ~x168 & x184 ;
  assign n356 = x168 & ~x184 ;
  assign n357 = ~x167 & x183 ;
  assign n358 = x167 & ~x183 ;
  assign n359 = ~x166 & x182 ;
  assign n360 = x166 & ~x182 ;
  assign n361 = ~x165 & x181 ;
  assign n362 = x165 & ~x181 ;
  assign n363 = ~x164 & x180 ;
  assign n364 = x164 & ~x180 ;
  assign n365 = ~x163 & x179 ;
  assign n366 = x163 & ~x179 ;
  assign n367 = ~x162 & x178 ;
  assign n368 = x162 & ~x178 ;
  assign n369 = ~x161 & x177 ;
  assign n370 = x161 & ~x177 ;
  assign n371 = x160 & ~x176 ;
  assign n372 = ~n370 & ~n371 ;
  assign n373 = ~n369 & ~n372 ;
  assign n374 = ~n368 & ~n373 ;
  assign n375 = ~n367 & ~n374 ;
  assign n376 = ~n366 & ~n375 ;
  assign n377 = ~n365 & ~n376 ;
  assign n378 = ~n364 & ~n377 ;
  assign n379 = ~n363 & ~n378 ;
  assign n380 = ~n362 & ~n379 ;
  assign n381 = ~n361 & ~n380 ;
  assign n382 = ~n360 & ~n381 ;
  assign n383 = ~n359 & ~n382 ;
  assign n384 = ~n358 & ~n383 ;
  assign n385 = ~n357 & ~n384 ;
  assign n386 = ~n356 & ~n385 ;
  assign n387 = ~n355 & ~n386 ;
  assign n388 = ~n354 & ~n387 ;
  assign n389 = ~n353 & ~n388 ;
  assign n390 = ~n352 & ~n389 ;
  assign n391 = ~n351 & ~n390 ;
  assign n392 = ~n350 & ~n391 ;
  assign n393 = ~n349 & ~n392 ;
  assign n394 = ~n348 & ~n393 ;
  assign n395 = ~n347 & ~n394 ;
  assign n396 = ~n346 & ~n395 ;
  assign n397 = ~n345 & ~n396 ;
  assign n398 = ~n344 & ~n397 ;
  assign n399 = ~n343 & ~n398 ;
  assign n400 = ~n342 & ~n399 ;
  assign n401 = ~n341 & ~n400 ;
  assign n402 = x177 & ~n401 ;
  assign n403 = x161 & n401 ;
  assign n404 = ~n402 & ~n403 ;
  assign n405 = n340 & ~n404 ;
  assign n406 = x176 & ~n401 ;
  assign n407 = x160 & n401 ;
  assign n408 = ~n406 & ~n407 ;
  assign n409 = x144 & ~n332 ;
  assign n410 = x128 & n332 ;
  assign n411 = ~n409 & ~n410 ;
  assign n412 = n408 & ~n411 ;
  assign n413 = ~n405 & n412 ;
  assign n414 = x178 & ~n401 ;
  assign n415 = x162 & n401 ;
  assign n416 = ~n414 & ~n415 ;
  assign n417 = x146 & ~n332 ;
  assign n418 = x130 & n332 ;
  assign n419 = ~n417 & ~n418 ;
  assign n420 = n416 & ~n419 ;
  assign n421 = ~n340 & n404 ;
  assign n422 = ~n420 & ~n421 ;
  assign n423 = ~n413 & n422 ;
  assign n424 = x147 & ~n332 ;
  assign n425 = x131 & n332 ;
  assign n426 = ~n424 & ~n425 ;
  assign n427 = x179 & ~n401 ;
  assign n428 = x163 & n401 ;
  assign n429 = ~n427 & ~n428 ;
  assign n430 = n426 & ~n429 ;
  assign n431 = ~n416 & n419 ;
  assign n432 = ~n430 & ~n431 ;
  assign n433 = ~n423 & n432 ;
  assign n434 = ~n426 & n429 ;
  assign n435 = x180 & ~n401 ;
  assign n436 = x164 & n401 ;
  assign n437 = ~n435 & ~n436 ;
  assign n438 = x148 & ~n332 ;
  assign n439 = x132 & n332 ;
  assign n440 = ~n438 & ~n439 ;
  assign n441 = n437 & ~n440 ;
  assign n442 = ~n434 & ~n441 ;
  assign n443 = ~n433 & n442 ;
  assign n444 = x181 & ~n401 ;
  assign n445 = x165 & n401 ;
  assign n446 = ~n444 & ~n445 ;
  assign n447 = x149 & ~n332 ;
  assign n448 = x133 & n332 ;
  assign n449 = ~n447 & ~n448 ;
  assign n450 = ~n446 & n449 ;
  assign n451 = ~n437 & n440 ;
  assign n452 = ~n450 & ~n451 ;
  assign n453 = ~n443 & n452 ;
  assign n454 = x182 & ~n401 ;
  assign n455 = x166 & n401 ;
  assign n456 = ~n454 & ~n455 ;
  assign n457 = x150 & ~n332 ;
  assign n458 = x134 & n332 ;
  assign n459 = ~n457 & ~n458 ;
  assign n460 = n456 & ~n459 ;
  assign n461 = n446 & ~n449 ;
  assign n462 = ~n460 & ~n461 ;
  assign n463 = ~n453 & n462 ;
  assign n464 = x151 & ~n332 ;
  assign n465 = x135 & n332 ;
  assign n466 = ~n464 & ~n465 ;
  assign n467 = x183 & ~n401 ;
  assign n468 = x167 & n401 ;
  assign n469 = ~n467 & ~n468 ;
  assign n470 = n466 & ~n469 ;
  assign n471 = ~n456 & n459 ;
  assign n472 = ~n470 & ~n471 ;
  assign n473 = ~n463 & n472 ;
  assign n474 = ~n466 & n469 ;
  assign n475 = x184 & ~n401 ;
  assign n476 = x168 & n401 ;
  assign n477 = ~n475 & ~n476 ;
  assign n478 = ~n335 & n477 ;
  assign n479 = ~n474 & ~n478 ;
  assign n480 = ~n473 & n479 ;
  assign n481 = n335 & ~n477 ;
  assign n482 = x185 & ~n401 ;
  assign n483 = x169 & n401 ;
  assign n484 = ~n482 & ~n483 ;
  assign n485 = x153 & ~n332 ;
  assign n486 = x137 & n332 ;
  assign n487 = ~n485 & ~n486 ;
  assign n488 = ~n484 & n487 ;
  assign n489 = ~n481 & ~n488 ;
  assign n490 = ~n480 & n489 ;
  assign n491 = n484 & ~n487 ;
  assign n492 = x154 & ~n332 ;
  assign n493 = x138 & n332 ;
  assign n494 = ~n492 & ~n493 ;
  assign n495 = x186 & ~n401 ;
  assign n496 = x170 & n401 ;
  assign n497 = ~n495 & ~n496 ;
  assign n498 = ~n494 & n497 ;
  assign n499 = ~n491 & ~n498 ;
  assign n500 = ~n490 & n499 ;
  assign n501 = x187 & ~n401 ;
  assign n502 = x171 & n401 ;
  assign n503 = ~n501 & ~n502 ;
  assign n504 = x155 & ~n332 ;
  assign n505 = x139 & n332 ;
  assign n506 = ~n504 & ~n505 ;
  assign n507 = ~n503 & n506 ;
  assign n508 = n494 & ~n497 ;
  assign n509 = ~n507 & ~n508 ;
  assign n510 = ~n500 & n509 ;
  assign n511 = x188 & ~n401 ;
  assign n512 = x172 & n401 ;
  assign n513 = ~n511 & ~n512 ;
  assign n514 = x156 & ~n332 ;
  assign n515 = x140 & n332 ;
  assign n516 = ~n514 & ~n515 ;
  assign n517 = n513 & ~n516 ;
  assign n518 = n503 & ~n506 ;
  assign n519 = ~n517 & ~n518 ;
  assign n520 = ~n510 & n519 ;
  assign n521 = ~n513 & n516 ;
  assign n522 = x189 & ~n401 ;
  assign n523 = x173 & n401 ;
  assign n524 = ~n522 & ~n523 ;
  assign n525 = x157 & ~n332 ;
  assign n526 = x141 & n332 ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = ~n524 & n527 ;
  assign n529 = ~n521 & ~n528 ;
  assign n530 = ~n520 & n529 ;
  assign n531 = n524 & ~n527 ;
  assign n532 = x158 & ~n332 ;
  assign n533 = x142 & n332 ;
  assign n534 = ~n532 & ~n533 ;
  assign n535 = x190 & ~n401 ;
  assign n536 = x174 & n401 ;
  assign n537 = ~n535 & ~n536 ;
  assign n538 = ~n534 & n537 ;
  assign n539 = ~n531 & ~n538 ;
  assign n540 = ~n530 & n539 ;
  assign n541 = n534 & ~n537 ;
  assign n542 = ~n540 & ~n541 ;
  assign n543 = ~n337 & ~n542 ;
  assign n544 = ~n336 & ~n543 ;
  assign n545 = ~n335 & n544 ;
  assign n546 = ~n477 & ~n544 ;
  assign n547 = ~n545 & ~n546 ;
  assign n548 = ~n259 & n262 ;
  assign n549 = ~n340 & n544 ;
  assign n550 = ~n404 & ~n544 ;
  assign n551 = ~n549 & ~n550 ;
  assign n552 = ~x207 & x223 ;
  assign n553 = x207 & ~x223 ;
  assign n554 = ~x206 & x222 ;
  assign n555 = x206 & ~x222 ;
  assign n556 = ~x205 & x221 ;
  assign n557 = x205 & ~x221 ;
  assign n558 = ~x204 & x220 ;
  assign n559 = x204 & ~x220 ;
  assign n560 = ~x203 & x219 ;
  assign n561 = x203 & ~x219 ;
  assign n562 = ~x202 & x218 ;
  assign n563 = x202 & ~x218 ;
  assign n564 = ~x201 & x217 ;
  assign n565 = x201 & ~x217 ;
  assign n566 = ~x200 & x216 ;
  assign n567 = x200 & ~x216 ;
  assign n568 = ~x199 & x215 ;
  assign n569 = x199 & ~x215 ;
  assign n570 = ~x198 & x214 ;
  assign n571 = x198 & ~x214 ;
  assign n572 = ~x197 & x213 ;
  assign n573 = x197 & ~x213 ;
  assign n574 = ~x196 & x212 ;
  assign n575 = x196 & ~x212 ;
  assign n576 = ~x195 & x211 ;
  assign n577 = x195 & ~x211 ;
  assign n578 = ~x194 & x210 ;
  assign n579 = x194 & ~x210 ;
  assign n580 = ~x193 & x209 ;
  assign n581 = x193 & ~x209 ;
  assign n582 = x192 & ~x208 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = ~n580 & ~n583 ;
  assign n585 = ~n579 & ~n584 ;
  assign n586 = ~n578 & ~n585 ;
  assign n587 = ~n577 & ~n586 ;
  assign n588 = ~n576 & ~n587 ;
  assign n589 = ~n575 & ~n588 ;
  assign n590 = ~n574 & ~n589 ;
  assign n591 = ~n573 & ~n590 ;
  assign n592 = ~n572 & ~n591 ;
  assign n593 = ~n571 & ~n592 ;
  assign n594 = ~n570 & ~n593 ;
  assign n595 = ~n569 & ~n594 ;
  assign n596 = ~n568 & ~n595 ;
  assign n597 = ~n567 & ~n596 ;
  assign n598 = ~n566 & ~n597 ;
  assign n599 = ~n565 & ~n598 ;
  assign n600 = ~n564 & ~n599 ;
  assign n601 = ~n563 & ~n600 ;
  assign n602 = ~n562 & ~n601 ;
  assign n603 = ~n561 & ~n602 ;
  assign n604 = ~n560 & ~n603 ;
  assign n605 = ~n559 & ~n604 ;
  assign n606 = ~n558 & ~n605 ;
  assign n607 = ~n557 & ~n606 ;
  assign n608 = ~n556 & ~n607 ;
  assign n609 = ~n555 & ~n608 ;
  assign n610 = ~n554 & ~n609 ;
  assign n611 = ~n553 & ~n610 ;
  assign n612 = ~n552 & ~n611 ;
  assign n613 = x209 & ~n612 ;
  assign n614 = x193 & n612 ;
  assign n615 = ~n613 & ~n614 ;
  assign n616 = n260 & ~n261 ;
  assign n617 = ~n260 & n261 ;
  assign n618 = ~x239 & x255 ;
  assign n619 = x239 & ~x255 ;
  assign n620 = ~x238 & x254 ;
  assign n621 = x238 & ~x254 ;
  assign n622 = ~x237 & x253 ;
  assign n623 = x237 & ~x253 ;
  assign n624 = ~x236 & x252 ;
  assign n625 = x236 & ~x252 ;
  assign n626 = ~x235 & x251 ;
  assign n627 = x235 & ~x251 ;
  assign n628 = ~x234 & x250 ;
  assign n629 = x234 & ~x250 ;
  assign n630 = ~x233 & x249 ;
  assign n631 = x233 & ~x249 ;
  assign n632 = ~x232 & x248 ;
  assign n633 = x232 & ~x248 ;
  assign n634 = ~x231 & x247 ;
  assign n635 = x231 & ~x247 ;
  assign n636 = ~x230 & x246 ;
  assign n637 = x230 & ~x246 ;
  assign n638 = ~x229 & x245 ;
  assign n639 = x229 & ~x245 ;
  assign n640 = ~x228 & x244 ;
  assign n641 = x228 & ~x244 ;
  assign n642 = ~x227 & x243 ;
  assign n643 = x227 & ~x243 ;
  assign n644 = ~x226 & x242 ;
  assign n645 = x226 & ~x242 ;
  assign n646 = ~x225 & x241 ;
  assign n647 = x225 & ~x241 ;
  assign n648 = x224 & ~x240 ;
  assign n649 = ~n647 & ~n648 ;
  assign n650 = ~n646 & ~n649 ;
  assign n651 = ~n645 & ~n650 ;
  assign n652 = ~n644 & ~n651 ;
  assign n653 = ~n643 & ~n652 ;
  assign n654 = ~n642 & ~n653 ;
  assign n655 = ~n641 & ~n654 ;
  assign n656 = ~n640 & ~n655 ;
  assign n657 = ~n639 & ~n656 ;
  assign n658 = ~n638 & ~n657 ;
  assign n659 = ~n637 & ~n658 ;
  assign n660 = ~n636 & ~n659 ;
  assign n661 = ~n635 & ~n660 ;
  assign n662 = ~n634 & ~n661 ;
  assign n663 = ~n633 & ~n662 ;
  assign n664 = ~n632 & ~n663 ;
  assign n665 = ~n631 & ~n664 ;
  assign n666 = ~n630 & ~n665 ;
  assign n667 = ~n629 & ~n666 ;
  assign n668 = ~n628 & ~n667 ;
  assign n669 = ~n627 & ~n668 ;
  assign n670 = ~n626 & ~n669 ;
  assign n671 = ~n625 & ~n670 ;
  assign n672 = ~n624 & ~n671 ;
  assign n673 = ~n623 & ~n672 ;
  assign n674 = ~n622 & ~n673 ;
  assign n675 = ~n621 & ~n674 ;
  assign n676 = ~n620 & ~n675 ;
  assign n677 = ~n619 & ~n676 ;
  assign n678 = ~n618 & ~n677 ;
  assign n679 = x254 & ~n678 ;
  assign n680 = x238 & n678 ;
  assign n681 = ~n679 & ~n680 ;
  assign n682 = x222 & ~n612 ;
  assign n683 = x206 & n612 ;
  assign n684 = ~n682 & ~n683 ;
  assign n685 = ~n681 & n684 ;
  assign n686 = x241 & ~n678 ;
  assign n687 = x225 & n678 ;
  assign n688 = ~n686 & ~n687 ;
  assign n689 = n615 & ~n688 ;
  assign n690 = x240 & ~n678 ;
  assign n691 = x224 & n678 ;
  assign n692 = ~n690 & ~n691 ;
  assign n693 = x208 & ~n612 ;
  assign n694 = x192 & n612 ;
  assign n695 = ~n693 & ~n694 ;
  assign n696 = n692 & ~n695 ;
  assign n697 = ~n689 & n696 ;
  assign n698 = x242 & ~n678 ;
  assign n699 = x226 & n678 ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = x210 & ~n612 ;
  assign n702 = x194 & n612 ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = n700 & ~n703 ;
  assign n705 = ~n615 & n688 ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = ~n697 & n706 ;
  assign n708 = x211 & ~n612 ;
  assign n709 = x195 & n612 ;
  assign n710 = ~n708 & ~n709 ;
  assign n711 = x243 & ~n678 ;
  assign n712 = x227 & n678 ;
  assign n713 = ~n711 & ~n712 ;
  assign n714 = n710 & ~n713 ;
  assign n715 = ~n700 & n703 ;
  assign n716 = ~n714 & ~n715 ;
  assign n717 = ~n707 & n716 ;
  assign n718 = x244 & ~n678 ;
  assign n719 = x228 & n678 ;
  assign n720 = ~n718 & ~n719 ;
  assign n721 = x212 & ~n612 ;
  assign n722 = x196 & n612 ;
  assign n723 = ~n721 & ~n722 ;
  assign n724 = n720 & ~n723 ;
  assign n725 = ~n710 & n713 ;
  assign n726 = ~n724 & ~n725 ;
  assign n727 = ~n717 & n726 ;
  assign n728 = ~n720 & n723 ;
  assign n729 = x245 & ~n678 ;
  assign n730 = x229 & n678 ;
  assign n731 = ~n729 & ~n730 ;
  assign n732 = x213 & ~n612 ;
  assign n733 = x197 & n612 ;
  assign n734 = ~n732 & ~n733 ;
  assign n735 = ~n731 & n734 ;
  assign n736 = ~n728 & ~n735 ;
  assign n737 = ~n727 & n736 ;
  assign n738 = n731 & ~n734 ;
  assign n739 = x214 & ~n612 ;
  assign n740 = x198 & n612 ;
  assign n741 = ~n739 & ~n740 ;
  assign n742 = x246 & ~n678 ;
  assign n743 = x230 & n678 ;
  assign n744 = ~n742 & ~n743 ;
  assign n745 = ~n741 & n744 ;
  assign n746 = ~n738 & ~n745 ;
  assign n747 = ~n737 & n746 ;
  assign n748 = n741 & ~n744 ;
  assign n749 = x215 & ~n612 ;
  assign n750 = x199 & n612 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = x247 & ~n678 ;
  assign n753 = x231 & n678 ;
  assign n754 = ~n752 & ~n753 ;
  assign n755 = n751 & ~n754 ;
  assign n756 = ~n748 & ~n755 ;
  assign n757 = ~n747 & n756 ;
  assign n758 = x248 & ~n678 ;
  assign n759 = x232 & n678 ;
  assign n760 = ~n758 & ~n759 ;
  assign n761 = x216 & ~n612 ;
  assign n762 = x200 & n612 ;
  assign n763 = ~n761 & ~n762 ;
  assign n764 = n760 & ~n763 ;
  assign n765 = ~n751 & n754 ;
  assign n766 = ~n764 & ~n765 ;
  assign n767 = ~n757 & n766 ;
  assign n768 = ~n760 & n763 ;
  assign n769 = x217 & ~n612 ;
  assign n770 = x201 & n612 ;
  assign n771 = ~n769 & ~n770 ;
  assign n772 = x249 & ~n678 ;
  assign n773 = x233 & n678 ;
  assign n774 = ~n772 & ~n773 ;
  assign n775 = n771 & ~n774 ;
  assign n776 = ~n768 & ~n775 ;
  assign n777 = ~n767 & n776 ;
  assign n778 = ~n771 & n774 ;
  assign n779 = x218 & ~n612 ;
  assign n780 = x202 & n612 ;
  assign n781 = ~n779 & ~n780 ;
  assign n782 = x250 & ~n678 ;
  assign n783 = x234 & n678 ;
  assign n784 = ~n782 & ~n783 ;
  assign n785 = ~n781 & n784 ;
  assign n786 = ~n778 & ~n785 ;
  assign n787 = ~n777 & n786 ;
  assign n788 = x219 & ~n612 ;
  assign n789 = x203 & n612 ;
  assign n790 = ~n788 & ~n789 ;
  assign n791 = x251 & ~n678 ;
  assign n792 = x235 & n678 ;
  assign n793 = ~n791 & ~n792 ;
  assign n794 = n790 & ~n793 ;
  assign n795 = n781 & ~n784 ;
  assign n796 = ~n794 & ~n795 ;
  assign n797 = ~n787 & n796 ;
  assign n798 = x252 & ~n678 ;
  assign n799 = x236 & n678 ;
  assign n800 = ~n798 & ~n799 ;
  assign n801 = x220 & ~n612 ;
  assign n802 = x204 & n612 ;
  assign n803 = ~n801 & ~n802 ;
  assign n804 = n800 & ~n803 ;
  assign n805 = ~n790 & n793 ;
  assign n806 = ~n804 & ~n805 ;
  assign n807 = ~n797 & n806 ;
  assign n808 = ~n800 & n803 ;
  assign n809 = x253 & ~n678 ;
  assign n810 = x237 & n678 ;
  assign n811 = ~n809 & ~n810 ;
  assign n812 = x221 & ~n612 ;
  assign n813 = x205 & n612 ;
  assign n814 = ~n812 & ~n813 ;
  assign n815 = ~n811 & n814 ;
  assign n816 = ~n808 & ~n815 ;
  assign n817 = ~n807 & n816 ;
  assign n818 = n681 & ~n684 ;
  assign n819 = n811 & ~n814 ;
  assign n820 = ~n818 & ~n819 ;
  assign n821 = ~n817 & n820 ;
  assign n822 = ~n685 & ~n821 ;
  assign n823 = ~n617 & ~n822 ;
  assign n824 = ~n616 & ~n823 ;
  assign n825 = ~n615 & n824 ;
  assign n826 = ~n688 & ~n824 ;
  assign n827 = ~n825 & ~n826 ;
  assign n828 = n551 & ~n827 ;
  assign n829 = ~n695 & n824 ;
  assign n830 = ~n692 & ~n824 ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = ~n411 & n544 ;
  assign n833 = ~n408 & ~n544 ;
  assign n834 = ~n832 & ~n833 ;
  assign n835 = n831 & ~n834 ;
  assign n836 = ~n828 & n835 ;
  assign n837 = ~n703 & n824 ;
  assign n838 = ~n700 & ~n824 ;
  assign n839 = ~n837 & ~n838 ;
  assign n840 = ~n419 & n544 ;
  assign n841 = ~n416 & ~n544 ;
  assign n842 = ~n840 & ~n841 ;
  assign n843 = n839 & ~n842 ;
  assign n844 = ~n551 & n827 ;
  assign n845 = ~n843 & ~n844 ;
  assign n846 = ~n836 & n845 ;
  assign n847 = ~n839 & n842 ;
  assign n848 = ~n710 & n824 ;
  assign n849 = ~n713 & ~n824 ;
  assign n850 = ~n848 & ~n849 ;
  assign n851 = ~n426 & n544 ;
  assign n852 = ~n429 & ~n544 ;
  assign n853 = ~n851 & ~n852 ;
  assign n854 = ~n850 & n853 ;
  assign n855 = ~n847 & ~n854 ;
  assign n856 = ~n846 & n855 ;
  assign n857 = ~n723 & n824 ;
  assign n858 = ~n720 & ~n824 ;
  assign n859 = ~n857 & ~n858 ;
  assign n860 = ~n440 & n544 ;
  assign n861 = ~n437 & ~n544 ;
  assign n862 = ~n860 & ~n861 ;
  assign n863 = n859 & ~n862 ;
  assign n864 = n850 & ~n853 ;
  assign n865 = ~n863 & ~n864 ;
  assign n866 = ~n856 & n865 ;
  assign n867 = ~n449 & n544 ;
  assign n868 = ~n446 & ~n544 ;
  assign n869 = ~n867 & ~n868 ;
  assign n870 = ~n734 & n824 ;
  assign n871 = ~n731 & ~n824 ;
  assign n872 = ~n870 & ~n871 ;
  assign n873 = n869 & ~n872 ;
  assign n874 = ~n859 & n862 ;
  assign n875 = ~n873 & ~n874 ;
  assign n876 = ~n866 & n875 ;
  assign n877 = ~n741 & n824 ;
  assign n878 = ~n744 & ~n824 ;
  assign n879 = ~n877 & ~n878 ;
  assign n880 = ~n459 & n544 ;
  assign n881 = ~n456 & ~n544 ;
  assign n882 = ~n880 & ~n881 ;
  assign n883 = n879 & ~n882 ;
  assign n884 = ~n869 & n872 ;
  assign n885 = ~n883 & ~n884 ;
  assign n886 = ~n876 & n885 ;
  assign n887 = ~n466 & n544 ;
  assign n888 = ~n469 & ~n544 ;
  assign n889 = ~n887 & ~n888 ;
  assign n890 = ~n751 & n824 ;
  assign n891 = ~n754 & ~n824 ;
  assign n892 = ~n890 & ~n891 ;
  assign n893 = n889 & ~n892 ;
  assign n894 = ~n879 & n882 ;
  assign n895 = ~n893 & ~n894 ;
  assign n896 = ~n886 & n895 ;
  assign n897 = ~n763 & n824 ;
  assign n898 = ~n760 & ~n824 ;
  assign n899 = ~n897 & ~n898 ;
  assign n900 = ~n547 & n899 ;
  assign n901 = ~n889 & n892 ;
  assign n902 = ~n900 & ~n901 ;
  assign n903 = ~n896 & n902 ;
  assign n904 = n484 & ~n544 ;
  assign n905 = n487 & n544 ;
  assign n906 = ~n904 & ~n905 ;
  assign n907 = ~n771 & n824 ;
  assign n908 = ~n774 & ~n824 ;
  assign n909 = ~n907 & ~n908 ;
  assign n910 = ~n906 & ~n909 ;
  assign n911 = n547 & ~n899 ;
  assign n912 = ~n910 & ~n911 ;
  assign n913 = ~n903 & n912 ;
  assign n914 = ~n781 & n824 ;
  assign n915 = ~n784 & ~n824 ;
  assign n916 = ~n914 & ~n915 ;
  assign n917 = ~n494 & n544 ;
  assign n918 = ~n497 & ~n544 ;
  assign n919 = ~n917 & ~n918 ;
  assign n920 = n916 & ~n919 ;
  assign n921 = n906 & n909 ;
  assign n922 = ~n920 & ~n921 ;
  assign n923 = ~n913 & n922 ;
  assign n924 = ~n916 & n919 ;
  assign n925 = ~n790 & n824 ;
  assign n926 = ~n793 & ~n824 ;
  assign n927 = ~n925 & ~n926 ;
  assign n928 = ~n506 & n544 ;
  assign n929 = ~n503 & ~n544 ;
  assign n930 = ~n928 & ~n929 ;
  assign n931 = ~n927 & n930 ;
  assign n932 = ~n924 & ~n931 ;
  assign n933 = ~n923 & n932 ;
  assign n934 = n927 & ~n930 ;
  assign n935 = ~n516 & n544 ;
  assign n936 = ~n513 & ~n544 ;
  assign n937 = ~n935 & ~n936 ;
  assign n938 = ~n803 & n824 ;
  assign n939 = ~n800 & ~n824 ;
  assign n940 = ~n938 & ~n939 ;
  assign n941 = ~n937 & n940 ;
  assign n942 = ~n934 & ~n941 ;
  assign n943 = ~n933 & n942 ;
  assign n944 = n937 & ~n940 ;
  assign n945 = ~n527 & n544 ;
  assign n946 = ~n524 & ~n544 ;
  assign n947 = ~n945 & ~n946 ;
  assign n948 = ~n814 & n824 ;
  assign n949 = ~n811 & ~n824 ;
  assign n950 = ~n948 & ~n949 ;
  assign n951 = n947 & ~n950 ;
  assign n952 = ~n944 & ~n951 ;
  assign n953 = ~n943 & n952 ;
  assign n954 = ~n947 & n950 ;
  assign n955 = ~n534 & n544 ;
  assign n956 = ~n537 & ~n544 ;
  assign n957 = ~n955 & ~n956 ;
  assign n958 = ~n684 & n824 ;
  assign n959 = ~n681 & ~n824 ;
  assign n960 = ~n958 & ~n959 ;
  assign n961 = ~n957 & n960 ;
  assign n962 = ~n954 & ~n961 ;
  assign n963 = ~n953 & n962 ;
  assign n964 = n259 & ~n262 ;
  assign n965 = n957 & ~n960 ;
  assign n966 = ~n964 & ~n965 ;
  assign n967 = ~n963 & n966 ;
  assign n968 = ~n548 & ~n967 ;
  assign n969 = ~n547 & ~n968 ;
  assign n970 = ~n899 & n968 ;
  assign n971 = ~n969 & ~n970 ;
  assign n972 = ~x15 & x31 ;
  assign n973 = x15 & ~x31 ;
  assign n974 = ~x14 & x30 ;
  assign n975 = x14 & ~x30 ;
  assign n976 = ~x13 & x29 ;
  assign n977 = x13 & ~x29 ;
  assign n978 = ~x12 & x28 ;
  assign n979 = x12 & ~x28 ;
  assign n980 = ~x11 & x27 ;
  assign n981 = x11 & ~x27 ;
  assign n982 = ~x10 & x26 ;
  assign n983 = x10 & ~x26 ;
  assign n984 = ~x9 & x25 ;
  assign n985 = x9 & ~x25 ;
  assign n986 = ~x8 & x24 ;
  assign n987 = x8 & ~x24 ;
  assign n988 = ~x7 & x23 ;
  assign n989 = x7 & ~x23 ;
  assign n990 = ~x6 & x22 ;
  assign n991 = x6 & ~x22 ;
  assign n992 = ~x5 & x21 ;
  assign n993 = x5 & ~x21 ;
  assign n994 = ~x4 & x20 ;
  assign n995 = x4 & ~x20 ;
  assign n996 = ~x3 & x19 ;
  assign n997 = x3 & ~x19 ;
  assign n998 = ~x2 & x18 ;
  assign n999 = x2 & ~x18 ;
  assign n1000 = ~x1 & x17 ;
  assign n1001 = x1 & ~x17 ;
  assign n1002 = x0 & ~x16 ;
  assign n1003 = ~n1001 & ~n1002 ;
  assign n1004 = ~n1000 & ~n1003 ;
  assign n1005 = ~n999 & ~n1004 ;
  assign n1006 = ~n998 & ~n1005 ;
  assign n1007 = ~n997 & ~n1006 ;
  assign n1008 = ~n996 & ~n1007 ;
  assign n1009 = ~n995 & ~n1008 ;
  assign n1010 = ~n994 & ~n1009 ;
  assign n1011 = ~n993 & ~n1010 ;
  assign n1012 = ~n992 & ~n1011 ;
  assign n1013 = ~n991 & ~n1012 ;
  assign n1014 = ~n990 & ~n1013 ;
  assign n1015 = ~n989 & ~n1014 ;
  assign n1016 = ~n988 & ~n1015 ;
  assign n1017 = ~n987 & ~n1016 ;
  assign n1018 = ~n986 & ~n1017 ;
  assign n1019 = ~n985 & ~n1018 ;
  assign n1020 = ~n984 & ~n1019 ;
  assign n1021 = ~n983 & ~n1020 ;
  assign n1022 = ~n982 & ~n1021 ;
  assign n1023 = ~n981 & ~n1022 ;
  assign n1024 = ~n980 & ~n1023 ;
  assign n1025 = ~n979 & ~n1024 ;
  assign n1026 = ~n978 & ~n1025 ;
  assign n1027 = ~n977 & ~n1026 ;
  assign n1028 = ~n976 & ~n1027 ;
  assign n1029 = ~n975 & ~n1028 ;
  assign n1030 = ~n974 & ~n1029 ;
  assign n1031 = ~n973 & ~n1030 ;
  assign n1032 = ~n972 & ~n1031 ;
  assign n1033 = x24 & ~n1032 ;
  assign n1034 = x8 & n1032 ;
  assign n1035 = ~n1033 & ~n1034 ;
  assign n1036 = n264 & ~n265 ;
  assign n1037 = ~n264 & n265 ;
  assign n1038 = x17 & ~n1032 ;
  assign n1039 = x1 & n1032 ;
  assign n1040 = ~n1038 & ~n1039 ;
  assign n1041 = ~x47 & x63 ;
  assign n1042 = x47 & ~x63 ;
  assign n1043 = ~x46 & x62 ;
  assign n1044 = x46 & ~x62 ;
  assign n1045 = ~x45 & x61 ;
  assign n1046 = x45 & ~x61 ;
  assign n1047 = ~x44 & x60 ;
  assign n1048 = x44 & ~x60 ;
  assign n1049 = ~x43 & x59 ;
  assign n1050 = x43 & ~x59 ;
  assign n1051 = ~x42 & x58 ;
  assign n1052 = x42 & ~x58 ;
  assign n1053 = ~x41 & x57 ;
  assign n1054 = x41 & ~x57 ;
  assign n1055 = ~x40 & x56 ;
  assign n1056 = x40 & ~x56 ;
  assign n1057 = ~x39 & x55 ;
  assign n1058 = x39 & ~x55 ;
  assign n1059 = ~x38 & x54 ;
  assign n1060 = x38 & ~x54 ;
  assign n1061 = ~x37 & x53 ;
  assign n1062 = x37 & ~x53 ;
  assign n1063 = ~x36 & x52 ;
  assign n1064 = x36 & ~x52 ;
  assign n1065 = ~x35 & x51 ;
  assign n1066 = x35 & ~x51 ;
  assign n1067 = ~x34 & x50 ;
  assign n1068 = x34 & ~x50 ;
  assign n1069 = ~x33 & x49 ;
  assign n1070 = x33 & ~x49 ;
  assign n1071 = x32 & ~x48 ;
  assign n1072 = ~n1070 & ~n1071 ;
  assign n1073 = ~n1069 & ~n1072 ;
  assign n1074 = ~n1068 & ~n1073 ;
  assign n1075 = ~n1067 & ~n1074 ;
  assign n1076 = ~n1066 & ~n1075 ;
  assign n1077 = ~n1065 & ~n1076 ;
  assign n1078 = ~n1064 & ~n1077 ;
  assign n1079 = ~n1063 & ~n1078 ;
  assign n1080 = ~n1062 & ~n1079 ;
  assign n1081 = ~n1061 & ~n1080 ;
  assign n1082 = ~n1060 & ~n1081 ;
  assign n1083 = ~n1059 & ~n1082 ;
  assign n1084 = ~n1058 & ~n1083 ;
  assign n1085 = ~n1057 & ~n1084 ;
  assign n1086 = ~n1056 & ~n1085 ;
  assign n1087 = ~n1055 & ~n1086 ;
  assign n1088 = ~n1054 & ~n1087 ;
  assign n1089 = ~n1053 & ~n1088 ;
  assign n1090 = ~n1052 & ~n1089 ;
  assign n1091 = ~n1051 & ~n1090 ;
  assign n1092 = ~n1050 & ~n1091 ;
  assign n1093 = ~n1049 & ~n1092 ;
  assign n1094 = ~n1048 & ~n1093 ;
  assign n1095 = ~n1047 & ~n1094 ;
  assign n1096 = ~n1046 & ~n1095 ;
  assign n1097 = ~n1045 & ~n1096 ;
  assign n1098 = ~n1044 & ~n1097 ;
  assign n1099 = ~n1043 & ~n1098 ;
  assign n1100 = ~n1042 & ~n1099 ;
  assign n1101 = ~n1041 & ~n1100 ;
  assign n1102 = x49 & ~n1101 ;
  assign n1103 = x33 & n1101 ;
  assign n1104 = ~n1102 & ~n1103 ;
  assign n1105 = n1040 & ~n1104 ;
  assign n1106 = x16 & ~n1032 ;
  assign n1107 = x0 & n1032 ;
  assign n1108 = ~n1106 & ~n1107 ;
  assign n1109 = x48 & ~n1101 ;
  assign n1110 = x32 & n1101 ;
  assign n1111 = ~n1109 & ~n1110 ;
  assign n1112 = ~n1108 & n1111 ;
  assign n1113 = ~n1105 & n1112 ;
  assign n1114 = x50 & ~n1101 ;
  assign n1115 = x34 & n1101 ;
  assign n1116 = ~n1114 & ~n1115 ;
  assign n1117 = x18 & ~n1032 ;
  assign n1118 = x2 & n1032 ;
  assign n1119 = ~n1117 & ~n1118 ;
  assign n1120 = n1116 & ~n1119 ;
  assign n1121 = ~n1040 & n1104 ;
  assign n1122 = ~n1120 & ~n1121 ;
  assign n1123 = ~n1113 & n1122 ;
  assign n1124 = x19 & ~n1032 ;
  assign n1125 = x3 & n1032 ;
  assign n1126 = ~n1124 & ~n1125 ;
  assign n1127 = x51 & ~n1101 ;
  assign n1128 = x35 & n1101 ;
  assign n1129 = ~n1127 & ~n1128 ;
  assign n1130 = n1126 & ~n1129 ;
  assign n1131 = ~n1116 & n1119 ;
  assign n1132 = ~n1130 & ~n1131 ;
  assign n1133 = ~n1123 & n1132 ;
  assign n1134 = ~n1126 & n1129 ;
  assign n1135 = x20 & ~n1032 ;
  assign n1136 = x4 & n1032 ;
  assign n1137 = ~n1135 & ~n1136 ;
  assign n1138 = x52 & ~n1101 ;
  assign n1139 = x36 & n1101 ;
  assign n1140 = ~n1138 & ~n1139 ;
  assign n1141 = ~n1137 & n1140 ;
  assign n1142 = ~n1134 & ~n1141 ;
  assign n1143 = ~n1133 & n1142 ;
  assign n1144 = n1137 & ~n1140 ;
  assign n1145 = x53 & ~n1101 ;
  assign n1146 = x37 & n1101 ;
  assign n1147 = ~n1145 & ~n1146 ;
  assign n1148 = x21 & ~n1032 ;
  assign n1149 = x5 & n1032 ;
  assign n1150 = ~n1148 & ~n1149 ;
  assign n1151 = ~n1147 & n1150 ;
  assign n1152 = ~n1144 & ~n1151 ;
  assign n1153 = ~n1143 & n1152 ;
  assign n1154 = n1147 & ~n1150 ;
  assign n1155 = x54 & ~n1101 ;
  assign n1156 = x38 & n1101 ;
  assign n1157 = ~n1155 & ~n1156 ;
  assign n1158 = x22 & ~n1032 ;
  assign n1159 = x6 & n1032 ;
  assign n1160 = ~n1158 & ~n1159 ;
  assign n1161 = n1157 & ~n1160 ;
  assign n1162 = ~n1154 & ~n1161 ;
  assign n1163 = ~n1153 & n1162 ;
  assign n1164 = ~n1157 & n1160 ;
  assign n1165 = x23 & ~n1032 ;
  assign n1166 = x7 & n1032 ;
  assign n1167 = ~n1165 & ~n1166 ;
  assign n1168 = x55 & ~n1101 ;
  assign n1169 = x39 & n1101 ;
  assign n1170 = ~n1168 & ~n1169 ;
  assign n1171 = n1167 & ~n1170 ;
  assign n1172 = ~n1164 & ~n1171 ;
  assign n1173 = ~n1163 & n1172 ;
  assign n1174 = ~n1167 & n1170 ;
  assign n1175 = x56 & ~n1101 ;
  assign n1176 = x40 & n1101 ;
  assign n1177 = ~n1175 & ~n1176 ;
  assign n1178 = ~n1035 & n1177 ;
  assign n1179 = ~n1174 & ~n1178 ;
  assign n1180 = ~n1173 & n1179 ;
  assign n1181 = n1035 & ~n1177 ;
  assign n1182 = x25 & ~n1032 ;
  assign n1183 = x9 & n1032 ;
  assign n1184 = ~n1182 & ~n1183 ;
  assign n1185 = x57 & ~n1101 ;
  assign n1186 = x41 & n1101 ;
  assign n1187 = ~n1185 & ~n1186 ;
  assign n1188 = n1184 & ~n1187 ;
  assign n1189 = ~n1181 & ~n1188 ;
  assign n1190 = ~n1180 & n1189 ;
  assign n1191 = ~n1184 & n1187 ;
  assign n1192 = x58 & ~n1101 ;
  assign n1193 = x42 & n1101 ;
  assign n1194 = ~n1192 & ~n1193 ;
  assign n1195 = x26 & ~n1032 ;
  assign n1196 = x10 & n1032 ;
  assign n1197 = ~n1195 & ~n1196 ;
  assign n1198 = n1194 & ~n1197 ;
  assign n1199 = ~n1191 & ~n1198 ;
  assign n1200 = ~n1190 & n1199 ;
  assign n1201 = x59 & ~n1101 ;
  assign n1202 = x43 & n1101 ;
  assign n1203 = ~n1201 & ~n1202 ;
  assign n1204 = x27 & ~n1032 ;
  assign n1205 = x11 & n1032 ;
  assign n1206 = ~n1204 & ~n1205 ;
  assign n1207 = ~n1203 & n1206 ;
  assign n1208 = ~n1194 & n1197 ;
  assign n1209 = ~n1207 & ~n1208 ;
  assign n1210 = ~n1200 & n1209 ;
  assign n1211 = x60 & ~n1101 ;
  assign n1212 = x44 & n1101 ;
  assign n1213 = ~n1211 & ~n1212 ;
  assign n1214 = x28 & ~n1032 ;
  assign n1215 = x12 & n1032 ;
  assign n1216 = ~n1214 & ~n1215 ;
  assign n1217 = n1213 & ~n1216 ;
  assign n1218 = n1203 & ~n1206 ;
  assign n1219 = ~n1217 & ~n1218 ;
  assign n1220 = ~n1210 & n1219 ;
  assign n1221 = ~n1213 & n1216 ;
  assign n1222 = x61 & ~n1101 ;
  assign n1223 = x45 & n1101 ;
  assign n1224 = ~n1222 & ~n1223 ;
  assign n1225 = x29 & ~n1032 ;
  assign n1226 = x13 & n1032 ;
  assign n1227 = ~n1225 & ~n1226 ;
  assign n1228 = ~n1224 & n1227 ;
  assign n1229 = ~n1221 & ~n1228 ;
  assign n1230 = ~n1220 & n1229 ;
  assign n1231 = n1224 & ~n1227 ;
  assign n1232 = x30 & ~n1032 ;
  assign n1233 = x14 & n1032 ;
  assign n1234 = ~n1232 & ~n1233 ;
  assign n1235 = x62 & ~n1101 ;
  assign n1236 = x46 & n1101 ;
  assign n1237 = ~n1235 & ~n1236 ;
  assign n1238 = ~n1234 & n1237 ;
  assign n1239 = ~n1231 & ~n1238 ;
  assign n1240 = ~n1230 & n1239 ;
  assign n1241 = n1234 & ~n1237 ;
  assign n1242 = ~n1240 & ~n1241 ;
  assign n1243 = ~n1037 & ~n1242 ;
  assign n1244 = ~n1036 & ~n1243 ;
  assign n1245 = ~n1035 & n1244 ;
  assign n1246 = ~n1177 & ~n1244 ;
  assign n1247 = ~n1245 & ~n1246 ;
  assign n1248 = ~n266 & n269 ;
  assign n1249 = ~n1040 & n1244 ;
  assign n1250 = ~n1104 & ~n1244 ;
  assign n1251 = ~n1249 & ~n1250 ;
  assign n1252 = ~x79 & x95 ;
  assign n1253 = x79 & ~x95 ;
  assign n1254 = ~x78 & x94 ;
  assign n1255 = x78 & ~x94 ;
  assign n1256 = ~x77 & x93 ;
  assign n1257 = x77 & ~x93 ;
  assign n1258 = ~x76 & x92 ;
  assign n1259 = x76 & ~x92 ;
  assign n1260 = ~x75 & x91 ;
  assign n1261 = x75 & ~x91 ;
  assign n1262 = ~x74 & x90 ;
  assign n1263 = x74 & ~x90 ;
  assign n1264 = ~x73 & x89 ;
  assign n1265 = x73 & ~x89 ;
  assign n1266 = ~x72 & x88 ;
  assign n1267 = x72 & ~x88 ;
  assign n1268 = ~x71 & x87 ;
  assign n1269 = x71 & ~x87 ;
  assign n1270 = ~x70 & x86 ;
  assign n1271 = x70 & ~x86 ;
  assign n1272 = ~x69 & x85 ;
  assign n1273 = x69 & ~x85 ;
  assign n1274 = ~x68 & x84 ;
  assign n1275 = x68 & ~x84 ;
  assign n1276 = ~x67 & x83 ;
  assign n1277 = x67 & ~x83 ;
  assign n1278 = ~x66 & x82 ;
  assign n1279 = x66 & ~x82 ;
  assign n1280 = ~x65 & x81 ;
  assign n1281 = x65 & ~x81 ;
  assign n1282 = x64 & ~x80 ;
  assign n1283 = ~n1281 & ~n1282 ;
  assign n1284 = ~n1280 & ~n1283 ;
  assign n1285 = ~n1279 & ~n1284 ;
  assign n1286 = ~n1278 & ~n1285 ;
  assign n1287 = ~n1277 & ~n1286 ;
  assign n1288 = ~n1276 & ~n1287 ;
  assign n1289 = ~n1275 & ~n1288 ;
  assign n1290 = ~n1274 & ~n1289 ;
  assign n1291 = ~n1273 & ~n1290 ;
  assign n1292 = ~n1272 & ~n1291 ;
  assign n1293 = ~n1271 & ~n1292 ;
  assign n1294 = ~n1270 & ~n1293 ;
  assign n1295 = ~n1269 & ~n1294 ;
  assign n1296 = ~n1268 & ~n1295 ;
  assign n1297 = ~n1267 & ~n1296 ;
  assign n1298 = ~n1266 & ~n1297 ;
  assign n1299 = ~n1265 & ~n1298 ;
  assign n1300 = ~n1264 & ~n1299 ;
  assign n1301 = ~n1263 & ~n1300 ;
  assign n1302 = ~n1262 & ~n1301 ;
  assign n1303 = ~n1261 & ~n1302 ;
  assign n1304 = ~n1260 & ~n1303 ;
  assign n1305 = ~n1259 & ~n1304 ;
  assign n1306 = ~n1258 & ~n1305 ;
  assign n1307 = ~n1257 & ~n1306 ;
  assign n1308 = ~n1256 & ~n1307 ;
  assign n1309 = ~n1255 & ~n1308 ;
  assign n1310 = ~n1254 & ~n1309 ;
  assign n1311 = ~n1253 & ~n1310 ;
  assign n1312 = ~n1252 & ~n1311 ;
  assign n1313 = x81 & ~n1312 ;
  assign n1314 = x65 & n1312 ;
  assign n1315 = ~n1313 & ~n1314 ;
  assign n1316 = n267 & ~n268 ;
  assign n1317 = ~n267 & n268 ;
  assign n1318 = ~x111 & x127 ;
  assign n1319 = x111 & ~x127 ;
  assign n1320 = ~x110 & x126 ;
  assign n1321 = x110 & ~x126 ;
  assign n1322 = ~x109 & x125 ;
  assign n1323 = x109 & ~x125 ;
  assign n1324 = ~x108 & x124 ;
  assign n1325 = x108 & ~x124 ;
  assign n1326 = ~x107 & x123 ;
  assign n1327 = x107 & ~x123 ;
  assign n1328 = ~x106 & x122 ;
  assign n1329 = x106 & ~x122 ;
  assign n1330 = ~x105 & x121 ;
  assign n1331 = x105 & ~x121 ;
  assign n1332 = ~x104 & x120 ;
  assign n1333 = x104 & ~x120 ;
  assign n1334 = ~x103 & x119 ;
  assign n1335 = x103 & ~x119 ;
  assign n1336 = ~x102 & x118 ;
  assign n1337 = x102 & ~x118 ;
  assign n1338 = ~x101 & x117 ;
  assign n1339 = x101 & ~x117 ;
  assign n1340 = ~x100 & x116 ;
  assign n1341 = x100 & ~x116 ;
  assign n1342 = ~x99 & x115 ;
  assign n1343 = x99 & ~x115 ;
  assign n1344 = ~x98 & x114 ;
  assign n1345 = x98 & ~x114 ;
  assign n1346 = ~x97 & x113 ;
  assign n1347 = x97 & ~x113 ;
  assign n1348 = x96 & ~x112 ;
  assign n1349 = ~n1347 & ~n1348 ;
  assign n1350 = ~n1346 & ~n1349 ;
  assign n1351 = ~n1345 & ~n1350 ;
  assign n1352 = ~n1344 & ~n1351 ;
  assign n1353 = ~n1343 & ~n1352 ;
  assign n1354 = ~n1342 & ~n1353 ;
  assign n1355 = ~n1341 & ~n1354 ;
  assign n1356 = ~n1340 & ~n1355 ;
  assign n1357 = ~n1339 & ~n1356 ;
  assign n1358 = ~n1338 & ~n1357 ;
  assign n1359 = ~n1337 & ~n1358 ;
  assign n1360 = ~n1336 & ~n1359 ;
  assign n1361 = ~n1335 & ~n1360 ;
  assign n1362 = ~n1334 & ~n1361 ;
  assign n1363 = ~n1333 & ~n1362 ;
  assign n1364 = ~n1332 & ~n1363 ;
  assign n1365 = ~n1331 & ~n1364 ;
  assign n1366 = ~n1330 & ~n1365 ;
  assign n1367 = ~n1329 & ~n1366 ;
  assign n1368 = ~n1328 & ~n1367 ;
  assign n1369 = ~n1327 & ~n1368 ;
  assign n1370 = ~n1326 & ~n1369 ;
  assign n1371 = ~n1325 & ~n1370 ;
  assign n1372 = ~n1324 & ~n1371 ;
  assign n1373 = ~n1323 & ~n1372 ;
  assign n1374 = ~n1322 & ~n1373 ;
  assign n1375 = ~n1321 & ~n1374 ;
  assign n1376 = ~n1320 & ~n1375 ;
  assign n1377 = ~n1319 & ~n1376 ;
  assign n1378 = ~n1318 & ~n1377 ;
  assign n1379 = x126 & ~n1378 ;
  assign n1380 = x110 & n1378 ;
  assign n1381 = ~n1379 & ~n1380 ;
  assign n1382 = x94 & ~n1312 ;
  assign n1383 = x78 & n1312 ;
  assign n1384 = ~n1382 & ~n1383 ;
  assign n1385 = ~n1381 & n1384 ;
  assign n1386 = x113 & ~n1378 ;
  assign n1387 = x97 & n1378 ;
  assign n1388 = ~n1386 & ~n1387 ;
  assign n1389 = n1315 & ~n1388 ;
  assign n1390 = x112 & ~n1378 ;
  assign n1391 = x96 & n1378 ;
  assign n1392 = ~n1390 & ~n1391 ;
  assign n1393 = x80 & ~n1312 ;
  assign n1394 = x64 & n1312 ;
  assign n1395 = ~n1393 & ~n1394 ;
  assign n1396 = n1392 & ~n1395 ;
  assign n1397 = ~n1389 & n1396 ;
  assign n1398 = x114 & ~n1378 ;
  assign n1399 = x98 & n1378 ;
  assign n1400 = ~n1398 & ~n1399 ;
  assign n1401 = x82 & ~n1312 ;
  assign n1402 = x66 & n1312 ;
  assign n1403 = ~n1401 & ~n1402 ;
  assign n1404 = n1400 & ~n1403 ;
  assign n1405 = ~n1315 & n1388 ;
  assign n1406 = ~n1404 & ~n1405 ;
  assign n1407 = ~n1397 & n1406 ;
  assign n1408 = x115 & ~n1378 ;
  assign n1409 = x99 & n1378 ;
  assign n1410 = ~n1408 & ~n1409 ;
  assign n1411 = x83 & ~n1312 ;
  assign n1412 = x67 & n1312 ;
  assign n1413 = ~n1411 & ~n1412 ;
  assign n1414 = ~n1410 & n1413 ;
  assign n1415 = ~n1400 & n1403 ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = ~n1407 & n1416 ;
  assign n1418 = x116 & ~n1378 ;
  assign n1419 = x100 & n1378 ;
  assign n1420 = ~n1418 & ~n1419 ;
  assign n1421 = x84 & ~n1312 ;
  assign n1422 = x68 & n1312 ;
  assign n1423 = ~n1421 & ~n1422 ;
  assign n1424 = n1420 & ~n1423 ;
  assign n1425 = n1410 & ~n1413 ;
  assign n1426 = ~n1424 & ~n1425 ;
  assign n1427 = ~n1417 & n1426 ;
  assign n1428 = x117 & ~n1378 ;
  assign n1429 = x101 & n1378 ;
  assign n1430 = ~n1428 & ~n1429 ;
  assign n1431 = x85 & ~n1312 ;
  assign n1432 = x69 & n1312 ;
  assign n1433 = ~n1431 & ~n1432 ;
  assign n1434 = ~n1430 & n1433 ;
  assign n1435 = ~n1420 & n1423 ;
  assign n1436 = ~n1434 & ~n1435 ;
  assign n1437 = ~n1427 & n1436 ;
  assign n1438 = n1430 & ~n1433 ;
  assign n1439 = x86 & ~n1312 ;
  assign n1440 = x70 & n1312 ;
  assign n1441 = ~n1439 & ~n1440 ;
  assign n1442 = x118 & ~n1378 ;
  assign n1443 = x102 & n1378 ;
  assign n1444 = ~n1442 & ~n1443 ;
  assign n1445 = ~n1441 & n1444 ;
  assign n1446 = ~n1438 & ~n1445 ;
  assign n1447 = ~n1437 & n1446 ;
  assign n1448 = x87 & ~n1312 ;
  assign n1449 = x71 & n1312 ;
  assign n1450 = ~n1448 & ~n1449 ;
  assign n1451 = x119 & ~n1378 ;
  assign n1452 = x103 & n1378 ;
  assign n1453 = ~n1451 & ~n1452 ;
  assign n1454 = n1450 & ~n1453 ;
  assign n1455 = n1441 & ~n1444 ;
  assign n1456 = ~n1454 & ~n1455 ;
  assign n1457 = ~n1447 & n1456 ;
  assign n1458 = ~n1450 & n1453 ;
  assign n1459 = x120 & ~n1378 ;
  assign n1460 = x104 & n1378 ;
  assign n1461 = ~n1459 & ~n1460 ;
  assign n1462 = x88 & ~n1312 ;
  assign n1463 = x72 & n1312 ;
  assign n1464 = ~n1462 & ~n1463 ;
  assign n1465 = n1461 & ~n1464 ;
  assign n1466 = ~n1458 & ~n1465 ;
  assign n1467 = ~n1457 & n1466 ;
  assign n1468 = ~n1461 & n1464 ;
  assign n1469 = x121 & ~n1378 ;
  assign n1470 = x105 & n1378 ;
  assign n1471 = ~n1469 & ~n1470 ;
  assign n1472 = x89 & ~n1312 ;
  assign n1473 = x73 & n1312 ;
  assign n1474 = ~n1472 & ~n1473 ;
  assign n1475 = ~n1471 & n1474 ;
  assign n1476 = ~n1468 & ~n1475 ;
  assign n1477 = ~n1467 & n1476 ;
  assign n1478 = n1471 & ~n1474 ;
  assign n1479 = x90 & ~n1312 ;
  assign n1480 = x74 & n1312 ;
  assign n1481 = ~n1479 & ~n1480 ;
  assign n1482 = x122 & ~n1378 ;
  assign n1483 = x106 & n1378 ;
  assign n1484 = ~n1482 & ~n1483 ;
  assign n1485 = ~n1481 & n1484 ;
  assign n1486 = ~n1478 & ~n1485 ;
  assign n1487 = ~n1477 & n1486 ;
  assign n1488 = x91 & ~n1312 ;
  assign n1489 = x75 & n1312 ;
  assign n1490 = ~n1488 & ~n1489 ;
  assign n1491 = x123 & ~n1378 ;
  assign n1492 = x107 & n1378 ;
  assign n1493 = ~n1491 & ~n1492 ;
  assign n1494 = n1490 & ~n1493 ;
  assign n1495 = n1481 & ~n1484 ;
  assign n1496 = ~n1494 & ~n1495 ;
  assign n1497 = ~n1487 & n1496 ;
  assign n1498 = x124 & ~n1378 ;
  assign n1499 = x108 & n1378 ;
  assign n1500 = ~n1498 & ~n1499 ;
  assign n1501 = x92 & ~n1312 ;
  assign n1502 = x76 & n1312 ;
  assign n1503 = ~n1501 & ~n1502 ;
  assign n1504 = n1500 & ~n1503 ;
  assign n1505 = ~n1490 & n1493 ;
  assign n1506 = ~n1504 & ~n1505 ;
  assign n1507 = ~n1497 & n1506 ;
  assign n1508 = ~n1500 & n1503 ;
  assign n1509 = x125 & ~n1378 ;
  assign n1510 = x109 & n1378 ;
  assign n1511 = ~n1509 & ~n1510 ;
  assign n1512 = x93 & ~n1312 ;
  assign n1513 = x77 & n1312 ;
  assign n1514 = ~n1512 & ~n1513 ;
  assign n1515 = ~n1511 & n1514 ;
  assign n1516 = ~n1508 & ~n1515 ;
  assign n1517 = ~n1507 & n1516 ;
  assign n1518 = n1381 & ~n1384 ;
  assign n1519 = n1511 & ~n1514 ;
  assign n1520 = ~n1518 & ~n1519 ;
  assign n1521 = ~n1517 & n1520 ;
  assign n1522 = ~n1385 & ~n1521 ;
  assign n1523 = ~n1317 & ~n1522 ;
  assign n1524 = ~n1316 & ~n1523 ;
  assign n1525 = ~n1315 & n1524 ;
  assign n1526 = ~n1388 & ~n1524 ;
  assign n1527 = ~n1525 & ~n1526 ;
  assign n1528 = n1251 & ~n1527 ;
  assign n1529 = ~n1395 & n1524 ;
  assign n1530 = ~n1392 & ~n1524 ;
  assign n1531 = ~n1529 & ~n1530 ;
  assign n1532 = ~n1108 & n1244 ;
  assign n1533 = ~n1111 & ~n1244 ;
  assign n1534 = ~n1532 & ~n1533 ;
  assign n1535 = n1531 & ~n1534 ;
  assign n1536 = ~n1528 & n1535 ;
  assign n1537 = ~n1403 & n1524 ;
  assign n1538 = ~n1400 & ~n1524 ;
  assign n1539 = ~n1537 & ~n1538 ;
  assign n1540 = ~n1119 & n1244 ;
  assign n1541 = ~n1116 & ~n1244 ;
  assign n1542 = ~n1540 & ~n1541 ;
  assign n1543 = n1539 & ~n1542 ;
  assign n1544 = ~n1251 & n1527 ;
  assign n1545 = ~n1543 & ~n1544 ;
  assign n1546 = ~n1536 & n1545 ;
  assign n1547 = ~n1539 & n1542 ;
  assign n1548 = ~n1126 & n1244 ;
  assign n1549 = ~n1129 & ~n1244 ;
  assign n1550 = ~n1548 & ~n1549 ;
  assign n1551 = n1410 & ~n1524 ;
  assign n1552 = n1413 & n1524 ;
  assign n1553 = ~n1551 & ~n1552 ;
  assign n1554 = n1550 & n1553 ;
  assign n1555 = ~n1547 & ~n1554 ;
  assign n1556 = ~n1546 & n1555 ;
  assign n1557 = ~n1137 & n1244 ;
  assign n1558 = ~n1140 & ~n1244 ;
  assign n1559 = ~n1557 & ~n1558 ;
  assign n1560 = ~n1423 & n1524 ;
  assign n1561 = ~n1420 & ~n1524 ;
  assign n1562 = ~n1560 & ~n1561 ;
  assign n1563 = ~n1559 & n1562 ;
  assign n1564 = ~n1550 & ~n1553 ;
  assign n1565 = ~n1563 & ~n1564 ;
  assign n1566 = ~n1556 & n1565 ;
  assign n1567 = ~n1150 & n1244 ;
  assign n1568 = ~n1147 & ~n1244 ;
  assign n1569 = ~n1567 & ~n1568 ;
  assign n1570 = ~n1433 & n1524 ;
  assign n1571 = ~n1430 & ~n1524 ;
  assign n1572 = ~n1570 & ~n1571 ;
  assign n1573 = n1569 & ~n1572 ;
  assign n1574 = n1559 & ~n1562 ;
  assign n1575 = ~n1573 & ~n1574 ;
  assign n1576 = ~n1566 & n1575 ;
  assign n1577 = ~n1441 & n1524 ;
  assign n1578 = ~n1444 & ~n1524 ;
  assign n1579 = ~n1577 & ~n1578 ;
  assign n1580 = ~n1160 & n1244 ;
  assign n1581 = ~n1157 & ~n1244 ;
  assign n1582 = ~n1580 & ~n1581 ;
  assign n1583 = n1579 & ~n1582 ;
  assign n1584 = ~n1569 & n1572 ;
  assign n1585 = ~n1583 & ~n1584 ;
  assign n1586 = ~n1576 & n1585 ;
  assign n1587 = ~n1167 & n1244 ;
  assign n1588 = ~n1170 & ~n1244 ;
  assign n1589 = ~n1587 & ~n1588 ;
  assign n1590 = ~n1450 & n1524 ;
  assign n1591 = ~n1453 & ~n1524 ;
  assign n1592 = ~n1590 & ~n1591 ;
  assign n1593 = n1589 & ~n1592 ;
  assign n1594 = ~n1579 & n1582 ;
  assign n1595 = ~n1593 & ~n1594 ;
  assign n1596 = ~n1586 & n1595 ;
  assign n1597 = ~n1464 & n1524 ;
  assign n1598 = ~n1461 & ~n1524 ;
  assign n1599 = ~n1597 & ~n1598 ;
  assign n1600 = ~n1247 & n1599 ;
  assign n1601 = ~n1589 & n1592 ;
  assign n1602 = ~n1600 & ~n1601 ;
  assign n1603 = ~n1596 & n1602 ;
  assign n1604 = ~n1184 & n1244 ;
  assign n1605 = ~n1187 & ~n1244 ;
  assign n1606 = ~n1604 & ~n1605 ;
  assign n1607 = ~n1474 & n1524 ;
  assign n1608 = ~n1471 & ~n1524 ;
  assign n1609 = ~n1607 & ~n1608 ;
  assign n1610 = n1606 & ~n1609 ;
  assign n1611 = n1247 & ~n1599 ;
  assign n1612 = ~n1610 & ~n1611 ;
  assign n1613 = ~n1603 & n1612 ;
  assign n1614 = ~n1481 & n1524 ;
  assign n1615 = ~n1484 & ~n1524 ;
  assign n1616 = ~n1614 & ~n1615 ;
  assign n1617 = n1194 & ~n1244 ;
  assign n1618 = n1197 & n1244 ;
  assign n1619 = ~n1617 & ~n1618 ;
  assign n1620 = n1616 & n1619 ;
  assign n1621 = ~n1606 & n1609 ;
  assign n1622 = ~n1620 & ~n1621 ;
  assign n1623 = ~n1613 & n1622 ;
  assign n1624 = ~n1616 & ~n1619 ;
  assign n1625 = ~n1490 & n1524 ;
  assign n1626 = ~n1493 & ~n1524 ;
  assign n1627 = ~n1625 & ~n1626 ;
  assign n1628 = ~n1206 & n1244 ;
  assign n1629 = ~n1203 & ~n1244 ;
  assign n1630 = ~n1628 & ~n1629 ;
  assign n1631 = ~n1627 & n1630 ;
  assign n1632 = ~n1624 & ~n1631 ;
  assign n1633 = ~n1623 & n1632 ;
  assign n1634 = n1627 & ~n1630 ;
  assign n1635 = ~n1216 & n1244 ;
  assign n1636 = ~n1213 & ~n1244 ;
  assign n1637 = ~n1635 & ~n1636 ;
  assign n1638 = ~n1503 & n1524 ;
  assign n1639 = ~n1500 & ~n1524 ;
  assign n1640 = ~n1638 & ~n1639 ;
  assign n1641 = ~n1637 & n1640 ;
  assign n1642 = ~n1634 & ~n1641 ;
  assign n1643 = ~n1633 & n1642 ;
  assign n1644 = n1637 & ~n1640 ;
  assign n1645 = ~n1227 & n1244 ;
  assign n1646 = ~n1224 & ~n1244 ;
  assign n1647 = ~n1645 & ~n1646 ;
  assign n1648 = ~n1514 & n1524 ;
  assign n1649 = ~n1511 & ~n1524 ;
  assign n1650 = ~n1648 & ~n1649 ;
  assign n1651 = n1647 & ~n1650 ;
  assign n1652 = ~n1644 & ~n1651 ;
  assign n1653 = ~n1643 & n1652 ;
  assign n1654 = ~n1647 & n1650 ;
  assign n1655 = ~n1234 & n1244 ;
  assign n1656 = ~n1237 & ~n1244 ;
  assign n1657 = ~n1655 & ~n1656 ;
  assign n1658 = ~n1384 & n1524 ;
  assign n1659 = ~n1381 & ~n1524 ;
  assign n1660 = ~n1658 & ~n1659 ;
  assign n1661 = ~n1657 & n1660 ;
  assign n1662 = ~n1654 & ~n1661 ;
  assign n1663 = ~n1653 & n1662 ;
  assign n1664 = n266 & ~n269 ;
  assign n1665 = n1657 & ~n1660 ;
  assign n1666 = ~n1664 & ~n1665 ;
  assign n1667 = ~n1663 & n1666 ;
  assign n1668 = ~n1248 & ~n1667 ;
  assign n1669 = ~n1247 & ~n1668 ;
  assign n1670 = ~n1599 & n1668 ;
  assign n1671 = ~n1669 & ~n1670 ;
  assign n1672 = n971 & ~n1671 ;
  assign n1673 = ~n1589 & ~n1668 ;
  assign n1674 = ~n1592 & n1668 ;
  assign n1675 = ~n1673 & ~n1674 ;
  assign n1676 = ~n889 & ~n968 ;
  assign n1677 = ~n892 & n968 ;
  assign n1678 = ~n1676 & ~n1677 ;
  assign n1679 = n1675 & ~n1678 ;
  assign n1680 = ~n1675 & n1678 ;
  assign n1681 = ~n882 & ~n968 ;
  assign n1682 = ~n879 & n968 ;
  assign n1683 = ~n1681 & ~n1682 ;
  assign n1684 = ~n1582 & ~n1668 ;
  assign n1685 = ~n1579 & n1668 ;
  assign n1686 = ~n1684 & ~n1685 ;
  assign n1687 = ~n1683 & n1686 ;
  assign n1688 = n1683 & ~n1686 ;
  assign n1689 = ~n1569 & ~n1668 ;
  assign n1690 = ~n1572 & n1668 ;
  assign n1691 = ~n1689 & ~n1690 ;
  assign n1692 = ~n869 & ~n968 ;
  assign n1693 = ~n872 & n968 ;
  assign n1694 = ~n1692 & ~n1693 ;
  assign n1695 = n1691 & ~n1694 ;
  assign n1696 = ~n1691 & n1694 ;
  assign n1697 = ~n862 & ~n968 ;
  assign n1698 = ~n859 & n968 ;
  assign n1699 = ~n1697 & ~n1698 ;
  assign n1700 = ~n1562 & n1668 ;
  assign n1701 = ~n1559 & ~n1668 ;
  assign n1702 = ~n1700 & ~n1701 ;
  assign n1703 = ~n1699 & n1702 ;
  assign n1704 = ~n1251 & ~n1668 ;
  assign n1705 = ~n1527 & n1668 ;
  assign n1706 = ~n1704 & ~n1705 ;
  assign n1707 = ~n827 & n968 ;
  assign n1708 = ~n551 & ~n968 ;
  assign n1709 = ~n1707 & ~n1708 ;
  assign n1710 = n1706 & ~n1709 ;
  assign n1711 = ~n834 & ~n968 ;
  assign n1712 = ~n831 & n968 ;
  assign n1713 = ~n1711 & ~n1712 ;
  assign n1714 = ~n1534 & ~n1668 ;
  assign n1715 = ~n1531 & n1668 ;
  assign n1716 = ~n1714 & ~n1715 ;
  assign n1717 = n1713 & ~n1716 ;
  assign n1718 = ~n1710 & n1717 ;
  assign n1719 = ~n842 & ~n968 ;
  assign n1720 = ~n839 & n968 ;
  assign n1721 = ~n1719 & ~n1720 ;
  assign n1722 = ~n1542 & ~n1668 ;
  assign n1723 = ~n1539 & n1668 ;
  assign n1724 = ~n1722 & ~n1723 ;
  assign n1725 = n1721 & ~n1724 ;
  assign n1726 = ~n1706 & n1709 ;
  assign n1727 = ~n1725 & ~n1726 ;
  assign n1728 = ~n1718 & n1727 ;
  assign n1729 = n853 & ~n968 ;
  assign n1730 = n850 & n968 ;
  assign n1731 = ~n1729 & ~n1730 ;
  assign n1732 = ~n1550 & ~n1668 ;
  assign n1733 = n1553 & n1668 ;
  assign n1734 = ~n1732 & ~n1733 ;
  assign n1735 = n1731 & n1734 ;
  assign n1736 = ~n1721 & n1724 ;
  assign n1737 = ~n1735 & ~n1736 ;
  assign n1738 = ~n1728 & n1737 ;
  assign n1739 = n1699 & ~n1702 ;
  assign n1740 = ~n1731 & ~n1734 ;
  assign n1741 = ~n1739 & ~n1740 ;
  assign n1742 = ~n1738 & n1741 ;
  assign n1743 = ~n1703 & ~n1742 ;
  assign n1744 = ~n1696 & ~n1743 ;
  assign n1745 = ~n1695 & ~n1744 ;
  assign n1746 = ~n1688 & ~n1745 ;
  assign n1747 = ~n1687 & ~n1746 ;
  assign n1748 = ~n1680 & ~n1747 ;
  assign n1749 = ~n1679 & ~n1748 ;
  assign n1750 = ~n1672 & ~n1749 ;
  assign n1751 = ~n971 & n1671 ;
  assign n1752 = ~n1606 & ~n1668 ;
  assign n1753 = ~n1609 & n1668 ;
  assign n1754 = ~n1752 & ~n1753 ;
  assign n1755 = n906 & ~n968 ;
  assign n1756 = ~n909 & n968 ;
  assign n1757 = ~n1755 & ~n1756 ;
  assign n1758 = n1754 & ~n1757 ;
  assign n1759 = ~n1751 & ~n1758 ;
  assign n1760 = ~n1750 & n1759 ;
  assign n1761 = ~n1754 & n1757 ;
  assign n1762 = n919 & ~n968 ;
  assign n1763 = n916 & n968 ;
  assign n1764 = ~n1762 & ~n1763 ;
  assign n1765 = n1619 & ~n1668 ;
  assign n1766 = ~n1616 & n1668 ;
  assign n1767 = ~n1765 & ~n1766 ;
  assign n1768 = ~n1764 & ~n1767 ;
  assign n1769 = ~n1761 & ~n1768 ;
  assign n1770 = ~n1760 & n1769 ;
  assign n1771 = n1764 & n1767 ;
  assign n1772 = n1630 & ~n1668 ;
  assign n1773 = n1627 & n1668 ;
  assign n1774 = ~n1772 & ~n1773 ;
  assign n1775 = n930 & ~n968 ;
  assign n1776 = n927 & n968 ;
  assign n1777 = ~n1775 & ~n1776 ;
  assign n1778 = ~n1774 & n1777 ;
  assign n1779 = ~n1771 & ~n1778 ;
  assign n1780 = ~n1770 & n1779 ;
  assign n1781 = n1774 & ~n1777 ;
  assign n1782 = ~n937 & ~n968 ;
  assign n1783 = ~n940 & n968 ;
  assign n1784 = ~n1782 & ~n1783 ;
  assign n1785 = ~n1637 & ~n1668 ;
  assign n1786 = ~n1640 & n1668 ;
  assign n1787 = ~n1785 & ~n1786 ;
  assign n1788 = n1784 & ~n1787 ;
  assign n1789 = ~n1781 & ~n1788 ;
  assign n1790 = ~n1780 & n1789 ;
  assign n1791 = ~n1784 & n1787 ;
  assign n1792 = ~n1647 & ~n1668 ;
  assign n1793 = ~n1650 & n1668 ;
  assign n1794 = ~n1792 & ~n1793 ;
  assign n1795 = ~n947 & ~n968 ;
  assign n1796 = ~n950 & n968 ;
  assign n1797 = ~n1795 & ~n1796 ;
  assign n1798 = n1794 & ~n1797 ;
  assign n1799 = ~n1791 & ~n1798 ;
  assign n1800 = ~n1790 & n1799 ;
  assign n1801 = ~n1794 & n1797 ;
  assign n1802 = ~n960 & n968 ;
  assign n1803 = ~n957 & ~n968 ;
  assign n1804 = ~n1802 & ~n1803 ;
  assign n1805 = ~n1660 & n1668 ;
  assign n1806 = ~n1657 & ~n1668 ;
  assign n1807 = ~n1805 & ~n1806 ;
  assign n1808 = n1804 & ~n1807 ;
  assign n1809 = ~n1801 & ~n1808 ;
  assign n1810 = ~n1800 & n1809 ;
  assign n1811 = ~n263 & n270 ;
  assign n1812 = ~n1804 & n1807 ;
  assign n1813 = ~n1811 & ~n1812 ;
  assign n1814 = ~n1810 & n1813 ;
  assign n1815 = ~n271 & ~n1814 ;
  assign n1816 = n1668 & ~n1815 ;
  assign n1817 = n968 & n1815 ;
  assign n1818 = ~n1816 & ~n1817 ;
  assign n1819 = ~n544 & n1818 ;
  assign n1820 = ~n824 & n968 ;
  assign n1821 = ~n1819 & ~n1820 ;
  assign n1822 = n1815 & ~n1821 ;
  assign n1823 = ~n1244 & n1818 ;
  assign n1824 = ~n1524 & n1668 ;
  assign n1825 = ~n1823 & ~n1824 ;
  assign n1826 = ~n1815 & ~n1825 ;
  assign n1827 = ~n1822 & ~n1826 ;
  assign n1828 = n332 & n1827 ;
  assign n1829 = n401 & ~n1827 ;
  assign n1830 = n1818 & ~n1829 ;
  assign n1831 = ~n1828 & n1830 ;
  assign n1832 = n612 & n1827 ;
  assign n1833 = n678 & ~n1827 ;
  assign n1834 = ~n1818 & ~n1833 ;
  assign n1835 = ~n1832 & n1834 ;
  assign n1836 = ~n1831 & ~n1835 ;
  assign n1837 = n1815 & ~n1836 ;
  assign n1838 = n1032 & n1827 ;
  assign n1839 = n1101 & ~n1827 ;
  assign n1840 = n1818 & ~n1839 ;
  assign n1841 = ~n1838 & n1840 ;
  assign n1842 = n1312 & n1827 ;
  assign n1843 = n1378 & ~n1827 ;
  assign n1844 = ~n1818 & ~n1843 ;
  assign n1845 = ~n1842 & n1844 ;
  assign n1846 = ~n1841 & ~n1845 ;
  assign n1847 = ~n1815 & ~n1846 ;
  assign n1848 = ~n1837 & ~n1847 ;
  assign n1849 = ~n1713 & n1815 ;
  assign n1850 = ~n1716 & ~n1815 ;
  assign n1851 = ~n1849 & ~n1850 ;
  assign n1852 = n1706 & ~n1815 ;
  assign n1853 = n1709 & n1815 ;
  assign n1854 = ~n1852 & ~n1853 ;
  assign n1855 = ~n1721 & n1815 ;
  assign n1856 = ~n1724 & ~n1815 ;
  assign n1857 = ~n1855 & ~n1856 ;
  assign n1858 = ~n1734 & ~n1815 ;
  assign n1859 = n1731 & n1815 ;
  assign n1860 = ~n1858 & ~n1859 ;
  assign n1861 = ~n1699 & n1815 ;
  assign n1862 = ~n1702 & ~n1815 ;
  assign n1863 = ~n1861 & ~n1862 ;
  assign n1864 = ~n1694 & n1815 ;
  assign n1865 = ~n1691 & ~n1815 ;
  assign n1866 = ~n1864 & ~n1865 ;
  assign n1867 = ~n1683 & n1815 ;
  assign n1868 = ~n1686 & ~n1815 ;
  assign n1869 = ~n1867 & ~n1868 ;
  assign n1870 = ~n1678 & n1815 ;
  assign n1871 = ~n1675 & ~n1815 ;
  assign n1872 = ~n1870 & ~n1871 ;
  assign n1873 = ~n971 & n1815 ;
  assign n1874 = ~n1671 & ~n1815 ;
  assign n1875 = ~n1873 & ~n1874 ;
  assign n1876 = ~n1757 & n1815 ;
  assign n1877 = ~n1754 & ~n1815 ;
  assign n1878 = ~n1876 & ~n1877 ;
  assign n1879 = ~n1767 & ~n1815 ;
  assign n1880 = n1764 & n1815 ;
  assign n1881 = ~n1879 & ~n1880 ;
  assign n1882 = n1774 & ~n1815 ;
  assign n1883 = n1777 & n1815 ;
  assign n1884 = ~n1882 & ~n1883 ;
  assign n1885 = ~n1784 & n1815 ;
  assign n1886 = ~n1787 & ~n1815 ;
  assign n1887 = ~n1885 & ~n1886 ;
  assign n1888 = ~n1797 & n1815 ;
  assign n1889 = ~n1794 & ~n1815 ;
  assign n1890 = ~n1888 & ~n1889 ;
  assign n1891 = ~n1804 & n1815 ;
  assign n1892 = ~n1807 & ~n1815 ;
  assign n1893 = ~n1891 & ~n1892 ;
  assign n1894 = n263 & n270 ;
  assign y0 = ~n1848 ;
  assign y1 = ~n1827 ;
  assign y2 = ~n1818 ;
  assign y3 = n1815 ;
  assign y4 = ~n1851 ;
  assign y5 = n1854 ;
  assign y6 = ~n1857 ;
  assign y7 = ~n1860 ;
  assign y8 = ~n1863 ;
  assign y9 = ~n1866 ;
  assign y10 = ~n1869 ;
  assign y11 = ~n1872 ;
  assign y12 = ~n1875 ;
  assign y13 = ~n1878 ;
  assign y14 = ~n1881 ;
  assign y15 = ~n1884 ;
  assign y16 = ~n1887 ;
  assign y17 = ~n1890 ;
  assign y18 = ~n1893 ;
  assign y19 = ~n1894 ;
endmodule
