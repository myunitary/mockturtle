module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 ;
  assign n33 = ~x0 & ~x1 ;
  assign n34 = ~x2 & ~x3 ;
  assign n35 = ~x4 & ~x5 ;
  assign n36 = n34 & n35 ;
  assign n37 = n33 & n36 ;
  assign n38 = ~x10 & ~x11 ;
  assign n39 = ~x13 & ~x14 ;
  assign n40 = n38 & n39 ;
  assign n41 = ~x6 & ~x7 ;
  assign n42 = ~x8 & ~x9 ;
  assign n43 = n41 & n42 ;
  assign n44 = n40 & n43 ;
  assign n45 = n37 & n44 ;
  assign n46 = ~x16 & ~x17 ;
  assign n47 = ~x18 & n46 ;
  assign n48 = ~x12 & ~x15 ;
  assign n49 = ~x19 & n48 ;
  assign n50 = n47 & n49 ;
  assign n51 = ~x21 & ~x22 ;
  assign n52 = ~x20 & ~x23 ;
  assign n53 = n51 & n52 ;
  assign n54 = ~x24 & ~x25 ;
  assign n55 = n53 & n54 ;
  assign n56 = n50 & n55 ;
  assign n57 = n45 & n56 ;
  assign n58 = ~x28 & ~x29 ;
  assign n59 = ~x30 & ~x31 ;
  assign n60 = n58 & n59 ;
  assign n64 = ~x26 & ~x27 ;
  assign n65 = n60 & n64 ;
  assign n66 = ~n57 & ~n65 ;
  assign n61 = x26 & ~x27 ;
  assign n62 = n60 & n61 ;
  assign n63 = n57 & ~n62 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n47 & n48 ;
  assign n69 = x24 & ~x25 ;
  assign n70 = ~x19 & n69 ;
  assign n71 = n53 & n70 ;
  assign n72 = n68 & n71 ;
  assign n73 = n45 & n72 ;
  assign n74 = ~x19 & n54 ;
  assign n75 = n53 & n74 ;
  assign n76 = n68 & n75 ;
  assign n77 = n45 & n76 ;
  assign n78 = n77 ^ n54 ;
  assign n79 = ~n73 & ~n78 ;
  assign n80 = ~n67 & ~n79 ;
  assign n81 = n33 & n48 ;
  assign n82 = n36 & n81 ;
  assign n83 = n44 & n82 ;
  assign n84 = x18 & n46 ;
  assign n85 = n83 & n84 ;
  assign n86 = n85 ^ x18 ;
  assign n87 = ~x19 & n53 ;
  assign n91 = ~n86 & n87 ;
  assign n88 = n68 & n87 ;
  assign n89 = n45 & n88 ;
  assign n90 = ~n86 & n89 ;
  assign n92 = n91 ^ n90 ;
  assign n93 = n83 ^ x16 ;
  assign n94 = ~x17 & ~n93 ;
  assign n95 = n92 & n94 ;
  assign n96 = n80 & n95 ;
  assign n115 = n92 & ~n93 ;
  assign n116 = n80 & n115 ;
  assign n122 = ~x17 & n116 ;
  assign n97 = ~n57 & n65 ;
  assign n98 = ~x24 & x25 ;
  assign n99 = n53 & n98 ;
  assign n100 = n50 & n99 ;
  assign n101 = n45 & n100 ;
  assign n102 = n101 ^ x25 ;
  assign n103 = n97 & ~n102 ;
  assign n104 = n45 & n68 ;
  assign n105 = x19 & ~n104 ;
  assign n106 = n45 & n50 ;
  assign n107 = ~x24 & n53 ;
  assign n108 = ~n106 & n107 ;
  assign n109 = ~n105 & n108 ;
  assign n110 = n103 & n109 ;
  assign n111 = ~x16 & n83 ;
  assign n117 = x17 & ~x18 ;
  assign n118 = n111 & n117 ;
  assign n119 = ~n116 & n118 ;
  assign n120 = n110 & n119 ;
  assign n112 = ~x17 & ~x18 ;
  assign n113 = ~n111 & n112 ;
  assign n114 = n110 & n113 ;
  assign n121 = n120 ^ n114 ;
  assign n123 = n122 ^ n121 ;
  assign n129 = n80 & n92 ;
  assign n124 = n46 & n83 ;
  assign n125 = ~x18 & ~n124 ;
  assign n126 = x17 & ~n111 ;
  assign n127 = n125 & ~n126 ;
  assign n128 = n110 & n127 ;
  assign n130 = n129 ^ n128 ;
  assign n131 = ~n96 & n130 ;
  assign n132 = n110 & n129 ;
  assign n134 = ~n110 & n129 ;
  assign n133 = n110 & ~n127 ;
  assign n135 = n134 ^ n133 ;
  assign n136 = n132 & n135 ;
  assign n137 = n136 ^ n135 ;
  assign n138 = ~x23 & n51 ;
  assign n141 = ~x20 & n138 ;
  assign n139 = n50 & n138 ;
  assign n140 = n45 & n139 ;
  assign n142 = n141 ^ n140 ;
  assign n146 = n80 & n142 ;
  assign n143 = n92 & n142 ;
  assign n144 = n80 & n143 ;
  assign n145 = ~n110 & n144 ;
  assign n147 = n146 ^ n145 ;
  assign n148 = n147 ^ n110 ;
  assign n149 = n110 & ~n146 ;
  assign n150 = ~x20 & n50 ;
  assign n151 = n45 & n150 ;
  assign n152 = n151 ^ x21 ;
  assign n153 = ~x22 & ~x23 ;
  assign n154 = ~x24 & n153 ;
  assign n155 = ~n102 & n154 ;
  assign n156 = n97 & n155 ;
  assign n157 = ~n152 & n156 ;
  assign n158 = n149 & n157 ;
  assign n159 = n158 ^ n157 ;
  assign n160 = n159 ^ n146 ;
  assign n165 = ~x24 & ~n152 ;
  assign n161 = n79 & ~n152 ;
  assign n162 = ~x24 & ~n102 ;
  assign n163 = n97 & n162 ;
  assign n164 = n161 & n163 ;
  assign n166 = n165 ^ n164 ;
  assign n167 = ~n146 & ~n166 ;
  assign n168 = ~x20 & ~x21 ;
  assign n169 = n50 & n168 ;
  assign n170 = n45 & n169 ;
  assign n171 = ~x23 & n170 ;
  assign n172 = n171 ^ n153 ;
  assign n180 = n80 & n172 ;
  assign n176 = ~x21 & ~x24 ;
  assign n177 = n172 & n176 ;
  assign n178 = ~n80 & n177 ;
  assign n173 = ~x24 & n151 ;
  assign n174 = n172 & n173 ;
  assign n175 = ~n80 & n174 ;
  assign n179 = n178 ^ n175 ;
  assign n181 = n180 ^ n179 ;
  assign n182 = n167 & n181 ;
  assign n183 = ~x22 & n170 ;
  assign n184 = x23 & ~n183 ;
  assign n185 = ~x24 & ~n89 ;
  assign n186 = n103 & n185 ;
  assign n187 = ~n184 & n186 ;
  assign n188 = ~n172 & n187 ;
  assign n189 = n80 & ~n187 ;
  assign n190 = n79 & n103 ;
  assign n191 = ~n67 & n79 ;
  assign n192 = ~n103 & n191 ;
  assign n193 = ~x26 & n33 ;
  assign n194 = n36 & n193 ;
  assign n195 = n44 & n194 ;
  assign n196 = n56 & n195 ;
  assign n197 = ~n61 & ~n196 ;
  assign n198 = ~x27 & n57 ;
  assign n199 = n60 & ~n198 ;
  assign n200 = ~n197 & n199 ;
  assign n201 = x27 & ~x28 ;
  assign n202 = ~n196 & n201 ;
  assign n203 = ~x27 & n196 ;
  assign n204 = x28 & n203 ;
  assign n205 = ~n202 & ~n204 ;
  assign n206 = ~x29 & n59 ;
  assign n207 = ~n205 & n206 ;
  assign n208 = x29 & ~n203 ;
  assign n209 = ~n58 & n59 ;
  assign n210 = ~n204 & n209 ;
  assign n211 = ~n208 & n210 ;
  assign n212 = ~x27 & ~x28 ;
  assign n213 = n196 & n212 ;
  assign n217 = x29 & n59 ;
  assign n218 = ~n213 & n217 ;
  assign n214 = x30 & ~x31 ;
  assign n215 = ~x29 & n214 ;
  assign n216 = n213 & n215 ;
  assign n219 = n218 ^ n216 ;
  assign n220 = ~x29 & ~n214 ;
  assign n221 = n212 & n220 ;
  assign n222 = n196 & n221 ;
  assign n223 = n222 ^ n214 ;
  assign n224 = ~x30 & x31 ;
  assign n225 = ~x29 & ~n224 ;
  assign n226 = n212 & n225 ;
  assign n227 = n196 & n226 ;
  assign n228 = n223 & ~n227 ;
  assign y0 = n96 ;
  assign y1 = n123 ;
  assign y2 = n131 ;
  assign y3 = n137 ;
  assign y4 = n148 ;
  assign y5 = n160 ;
  assign y6 = n182 ;
  assign y7 = n188 ;
  assign y8 = n189 ;
  assign y9 = n190 ;
  assign y10 = n192 ;
  assign y11 = n200 ;
  assign y12 = n207 ;
  assign y13 = n211 ;
  assign y14 = n219 ;
  assign y15 = n228 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
  assign y30 = 1'b0 ;
  assign y31 = 1'b0 ;
endmodule
