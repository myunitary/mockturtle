module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 ;
  assign n94 = x0 & ~x8 ;
  assign n49 = x8 ^ x0 ;
  assign n92 = x1 & ~x9 ;
  assign n93 = ~n49 & n92 ;
  assign n95 = n94 ^ n93 ;
  assign n50 = x9 ^ x1 ;
  assign n51 = n49 & n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n52 ^ n50 ;
  assign n89 = x2 & ~x10 ;
  assign n54 = x10 ^ x2 ;
  assign n85 = x3 & x11 ;
  assign n86 = n85 ^ x3 ;
  assign n87 = n54 & n86 ;
  assign n88 = n87 ^ n86 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = ~n53 & n90 ;
  assign n96 = n95 ^ n91 ;
  assign n55 = x11 ^ x3 ;
  assign n56 = n54 & n55 ;
  assign n57 = n56 ^ n54 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = ~n53 & ~n58 ;
  assign n81 = x4 & ~x12 ;
  assign n60 = x12 ^ x4 ;
  assign n79 = x5 & ~x13 ;
  assign n80 = ~n60 & n79 ;
  assign n82 = n81 ^ n80 ;
  assign n61 = x13 ^ x5 ;
  assign n62 = n60 & n61 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = n63 ^ n61 ;
  assign n76 = x6 & ~x14 ;
  assign n65 = x14 ^ x6 ;
  assign n72 = x7 & x15 ;
  assign n73 = n72 ^ x7 ;
  assign n74 = n65 & n73 ;
  assign n75 = n74 ^ n73 ;
  assign n77 = n76 ^ n75 ;
  assign n78 = ~n64 & n77 ;
  assign n83 = n82 ^ n78 ;
  assign n84 = n59 & n83 ;
  assign n97 = n96 ^ n84 ;
  assign n66 = x15 ^ x7 ;
  assign n67 = n65 & n66 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = n68 ^ n66 ;
  assign n70 = ~n64 & ~n69 ;
  assign n71 = n59 & n70 ;
  assign n98 = n97 ^ n71 ;
  assign n443 = x0 & ~n98 ;
  assign n100 = x8 & n98 ;
  assign n444 = n443 ^ n100 ;
  assign n101 = n100 ^ x8 ;
  assign n99 = x0 & n98 ;
  assign n102 = n101 ^ n99 ;
  assign n191 = ~x16 & n102 ;
  assign n103 = n102 ^ x16 ;
  assign n105 = x9 & n98 ;
  assign n106 = n105 ^ x9 ;
  assign n104 = x1 & n98 ;
  assign n107 = n106 ^ n104 ;
  assign n189 = ~x17 & n107 ;
  assign n190 = ~n103 & n189 ;
  assign n192 = n191 ^ n190 ;
  assign n108 = n107 ^ x17 ;
  assign n109 = n103 & n108 ;
  assign n110 = n109 ^ n103 ;
  assign n111 = n110 ^ n108 ;
  assign n113 = x10 & n98 ;
  assign n114 = n113 ^ x10 ;
  assign n112 = x2 & n98 ;
  assign n115 = n114 ^ n112 ;
  assign n186 = ~x18 & n115 ;
  assign n116 = n115 ^ x18 ;
  assign n118 = x11 & n98 ;
  assign n119 = n118 ^ x11 ;
  assign n117 = x3 & n98 ;
  assign n120 = n119 ^ n117 ;
  assign n182 = x19 & n120 ;
  assign n183 = n182 ^ n120 ;
  assign n184 = n116 & n183 ;
  assign n185 = n184 ^ n183 ;
  assign n187 = n186 ^ n185 ;
  assign n188 = ~n111 & n187 ;
  assign n193 = n192 ^ n188 ;
  assign n121 = n120 ^ x19 ;
  assign n122 = n116 & n121 ;
  assign n123 = n122 ^ n116 ;
  assign n124 = n123 ^ n121 ;
  assign n125 = ~n111 & ~n124 ;
  assign n127 = x12 & n98 ;
  assign n128 = n127 ^ x12 ;
  assign n126 = x4 & n98 ;
  assign n129 = n128 ^ n126 ;
  assign n178 = ~x20 & n129 ;
  assign n130 = n129 ^ x20 ;
  assign n132 = x13 & n98 ;
  assign n133 = n132 ^ x13 ;
  assign n131 = x5 & n98 ;
  assign n134 = n133 ^ n131 ;
  assign n174 = x21 & n134 ;
  assign n175 = n174 ^ n134 ;
  assign n176 = n130 & n175 ;
  assign n177 = n176 ^ n175 ;
  assign n179 = n178 ^ n177 ;
  assign n135 = n134 ^ x21 ;
  assign n136 = n130 & n135 ;
  assign n137 = n136 ^ n130 ;
  assign n138 = n137 ^ n135 ;
  assign n140 = x14 & n98 ;
  assign n141 = n140 ^ x14 ;
  assign n139 = x6 & n98 ;
  assign n142 = n141 ^ n139 ;
  assign n170 = x22 & n142 ;
  assign n171 = n170 ^ n142 ;
  assign n143 = n142 ^ x22 ;
  assign n156 = x15 & n59 ;
  assign n157 = n83 & n156 ;
  assign n153 = x15 & n71 ;
  assign n154 = n153 ^ x15 ;
  assign n152 = x15 & n96 ;
  assign n155 = n154 ^ n152 ;
  assign n158 = n157 ^ n155 ;
  assign n149 = x7 & n59 ;
  assign n150 = n83 & n149 ;
  assign n146 = x7 & n71 ;
  assign n147 = n146 ^ x7 ;
  assign n144 = x7 & n96 ;
  assign n145 = n144 ^ x7 ;
  assign n148 = n147 ^ n145 ;
  assign n151 = n150 ^ n148 ;
  assign n159 = n158 ^ n151 ;
  assign n166 = x23 & n159 ;
  assign n167 = n166 ^ n159 ;
  assign n168 = n143 & n167 ;
  assign n169 = n168 ^ n167 ;
  assign n172 = n171 ^ n169 ;
  assign n173 = ~n138 & n172 ;
  assign n180 = n179 ^ n173 ;
  assign n181 = n125 & n180 ;
  assign n194 = n193 ^ n181 ;
  assign n160 = n159 ^ x23 ;
  assign n161 = n143 & n160 ;
  assign n162 = n161 ^ n143 ;
  assign n163 = n162 ^ n160 ;
  assign n164 = ~n138 & ~n163 ;
  assign n165 = n125 & n164 ;
  assign n195 = n194 ^ n165 ;
  assign n198 = n102 & n195 ;
  assign n445 = n198 ^ n102 ;
  assign n196 = x16 & n195 ;
  assign n446 = n445 ^ n196 ;
  assign n536 = n444 & ~n446 ;
  assign n447 = n446 ^ n444 ;
  assign n448 = x1 & ~n98 ;
  assign n449 = n448 ^ n105 ;
  assign n203 = n107 & n195 ;
  assign n450 = n203 ^ n107 ;
  assign n201 = x17 & n195 ;
  assign n451 = n450 ^ n201 ;
  assign n534 = n449 & ~n451 ;
  assign n535 = ~n447 & n534 ;
  assign n537 = n536 ^ n535 ;
  assign n452 = n451 ^ n449 ;
  assign n453 = n447 & n452 ;
  assign n454 = n453 ^ n447 ;
  assign n455 = n454 ^ n452 ;
  assign n211 = n115 & n195 ;
  assign n456 = n211 ^ n115 ;
  assign n209 = x18 & n195 ;
  assign n457 = n456 ^ n209 ;
  assign n458 = x2 & ~n98 ;
  assign n459 = n458 ^ n113 ;
  assign n531 = ~n457 & n459 ;
  assign n460 = n459 ^ n457 ;
  assign n216 = n120 & n195 ;
  assign n461 = n216 ^ n120 ;
  assign n214 = x19 & n195 ;
  assign n462 = n461 ^ n214 ;
  assign n463 = x3 & ~n98 ;
  assign n464 = n463 ^ n118 ;
  assign n527 = n462 & n464 ;
  assign n528 = n527 ^ n464 ;
  assign n529 = n460 & n528 ;
  assign n530 = n529 ^ n528 ;
  assign n532 = n531 ^ n530 ;
  assign n533 = ~n455 & n532 ;
  assign n538 = n537 ^ n533 ;
  assign n465 = n464 ^ n462 ;
  assign n466 = n460 & n465 ;
  assign n467 = n466 ^ n460 ;
  assign n468 = n467 ^ n465 ;
  assign n469 = ~n455 & ~n468 ;
  assign n225 = n129 & n195 ;
  assign n470 = n225 ^ n129 ;
  assign n223 = x20 & n195 ;
  assign n471 = n470 ^ n223 ;
  assign n472 = x4 & ~n98 ;
  assign n473 = n472 ^ n127 ;
  assign n523 = ~n471 & n473 ;
  assign n474 = n473 ^ n471 ;
  assign n230 = n134 & n195 ;
  assign n475 = n230 ^ n134 ;
  assign n228 = x21 & n195 ;
  assign n476 = n475 ^ n228 ;
  assign n477 = x5 & ~n98 ;
  assign n478 = n477 ^ n132 ;
  assign n519 = n476 & n478 ;
  assign n520 = n519 ^ n478 ;
  assign n521 = n474 & n520 ;
  assign n522 = n521 ^ n520 ;
  assign n524 = n523 ^ n522 ;
  assign n479 = n478 ^ n476 ;
  assign n480 = n474 & n479 ;
  assign n481 = n480 ^ n474 ;
  assign n482 = n481 ^ n479 ;
  assign n485 = x6 & ~n98 ;
  assign n486 = n485 ^ n140 ;
  assign n515 = ~n142 & n486 ;
  assign n516 = ~n195 & n515 ;
  assign n491 = x7 & ~n98 ;
  assign n490 = x15 & n98 ;
  assign n492 = n491 ^ n490 ;
  assign n503 = ~n159 & n492 ;
  assign n504 = n195 & n503 ;
  assign n505 = n504 ^ n503 ;
  assign n501 = ~x23 & n492 ;
  assign n502 = n195 & n501 ;
  assign n506 = n505 ^ n502 ;
  assign n512 = n486 & n506 ;
  assign n238 = n142 & n195 ;
  assign n483 = n238 ^ n142 ;
  assign n509 = n483 ^ n195 ;
  assign n510 = n506 & ~n509 ;
  assign n236 = x22 & n195 ;
  assign n507 = n236 ^ n195 ;
  assign n508 = n506 & n507 ;
  assign n511 = n510 ^ n508 ;
  assign n513 = n512 ^ n511 ;
  assign n499 = ~x22 & n486 ;
  assign n500 = n195 & n499 ;
  assign n514 = n513 ^ n500 ;
  assign n517 = n516 ^ n514 ;
  assign n518 = ~n482 & n517 ;
  assign n525 = n524 ^ n518 ;
  assign n526 = n469 & n525 ;
  assign n539 = n538 ^ n526 ;
  assign n484 = n483 ^ n236 ;
  assign n487 = n486 ^ n484 ;
  assign n243 = n159 & n195 ;
  assign n488 = n243 ^ n159 ;
  assign n241 = x23 & n195 ;
  assign n489 = n488 ^ n241 ;
  assign n493 = n492 ^ n489 ;
  assign n494 = n487 & n493 ;
  assign n495 = n494 ^ n487 ;
  assign n496 = n495 ^ n493 ;
  assign n497 = ~n482 & ~n496 ;
  assign n498 = n469 & n497 ;
  assign n540 = n539 ^ n498 ;
  assign n809 = n444 & ~n540 ;
  assign n808 = n446 & n540 ;
  assign n810 = n809 ^ n808 ;
  assign n542 = n446 & ~n540 ;
  assign n541 = n444 & n540 ;
  assign n543 = n542 ^ n541 ;
  assign n197 = n196 ^ x16 ;
  assign n199 = n198 ^ n197 ;
  assign n287 = ~x24 & n199 ;
  assign n200 = n199 ^ x24 ;
  assign n202 = n201 ^ x17 ;
  assign n204 = n203 ^ n202 ;
  assign n285 = ~x25 & n204 ;
  assign n286 = ~n200 & n285 ;
  assign n288 = n287 ^ n286 ;
  assign n205 = n204 ^ x25 ;
  assign n206 = n200 & n205 ;
  assign n207 = n206 ^ n200 ;
  assign n208 = n207 ^ n205 ;
  assign n210 = n209 ^ x18 ;
  assign n212 = n211 ^ n210 ;
  assign n282 = ~x26 & n212 ;
  assign n213 = n212 ^ x26 ;
  assign n215 = n214 ^ x19 ;
  assign n217 = n216 ^ n215 ;
  assign n278 = x27 & n217 ;
  assign n279 = n278 ^ n217 ;
  assign n280 = n213 & n279 ;
  assign n281 = n280 ^ n279 ;
  assign n283 = n282 ^ n281 ;
  assign n284 = ~n208 & n283 ;
  assign n289 = n288 ^ n284 ;
  assign n218 = n217 ^ x27 ;
  assign n219 = n213 & n218 ;
  assign n220 = n219 ^ n213 ;
  assign n221 = n220 ^ n218 ;
  assign n222 = ~n208 & ~n221 ;
  assign n224 = n223 ^ x20 ;
  assign n226 = n225 ^ n224 ;
  assign n274 = ~x28 & n226 ;
  assign n227 = n226 ^ x28 ;
  assign n229 = n228 ^ x21 ;
  assign n231 = n230 ^ n229 ;
  assign n270 = x29 & n231 ;
  assign n271 = n270 ^ n231 ;
  assign n272 = n227 & n271 ;
  assign n273 = n272 ^ n271 ;
  assign n275 = n274 ^ n273 ;
  assign n232 = n231 ^ x29 ;
  assign n233 = n227 & n232 ;
  assign n234 = n233 ^ n227 ;
  assign n235 = n234 ^ n232 ;
  assign n266 = ~x30 & n142 ;
  assign n267 = n195 & n266 ;
  assign n256 = ~x31 & n159 ;
  assign n257 = n195 & n256 ;
  assign n253 = x23 & ~x31 ;
  assign n254 = n195 & n253 ;
  assign n255 = n254 ^ n253 ;
  assign n258 = n257 ^ n255 ;
  assign n262 = x30 & n258 ;
  assign n263 = n262 ^ n258 ;
  assign n237 = n236 ^ x22 ;
  assign n260 = n237 & n258 ;
  assign n259 = n238 & n258 ;
  assign n261 = n260 ^ n259 ;
  assign n264 = n263 ^ n261 ;
  assign n251 = x22 & ~x30 ;
  assign n252 = ~n195 & n251 ;
  assign n265 = n264 ^ n252 ;
  assign n268 = n267 ^ n265 ;
  assign n269 = ~n235 & n268 ;
  assign n276 = n275 ^ n269 ;
  assign n277 = n222 & n276 ;
  assign n290 = n289 ^ n277 ;
  assign n239 = n238 ^ n237 ;
  assign n240 = n239 ^ x30 ;
  assign n242 = n241 ^ x23 ;
  assign n244 = n243 ^ n242 ;
  assign n245 = n244 ^ x31 ;
  assign n246 = n240 & n245 ;
  assign n247 = n246 ^ n240 ;
  assign n248 = n247 ^ n245 ;
  assign n249 = ~n235 & ~n248 ;
  assign n250 = n222 & n249 ;
  assign n291 = n290 ^ n250 ;
  assign n545 = n199 & ~n291 ;
  assign n544 = x24 & n291 ;
  assign n546 = n545 ^ n544 ;
  assign n625 = n543 & ~n546 ;
  assign n547 = n546 ^ n543 ;
  assign n549 = n451 & ~n540 ;
  assign n548 = n449 & n540 ;
  assign n550 = n549 ^ n548 ;
  assign n552 = n204 & ~n291 ;
  assign n551 = x25 & n291 ;
  assign n553 = n552 ^ n551 ;
  assign n623 = n550 & ~n553 ;
  assign n624 = ~n547 & n623 ;
  assign n626 = n625 ^ n624 ;
  assign n554 = n553 ^ n550 ;
  assign n555 = ~n547 & ~n554 ;
  assign n557 = n212 & ~n291 ;
  assign n556 = x26 & n291 ;
  assign n558 = n557 ^ n556 ;
  assign n560 = n457 & ~n540 ;
  assign n559 = n459 & n540 ;
  assign n561 = n560 ^ n559 ;
  assign n620 = ~n558 & n561 ;
  assign n562 = n561 ^ n558 ;
  assign n564 = n217 & ~n291 ;
  assign n563 = x27 & n291 ;
  assign n565 = n564 ^ n563 ;
  assign n567 = n462 & ~n540 ;
  assign n566 = n464 & n540 ;
  assign n568 = n567 ^ n566 ;
  assign n618 = ~n565 & n568 ;
  assign n619 = ~n562 & n618 ;
  assign n621 = n620 ^ n619 ;
  assign n622 = n555 & n621 ;
  assign n627 = n626 ^ n622 ;
  assign n569 = n568 ^ n565 ;
  assign n570 = ~n562 & ~n569 ;
  assign n571 = n555 & n570 ;
  assign n573 = n226 & ~n291 ;
  assign n572 = x28 & n291 ;
  assign n574 = n573 ^ n572 ;
  assign n576 = n471 & ~n540 ;
  assign n575 = n473 & n540 ;
  assign n577 = n576 ^ n575 ;
  assign n614 = ~n574 & n577 ;
  assign n578 = n577 ^ n574 ;
  assign n580 = n231 & ~n291 ;
  assign n579 = x29 & n291 ;
  assign n581 = n580 ^ n579 ;
  assign n583 = n476 & ~n540 ;
  assign n582 = n478 & n540 ;
  assign n584 = n583 ^ n582 ;
  assign n612 = ~n581 & n584 ;
  assign n613 = ~n578 & n612 ;
  assign n615 = n614 ^ n613 ;
  assign n585 = n584 ^ n581 ;
  assign n586 = ~n578 & ~n585 ;
  assign n588 = n239 & ~n291 ;
  assign n587 = x30 & n291 ;
  assign n589 = n588 ^ n587 ;
  assign n591 = n484 & ~n540 ;
  assign n590 = n486 & n540 ;
  assign n592 = n591 ^ n590 ;
  assign n609 = ~n589 & n592 ;
  assign n593 = n592 ^ n589 ;
  assign n595 = n489 & n540 ;
  assign n596 = n595 ^ n489 ;
  assign n594 = n492 & n540 ;
  assign n597 = n596 ^ n594 ;
  assign n325 = n244 & n291 ;
  assign n599 = n325 ^ n244 ;
  assign n598 = x31 & n291 ;
  assign n600 = n599 ^ n598 ;
  assign n605 = n597 & n600 ;
  assign n606 = n605 ^ n597 ;
  assign n607 = n593 & n606 ;
  assign n608 = n607 ^ n606 ;
  assign n610 = n609 ^ n608 ;
  assign n611 = n586 & n610 ;
  assign n616 = n615 ^ n611 ;
  assign n617 = n571 & n616 ;
  assign n628 = n627 ^ n617 ;
  assign n601 = n600 ^ n597 ;
  assign n602 = ~n593 & ~n601 ;
  assign n603 = n586 & n602 ;
  assign n604 = n571 & n603 ;
  assign n629 = n628 ^ n604 ;
  assign n812 = n543 & ~n629 ;
  assign n811 = n546 & n629 ;
  assign n813 = n812 ^ n811 ;
  assign n901 = n810 & ~n813 ;
  assign n814 = n813 ^ n810 ;
  assign n816 = n449 & ~n540 ;
  assign n815 = n451 & n540 ;
  assign n817 = n816 ^ n815 ;
  assign n819 = n550 & ~n629 ;
  assign n818 = n553 & n629 ;
  assign n820 = n819 ^ n818 ;
  assign n899 = n817 & ~n820 ;
  assign n900 = ~n814 & n899 ;
  assign n902 = n901 ^ n900 ;
  assign n821 = n820 ^ n817 ;
  assign n822 = ~n814 & ~n821 ;
  assign n824 = n561 & ~n629 ;
  assign n823 = n558 & n629 ;
  assign n825 = n824 ^ n823 ;
  assign n827 = n459 & ~n540 ;
  assign n826 = n457 & n540 ;
  assign n828 = n827 ^ n826 ;
  assign n896 = ~n825 & n828 ;
  assign n829 = n828 ^ n825 ;
  assign n831 = n568 & ~n629 ;
  assign n830 = n565 & n629 ;
  assign n832 = n831 ^ n830 ;
  assign n834 = n464 & ~n540 ;
  assign n833 = n462 & n540 ;
  assign n835 = n834 ^ n833 ;
  assign n894 = ~n832 & n835 ;
  assign n895 = ~n829 & n894 ;
  assign n897 = n896 ^ n895 ;
  assign n898 = n822 & n897 ;
  assign n903 = n902 ^ n898 ;
  assign n836 = n835 ^ n832 ;
  assign n837 = ~n829 & ~n836 ;
  assign n838 = n822 & n837 ;
  assign n840 = n577 & ~n629 ;
  assign n839 = n574 & n629 ;
  assign n841 = n840 ^ n839 ;
  assign n843 = n473 & ~n540 ;
  assign n842 = n471 & n540 ;
  assign n844 = n843 ^ n842 ;
  assign n890 = ~n841 & n844 ;
  assign n845 = n844 ^ n841 ;
  assign n847 = n584 & ~n629 ;
  assign n846 = n581 & n629 ;
  assign n848 = n847 ^ n846 ;
  assign n850 = n478 & ~n540 ;
  assign n849 = n476 & n540 ;
  assign n851 = n850 ^ n849 ;
  assign n888 = ~n848 & n851 ;
  assign n889 = ~n845 & n888 ;
  assign n891 = n890 ^ n889 ;
  assign n852 = n851 ^ n848 ;
  assign n853 = ~n845 & ~n852 ;
  assign n858 = n486 & ~n540 ;
  assign n857 = n484 & n540 ;
  assign n859 = n858 ^ n857 ;
  assign n884 = ~n592 & n859 ;
  assign n885 = ~n629 & n884 ;
  assign n863 = n492 & ~n540 ;
  assign n864 = n863 ^ n595 ;
  assign n873 = ~n600 & n864 ;
  assign n874 = n629 & n873 ;
  assign n871 = ~n597 & n864 ;
  assign n872 = ~n629 & n871 ;
  assign n875 = n874 ^ n872 ;
  assign n881 = n859 & n875 ;
  assign n878 = ~n592 & ~n629 ;
  assign n879 = n875 & n878 ;
  assign n876 = ~n589 & n629 ;
  assign n877 = n875 & n876 ;
  assign n880 = n879 ^ n877 ;
  assign n882 = n881 ^ n880 ;
  assign n869 = ~n589 & n859 ;
  assign n870 = n629 & n869 ;
  assign n883 = n882 ^ n870 ;
  assign n886 = n885 ^ n883 ;
  assign n887 = n853 & n886 ;
  assign n892 = n891 ^ n887 ;
  assign n893 = n838 & n892 ;
  assign n904 = n903 ^ n893 ;
  assign n855 = n592 & ~n629 ;
  assign n854 = n589 & n629 ;
  assign n856 = n855 ^ n854 ;
  assign n860 = n859 ^ n856 ;
  assign n861 = n597 & ~n629 ;
  assign n684 = n600 & n629 ;
  assign n862 = n861 ^ n684 ;
  assign n865 = n864 ^ n862 ;
  assign n866 = ~n860 & ~n865 ;
  assign n867 = n853 & n866 ;
  assign n868 = n838 & n867 ;
  assign n905 = n904 ^ n868 ;
  assign n1084 = n810 & ~n905 ;
  assign n1083 = n813 & n905 ;
  assign n1085 = n1084 ^ n1083 ;
  assign n907 = n813 & ~n905 ;
  assign n906 = n810 & n905 ;
  assign n908 = n907 ^ n906 ;
  assign n631 = n546 & ~n629 ;
  assign n630 = n543 & n629 ;
  assign n632 = n631 ^ n630 ;
  assign n293 = x24 & ~n291 ;
  assign n292 = n199 & n291 ;
  assign n294 = n293 ^ n292 ;
  assign n361 = ~x32 & n294 ;
  assign n295 = n294 ^ x32 ;
  assign n297 = x25 & ~n291 ;
  assign n296 = n204 & n291 ;
  assign n298 = n297 ^ n296 ;
  assign n359 = ~x33 & n298 ;
  assign n360 = ~n295 & n359 ;
  assign n362 = n361 ^ n360 ;
  assign n299 = n298 ^ x33 ;
  assign n300 = ~n295 & ~n299 ;
  assign n302 = x26 & ~n291 ;
  assign n301 = n212 & n291 ;
  assign n303 = n302 ^ n301 ;
  assign n356 = ~x34 & n303 ;
  assign n304 = n303 ^ x34 ;
  assign n306 = x27 & ~n291 ;
  assign n305 = n217 & n291 ;
  assign n307 = n306 ^ n305 ;
  assign n354 = ~x35 & n307 ;
  assign n355 = ~n304 & n354 ;
  assign n357 = n356 ^ n355 ;
  assign n358 = n300 & n357 ;
  assign n363 = n362 ^ n358 ;
  assign n308 = n307 ^ x35 ;
  assign n309 = ~n304 & ~n308 ;
  assign n310 = n300 & n309 ;
  assign n312 = x28 & ~n291 ;
  assign n311 = n226 & n291 ;
  assign n313 = n312 ^ n311 ;
  assign n350 = ~x36 & n313 ;
  assign n314 = n313 ^ x36 ;
  assign n316 = x29 & ~n291 ;
  assign n315 = n231 & n291 ;
  assign n317 = n316 ^ n315 ;
  assign n348 = ~x37 & n317 ;
  assign n349 = ~n314 & n348 ;
  assign n351 = n350 ^ n349 ;
  assign n318 = n317 ^ x37 ;
  assign n319 = ~n314 & ~n318 ;
  assign n344 = ~x38 & n239 ;
  assign n345 = n291 & n344 ;
  assign n335 = ~x39 & n244 ;
  assign n336 = n291 & n335 ;
  assign n333 = x31 & ~x39 ;
  assign n334 = ~n291 & n333 ;
  assign n337 = n336 ^ n334 ;
  assign n341 = ~x38 & n337 ;
  assign n321 = x30 & ~n291 ;
  assign n339 = n321 & n337 ;
  assign n320 = n239 & n291 ;
  assign n338 = n320 & n337 ;
  assign n340 = n339 ^ n338 ;
  assign n342 = n341 ^ n340 ;
  assign n331 = x30 & ~x38 ;
  assign n332 = ~n291 & n331 ;
  assign n343 = n342 ^ n332 ;
  assign n346 = n345 ^ n343 ;
  assign n347 = n319 & n346 ;
  assign n352 = n351 ^ n347 ;
  assign n353 = n310 & n352 ;
  assign n364 = n363 ^ n353 ;
  assign n322 = n321 ^ n320 ;
  assign n323 = n322 ^ x38 ;
  assign n324 = x31 & ~n291 ;
  assign n326 = n325 ^ n324 ;
  assign n327 = n326 ^ x39 ;
  assign n328 = ~n323 & ~n327 ;
  assign n329 = n319 & n328 ;
  assign n330 = n310 & n329 ;
  assign n365 = n364 ^ n330 ;
  assign n634 = n294 & ~n365 ;
  assign n633 = x32 & n365 ;
  assign n635 = n634 ^ n633 ;
  assign n714 = n632 & ~n635 ;
  assign n636 = n635 ^ n632 ;
  assign n638 = n553 & ~n629 ;
  assign n637 = n550 & n629 ;
  assign n639 = n638 ^ n637 ;
  assign n641 = n298 & ~n365 ;
  assign n640 = x33 & n365 ;
  assign n642 = n641 ^ n640 ;
  assign n712 = n639 & ~n642 ;
  assign n713 = ~n636 & n712 ;
  assign n715 = n714 ^ n713 ;
  assign n643 = n642 ^ n639 ;
  assign n644 = ~n636 & ~n643 ;
  assign n646 = n303 & ~n365 ;
  assign n645 = x34 & n365 ;
  assign n647 = n646 ^ n645 ;
  assign n649 = n558 & ~n629 ;
  assign n648 = n561 & n629 ;
  assign n650 = n649 ^ n648 ;
  assign n709 = ~n647 & n650 ;
  assign n651 = n650 ^ n647 ;
  assign n653 = n307 & ~n365 ;
  assign n652 = x35 & n365 ;
  assign n654 = n653 ^ n652 ;
  assign n656 = n565 & ~n629 ;
  assign n655 = n568 & n629 ;
  assign n657 = n656 ^ n655 ;
  assign n707 = ~n654 & n657 ;
  assign n708 = ~n651 & n707 ;
  assign n710 = n709 ^ n708 ;
  assign n711 = n644 & n710 ;
  assign n716 = n715 ^ n711 ;
  assign n658 = n657 ^ n654 ;
  assign n659 = ~n651 & ~n658 ;
  assign n660 = n644 & n659 ;
  assign n662 = n313 & ~n365 ;
  assign n661 = x36 & n365 ;
  assign n663 = n662 ^ n661 ;
  assign n665 = n574 & ~n629 ;
  assign n664 = n577 & n629 ;
  assign n666 = n665 ^ n664 ;
  assign n703 = ~n663 & n666 ;
  assign n667 = n666 ^ n663 ;
  assign n669 = n317 & ~n365 ;
  assign n668 = x37 & n365 ;
  assign n670 = n669 ^ n668 ;
  assign n672 = n581 & ~n629 ;
  assign n671 = n584 & n629 ;
  assign n673 = n672 ^ n671 ;
  assign n701 = ~n670 & n673 ;
  assign n702 = ~n667 & n701 ;
  assign n704 = n703 ^ n702 ;
  assign n674 = n673 ^ n670 ;
  assign n675 = ~n667 & ~n674 ;
  assign n677 = n322 & ~n365 ;
  assign n676 = x38 & n365 ;
  assign n678 = n677 ^ n676 ;
  assign n680 = n589 & ~n629 ;
  assign n679 = n592 & n629 ;
  assign n681 = n680 ^ n679 ;
  assign n698 = ~n678 & n681 ;
  assign n682 = n681 ^ n678 ;
  assign n685 = n684 ^ n600 ;
  assign n683 = n597 & n629 ;
  assign n686 = n685 ^ n683 ;
  assign n688 = n326 & ~n365 ;
  assign n687 = x39 & n365 ;
  assign n689 = n688 ^ n687 ;
  assign n694 = n686 & n689 ;
  assign n695 = n694 ^ n686 ;
  assign n696 = n682 & n695 ;
  assign n697 = n696 ^ n695 ;
  assign n699 = n698 ^ n697 ;
  assign n700 = n675 & n699 ;
  assign n705 = n704 ^ n700 ;
  assign n706 = n660 & n705 ;
  assign n717 = n716 ^ n706 ;
  assign n690 = n689 ^ n686 ;
  assign n691 = ~n682 & ~n690 ;
  assign n692 = n675 & n691 ;
  assign n693 = n660 & n692 ;
  assign n718 = n717 ^ n693 ;
  assign n910 = n632 & ~n718 ;
  assign n909 = n635 & n718 ;
  assign n911 = n910 ^ n909 ;
  assign n988 = n908 & ~n911 ;
  assign n912 = n911 ^ n908 ;
  assign n914 = n820 & ~n905 ;
  assign n913 = n817 & n905 ;
  assign n915 = n914 ^ n913 ;
  assign n917 = n639 & ~n718 ;
  assign n916 = n642 & n718 ;
  assign n918 = n917 ^ n916 ;
  assign n986 = n915 & ~n918 ;
  assign n987 = ~n912 & n986 ;
  assign n989 = n988 ^ n987 ;
  assign n919 = n918 ^ n915 ;
  assign n920 = ~n912 & ~n919 ;
  assign n922 = n650 & ~n718 ;
  assign n921 = n647 & n718 ;
  assign n923 = n922 ^ n921 ;
  assign n925 = n825 & ~n905 ;
  assign n924 = n828 & n905 ;
  assign n926 = n925 ^ n924 ;
  assign n983 = ~n923 & n926 ;
  assign n927 = n926 ^ n923 ;
  assign n929 = n657 & ~n718 ;
  assign n928 = n654 & n718 ;
  assign n930 = n929 ^ n928 ;
  assign n932 = n832 & ~n905 ;
  assign n931 = n835 & n905 ;
  assign n933 = n932 ^ n931 ;
  assign n981 = ~n930 & n933 ;
  assign n982 = ~n927 & n981 ;
  assign n984 = n983 ^ n982 ;
  assign n985 = n920 & n984 ;
  assign n990 = n989 ^ n985 ;
  assign n934 = n933 ^ n930 ;
  assign n935 = ~n927 & ~n934 ;
  assign n936 = n920 & n935 ;
  assign n938 = n666 & ~n718 ;
  assign n937 = n663 & n718 ;
  assign n939 = n938 ^ n937 ;
  assign n941 = n841 & ~n905 ;
  assign n940 = n844 & n905 ;
  assign n942 = n941 ^ n940 ;
  assign n977 = ~n939 & n942 ;
  assign n943 = n942 ^ n939 ;
  assign n945 = n673 & ~n718 ;
  assign n944 = n670 & n718 ;
  assign n946 = n945 ^ n944 ;
  assign n948 = n848 & ~n905 ;
  assign n947 = n851 & n905 ;
  assign n949 = n948 ^ n947 ;
  assign n975 = ~n946 & n949 ;
  assign n976 = ~n943 & n975 ;
  assign n978 = n977 ^ n976 ;
  assign n950 = n949 ^ n946 ;
  assign n951 = ~n943 & ~n950 ;
  assign n953 = n681 & ~n718 ;
  assign n952 = n678 & n718 ;
  assign n954 = n953 ^ n952 ;
  assign n956 = n856 & ~n905 ;
  assign n955 = n859 & n905 ;
  assign n957 = n956 ^ n955 ;
  assign n972 = ~n954 & n957 ;
  assign n958 = n957 ^ n954 ;
  assign n960 = n862 & ~n905 ;
  assign n959 = n864 & n905 ;
  assign n961 = n960 ^ n959 ;
  assign n774 = n686 & n718 ;
  assign n962 = n774 ^ n686 ;
  assign n772 = n689 & n718 ;
  assign n963 = n962 ^ n772 ;
  assign n968 = n961 & n963 ;
  assign n969 = n968 ^ n961 ;
  assign n970 = n958 & n969 ;
  assign n971 = n970 ^ n969 ;
  assign n973 = n972 ^ n971 ;
  assign n974 = n951 & n973 ;
  assign n979 = n978 ^ n974 ;
  assign n980 = n936 & n979 ;
  assign n991 = n990 ^ n980 ;
  assign n964 = n963 ^ n961 ;
  assign n965 = ~n958 & ~n964 ;
  assign n966 = n951 & n965 ;
  assign n967 = n936 & n966 ;
  assign n992 = n991 ^ n967 ;
  assign n1087 = n908 & ~n992 ;
  assign n1086 = n911 & n992 ;
  assign n1088 = n1087 ^ n1086 ;
  assign n1177 = n1085 & ~n1088 ;
  assign n1089 = n1088 ^ n1085 ;
  assign n1091 = n817 & ~n905 ;
  assign n1090 = n820 & n905 ;
  assign n1092 = n1091 ^ n1090 ;
  assign n1094 = n915 & ~n992 ;
  assign n1093 = n918 & n992 ;
  assign n1095 = n1094 ^ n1093 ;
  assign n1175 = n1092 & ~n1095 ;
  assign n1176 = ~n1089 & n1175 ;
  assign n1178 = n1177 ^ n1176 ;
  assign n1096 = n1095 ^ n1092 ;
  assign n1097 = ~n1089 & ~n1096 ;
  assign n1099 = n926 & ~n992 ;
  assign n1098 = n923 & n992 ;
  assign n1100 = n1099 ^ n1098 ;
  assign n1102 = n828 & ~n905 ;
  assign n1101 = n825 & n905 ;
  assign n1103 = n1102 ^ n1101 ;
  assign n1172 = ~n1100 & n1103 ;
  assign n1104 = n1103 ^ n1100 ;
  assign n1106 = n933 & ~n992 ;
  assign n1105 = n930 & n992 ;
  assign n1107 = n1106 ^ n1105 ;
  assign n1109 = n835 & ~n905 ;
  assign n1108 = n832 & n905 ;
  assign n1110 = n1109 ^ n1108 ;
  assign n1170 = ~n1107 & n1110 ;
  assign n1171 = ~n1104 & n1170 ;
  assign n1173 = n1172 ^ n1171 ;
  assign n1174 = n1097 & n1173 ;
  assign n1179 = n1178 ^ n1174 ;
  assign n1111 = n1110 ^ n1107 ;
  assign n1112 = ~n1104 & ~n1111 ;
  assign n1113 = n1097 & n1112 ;
  assign n1115 = n942 & ~n992 ;
  assign n1114 = n939 & n992 ;
  assign n1116 = n1115 ^ n1114 ;
  assign n1118 = n844 & ~n905 ;
  assign n1117 = n841 & n905 ;
  assign n1119 = n1118 ^ n1117 ;
  assign n1166 = ~n1116 & n1119 ;
  assign n1120 = n1119 ^ n1116 ;
  assign n1122 = n949 & ~n992 ;
  assign n1121 = n946 & n992 ;
  assign n1123 = n1122 ^ n1121 ;
  assign n1125 = n851 & ~n905 ;
  assign n1124 = n848 & n905 ;
  assign n1126 = n1125 ^ n1124 ;
  assign n1164 = ~n1123 & n1126 ;
  assign n1165 = ~n1120 & n1164 ;
  assign n1167 = n1166 ^ n1165 ;
  assign n1127 = n1126 ^ n1123 ;
  assign n1128 = ~n1120 & ~n1127 ;
  assign n1133 = n859 & ~n905 ;
  assign n1132 = n856 & n905 ;
  assign n1134 = n1133 ^ n1132 ;
  assign n1160 = ~n957 & n1134 ;
  assign n1161 = ~n992 & n1160 ;
  assign n1139 = n864 & ~n905 ;
  assign n1138 = n862 & n905 ;
  assign n1140 = n1139 ^ n1138 ;
  assign n1149 = ~n963 & n1140 ;
  assign n1150 = n992 & n1149 ;
  assign n1147 = ~n961 & n1140 ;
  assign n1148 = ~n992 & n1147 ;
  assign n1151 = n1150 ^ n1148 ;
  assign n1157 = n1134 & n1151 ;
  assign n1154 = ~n957 & ~n992 ;
  assign n1155 = n1151 & n1154 ;
  assign n1152 = ~n954 & n992 ;
  assign n1153 = n1151 & n1152 ;
  assign n1156 = n1155 ^ n1153 ;
  assign n1158 = n1157 ^ n1156 ;
  assign n1145 = ~n954 & n1134 ;
  assign n1146 = n992 & n1145 ;
  assign n1159 = n1158 ^ n1146 ;
  assign n1162 = n1161 ^ n1159 ;
  assign n1163 = n1128 & n1162 ;
  assign n1168 = n1167 ^ n1163 ;
  assign n1169 = n1113 & n1168 ;
  assign n1180 = n1179 ^ n1169 ;
  assign n1130 = n957 & ~n992 ;
  assign n1129 = n954 & n992 ;
  assign n1131 = n1130 ^ n1129 ;
  assign n1135 = n1134 ^ n1131 ;
  assign n1136 = n961 & ~n992 ;
  assign n1048 = n963 & n992 ;
  assign n1137 = n1136 ^ n1048 ;
  assign n1141 = n1140 ^ n1137 ;
  assign n1142 = ~n1135 & ~n1141 ;
  assign n1143 = n1128 & n1142 ;
  assign n1144 = n1113 & n1143 ;
  assign n1181 = n1180 ^ n1144 ;
  assign n1273 = n1085 & ~n1181 ;
  assign n1272 = n1088 & n1181 ;
  assign n1274 = n1273 ^ n1272 ;
  assign n1183 = n1088 & ~n1181 ;
  assign n1182 = n1085 & n1181 ;
  assign n1184 = n1183 ^ n1182 ;
  assign n994 = n911 & ~n992 ;
  assign n993 = n908 & n992 ;
  assign n995 = n994 ^ n993 ;
  assign n720 = n635 & ~n718 ;
  assign n719 = n632 & n718 ;
  assign n721 = n720 ^ n719 ;
  assign n367 = x32 & ~n365 ;
  assign n366 = n294 & n365 ;
  assign n368 = n367 ^ n366 ;
  assign n435 = ~x40 & n368 ;
  assign n369 = n368 ^ x40 ;
  assign n371 = x33 & ~n365 ;
  assign n370 = n298 & n365 ;
  assign n372 = n371 ^ n370 ;
  assign n433 = ~x41 & n372 ;
  assign n434 = ~n369 & n433 ;
  assign n436 = n435 ^ n434 ;
  assign n373 = n372 ^ x41 ;
  assign n374 = ~n369 & ~n373 ;
  assign n376 = x34 & ~n365 ;
  assign n375 = n303 & n365 ;
  assign n377 = n376 ^ n375 ;
  assign n430 = ~x42 & n377 ;
  assign n378 = n377 ^ x42 ;
  assign n380 = x35 & ~n365 ;
  assign n379 = n307 & n365 ;
  assign n381 = n380 ^ n379 ;
  assign n428 = ~x43 & n381 ;
  assign n429 = ~n378 & n428 ;
  assign n431 = n430 ^ n429 ;
  assign n432 = n374 & n431 ;
  assign n437 = n436 ^ n432 ;
  assign n382 = n381 ^ x43 ;
  assign n383 = ~n378 & ~n382 ;
  assign n384 = n374 & n383 ;
  assign n386 = x36 & ~n365 ;
  assign n385 = n313 & n365 ;
  assign n387 = n386 ^ n385 ;
  assign n424 = ~x44 & n387 ;
  assign n388 = n387 ^ x44 ;
  assign n390 = x37 & ~n365 ;
  assign n389 = n317 & n365 ;
  assign n391 = n390 ^ n389 ;
  assign n422 = ~x45 & n391 ;
  assign n423 = ~n388 & n422 ;
  assign n425 = n424 ^ n423 ;
  assign n392 = n391 ^ x45 ;
  assign n393 = ~n388 & ~n392 ;
  assign n418 = ~x46 & n322 ;
  assign n419 = n365 & n418 ;
  assign n409 = ~x47 & n326 ;
  assign n410 = n365 & n409 ;
  assign n407 = x39 & ~x47 ;
  assign n408 = ~n365 & n407 ;
  assign n411 = n410 ^ n408 ;
  assign n415 = ~x46 & n411 ;
  assign n395 = x38 & ~n365 ;
  assign n413 = n395 & n411 ;
  assign n394 = n322 & n365 ;
  assign n412 = n394 & n411 ;
  assign n414 = n413 ^ n412 ;
  assign n416 = n415 ^ n414 ;
  assign n405 = x38 & ~x46 ;
  assign n406 = ~n365 & n405 ;
  assign n417 = n416 ^ n406 ;
  assign n420 = n419 ^ n417 ;
  assign n421 = n393 & n420 ;
  assign n426 = n425 ^ n421 ;
  assign n427 = n384 & n426 ;
  assign n438 = n437 ^ n427 ;
  assign n396 = n395 ^ n394 ;
  assign n397 = n396 ^ x46 ;
  assign n399 = x39 & ~n365 ;
  assign n398 = n326 & n365 ;
  assign n400 = n399 ^ n398 ;
  assign n401 = n400 ^ x47 ;
  assign n402 = ~n397 & ~n401 ;
  assign n403 = n393 & n402 ;
  assign n404 = n384 & n403 ;
  assign n439 = n438 ^ n404 ;
  assign n441 = n368 & ~n439 ;
  assign n440 = x40 & n439 ;
  assign n442 = n441 ^ n440 ;
  assign n800 = ~n442 & n721 ;
  assign n722 = n721 ^ n442 ;
  assign n724 = n372 & ~n439 ;
  assign n723 = x41 & n439 ;
  assign n725 = n724 ^ n723 ;
  assign n727 = n642 & ~n718 ;
  assign n726 = n639 & n718 ;
  assign n728 = n727 ^ n726 ;
  assign n798 = ~n725 & n728 ;
  assign n799 = ~n722 & n798 ;
  assign n801 = n800 ^ n799 ;
  assign n729 = n728 ^ n725 ;
  assign n730 = ~n722 & ~n729 ;
  assign n732 = n377 & ~n439 ;
  assign n731 = x42 & n439 ;
  assign n733 = n732 ^ n731 ;
  assign n735 = n647 & ~n718 ;
  assign n734 = n650 & n718 ;
  assign n736 = n735 ^ n734 ;
  assign n795 = ~n733 & n736 ;
  assign n737 = n736 ^ n733 ;
  assign n739 = n381 & ~n439 ;
  assign n738 = x43 & n439 ;
  assign n740 = n739 ^ n738 ;
  assign n742 = n654 & ~n718 ;
  assign n741 = n657 & n718 ;
  assign n743 = n742 ^ n741 ;
  assign n793 = ~n740 & n743 ;
  assign n794 = ~n737 & n793 ;
  assign n796 = n795 ^ n794 ;
  assign n797 = n730 & n796 ;
  assign n802 = n801 ^ n797 ;
  assign n744 = n743 ^ n740 ;
  assign n745 = ~n737 & ~n744 ;
  assign n746 = n730 & n745 ;
  assign n748 = n387 & ~n439 ;
  assign n747 = x44 & n439 ;
  assign n749 = n748 ^ n747 ;
  assign n751 = n663 & ~n718 ;
  assign n750 = n666 & n718 ;
  assign n752 = n751 ^ n750 ;
  assign n789 = ~n749 & n752 ;
  assign n753 = n752 ^ n749 ;
  assign n755 = n391 & ~n439 ;
  assign n754 = x45 & n439 ;
  assign n756 = n755 ^ n754 ;
  assign n758 = n670 & ~n718 ;
  assign n757 = n673 & n718 ;
  assign n759 = n758 ^ n757 ;
  assign n787 = ~n756 & n759 ;
  assign n788 = ~n753 & n787 ;
  assign n790 = n789 ^ n788 ;
  assign n760 = n759 ^ n756 ;
  assign n761 = ~n753 & ~n760 ;
  assign n763 = n396 & ~n439 ;
  assign n762 = x46 & n439 ;
  assign n764 = n763 ^ n762 ;
  assign n766 = n678 & ~n718 ;
  assign n765 = n681 & n718 ;
  assign n767 = n766 ^ n765 ;
  assign n784 = ~n764 & n767 ;
  assign n768 = n767 ^ n764 ;
  assign n770 = n400 & ~n439 ;
  assign n769 = x47 & n439 ;
  assign n771 = n770 ^ n769 ;
  assign n773 = n772 ^ n689 ;
  assign n775 = n774 ^ n773 ;
  assign n780 = n771 & n775 ;
  assign n781 = n780 ^ n775 ;
  assign n782 = n768 & n781 ;
  assign n783 = n782 ^ n781 ;
  assign n785 = n784 ^ n783 ;
  assign n786 = n761 & n785 ;
  assign n791 = n790 ^ n786 ;
  assign n792 = n746 & n791 ;
  assign n803 = n802 ^ n792 ;
  assign n776 = n775 ^ n771 ;
  assign n777 = ~n768 & ~n776 ;
  assign n778 = n761 & n777 ;
  assign n779 = n746 & n778 ;
  assign n804 = n803 ^ n779 ;
  assign n806 = n721 & ~n804 ;
  assign n805 = n442 & n804 ;
  assign n807 = n806 ^ n805 ;
  assign n1075 = ~n807 & n995 ;
  assign n996 = n995 ^ n807 ;
  assign n998 = n728 & ~n804 ;
  assign n997 = n725 & n804 ;
  assign n999 = n998 ^ n997 ;
  assign n1001 = n918 & ~n992 ;
  assign n1000 = n915 & n992 ;
  assign n1002 = n1001 ^ n1000 ;
  assign n1073 = ~n999 & n1002 ;
  assign n1074 = ~n996 & n1073 ;
  assign n1076 = n1075 ^ n1074 ;
  assign n1003 = n1002 ^ n999 ;
  assign n1004 = ~n996 & ~n1003 ;
  assign n1006 = n736 & ~n804 ;
  assign n1005 = n733 & n804 ;
  assign n1007 = n1006 ^ n1005 ;
  assign n1009 = n923 & ~n992 ;
  assign n1008 = n926 & n992 ;
  assign n1010 = n1009 ^ n1008 ;
  assign n1070 = ~n1007 & n1010 ;
  assign n1011 = n1010 ^ n1007 ;
  assign n1013 = n743 & ~n804 ;
  assign n1012 = n740 & n804 ;
  assign n1014 = n1013 ^ n1012 ;
  assign n1016 = n930 & ~n992 ;
  assign n1015 = n933 & n992 ;
  assign n1017 = n1016 ^ n1015 ;
  assign n1068 = ~n1014 & n1017 ;
  assign n1069 = ~n1011 & n1068 ;
  assign n1071 = n1070 ^ n1069 ;
  assign n1072 = n1004 & n1071 ;
  assign n1077 = n1076 ^ n1072 ;
  assign n1018 = n1017 ^ n1014 ;
  assign n1019 = ~n1011 & ~n1018 ;
  assign n1020 = n1004 & n1019 ;
  assign n1022 = n752 & ~n804 ;
  assign n1021 = n749 & n804 ;
  assign n1023 = n1022 ^ n1021 ;
  assign n1025 = n939 & ~n992 ;
  assign n1024 = n942 & n992 ;
  assign n1026 = n1025 ^ n1024 ;
  assign n1064 = ~n1023 & n1026 ;
  assign n1027 = n1026 ^ n1023 ;
  assign n1029 = n759 & ~n804 ;
  assign n1028 = n756 & n804 ;
  assign n1030 = n1029 ^ n1028 ;
  assign n1032 = n946 & ~n992 ;
  assign n1031 = n949 & n992 ;
  assign n1033 = n1032 ^ n1031 ;
  assign n1062 = ~n1030 & n1033 ;
  assign n1063 = ~n1027 & n1062 ;
  assign n1065 = n1064 ^ n1063 ;
  assign n1034 = n1033 ^ n1030 ;
  assign n1035 = ~n1027 & ~n1034 ;
  assign n1037 = n767 & ~n804 ;
  assign n1036 = n764 & n804 ;
  assign n1038 = n1037 ^ n1036 ;
  assign n1040 = n954 & ~n992 ;
  assign n1039 = n957 & n992 ;
  assign n1041 = n1040 ^ n1039 ;
  assign n1059 = ~n1038 & n1041 ;
  assign n1042 = n1041 ^ n1038 ;
  assign n1044 = n775 & n804 ;
  assign n1045 = n1044 ^ n775 ;
  assign n1043 = n771 & n804 ;
  assign n1046 = n1045 ^ n1043 ;
  assign n1049 = n1048 ^ n963 ;
  assign n1047 = n961 & n992 ;
  assign n1050 = n1049 ^ n1047 ;
  assign n1055 = n1046 & n1050 ;
  assign n1056 = n1055 ^ n1050 ;
  assign n1057 = n1042 & n1056 ;
  assign n1058 = n1057 ^ n1056 ;
  assign n1060 = n1059 ^ n1058 ;
  assign n1061 = n1035 & n1060 ;
  assign n1066 = n1065 ^ n1061 ;
  assign n1067 = n1020 & n1066 ;
  assign n1078 = n1077 ^ n1067 ;
  assign n1051 = n1050 ^ n1046 ;
  assign n1052 = ~n1042 & ~n1051 ;
  assign n1053 = n1035 & n1052 ;
  assign n1054 = n1020 & n1053 ;
  assign n1079 = n1078 ^ n1054 ;
  assign n1081 = n995 & ~n1079 ;
  assign n1080 = n807 & n1079 ;
  assign n1082 = n1081 ^ n1080 ;
  assign n1263 = ~n1082 & n1184 ;
  assign n1185 = n1184 ^ n1082 ;
  assign n1187 = n1002 & ~n1079 ;
  assign n1186 = n999 & n1079 ;
  assign n1188 = n1187 ^ n1186 ;
  assign n1190 = n1095 & ~n1181 ;
  assign n1189 = n1092 & n1181 ;
  assign n1191 = n1190 ^ n1189 ;
  assign n1261 = ~n1188 & n1191 ;
  assign n1262 = ~n1185 & n1261 ;
  assign n1264 = n1263 ^ n1262 ;
  assign n1192 = n1191 ^ n1188 ;
  assign n1193 = ~n1185 & ~n1192 ;
  assign n1195 = n1010 & ~n1079 ;
  assign n1194 = n1007 & n1079 ;
  assign n1196 = n1195 ^ n1194 ;
  assign n1198 = n1100 & ~n1181 ;
  assign n1197 = n1103 & n1181 ;
  assign n1199 = n1198 ^ n1197 ;
  assign n1258 = ~n1196 & n1199 ;
  assign n1200 = n1199 ^ n1196 ;
  assign n1202 = n1017 & ~n1079 ;
  assign n1201 = n1014 & n1079 ;
  assign n1203 = n1202 ^ n1201 ;
  assign n1205 = n1107 & ~n1181 ;
  assign n1204 = n1110 & n1181 ;
  assign n1206 = n1205 ^ n1204 ;
  assign n1256 = ~n1203 & n1206 ;
  assign n1257 = ~n1200 & n1256 ;
  assign n1259 = n1258 ^ n1257 ;
  assign n1260 = n1193 & n1259 ;
  assign n1265 = n1264 ^ n1260 ;
  assign n1207 = n1206 ^ n1203 ;
  assign n1208 = ~n1200 & ~n1207 ;
  assign n1209 = n1193 & n1208 ;
  assign n1211 = n1026 & ~n1079 ;
  assign n1210 = n1023 & n1079 ;
  assign n1212 = n1211 ^ n1210 ;
  assign n1214 = n1116 & ~n1181 ;
  assign n1213 = n1119 & n1181 ;
  assign n1215 = n1214 ^ n1213 ;
  assign n1252 = ~n1212 & n1215 ;
  assign n1216 = n1215 ^ n1212 ;
  assign n1218 = n1033 & ~n1079 ;
  assign n1217 = n1030 & n1079 ;
  assign n1219 = n1218 ^ n1217 ;
  assign n1221 = n1123 & ~n1181 ;
  assign n1220 = n1126 & n1181 ;
  assign n1222 = n1221 ^ n1220 ;
  assign n1250 = ~n1219 & n1222 ;
  assign n1251 = ~n1216 & n1250 ;
  assign n1253 = n1252 ^ n1251 ;
  assign n1223 = n1222 ^ n1219 ;
  assign n1224 = ~n1216 & ~n1223 ;
  assign n1226 = n1041 & ~n1079 ;
  assign n1225 = n1038 & n1079 ;
  assign n1227 = n1226 ^ n1225 ;
  assign n1229 = n1131 & ~n1181 ;
  assign n1228 = n1134 & n1181 ;
  assign n1230 = n1229 ^ n1228 ;
  assign n1247 = ~n1227 & n1230 ;
  assign n1231 = n1230 ^ n1227 ;
  assign n1233 = n1050 & n1079 ;
  assign n1234 = n1233 ^ n1050 ;
  assign n1232 = n1046 & n1079 ;
  assign n1235 = n1234 ^ n1232 ;
  assign n1237 = n1137 & ~n1181 ;
  assign n1236 = n1140 & n1181 ;
  assign n1238 = n1237 ^ n1236 ;
  assign n1243 = n1235 & n1238 ;
  assign n1244 = n1243 ^ n1238 ;
  assign n1245 = n1231 & n1244 ;
  assign n1246 = n1245 ^ n1244 ;
  assign n1248 = n1247 ^ n1246 ;
  assign n1249 = n1224 & n1248 ;
  assign n1254 = n1253 ^ n1249 ;
  assign n1255 = n1209 & n1254 ;
  assign n1266 = n1265 ^ n1255 ;
  assign n1239 = n1238 ^ n1235 ;
  assign n1240 = ~n1231 & ~n1239 ;
  assign n1241 = n1224 & n1240 ;
  assign n1242 = n1209 & n1241 ;
  assign n1267 = n1266 ^ n1242 ;
  assign n1269 = n1184 & n1267 ;
  assign n1270 = n1269 ^ n1184 ;
  assign n1268 = n1082 & n1267 ;
  assign n1271 = n1270 ^ n1268 ;
  assign n1384 = ~n1271 & n1274 ;
  assign n1275 = n1274 ^ n1271 ;
  assign n1277 = n1191 & n1267 ;
  assign n1278 = n1277 ^ n1191 ;
  assign n1276 = n1188 & n1267 ;
  assign n1279 = n1278 ^ n1276 ;
  assign n1281 = n1092 & ~n1181 ;
  assign n1280 = n1095 & n1181 ;
  assign n1282 = n1281 ^ n1280 ;
  assign n1382 = ~n1279 & n1282 ;
  assign n1383 = ~n1275 & n1382 ;
  assign n1385 = n1384 ^ n1383 ;
  assign n1283 = n1282 ^ n1279 ;
  assign n1284 = n1275 & n1283 ;
  assign n1285 = n1284 ^ n1275 ;
  assign n1286 = n1285 ^ n1283 ;
  assign n1288 = n1199 & n1267 ;
  assign n1289 = n1288 ^ n1199 ;
  assign n1287 = n1196 & n1267 ;
  assign n1290 = n1289 ^ n1287 ;
  assign n1292 = n1103 & ~n1181 ;
  assign n1291 = n1100 & n1181 ;
  assign n1293 = n1292 ^ n1291 ;
  assign n1379 = ~n1290 & n1293 ;
  assign n1294 = n1293 ^ n1290 ;
  assign n1296 = n1206 & n1267 ;
  assign n1297 = n1296 ^ n1206 ;
  assign n1295 = n1203 & n1267 ;
  assign n1298 = n1297 ^ n1295 ;
  assign n1300 = n1110 & ~n1181 ;
  assign n1299 = n1107 & n1181 ;
  assign n1301 = n1300 ^ n1299 ;
  assign n1375 = n1298 & n1301 ;
  assign n1376 = n1375 ^ n1301 ;
  assign n1377 = n1294 & n1376 ;
  assign n1378 = n1377 ^ n1376 ;
  assign n1380 = n1379 ^ n1378 ;
  assign n1381 = ~n1286 & n1380 ;
  assign n1386 = n1385 ^ n1381 ;
  assign n1302 = n1301 ^ n1298 ;
  assign n1303 = n1294 & n1302 ;
  assign n1304 = n1303 ^ n1294 ;
  assign n1305 = n1304 ^ n1302 ;
  assign n1306 = ~n1286 & ~n1305 ;
  assign n1308 = n1215 & n1267 ;
  assign n1309 = n1308 ^ n1215 ;
  assign n1307 = n1212 & n1267 ;
  assign n1310 = n1309 ^ n1307 ;
  assign n1312 = n1119 & ~n1181 ;
  assign n1311 = n1116 & n1181 ;
  assign n1313 = n1312 ^ n1311 ;
  assign n1371 = ~n1310 & n1313 ;
  assign n1314 = n1313 ^ n1310 ;
  assign n1316 = n1222 & n1267 ;
  assign n1317 = n1316 ^ n1222 ;
  assign n1315 = n1219 & n1267 ;
  assign n1318 = n1317 ^ n1315 ;
  assign n1320 = n1126 & ~n1181 ;
  assign n1319 = n1123 & n1181 ;
  assign n1321 = n1320 ^ n1319 ;
  assign n1367 = n1318 & n1321 ;
  assign n1368 = n1367 ^ n1321 ;
  assign n1369 = n1314 & n1368 ;
  assign n1370 = n1369 ^ n1368 ;
  assign n1372 = n1371 ^ n1370 ;
  assign n1322 = n1321 ^ n1318 ;
  assign n1323 = n1314 & n1322 ;
  assign n1324 = n1323 ^ n1314 ;
  assign n1325 = n1324 ^ n1322 ;
  assign n1331 = n1134 & ~n1181 ;
  assign n1330 = n1131 & n1181 ;
  assign n1332 = n1331 ^ n1330 ;
  assign n1363 = ~n1230 & n1332 ;
  assign n1364 = ~n1267 & n1363 ;
  assign n1339 = n1140 & ~n1181 ;
  assign n1338 = n1137 & n1181 ;
  assign n1340 = n1339 ^ n1338 ;
  assign n1351 = ~n1238 & n1340 ;
  assign n1352 = n1267 & n1351 ;
  assign n1353 = n1352 ^ n1351 ;
  assign n1349 = ~n1235 & n1340 ;
  assign n1350 = n1267 & n1349 ;
  assign n1354 = n1353 ^ n1350 ;
  assign n1360 = n1332 & n1354 ;
  assign n1327 = n1230 & n1267 ;
  assign n1328 = n1327 ^ n1230 ;
  assign n1357 = n1328 ^ n1267 ;
  assign n1358 = n1354 & ~n1357 ;
  assign n1326 = n1227 & n1267 ;
  assign n1355 = n1326 ^ n1267 ;
  assign n1356 = n1354 & n1355 ;
  assign n1359 = n1358 ^ n1356 ;
  assign n1361 = n1360 ^ n1359 ;
  assign n1347 = ~n1227 & n1332 ;
  assign n1348 = n1267 & n1347 ;
  assign n1362 = n1361 ^ n1348 ;
  assign n1365 = n1364 ^ n1362 ;
  assign n1366 = ~n1325 & n1365 ;
  assign n1373 = n1372 ^ n1366 ;
  assign n1374 = n1306 & n1373 ;
  assign n1387 = n1386 ^ n1374 ;
  assign n1329 = n1328 ^ n1326 ;
  assign n1333 = n1332 ^ n1329 ;
  assign n1335 = n1238 & n1267 ;
  assign n1336 = n1335 ^ n1238 ;
  assign n1334 = n1235 & n1267 ;
  assign n1337 = n1336 ^ n1334 ;
  assign n1341 = n1340 ^ n1337 ;
  assign n1342 = n1333 & n1341 ;
  assign n1343 = n1342 ^ n1333 ;
  assign n1344 = n1343 ^ n1341 ;
  assign n1345 = ~n1325 & ~n1344 ;
  assign n1346 = n1306 & n1345 ;
  assign n1388 = n1387 ^ n1346 ;
  assign n1390 = n1274 & n1388 ;
  assign n1391 = n1390 ^ n1274 ;
  assign n1389 = n1271 & n1388 ;
  assign n1392 = n1391 ^ n1389 ;
  assign n1394 = n1282 & n1388 ;
  assign n1395 = n1394 ^ n1282 ;
  assign n1393 = n1279 & n1388 ;
  assign n1396 = n1395 ^ n1393 ;
  assign n1398 = n1293 & n1388 ;
  assign n1399 = n1398 ^ n1293 ;
  assign n1397 = n1290 & n1388 ;
  assign n1400 = n1399 ^ n1397 ;
  assign n1402 = n1301 & n1388 ;
  assign n1403 = n1402 ^ n1301 ;
  assign n1401 = n1298 & n1388 ;
  assign n1404 = n1403 ^ n1401 ;
  assign n1406 = n1313 & n1388 ;
  assign n1407 = n1406 ^ n1313 ;
  assign n1405 = n1310 & n1388 ;
  assign n1408 = n1407 ^ n1405 ;
  assign n1410 = n1321 & n1388 ;
  assign n1411 = n1410 ^ n1321 ;
  assign n1409 = n1318 & n1388 ;
  assign n1412 = n1411 ^ n1409 ;
  assign n1414 = n1332 & n1388 ;
  assign n1415 = n1414 ^ n1332 ;
  assign n1413 = n1329 & n1388 ;
  assign n1416 = n1415 ^ n1413 ;
  assign n1418 = n1340 & n1388 ;
  assign n1419 = n1418 ^ n1340 ;
  assign n1417 = n1337 & n1388 ;
  assign n1420 = n1419 ^ n1417 ;
  assign n1421 = n1389 ^ n1271 ;
  assign n1422 = n1421 ^ n1390 ;
  assign n1423 = n1393 ^ n1279 ;
  assign n1424 = n1423 ^ n1394 ;
  assign n1425 = n1397 ^ n1290 ;
  assign n1426 = n1425 ^ n1398 ;
  assign n1427 = n1401 ^ n1298 ;
  assign n1428 = n1427 ^ n1402 ;
  assign n1429 = n1405 ^ n1310 ;
  assign n1430 = n1429 ^ n1406 ;
  assign n1431 = n1409 ^ n1318 ;
  assign n1432 = n1431 ^ n1410 ;
  assign n1433 = n1413 ^ n1329 ;
  assign n1434 = n1433 ^ n1414 ;
  assign n1435 = n1417 ^ n1337 ;
  assign n1436 = n1435 ^ n1418 ;
  assign n1437 = n1082 & ~n1267 ;
  assign n1438 = n1437 ^ n1269 ;
  assign n1439 = n1188 & ~n1267 ;
  assign n1440 = n1439 ^ n1277 ;
  assign n1441 = n1196 & ~n1267 ;
  assign n1442 = n1441 ^ n1288 ;
  assign n1443 = n1203 & ~n1267 ;
  assign n1444 = n1443 ^ n1296 ;
  assign n1445 = n1212 & ~n1267 ;
  assign n1446 = n1445 ^ n1308 ;
  assign n1447 = n1219 & ~n1267 ;
  assign n1448 = n1447 ^ n1316 ;
  assign n1449 = n1227 & ~n1267 ;
  assign n1450 = n1449 ^ n1327 ;
  assign n1451 = n1235 & ~n1267 ;
  assign n1452 = n1451 ^ n1335 ;
  assign n1454 = n807 & ~n1079 ;
  assign n1453 = n995 & n1079 ;
  assign n1455 = n1454 ^ n1453 ;
  assign n1457 = n999 & ~n1079 ;
  assign n1456 = n1002 & n1079 ;
  assign n1458 = n1457 ^ n1456 ;
  assign n1460 = n1007 & ~n1079 ;
  assign n1459 = n1010 & n1079 ;
  assign n1461 = n1460 ^ n1459 ;
  assign n1463 = n1014 & ~n1079 ;
  assign n1462 = n1017 & n1079 ;
  assign n1464 = n1463 ^ n1462 ;
  assign n1466 = n1023 & ~n1079 ;
  assign n1465 = n1026 & n1079 ;
  assign n1467 = n1466 ^ n1465 ;
  assign n1469 = n1030 & ~n1079 ;
  assign n1468 = n1033 & n1079 ;
  assign n1470 = n1469 ^ n1468 ;
  assign n1472 = n1038 & ~n1079 ;
  assign n1471 = n1041 & n1079 ;
  assign n1473 = n1472 ^ n1471 ;
  assign n1474 = n1046 & ~n1079 ;
  assign n1475 = n1474 ^ n1233 ;
  assign n1477 = n442 & ~n804 ;
  assign n1476 = n721 & n804 ;
  assign n1478 = n1477 ^ n1476 ;
  assign n1480 = n725 & ~n804 ;
  assign n1479 = n728 & n804 ;
  assign n1481 = n1480 ^ n1479 ;
  assign n1483 = n733 & ~n804 ;
  assign n1482 = n736 & n804 ;
  assign n1484 = n1483 ^ n1482 ;
  assign n1486 = n740 & ~n804 ;
  assign n1485 = n743 & n804 ;
  assign n1487 = n1486 ^ n1485 ;
  assign n1489 = n749 & ~n804 ;
  assign n1488 = n752 & n804 ;
  assign n1490 = n1489 ^ n1488 ;
  assign n1492 = n756 & ~n804 ;
  assign n1491 = n759 & n804 ;
  assign n1493 = n1492 ^ n1491 ;
  assign n1495 = n764 & ~n804 ;
  assign n1494 = n767 & n804 ;
  assign n1496 = n1495 ^ n1494 ;
  assign n1497 = n771 & ~n804 ;
  assign n1498 = n1497 ^ n1044 ;
  assign n1500 = x40 & ~n439 ;
  assign n1499 = n368 & n439 ;
  assign n1501 = n1500 ^ n1499 ;
  assign n1503 = x41 & ~n439 ;
  assign n1502 = n372 & n439 ;
  assign n1504 = n1503 ^ n1502 ;
  assign n1506 = x42 & ~n439 ;
  assign n1505 = n377 & n439 ;
  assign n1507 = n1506 ^ n1505 ;
  assign n1509 = x43 & ~n439 ;
  assign n1508 = n381 & n439 ;
  assign n1510 = n1509 ^ n1508 ;
  assign n1512 = x44 & ~n439 ;
  assign n1511 = n387 & n439 ;
  assign n1513 = n1512 ^ n1511 ;
  assign n1515 = x45 & ~n439 ;
  assign n1514 = n391 & n439 ;
  assign n1516 = n1515 ^ n1514 ;
  assign n1518 = x46 & ~n439 ;
  assign n1517 = n396 & n439 ;
  assign n1519 = n1518 ^ n1517 ;
  assign n1521 = x47 & ~n439 ;
  assign n1520 = n400 & n439 ;
  assign n1522 = n1521 ^ n1520 ;
  assign y0 = n1392 ;
  assign y1 = n1396 ;
  assign y2 = n1400 ;
  assign y3 = n1404 ;
  assign y4 = n1408 ;
  assign y5 = n1412 ;
  assign y6 = n1416 ;
  assign y7 = n1420 ;
  assign y8 = n1422 ;
  assign y9 = n1424 ;
  assign y10 = n1426 ;
  assign y11 = n1428 ;
  assign y12 = n1430 ;
  assign y13 = n1432 ;
  assign y14 = n1434 ;
  assign y15 = n1436 ;
  assign y16 = n1438 ;
  assign y17 = n1440 ;
  assign y18 = n1442 ;
  assign y19 = n1444 ;
  assign y20 = n1446 ;
  assign y21 = n1448 ;
  assign y22 = n1450 ;
  assign y23 = n1452 ;
  assign y24 = n1455 ;
  assign y25 = n1458 ;
  assign y26 = n1461 ;
  assign y27 = n1464 ;
  assign y28 = n1467 ;
  assign y29 = n1470 ;
  assign y30 = n1473 ;
  assign y31 = n1475 ;
  assign y32 = n1478 ;
  assign y33 = n1481 ;
  assign y34 = n1484 ;
  assign y35 = n1487 ;
  assign y36 = n1490 ;
  assign y37 = n1493 ;
  assign y38 = n1496 ;
  assign y39 = n1498 ;
  assign y40 = n1501 ;
  assign y41 = n1504 ;
  assign y42 = n1507 ;
  assign y43 = n1510 ;
  assign y44 = n1513 ;
  assign y45 = n1516 ;
  assign y46 = n1519 ;
  assign y47 = n1522 ;
endmodule
