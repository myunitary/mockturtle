module bitonic_sort_inc_1_4 (in_array_0, in_array_1, in_array_2, in_array_3, out_array_0, out_array_1, out_array_2, out_array_3);
input in_array_0, in_array_1, in_array_2, in_array_3;
output out_array_0, out_array_1, out_array_2, out_array_3;
wire _00_, _01_, _02_, _02__neg, _03_, _04_, _05_, _06_, _06__neg, _07_, _08_, _09_, _10_, _11_, _12_, _13_, _14_, _15_, _16_, _16__neg;
assign _16__neg = in_array_1 | in_array_0;
assign _16_ = ~_16__neg;
assign _00_ = ~_16_;
assign _01_ = in_array_3 & in_array_2;
assign _02__neg = _01_ | _16_;
assign _02_ = ~_02__neg;
assign _03_ = _02_ ^ _00_;
assign _04_ = in_array_1 & in_array_0;
assign _05_ = ~_04_;
assign _06__neg = in_array_3 | in_array_2;
assign _06_ = ~_06__neg;
assign _07_ = _06_ & _04_;
assign _08_ = _07_ ^ _05_;
assign _09_ = _08_ & _03_;
assign out_array_3 = _09_ ^ _03_;
assign _10_ = _02_ ^ _01_;
assign _11_ = _07_ ^ _06_;
assign _12_ = _11_ & _10_;
assign out_array_1 = _12_ ^ _10_;
assign _13_ = _07_ ^ _04_;
assign out_array_2 = _09_ ^ _13_;
assign _14_ = ~_06_;
assign _15_ = _07_ ^ _14_;
assign out_array_0 = _12_ ^ _15_;
endmodule
