module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 ;
  assign n192 = x33 ^ x1 ;
  assign n193 = ~x0 & x32 ;
  assign n194 = ~n192 & n193 ;
  assign n191 = ~x1 & x33 ;
  assign n195 = n194 ^ n191 ;
  assign n187 = x35 ^ x3 ;
  assign n196 = x34 ^ x2 ;
  assign n197 = ~n187 & ~n196 ;
  assign n198 = n195 & n197 ;
  assign n188 = ~x2 & x34 ;
  assign n189 = ~n187 & n188 ;
  assign n186 = ~x3 & x35 ;
  assign n190 = n189 ^ n186 ;
  assign n199 = n198 ^ n190 ;
  assign n173 = x39 ^ x7 ;
  assign n177 = x38 ^ x6 ;
  assign n178 = ~n173 & ~n177 ;
  assign n180 = x37 ^ x5 ;
  assign n200 = x36 ^ x4 ;
  assign n201 = ~n180 & ~n200 ;
  assign n202 = n178 & n201 ;
  assign n203 = n199 & n202 ;
  assign n181 = ~x4 & x36 ;
  assign n182 = ~n180 & n181 ;
  assign n179 = ~x5 & x37 ;
  assign n183 = n182 ^ n179 ;
  assign n184 = n178 & n183 ;
  assign n174 = ~x6 & x38 ;
  assign n175 = ~n173 & n174 ;
  assign n172 = ~x7 & x39 ;
  assign n176 = n175 ^ n172 ;
  assign n185 = n184 ^ n176 ;
  assign n204 = n203 ^ n185 ;
  assign n140 = x47 ^ x15 ;
  assign n144 = x46 ^ x14 ;
  assign n145 = ~n140 & ~n144 ;
  assign n147 = x45 ^ x13 ;
  assign n153 = x44 ^ x12 ;
  assign n154 = ~n147 & ~n153 ;
  assign n155 = n145 & n154 ;
  assign n157 = x43 ^ x11 ;
  assign n161 = x42 ^ x10 ;
  assign n162 = ~n157 & ~n161 ;
  assign n164 = x41 ^ x9 ;
  assign n205 = x40 ^ x8 ;
  assign n206 = ~n164 & ~n205 ;
  assign n207 = n162 & n206 ;
  assign n208 = n155 & n207 ;
  assign n209 = n204 & n208 ;
  assign n165 = ~x8 & x40 ;
  assign n166 = ~n164 & n165 ;
  assign n163 = ~x9 & x41 ;
  assign n167 = n166 ^ n163 ;
  assign n168 = n162 & n167 ;
  assign n158 = ~x10 & x42 ;
  assign n159 = ~n157 & n158 ;
  assign n156 = ~x11 & x43 ;
  assign n160 = n159 ^ n156 ;
  assign n169 = n168 ^ n160 ;
  assign n170 = n155 & n169 ;
  assign n148 = ~x12 & x44 ;
  assign n149 = ~n147 & n148 ;
  assign n146 = ~x13 & x45 ;
  assign n150 = n149 ^ n146 ;
  assign n151 = n145 & n150 ;
  assign n141 = ~x14 & x46 ;
  assign n142 = ~n140 & n141 ;
  assign n139 = ~x15 & x47 ;
  assign n143 = n142 ^ n139 ;
  assign n152 = n151 ^ n143 ;
  assign n171 = n170 ^ n152 ;
  assign n210 = n209 ^ n171 ;
  assign n65 = x32 ^ x0 ;
  assign n67 = x63 ^ x31 ;
  assign n71 = x62 ^ x30 ;
  assign n72 = ~n67 & ~n71 ;
  assign n74 = x61 ^ x29 ;
  assign n80 = x60 ^ x28 ;
  assign n81 = ~n74 & ~n80 ;
  assign n82 = n72 & n81 ;
  assign n84 = x59 ^ x27 ;
  assign n88 = x58 ^ x26 ;
  assign n89 = ~n84 & ~n88 ;
  assign n91 = x57 ^ x25 ;
  assign n99 = x56 ^ x24 ;
  assign n100 = ~n91 & ~n99 ;
  assign n101 = n89 & n100 ;
  assign n102 = n82 & n101 ;
  assign n104 = x55 ^ x23 ;
  assign n108 = x54 ^ x22 ;
  assign n109 = ~n104 & ~n108 ;
  assign n111 = x53 ^ x21 ;
  assign n117 = x52 ^ x20 ;
  assign n118 = ~n111 & ~n117 ;
  assign n119 = n109 & n118 ;
  assign n121 = x51 ^ x19 ;
  assign n125 = x50 ^ x18 ;
  assign n126 = ~n121 & ~n125 ;
  assign n128 = x49 ^ x17 ;
  assign n211 = x48 ^ x16 ;
  assign n212 = ~n128 & ~n211 ;
  assign n213 = n126 & n212 ;
  assign n214 = n119 & n213 ;
  assign n215 = n102 & n214 ;
  assign n216 = n65 & n215 ;
  assign n217 = n210 & n216 ;
  assign n129 = ~x16 & x48 ;
  assign n130 = ~n128 & n129 ;
  assign n127 = ~x17 & x49 ;
  assign n131 = n130 ^ n127 ;
  assign n132 = n126 & n131 ;
  assign n122 = ~x18 & x50 ;
  assign n123 = ~n121 & n122 ;
  assign n120 = ~x19 & x51 ;
  assign n124 = n123 ^ n120 ;
  assign n133 = n132 ^ n124 ;
  assign n134 = n119 & n133 ;
  assign n112 = ~x20 & x52 ;
  assign n113 = ~n111 & n112 ;
  assign n110 = ~x21 & x53 ;
  assign n114 = n113 ^ n110 ;
  assign n115 = n109 & n114 ;
  assign n105 = ~x22 & x54 ;
  assign n106 = ~n104 & n105 ;
  assign n103 = ~x23 & x55 ;
  assign n107 = n106 ^ n103 ;
  assign n116 = n115 ^ n107 ;
  assign n135 = n134 ^ n116 ;
  assign n136 = n102 & n135 ;
  assign n92 = ~x24 & x56 ;
  assign n93 = ~n91 & n92 ;
  assign n90 = ~x25 & x57 ;
  assign n94 = n93 ^ n90 ;
  assign n95 = n89 & n94 ;
  assign n85 = ~x26 & x58 ;
  assign n86 = ~n84 & n85 ;
  assign n83 = ~x27 & x59 ;
  assign n87 = n86 ^ n83 ;
  assign n96 = n95 ^ n87 ;
  assign n97 = n82 & n96 ;
  assign n75 = ~x28 & x60 ;
  assign n76 = ~n74 & n75 ;
  assign n73 = ~x29 & x61 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = n72 & n77 ;
  assign n68 = ~x30 & x62 ;
  assign n69 = ~n67 & n68 ;
  assign n66 = ~x31 & x63 ;
  assign n70 = n69 ^ n66 ;
  assign n79 = n78 ^ n70 ;
  assign n98 = n97 ^ n79 ;
  assign n137 = n136 ^ n98 ;
  assign n138 = n65 & n137 ;
  assign n218 = n217 ^ n138 ;
  assign n219 = n218 ^ x32 ;
  assign n221 = n192 & n215 ;
  assign n222 = n210 & n221 ;
  assign n220 = n137 & n192 ;
  assign n223 = n222 ^ n220 ;
  assign n224 = n223 ^ x33 ;
  assign n226 = n196 & n215 ;
  assign n227 = n210 & n226 ;
  assign n225 = n137 & n196 ;
  assign n228 = n227 ^ n225 ;
  assign n229 = n228 ^ x34 ;
  assign n231 = n187 & n215 ;
  assign n232 = n210 & n231 ;
  assign n230 = n137 & n187 ;
  assign n233 = n232 ^ n230 ;
  assign n234 = n233 ^ x35 ;
  assign n236 = n200 & n215 ;
  assign n237 = n210 & n236 ;
  assign n235 = n137 & n200 ;
  assign n238 = n237 ^ n235 ;
  assign n239 = n238 ^ x36 ;
  assign n241 = n180 & n215 ;
  assign n242 = n210 & n241 ;
  assign n240 = n137 & n180 ;
  assign n243 = n242 ^ n240 ;
  assign n244 = n243 ^ x37 ;
  assign n246 = n177 & n215 ;
  assign n247 = n210 & n246 ;
  assign n245 = n137 & n177 ;
  assign n248 = n247 ^ n245 ;
  assign n249 = n248 ^ x38 ;
  assign n251 = n173 & n215 ;
  assign n252 = n210 & n251 ;
  assign n250 = n137 & n173 ;
  assign n253 = n252 ^ n250 ;
  assign n254 = n253 ^ x39 ;
  assign n256 = n205 & n215 ;
  assign n257 = n210 & n256 ;
  assign n255 = n137 & n205 ;
  assign n258 = n257 ^ n255 ;
  assign n259 = n258 ^ x40 ;
  assign n261 = n164 & n215 ;
  assign n262 = n210 & n261 ;
  assign n260 = n137 & n164 ;
  assign n263 = n262 ^ n260 ;
  assign n264 = n263 ^ x41 ;
  assign n266 = n161 & n215 ;
  assign n267 = n210 & n266 ;
  assign n265 = n137 & n161 ;
  assign n268 = n267 ^ n265 ;
  assign n269 = n268 ^ x42 ;
  assign n271 = n157 & n215 ;
  assign n272 = n210 & n271 ;
  assign n270 = n137 & n157 ;
  assign n273 = n272 ^ n270 ;
  assign n274 = n273 ^ x43 ;
  assign n276 = n153 & n215 ;
  assign n277 = n210 & n276 ;
  assign n275 = n137 & n153 ;
  assign n278 = n277 ^ n275 ;
  assign n279 = n278 ^ x44 ;
  assign n281 = n147 & n215 ;
  assign n282 = n210 & n281 ;
  assign n280 = n137 & n147 ;
  assign n283 = n282 ^ n280 ;
  assign n284 = n283 ^ x45 ;
  assign n286 = n144 & n215 ;
  assign n287 = n210 & n286 ;
  assign n285 = n137 & n144 ;
  assign n288 = n287 ^ n285 ;
  assign n289 = n288 ^ x46 ;
  assign n291 = n140 & n215 ;
  assign n292 = n210 & n291 ;
  assign n290 = n137 & n140 ;
  assign n293 = n292 ^ n290 ;
  assign n294 = n293 ^ x47 ;
  assign n296 = n211 & n215 ;
  assign n297 = n210 & n296 ;
  assign n295 = n137 & n211 ;
  assign n298 = n297 ^ n295 ;
  assign n299 = n298 ^ x48 ;
  assign n301 = n128 & n215 ;
  assign n302 = n210 & n301 ;
  assign n300 = n128 & n137 ;
  assign n303 = n302 ^ n300 ;
  assign n304 = n303 ^ x49 ;
  assign n306 = n125 & n215 ;
  assign n307 = n210 & n306 ;
  assign n305 = n125 & n137 ;
  assign n308 = n307 ^ n305 ;
  assign n309 = n308 ^ x50 ;
  assign n311 = n121 & n215 ;
  assign n312 = n210 & n311 ;
  assign n310 = n121 & n137 ;
  assign n313 = n312 ^ n310 ;
  assign n314 = n313 ^ x51 ;
  assign n316 = n117 & n215 ;
  assign n317 = n210 & n316 ;
  assign n315 = n117 & n137 ;
  assign n318 = n317 ^ n315 ;
  assign n319 = n318 ^ x52 ;
  assign n321 = n111 & n215 ;
  assign n322 = n210 & n321 ;
  assign n320 = n111 & n137 ;
  assign n323 = n322 ^ n320 ;
  assign n324 = n323 ^ x53 ;
  assign n326 = n108 & n215 ;
  assign n327 = n210 & n326 ;
  assign n325 = n108 & n137 ;
  assign n328 = n327 ^ n325 ;
  assign n329 = n328 ^ x54 ;
  assign n331 = n104 & n215 ;
  assign n332 = n210 & n331 ;
  assign n330 = n104 & n137 ;
  assign n333 = n332 ^ n330 ;
  assign n334 = n333 ^ x55 ;
  assign n336 = n99 & n215 ;
  assign n337 = n210 & n336 ;
  assign n335 = n99 & n137 ;
  assign n338 = n337 ^ n335 ;
  assign n339 = n338 ^ x56 ;
  assign n341 = n91 & n215 ;
  assign n342 = n210 & n341 ;
  assign n340 = n91 & n137 ;
  assign n343 = n342 ^ n340 ;
  assign n344 = n343 ^ x57 ;
  assign n346 = n88 & n215 ;
  assign n347 = n210 & n346 ;
  assign n345 = n88 & n137 ;
  assign n348 = n347 ^ n345 ;
  assign n349 = n348 ^ x58 ;
  assign n351 = n84 & n215 ;
  assign n352 = n210 & n351 ;
  assign n350 = n84 & n137 ;
  assign n353 = n352 ^ n350 ;
  assign n354 = n353 ^ x59 ;
  assign n356 = n80 & n215 ;
  assign n357 = n210 & n356 ;
  assign n355 = n80 & n137 ;
  assign n358 = n357 ^ n355 ;
  assign n359 = n358 ^ x60 ;
  assign n361 = n74 & n215 ;
  assign n362 = n210 & n361 ;
  assign n360 = n74 & n137 ;
  assign n363 = n362 ^ n360 ;
  assign n364 = n363 ^ x61 ;
  assign n366 = n71 & n215 ;
  assign n367 = n210 & n366 ;
  assign n365 = n71 & n137 ;
  assign n368 = n367 ^ n365 ;
  assign n369 = n368 ^ x62 ;
  assign n371 = n67 & n215 ;
  assign n372 = n210 & n371 ;
  assign n370 = n67 & n137 ;
  assign n373 = n372 ^ n370 ;
  assign n374 = n373 ^ x63 ;
  assign y0 = n219 ;
  assign y1 = n224 ;
  assign y2 = n229 ;
  assign y3 = n234 ;
  assign y4 = n239 ;
  assign y5 = n244 ;
  assign y6 = n249 ;
  assign y7 = n254 ;
  assign y8 = n259 ;
  assign y9 = n264 ;
  assign y10 = n269 ;
  assign y11 = n274 ;
  assign y12 = n279 ;
  assign y13 = n284 ;
  assign y14 = n289 ;
  assign y15 = n294 ;
  assign y16 = n299 ;
  assign y17 = n304 ;
  assign y18 = n309 ;
  assign y19 = n314 ;
  assign y20 = n319 ;
  assign y21 = n324 ;
  assign y22 = n329 ;
  assign y23 = n334 ;
  assign y24 = n339 ;
  assign y25 = n344 ;
  assign y26 = n349 ;
  assign y27 = n354 ;
  assign y28 = n359 ;
  assign y29 = n364 ;
  assign y30 = n369 ;
  assign y31 = n374 ;
endmodule
