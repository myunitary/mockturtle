module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 ;
  assign n33 = ~x0 & x1 ;
  assign n34 = ~x0 & ~x1 ;
  assign n35 = x2 & n34 ;
  assign n36 = ~x2 & x3 ;
  assign n37 = n34 & n36 ;
  assign n38 = ~x2 & ~x3 ;
  assign n39 = n34 & n38 ;
  assign n40 = x4 & n39 ;
  assign n41 = ~x4 & x5 ;
  assign n42 = n39 & n41 ;
  assign n43 = ~x4 & ~x5 ;
  assign n44 = n39 & n43 ;
  assign n45 = x6 & n44 ;
  assign n46 = ~x6 & x7 ;
  assign n47 = n44 & n46 ;
  assign n48 = ~x6 & ~x7 ;
  assign n49 = n43 & n48 ;
  assign n50 = n39 & n49 ;
  assign n51 = x8 & n50 ;
  assign n52 = ~x8 & x9 ;
  assign n53 = n50 & n52 ;
  assign n54 = ~x8 & ~x9 ;
  assign n55 = n50 & n54 ;
  assign n56 = x10 & n55 ;
  assign n57 = ~x10 & x11 ;
  assign n58 = n55 & n57 ;
  assign n59 = ~x10 & ~x11 ;
  assign n60 = n54 & n59 ;
  assign n61 = n50 & n60 ;
  assign n62 = x12 & n61 ;
  assign n63 = ~x12 & x13 ;
  assign n64 = n61 & n63 ;
  assign n65 = ~x12 & ~x13 ;
  assign n66 = x14 & n65 ;
  assign n67 = n61 & n66 ;
  assign n68 = ~x14 & x15 ;
  assign n69 = n65 & n68 ;
  assign n70 = n61 & n69 ;
  assign n71 = ~x14 & ~x15 ;
  assign n72 = n65 & n71 ;
  assign n73 = n60 & n72 ;
  assign n74 = n50 & n73 ;
  assign n75 = x16 & n74 ;
  assign n76 = ~x16 & x17 ;
  assign n77 = n74 & n76 ;
  assign n78 = ~x16 & ~x17 ;
  assign n79 = x18 & n78 ;
  assign n80 = n74 & n79 ;
  assign n81 = ~x18 & n78 ;
  assign n82 = x19 & n81 ;
  assign n83 = n74 & n82 ;
  assign n84 = ~x18 & ~x19 ;
  assign n85 = n78 & n84 ;
  assign n86 = x20 & n85 ;
  assign n87 = n74 & n86 ;
  assign n88 = ~x20 & x21 ;
  assign n89 = n85 & n88 ;
  assign n90 = n74 & n89 ;
  assign n91 = ~x20 & ~x21 ;
  assign n92 = x22 & n91 ;
  assign n93 = n85 & n92 ;
  assign n94 = n74 & n93 ;
  assign n95 = ~x22 & n91 ;
  assign n96 = x23 & n95 ;
  assign n97 = n85 & n96 ;
  assign n98 = n74 & n97 ;
  assign n99 = ~x22 & ~x23 ;
  assign n100 = n91 & n99 ;
  assign n101 = n85 & n100 ;
  assign n102 = x24 & n101 ;
  assign n103 = n74 & n102 ;
  assign n104 = ~x24 & x25 ;
  assign n105 = n101 & n104 ;
  assign n106 = n74 & n105 ;
  assign n107 = ~x24 & ~x25 ;
  assign n108 = x26 & n107 ;
  assign n109 = n101 & n108 ;
  assign n110 = n74 & n109 ;
  assign n111 = ~x26 & n107 ;
  assign n112 = x27 & n111 ;
  assign n113 = n101 & n112 ;
  assign n114 = n74 & n113 ;
  assign n115 = ~x26 & ~x27 ;
  assign n116 = n107 & n115 ;
  assign n117 = x28 & n116 ;
  assign n118 = n101 & n117 ;
  assign n119 = n74 & n118 ;
  assign n120 = ~x28 & x29 ;
  assign n121 = n116 & n120 ;
  assign n122 = n101 & n121 ;
  assign n123 = n74 & n122 ;
  assign n124 = ~x29 & x30 ;
  assign n125 = ~x28 & n124 ;
  assign n126 = n116 & n125 ;
  assign n127 = n101 & n126 ;
  assign n128 = n74 & n127 ;
  assign n129 = ~x29 & ~x30 ;
  assign n130 = ~x28 & x31 ;
  assign n131 = n129 & n130 ;
  assign n132 = n116 & n131 ;
  assign n133 = n101 & n132 ;
  assign n134 = n74 & n133 ;
  assign y0 = x0 ;
  assign y1 = n33 ;
  assign y2 = n35 ;
  assign y3 = n37 ;
  assign y4 = n40 ;
  assign y5 = n42 ;
  assign y6 = n45 ;
  assign y7 = n47 ;
  assign y8 = n51 ;
  assign y9 = n53 ;
  assign y10 = n56 ;
  assign y11 = n58 ;
  assign y12 = n62 ;
  assign y13 = n64 ;
  assign y14 = n67 ;
  assign y15 = n70 ;
  assign y16 = n75 ;
  assign y17 = n77 ;
  assign y18 = n80 ;
  assign y19 = n83 ;
  assign y20 = n87 ;
  assign y21 = n90 ;
  assign y22 = n94 ;
  assign y23 = n98 ;
  assign y24 = n103 ;
  assign y25 = n106 ;
  assign y26 = n110 ;
  assign y27 = n114 ;
  assign y28 = n119 ;
  assign y29 = n123 ;
  assign y30 = n128 ;
  assign y31 = n134 ;
endmodule
