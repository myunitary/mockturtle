// Benchmark "/tmp/tmp" written by ABC on Wed Nov 12 17:45:18 2025

module multiplier_opt ( 
    n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
    n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127  );
  input  n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
    n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
    n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127;
  wire new_n129, new_n130, new_n131, new_n132, new_n133, new_n134, new_n135,
    new_n136, new_n137, new_n138, new_n139, new_n140, new_n141, new_n142,
    new_n143, new_n144, new_n145, new_n146, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n182, new_n183, new_n184,
    new_n185, new_n186, new_n187, new_n188, new_n189, new_n190, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510, new_n1511, new_n1512,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1564, new_n1565, new_n1566,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1584,
    new_n1585, new_n1586, new_n1587, new_n1588, new_n1589, new_n1590,
    new_n1591, new_n1592, new_n1593, new_n1594, new_n1595, new_n1596,
    new_n1597, new_n1598, new_n1599, new_n1600, new_n1601, new_n1602,
    new_n1603, new_n1604, new_n1605, new_n1606, new_n1607, new_n1608,
    new_n1609, new_n1610, new_n1611, new_n1612, new_n1613, new_n1614,
    new_n1615, new_n1616, new_n1617, new_n1618, new_n1619, new_n1620,
    new_n1621, new_n1622, new_n1623, new_n1624, new_n1625, new_n1626,
    new_n1627, new_n1628, new_n1629, new_n1630, new_n1631, new_n1632,
    new_n1633, new_n1634, new_n1635, new_n1636, new_n1637, new_n1638,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1644,
    new_n1645, new_n1646, new_n1647, new_n1648, new_n1649, new_n1650,
    new_n1651, new_n1652, new_n1653, new_n1654, new_n1655, new_n1656,
    new_n1657, new_n1658, new_n1659, new_n1660, new_n1661, new_n1662,
    new_n1663, new_n1664, new_n1665, new_n1666, new_n1667, new_n1668,
    new_n1669, new_n1670, new_n1671, new_n1672, new_n1673, new_n1674,
    new_n1675, new_n1676, new_n1677, new_n1678, new_n1679, new_n1680,
    new_n1681, new_n1682, new_n1683, new_n1684, new_n1685, new_n1686,
    new_n1687, new_n1688, new_n1689, new_n1690, new_n1691, new_n1692,
    new_n1693, new_n1694, new_n1695, new_n1696, new_n1697, new_n1698,
    new_n1699, new_n1700, new_n1701, new_n1702, new_n1703, new_n1704,
    new_n1705, new_n1706, new_n1707, new_n1708, new_n1709, new_n1710,
    new_n1711, new_n1712, new_n1713, new_n1714, new_n1715, new_n1716,
    new_n1717, new_n1718, new_n1719, new_n1720, new_n1721, new_n1722,
    new_n1723, new_n1724, new_n1725, new_n1726, new_n1727, new_n1728,
    new_n1729, new_n1730, new_n1731, new_n1732, new_n1733, new_n1734,
    new_n1735, new_n1736, new_n1737, new_n1738, new_n1739, new_n1740,
    new_n1741, new_n1742, new_n1743, new_n1744, new_n1745, new_n1746,
    new_n1747, new_n1748, new_n1749, new_n1750, new_n1751, new_n1752,
    new_n1753, new_n1754, new_n1755, new_n1756, new_n1757, new_n1758,
    new_n1759, new_n1760, new_n1761, new_n1762, new_n1763, new_n1764,
    new_n1765, new_n1766, new_n1767, new_n1768, new_n1769, new_n1770,
    new_n1771, new_n1772, new_n1773, new_n1774, new_n1775, new_n1776,
    new_n1777, new_n1778, new_n1779, new_n1780, new_n1781, new_n1782,
    new_n1783, new_n1784, new_n1785, new_n1786, new_n1787, new_n1788,
    new_n1789, new_n1790, new_n1791, new_n1792, new_n1793, new_n1794,
    new_n1795, new_n1796, new_n1797, new_n1798, new_n1799, new_n1800,
    new_n1801, new_n1802, new_n1803, new_n1804, new_n1805, new_n1806,
    new_n1807, new_n1808, new_n1809, new_n1810, new_n1811, new_n1812,
    new_n1813, new_n1814, new_n1815, new_n1816, new_n1817, new_n1818,
    new_n1819, new_n1820, new_n1821, new_n1822, new_n1823, new_n1824,
    new_n1825, new_n1826, new_n1827, new_n1828, new_n1829, new_n1830,
    new_n1831, new_n1832, new_n1833, new_n1834, new_n1835, new_n1836,
    new_n1837, new_n1838, new_n1839, new_n1840, new_n1841, new_n1842,
    new_n1843, new_n1844, new_n1845, new_n1846, new_n1847, new_n1848,
    new_n1849, new_n1850, new_n1851, new_n1852, new_n1853, new_n1854,
    new_n1855, new_n1856, new_n1857, new_n1858, new_n1859, new_n1860,
    new_n1861, new_n1862, new_n1863, new_n1864, new_n1865, new_n1866,
    new_n1867, new_n1868, new_n1869, new_n1870, new_n1871, new_n1872,
    new_n1873, new_n1874, new_n1875, new_n1876, new_n1877, new_n1878,
    new_n1879, new_n1880, new_n1881, new_n1882, new_n1883, new_n1884,
    new_n1885, new_n1886, new_n1887, new_n1888, new_n1889, new_n1890,
    new_n1891, new_n1892, new_n1893, new_n1894, new_n1895, new_n1896,
    new_n1897, new_n1898, new_n1899, new_n1900, new_n1901, new_n1902,
    new_n1903, new_n1904, new_n1905, new_n1906, new_n1907, new_n1908,
    new_n1909, new_n1910, new_n1911, new_n1912, new_n1913, new_n1914,
    new_n1915, new_n1916, new_n1917, new_n1918, new_n1919, new_n1920,
    new_n1921, new_n1922, new_n1923, new_n1924, new_n1925, new_n1926,
    new_n1927, new_n1928, new_n1929, new_n1930, new_n1931, new_n1932,
    new_n1933, new_n1934, new_n1935, new_n1936, new_n1937, new_n1938,
    new_n1939, new_n1940, new_n1941, new_n1942, new_n1943, new_n1944,
    new_n1945, new_n1946, new_n1947, new_n1948, new_n1949, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986,
    new_n1987, new_n1988, new_n1989, new_n1990, new_n1991, new_n1992,
    new_n1993, new_n1994, new_n1995, new_n1996, new_n1997, new_n1998,
    new_n1999, new_n2000, new_n2001, new_n2002, new_n2003, new_n2004,
    new_n2005, new_n2006, new_n2007, new_n2008, new_n2009, new_n2010,
    new_n2011, new_n2012, new_n2013, new_n2014, new_n2015, new_n2016,
    new_n2017, new_n2018, new_n2019, new_n2020, new_n2021, new_n2022,
    new_n2023, new_n2024, new_n2025, new_n2026, new_n2027, new_n2028,
    new_n2029, new_n2030, new_n2031, new_n2032, new_n2033, new_n2034,
    new_n2035, new_n2036, new_n2037, new_n2038, new_n2039, new_n2040,
    new_n2041, new_n2042, new_n2043, new_n2044, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058,
    new_n2059, new_n2060, new_n2061, new_n2062, new_n2063, new_n2064,
    new_n2065, new_n2066, new_n2067, new_n2068, new_n2069, new_n2070,
    new_n2071, new_n2072, new_n2073, new_n2074, new_n2075, new_n2076,
    new_n2077, new_n2078, new_n2079, new_n2080, new_n2081, new_n2082,
    new_n2083, new_n2084, new_n2085, new_n2086, new_n2087, new_n2088,
    new_n2089, new_n2090, new_n2091, new_n2092, new_n2093, new_n2094,
    new_n2095, new_n2096, new_n2097, new_n2098, new_n2099, new_n2100,
    new_n2101, new_n2102, new_n2103, new_n2104, new_n2105, new_n2106,
    new_n2107, new_n2108, new_n2109, new_n2110, new_n2111, new_n2112,
    new_n2113, new_n2114, new_n2115, new_n2116, new_n2117, new_n2118,
    new_n2119, new_n2120, new_n2121, new_n2122, new_n2123, new_n2124,
    new_n2125, new_n2126, new_n2127, new_n2128, new_n2129, new_n2130,
    new_n2131, new_n2132, new_n2133, new_n2134, new_n2135, new_n2136,
    new_n2137, new_n2138, new_n2139, new_n2140, new_n2141, new_n2142,
    new_n2143, new_n2144, new_n2145, new_n2146, new_n2147, new_n2148,
    new_n2149, new_n2150, new_n2151, new_n2152, new_n2153, new_n2154,
    new_n2155, new_n2156, new_n2157, new_n2158, new_n2159, new_n2160,
    new_n2161, new_n2162, new_n2163, new_n2164, new_n2165, new_n2166,
    new_n2167, new_n2168, new_n2169, new_n2170, new_n2171, new_n2172,
    new_n2173, new_n2174, new_n2175, new_n2176, new_n2177, new_n2178,
    new_n2179, new_n2180, new_n2181, new_n2182, new_n2183, new_n2184,
    new_n2185, new_n2186, new_n2187, new_n2188, new_n2189, new_n2190,
    new_n2191, new_n2192, new_n2193, new_n2194, new_n2195, new_n2196,
    new_n2197, new_n2198, new_n2199, new_n2200, new_n2201, new_n2202,
    new_n2203, new_n2204, new_n2205, new_n2206, new_n2207, new_n2208,
    new_n2209, new_n2210, new_n2211, new_n2212, new_n2213, new_n2214,
    new_n2215, new_n2216, new_n2217, new_n2218, new_n2219, new_n2220,
    new_n2221, new_n2222, new_n2223, new_n2224, new_n2225, new_n2226,
    new_n2227, new_n2228, new_n2229, new_n2230, new_n2231, new_n2232,
    new_n2233, new_n2234, new_n2235, new_n2236, new_n2237, new_n2238,
    new_n2239, new_n2240, new_n2241, new_n2242, new_n2243, new_n2244,
    new_n2245, new_n2246, new_n2247, new_n2248, new_n2249, new_n2250,
    new_n2251, new_n2252, new_n2253, new_n2254, new_n2255, new_n2256,
    new_n2257, new_n2258, new_n2259, new_n2260, new_n2261, new_n2262,
    new_n2263, new_n2264, new_n2265, new_n2266, new_n2267, new_n2268,
    new_n2269, new_n2270, new_n2271, new_n2272, new_n2273, new_n2274,
    new_n2275, new_n2276, new_n2277, new_n2278, new_n2279, new_n2280,
    new_n2281, new_n2282, new_n2283, new_n2284, new_n2285, new_n2286,
    new_n2287, new_n2288, new_n2289, new_n2290, new_n2291, new_n2292,
    new_n2293, new_n2294, new_n2295, new_n2296, new_n2297, new_n2298,
    new_n2299, new_n2300, new_n2301, new_n2302, new_n2303, new_n2304,
    new_n2305, new_n2306, new_n2307, new_n2308, new_n2309, new_n2310,
    new_n2311, new_n2312, new_n2313, new_n2314, new_n2315, new_n2316,
    new_n2317, new_n2318, new_n2319, new_n2320, new_n2321, new_n2322,
    new_n2323, new_n2324, new_n2325, new_n2326, new_n2327, new_n2328,
    new_n2329, new_n2330, new_n2331, new_n2332, new_n2333, new_n2334,
    new_n2335, new_n2336, new_n2337, new_n2338, new_n2339, new_n2340,
    new_n2341, new_n2342, new_n2343, new_n2344, new_n2345, new_n2346,
    new_n2347, new_n2348, new_n2349, new_n2350, new_n2351, new_n2352,
    new_n2353, new_n2354, new_n2355, new_n2356, new_n2357, new_n2358,
    new_n2359, new_n2360, new_n2361, new_n2362, new_n2363, new_n2364,
    new_n2365, new_n2366, new_n2367, new_n2368, new_n2369, new_n2370,
    new_n2371, new_n2372, new_n2373, new_n2374, new_n2375, new_n2376,
    new_n2377, new_n2378, new_n2379, new_n2380, new_n2381, new_n2382,
    new_n2383, new_n2384, new_n2385, new_n2386, new_n2387, new_n2388,
    new_n2389, new_n2390, new_n2391, new_n2392, new_n2393, new_n2394,
    new_n2395, new_n2396, new_n2397, new_n2398, new_n2399, new_n2400,
    new_n2401, new_n2402, new_n2403, new_n2404, new_n2405, new_n2406,
    new_n2407, new_n2408, new_n2409, new_n2410, new_n2411, new_n2412,
    new_n2413, new_n2414, new_n2415, new_n2416, new_n2417, new_n2418,
    new_n2419, new_n2420, new_n2421, new_n2422, new_n2423, new_n2424,
    new_n2425, new_n2426, new_n2427, new_n2428, new_n2429, new_n2430,
    new_n2431, new_n2432, new_n2433, new_n2434, new_n2435, new_n2436,
    new_n2437, new_n2438, new_n2439, new_n2440, new_n2441, new_n2442,
    new_n2443, new_n2444, new_n2445, new_n2446, new_n2447, new_n2448,
    new_n2449, new_n2450, new_n2451, new_n2452, new_n2453, new_n2454,
    new_n2455, new_n2456, new_n2457, new_n2458, new_n2459, new_n2460,
    new_n2461, new_n2462, new_n2463, new_n2464, new_n2465, new_n2466,
    new_n2467, new_n2468, new_n2469, new_n2470, new_n2471, new_n2472,
    new_n2473, new_n2474, new_n2475, new_n2476, new_n2477, new_n2478,
    new_n2479, new_n2480, new_n2481, new_n2482, new_n2483, new_n2484,
    new_n2485, new_n2486, new_n2487, new_n2488, new_n2489, new_n2490,
    new_n2491, new_n2492, new_n2493, new_n2494, new_n2495, new_n2496,
    new_n2497, new_n2498, new_n2499, new_n2500, new_n2501, new_n2502,
    new_n2503, new_n2504, new_n2505, new_n2506, new_n2507, new_n2508,
    new_n2509, new_n2510, new_n2511, new_n2512, new_n2513, new_n2514,
    new_n2515, new_n2516, new_n2517, new_n2518, new_n2519, new_n2520,
    new_n2521, new_n2522, new_n2523, new_n2524, new_n2525, new_n2526,
    new_n2527, new_n2528, new_n2529, new_n2530, new_n2531, new_n2532,
    new_n2533, new_n2534, new_n2535, new_n2536, new_n2537, new_n2538,
    new_n2539, new_n2540, new_n2541, new_n2542, new_n2543, new_n2544,
    new_n2545, new_n2546, new_n2547, new_n2548, new_n2549, new_n2550,
    new_n2551, new_n2552, new_n2553, new_n2554, new_n2555, new_n2556,
    new_n2557, new_n2558, new_n2559, new_n2560, new_n2561, new_n2562,
    new_n2563, new_n2564, new_n2565, new_n2566, new_n2567, new_n2568,
    new_n2569, new_n2570, new_n2571, new_n2572, new_n2573, new_n2574,
    new_n2575, new_n2576, new_n2577, new_n2578, new_n2579, new_n2580,
    new_n2581, new_n2582, new_n2583, new_n2584, new_n2585, new_n2586,
    new_n2587, new_n2588, new_n2589, new_n2590, new_n2591, new_n2592,
    new_n2593, new_n2594, new_n2595, new_n2596, new_n2597, new_n2598,
    new_n2599, new_n2600, new_n2601, new_n2602, new_n2603, new_n2604,
    new_n2605, new_n2606, new_n2607, new_n2608, new_n2609, new_n2610,
    new_n2611, new_n2612, new_n2613, new_n2614, new_n2615, new_n2616,
    new_n2617, new_n2618, new_n2619, new_n2620, new_n2621, new_n2622,
    new_n2623, new_n2624, new_n2625, new_n2626, new_n2627, new_n2628,
    new_n2629, new_n2630, new_n2631, new_n2632, new_n2633, new_n2634,
    new_n2635, new_n2636, new_n2637, new_n2638, new_n2639, new_n2640,
    new_n2641, new_n2642, new_n2643, new_n2644, new_n2645, new_n2646,
    new_n2647, new_n2648, new_n2649, new_n2650, new_n2651, new_n2652,
    new_n2653, new_n2654, new_n2655, new_n2656, new_n2657, new_n2658,
    new_n2659, new_n2660, new_n2661, new_n2662, new_n2663, new_n2664,
    new_n2665, new_n2666, new_n2667, new_n2668, new_n2669, new_n2670,
    new_n2671, new_n2672, new_n2673, new_n2674, new_n2675, new_n2676,
    new_n2677, new_n2678, new_n2679, new_n2680, new_n2681, new_n2682,
    new_n2683, new_n2684, new_n2685, new_n2686, new_n2687, new_n2688,
    new_n2689, new_n2690, new_n2691, new_n2692, new_n2693, new_n2694,
    new_n2695, new_n2696, new_n2697, new_n2698, new_n2699, new_n2700,
    new_n2701, new_n2702, new_n2703, new_n2704, new_n2705, new_n2706,
    new_n2707, new_n2708, new_n2709, new_n2710, new_n2711, new_n2712,
    new_n2713, new_n2714, new_n2715, new_n2716, new_n2717, new_n2718,
    new_n2719, new_n2720, new_n2721, new_n2722, new_n2723, new_n2724,
    new_n2725, new_n2726, new_n2727, new_n2728, new_n2729, new_n2730,
    new_n2731, new_n2732, new_n2733, new_n2734, new_n2735, new_n2736,
    new_n2737, new_n2738, new_n2739, new_n2740, new_n2741, new_n2742,
    new_n2743, new_n2744, new_n2745, new_n2746, new_n2747, new_n2748,
    new_n2749, new_n2750, new_n2751, new_n2752, new_n2753, new_n2754,
    new_n2755, new_n2756, new_n2757, new_n2758, new_n2759, new_n2760,
    new_n2761, new_n2762, new_n2763, new_n2764, new_n2765, new_n2766,
    new_n2767, new_n2768, new_n2769, new_n2770, new_n2771, new_n2772,
    new_n2773, new_n2774, new_n2775, new_n2776, new_n2777, new_n2778,
    new_n2779, new_n2780, new_n2781, new_n2782, new_n2783, new_n2784,
    new_n2785, new_n2786, new_n2787, new_n2788, new_n2789, new_n2790,
    new_n2791, new_n2792, new_n2793, new_n2794, new_n2795, new_n2796,
    new_n2797, new_n2798, new_n2799, new_n2800, new_n2801, new_n2802,
    new_n2803, new_n2804, new_n2805, new_n2806, new_n2807, new_n2808,
    new_n2809, new_n2810, new_n2811, new_n2812, new_n2813, new_n2814,
    new_n2815, new_n2816, new_n2817, new_n2818, new_n2819, new_n2820,
    new_n2821, new_n2822, new_n2823, new_n2824, new_n2825, new_n2826,
    new_n2827, new_n2828, new_n2829, new_n2830, new_n2831, new_n2832,
    new_n2833, new_n2834, new_n2835, new_n2836, new_n2837, new_n2838,
    new_n2839, new_n2840, new_n2841, new_n2842, new_n2843, new_n2844,
    new_n2845, new_n2846, new_n2847, new_n2848, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2853, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858, new_n2859, new_n2860, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874,
    new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886,
    new_n2887, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944, new_n2945, new_n2946,
    new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978, new_n2979, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017, new_n3018,
    new_n3019, new_n3020, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125, new_n3126,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156,
    new_n3157, new_n3158, new_n3159, new_n3160, new_n3161, new_n3162,
    new_n3163, new_n3164, new_n3165, new_n3166, new_n3167, new_n3168,
    new_n3169, new_n3170, new_n3171, new_n3172, new_n3173, new_n3174,
    new_n3175, new_n3176, new_n3177, new_n3178, new_n3179, new_n3180,
    new_n3181, new_n3182, new_n3183, new_n3184, new_n3185, new_n3186,
    new_n3187, new_n3188, new_n3189, new_n3190, new_n3191, new_n3192,
    new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198,
    new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204,
    new_n3205, new_n3206, new_n3207, new_n3208, new_n3209, new_n3210,
    new_n3211, new_n3212, new_n3213, new_n3214, new_n3215, new_n3216,
    new_n3217, new_n3218, new_n3219, new_n3220, new_n3221, new_n3222,
    new_n3223, new_n3224, new_n3225, new_n3226, new_n3227, new_n3228,
    new_n3229, new_n3230, new_n3231, new_n3232, new_n3233, new_n3234,
    new_n3235, new_n3236, new_n3237, new_n3238, new_n3239, new_n3240,
    new_n3241, new_n3242, new_n3243, new_n3244, new_n3245, new_n3246,
    new_n3247, new_n3248, new_n3249, new_n3250, new_n3251, new_n3252,
    new_n3253, new_n3254, new_n3255, new_n3256, new_n3257, new_n3258,
    new_n3259, new_n3260, new_n3261, new_n3262, new_n3263, new_n3264,
    new_n3265, new_n3266, new_n3267, new_n3268, new_n3269, new_n3270,
    new_n3271, new_n3272, new_n3273, new_n3274, new_n3275, new_n3276,
    new_n3277, new_n3278, new_n3279, new_n3280, new_n3281, new_n3282,
    new_n3283, new_n3284, new_n3285, new_n3286, new_n3287, new_n3288,
    new_n3289, new_n3290, new_n3291, new_n3292, new_n3293, new_n3294,
    new_n3295, new_n3296, new_n3297, new_n3298, new_n3299, new_n3300,
    new_n3301, new_n3302, new_n3303, new_n3304, new_n3305, new_n3306,
    new_n3307, new_n3308, new_n3309, new_n3310, new_n3311, new_n3312,
    new_n3313, new_n3314, new_n3315, new_n3316, new_n3317, new_n3318,
    new_n3319, new_n3320, new_n3321, new_n3322, new_n3323, new_n3324,
    new_n3325, new_n3326, new_n3327, new_n3328, new_n3329, new_n3330,
    new_n3331, new_n3332, new_n3333, new_n3334, new_n3335, new_n3336,
    new_n3337, new_n3338, new_n3339, new_n3340, new_n3341, new_n3342,
    new_n3343, new_n3344, new_n3345, new_n3346, new_n3347, new_n3348,
    new_n3349, new_n3350, new_n3351, new_n3352, new_n3353, new_n3354,
    new_n3355, new_n3356, new_n3357, new_n3358, new_n3359, new_n3360,
    new_n3361, new_n3362, new_n3363, new_n3364, new_n3365, new_n3366,
    new_n3367, new_n3368, new_n3369, new_n3370, new_n3371, new_n3372,
    new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378,
    new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384,
    new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390,
    new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396,
    new_n3397, new_n3398, new_n3399, new_n3400, new_n3401, new_n3402,
    new_n3403, new_n3404, new_n3405, new_n3406, new_n3407, new_n3408,
    new_n3409, new_n3410, new_n3411, new_n3412, new_n3413, new_n3414,
    new_n3415, new_n3416, new_n3417, new_n3418, new_n3419, new_n3420,
    new_n3421, new_n3422, new_n3423, new_n3424, new_n3425, new_n3426,
    new_n3427, new_n3428, new_n3429, new_n3430, new_n3431, new_n3432,
    new_n3433, new_n3434, new_n3435, new_n3436, new_n3437, new_n3438,
    new_n3439, new_n3440, new_n3441, new_n3442, new_n3443, new_n3444,
    new_n3445, new_n3446, new_n3447, new_n3448, new_n3449, new_n3450,
    new_n3451, new_n3452, new_n3453, new_n3454, new_n3455, new_n3456,
    new_n3457, new_n3458, new_n3459, new_n3460, new_n3461, new_n3462,
    new_n3463, new_n3464, new_n3465, new_n3466, new_n3467, new_n3468,
    new_n3469, new_n3470, new_n3471, new_n3472, new_n3473, new_n3474,
    new_n3475, new_n3476, new_n3477, new_n3478, new_n3479, new_n3480,
    new_n3481, new_n3482, new_n3483, new_n3484, new_n3485, new_n3486,
    new_n3487, new_n3488, new_n3489, new_n3490, new_n3491, new_n3492,
    new_n3493, new_n3494, new_n3495, new_n3496, new_n3497, new_n3498,
    new_n3499, new_n3500, new_n3501, new_n3502, new_n3503, new_n3504,
    new_n3505, new_n3506, new_n3507, new_n3508, new_n3509, new_n3510,
    new_n3511, new_n3512, new_n3513, new_n3514, new_n3515, new_n3516,
    new_n3517, new_n3518, new_n3519, new_n3520, new_n3521, new_n3522,
    new_n3523, new_n3524, new_n3525, new_n3526, new_n3527, new_n3528,
    new_n3529, new_n3530, new_n3531, new_n3532, new_n3533, new_n3534,
    new_n3535, new_n3536, new_n3537, new_n3538, new_n3539, new_n3540,
    new_n3541, new_n3542, new_n3543, new_n3544, new_n3545, new_n3546,
    new_n3547, new_n3548, new_n3549, new_n3550, new_n3551, new_n3552,
    new_n3553, new_n3554, new_n3555, new_n3556, new_n3557, new_n3558,
    new_n3559, new_n3560, new_n3561, new_n3562, new_n3563, new_n3564,
    new_n3565, new_n3566, new_n3567, new_n3568, new_n3569, new_n3570,
    new_n3571, new_n3572, new_n3573, new_n3574, new_n3575, new_n3576,
    new_n3577, new_n3578, new_n3579, new_n3580, new_n3581, new_n3582,
    new_n3583, new_n3584, new_n3585, new_n3586, new_n3587, new_n3588,
    new_n3589, new_n3590, new_n3591, new_n3592, new_n3593, new_n3594,
    new_n3595, new_n3596, new_n3597, new_n3598, new_n3599, new_n3600,
    new_n3601, new_n3602, new_n3603, new_n3604, new_n3605, new_n3606,
    new_n3607, new_n3608, new_n3609, new_n3610, new_n3611, new_n3612,
    new_n3613, new_n3614, new_n3615, new_n3616, new_n3617, new_n3618,
    new_n3619, new_n3620, new_n3621, new_n3622, new_n3623, new_n3624,
    new_n3625, new_n3626, new_n3627, new_n3628, new_n3629, new_n3630,
    new_n3631, new_n3632, new_n3633, new_n3634, new_n3635, new_n3636,
    new_n3637, new_n3638, new_n3639, new_n3640, new_n3641, new_n3642,
    new_n3643, new_n3644, new_n3645, new_n3646, new_n3647, new_n3648,
    new_n3649, new_n3650, new_n3651, new_n3652, new_n3653, new_n3654,
    new_n3655, new_n3656, new_n3657, new_n3658, new_n3659, new_n3660,
    new_n3661, new_n3662, new_n3663, new_n3664, new_n3665, new_n3666,
    new_n3667, new_n3668, new_n3669, new_n3670, new_n3671, new_n3672,
    new_n3673, new_n3674, new_n3675, new_n3676, new_n3677, new_n3678,
    new_n3679, new_n3680, new_n3681, new_n3682, new_n3683, new_n3684,
    new_n3685, new_n3686, new_n3687, new_n3688, new_n3689, new_n3690,
    new_n3691, new_n3692, new_n3693, new_n3694, new_n3695, new_n3696,
    new_n3697, new_n3698, new_n3699, new_n3700, new_n3701, new_n3702,
    new_n3703, new_n3704, new_n3705, new_n3706, new_n3707, new_n3708,
    new_n3709, new_n3710, new_n3711, new_n3712, new_n3713, new_n3714,
    new_n3715, new_n3716, new_n3717, new_n3718, new_n3719, new_n3720,
    new_n3721, new_n3722, new_n3723, new_n3724, new_n3725, new_n3726,
    new_n3727, new_n3728, new_n3729, new_n3730, new_n3731, new_n3732,
    new_n3733, new_n3734, new_n3735, new_n3736, new_n3737, new_n3738,
    new_n3739, new_n3740, new_n3741, new_n3742, new_n3743, new_n3744,
    new_n3745, new_n3746, new_n3747, new_n3748, new_n3749, new_n3750,
    new_n3751, new_n3752, new_n3753, new_n3754, new_n3755, new_n3756,
    new_n3757, new_n3758, new_n3759, new_n3760, new_n3761, new_n3762,
    new_n3763, new_n3764, new_n3765, new_n3766, new_n3767, new_n3768,
    new_n3769, new_n3770, new_n3771, new_n3772, new_n3773, new_n3774,
    new_n3775, new_n3776, new_n3777, new_n3778, new_n3779, new_n3780,
    new_n3781, new_n3782, new_n3783, new_n3784, new_n3785, new_n3786,
    new_n3787, new_n3788, new_n3789, new_n3790, new_n3791, new_n3792,
    new_n3793, new_n3794, new_n3795, new_n3796, new_n3797, new_n3798,
    new_n3799, new_n3800, new_n3801, new_n3802, new_n3803, new_n3804,
    new_n3805, new_n3806, new_n3807, new_n3808, new_n3809, new_n3810,
    new_n3811, new_n3812, new_n3813, new_n3814, new_n3815, new_n3816,
    new_n3817, new_n3818, new_n3819, new_n3820, new_n3821, new_n3822,
    new_n3823, new_n3824, new_n3825, new_n3826, new_n3827, new_n3828,
    new_n3829, new_n3830, new_n3831, new_n3832, new_n3833, new_n3834,
    new_n3835, new_n3836, new_n3837, new_n3838, new_n3839, new_n3840,
    new_n3841, new_n3842, new_n3843, new_n3844, new_n3845, new_n3846,
    new_n3847, new_n3848, new_n3849, new_n3850, new_n3851, new_n3852,
    new_n3853, new_n3854, new_n3855, new_n3856, new_n3857, new_n3858,
    new_n3859, new_n3860, new_n3861, new_n3862, new_n3863, new_n3864,
    new_n3865, new_n3866, new_n3867, new_n3868, new_n3869, new_n3870,
    new_n3871, new_n3872, new_n3873, new_n3874, new_n3875, new_n3876,
    new_n3877, new_n3878, new_n3879, new_n3880, new_n3881, new_n3882,
    new_n3883, new_n3884, new_n3885, new_n3886, new_n3887, new_n3888,
    new_n3889, new_n3890, new_n3891, new_n3892, new_n3893, new_n3894,
    new_n3895, new_n3896, new_n3897, new_n3898, new_n3899, new_n3900,
    new_n3901, new_n3902, new_n3903, new_n3904, new_n3905, new_n3906,
    new_n3907, new_n3908, new_n3909, new_n3910, new_n3911, new_n3912,
    new_n3913, new_n3914, new_n3915, new_n3916, new_n3917, new_n3918,
    new_n3919, new_n3920, new_n3921, new_n3922, new_n3923, new_n3924,
    new_n3925, new_n3926, new_n3927, new_n3928, new_n3929, new_n3930,
    new_n3931, new_n3932, new_n3933, new_n3934, new_n3935, new_n3936,
    new_n3937, new_n3938, new_n3939, new_n3940, new_n3941, new_n3942,
    new_n3943, new_n3944, new_n3945, new_n3946, new_n3947, new_n3948,
    new_n3949, new_n3950, new_n3951, new_n3952, new_n3953, new_n3954,
    new_n3955, new_n3956, new_n3957, new_n3958, new_n3959, new_n3960,
    new_n3961, new_n3962, new_n3963, new_n3964, new_n3965, new_n3966,
    new_n3967, new_n3968, new_n3969, new_n3970, new_n3971, new_n3972,
    new_n3973, new_n3974, new_n3975, new_n3976, new_n3977, new_n3978,
    new_n3979, new_n3980, new_n3981, new_n3982, new_n3983, new_n3984,
    new_n3985, new_n3986, new_n3987, new_n3988, new_n3989, new_n3990,
    new_n3991, new_n3992, new_n3993, new_n3994, new_n3995, new_n3996,
    new_n3997, new_n3998, new_n3999, new_n4000, new_n4001, new_n4002,
    new_n4003, new_n4004, new_n4005, new_n4006, new_n4007, new_n4008,
    new_n4009, new_n4010, new_n4011, new_n4012, new_n4013, new_n4014,
    new_n4015, new_n4016, new_n4017, new_n4018, new_n4019, new_n4020,
    new_n4021, new_n4022, new_n4023, new_n4024, new_n4025, new_n4026,
    new_n4027, new_n4028, new_n4029, new_n4030, new_n4031, new_n4032,
    new_n4033, new_n4034, new_n4035, new_n4036, new_n4037, new_n4038,
    new_n4039, new_n4040, new_n4041, new_n4042, new_n4043, new_n4044,
    new_n4045, new_n4046, new_n4047, new_n4048, new_n4049, new_n4050,
    new_n4051, new_n4052, new_n4053, new_n4054, new_n4055, new_n4056,
    new_n4057, new_n4058, new_n4059, new_n4060, new_n4061, new_n4062,
    new_n4063, new_n4064, new_n4065, new_n4066, new_n4067, new_n4068,
    new_n4069, new_n4070, new_n4071, new_n4072, new_n4073, new_n4074,
    new_n4075, new_n4076, new_n4077, new_n4078, new_n4079, new_n4080,
    new_n4081, new_n4082, new_n4083, new_n4084, new_n4085, new_n4086,
    new_n4087, new_n4088, new_n4089, new_n4090, new_n4091, new_n4092,
    new_n4093, new_n4094, new_n4095, new_n4096, new_n4097, new_n4098,
    new_n4099, new_n4100, new_n4101, new_n4102, new_n4103, new_n4104,
    new_n4105, new_n4106, new_n4107, new_n4108, new_n4109, new_n4110,
    new_n4111, new_n4112, new_n4113, new_n4114, new_n4115, new_n4116,
    new_n4117, new_n4118, new_n4119, new_n4120, new_n4121, new_n4122,
    new_n4123, new_n4124, new_n4125, new_n4126, new_n4127, new_n4128,
    new_n4129, new_n4130, new_n4131, new_n4132, new_n4133, new_n4134,
    new_n4135, new_n4136, new_n4137, new_n4138, new_n4139, new_n4140,
    new_n4141, new_n4142, new_n4143, new_n4144, new_n4145, new_n4146,
    new_n4147, new_n4148, new_n4149, new_n4150, new_n4151, new_n4152,
    new_n4153, new_n4154, new_n4155, new_n4156, new_n4157, new_n4158,
    new_n4159, new_n4160, new_n4161, new_n4162, new_n4163, new_n4164,
    new_n4165, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170,
    new_n4171, new_n4172, new_n4173, new_n4174, new_n4175, new_n4176,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200,
    new_n4201, new_n4202, new_n4203, new_n4204, new_n4205, new_n4206,
    new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221, new_n4222, new_n4223, new_n4224,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230,
    new_n4231, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254,
    new_n4255, new_n4256, new_n4257, new_n4258, new_n4259, new_n4260,
    new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266,
    new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272,
    new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278,
    new_n4279, new_n4280, new_n4281, new_n4282, new_n4283, new_n4284,
    new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290,
    new_n4291, new_n4292, new_n4293, new_n4294, new_n4295, new_n4296,
    new_n4297, new_n4298, new_n4299, new_n4300, new_n4301, new_n4302,
    new_n4303, new_n4304, new_n4305, new_n4306, new_n4307, new_n4308,
    new_n4309, new_n4310, new_n4311, new_n4312, new_n4313, new_n4314,
    new_n4315, new_n4316, new_n4317, new_n4318, new_n4319, new_n4320,
    new_n4321, new_n4322, new_n4323, new_n4324, new_n4325, new_n4326,
    new_n4327, new_n4328, new_n4329, new_n4330, new_n4331, new_n4332,
    new_n4333, new_n4334, new_n4335, new_n4336, new_n4337, new_n4338,
    new_n4339, new_n4340, new_n4341, new_n4342, new_n4343, new_n4344,
    new_n4345, new_n4346, new_n4347, new_n4348, new_n4349, new_n4350,
    new_n4351, new_n4352, new_n4353, new_n4354, new_n4355, new_n4356,
    new_n4357, new_n4358, new_n4359, new_n4360, new_n4361, new_n4362,
    new_n4363, new_n4364, new_n4365, new_n4366, new_n4367, new_n4368,
    new_n4369, new_n4370, new_n4371, new_n4372, new_n4373, new_n4374,
    new_n4375, new_n4376, new_n4377, new_n4378, new_n4379, new_n4380,
    new_n4381, new_n4382, new_n4383, new_n4384, new_n4385, new_n4386,
    new_n4387, new_n4388, new_n4389, new_n4390, new_n4391, new_n4392,
    new_n4393, new_n4394, new_n4395, new_n4396, new_n4397, new_n4398,
    new_n4399, new_n4400, new_n4401, new_n4402, new_n4403, new_n4404,
    new_n4405, new_n4406, new_n4407, new_n4408, new_n4409, new_n4410,
    new_n4411, new_n4412, new_n4413, new_n4414, new_n4415, new_n4416,
    new_n4417, new_n4418, new_n4419, new_n4420, new_n4421, new_n4422,
    new_n4423, new_n4424, new_n4425, new_n4426, new_n4427, new_n4428,
    new_n4429, new_n4430, new_n4431, new_n4432, new_n4433, new_n4434,
    new_n4435, new_n4436, new_n4437, new_n4438, new_n4439, new_n4440,
    new_n4441, new_n4442, new_n4443, new_n4444, new_n4445, new_n4446,
    new_n4447, new_n4448, new_n4449, new_n4450, new_n4451, new_n4452,
    new_n4453, new_n4454, new_n4455, new_n4456, new_n4457, new_n4458,
    new_n4459, new_n4460, new_n4461, new_n4462, new_n4463, new_n4464,
    new_n4465, new_n4466, new_n4467, new_n4468, new_n4469, new_n4470,
    new_n4471, new_n4472, new_n4473, new_n4474, new_n4475, new_n4476,
    new_n4477, new_n4478, new_n4479, new_n4480, new_n4481, new_n4482,
    new_n4483, new_n4484, new_n4485, new_n4486, new_n4487, new_n4488,
    new_n4489, new_n4490, new_n4491, new_n4492, new_n4493, new_n4494,
    new_n4495, new_n4496, new_n4497, new_n4498, new_n4499, new_n4500,
    new_n4501, new_n4502, new_n4503, new_n4504, new_n4505, new_n4506,
    new_n4507, new_n4508, new_n4509, new_n4510, new_n4511, new_n4512,
    new_n4513, new_n4514, new_n4515, new_n4516, new_n4517, new_n4518,
    new_n4519, new_n4520, new_n4521, new_n4522, new_n4523, new_n4524,
    new_n4525, new_n4526, new_n4527, new_n4528, new_n4529, new_n4530,
    new_n4531, new_n4532, new_n4533, new_n4534, new_n4535, new_n4536,
    new_n4537, new_n4538, new_n4539, new_n4540, new_n4541, new_n4542,
    new_n4543, new_n4544, new_n4545, new_n4546, new_n4547, new_n4548,
    new_n4549, new_n4550, new_n4551, new_n4552, new_n4553, new_n4554,
    new_n4555, new_n4556, new_n4557, new_n4558, new_n4559, new_n4560,
    new_n4561, new_n4562, new_n4563, new_n4564, new_n4565, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4574, new_n4575, new_n4576, new_n4577, new_n4578,
    new_n4579, new_n4580, new_n4581, new_n4582, new_n4583, new_n4584,
    new_n4585, new_n4586, new_n4587, new_n4588, new_n4589, new_n4590,
    new_n4591, new_n4592, new_n4593, new_n4594, new_n4595, new_n4596,
    new_n4597, new_n4598, new_n4599, new_n4600, new_n4601, new_n4602,
    new_n4603, new_n4604, new_n4605, new_n4606, new_n4607, new_n4608,
    new_n4609, new_n4610, new_n4611, new_n4612, new_n4613, new_n4614,
    new_n4615, new_n4616, new_n4617, new_n4618, new_n4619, new_n4620,
    new_n4621, new_n4622, new_n4623, new_n4624, new_n4625, new_n4626,
    new_n4627, new_n4628, new_n4629, new_n4630, new_n4631, new_n4632,
    new_n4633, new_n4634, new_n4635, new_n4636, new_n4637, new_n4638,
    new_n4639, new_n4640, new_n4641, new_n4642, new_n4643, new_n4644,
    new_n4645, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650,
    new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656,
    new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662,
    new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668,
    new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674,
    new_n4675, new_n4676, new_n4677, new_n4678, new_n4679, new_n4680,
    new_n4681, new_n4682, new_n4683, new_n4684, new_n4685, new_n4686,
    new_n4687, new_n4688, new_n4689, new_n4690, new_n4691, new_n4692,
    new_n4693, new_n4694, new_n4695, new_n4696, new_n4697, new_n4698,
    new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704,
    new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710,
    new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716,
    new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722,
    new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728,
    new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743, new_n4744, new_n4745, new_n4746,
    new_n4747, new_n4748, new_n4749, new_n4750, new_n4751, new_n4752,
    new_n4753, new_n4754, new_n4755, new_n4756, new_n4757, new_n4758,
    new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764,
    new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770,
    new_n4771, new_n4772, new_n4773, new_n4774, new_n4775, new_n4776,
    new_n4777, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782,
    new_n4783, new_n4784, new_n4785, new_n4786, new_n4787, new_n4788,
    new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794,
    new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800,
    new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806,
    new_n4807, new_n4808, new_n4809, new_n4810, new_n4811, new_n4812,
    new_n4813, new_n4814, new_n4815, new_n4816, new_n4817, new_n4818,
    new_n4819, new_n4820, new_n4821, new_n4822, new_n4823, new_n4824,
    new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4830,
    new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836,
    new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842,
    new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848,
    new_n4849, new_n4850, new_n4851, new_n4852, new_n4853, new_n4854,
    new_n4855, new_n4856, new_n4857, new_n4858, new_n4859, new_n4860,
    new_n4861, new_n4862, new_n4863, new_n4864, new_n4865, new_n4866,
    new_n4867, new_n4868, new_n4869, new_n4870, new_n4871, new_n4872,
    new_n4873, new_n4874, new_n4875, new_n4876, new_n4877, new_n4878,
    new_n4879, new_n4880, new_n4881, new_n4882, new_n4883, new_n4884,
    new_n4885, new_n4886, new_n4887, new_n4888, new_n4889, new_n4890,
    new_n4891, new_n4892, new_n4893, new_n4894, new_n4895, new_n4896,
    new_n4897, new_n4898, new_n4899, new_n4900, new_n4901, new_n4902,
    new_n4903, new_n4904, new_n4905, new_n4906, new_n4907, new_n4908,
    new_n4909, new_n4910, new_n4911, new_n4912, new_n4913, new_n4914,
    new_n4915, new_n4916, new_n4917, new_n4918, new_n4919, new_n4920,
    new_n4921, new_n4922, new_n4923, new_n4924, new_n4925, new_n4926,
    new_n4927, new_n4928, new_n4929, new_n4930, new_n4931, new_n4932,
    new_n4933, new_n4934, new_n4935, new_n4936, new_n4937, new_n4938,
    new_n4939, new_n4940, new_n4941, new_n4942, new_n4943, new_n4944,
    new_n4945, new_n4946, new_n4947, new_n4948, new_n4949, new_n4950,
    new_n4951, new_n4952, new_n4953, new_n4954, new_n4955, new_n4956,
    new_n4957, new_n4958, new_n4959, new_n4960, new_n4961, new_n4962,
    new_n4963, new_n4964, new_n4965, new_n4966, new_n4967, new_n4968,
    new_n4969, new_n4970, new_n4971, new_n4972, new_n4973, new_n4974,
    new_n4975, new_n4976, new_n4977, new_n4978, new_n4979, new_n4980,
    new_n4981, new_n4982, new_n4983, new_n4984, new_n4985, new_n4986,
    new_n4987, new_n4988, new_n4989, new_n4990, new_n4991, new_n4992,
    new_n4993, new_n4994, new_n4995, new_n4996, new_n4997, new_n4998,
    new_n4999, new_n5000, new_n5001, new_n5002, new_n5003, new_n5004,
    new_n5005, new_n5006, new_n5007, new_n5008, new_n5009, new_n5010,
    new_n5011, new_n5012, new_n5013, new_n5014, new_n5015, new_n5016,
    new_n5017, new_n5018, new_n5019, new_n5020, new_n5021, new_n5022,
    new_n5023, new_n5024, new_n5025, new_n5026, new_n5027, new_n5028,
    new_n5029, new_n5030, new_n5031, new_n5032, new_n5033, new_n5034,
    new_n5035, new_n5036, new_n5037, new_n5038, new_n5039, new_n5040,
    new_n5041, new_n5042, new_n5043, new_n5044, new_n5045, new_n5046,
    new_n5047, new_n5048, new_n5049, new_n5050, new_n5051, new_n5052,
    new_n5053, new_n5054, new_n5055, new_n5056, new_n5057, new_n5058,
    new_n5059, new_n5060, new_n5061, new_n5062, new_n5063, new_n5064,
    new_n5065, new_n5066, new_n5067, new_n5068, new_n5069, new_n5070,
    new_n5071, new_n5072, new_n5073, new_n5074, new_n5075, new_n5076,
    new_n5077, new_n5078, new_n5079, new_n5080, new_n5081, new_n5082,
    new_n5083, new_n5084, new_n5085, new_n5086, new_n5087, new_n5088,
    new_n5089, new_n5090, new_n5091, new_n5092, new_n5093, new_n5094,
    new_n5095, new_n5096, new_n5097, new_n5098, new_n5099, new_n5100,
    new_n5101, new_n5102, new_n5103, new_n5104, new_n5105, new_n5106,
    new_n5107, new_n5108, new_n5109, new_n5110, new_n5111, new_n5112,
    new_n5113, new_n5114, new_n5115, new_n5116, new_n5117, new_n5118,
    new_n5119, new_n5120, new_n5121, new_n5122, new_n5123, new_n5124,
    new_n5125, new_n5126, new_n5127, new_n5128, new_n5129, new_n5130,
    new_n5131, new_n5132, new_n5133, new_n5134, new_n5135, new_n5136,
    new_n5137, new_n5138, new_n5139, new_n5140, new_n5141, new_n5142,
    new_n5143, new_n5144, new_n5145, new_n5146, new_n5147, new_n5148,
    new_n5149, new_n5150, new_n5151, new_n5152, new_n5153, new_n5154,
    new_n5155, new_n5156, new_n5157, new_n5158, new_n5159, new_n5160,
    new_n5161, new_n5162, new_n5163, new_n5164, new_n5165, new_n5166,
    new_n5167, new_n5168, new_n5169, new_n5170, new_n5171, new_n5172,
    new_n5173, new_n5174, new_n5175, new_n5176, new_n5177, new_n5178,
    new_n5179, new_n5180, new_n5181, new_n5182, new_n5183, new_n5184,
    new_n5185, new_n5186, new_n5187, new_n5188, new_n5189, new_n5190,
    new_n5191, new_n5192, new_n5193, new_n5194, new_n5195, new_n5196,
    new_n5197, new_n5198, new_n5199, new_n5200, new_n5201, new_n5202,
    new_n5203, new_n5204, new_n5205, new_n5206, new_n5207, new_n5208,
    new_n5209, new_n5210, new_n5211, new_n5212, new_n5213, new_n5214,
    new_n5215, new_n5216, new_n5217, new_n5218, new_n5219, new_n5220,
    new_n5221, new_n5222, new_n5223, new_n5224, new_n5225, new_n5226,
    new_n5227, new_n5228, new_n5229, new_n5230, new_n5231, new_n5232,
    new_n5233, new_n5234, new_n5235, new_n5236, new_n5237, new_n5238,
    new_n5239, new_n5240, new_n5241, new_n5242, new_n5243, new_n5244,
    new_n5245, new_n5246, new_n5247, new_n5248, new_n5249, new_n5250,
    new_n5251, new_n5252, new_n5253, new_n5254, new_n5255, new_n5256,
    new_n5257, new_n5258, new_n5259, new_n5260, new_n5261, new_n5262,
    new_n5263, new_n5264, new_n5265, new_n5266, new_n5267, new_n5268,
    new_n5269, new_n5270, new_n5271, new_n5272, new_n5273, new_n5274,
    new_n5275, new_n5276, new_n5277, new_n5278, new_n5279, new_n5280,
    new_n5281, new_n5282, new_n5283, new_n5284, new_n5285, new_n5286,
    new_n5287, new_n5288, new_n5289, new_n5290, new_n5291, new_n5292,
    new_n5293, new_n5294, new_n5295, new_n5296, new_n5297, new_n5298,
    new_n5299, new_n5300, new_n5301, new_n5302, new_n5303, new_n5304,
    new_n5305, new_n5306, new_n5307, new_n5308, new_n5309, new_n5310,
    new_n5311, new_n5312, new_n5313, new_n5314, new_n5315, new_n5316,
    new_n5317, new_n5318, new_n5319, new_n5320, new_n5321, new_n5322,
    new_n5323, new_n5324, new_n5325, new_n5326, new_n5327, new_n5328,
    new_n5329, new_n5330, new_n5331, new_n5332, new_n5333, new_n5334,
    new_n5335, new_n5336, new_n5337, new_n5338, new_n5339, new_n5340,
    new_n5341, new_n5342, new_n5343, new_n5344, new_n5345, new_n5346,
    new_n5347, new_n5348, new_n5349, new_n5350, new_n5351, new_n5352,
    new_n5353, new_n5354, new_n5355, new_n5356, new_n5357, new_n5358,
    new_n5359, new_n5360, new_n5361, new_n5362, new_n5363, new_n5364,
    new_n5365, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370,
    new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376,
    new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382,
    new_n5383, new_n5384, new_n5385, new_n5386, new_n5387, new_n5388,
    new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394,
    new_n5395, new_n5396, new_n5397, new_n5398, new_n5399, new_n5400,
    new_n5401, new_n5402, new_n5403, new_n5404, new_n5405, new_n5406,
    new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412,
    new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418,
    new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424,
    new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430,
    new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436,
    new_n5437, new_n5438, new_n5439, new_n5440, new_n5441, new_n5442,
    new_n5443, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448,
    new_n5449, new_n5450, new_n5451, new_n5452, new_n5453, new_n5454,
    new_n5455, new_n5456, new_n5457, new_n5458, new_n5459, new_n5460,
    new_n5461, new_n5462, new_n5463, new_n5464, new_n5465, new_n5466,
    new_n5467, new_n5468, new_n5469, new_n5470, new_n5471, new_n5472,
    new_n5473, new_n5474, new_n5475, new_n5476, new_n5477, new_n5478,
    new_n5479, new_n5480, new_n5481, new_n5482, new_n5483, new_n5484,
    new_n5485, new_n5486, new_n5487, new_n5488, new_n5489, new_n5490,
    new_n5491, new_n5492, new_n5493, new_n5494, new_n5495, new_n5496,
    new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502,
    new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508,
    new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514,
    new_n5515, new_n5516, new_n5517, new_n5518, new_n5519, new_n5520,
    new_n5521, new_n5522, new_n5523, new_n5524, new_n5525, new_n5526,
    new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532,
    new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538,
    new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544,
    new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550,
    new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556,
    new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562,
    new_n5563, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586,
    new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592,
    new_n5593, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598,
    new_n5599, new_n5600, new_n5601, new_n5602, new_n5603, new_n5604,
    new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610,
    new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5616,
    new_n5617, new_n5618, new_n5619, new_n5620, new_n5621, new_n5622,
    new_n5623, new_n5624, new_n5625, new_n5626, new_n5627, new_n5628,
    new_n5629, new_n5630, new_n5631, new_n5632, new_n5633, new_n5634,
    new_n5635, new_n5636, new_n5637, new_n5638, new_n5639, new_n5640,
    new_n5641, new_n5642, new_n5643, new_n5644, new_n5645, new_n5646,
    new_n5647, new_n5648, new_n5649, new_n5650, new_n5651, new_n5652,
    new_n5653, new_n5654, new_n5655, new_n5656, new_n5657, new_n5658,
    new_n5659, new_n5660, new_n5661, new_n5662, new_n5663, new_n5664,
    new_n5665, new_n5666, new_n5667, new_n5668, new_n5669, new_n5670,
    new_n5671, new_n5672, new_n5673, new_n5674, new_n5675, new_n5676,
    new_n5677, new_n5678, new_n5679, new_n5680, new_n5681, new_n5682,
    new_n5683, new_n5684, new_n5685, new_n5686, new_n5687, new_n5688,
    new_n5689, new_n5690, new_n5691, new_n5692, new_n5693, new_n5694,
    new_n5695, new_n5696, new_n5697, new_n5698, new_n5699, new_n5700,
    new_n5701, new_n5702, new_n5703, new_n5704, new_n5705, new_n5706,
    new_n5707, new_n5708, new_n5709, new_n5710, new_n5711, new_n5712,
    new_n5713, new_n5714, new_n5715, new_n5716, new_n5717, new_n5718,
    new_n5719, new_n5720, new_n5721, new_n5722, new_n5723, new_n5724,
    new_n5725, new_n5726, new_n5727, new_n5728, new_n5729, new_n5730,
    new_n5731, new_n5732, new_n5733, new_n5734, new_n5735, new_n5736,
    new_n5737, new_n5738, new_n5739, new_n5740, new_n5741, new_n5742,
    new_n5743, new_n5744, new_n5745, new_n5746, new_n5747, new_n5748,
    new_n5749, new_n5750, new_n5751, new_n5752, new_n5753, new_n5754,
    new_n5755, new_n5756, new_n5757, new_n5758, new_n5759, new_n5760,
    new_n5761, new_n5762, new_n5763, new_n5764, new_n5765, new_n5766,
    new_n5767, new_n5768, new_n5769, new_n5770, new_n5771, new_n5772,
    new_n5773, new_n5774, new_n5775, new_n5776, new_n5777, new_n5778,
    new_n5779, new_n5780, new_n5781, new_n5782, new_n5783, new_n5784,
    new_n5785, new_n5786, new_n5787, new_n5788, new_n5789, new_n5790,
    new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796,
    new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5806, new_n5807, new_n5808,
    new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850,
    new_n5851, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856,
    new_n5857, new_n5858, new_n5859, new_n5860, new_n5861, new_n5862,
    new_n5863, new_n5864, new_n5865, new_n5866, new_n5867, new_n5868,
    new_n5869, new_n5870, new_n5871, new_n5872, new_n5873, new_n5874,
    new_n5875, new_n5876, new_n5877, new_n5878, new_n5879, new_n5880,
    new_n5881, new_n5882, new_n5883, new_n5884, new_n5885, new_n5886,
    new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892,
    new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898,
    new_n5899, new_n5900, new_n5901, new_n5902, new_n5903, new_n5904,
    new_n5905, new_n5906, new_n5907, new_n5908, new_n5909, new_n5910,
    new_n5911, new_n5912, new_n5913, new_n5914, new_n5915, new_n5916,
    new_n5917, new_n5918, new_n5919, new_n5920, new_n5921, new_n5922,
    new_n5923, new_n5924, new_n5925, new_n5926, new_n5927, new_n5928,
    new_n5929, new_n5930, new_n5931, new_n5932, new_n5933, new_n5934,
    new_n5935, new_n5936, new_n5937, new_n5938, new_n5939, new_n5940,
    new_n5941, new_n5942, new_n5943, new_n5944, new_n5945, new_n5946,
    new_n5947, new_n5948, new_n5949, new_n5950, new_n5951, new_n5952,
    new_n5953, new_n5954, new_n5955, new_n5956, new_n5957, new_n5958,
    new_n5959, new_n5960, new_n5961, new_n5962, new_n5963, new_n5964,
    new_n5965, new_n5966, new_n5967, new_n5968, new_n5969, new_n5970,
    new_n5971, new_n5972, new_n5973, new_n5974, new_n5975, new_n5976,
    new_n5977, new_n5978, new_n5979, new_n5980, new_n5981, new_n5982,
    new_n5983, new_n5984, new_n5985, new_n5986, new_n5987, new_n5988,
    new_n5989, new_n5990, new_n5991, new_n5992, new_n5993, new_n5994,
    new_n5995, new_n5996, new_n5997, new_n5998, new_n5999, new_n6000,
    new_n6001, new_n6002, new_n6003, new_n6004, new_n6005, new_n6006,
    new_n6007, new_n6008, new_n6009, new_n6010, new_n6011, new_n6012,
    new_n6013, new_n6014, new_n6015, new_n6016, new_n6017, new_n6018,
    new_n6019, new_n6020, new_n6021, new_n6022, new_n6023, new_n6024,
    new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030,
    new_n6031, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036,
    new_n6037, new_n6038, new_n6039, new_n6040, new_n6041, new_n6042,
    new_n6043, new_n6044, new_n6045, new_n6046, new_n6047, new_n6048,
    new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6054,
    new_n6055, new_n6056, new_n6057, new_n6058, new_n6059, new_n6060,
    new_n6061, new_n6062, new_n6063, new_n6064, new_n6065, new_n6066,
    new_n6067, new_n6068, new_n6069, new_n6070, new_n6071, new_n6072,
    new_n6073, new_n6074, new_n6075, new_n6076, new_n6077, new_n6078,
    new_n6079, new_n6080, new_n6081, new_n6082, new_n6083, new_n6084,
    new_n6085, new_n6086, new_n6087, new_n6088, new_n6089, new_n6090,
    new_n6091, new_n6092, new_n6093, new_n6094, new_n6095, new_n6096,
    new_n6097, new_n6098, new_n6099, new_n6100, new_n6101, new_n6102,
    new_n6103, new_n6104, new_n6105, new_n6106, new_n6107, new_n6108,
    new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114,
    new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120,
    new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126,
    new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384,
    new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407, new_n6408,
    new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427, new_n6428, new_n6429, new_n6430, new_n6431, new_n6432,
    new_n6433, new_n6434, new_n6435, new_n6436, new_n6437, new_n6438,
    new_n6439, new_n6440, new_n6441, new_n6442, new_n6443, new_n6444,
    new_n6445, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456,
    new_n6457, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476, new_n6477, new_n6478, new_n6479, new_n6480,
    new_n6481, new_n6482, new_n6483, new_n6484, new_n6485, new_n6486,
    new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492,
    new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6498,
    new_n6499, new_n6500, new_n6501, new_n6502, new_n6503, new_n6504,
    new_n6505, new_n6506, new_n6507, new_n6508, new_n6509, new_n6510,
    new_n6511, new_n6512, new_n6513, new_n6514, new_n6515, new_n6516,
    new_n6517, new_n6518, new_n6519, new_n6520, new_n6521, new_n6522,
    new_n6523, new_n6524, new_n6525, new_n6526, new_n6527, new_n6528,
    new_n6529, new_n6530, new_n6531, new_n6532, new_n6533, new_n6534,
    new_n6535, new_n6536, new_n6537, new_n6538, new_n6539, new_n6540,
    new_n6541, new_n6542, new_n6543, new_n6544, new_n6545, new_n6546,
    new_n6547, new_n6548, new_n6549, new_n6550, new_n6551, new_n6552,
    new_n6553, new_n6554, new_n6555, new_n6556, new_n6557, new_n6558,
    new_n6559, new_n6560, new_n6561, new_n6562, new_n6563, new_n6564,
    new_n6565, new_n6566, new_n6567, new_n6568, new_n6569, new_n6570,
    new_n6571, new_n6572, new_n6573, new_n6574, new_n6575, new_n6576,
    new_n6577, new_n6578, new_n6579, new_n6580, new_n6581, new_n6582,
    new_n6583, new_n6584, new_n6585, new_n6586, new_n6587, new_n6588,
    new_n6589, new_n6590, new_n6591, new_n6592, new_n6593, new_n6594,
    new_n6595, new_n6596, new_n6597, new_n6598, new_n6599, new_n6600,
    new_n6601, new_n6602, new_n6603, new_n6604, new_n6605, new_n6606,
    new_n6607, new_n6608, new_n6609, new_n6610, new_n6611, new_n6612,
    new_n6613, new_n6614, new_n6615, new_n6616, new_n6617, new_n6618,
    new_n6619, new_n6620, new_n6621, new_n6622, new_n6623, new_n6624,
    new_n6625, new_n6626, new_n6627, new_n6628, new_n6629, new_n6630,
    new_n6631, new_n6632, new_n6633, new_n6634, new_n6635, new_n6636,
    new_n6637, new_n6638, new_n6639, new_n6640, new_n6641, new_n6642,
    new_n6643, new_n6644, new_n6645, new_n6646, new_n6647, new_n6648,
    new_n6649, new_n6650, new_n6651, new_n6652, new_n6653, new_n6654,
    new_n6655, new_n6656, new_n6657, new_n6658, new_n6659, new_n6660,
    new_n6661, new_n6662, new_n6663, new_n6664, new_n6665, new_n6666,
    new_n6667, new_n6668, new_n6669, new_n6670, new_n6671, new_n6672,
    new_n6673, new_n6674, new_n6675, new_n6676, new_n6677, new_n6678,
    new_n6679, new_n6680, new_n6681, new_n6682, new_n6683, new_n6684,
    new_n6685, new_n6686, new_n6687, new_n6688, new_n6689, new_n6690,
    new_n6691, new_n6692, new_n6693, new_n6694, new_n6695, new_n6696,
    new_n6697, new_n6698, new_n6699, new_n6700, new_n6701, new_n6702,
    new_n6703, new_n6704, new_n6705, new_n6706, new_n6707, new_n6708,
    new_n6709, new_n6710, new_n6711, new_n6712, new_n6713, new_n6714,
    new_n6715, new_n6716, new_n6717, new_n6718, new_n6719, new_n6720,
    new_n6721, new_n6722, new_n6723, new_n6724, new_n6725, new_n6726,
    new_n6727, new_n6728, new_n6729, new_n6730, new_n6731, new_n6732,
    new_n6733, new_n6734, new_n6735, new_n6736, new_n6737, new_n6738,
    new_n6739, new_n6740, new_n6741, new_n6742, new_n6743, new_n6744,
    new_n6745, new_n6746, new_n6747, new_n6748, new_n6749, new_n6750,
    new_n6751, new_n6752, new_n6753, new_n6754, new_n6755, new_n6756,
    new_n6757, new_n6758, new_n6759, new_n6760, new_n6761, new_n6762,
    new_n6763, new_n6764, new_n6765, new_n6766, new_n6767, new_n6768,
    new_n6769, new_n6770, new_n6771, new_n6772, new_n6773, new_n6774,
    new_n6775, new_n6776, new_n6777, new_n6778, new_n6779, new_n6780,
    new_n6781, new_n6782, new_n6783, new_n6784, new_n6785, new_n6786,
    new_n6787, new_n6788, new_n6789, new_n6790, new_n6791, new_n6792,
    new_n6793, new_n6794, new_n6795, new_n6796, new_n6797, new_n6798,
    new_n6799, new_n6800, new_n6801, new_n6802, new_n6803, new_n6804,
    new_n6805, new_n6806, new_n6807, new_n6808, new_n6809, new_n6810,
    new_n6811, new_n6812, new_n6813, new_n6814, new_n6815, new_n6816,
    new_n6817, new_n6818, new_n6819, new_n6820, new_n6821, new_n6822,
    new_n6823, new_n6824, new_n6825, new_n6826, new_n6827, new_n6828,
    new_n6829, new_n6830, new_n6831, new_n6832, new_n6833, new_n6834,
    new_n6835, new_n6836, new_n6837, new_n6838, new_n6839, new_n6840,
    new_n6841, new_n6842, new_n6843, new_n6844, new_n6845, new_n6846,
    new_n6847, new_n6848, new_n6849, new_n6850, new_n6851, new_n6852,
    new_n6853, new_n6854, new_n6855, new_n6856, new_n6857, new_n6858,
    new_n6859, new_n6860, new_n6861, new_n6862, new_n6863, new_n6864,
    new_n6865, new_n6866, new_n6867, new_n6868, new_n6869, new_n6870,
    new_n6871, new_n6872, new_n6873, new_n6874, new_n6875, new_n6876,
    new_n6877, new_n6878, new_n6879, new_n6880, new_n6881, new_n6882,
    new_n6883, new_n6884, new_n6885, new_n6886, new_n6887, new_n6888,
    new_n6889, new_n6890, new_n6891, new_n6892, new_n6893, new_n6894,
    new_n6895, new_n6896, new_n6897, new_n6898, new_n6899, new_n6900,
    new_n6901, new_n6902, new_n6903, new_n6904, new_n6905, new_n6906,
    new_n6907, new_n6908, new_n6909, new_n6910, new_n6911, new_n6912,
    new_n6913, new_n6914, new_n6915, new_n6916, new_n6917, new_n6918,
    new_n6919, new_n6920, new_n6921, new_n6922, new_n6923, new_n6924,
    new_n6925, new_n6926, new_n6927, new_n6928, new_n6929, new_n6930,
    new_n6931, new_n6932, new_n6933, new_n6934, new_n6935, new_n6936,
    new_n6937, new_n6938, new_n6939, new_n6940, new_n6941, new_n6942,
    new_n6943, new_n6944, new_n6945, new_n6946, new_n6947, new_n6948,
    new_n6949, new_n6950, new_n6951, new_n6952, new_n6953, new_n6954,
    new_n6955, new_n6956, new_n6957, new_n6958, new_n6959, new_n6960,
    new_n6961, new_n6962, new_n6963, new_n6964, new_n6965, new_n6966,
    new_n6967, new_n6968, new_n6969, new_n6970, new_n6971, new_n6972,
    new_n6973, new_n6974, new_n6975, new_n6976, new_n6977, new_n6978,
    new_n6979, new_n6980, new_n6981, new_n6982, new_n6983, new_n6984,
    new_n6985, new_n6986, new_n6987, new_n6988, new_n6989, new_n6990,
    new_n6991, new_n6992, new_n6993, new_n6994, new_n6995, new_n6996,
    new_n6997, new_n6998, new_n6999, new_n7000, new_n7001, new_n7002,
    new_n7003, new_n7004, new_n7005, new_n7006, new_n7007, new_n7008,
    new_n7009, new_n7010, new_n7011, new_n7012, new_n7013, new_n7014,
    new_n7015, new_n7016, new_n7017, new_n7018, new_n7019, new_n7020,
    new_n7021, new_n7022, new_n7023, new_n7024, new_n7025, new_n7026,
    new_n7027, new_n7028, new_n7029, new_n7030, new_n7031, new_n7032,
    new_n7033, new_n7034, new_n7035, new_n7036, new_n7037, new_n7038,
    new_n7039, new_n7040, new_n7041, new_n7042, new_n7043, new_n7044,
    new_n7045, new_n7046, new_n7047, new_n7048, new_n7049, new_n7050,
    new_n7051, new_n7052, new_n7053, new_n7054, new_n7055, new_n7056,
    new_n7057, new_n7058, new_n7059, new_n7060, new_n7061, new_n7062,
    new_n7063, new_n7064, new_n7065, new_n7066, new_n7067, new_n7068,
    new_n7069, new_n7070, new_n7071, new_n7072, new_n7073, new_n7074,
    new_n7075, new_n7076, new_n7077, new_n7078, new_n7079, new_n7080,
    new_n7081, new_n7082, new_n7083, new_n7084, new_n7085, new_n7086,
    new_n7087, new_n7088, new_n7089, new_n7090, new_n7091, new_n7092,
    new_n7093, new_n7094, new_n7095, new_n7096, new_n7097, new_n7098,
    new_n7099, new_n7100, new_n7101, new_n7102, new_n7103, new_n7104,
    new_n7105, new_n7106, new_n7107, new_n7108, new_n7109, new_n7110,
    new_n7111, new_n7112, new_n7113, new_n7114, new_n7115, new_n7116,
    new_n7117, new_n7118, new_n7119, new_n7120, new_n7121, new_n7122,
    new_n7123, new_n7124, new_n7125, new_n7126, new_n7127, new_n7128,
    new_n7129, new_n7130, new_n7131, new_n7132, new_n7133, new_n7134,
    new_n7135, new_n7136, new_n7137, new_n7138, new_n7139, new_n7140,
    new_n7141, new_n7142, new_n7143, new_n7144, new_n7145, new_n7146,
    new_n7147, new_n7148, new_n7149, new_n7150, new_n7151, new_n7152,
    new_n7153, new_n7154, new_n7155, new_n7156, new_n7157, new_n7158,
    new_n7159, new_n7160, new_n7161, new_n7162, new_n7163, new_n7164,
    new_n7165, new_n7166, new_n7167, new_n7168, new_n7169, new_n7170,
    new_n7171, new_n7172, new_n7173, new_n7174, new_n7175, new_n7176,
    new_n7177, new_n7178, new_n7179, new_n7180, new_n7181, new_n7182,
    new_n7183, new_n7184, new_n7185, new_n7186, new_n7187, new_n7188,
    new_n7189, new_n7190, new_n7191, new_n7192, new_n7193, new_n7194,
    new_n7195, new_n7196, new_n7197, new_n7198, new_n7199, new_n7200,
    new_n7201, new_n7202, new_n7203, new_n7204, new_n7205, new_n7206,
    new_n7207, new_n7208, new_n7209, new_n7210, new_n7211, new_n7212,
    new_n7213, new_n7214, new_n7215, new_n7216, new_n7217, new_n7218,
    new_n7219, new_n7220, new_n7221, new_n7222, new_n7223, new_n7224,
    new_n7225, new_n7226, new_n7227, new_n7228, new_n7229, new_n7230,
    new_n7231, new_n7232, new_n7233, new_n7234, new_n7235, new_n7236,
    new_n7237, new_n7238, new_n7239, new_n7240, new_n7241, new_n7242,
    new_n7243, new_n7244, new_n7245, new_n7246, new_n7247, new_n7248,
    new_n7249, new_n7250, new_n7251, new_n7252, new_n7253, new_n7254,
    new_n7255, new_n7256, new_n7257, new_n7258, new_n7259, new_n7260,
    new_n7261, new_n7262, new_n7263, new_n7264, new_n7265, new_n7266,
    new_n7267, new_n7268, new_n7269, new_n7270, new_n7271, new_n7272,
    new_n7273, new_n7274, new_n7275, new_n7276, new_n7277, new_n7278,
    new_n7279, new_n7280, new_n7281, new_n7282, new_n7283, new_n7284,
    new_n7285, new_n7286, new_n7287, new_n7288, new_n7289, new_n7290,
    new_n7291, new_n7292, new_n7293, new_n7294, new_n7295, new_n7296,
    new_n7297, new_n7298, new_n7299, new_n7300, new_n7301, new_n7302,
    new_n7303, new_n7304, new_n7305, new_n7306, new_n7307, new_n7308,
    new_n7309, new_n7310, new_n7311, new_n7312, new_n7313, new_n7314,
    new_n7315, new_n7316, new_n7317, new_n7318, new_n7319, new_n7320,
    new_n7321, new_n7322, new_n7323, new_n7324, new_n7325, new_n7326,
    new_n7327, new_n7328, new_n7329, new_n7330, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335, new_n7336, new_n7337, new_n7338,
    new_n7339, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346, new_n7347, new_n7348, new_n7349, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428,
    new_n7429, new_n7430, new_n7431, new_n7432, new_n7433, new_n7434,
    new_n7435, new_n7436, new_n7437, new_n7438, new_n7439, new_n7440,
    new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446,
    new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452,
    new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458,
    new_n7459, new_n7460, new_n7461, new_n7462, new_n7463, new_n7464,
    new_n7465, new_n7466, new_n7467, new_n7468, new_n7469, new_n7470,
    new_n7471, new_n7472, new_n7473, new_n7474, new_n7475, new_n7476,
    new_n7477, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482,
    new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488,
    new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494,
    new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500,
    new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506,
    new_n7507, new_n7508, new_n7509, new_n7510, new_n7511, new_n7512,
    new_n7513, new_n7514, new_n7515, new_n7516, new_n7517, new_n7518,
    new_n7519, new_n7520, new_n7521, new_n7522, new_n7523, new_n7524,
    new_n7525, new_n7526, new_n7527, new_n7528, new_n7529, new_n7530,
    new_n7531, new_n7532, new_n7533, new_n7534, new_n7535, new_n7536,
    new_n7537, new_n7538, new_n7539, new_n7540, new_n7541, new_n7542,
    new_n7543, new_n7544, new_n7545, new_n7546, new_n7547, new_n7548,
    new_n7549, new_n7550, new_n7551, new_n7552, new_n7553, new_n7554,
    new_n7555, new_n7556, new_n7557, new_n7558, new_n7559, new_n7560,
    new_n7561, new_n7562, new_n7563, new_n7564, new_n7565, new_n7566,
    new_n7567, new_n7568, new_n7569, new_n7570, new_n7571, new_n7572,
    new_n7573, new_n7574, new_n7575, new_n7576, new_n7577, new_n7578,
    new_n7579, new_n7580, new_n7581, new_n7582, new_n7583, new_n7584,
    new_n7585, new_n7586, new_n7587, new_n7588, new_n7589, new_n7590,
    new_n7591, new_n7592, new_n7593, new_n7594, new_n7595, new_n7596,
    new_n7597, new_n7598, new_n7599, new_n7600, new_n7601, new_n7602,
    new_n7603, new_n7604, new_n7605, new_n7606, new_n7607, new_n7608,
    new_n7609, new_n7610, new_n7611, new_n7612, new_n7613, new_n7614,
    new_n7615, new_n7616, new_n7617, new_n7618, new_n7619, new_n7620,
    new_n7621, new_n7622, new_n7623, new_n7624, new_n7625, new_n7626,
    new_n7627, new_n7628, new_n7629, new_n7630, new_n7631, new_n7632,
    new_n7633, new_n7634, new_n7635, new_n7636, new_n7637, new_n7638,
    new_n7639, new_n7640, new_n7641, new_n7642, new_n7643, new_n7644,
    new_n7645, new_n7646, new_n7647, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674,
    new_n7675, new_n7676, new_n7677, new_n7678, new_n7679, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692,
    new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730, new_n7731, new_n7732, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770,
    new_n7771, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806,
    new_n7807, new_n7808, new_n7809, new_n7810, new_n7811, new_n7812,
    new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818,
    new_n7819, new_n7820, new_n7821, new_n7822, new_n7823, new_n7824,
    new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830,
    new_n7831, new_n7832, new_n7833, new_n7834, new_n7835, new_n7836,
    new_n7837, new_n7838, new_n7839, new_n7840, new_n7841, new_n7842,
    new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848,
    new_n7849, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884,
    new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890,
    new_n7891, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896,
    new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902,
    new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7909, new_n7910, new_n7911, new_n7912, new_n7913, new_n7914,
    new_n7915, new_n7916, new_n7917, new_n7918, new_n7919, new_n7920,
    new_n7921, new_n7922, new_n7923, new_n7924, new_n7925, new_n7926,
    new_n7927, new_n7928, new_n7929, new_n7930, new_n7931, new_n7932,
    new_n7933, new_n7934, new_n7935, new_n7936, new_n7937, new_n7938,
    new_n7939, new_n7940, new_n7941, new_n7942, new_n7943, new_n7944,
    new_n7945, new_n7946, new_n7947, new_n7948, new_n7949, new_n7950,
    new_n7951, new_n7952, new_n7953, new_n7954, new_n7955, new_n7956,
    new_n7957, new_n7958, new_n7959, new_n7960, new_n7961, new_n7962,
    new_n7963, new_n7964, new_n7965, new_n7966, new_n7967, new_n7968,
    new_n7969, new_n7970, new_n7971, new_n7972, new_n7973, new_n7974,
    new_n7975, new_n7976, new_n7977, new_n7978, new_n7979, new_n7980,
    new_n7981, new_n7982, new_n7983, new_n7984, new_n7985, new_n7986,
    new_n7987, new_n7988, new_n7989, new_n7990, new_n7991, new_n7992,
    new_n7993, new_n7994, new_n7995, new_n7996, new_n7997, new_n7998,
    new_n7999, new_n8000, new_n8001, new_n8002, new_n8003, new_n8004,
    new_n8005, new_n8006, new_n8007, new_n8008, new_n8009, new_n8010,
    new_n8011, new_n8012, new_n8013, new_n8014, new_n8015, new_n8016,
    new_n8017, new_n8018, new_n8019, new_n8020, new_n8021, new_n8022,
    new_n8023, new_n8024, new_n8025, new_n8026, new_n8027, new_n8028,
    new_n8029, new_n8030, new_n8031, new_n8032, new_n8033, new_n8034,
    new_n8035, new_n8036, new_n8037, new_n8038, new_n8039, new_n8040,
    new_n8041, new_n8042, new_n8043, new_n8044, new_n8045, new_n8046,
    new_n8047, new_n8048, new_n8049, new_n8050, new_n8051, new_n8052,
    new_n8053, new_n8054, new_n8055, new_n8056, new_n8057, new_n8058,
    new_n8059, new_n8060, new_n8061, new_n8062, new_n8063, new_n8064,
    new_n8065, new_n8066, new_n8067, new_n8068, new_n8069, new_n8070,
    new_n8071, new_n8072, new_n8073, new_n8074, new_n8075, new_n8076,
    new_n8077, new_n8078, new_n8079, new_n8080, new_n8081, new_n8082,
    new_n8083, new_n8084, new_n8085, new_n8086, new_n8087, new_n8088,
    new_n8089, new_n8090, new_n8091, new_n8092, new_n8093, new_n8094,
    new_n8095, new_n8096, new_n8097, new_n8098, new_n8099, new_n8100,
    new_n8101, new_n8102, new_n8103, new_n8104, new_n8105, new_n8106,
    new_n8107, new_n8108, new_n8109, new_n8110, new_n8111, new_n8112,
    new_n8113, new_n8114, new_n8115, new_n8116, new_n8117, new_n8118,
    new_n8119, new_n8120, new_n8121, new_n8122, new_n8123, new_n8124,
    new_n8125, new_n8126, new_n8127, new_n8128, new_n8129, new_n8130,
    new_n8131, new_n8132, new_n8133, new_n8134, new_n8135, new_n8136,
    new_n8137, new_n8138, new_n8139, new_n8140, new_n8141, new_n8142,
    new_n8143, new_n8144, new_n8145, new_n8146, new_n8147, new_n8148,
    new_n8149, new_n8150, new_n8151, new_n8152, new_n8153, new_n8154,
    new_n8155, new_n8156, new_n8157, new_n8158, new_n8159, new_n8160,
    new_n8161, new_n8162, new_n8163, new_n8164, new_n8165, new_n8166,
    new_n8167, new_n8168, new_n8169, new_n8170, new_n8171, new_n8172,
    new_n8173, new_n8174, new_n8175, new_n8176, new_n8177, new_n8178,
    new_n8179, new_n8180, new_n8181, new_n8182, new_n8183, new_n8184,
    new_n8185, new_n8186, new_n8187, new_n8188, new_n8189, new_n8190,
    new_n8191, new_n8192, new_n8193, new_n8194, new_n8195, new_n8196,
    new_n8197, new_n8198, new_n8199, new_n8200, new_n8201, new_n8202,
    new_n8203, new_n8204, new_n8205, new_n8206, new_n8207, new_n8208,
    new_n8209, new_n8210, new_n8211, new_n8212, new_n8213, new_n8214,
    new_n8215, new_n8216, new_n8217, new_n8218, new_n8219, new_n8220,
    new_n8221, new_n8222, new_n8223, new_n8224, new_n8225, new_n8226,
    new_n8227, new_n8228, new_n8229, new_n8230, new_n8231, new_n8232,
    new_n8233, new_n8234, new_n8235, new_n8236, new_n8237, new_n8238,
    new_n8239, new_n8240, new_n8241, new_n8242, new_n8243, new_n8244,
    new_n8245, new_n8246, new_n8247, new_n8248, new_n8249, new_n8250,
    new_n8251, new_n8252, new_n8253, new_n8254, new_n8255, new_n8256,
    new_n8257, new_n8258, new_n8259, new_n8260, new_n8261, new_n8262,
    new_n8263, new_n8264, new_n8265, new_n8266, new_n8267, new_n8268,
    new_n8269, new_n8270, new_n8271, new_n8272, new_n8273, new_n8274,
    new_n8275, new_n8276, new_n8277, new_n8278, new_n8279, new_n8280,
    new_n8281, new_n8282, new_n8283, new_n8284, new_n8285, new_n8286,
    new_n8287, new_n8288, new_n8289, new_n8290, new_n8291, new_n8292,
    new_n8293, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298,
    new_n8299, new_n8300, new_n8301, new_n8302, new_n8303, new_n8304,
    new_n8305, new_n8306, new_n8307, new_n8308, new_n8309, new_n8310,
    new_n8311, new_n8312, new_n8313, new_n8314, new_n8315, new_n8316,
    new_n8317, new_n8318, new_n8319, new_n8320, new_n8321, new_n8322,
    new_n8323, new_n8324, new_n8325, new_n8326, new_n8327, new_n8328,
    new_n8329, new_n8330, new_n8331, new_n8332, new_n8333, new_n8334,
    new_n8335, new_n8336, new_n8337, new_n8338, new_n8339, new_n8340,
    new_n8341, new_n8342, new_n8343, new_n8344, new_n8345, new_n8346,
    new_n8347, new_n8348, new_n8349, new_n8350, new_n8351, new_n8352,
    new_n8353, new_n8354, new_n8355, new_n8356, new_n8357, new_n8358,
    new_n8359, new_n8360, new_n8361, new_n8362, new_n8363, new_n8364,
    new_n8365, new_n8366, new_n8367, new_n8368, new_n8369, new_n8370,
    new_n8371, new_n8372, new_n8373, new_n8374, new_n8375, new_n8376,
    new_n8377, new_n8378, new_n8379, new_n8380, new_n8381, new_n8382,
    new_n8383, new_n8384, new_n8385, new_n8386, new_n8387, new_n8388,
    new_n8389, new_n8390, new_n8391, new_n8392, new_n8393, new_n8394,
    new_n8395, new_n8396, new_n8397, new_n8398, new_n8399, new_n8400,
    new_n8401, new_n8402, new_n8403, new_n8404, new_n8405, new_n8406,
    new_n8407, new_n8408, new_n8409, new_n8410, new_n8411, new_n8412,
    new_n8413, new_n8414, new_n8415, new_n8416, new_n8417, new_n8418,
    new_n8419, new_n8420, new_n8421, new_n8422, new_n8423, new_n8424,
    new_n8425, new_n8426, new_n8427, new_n8428, new_n8429, new_n8430,
    new_n8431, new_n8432, new_n8433, new_n8434, new_n8435, new_n8436,
    new_n8437, new_n8438, new_n8439, new_n8440, new_n8441, new_n8442,
    new_n8443, new_n8444, new_n8445, new_n8446, new_n8447, new_n8448,
    new_n8449, new_n8450, new_n8451, new_n8452, new_n8453, new_n8454,
    new_n8455, new_n8456, new_n8457, new_n8458, new_n8459, new_n8460,
    new_n8461, new_n8462, new_n8463, new_n8464, new_n8465, new_n8466,
    new_n8467, new_n8468, new_n8469, new_n8470, new_n8471, new_n8472,
    new_n8473, new_n8474, new_n8475, new_n8476, new_n8477, new_n8478,
    new_n8479, new_n8480, new_n8481, new_n8482, new_n8483, new_n8484,
    new_n8485, new_n8486, new_n8487, new_n8488, new_n8489, new_n8490,
    new_n8491, new_n8492, new_n8493, new_n8494, new_n8495, new_n8496,
    new_n8497, new_n8498, new_n8499, new_n8500, new_n8501, new_n8502,
    new_n8503, new_n8504, new_n8505, new_n8506, new_n8507, new_n8508,
    new_n8509, new_n8510, new_n8511, new_n8512, new_n8513, new_n8514,
    new_n8515, new_n8516, new_n8517, new_n8518, new_n8519, new_n8520,
    new_n8521, new_n8522, new_n8523, new_n8524, new_n8525, new_n8526,
    new_n8527, new_n8528, new_n8529, new_n8530, new_n8531, new_n8532,
    new_n8533, new_n8534, new_n8535, new_n8536, new_n8537, new_n8538,
    new_n8539, new_n8540, new_n8541, new_n8542, new_n8543, new_n8544,
    new_n8545, new_n8546, new_n8547, new_n8548, new_n8549, new_n8550,
    new_n8551, new_n8552, new_n8553, new_n8554, new_n8555, new_n8556,
    new_n8557, new_n8558, new_n8559, new_n8560, new_n8561, new_n8562,
    new_n8563, new_n8564, new_n8565, new_n8566, new_n8567, new_n8568,
    new_n8569, new_n8570, new_n8571, new_n8572, new_n8573, new_n8574,
    new_n8575, new_n8576, new_n8577, new_n8578, new_n8579, new_n8580,
    new_n8581, new_n8582, new_n8583, new_n8584, new_n8585, new_n8586,
    new_n8587, new_n8588, new_n8589, new_n8590, new_n8591, new_n8592,
    new_n8593, new_n8594, new_n8595, new_n8596, new_n8597, new_n8598,
    new_n8599, new_n8600, new_n8601, new_n8602, new_n8603, new_n8604,
    new_n8605, new_n8606, new_n8607, new_n8608, new_n8609, new_n8610,
    new_n8611, new_n8612, new_n8613, new_n8614, new_n8615, new_n8616,
    new_n8617, new_n8618, new_n8619, new_n8620, new_n8621, new_n8622,
    new_n8623, new_n8624, new_n8625, new_n8626, new_n8627, new_n8628,
    new_n8629, new_n8630, new_n8631, new_n8632, new_n8633, new_n8634,
    new_n8635, new_n8636, new_n8637, new_n8638, new_n8639, new_n8640,
    new_n8641, new_n8642, new_n8643, new_n8644, new_n8645, new_n8646,
    new_n8647, new_n8648, new_n8649, new_n8650, new_n8651, new_n8652,
    new_n8653, new_n8654, new_n8655, new_n8656, new_n8657, new_n8658,
    new_n8659, new_n8660, new_n8661, new_n8662, new_n8663, new_n8664,
    new_n8665, new_n8666, new_n8667, new_n8668, new_n8669, new_n8670,
    new_n8671, new_n8672, new_n8673, new_n8674, new_n8675, new_n8676,
    new_n8677, new_n8678, new_n8679, new_n8680, new_n8681, new_n8682,
    new_n8683, new_n8684, new_n8685, new_n8686, new_n8687, new_n8688,
    new_n8689, new_n8690, new_n8691, new_n8692, new_n8693, new_n8694,
    new_n8695, new_n8696, new_n8697, new_n8698, new_n8699, new_n8700,
    new_n8701, new_n8702, new_n8703, new_n8704, new_n8705, new_n8706,
    new_n8707, new_n8708, new_n8709, new_n8710, new_n8711, new_n8712,
    new_n8713, new_n8714, new_n8715, new_n8716, new_n8717, new_n8718,
    new_n8719, new_n8720, new_n8721, new_n8722, new_n8723, new_n8724,
    new_n8725, new_n8726, new_n8727, new_n8728, new_n8729, new_n8730,
    new_n8731, new_n8732, new_n8733, new_n8734, new_n8735, new_n8736,
    new_n8737, new_n8738, new_n8739, new_n8740, new_n8741, new_n8742,
    new_n8743, new_n8744, new_n8745, new_n8746, new_n8747, new_n8748,
    new_n8749, new_n8750, new_n8751, new_n8752, new_n8753, new_n8754,
    new_n8755, new_n8756, new_n8757, new_n8758, new_n8759, new_n8760,
    new_n8761, new_n8762, new_n8763, new_n8764, new_n8765, new_n8766,
    new_n8767, new_n8768, new_n8769, new_n8770, new_n8771, new_n8772,
    new_n8773, new_n8774, new_n8775, new_n8776, new_n8777, new_n8778,
    new_n8779, new_n8780, new_n8781, new_n8782, new_n8783, new_n8784,
    new_n8785, new_n8786, new_n8787, new_n8788, new_n8789, new_n8790,
    new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796,
    new_n8797, new_n8798, new_n8799, new_n8800, new_n8801, new_n8802,
    new_n8803, new_n8804, new_n8805, new_n8806, new_n8807, new_n8808,
    new_n8809, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814,
    new_n8815, new_n8816, new_n8817, new_n8818, new_n8819, new_n8820,
    new_n8821, new_n8822, new_n8823, new_n8824, new_n8825, new_n8826,
    new_n8827, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832,
    new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838,
    new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844,
    new_n8845, new_n8846, new_n8847, new_n8848, new_n8849, new_n8850,
    new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856,
    new_n8857, new_n8858, new_n8859, new_n8860, new_n8861, new_n8862,
    new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868,
    new_n8869, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874,
    new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880,
    new_n8881, new_n8882, new_n8883, new_n8884, new_n8885, new_n8886,
    new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8908, new_n8909, new_n8910,
    new_n8911, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042,
    new_n9043, new_n9044, new_n9045, new_n9046, new_n9047, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9060,
    new_n9061, new_n9062, new_n9063, new_n9064, new_n9065, new_n9066,
    new_n9067, new_n9068, new_n9069, new_n9070, new_n9071, new_n9072,
    new_n9073, new_n9074, new_n9075, new_n9076, new_n9077, new_n9078,
    new_n9079, new_n9080, new_n9081, new_n9082, new_n9083, new_n9084,
    new_n9085, new_n9086, new_n9087, new_n9088, new_n9089, new_n9090,
    new_n9091, new_n9092, new_n9093, new_n9094, new_n9095, new_n9096,
    new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102,
    new_n9103, new_n9104, new_n9105, new_n9106, new_n9107, new_n9108,
    new_n9109, new_n9110, new_n9111, new_n9112, new_n9113, new_n9114,
    new_n9115, new_n9116, new_n9117, new_n9118, new_n9119, new_n9120,
    new_n9121, new_n9122, new_n9123, new_n9124, new_n9125, new_n9126,
    new_n9127, new_n9128, new_n9129, new_n9130, new_n9131, new_n9132,
    new_n9133, new_n9134, new_n9135, new_n9136, new_n9137, new_n9138,
    new_n9139, new_n9140, new_n9141, new_n9142, new_n9143, new_n9144,
    new_n9145, new_n9146, new_n9147, new_n9148, new_n9149, new_n9150,
    new_n9151, new_n9152, new_n9153, new_n9154, new_n9155, new_n9156,
    new_n9157, new_n9158, new_n9159, new_n9160, new_n9161, new_n9162,
    new_n9163, new_n9164, new_n9165, new_n9166, new_n9167, new_n9168,
    new_n9169, new_n9170, new_n9171, new_n9172, new_n9173, new_n9174,
    new_n9175, new_n9176, new_n9177, new_n9178, new_n9179, new_n9180,
    new_n9181, new_n9182, new_n9183, new_n9184, new_n9185, new_n9186,
    new_n9187, new_n9188, new_n9189, new_n9190, new_n9191, new_n9192,
    new_n9193, new_n9194, new_n9195, new_n9196, new_n9197, new_n9198,
    new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204,
    new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210,
    new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216,
    new_n9217, new_n9218, new_n9219, new_n9220, new_n9221, new_n9222,
    new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228,
    new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234,
    new_n9235, new_n9236, new_n9237, new_n9238, new_n9239, new_n9240,
    new_n9241, new_n9242, new_n9243, new_n9244, new_n9245, new_n9246,
    new_n9247, new_n9248, new_n9249, new_n9250, new_n9251, new_n9252,
    new_n9253, new_n9254, new_n9255, new_n9256, new_n9257, new_n9258,
    new_n9259, new_n9260, new_n9261, new_n9262, new_n9263, new_n9264,
    new_n9265, new_n9266, new_n9267, new_n9268, new_n9269, new_n9270,
    new_n9271, new_n9272, new_n9273, new_n9274, new_n9275, new_n9276,
    new_n9277, new_n9278, new_n9279, new_n9280, new_n9281, new_n9282,
    new_n9283, new_n9284, new_n9285, new_n9286, new_n9287, new_n9288,
    new_n9289, new_n9290, new_n9291, new_n9292, new_n9293, new_n9294,
    new_n9295, new_n9296, new_n9297, new_n9298, new_n9299, new_n9300,
    new_n9301, new_n9302, new_n9303, new_n9304, new_n9305, new_n9306,
    new_n9307, new_n9308, new_n9309, new_n9310, new_n9311, new_n9312,
    new_n9313, new_n9314, new_n9315, new_n9316, new_n9317, new_n9318,
    new_n9319, new_n9320, new_n9321, new_n9322, new_n9323, new_n9324,
    new_n9325, new_n9326, new_n9327, new_n9328, new_n9329, new_n9330,
    new_n9331, new_n9332, new_n9333, new_n9334, new_n9335, new_n9336,
    new_n9337, new_n9338, new_n9339, new_n9340, new_n9341, new_n9342,
    new_n9343, new_n9344, new_n9345, new_n9346, new_n9347, new_n9348,
    new_n9349, new_n9350, new_n9351, new_n9352, new_n9353, new_n9354,
    new_n9355, new_n9356, new_n9357, new_n9358, new_n9359, new_n9360,
    new_n9361, new_n9362, new_n9363, new_n9364, new_n9365, new_n9366,
    new_n9367, new_n9368, new_n9369, new_n9370, new_n9371, new_n9372,
    new_n9373, new_n9374, new_n9375, new_n9376, new_n9377, new_n9378,
    new_n9379, new_n9380, new_n9381, new_n9382, new_n9383, new_n9384,
    new_n9385, new_n9386, new_n9387, new_n9388, new_n9389, new_n9390,
    new_n9391, new_n9392, new_n9393, new_n9394, new_n9395, new_n9396,
    new_n9397, new_n9398, new_n9399, new_n9400, new_n9401, new_n9402,
    new_n9403, new_n9404, new_n9405, new_n9406, new_n9407, new_n9408,
    new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414,
    new_n9415, new_n9416, new_n9417, new_n9418, new_n9419, new_n9420,
    new_n9421, new_n9422, new_n9423, new_n9424, new_n9425, new_n9426,
    new_n9427, new_n9428, new_n9429, new_n9430, new_n9431, new_n9432,
    new_n9433, new_n9434, new_n9435, new_n9436, new_n9437, new_n9438,
    new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444,
    new_n9445, new_n9446, new_n9447, new_n9448, new_n9449, new_n9450,
    new_n9451, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456,
    new_n9457, new_n9458, new_n9459, new_n9460, new_n9461, new_n9462,
    new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468,
    new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9474,
    new_n9475, new_n9476, new_n9477, new_n9478, new_n9479, new_n9480,
    new_n9481, new_n9482, new_n9483, new_n9484, new_n9485, new_n9486,
    new_n9487, new_n9488, new_n9489, new_n9490, new_n9491, new_n9492,
    new_n9493, new_n9494, new_n9495, new_n9496, new_n9497, new_n9498,
    new_n9499, new_n9500, new_n9501, new_n9502, new_n9503, new_n9504,
    new_n9505, new_n9506, new_n9507, new_n9508, new_n9509, new_n9510,
    new_n9511, new_n9512, new_n9513, new_n9514, new_n9515, new_n9516,
    new_n9517, new_n9518, new_n9519, new_n9520, new_n9521, new_n9522,
    new_n9523, new_n9524, new_n9525, new_n9526, new_n9527, new_n9528,
    new_n9529, new_n9530, new_n9531, new_n9532, new_n9533, new_n9534,
    new_n9535, new_n9536, new_n9537, new_n9538, new_n9539, new_n9540,
    new_n9541, new_n9542, new_n9543, new_n9544, new_n9545, new_n9546,
    new_n9547, new_n9548, new_n9549, new_n9550, new_n9551, new_n9552,
    new_n9553, new_n9554, new_n9555, new_n9556, new_n9557, new_n9558,
    new_n9559, new_n9560, new_n9561, new_n9562, new_n9563, new_n9564,
    new_n9565, new_n9566, new_n9567, new_n9568, new_n9569, new_n9570,
    new_n9571, new_n9572, new_n9573, new_n9574, new_n9575, new_n9576,
    new_n9577, new_n9578, new_n9579, new_n9580, new_n9581, new_n9582,
    new_n9583, new_n9584, new_n9585, new_n9586, new_n9587, new_n9588,
    new_n9589, new_n9590, new_n9591, new_n9592, new_n9593, new_n9594,
    new_n9595, new_n9596, new_n9597, new_n9598, new_n9599, new_n9600,
    new_n9601, new_n9602, new_n9603, new_n9604, new_n9605, new_n9606,
    new_n9607, new_n9608, new_n9609, new_n9610, new_n9611, new_n9612,
    new_n9613, new_n9614, new_n9615, new_n9616, new_n9617, new_n9618,
    new_n9619, new_n9620, new_n9621, new_n9622, new_n9623, new_n9624,
    new_n9625, new_n9626, new_n9627, new_n9628, new_n9629, new_n9630,
    new_n9631, new_n9632, new_n9633, new_n9634, new_n9635, new_n9636,
    new_n9637, new_n9638, new_n9639, new_n9640, new_n9641, new_n9642,
    new_n9643, new_n9644, new_n9645, new_n9646, new_n9647, new_n9648,
    new_n9649, new_n9650, new_n9651, new_n9652, new_n9653, new_n9654,
    new_n9655, new_n9656, new_n9657, new_n9658, new_n9659, new_n9660,
    new_n9661, new_n9662, new_n9663, new_n9664, new_n9665, new_n9666,
    new_n9667, new_n9668, new_n9669, new_n9670, new_n9671, new_n9672,
    new_n9673, new_n9674, new_n9675, new_n9676, new_n9677, new_n9678,
    new_n9679, new_n9680, new_n9681, new_n9682, new_n9683, new_n9684,
    new_n9685, new_n9686, new_n9687, new_n9688, new_n9689, new_n9690,
    new_n9691, new_n9692, new_n9693, new_n9694, new_n9695, new_n9696,
    new_n9697, new_n9698, new_n9699, new_n9700, new_n9701, new_n9702,
    new_n9703, new_n9704, new_n9705, new_n9706, new_n9707, new_n9708,
    new_n9709, new_n9710, new_n9711, new_n9712, new_n9713, new_n9714,
    new_n9715, new_n9716, new_n9717, new_n9718, new_n9719, new_n9720,
    new_n9721, new_n9722, new_n9723, new_n9724, new_n9725, new_n9726,
    new_n9727, new_n9728, new_n9729, new_n9730, new_n9731, new_n9732,
    new_n9733, new_n9734, new_n9735, new_n9736, new_n9737, new_n9738,
    new_n9739, new_n9740, new_n9741, new_n9742, new_n9743, new_n9744,
    new_n9745, new_n9746, new_n9747, new_n9748, new_n9749, new_n9750,
    new_n9751, new_n9752, new_n9753, new_n9754, new_n9755, new_n9756,
    new_n9757, new_n9758, new_n9759, new_n9760, new_n9761, new_n9762,
    new_n9763, new_n9764, new_n9765, new_n9766, new_n9767, new_n9768,
    new_n9769, new_n9770, new_n9771, new_n9772, new_n9773, new_n9774,
    new_n9775, new_n9776, new_n9777, new_n9778, new_n9779, new_n9780,
    new_n9781, new_n9782, new_n9783, new_n9784, new_n9785, new_n9786,
    new_n9787, new_n9788, new_n9789, new_n9790, new_n9791, new_n9792,
    new_n9793, new_n9794, new_n9795, new_n9796, new_n9797, new_n9798,
    new_n9799, new_n9800, new_n9801, new_n9802, new_n9803, new_n9804,
    new_n9805, new_n9806, new_n9807, new_n9808, new_n9809, new_n9810,
    new_n9811, new_n9812, new_n9813, new_n9814, new_n9815, new_n9816,
    new_n9817, new_n9818, new_n9819, new_n9820, new_n9821, new_n9822,
    new_n9823, new_n9824, new_n9825, new_n9826, new_n9827, new_n9828,
    new_n9829, new_n9830, new_n9831, new_n9832, new_n9833, new_n9834,
    new_n9835, new_n9836, new_n9837, new_n9838, new_n9839, new_n9840,
    new_n9841, new_n9842, new_n9843, new_n9844, new_n9845, new_n9846,
    new_n9847, new_n9848, new_n9849, new_n9850, new_n9851, new_n9852,
    new_n9853, new_n9854, new_n9855, new_n9856, new_n9857, new_n9858,
    new_n9859, new_n9860, new_n9861, new_n9862, new_n9863, new_n9864,
    new_n9865, new_n9866, new_n9867, new_n9868, new_n9869, new_n9870,
    new_n9871, new_n9872, new_n9873, new_n9874, new_n9875, new_n9876,
    new_n9877, new_n9878, new_n9879, new_n9880, new_n9881, new_n9882,
    new_n9883, new_n9884, new_n9885, new_n9886, new_n9887, new_n9888,
    new_n9889, new_n9890, new_n9891, new_n9892, new_n9893, new_n9894,
    new_n9895, new_n9896, new_n9897, new_n9898, new_n9899, new_n9900,
    new_n9901, new_n9902, new_n9903, new_n9904, new_n9905, new_n9906,
    new_n9907, new_n9908, new_n9909, new_n9910, new_n9911, new_n9912,
    new_n9913, new_n9914, new_n9915, new_n9916, new_n9917, new_n9918,
    new_n9919, new_n9920, new_n9921, new_n9922, new_n9923, new_n9924,
    new_n9925, new_n9926, new_n9927, new_n9928, new_n9929, new_n9930,
    new_n9931, new_n9932, new_n9933, new_n9934, new_n9935, new_n9936,
    new_n9937, new_n9938, new_n9939, new_n9940, new_n9941, new_n9942,
    new_n9943, new_n9944, new_n9945, new_n9946, new_n9947, new_n9948,
    new_n9949, new_n9950, new_n9951, new_n9952, new_n9953, new_n9954,
    new_n9955, new_n9956, new_n9957, new_n9958, new_n9959, new_n9960,
    new_n9961, new_n9962, new_n9963, new_n9964, new_n9965, new_n9966,
    new_n9967, new_n9968, new_n9969, new_n9970, new_n9971, new_n9972,
    new_n9973, new_n9974, new_n9975, new_n9976, new_n9977, new_n9978,
    new_n9979, new_n9980, new_n9981, new_n9982, new_n9983, new_n9984,
    new_n9985, new_n9986, new_n9987, new_n9988, new_n9989, new_n9990,
    new_n9991, new_n9992, new_n9993, new_n9994, new_n9995, new_n9996,
    new_n9997, new_n9998, new_n9999, new_n10000, new_n10001, new_n10002,
    new_n10003, new_n10004, new_n10005, new_n10006, new_n10007, new_n10008,
    new_n10009, new_n10010, new_n10011, new_n10012, new_n10013, new_n10014,
    new_n10015, new_n10016, new_n10017, new_n10018, new_n10019, new_n10020,
    new_n10021, new_n10022, new_n10023, new_n10024, new_n10025, new_n10026,
    new_n10027, new_n10028, new_n10029, new_n10030, new_n10031, new_n10032,
    new_n10033, new_n10034, new_n10035, new_n10036, new_n10037, new_n10038,
    new_n10039, new_n10040, new_n10041, new_n10042, new_n10043, new_n10044,
    new_n10045, new_n10046, new_n10047, new_n10048, new_n10049, new_n10050,
    new_n10051, new_n10052, new_n10053, new_n10054, new_n10055, new_n10056,
    new_n10057, new_n10058, new_n10059, new_n10060, new_n10061, new_n10062,
    new_n10063, new_n10064, new_n10065, new_n10066, new_n10067, new_n10068,
    new_n10069, new_n10070, new_n10071, new_n10072, new_n10073, new_n10074,
    new_n10075, new_n10076, new_n10077, new_n10078, new_n10079, new_n10080,
    new_n10081, new_n10082, new_n10083, new_n10084, new_n10085, new_n10086,
    new_n10087, new_n10088, new_n10089, new_n10090, new_n10091, new_n10092,
    new_n10093, new_n10094, new_n10095, new_n10096, new_n10097, new_n10098,
    new_n10099, new_n10100, new_n10101, new_n10102, new_n10103, new_n10104,
    new_n10105, new_n10106, new_n10107, new_n10108, new_n10109, new_n10110,
    new_n10111, new_n10112, new_n10113, new_n10114, new_n10115, new_n10116,
    new_n10117, new_n10118, new_n10119, new_n10120, new_n10121, new_n10122,
    new_n10123, new_n10124, new_n10125, new_n10126, new_n10127, new_n10128,
    new_n10129, new_n10130, new_n10131, new_n10132, new_n10133, new_n10134,
    new_n10135, new_n10136, new_n10137, new_n10138, new_n10139, new_n10140,
    new_n10141, new_n10142, new_n10143, new_n10144, new_n10145, new_n10146,
    new_n10147, new_n10148, new_n10149, new_n10150, new_n10151, new_n10152,
    new_n10153, new_n10154, new_n10155, new_n10156, new_n10157, new_n10158,
    new_n10159, new_n10160, new_n10161, new_n10162, new_n10163, new_n10164,
    new_n10165, new_n10166, new_n10167, new_n10168, new_n10169, new_n10170,
    new_n10171, new_n10172, new_n10173, new_n10174, new_n10175, new_n10176,
    new_n10177, new_n10178, new_n10179, new_n10180, new_n10181, new_n10182,
    new_n10183, new_n10184, new_n10185, new_n10186, new_n10187, new_n10188,
    new_n10189, new_n10190, new_n10191, new_n10192, new_n10193, new_n10194,
    new_n10195, new_n10196, new_n10197, new_n10198, new_n10199, new_n10200,
    new_n10201, new_n10202, new_n10203, new_n10204, new_n10205, new_n10206,
    new_n10207, new_n10208, new_n10209, new_n10210, new_n10211, new_n10212,
    new_n10213, new_n10214, new_n10215, new_n10216, new_n10217, new_n10218,
    new_n10219, new_n10220, new_n10221, new_n10222, new_n10223, new_n10224,
    new_n10225, new_n10226, new_n10227, new_n10228, new_n10229, new_n10230,
    new_n10231, new_n10232, new_n10233, new_n10234, new_n10235, new_n10236,
    new_n10237, new_n10238, new_n10239, new_n10240, new_n10241, new_n10242,
    new_n10243, new_n10244, new_n10245, new_n10246, new_n10247, new_n10248,
    new_n10249, new_n10250, new_n10251, new_n10252, new_n10253, new_n10254,
    new_n10255, new_n10256, new_n10257, new_n10258, new_n10259, new_n10260,
    new_n10261, new_n10262, new_n10263, new_n10264, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10275, new_n10276, new_n10277, new_n10278,
    new_n10279, new_n10280, new_n10281, new_n10282, new_n10283, new_n10284,
    new_n10285, new_n10286, new_n10287, new_n10288, new_n10289, new_n10290,
    new_n10291, new_n10292, new_n10293, new_n10294, new_n10295, new_n10296,
    new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302,
    new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308,
    new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314,
    new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320,
    new_n10321, new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327, new_n10328, new_n10329, new_n10330, new_n10331, new_n10332,
    new_n10333, new_n10334, new_n10335, new_n10336, new_n10337, new_n10338,
    new_n10339, new_n10340, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345, new_n10346, new_n10347, new_n10348, new_n10349, new_n10350,
    new_n10351, new_n10352, new_n10353, new_n10354, new_n10355, new_n10356,
    new_n10357, new_n10358, new_n10359, new_n10360, new_n10361, new_n10362,
    new_n10363, new_n10364, new_n10365, new_n10366, new_n10367, new_n10368,
    new_n10369, new_n10370, new_n10371, new_n10372, new_n10373, new_n10374,
    new_n10375, new_n10376, new_n10377, new_n10378, new_n10379, new_n10380,
    new_n10381, new_n10382, new_n10383, new_n10384, new_n10385, new_n10386,
    new_n10387, new_n10388, new_n10389, new_n10390, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403, new_n10404,
    new_n10405, new_n10406, new_n10407, new_n10408, new_n10409, new_n10410,
    new_n10411, new_n10412, new_n10413, new_n10414, new_n10415, new_n10416,
    new_n10417, new_n10418, new_n10419, new_n10420, new_n10421, new_n10422,
    new_n10423, new_n10424, new_n10425, new_n10426, new_n10427, new_n10428,
    new_n10429, new_n10430, new_n10431, new_n10432, new_n10433, new_n10434,
    new_n10435, new_n10436, new_n10437, new_n10438, new_n10439, new_n10440,
    new_n10441, new_n10442, new_n10443, new_n10444, new_n10445, new_n10446,
    new_n10447, new_n10448, new_n10449, new_n10450, new_n10451, new_n10452,
    new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458,
    new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464,
    new_n10465, new_n10466, new_n10467, new_n10468, new_n10469, new_n10470,
    new_n10471, new_n10472, new_n10473, new_n10474, new_n10475, new_n10476,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510, new_n10511, new_n10512,
    new_n10513, new_n10514, new_n10515, new_n10516, new_n10517, new_n10518,
    new_n10519, new_n10520, new_n10521, new_n10522, new_n10523, new_n10524,
    new_n10525, new_n10526, new_n10527, new_n10528, new_n10529, new_n10530,
    new_n10531, new_n10532, new_n10533, new_n10534, new_n10535, new_n10536,
    new_n10537, new_n10538, new_n10539, new_n10540, new_n10541, new_n10542,
    new_n10543, new_n10544, new_n10545, new_n10546, new_n10547, new_n10548,
    new_n10549, new_n10550, new_n10551, new_n10552, new_n10553, new_n10554,
    new_n10555, new_n10556, new_n10557, new_n10558, new_n10559, new_n10560,
    new_n10561, new_n10562, new_n10563, new_n10564, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572,
    new_n10573, new_n10574, new_n10575, new_n10576, new_n10577, new_n10578,
    new_n10579, new_n10580, new_n10581, new_n10582, new_n10583, new_n10584,
    new_n10585, new_n10586, new_n10587, new_n10588, new_n10589, new_n10590,
    new_n10591, new_n10592, new_n10593, new_n10594, new_n10595, new_n10596,
    new_n10597, new_n10598, new_n10599, new_n10600, new_n10601, new_n10602,
    new_n10603, new_n10604, new_n10605, new_n10606, new_n10607, new_n10608,
    new_n10609, new_n10610, new_n10611, new_n10612, new_n10613, new_n10614,
    new_n10615, new_n10616, new_n10617, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628, new_n10629, new_n10630, new_n10631, new_n10632,
    new_n10633, new_n10634, new_n10635, new_n10636, new_n10637, new_n10638,
    new_n10639, new_n10640, new_n10641, new_n10642, new_n10643, new_n10644,
    new_n10645, new_n10646, new_n10647, new_n10648, new_n10649, new_n10650,
    new_n10651, new_n10652, new_n10653, new_n10654, new_n10655, new_n10656,
    new_n10657, new_n10658, new_n10659, new_n10660, new_n10661, new_n10662,
    new_n10663, new_n10664, new_n10665, new_n10666, new_n10667, new_n10668,
    new_n10669, new_n10670, new_n10671, new_n10672, new_n10673, new_n10674,
    new_n10675, new_n10676, new_n10677, new_n10678, new_n10679, new_n10680,
    new_n10681, new_n10682, new_n10683, new_n10684, new_n10685, new_n10686,
    new_n10687, new_n10688, new_n10689, new_n10690, new_n10691, new_n10692,
    new_n10693, new_n10694, new_n10695, new_n10696, new_n10697, new_n10698,
    new_n10699, new_n10700, new_n10701, new_n10702, new_n10703, new_n10704,
    new_n10705, new_n10706, new_n10707, new_n10708, new_n10709, new_n10710,
    new_n10711, new_n10712, new_n10713, new_n10714, new_n10715, new_n10716,
    new_n10717, new_n10718, new_n10719, new_n10720, new_n10721, new_n10722,
    new_n10723, new_n10724, new_n10725, new_n10726, new_n10727, new_n10728,
    new_n10729, new_n10730, new_n10731, new_n10732, new_n10733, new_n10734,
    new_n10735, new_n10736, new_n10737, new_n10738, new_n10739, new_n10740,
    new_n10741, new_n10742, new_n10743, new_n10744, new_n10745, new_n10746,
    new_n10747, new_n10748, new_n10749, new_n10750, new_n10751, new_n10752,
    new_n10753, new_n10754, new_n10755, new_n10756, new_n10757, new_n10758,
    new_n10759, new_n10760, new_n10761, new_n10762, new_n10763, new_n10764,
    new_n10765, new_n10766, new_n10767, new_n10768, new_n10769, new_n10770,
    new_n10771, new_n10772, new_n10773, new_n10774, new_n10775, new_n10776,
    new_n10777, new_n10778, new_n10779, new_n10780, new_n10781, new_n10782,
    new_n10783, new_n10784, new_n10785, new_n10786, new_n10787, new_n10788,
    new_n10789, new_n10790, new_n10791, new_n10792, new_n10793, new_n10794,
    new_n10795, new_n10796, new_n10797, new_n10798, new_n10799, new_n10800,
    new_n10801, new_n10802, new_n10803, new_n10804, new_n10805, new_n10806,
    new_n10807, new_n10808, new_n10809, new_n10810, new_n10811, new_n10812,
    new_n10813, new_n10814, new_n10815, new_n10816, new_n10817, new_n10818,
    new_n10819, new_n10820, new_n10821, new_n10822, new_n10823, new_n10824,
    new_n10825, new_n10826, new_n10827, new_n10828, new_n10829, new_n10830,
    new_n10831, new_n10832, new_n10833, new_n10834, new_n10835, new_n10836,
    new_n10837, new_n10838, new_n10839, new_n10840, new_n10841, new_n10842,
    new_n10843, new_n10844, new_n10845, new_n10846, new_n10847, new_n10848,
    new_n10849, new_n10850, new_n10851, new_n10852, new_n10853, new_n10854,
    new_n10855, new_n10856, new_n10857, new_n10858, new_n10859, new_n10860,
    new_n10861, new_n10862, new_n10863, new_n10864, new_n10865, new_n10866,
    new_n10867, new_n10868, new_n10869, new_n10870, new_n10871, new_n10872,
    new_n10873, new_n10874, new_n10875, new_n10876, new_n10877, new_n10878,
    new_n10879, new_n10880, new_n10881, new_n10882, new_n10883, new_n10884,
    new_n10885, new_n10886, new_n10887, new_n10888, new_n10889, new_n10890,
    new_n10891, new_n10892, new_n10893, new_n10894, new_n10895, new_n10896,
    new_n10897, new_n10898, new_n10899, new_n10900, new_n10901, new_n10902,
    new_n10903, new_n10904, new_n10905, new_n10906, new_n10907, new_n10908,
    new_n10909, new_n10910, new_n10911, new_n10912, new_n10913, new_n10914,
    new_n10915, new_n10916, new_n10917, new_n10918, new_n10919, new_n10920,
    new_n10921, new_n10922, new_n10923, new_n10924, new_n10925, new_n10926,
    new_n10927, new_n10928, new_n10929, new_n10930, new_n10931, new_n10932,
    new_n10933, new_n10934, new_n10935, new_n10936, new_n10937, new_n10938,
    new_n10939, new_n10940, new_n10941, new_n10942, new_n10943, new_n10944,
    new_n10945, new_n10946, new_n10947, new_n10948, new_n10949, new_n10950,
    new_n10951, new_n10952, new_n10953, new_n10954, new_n10955, new_n10956,
    new_n10957, new_n10958, new_n10959, new_n10960, new_n10961, new_n10962,
    new_n10963, new_n10964, new_n10965, new_n10966, new_n10967, new_n10968,
    new_n10969, new_n10970, new_n10971, new_n10972, new_n10973, new_n10974,
    new_n10975, new_n10976, new_n10977, new_n10978, new_n10979, new_n10980,
    new_n10981, new_n10982, new_n10983, new_n10984, new_n10985, new_n10986,
    new_n10987, new_n10988, new_n10989, new_n10990, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005, new_n11006, new_n11007, new_n11008, new_n11009, new_n11010,
    new_n11011, new_n11012, new_n11013, new_n11014, new_n11015, new_n11016,
    new_n11017, new_n11018, new_n11019, new_n11020, new_n11021, new_n11022,
    new_n11023, new_n11024, new_n11025, new_n11026, new_n11027, new_n11028,
    new_n11029, new_n11030, new_n11031, new_n11032, new_n11033, new_n11034,
    new_n11035, new_n11036, new_n11037, new_n11038, new_n11039, new_n11040,
    new_n11041, new_n11042, new_n11043, new_n11044, new_n11045, new_n11046,
    new_n11047, new_n11048, new_n11049, new_n11050, new_n11051, new_n11052,
    new_n11053, new_n11054, new_n11055, new_n11056, new_n11057, new_n11058,
    new_n11059, new_n11060, new_n11061, new_n11062, new_n11063, new_n11064,
    new_n11065, new_n11066, new_n11067, new_n11068, new_n11069, new_n11070,
    new_n11071, new_n11072, new_n11073, new_n11074, new_n11075, new_n11076,
    new_n11077, new_n11078, new_n11079, new_n11080, new_n11081, new_n11082,
    new_n11083, new_n11084, new_n11085, new_n11086, new_n11087, new_n11088,
    new_n11089, new_n11090, new_n11091, new_n11092, new_n11093, new_n11094,
    new_n11095, new_n11096, new_n11097, new_n11098, new_n11099, new_n11100,
    new_n11101, new_n11102, new_n11103, new_n11104, new_n11105, new_n11106,
    new_n11107, new_n11108, new_n11109, new_n11110, new_n11111, new_n11112,
    new_n11113, new_n11114, new_n11115, new_n11116, new_n11117, new_n11118,
    new_n11119, new_n11120, new_n11121, new_n11122, new_n11123, new_n11124,
    new_n11125, new_n11126, new_n11127, new_n11128, new_n11129, new_n11130,
    new_n11131, new_n11132, new_n11133, new_n11134, new_n11135, new_n11136,
    new_n11137, new_n11138, new_n11139, new_n11140, new_n11141, new_n11142,
    new_n11143, new_n11144, new_n11145, new_n11146, new_n11147, new_n11148,
    new_n11149, new_n11150, new_n11151, new_n11152, new_n11153, new_n11154,
    new_n11155, new_n11156, new_n11157, new_n11158, new_n11159, new_n11160,
    new_n11161, new_n11162, new_n11163, new_n11164, new_n11165, new_n11166,
    new_n11167, new_n11168, new_n11169, new_n11170, new_n11171, new_n11172,
    new_n11173, new_n11174, new_n11175, new_n11176, new_n11177, new_n11178,
    new_n11179, new_n11180, new_n11181, new_n11182, new_n11183, new_n11184,
    new_n11185, new_n11186, new_n11187, new_n11188, new_n11189, new_n11190,
    new_n11191, new_n11192, new_n11193, new_n11194, new_n11195, new_n11196,
    new_n11197, new_n11198, new_n11199, new_n11200, new_n11201, new_n11202,
    new_n11203, new_n11204, new_n11205, new_n11206, new_n11207, new_n11208,
    new_n11209, new_n11210, new_n11211, new_n11212, new_n11213, new_n11214,
    new_n11215, new_n11216, new_n11217, new_n11218, new_n11219, new_n11220,
    new_n11221, new_n11222, new_n11223, new_n11224, new_n11225, new_n11226,
    new_n11227, new_n11228, new_n11229, new_n11230, new_n11231, new_n11232,
    new_n11233, new_n11234, new_n11235, new_n11236, new_n11237, new_n11238,
    new_n11239, new_n11240, new_n11241, new_n11242, new_n11243, new_n11244,
    new_n11245, new_n11246, new_n11247, new_n11248, new_n11249, new_n11250,
    new_n11251, new_n11252, new_n11253, new_n11254, new_n11255, new_n11256,
    new_n11257, new_n11258, new_n11259, new_n11260, new_n11261, new_n11262,
    new_n11263, new_n11264, new_n11265, new_n11266, new_n11267, new_n11268,
    new_n11269, new_n11270, new_n11271, new_n11272, new_n11273, new_n11274,
    new_n11275, new_n11276, new_n11277, new_n11278, new_n11279, new_n11280,
    new_n11281, new_n11282, new_n11283, new_n11284, new_n11285, new_n11286,
    new_n11287, new_n11288, new_n11289, new_n11290, new_n11291, new_n11292,
    new_n11293, new_n11294, new_n11295, new_n11296, new_n11297, new_n11298,
    new_n11299, new_n11300, new_n11301, new_n11302, new_n11303, new_n11304,
    new_n11305, new_n11306, new_n11307, new_n11308, new_n11309, new_n11310,
    new_n11311, new_n11312, new_n11313, new_n11314, new_n11315, new_n11316,
    new_n11317, new_n11318, new_n11319, new_n11320, new_n11321, new_n11322,
    new_n11323, new_n11324, new_n11325, new_n11326, new_n11327, new_n11328,
    new_n11329, new_n11330, new_n11331, new_n11332, new_n11333, new_n11334,
    new_n11335, new_n11336, new_n11337, new_n11338, new_n11339, new_n11340,
    new_n11341, new_n11342, new_n11343, new_n11344, new_n11345, new_n11346,
    new_n11347, new_n11348, new_n11349, new_n11350, new_n11351, new_n11352,
    new_n11353, new_n11354, new_n11355, new_n11356, new_n11357, new_n11358,
    new_n11359, new_n11360, new_n11361, new_n11362, new_n11363, new_n11364,
    new_n11365, new_n11366, new_n11367, new_n11368, new_n11369, new_n11370,
    new_n11371, new_n11372, new_n11373, new_n11374, new_n11375, new_n11376,
    new_n11377, new_n11378, new_n11379, new_n11380, new_n11381, new_n11382,
    new_n11383, new_n11384, new_n11385, new_n11386, new_n11387, new_n11388,
    new_n11389, new_n11390, new_n11391, new_n11392, new_n11393, new_n11394,
    new_n11395, new_n11396, new_n11397, new_n11398, new_n11399, new_n11400,
    new_n11401, new_n11402, new_n11403, new_n11404, new_n11405, new_n11406,
    new_n11407, new_n11408, new_n11409, new_n11410, new_n11411, new_n11412,
    new_n11413, new_n11414, new_n11415, new_n11416, new_n11417, new_n11418,
    new_n11419, new_n11420, new_n11421, new_n11422, new_n11423, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472,
    new_n11473, new_n11474, new_n11475, new_n11476, new_n11477, new_n11478,
    new_n11479, new_n11480, new_n11481, new_n11482, new_n11483, new_n11484,
    new_n11485, new_n11486, new_n11487, new_n11488, new_n11489, new_n11490,
    new_n11491, new_n11492, new_n11493, new_n11494, new_n11495, new_n11496,
    new_n11497, new_n11498, new_n11499, new_n11500, new_n11501, new_n11502,
    new_n11503, new_n11504, new_n11505, new_n11506, new_n11507, new_n11508,
    new_n11509, new_n11510, new_n11511, new_n11512, new_n11513, new_n11514,
    new_n11515, new_n11516, new_n11517, new_n11518, new_n11519, new_n11520,
    new_n11521, new_n11522, new_n11523, new_n11524, new_n11525, new_n11526,
    new_n11527, new_n11528, new_n11529, new_n11530, new_n11531, new_n11532,
    new_n11533, new_n11534, new_n11535, new_n11536, new_n11537, new_n11538,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548, new_n11549, new_n11550,
    new_n11551, new_n11552, new_n11553, new_n11554, new_n11555, new_n11556,
    new_n11557, new_n11558, new_n11559, new_n11560, new_n11561, new_n11562,
    new_n11563, new_n11564, new_n11565, new_n11566, new_n11567, new_n11568,
    new_n11569, new_n11570, new_n11571, new_n11572, new_n11573, new_n11574,
    new_n11575, new_n11576, new_n11577, new_n11578, new_n11579, new_n11580,
    new_n11581, new_n11582, new_n11583, new_n11584, new_n11585, new_n11586,
    new_n11587, new_n11588, new_n11589, new_n11590, new_n11591, new_n11592,
    new_n11593, new_n11594, new_n11595, new_n11596, new_n11597, new_n11598,
    new_n11599, new_n11600, new_n11601, new_n11602, new_n11603, new_n11604,
    new_n11605, new_n11606, new_n11607, new_n11608, new_n11609, new_n11610,
    new_n11611, new_n11612, new_n11613, new_n11614, new_n11615, new_n11616,
    new_n11617, new_n11618, new_n11619, new_n11620, new_n11621, new_n11622,
    new_n11623, new_n11624, new_n11625, new_n11626, new_n11627, new_n11628,
    new_n11629, new_n11630, new_n11631, new_n11632, new_n11633, new_n11634,
    new_n11635, new_n11636, new_n11637, new_n11638, new_n11639, new_n11640,
    new_n11641, new_n11642, new_n11643, new_n11644, new_n11645, new_n11646,
    new_n11647, new_n11648, new_n11649, new_n11650, new_n11651, new_n11652,
    new_n11653, new_n11654, new_n11655, new_n11656, new_n11657, new_n11658,
    new_n11659, new_n11660, new_n11661, new_n11662, new_n11663, new_n11664,
    new_n11665, new_n11666, new_n11667, new_n11668, new_n11669, new_n11670,
    new_n11671, new_n11672, new_n11673, new_n11674, new_n11675, new_n11676,
    new_n11677, new_n11678, new_n11679, new_n11680, new_n11681, new_n11682,
    new_n11683, new_n11684, new_n11685, new_n11686, new_n11687, new_n11688,
    new_n11689, new_n11690, new_n11691, new_n11692, new_n11693, new_n11694,
    new_n11695, new_n11696, new_n11697, new_n11698, new_n11699, new_n11700,
    new_n11701, new_n11702, new_n11703, new_n11704, new_n11705, new_n11706,
    new_n11707, new_n11708, new_n11709, new_n11710, new_n11711, new_n11712,
    new_n11713, new_n11714, new_n11715, new_n11716, new_n11717, new_n11718,
    new_n11719, new_n11720, new_n11721, new_n11722, new_n11723, new_n11724,
    new_n11725, new_n11726, new_n11727, new_n11728, new_n11729, new_n11730,
    new_n11731, new_n11732, new_n11733, new_n11734, new_n11735, new_n11736,
    new_n11737, new_n11738, new_n11739, new_n11740, new_n11741, new_n11742,
    new_n11743, new_n11744, new_n11745, new_n11746, new_n11747, new_n11748,
    new_n11749, new_n11750, new_n11751, new_n11752, new_n11753, new_n11754,
    new_n11755, new_n11756, new_n11757, new_n11758, new_n11759, new_n11760,
    new_n11761, new_n11762, new_n11763, new_n11764, new_n11765, new_n11766,
    new_n11767, new_n11768, new_n11769, new_n11770, new_n11771, new_n11772,
    new_n11773, new_n11774, new_n11775, new_n11776, new_n11777, new_n11778,
    new_n11779, new_n11780, new_n11781, new_n11782, new_n11783, new_n11784,
    new_n11785, new_n11786, new_n11787, new_n11788, new_n11789, new_n11790,
    new_n11791, new_n11792, new_n11793, new_n11794, new_n11795, new_n11796,
    new_n11797, new_n11798, new_n11799, new_n11800, new_n11801, new_n11802,
    new_n11803, new_n11804, new_n11805, new_n11806, new_n11807, new_n11808,
    new_n11809, new_n11810, new_n11811, new_n11812, new_n11813, new_n11814,
    new_n11815, new_n11816, new_n11817, new_n11818, new_n11819, new_n11820,
    new_n11821, new_n11822, new_n11823, new_n11824, new_n11825, new_n11826,
    new_n11827, new_n11828, new_n11829, new_n11830, new_n11831, new_n11832,
    new_n11833, new_n11834, new_n11835, new_n11836, new_n11837, new_n11838,
    new_n11839, new_n11840, new_n11841, new_n11842, new_n11843, new_n11844,
    new_n11845, new_n11846, new_n11847, new_n11848, new_n11849, new_n11850,
    new_n11851, new_n11852, new_n11853, new_n11854, new_n11855, new_n11856,
    new_n11857, new_n11858, new_n11859, new_n11860, new_n11861, new_n11862,
    new_n11863, new_n11864, new_n11865, new_n11866, new_n11867, new_n11868,
    new_n11869, new_n11870, new_n11871, new_n11872, new_n11873, new_n11874,
    new_n11875, new_n11876, new_n11877, new_n11878, new_n11879, new_n11880,
    new_n11881, new_n11882, new_n11883, new_n11884, new_n11885, new_n11886,
    new_n11887, new_n11888, new_n11889, new_n11890, new_n11891, new_n11892,
    new_n11893, new_n11894, new_n11895, new_n11896, new_n11897, new_n11898,
    new_n11899, new_n11900, new_n11901, new_n11902, new_n11903, new_n11904,
    new_n11905, new_n11906, new_n11907, new_n11908, new_n11909, new_n11910,
    new_n11911, new_n11912, new_n11913, new_n11914, new_n11915, new_n11916,
    new_n11917, new_n11918, new_n11919, new_n11920, new_n11921, new_n11922,
    new_n11923, new_n11924, new_n11925, new_n11926, new_n11927, new_n11928,
    new_n11929, new_n11930, new_n11931, new_n11932, new_n11933, new_n11934,
    new_n11935, new_n11936, new_n11937, new_n11938, new_n11939, new_n11940,
    new_n11941, new_n11942, new_n11943, new_n11944, new_n11945, new_n11946,
    new_n11947, new_n11948, new_n11949, new_n11950, new_n11951, new_n11952,
    new_n11953, new_n11954, new_n11955, new_n11956, new_n11957, new_n11958,
    new_n11959, new_n11960, new_n11961, new_n11962, new_n11963, new_n11964,
    new_n11965, new_n11966, new_n11967, new_n11968, new_n11969, new_n11970,
    new_n11971, new_n11972, new_n11973, new_n11974, new_n11975, new_n11976,
    new_n11977, new_n11978, new_n11979, new_n11980, new_n11981, new_n11982,
    new_n11983, new_n11984, new_n11985, new_n11986, new_n11987, new_n11988,
    new_n11989, new_n11990, new_n11991, new_n11992, new_n11993, new_n11994,
    new_n11995, new_n11996, new_n11997, new_n11998, new_n11999, new_n12000,
    new_n12001, new_n12002, new_n12003, new_n12004, new_n12005, new_n12006,
    new_n12007, new_n12008, new_n12009, new_n12010, new_n12011, new_n12012,
    new_n12013, new_n12014, new_n12015, new_n12016, new_n12017, new_n12018,
    new_n12019, new_n12020, new_n12021, new_n12022, new_n12023, new_n12024,
    new_n12025, new_n12026, new_n12027, new_n12028, new_n12029, new_n12030,
    new_n12031, new_n12032, new_n12033, new_n12034, new_n12035, new_n12036,
    new_n12037, new_n12038, new_n12039, new_n12040, new_n12041, new_n12042,
    new_n12043, new_n12044, new_n12045, new_n12046, new_n12047, new_n12048,
    new_n12049, new_n12050, new_n12051, new_n12052, new_n12053, new_n12054,
    new_n12055, new_n12056, new_n12057, new_n12058, new_n12059, new_n12060,
    new_n12061, new_n12062, new_n12063, new_n12064, new_n12065, new_n12066,
    new_n12067, new_n12068, new_n12069, new_n12070, new_n12071, new_n12072,
    new_n12073, new_n12074, new_n12075, new_n12076, new_n12077, new_n12078,
    new_n12079, new_n12080, new_n12081, new_n12082, new_n12083, new_n12084,
    new_n12085, new_n12086, new_n12087, new_n12088, new_n12089, new_n12090,
    new_n12091, new_n12092, new_n12093, new_n12094, new_n12095, new_n12096,
    new_n12097, new_n12098, new_n12099, new_n12100, new_n12101, new_n12102,
    new_n12103, new_n12104, new_n12105, new_n12106, new_n12107, new_n12108,
    new_n12109, new_n12110, new_n12111, new_n12112, new_n12113, new_n12114,
    new_n12115, new_n12116, new_n12117, new_n12118, new_n12119, new_n12120,
    new_n12121, new_n12122, new_n12123, new_n12124, new_n12125, new_n12126,
    new_n12127, new_n12128, new_n12129, new_n12130, new_n12131, new_n12132,
    new_n12133, new_n12134, new_n12135, new_n12136, new_n12137, new_n12138,
    new_n12139, new_n12140, new_n12141, new_n12142, new_n12143, new_n12144,
    new_n12145, new_n12146, new_n12147, new_n12148, new_n12149, new_n12150,
    new_n12151, new_n12152, new_n12153, new_n12154, new_n12155, new_n12156,
    new_n12157, new_n12158, new_n12159, new_n12160, new_n12161, new_n12162,
    new_n12163, new_n12164, new_n12165, new_n12166, new_n12167, new_n12168,
    new_n12169, new_n12170, new_n12171, new_n12172, new_n12173, new_n12174,
    new_n12175, new_n12176, new_n12177, new_n12178, new_n12179, new_n12180,
    new_n12181, new_n12182, new_n12183, new_n12184, new_n12185, new_n12186,
    new_n12187, new_n12188, new_n12189, new_n12190, new_n12191, new_n12192,
    new_n12193, new_n12194, new_n12195, new_n12196, new_n12197, new_n12198,
    new_n12199, new_n12200, new_n12201, new_n12202, new_n12203, new_n12204,
    new_n12205, new_n12206, new_n12207, new_n12208, new_n12209, new_n12210,
    new_n12211, new_n12212, new_n12213, new_n12214, new_n12215, new_n12216,
    new_n12217, new_n12218, new_n12219, new_n12220, new_n12221, new_n12222,
    new_n12223, new_n12224, new_n12225, new_n12226, new_n12227, new_n12228,
    new_n12229, new_n12230, new_n12231, new_n12232, new_n12233, new_n12234,
    new_n12235, new_n12236, new_n12237, new_n12238, new_n12239, new_n12240,
    new_n12241, new_n12242, new_n12243, new_n12244, new_n12245, new_n12246,
    new_n12247, new_n12248, new_n12249, new_n12250, new_n12251, new_n12252,
    new_n12253, new_n12254, new_n12255, new_n12256, new_n12257, new_n12258,
    new_n12259, new_n12260, new_n12261, new_n12262, new_n12263, new_n12264,
    new_n12265, new_n12266, new_n12267, new_n12268, new_n12269, new_n12270,
    new_n12271, new_n12272, new_n12273, new_n12274, new_n12275, new_n12276,
    new_n12277, new_n12278, new_n12279, new_n12280, new_n12281, new_n12282,
    new_n12283, new_n12284, new_n12285, new_n12286, new_n12287, new_n12288,
    new_n12289, new_n12290, new_n12291, new_n12292, new_n12293, new_n12294,
    new_n12295, new_n12296, new_n12297, new_n12298, new_n12299, new_n12300,
    new_n12301, new_n12302, new_n12303, new_n12304, new_n12305, new_n12306,
    new_n12307, new_n12308, new_n12309, new_n12310, new_n12311, new_n12312,
    new_n12313, new_n12314, new_n12315, new_n12316, new_n12317, new_n12318,
    new_n12319, new_n12320, new_n12321, new_n12322, new_n12323, new_n12324,
    new_n12325, new_n12326, new_n12327, new_n12328, new_n12329, new_n12330,
    new_n12331, new_n12332, new_n12333, new_n12334, new_n12335, new_n12336,
    new_n12337, new_n12338, new_n12339, new_n12340, new_n12341, new_n12342,
    new_n12343, new_n12344, new_n12345, new_n12346, new_n12347, new_n12348,
    new_n12349, new_n12350, new_n12351, new_n12352, new_n12353, new_n12354,
    new_n12355, new_n12356, new_n12357, new_n12358, new_n12359, new_n12360,
    new_n12361, new_n12362, new_n12363, new_n12364, new_n12365, new_n12366,
    new_n12367, new_n12368, new_n12369, new_n12370, new_n12371, new_n12372,
    new_n12373, new_n12374, new_n12375, new_n12376, new_n12377, new_n12378,
    new_n12379, new_n12380, new_n12381, new_n12382, new_n12383, new_n12384,
    new_n12385, new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391, new_n12392, new_n12393, new_n12394, new_n12395, new_n12396,
    new_n12397, new_n12398, new_n12399, new_n12400, new_n12401, new_n12402,
    new_n12403, new_n12404, new_n12405, new_n12406, new_n12407, new_n12408,
    new_n12409, new_n12410, new_n12411, new_n12412, new_n12413, new_n12414,
    new_n12415, new_n12416, new_n12417, new_n12418, new_n12419, new_n12420,
    new_n12421, new_n12422, new_n12423, new_n12424, new_n12425, new_n12426,
    new_n12427, new_n12428, new_n12429, new_n12430, new_n12431, new_n12432,
    new_n12433, new_n12434, new_n12435, new_n12436, new_n12437, new_n12438,
    new_n12439, new_n12440, new_n12441, new_n12442, new_n12443, new_n12444,
    new_n12445, new_n12446, new_n12447, new_n12448, new_n12449, new_n12450,
    new_n12451, new_n12452, new_n12453, new_n12454, new_n12455, new_n12456,
    new_n12457, new_n12458, new_n12459, new_n12460, new_n12461, new_n12462,
    new_n12463, new_n12464, new_n12465, new_n12466, new_n12467, new_n12468,
    new_n12469, new_n12470, new_n12471, new_n12472, new_n12473, new_n12474,
    new_n12475, new_n12476, new_n12477, new_n12478, new_n12479, new_n12480,
    new_n12481, new_n12482, new_n12483, new_n12484, new_n12485, new_n12486,
    new_n12487, new_n12488, new_n12489, new_n12490, new_n12491, new_n12492,
    new_n12493, new_n12494, new_n12495, new_n12496, new_n12497, new_n12498,
    new_n12499, new_n12500, new_n12501, new_n12502, new_n12503, new_n12504,
    new_n12505, new_n12506, new_n12507, new_n12508, new_n12509, new_n12510,
    new_n12511, new_n12512, new_n12513, new_n12514, new_n12515, new_n12516,
    new_n12517, new_n12518, new_n12519, new_n12520, new_n12521, new_n12522,
    new_n12523, new_n12524, new_n12525, new_n12526, new_n12527, new_n12528,
    new_n12529, new_n12530, new_n12531, new_n12532, new_n12533, new_n12534,
    new_n12535, new_n12536, new_n12537, new_n12538, new_n12539, new_n12540,
    new_n12541, new_n12542, new_n12543, new_n12544, new_n12545, new_n12546,
    new_n12547, new_n12548, new_n12549, new_n12550, new_n12551, new_n12552,
    new_n12553, new_n12554, new_n12555, new_n12556, new_n12557, new_n12558,
    new_n12559, new_n12560, new_n12561, new_n12562, new_n12563, new_n12564,
    new_n12565, new_n12566, new_n12567, new_n12568, new_n12569, new_n12570,
    new_n12571, new_n12572, new_n12573, new_n12574, new_n12575, new_n12576,
    new_n12577, new_n12578, new_n12579, new_n12580, new_n12581, new_n12582,
    new_n12583, new_n12584, new_n12585, new_n12586, new_n12587, new_n12588,
    new_n12589, new_n12590, new_n12591, new_n12592, new_n12593, new_n12594,
    new_n12595, new_n12596, new_n12597, new_n12598, new_n12599, new_n12600,
    new_n12601, new_n12602, new_n12603, new_n12604, new_n12605, new_n12606,
    new_n12607, new_n12608, new_n12609, new_n12610, new_n12611, new_n12612,
    new_n12613, new_n12614, new_n12615, new_n12616, new_n12617, new_n12618,
    new_n12619, new_n12620, new_n12621, new_n12622, new_n12623, new_n12624,
    new_n12625, new_n12626, new_n12627, new_n12628, new_n12629, new_n12630,
    new_n12631, new_n12632, new_n12633, new_n12634, new_n12635, new_n12636,
    new_n12637, new_n12638, new_n12639, new_n12640, new_n12641, new_n12642,
    new_n12643, new_n12644, new_n12645, new_n12646, new_n12647, new_n12648,
    new_n12649, new_n12650, new_n12651, new_n12652, new_n12653, new_n12654,
    new_n12655, new_n12656, new_n12657, new_n12658, new_n12659, new_n12660,
    new_n12661, new_n12662, new_n12663, new_n12664, new_n12665, new_n12666,
    new_n12667, new_n12668, new_n12669, new_n12670, new_n12671, new_n12672,
    new_n12673, new_n12674, new_n12675, new_n12676, new_n12677, new_n12678,
    new_n12679, new_n12680, new_n12681, new_n12682, new_n12683, new_n12684,
    new_n12685, new_n12686, new_n12687, new_n12688, new_n12689, new_n12690,
    new_n12691, new_n12692, new_n12693, new_n12694, new_n12695, new_n12696,
    new_n12697, new_n12698, new_n12699, new_n12700, new_n12701, new_n12702,
    new_n12703, new_n12704, new_n12705, new_n12706, new_n12707, new_n12708,
    new_n12709, new_n12710, new_n12711, new_n12712, new_n12713, new_n12714,
    new_n12715, new_n12716, new_n12717, new_n12718, new_n12719, new_n12720,
    new_n12721, new_n12722, new_n12723, new_n12724, new_n12725, new_n12726,
    new_n12727, new_n12728, new_n12729, new_n12730, new_n12731, new_n12732,
    new_n12733, new_n12734, new_n12735, new_n12736, new_n12737, new_n12738,
    new_n12739, new_n12740, new_n12741, new_n12742, new_n12743, new_n12744,
    new_n12745, new_n12746, new_n12747, new_n12748, new_n12749, new_n12750,
    new_n12751, new_n12752, new_n12753, new_n12754, new_n12755, new_n12756,
    new_n12757, new_n12758, new_n12759, new_n12760, new_n12761, new_n12762,
    new_n12763, new_n12764, new_n12765, new_n12766, new_n12767, new_n12768,
    new_n12769, new_n12770, new_n12771, new_n12772, new_n12773, new_n12774,
    new_n12775, new_n12776, new_n12777, new_n12778, new_n12779, new_n12780,
    new_n12781, new_n12782, new_n12783, new_n12784, new_n12785, new_n12786,
    new_n12787, new_n12788, new_n12789, new_n12790, new_n12791, new_n12792,
    new_n12793, new_n12794, new_n12795, new_n12796, new_n12797, new_n12798,
    new_n12799, new_n12800, new_n12801, new_n12802, new_n12803, new_n12804,
    new_n12805, new_n12806, new_n12807, new_n12808, new_n12809, new_n12810,
    new_n12811, new_n12812, new_n12813, new_n12814, new_n12815, new_n12816,
    new_n12817, new_n12818, new_n12819, new_n12820, new_n12821, new_n12822,
    new_n12823, new_n12824, new_n12825, new_n12826, new_n12827, new_n12828,
    new_n12829, new_n12830, new_n12831, new_n12832, new_n12833, new_n12834,
    new_n12835, new_n12836, new_n12837, new_n12838, new_n12839, new_n12840,
    new_n12841, new_n12842, new_n12843, new_n12844, new_n12845, new_n12846,
    new_n12847, new_n12848, new_n12849, new_n12850, new_n12851, new_n12852,
    new_n12853, new_n12854, new_n12855, new_n12856, new_n12857, new_n12858,
    new_n12859, new_n12860, new_n12861, new_n12862, new_n12863, new_n12864,
    new_n12865, new_n12866, new_n12867, new_n12868, new_n12869, new_n12870,
    new_n12871, new_n12872, new_n12873, new_n12874, new_n12875, new_n12876,
    new_n12877, new_n12878, new_n12879, new_n12880, new_n12881, new_n12882,
    new_n12883, new_n12884, new_n12885, new_n12886, new_n12887, new_n12888,
    new_n12889, new_n12890, new_n12891, new_n12892, new_n12893, new_n12894,
    new_n12895, new_n12896, new_n12897, new_n12898, new_n12899, new_n12900,
    new_n12901, new_n12902, new_n12903, new_n12904, new_n12905, new_n12906,
    new_n12907, new_n12908, new_n12909, new_n12910, new_n12911, new_n12912,
    new_n12913, new_n12914, new_n12915, new_n12916, new_n12917, new_n12918,
    new_n12919, new_n12920, new_n12921, new_n12922, new_n12923, new_n12924,
    new_n12925, new_n12926, new_n12927, new_n12928, new_n12929, new_n12930,
    new_n12931, new_n12932, new_n12933, new_n12934, new_n12935, new_n12936,
    new_n12937, new_n12938, new_n12939, new_n12940, new_n12941, new_n12942,
    new_n12943, new_n12944, new_n12945, new_n12946, new_n12947, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956, new_n12957, new_n12958, new_n12959, new_n12960,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972,
    new_n12973, new_n12974, new_n12975, new_n12976, new_n12977, new_n12978,
    new_n12979, new_n12980, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985, new_n12986, new_n12987, new_n12988, new_n12989, new_n12990,
    new_n12991, new_n12992, new_n12993, new_n12994, new_n12995, new_n12996,
    new_n12997, new_n12998, new_n12999, new_n13000, new_n13001, new_n13002,
    new_n13003, new_n13004, new_n13005, new_n13006, new_n13007, new_n13008,
    new_n13009, new_n13010, new_n13011, new_n13012, new_n13013, new_n13014,
    new_n13015, new_n13016, new_n13017, new_n13018, new_n13019, new_n13020,
    new_n13021, new_n13022, new_n13023, new_n13024, new_n13025, new_n13026,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043, new_n13044,
    new_n13045, new_n13046, new_n13047, new_n13048, new_n13049, new_n13050,
    new_n13051, new_n13052, new_n13053, new_n13054, new_n13055, new_n13056,
    new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062,
    new_n13063, new_n13064, new_n13065, new_n13066, new_n13067, new_n13068,
    new_n13069, new_n13070, new_n13071, new_n13072, new_n13073, new_n13074,
    new_n13075, new_n13076, new_n13077, new_n13078, new_n13079, new_n13080,
    new_n13081, new_n13082, new_n13083, new_n13084, new_n13085, new_n13086,
    new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092,
    new_n13093, new_n13094, new_n13095, new_n13096, new_n13097, new_n13098,
    new_n13099, new_n13100, new_n13101, new_n13102, new_n13103, new_n13104,
    new_n13105, new_n13106, new_n13107, new_n13108, new_n13109, new_n13110,
    new_n13111, new_n13112, new_n13113, new_n13114, new_n13115, new_n13116,
    new_n13117, new_n13118, new_n13119, new_n13120, new_n13121, new_n13122,
    new_n13123, new_n13124, new_n13125, new_n13126, new_n13127, new_n13128,
    new_n13129, new_n13130, new_n13131, new_n13132, new_n13133, new_n13134,
    new_n13135, new_n13136, new_n13137, new_n13138, new_n13139, new_n13140,
    new_n13141, new_n13142, new_n13143, new_n13144, new_n13145, new_n13146,
    new_n13147, new_n13148, new_n13149, new_n13150, new_n13151, new_n13152,
    new_n13153, new_n13154, new_n13155, new_n13156, new_n13157, new_n13158,
    new_n13159, new_n13160, new_n13161, new_n13162, new_n13163, new_n13164,
    new_n13165, new_n13166, new_n13167, new_n13168, new_n13169, new_n13170,
    new_n13171, new_n13172, new_n13173, new_n13174, new_n13175, new_n13176,
    new_n13177, new_n13178, new_n13179, new_n13180, new_n13181, new_n13182,
    new_n13183, new_n13184, new_n13185, new_n13186, new_n13187, new_n13188,
    new_n13189, new_n13190, new_n13191, new_n13192, new_n13193, new_n13194,
    new_n13195, new_n13196, new_n13197, new_n13198, new_n13199, new_n13200,
    new_n13201, new_n13202, new_n13203, new_n13204, new_n13205, new_n13206,
    new_n13207, new_n13208, new_n13209, new_n13210, new_n13211, new_n13212,
    new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218,
    new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224,
    new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230,
    new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236,
    new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13255, new_n13256, new_n13257, new_n13258, new_n13259, new_n13260,
    new_n13261, new_n13262, new_n13263, new_n13264, new_n13265, new_n13266,
    new_n13267, new_n13268, new_n13269, new_n13270, new_n13271, new_n13272,
    new_n13273, new_n13274, new_n13275, new_n13276, new_n13277, new_n13278,
    new_n13279, new_n13280, new_n13281, new_n13282, new_n13283, new_n13284,
    new_n13285, new_n13286, new_n13287, new_n13288, new_n13289, new_n13290,
    new_n13291, new_n13292, new_n13293, new_n13294, new_n13295, new_n13296,
    new_n13297, new_n13298, new_n13299, new_n13300, new_n13301, new_n13302,
    new_n13303, new_n13304, new_n13305, new_n13306, new_n13307, new_n13308,
    new_n13309, new_n13310, new_n13311, new_n13312, new_n13313, new_n13314,
    new_n13315, new_n13316, new_n13317, new_n13318, new_n13319, new_n13320,
    new_n13321, new_n13322, new_n13323, new_n13324, new_n13325, new_n13326,
    new_n13327, new_n13328, new_n13329, new_n13330, new_n13331, new_n13332,
    new_n13333, new_n13334, new_n13335, new_n13336, new_n13337, new_n13338,
    new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344,
    new_n13345, new_n13346, new_n13347, new_n13348, new_n13349, new_n13350,
    new_n13351, new_n13352, new_n13353, new_n13354, new_n13355, new_n13356,
    new_n13357, new_n13358, new_n13359, new_n13360, new_n13361, new_n13362,
    new_n13363, new_n13364, new_n13365, new_n13366, new_n13367, new_n13368,
    new_n13369, new_n13370, new_n13371, new_n13372, new_n13373, new_n13374,
    new_n13375, new_n13376, new_n13377, new_n13378, new_n13379, new_n13380,
    new_n13381, new_n13382, new_n13383, new_n13384, new_n13385, new_n13386,
    new_n13387, new_n13388, new_n13389, new_n13390, new_n13391, new_n13392,
    new_n13393, new_n13394, new_n13395, new_n13396, new_n13397, new_n13398,
    new_n13399, new_n13400, new_n13401, new_n13402, new_n13403, new_n13404,
    new_n13405, new_n13406, new_n13407, new_n13408, new_n13409, new_n13410,
    new_n13411, new_n13412, new_n13413, new_n13414, new_n13415, new_n13416,
    new_n13417, new_n13418, new_n13419, new_n13420, new_n13421, new_n13422,
    new_n13423, new_n13424, new_n13425, new_n13426, new_n13427, new_n13428,
    new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434,
    new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440,
    new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446,
    new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452,
    new_n13453, new_n13454, new_n13455, new_n13456, new_n13457, new_n13458,
    new_n13459, new_n13460, new_n13461, new_n13462, new_n13463, new_n13464,
    new_n13465, new_n13466, new_n13467, new_n13468, new_n13469, new_n13470,
    new_n13471, new_n13472, new_n13473, new_n13474, new_n13475, new_n13476,
    new_n13477, new_n13478, new_n13479, new_n13480, new_n13481, new_n13482,
    new_n13483, new_n13484, new_n13485, new_n13486, new_n13487, new_n13488,
    new_n13489, new_n13490, new_n13491, new_n13492, new_n13493, new_n13494,
    new_n13495, new_n13496, new_n13497, new_n13498, new_n13499, new_n13500,
    new_n13501, new_n13502, new_n13503, new_n13504, new_n13505, new_n13506,
    new_n13507, new_n13508, new_n13509, new_n13510, new_n13511, new_n13512,
    new_n13513, new_n13514, new_n13515, new_n13516, new_n13517, new_n13518,
    new_n13519, new_n13520, new_n13521, new_n13522, new_n13523, new_n13524,
    new_n13525, new_n13526, new_n13527, new_n13528, new_n13529, new_n13530,
    new_n13531, new_n13532, new_n13533, new_n13534, new_n13535, new_n13536,
    new_n13537, new_n13538, new_n13539, new_n13540, new_n13541, new_n13542,
    new_n13543, new_n13544, new_n13545, new_n13546, new_n13547, new_n13548,
    new_n13549, new_n13550, new_n13551, new_n13552, new_n13553, new_n13554,
    new_n13555, new_n13556, new_n13557, new_n13558, new_n13559, new_n13560,
    new_n13561, new_n13562, new_n13563, new_n13564, new_n13565, new_n13566,
    new_n13567, new_n13568, new_n13569, new_n13570, new_n13571, new_n13572,
    new_n13573, new_n13574, new_n13575, new_n13576, new_n13577, new_n13578,
    new_n13579, new_n13580, new_n13581, new_n13582, new_n13583, new_n13584,
    new_n13585, new_n13586, new_n13587, new_n13588, new_n13589, new_n13590,
    new_n13591, new_n13592, new_n13593, new_n13594, new_n13595, new_n13596,
    new_n13597, new_n13598, new_n13599, new_n13600, new_n13601, new_n13602,
    new_n13603, new_n13604, new_n13605, new_n13606, new_n13607, new_n13608,
    new_n13609, new_n13610, new_n13611, new_n13612, new_n13613, new_n13614,
    new_n13615, new_n13616, new_n13617, new_n13618, new_n13619, new_n13620,
    new_n13621, new_n13622, new_n13623, new_n13624, new_n13625, new_n13626,
    new_n13627, new_n13628, new_n13629, new_n13630, new_n13631, new_n13632,
    new_n13633, new_n13634, new_n13635, new_n13636, new_n13637, new_n13638,
    new_n13639, new_n13640, new_n13641, new_n13642, new_n13643, new_n13644,
    new_n13645, new_n13646, new_n13647, new_n13648, new_n13649, new_n13650,
    new_n13651, new_n13652, new_n13653, new_n13654, new_n13655, new_n13656,
    new_n13657, new_n13658, new_n13659, new_n13660, new_n13661, new_n13662,
    new_n13663, new_n13664, new_n13665, new_n13666, new_n13667, new_n13668,
    new_n13669, new_n13670, new_n13671, new_n13672, new_n13673, new_n13674,
    new_n13675, new_n13676, new_n13677, new_n13678, new_n13679, new_n13680,
    new_n13681, new_n13682, new_n13683, new_n13684, new_n13685, new_n13686,
    new_n13687, new_n13688, new_n13689, new_n13690, new_n13691, new_n13692,
    new_n13693, new_n13694, new_n13695, new_n13696, new_n13697, new_n13698,
    new_n13699, new_n13700, new_n13701, new_n13702, new_n13703, new_n13704,
    new_n13705, new_n13706, new_n13707, new_n13708, new_n13709, new_n13710,
    new_n13711, new_n13712, new_n13713, new_n13714, new_n13715, new_n13716,
    new_n13717, new_n13718, new_n13719, new_n13720, new_n13721, new_n13722,
    new_n13723, new_n13724, new_n13725, new_n13726, new_n13727, new_n13728,
    new_n13729, new_n13730, new_n13731, new_n13732, new_n13733, new_n13734,
    new_n13735, new_n13736, new_n13737, new_n13738, new_n13739, new_n13740,
    new_n13741, new_n13742, new_n13743, new_n13744, new_n13745, new_n13746,
    new_n13747, new_n13748, new_n13749, new_n13750, new_n13751, new_n13752,
    new_n13753, new_n13754, new_n13755, new_n13756, new_n13757, new_n13758,
    new_n13759, new_n13760, new_n13761, new_n13762, new_n13763, new_n13764,
    new_n13765, new_n13766, new_n13767, new_n13768, new_n13769, new_n13770,
    new_n13771, new_n13772, new_n13773, new_n13774, new_n13775, new_n13776,
    new_n13777, new_n13778, new_n13779, new_n13780, new_n13781, new_n13782,
    new_n13783, new_n13784, new_n13785, new_n13786, new_n13787, new_n13788,
    new_n13789, new_n13790, new_n13791, new_n13792, new_n13793, new_n13794,
    new_n13795, new_n13796, new_n13797, new_n13798, new_n13799, new_n13800,
    new_n13801, new_n13802, new_n13803, new_n13804, new_n13805, new_n13806,
    new_n13807, new_n13808, new_n13809, new_n13810, new_n13811, new_n13812,
    new_n13813, new_n13814, new_n13815, new_n13816, new_n13817, new_n13818,
    new_n13819, new_n13820, new_n13821, new_n13822, new_n13823, new_n13824,
    new_n13825, new_n13826, new_n13827, new_n13828, new_n13829, new_n13830,
    new_n13831, new_n13832, new_n13833, new_n13834, new_n13835, new_n13836,
    new_n13837, new_n13838, new_n13839, new_n13840, new_n13841, new_n13842,
    new_n13843, new_n13844, new_n13845, new_n13846, new_n13847, new_n13848,
    new_n13849, new_n13850, new_n13851, new_n13852, new_n13853, new_n13854,
    new_n13855, new_n13856, new_n13857, new_n13858, new_n13859, new_n13860,
    new_n13861, new_n13862, new_n13863, new_n13864, new_n13865, new_n13866,
    new_n13867, new_n13868, new_n13869, new_n13870, new_n13871, new_n13872,
    new_n13873, new_n13874, new_n13875, new_n13876, new_n13877, new_n13878,
    new_n13879, new_n13880, new_n13881, new_n13882, new_n13883, new_n13884,
    new_n13885, new_n13886, new_n13887, new_n13888, new_n13889, new_n13890,
    new_n13891, new_n13892, new_n13893, new_n13894, new_n13895, new_n13896,
    new_n13897, new_n13898, new_n13899, new_n13900, new_n13901, new_n13902,
    new_n13903, new_n13904, new_n13905, new_n13906, new_n13907, new_n13908,
    new_n13909, new_n13910, new_n13911, new_n13912, new_n13913, new_n13914,
    new_n13915, new_n13916, new_n13917, new_n13918, new_n13919, new_n13920,
    new_n13921, new_n13922, new_n13923, new_n13924, new_n13925, new_n13926,
    new_n13927, new_n13928, new_n13929, new_n13930, new_n13931, new_n13932,
    new_n13933, new_n13934, new_n13935, new_n13936, new_n13937, new_n13938,
    new_n13939, new_n13940, new_n13941, new_n13942, new_n13943, new_n13944,
    new_n13945, new_n13946, new_n13947, new_n13948, new_n13949, new_n13950,
    new_n13951, new_n13952, new_n13953, new_n13954, new_n13955, new_n13956,
    new_n13957, new_n13958, new_n13959, new_n13960, new_n13961, new_n13962,
    new_n13963, new_n13964, new_n13965, new_n13966, new_n13967, new_n13968,
    new_n13969, new_n13970, new_n13971, new_n13972, new_n13973, new_n13974,
    new_n13975, new_n13976, new_n13977, new_n13978, new_n13979, new_n13980,
    new_n13981, new_n13982, new_n13983, new_n13984, new_n13985, new_n13986,
    new_n13987, new_n13988, new_n13989, new_n13990, new_n13991, new_n13992,
    new_n13993, new_n13994, new_n13995, new_n13996, new_n13997, new_n13998,
    new_n13999, new_n14000, new_n14001, new_n14002, new_n14003, new_n14004,
    new_n14005, new_n14006, new_n14007, new_n14008, new_n14009, new_n14010,
    new_n14011, new_n14012, new_n14013, new_n14014, new_n14015, new_n14016,
    new_n14017, new_n14018, new_n14019, new_n14020, new_n14021, new_n14022,
    new_n14023, new_n14024, new_n14025, new_n14026, new_n14027, new_n14028,
    new_n14029, new_n14030, new_n14031, new_n14032, new_n14033, new_n14034,
    new_n14035, new_n14036, new_n14037, new_n14038, new_n14039, new_n14040,
    new_n14041, new_n14042, new_n14043, new_n14044, new_n14045, new_n14046,
    new_n14047, new_n14048, new_n14049, new_n14050, new_n14051, new_n14052,
    new_n14053, new_n14054, new_n14055, new_n14056, new_n14057, new_n14058,
    new_n14059, new_n14060, new_n14061, new_n14062, new_n14063, new_n14064,
    new_n14065, new_n14066, new_n14067, new_n14068, new_n14069, new_n14070,
    new_n14071, new_n14072, new_n14073, new_n14074, new_n14075, new_n14076,
    new_n14077, new_n14078, new_n14079, new_n14080, new_n14081, new_n14082,
    new_n14083, new_n14084, new_n14085, new_n14086, new_n14087, new_n14088,
    new_n14089, new_n14090, new_n14091, new_n14092, new_n14093, new_n14094,
    new_n14095, new_n14096, new_n14097, new_n14098, new_n14099, new_n14100,
    new_n14101, new_n14102, new_n14103, new_n14104, new_n14105, new_n14106,
    new_n14107, new_n14108, new_n14109, new_n14110, new_n14111, new_n14112,
    new_n14113, new_n14114, new_n14115, new_n14116, new_n14117, new_n14118,
    new_n14119, new_n14120, new_n14121, new_n14122, new_n14123, new_n14124,
    new_n14125, new_n14126, new_n14127, new_n14128, new_n14129, new_n14130,
    new_n14131, new_n14132, new_n14133, new_n14134, new_n14135, new_n14136,
    new_n14137, new_n14138, new_n14139, new_n14140, new_n14141, new_n14142,
    new_n14143, new_n14144, new_n14145, new_n14146, new_n14147, new_n14148,
    new_n14149, new_n14150, new_n14151, new_n14152, new_n14153, new_n14154,
    new_n14155, new_n14156, new_n14157, new_n14158, new_n14159, new_n14160,
    new_n14161, new_n14162, new_n14163, new_n14164, new_n14165, new_n14166,
    new_n14167, new_n14168, new_n14169, new_n14170, new_n14171, new_n14172,
    new_n14173, new_n14174, new_n14175, new_n14176, new_n14177, new_n14178,
    new_n14179, new_n14180, new_n14181, new_n14182, new_n14183, new_n14184,
    new_n14185, new_n14186, new_n14187, new_n14188, new_n14189, new_n14190,
    new_n14191, new_n14192, new_n14193, new_n14194, new_n14195, new_n14196,
    new_n14197, new_n14198, new_n14199, new_n14200, new_n14201, new_n14202,
    new_n14203, new_n14204, new_n14205, new_n14206, new_n14207, new_n14208,
    new_n14209, new_n14210, new_n14211, new_n14212, new_n14213, new_n14214,
    new_n14215, new_n14216, new_n14217, new_n14218, new_n14219, new_n14220,
    new_n14221, new_n14222, new_n14223, new_n14224, new_n14225, new_n14226,
    new_n14227, new_n14228, new_n14229, new_n14230, new_n14231, new_n14232,
    new_n14233, new_n14234, new_n14235, new_n14236, new_n14237, new_n14238,
    new_n14239, new_n14240, new_n14241, new_n14242, new_n14243, new_n14244,
    new_n14245, new_n14246, new_n14247, new_n14248, new_n14249, new_n14250,
    new_n14251, new_n14252, new_n14253, new_n14254, new_n14255, new_n14256,
    new_n14257, new_n14258, new_n14259, new_n14260, new_n14261, new_n14262,
    new_n14263, new_n14264, new_n14265, new_n14266, new_n14267, new_n14268,
    new_n14269, new_n14270, new_n14271, new_n14272, new_n14273, new_n14274,
    new_n14275, new_n14276, new_n14277, new_n14278, new_n14279, new_n14280,
    new_n14281, new_n14282, new_n14283, new_n14284, new_n14285, new_n14286,
    new_n14287, new_n14288, new_n14289, new_n14290, new_n14291, new_n14292,
    new_n14293, new_n14294, new_n14295, new_n14296, new_n14297, new_n14298,
    new_n14299, new_n14300, new_n14301, new_n14302, new_n14303, new_n14304,
    new_n14305, new_n14306, new_n14307, new_n14308, new_n14309, new_n14310,
    new_n14311, new_n14312, new_n14313, new_n14314, new_n14315, new_n14316,
    new_n14317, new_n14318, new_n14319, new_n14320, new_n14321, new_n14322,
    new_n14323, new_n14324, new_n14325, new_n14326, new_n14327, new_n14328,
    new_n14329, new_n14330, new_n14331, new_n14332, new_n14333, new_n14334,
    new_n14335, new_n14336, new_n14337, new_n14338, new_n14339, new_n14340,
    new_n14341, new_n14342, new_n14343, new_n14344, new_n14345, new_n14346,
    new_n14347, new_n14348, new_n14349, new_n14350, new_n14351, new_n14352,
    new_n14353, new_n14354, new_n14355, new_n14356, new_n14357, new_n14358,
    new_n14359, new_n14360, new_n14361, new_n14362, new_n14363, new_n14364,
    new_n14365, new_n14366, new_n14367, new_n14368, new_n14369, new_n14370,
    new_n14371, new_n14372, new_n14373, new_n14374, new_n14375, new_n14376,
    new_n14377, new_n14378, new_n14379, new_n14380, new_n14381, new_n14382,
    new_n14383, new_n14384, new_n14385, new_n14386, new_n14387, new_n14388,
    new_n14389, new_n14390, new_n14391, new_n14392, new_n14393, new_n14394,
    new_n14395, new_n14396, new_n14397, new_n14398, new_n14399, new_n14400,
    new_n14401, new_n14402, new_n14403, new_n14404, new_n14405, new_n14406,
    new_n14407, new_n14408, new_n14409, new_n14410, new_n14411, new_n14412,
    new_n14413, new_n14414, new_n14415, new_n14416, new_n14417, new_n14418,
    new_n14419, new_n14420, new_n14421, new_n14422, new_n14423, new_n14424,
    new_n14425, new_n14426, new_n14427, new_n14428, new_n14429, new_n14430,
    new_n14431, new_n14432, new_n14433, new_n14434, new_n14435, new_n14436,
    new_n14437, new_n14438, new_n14439, new_n14440, new_n14441, new_n14442,
    new_n14443, new_n14444, new_n14445, new_n14446, new_n14447, new_n14448,
    new_n14449, new_n14450, new_n14451, new_n14452, new_n14453, new_n14454,
    new_n14455, new_n14456, new_n14457, new_n14458, new_n14459, new_n14460,
    new_n14461, new_n14462, new_n14463, new_n14464, new_n14465, new_n14466,
    new_n14467, new_n14468, new_n14469, new_n14470, new_n14471, new_n14472,
    new_n14473, new_n14474, new_n14475, new_n14476, new_n14477, new_n14478,
    new_n14479, new_n14480, new_n14481, new_n14482, new_n14483, new_n14484,
    new_n14485, new_n14486, new_n14487, new_n14488, new_n14489, new_n14490,
    new_n14491, new_n14492, new_n14493, new_n14494, new_n14495, new_n14496,
    new_n14497, new_n14498, new_n14499, new_n14500, new_n14501, new_n14502,
    new_n14503, new_n14504, new_n14505, new_n14506, new_n14507, new_n14508,
    new_n14509, new_n14510, new_n14511, new_n14512, new_n14513, new_n14514,
    new_n14515, new_n14516, new_n14517, new_n14518, new_n14519, new_n14520,
    new_n14521, new_n14522, new_n14523, new_n14524, new_n14525, new_n14526,
    new_n14527, new_n14528, new_n14529, new_n14530, new_n14531, new_n14532,
    new_n14533, new_n14534, new_n14535, new_n14536, new_n14537, new_n14538,
    new_n14539, new_n14540, new_n14541, new_n14542, new_n14543, new_n14544,
    new_n14545, new_n14546, new_n14547, new_n14548, new_n14549, new_n14550,
    new_n14551, new_n14552, new_n14553, new_n14554, new_n14555, new_n14556,
    new_n14557, new_n14558, new_n14559, new_n14560, new_n14561, new_n14562,
    new_n14563, new_n14564, new_n14565, new_n14566, new_n14567, new_n14568,
    new_n14569, new_n14570, new_n14571, new_n14572, new_n14573, new_n14574,
    new_n14575, new_n14576, new_n14577, new_n14578, new_n14579, new_n14580,
    new_n14581, new_n14582, new_n14583, new_n14584, new_n14585, new_n14586,
    new_n14587, new_n14588, new_n14589, new_n14590, new_n14591, new_n14592,
    new_n14593, new_n14594, new_n14595, new_n14596, new_n14597, new_n14598,
    new_n14599, new_n14600, new_n14601, new_n14602, new_n14603, new_n14604,
    new_n14605, new_n14606, new_n14607, new_n14608, new_n14609, new_n14610,
    new_n14611, new_n14612, new_n14613, new_n14614, new_n14615, new_n14616,
    new_n14617, new_n14618, new_n14619, new_n14620, new_n14621, new_n14622,
    new_n14623, new_n14624, new_n14625, new_n14626, new_n14627, new_n14628,
    new_n14629, new_n14630, new_n14631, new_n14632, new_n14633, new_n14634,
    new_n14635, new_n14636, new_n14637, new_n14638, new_n14639, new_n14640,
    new_n14641, new_n14642, new_n14643, new_n14644, new_n14645, new_n14646,
    new_n14647, new_n14648, new_n14649, new_n14650, new_n14651, new_n14652,
    new_n14653, new_n14654, new_n14655, new_n14656, new_n14657, new_n14658,
    new_n14659, new_n14660, new_n14661, new_n14662, new_n14663, new_n14664,
    new_n14665, new_n14666, new_n14667, new_n14668, new_n14669, new_n14670,
    new_n14671, new_n14672, new_n14673, new_n14674, new_n14675, new_n14676,
    new_n14677, new_n14678, new_n14679, new_n14680, new_n14681, new_n14682,
    new_n14683, new_n14684, new_n14685, new_n14686, new_n14687, new_n14688,
    new_n14689, new_n14690, new_n14691, new_n14692, new_n14693, new_n14694,
    new_n14695, new_n14696, new_n14697, new_n14698, new_n14699, new_n14700,
    new_n14701, new_n14702, new_n14703, new_n14704, new_n14705, new_n14706,
    new_n14707, new_n14708, new_n14709, new_n14710, new_n14711, new_n14712,
    new_n14713, new_n14714, new_n14715, new_n14716, new_n14717, new_n14718,
    new_n14719, new_n14720, new_n14721, new_n14722, new_n14723, new_n14724,
    new_n14725, new_n14726, new_n14727, new_n14728, new_n14729, new_n14730,
    new_n14731, new_n14732, new_n14733, new_n14734, new_n14735, new_n14736,
    new_n14737, new_n14738, new_n14739, new_n14740, new_n14741, new_n14742,
    new_n14743, new_n14744, new_n14745, new_n14746, new_n14747, new_n14748,
    new_n14749, new_n14750, new_n14751, new_n14752, new_n14753, new_n14754,
    new_n14755, new_n14756, new_n14757, new_n14758, new_n14759, new_n14760,
    new_n14761, new_n14762, new_n14763, new_n14764, new_n14765, new_n14766,
    new_n14767, new_n14768, new_n14769, new_n14770, new_n14771, new_n14772,
    new_n14773, new_n14774, new_n14775, new_n14776, new_n14777, new_n14778,
    new_n14779, new_n14780, new_n14781, new_n14782, new_n14783, new_n14784,
    new_n14785, new_n14786, new_n14787, new_n14788, new_n14789, new_n14790,
    new_n14791, new_n14792, new_n14793, new_n14794, new_n14795, new_n14796,
    new_n14797, new_n14798, new_n14799, new_n14800, new_n14801, new_n14802,
    new_n14803, new_n14804, new_n14805, new_n14806, new_n14807, new_n14808,
    new_n14809, new_n14810, new_n14811, new_n14812, new_n14813, new_n14814,
    new_n14815, new_n14816, new_n14817, new_n14818, new_n14819, new_n14820,
    new_n14821, new_n14822, new_n14823, new_n14824, new_n14825, new_n14826,
    new_n14827, new_n14828, new_n14829, new_n14830, new_n14831, new_n14832,
    new_n14833, new_n14834, new_n14835, new_n14836, new_n14837, new_n14838,
    new_n14839, new_n14840, new_n14841, new_n14842, new_n14843, new_n14844,
    new_n14845, new_n14846, new_n14847, new_n14848, new_n14849, new_n14850,
    new_n14851, new_n14852, new_n14853, new_n14854, new_n14855, new_n14856,
    new_n14857, new_n14858, new_n14859, new_n14860, new_n14861, new_n14862,
    new_n14863, new_n14864, new_n14865, new_n14866, new_n14867, new_n14868,
    new_n14869, new_n14870, new_n14871, new_n14872, new_n14873, new_n14874,
    new_n14875, new_n14876, new_n14877, new_n14878, new_n14879, new_n14880,
    new_n14881, new_n14882, new_n14883, new_n14884, new_n14885, new_n14886,
    new_n14887, new_n14888, new_n14889, new_n14890, new_n14891, new_n14892,
    new_n14893, new_n14894, new_n14895, new_n14896, new_n14897, new_n14898,
    new_n14899, new_n14900, new_n14901, new_n14902, new_n14903, new_n14904,
    new_n14905, new_n14906, new_n14907, new_n14908, new_n14909, new_n14910,
    new_n14911, new_n14912, new_n14913, new_n14914, new_n14915, new_n14916,
    new_n14917, new_n14918, new_n14919, new_n14920, new_n14921, new_n14922,
    new_n14923, new_n14924, new_n14925, new_n14926, new_n14927, new_n14928,
    new_n14929, new_n14930, new_n14931, new_n14932, new_n14933, new_n14934,
    new_n14935, new_n14936, new_n14937, new_n14938, new_n14939, new_n14940,
    new_n14941, new_n14942, new_n14943, new_n14944, new_n14945, new_n14946,
    new_n14947, new_n14948, new_n14949, new_n14950, new_n14951, new_n14952,
    new_n14953, new_n14954, new_n14955, new_n14956, new_n14957, new_n14958,
    new_n14959, new_n14960, new_n14961, new_n14962, new_n14963, new_n14964,
    new_n14965, new_n14966, new_n14967, new_n14968, new_n14969, new_n14970,
    new_n14971, new_n14972, new_n14973, new_n14974, new_n14975, new_n14976,
    new_n14977, new_n14978, new_n14979, new_n14980, new_n14981, new_n14982,
    new_n14983, new_n14984, new_n14985, new_n14986, new_n14987, new_n14988,
    new_n14989, new_n14990, new_n14991, new_n14992, new_n14993, new_n14994,
    new_n14995, new_n14996, new_n14997, new_n14998, new_n14999, new_n15000,
    new_n15001, new_n15002, new_n15003, new_n15004, new_n15005, new_n15006,
    new_n15007, new_n15008, new_n15009, new_n15010, new_n15011, new_n15012,
    new_n15013, new_n15014, new_n15015, new_n15016, new_n15017, new_n15018,
    new_n15019, new_n15020, new_n15021, new_n15022, new_n15023, new_n15024,
    new_n15025, new_n15026, new_n15027, new_n15028, new_n15029, new_n15030,
    new_n15031, new_n15032, new_n15033, new_n15034, new_n15035, new_n15036,
    new_n15037, new_n15038, new_n15039, new_n15040, new_n15041, new_n15042,
    new_n15043, new_n15044, new_n15045, new_n15046, new_n15047, new_n15048,
    new_n15049, new_n15050, new_n15051, new_n15052, new_n15053, new_n15054,
    new_n15055, new_n15056, new_n15057, new_n15058, new_n15059, new_n15060,
    new_n15061, new_n15062, new_n15063, new_n15064, new_n15065, new_n15066,
    new_n15067, new_n15068, new_n15069, new_n15070, new_n15071, new_n15072,
    new_n15073, new_n15074, new_n15075, new_n15076, new_n15077, new_n15078,
    new_n15079, new_n15080, new_n15081, new_n15082, new_n15083, new_n15084,
    new_n15085, new_n15086, new_n15087, new_n15088, new_n15089, new_n15090,
    new_n15091, new_n15092, new_n15093, new_n15094, new_n15095, new_n15096,
    new_n15097, new_n15098, new_n15099, new_n15100, new_n15101, new_n15102,
    new_n15103, new_n15104, new_n15105, new_n15106, new_n15107, new_n15108,
    new_n15109, new_n15110, new_n15111, new_n15112, new_n15113, new_n15114,
    new_n15115, new_n15116, new_n15117, new_n15118, new_n15119, new_n15120,
    new_n15121, new_n15122, new_n15123, new_n15124, new_n15125, new_n15126,
    new_n15127, new_n15128, new_n15129, new_n15130, new_n15131, new_n15132,
    new_n15133, new_n15134, new_n15135, new_n15136, new_n15137, new_n15138,
    new_n15139, new_n15140, new_n15141, new_n15142, new_n15143, new_n15144,
    new_n15145, new_n15146, new_n15147, new_n15148, new_n15149, new_n15150,
    new_n15151, new_n15152, new_n15153, new_n15154, new_n15155, new_n15156,
    new_n15157, new_n15158, new_n15159, new_n15160, new_n15161, new_n15162,
    new_n15163, new_n15164, new_n15165, new_n15166, new_n15167, new_n15168,
    new_n15169, new_n15170, new_n15171, new_n15172, new_n15173, new_n15174,
    new_n15175, new_n15176, new_n15177, new_n15178, new_n15179, new_n15180,
    new_n15181, new_n15182, new_n15183, new_n15184, new_n15185, new_n15186,
    new_n15187, new_n15188, new_n15189, new_n15190, new_n15191, new_n15192,
    new_n15193, new_n15194, new_n15195, new_n15196, new_n15197, new_n15198,
    new_n15199, new_n15200, new_n15201, new_n15202, new_n15203, new_n15204,
    new_n15205, new_n15206, new_n15207, new_n15208, new_n15209, new_n15210,
    new_n15211, new_n15212, new_n15213, new_n15214, new_n15215, new_n15216,
    new_n15217, new_n15218, new_n15219, new_n15220, new_n15221, new_n15222,
    new_n15223, new_n15224, new_n15225, new_n15226, new_n15227, new_n15228,
    new_n15229, new_n15230, new_n15231, new_n15232, new_n15233, new_n15234,
    new_n15235, new_n15236, new_n15237, new_n15238, new_n15239, new_n15240,
    new_n15241, new_n15242, new_n15243, new_n15244, new_n15245, new_n15246,
    new_n15247, new_n15248, new_n15249, new_n15250, new_n15251, new_n15252,
    new_n15253, new_n15254, new_n15255, new_n15256, new_n15257, new_n15258,
    new_n15259, new_n15260, new_n15261, new_n15262, new_n15263, new_n15264,
    new_n15265, new_n15266, new_n15267, new_n15268, new_n15269, new_n15270,
    new_n15271, new_n15272, new_n15273, new_n15274, new_n15275, new_n15276,
    new_n15277, new_n15278, new_n15279, new_n15280, new_n15281, new_n15282,
    new_n15283, new_n15284, new_n15285, new_n15286, new_n15287, new_n15288,
    new_n15289, new_n15290, new_n15291, new_n15292, new_n15293, new_n15294,
    new_n15295, new_n15296, new_n15297, new_n15298, new_n15299, new_n15300,
    new_n15301, new_n15302, new_n15303, new_n15304, new_n15305, new_n15306,
    new_n15307, new_n15308, new_n15309, new_n15310, new_n15311, new_n15312,
    new_n15313, new_n15314, new_n15315, new_n15316, new_n15317, new_n15318,
    new_n15319, new_n15320, new_n15321, new_n15322, new_n15323, new_n15324,
    new_n15325, new_n15326, new_n15327, new_n15328, new_n15329, new_n15330,
    new_n15331, new_n15332, new_n15333, new_n15334, new_n15335, new_n15336,
    new_n15337, new_n15338, new_n15339, new_n15340, new_n15341, new_n15342,
    new_n15343, new_n15344, new_n15345, new_n15346, new_n15347, new_n15348,
    new_n15349, new_n15350, new_n15351, new_n15352, new_n15353, new_n15354,
    new_n15355, new_n15356, new_n15357, new_n15358, new_n15359, new_n15360,
    new_n15361, new_n15362, new_n15363, new_n15364, new_n15365, new_n15366,
    new_n15367, new_n15368, new_n15369, new_n15370, new_n15371, new_n15372,
    new_n15373, new_n15374, new_n15375, new_n15376, new_n15377, new_n15378,
    new_n15379, new_n15380, new_n15381, new_n15382, new_n15383, new_n15384,
    new_n15385, new_n15386, new_n15387, new_n15388, new_n15389, new_n15390,
    new_n15391, new_n15392, new_n15393, new_n15394, new_n15395, new_n15396,
    new_n15397, new_n15398, new_n15399, new_n15400, new_n15401, new_n15402,
    new_n15403, new_n15404, new_n15405, new_n15406, new_n15407, new_n15408,
    new_n15409, new_n15410, new_n15411, new_n15412, new_n15413, new_n15414,
    new_n15415, new_n15416, new_n15417, new_n15418, new_n15419, new_n15420,
    new_n15421, new_n15422, new_n15423, new_n15424, new_n15425, new_n15426,
    new_n15427, new_n15428, new_n15429, new_n15430, new_n15431, new_n15432,
    new_n15433, new_n15434, new_n15435, new_n15436, new_n15437, new_n15438,
    new_n15439, new_n15440, new_n15441, new_n15442, new_n15443, new_n15444,
    new_n15445, new_n15446, new_n15447, new_n15448, new_n15449, new_n15450,
    new_n15451, new_n15452, new_n15453, new_n15454, new_n15455, new_n15456,
    new_n15457, new_n15458, new_n15459, new_n15460, new_n15461, new_n15462,
    new_n15463, new_n15464, new_n15465, new_n15466, new_n15467, new_n15468,
    new_n15469, new_n15470, new_n15471, new_n15472, new_n15473, new_n15474,
    new_n15475, new_n15476, new_n15477, new_n15478, new_n15479, new_n15480,
    new_n15481, new_n15482, new_n15483, new_n15484, new_n15485, new_n15486,
    new_n15487, new_n15488, new_n15489, new_n15490, new_n15491, new_n15492,
    new_n15493, new_n15494, new_n15495, new_n15496, new_n15497, new_n15498,
    new_n15499, new_n15500, new_n15501, new_n15502, new_n15503, new_n15504,
    new_n15505, new_n15506, new_n15507, new_n15508, new_n15509, new_n15510,
    new_n15511, new_n15512, new_n15513, new_n15514, new_n15515, new_n15516,
    new_n15517, new_n15518, new_n15519, new_n15520, new_n15521, new_n15522,
    new_n15523, new_n15524, new_n15525, new_n15526, new_n15527, new_n15528,
    new_n15529, new_n15530, new_n15531, new_n15532, new_n15533, new_n15534,
    new_n15535, new_n15536, new_n15537, new_n15538, new_n15539, new_n15540,
    new_n15541, new_n15542, new_n15543, new_n15544, new_n15545, new_n15546,
    new_n15547, new_n15548, new_n15549, new_n15550, new_n15551, new_n15552,
    new_n15553, new_n15554, new_n15555, new_n15556, new_n15557, new_n15558,
    new_n15559, new_n15560, new_n15561, new_n15562, new_n15563, new_n15564,
    new_n15565, new_n15566, new_n15567, new_n15568, new_n15569, new_n15570,
    new_n15571, new_n15572, new_n15573, new_n15574, new_n15575, new_n15576,
    new_n15577, new_n15578, new_n15579, new_n15580, new_n15581, new_n15582,
    new_n15583, new_n15584, new_n15585, new_n15586, new_n15587, new_n15588,
    new_n15589, new_n15590, new_n15591, new_n15592, new_n15593, new_n15594,
    new_n15595, new_n15596, new_n15597, new_n15598, new_n15599, new_n15600,
    new_n15601, new_n15602, new_n15603, new_n15604, new_n15605, new_n15606,
    new_n15607, new_n15608, new_n15609, new_n15610, new_n15611, new_n15612,
    new_n15613, new_n15614, new_n15615, new_n15616, new_n15617, new_n15618,
    new_n15619, new_n15620, new_n15621, new_n15622, new_n15623, new_n15624,
    new_n15625, new_n15626, new_n15627, new_n15628, new_n15629, new_n15630,
    new_n15631, new_n15632, new_n15633, new_n15634, new_n15635, new_n15636,
    new_n15637, new_n15638, new_n15639, new_n15640, new_n15641, new_n15642,
    new_n15643, new_n15644, new_n15645, new_n15646, new_n15647, new_n15648,
    new_n15649, new_n15650, new_n15651, new_n15652, new_n15653, new_n15654,
    new_n15655, new_n15656, new_n15657, new_n15658, new_n15659, new_n15660,
    new_n15661, new_n15662, new_n15663, new_n15664, new_n15665, new_n15666,
    new_n15667, new_n15668, new_n15669, new_n15670, new_n15671, new_n15672,
    new_n15673, new_n15674, new_n15675, new_n15676, new_n15677, new_n15678,
    new_n15679, new_n15680, new_n15681, new_n15682, new_n15683, new_n15684,
    new_n15685, new_n15686, new_n15687, new_n15688, new_n15689, new_n15690,
    new_n15691, new_n15692, new_n15693, new_n15694, new_n15695, new_n15696,
    new_n15697, new_n15698, new_n15699, new_n15700, new_n15701, new_n15702,
    new_n15703, new_n15704, new_n15705, new_n15706, new_n15707, new_n15708,
    new_n15709, new_n15710, new_n15711, new_n15712, new_n15713, new_n15714,
    new_n15715, new_n15716, new_n15717, new_n15718, new_n15719, new_n15720,
    new_n15721, new_n15722, new_n15723, new_n15724, new_n15725, new_n15726,
    new_n15727, new_n15728, new_n15729, new_n15730, new_n15731, new_n15732,
    new_n15733, new_n15734, new_n15735, new_n15736, new_n15737, new_n15738,
    new_n15739, new_n15740, new_n15741, new_n15742, new_n15743, new_n15744,
    new_n15745, new_n15746, new_n15747, new_n15748, new_n15749, new_n15750,
    new_n15751, new_n15752, new_n15753, new_n15754, new_n15755, new_n15756,
    new_n15757, new_n15758, new_n15759, new_n15760, new_n15761, new_n15762,
    new_n15763, new_n15764, new_n15765, new_n15766, new_n15767, new_n15768,
    new_n15769, new_n15770, new_n15771, new_n15772, new_n15773, new_n15774,
    new_n15775, new_n15776, new_n15777, new_n15778, new_n15779, new_n15780,
    new_n15781, new_n15782, new_n15783, new_n15784, new_n15785, new_n15786,
    new_n15787, new_n15788, new_n15789, new_n15790, new_n15791, new_n15792,
    new_n15793, new_n15794, new_n15795, new_n15796, new_n15797, new_n15798,
    new_n15799, new_n15800, new_n15801, new_n15802, new_n15803, new_n15804,
    new_n15805, new_n15806, new_n15807, new_n15808, new_n15809, new_n15810,
    new_n15811, new_n15812, new_n15813, new_n15814, new_n15815, new_n15816,
    new_n15817, new_n15818, new_n15819, new_n15820, new_n15821, new_n15822,
    new_n15823, new_n15824, new_n15825, new_n15826, new_n15827, new_n15828,
    new_n15829, new_n15830, new_n15831, new_n15832, new_n15833, new_n15834,
    new_n15835, new_n15836, new_n15837, new_n15838, new_n15839, new_n15840,
    new_n15841, new_n15842, new_n15843, new_n15844, new_n15845, new_n15846,
    new_n15847, new_n15848, new_n15849, new_n15850, new_n15851, new_n15852,
    new_n15853, new_n15854, new_n15855, new_n15856, new_n15857, new_n15858,
    new_n15859, new_n15860, new_n15861, new_n15862, new_n15863, new_n15864,
    new_n15865, new_n15866, new_n15867, new_n15868, new_n15869, new_n15870,
    new_n15871, new_n15872, new_n15873, new_n15874, new_n15875, new_n15876,
    new_n15877, new_n15878, new_n15879, new_n15880, new_n15881, new_n15882,
    new_n15883, new_n15884, new_n15885, new_n15886, new_n15887, new_n15888,
    new_n15889, new_n15890, new_n15891, new_n15892, new_n15893, new_n15894,
    new_n15895, new_n15896, new_n15897, new_n15898, new_n15899, new_n15900,
    new_n15901, new_n15902, new_n15903, new_n15904, new_n15905, new_n15906,
    new_n15907, new_n15908, new_n15909, new_n15910, new_n15911, new_n15912,
    new_n15913, new_n15914, new_n15915, new_n15916, new_n15917, new_n15918,
    new_n15919, new_n15920, new_n15921, new_n15922, new_n15923, new_n15924,
    new_n15925, new_n15926, new_n15927, new_n15928, new_n15929, new_n15930,
    new_n15931, new_n15932, new_n15933, new_n15934, new_n15935, new_n15936,
    new_n15937, new_n15938, new_n15939, new_n15940, new_n15941, new_n15942,
    new_n15943, new_n15944, new_n15945, new_n15946, new_n15947, new_n15948,
    new_n15949, new_n15950, new_n15951, new_n15952, new_n15953, new_n15954,
    new_n15955, new_n15956, new_n15957, new_n15958, new_n15959, new_n15960,
    new_n15961, new_n15962, new_n15963, new_n15964, new_n15965, new_n15966,
    new_n15967, new_n15968, new_n15969, new_n15970, new_n15971, new_n15972,
    new_n15973, new_n15974, new_n15975, new_n15976, new_n15977, new_n15978,
    new_n15979, new_n15980, new_n15981, new_n15982, new_n15983, new_n15984,
    new_n15985, new_n15986, new_n15987, new_n15988, new_n15989, new_n15990,
    new_n15991, new_n15992, new_n15993, new_n15994, new_n15995, new_n15996,
    new_n15997, new_n15998, new_n15999, new_n16000, new_n16001, new_n16002,
    new_n16003, new_n16004, new_n16005, new_n16006, new_n16007, new_n16008,
    new_n16009, new_n16010, new_n16011, new_n16012, new_n16013, new_n16014,
    new_n16015, new_n16016, new_n16017, new_n16018, new_n16019, new_n16020,
    new_n16021, new_n16022, new_n16023, new_n16024, new_n16025, new_n16026,
    new_n16027, new_n16028, new_n16029, new_n16030, new_n16031, new_n16032,
    new_n16033, new_n16034, new_n16035, new_n16036, new_n16037, new_n16038,
    new_n16039, new_n16040, new_n16041, new_n16042, new_n16043, new_n16044,
    new_n16045, new_n16046, new_n16047, new_n16048, new_n16049, new_n16050,
    new_n16051, new_n16052, new_n16053, new_n16054, new_n16055, new_n16056,
    new_n16057, new_n16058, new_n16059, new_n16060, new_n16061, new_n16062,
    new_n16063, new_n16064, new_n16065, new_n16066, new_n16067, new_n16068,
    new_n16069, new_n16070, new_n16071, new_n16072, new_n16073, new_n16074,
    new_n16075, new_n16076, new_n16077, new_n16078, new_n16079, new_n16080,
    new_n16081, new_n16082, new_n16083, new_n16084, new_n16085, new_n16086,
    new_n16087, new_n16088, new_n16089, new_n16090, new_n16091, new_n16092,
    new_n16093, new_n16094, new_n16095, new_n16096, new_n16097, new_n16098,
    new_n16099, new_n16100, new_n16101, new_n16102, new_n16103, new_n16104,
    new_n16105, new_n16106, new_n16107, new_n16108, new_n16109, new_n16110,
    new_n16111, new_n16112, new_n16113, new_n16114, new_n16115, new_n16116,
    new_n16117, new_n16118, new_n16119, new_n16120, new_n16121, new_n16122,
    new_n16123, new_n16124, new_n16125, new_n16126, new_n16127, new_n16128,
    new_n16129, new_n16130, new_n16131, new_n16132, new_n16133, new_n16134,
    new_n16135, new_n16136, new_n16137, new_n16138, new_n16139, new_n16140,
    new_n16141, new_n16142, new_n16143, new_n16144, new_n16145, new_n16146,
    new_n16147, new_n16148, new_n16149, new_n16150, new_n16151, new_n16152,
    new_n16153, new_n16154, new_n16155, new_n16156, new_n16157, new_n16158,
    new_n16159, new_n16160, new_n16161, new_n16162, new_n16163, new_n16164,
    new_n16165, new_n16166, new_n16167, new_n16168, new_n16169, new_n16170,
    new_n16171, new_n16172, new_n16173, new_n16174, new_n16175, new_n16176,
    new_n16177, new_n16178, new_n16179, new_n16180, new_n16181, new_n16182,
    new_n16183, new_n16184, new_n16185, new_n16186, new_n16187, new_n16188,
    new_n16189, new_n16190, new_n16191, new_n16192, new_n16193, new_n16194,
    new_n16195, new_n16196, new_n16197, new_n16198, new_n16199, new_n16200,
    new_n16201, new_n16202, new_n16203, new_n16204, new_n16205, new_n16206,
    new_n16207, new_n16208, new_n16209, new_n16210, new_n16211, new_n16212,
    new_n16213, new_n16214, new_n16215, new_n16216, new_n16217, new_n16218,
    new_n16219, new_n16220, new_n16221, new_n16222, new_n16223, new_n16224,
    new_n16225, new_n16226, new_n16227, new_n16228, new_n16229, new_n16230,
    new_n16231, new_n16232, new_n16233, new_n16234, new_n16235, new_n16236,
    new_n16237, new_n16238, new_n16239, new_n16240, new_n16241, new_n16242,
    new_n16243, new_n16244, new_n16245, new_n16246, new_n16247, new_n16248,
    new_n16249, new_n16250, new_n16251, new_n16252, new_n16253, new_n16254,
    new_n16255, new_n16256, new_n16257, new_n16258, new_n16259, new_n16260,
    new_n16261, new_n16262, new_n16263, new_n16264, new_n16265, new_n16266,
    new_n16267, new_n16268, new_n16269, new_n16270, new_n16271, new_n16272,
    new_n16273, new_n16274, new_n16275, new_n16276, new_n16277, new_n16278,
    new_n16279, new_n16280, new_n16281, new_n16282, new_n16283, new_n16284,
    new_n16285, new_n16286, new_n16287, new_n16288, new_n16289, new_n16290,
    new_n16291, new_n16292, new_n16293, new_n16294, new_n16295, new_n16296,
    new_n16297, new_n16298, new_n16299, new_n16300, new_n16301, new_n16302,
    new_n16303, new_n16304, new_n16305, new_n16306, new_n16307, new_n16308,
    new_n16309, new_n16310, new_n16311, new_n16312, new_n16313, new_n16314,
    new_n16315, new_n16316, new_n16317, new_n16318, new_n16319, new_n16320,
    new_n16321, new_n16322, new_n16323, new_n16324, new_n16325, new_n16326,
    new_n16327, new_n16328, new_n16329, new_n16330, new_n16331, new_n16332,
    new_n16333, new_n16334, new_n16335, new_n16336, new_n16337, new_n16338,
    new_n16339, new_n16340, new_n16341, new_n16342, new_n16343, new_n16344,
    new_n16345, new_n16346, new_n16347, new_n16348, new_n16349, new_n16350,
    new_n16351, new_n16352, new_n16353, new_n16354, new_n16355, new_n16356,
    new_n16357, new_n16358, new_n16359, new_n16360, new_n16361, new_n16362,
    new_n16363, new_n16364, new_n16365, new_n16366, new_n16367, new_n16368,
    new_n16369, new_n16370, new_n16371, new_n16372, new_n16373, new_n16374,
    new_n16375, new_n16376, new_n16377, new_n16378, new_n16379, new_n16380,
    new_n16381, new_n16382, new_n16383, new_n16384, new_n16385, new_n16386,
    new_n16387, new_n16388, new_n16389, new_n16390, new_n16391, new_n16392,
    new_n16393, new_n16394, new_n16395, new_n16396, new_n16397, new_n16398,
    new_n16399, new_n16400, new_n16401, new_n16402, new_n16403, new_n16404,
    new_n16405, new_n16406, new_n16407, new_n16408, new_n16409, new_n16410,
    new_n16411, new_n16412, new_n16413, new_n16414, new_n16415, new_n16416,
    new_n16417, new_n16418, new_n16419, new_n16420, new_n16421, new_n16422,
    new_n16423, new_n16424, new_n16425, new_n16426, new_n16427, new_n16428,
    new_n16429, new_n16430, new_n16431, new_n16432, new_n16433, new_n16434,
    new_n16435, new_n16436, new_n16437, new_n16438, new_n16439, new_n16440,
    new_n16441, new_n16442, new_n16443, new_n16444, new_n16445, new_n16446,
    new_n16447, new_n16448, new_n16449, new_n16450, new_n16451, new_n16452,
    new_n16453, new_n16454, new_n16455, new_n16456, new_n16457, new_n16458,
    new_n16459, new_n16460, new_n16461, new_n16462, new_n16463, new_n16464,
    new_n16465, new_n16466, new_n16467, new_n16468, new_n16469, new_n16470,
    new_n16471, new_n16472, new_n16473, new_n16474, new_n16475, new_n16476,
    new_n16477, new_n16478, new_n16479, new_n16480, new_n16481, new_n16482,
    new_n16483, new_n16484, new_n16485, new_n16486, new_n16487, new_n16488,
    new_n16489, new_n16490, new_n16491, new_n16492, new_n16493, new_n16494,
    new_n16495, new_n16496, new_n16497, new_n16498, new_n16499, new_n16500,
    new_n16501, new_n16502, new_n16503, new_n16504, new_n16505, new_n16506,
    new_n16507, new_n16508, new_n16509, new_n16510, new_n16511, new_n16512,
    new_n16513, new_n16514, new_n16515, new_n16516, new_n16517, new_n16518,
    new_n16519, new_n16520, new_n16521, new_n16522, new_n16523, new_n16524,
    new_n16525, new_n16526, new_n16527, new_n16528, new_n16529, new_n16530,
    new_n16531, new_n16532, new_n16533, new_n16534, new_n16535, new_n16536,
    new_n16537, new_n16538, new_n16539, new_n16540, new_n16541, new_n16542,
    new_n16543, new_n16544, new_n16545, new_n16546, new_n16547, new_n16548,
    new_n16549, new_n16550, new_n16551, new_n16552, new_n16553, new_n16554,
    new_n16555, new_n16556, new_n16557, new_n16558, new_n16559, new_n16560,
    new_n16561, new_n16562, new_n16563, new_n16564, new_n16565, new_n16566,
    new_n16567, new_n16568, new_n16569, new_n16570, new_n16571, new_n16572,
    new_n16573, new_n16574, new_n16575, new_n16576, new_n16577, new_n16578,
    new_n16579, new_n16580, new_n16581, new_n16582, new_n16583, new_n16584,
    new_n16585, new_n16586, new_n16587, new_n16588, new_n16589, new_n16590,
    new_n16591, new_n16592, new_n16593, new_n16594, new_n16595, new_n16596,
    new_n16597, new_n16598, new_n16599, new_n16600, new_n16601, new_n16602,
    new_n16603, new_n16604, new_n16605, new_n16606, new_n16607, new_n16608,
    new_n16609, new_n16610, new_n16611, new_n16612, new_n16613, new_n16614,
    new_n16615, new_n16616, new_n16617, new_n16618, new_n16619, new_n16620,
    new_n16621, new_n16622, new_n16623, new_n16624, new_n16625, new_n16626,
    new_n16627, new_n16628, new_n16629, new_n16630, new_n16631, new_n16632,
    new_n16633, new_n16634, new_n16635, new_n16636, new_n16637, new_n16638,
    new_n16639, new_n16640, new_n16641, new_n16642, new_n16643, new_n16644,
    new_n16645, new_n16646, new_n16647, new_n16648, new_n16649, new_n16650,
    new_n16651, new_n16652, new_n16653, new_n16654, new_n16655, new_n16656,
    new_n16657, new_n16658, new_n16659, new_n16660, new_n16661, new_n16662,
    new_n16663, new_n16664, new_n16665, new_n16666, new_n16667, new_n16668,
    new_n16669, new_n16670, new_n16671, new_n16672, new_n16673, new_n16674,
    new_n16675, new_n16676, new_n16677, new_n16678, new_n16679, new_n16680,
    new_n16681, new_n16682, new_n16683, new_n16684, new_n16685, new_n16686,
    new_n16687, new_n16688, new_n16689, new_n16690, new_n16691, new_n16692,
    new_n16693, new_n16694, new_n16695, new_n16696, new_n16697, new_n16698,
    new_n16699, new_n16700, new_n16701, new_n16702, new_n16703, new_n16704,
    new_n16705, new_n16706, new_n16707, new_n16708, new_n16709, new_n16710,
    new_n16711, new_n16712, new_n16713, new_n16714, new_n16715, new_n16716,
    new_n16717, new_n16718, new_n16719, new_n16720, new_n16721, new_n16722,
    new_n16723, new_n16724, new_n16725, new_n16726, new_n16727, new_n16728,
    new_n16729, new_n16730, new_n16731, new_n16732, new_n16733, new_n16734,
    new_n16735, new_n16736, new_n16737, new_n16738, new_n16739, new_n16740,
    new_n16741, new_n16742, new_n16743, new_n16744, new_n16745, new_n16746,
    new_n16747, new_n16748, new_n16749, new_n16750, new_n16751, new_n16752,
    new_n16753, new_n16754, new_n16755, new_n16756, new_n16757, new_n16758,
    new_n16759, new_n16760, new_n16761, new_n16762, new_n16763, new_n16764,
    new_n16765, new_n16766, new_n16767, new_n16768, new_n16769, new_n16770,
    new_n16771, new_n16772, new_n16773, new_n16774, new_n16775, new_n16776,
    new_n16777, new_n16778, new_n16779, new_n16780, new_n16781, new_n16782,
    new_n16783, new_n16784, new_n16785, new_n16786, new_n16787, new_n16788,
    new_n16789, new_n16790, new_n16791, new_n16792, new_n16793, new_n16794,
    new_n16795, new_n16796, new_n16797, new_n16798, new_n16799, new_n16800,
    new_n16801, new_n16802, new_n16803, new_n16804, new_n16805, new_n16806,
    new_n16807, new_n16808, new_n16809, new_n16810, new_n16811, new_n16812,
    new_n16813, new_n16814, new_n16815, new_n16816, new_n16817, new_n16818,
    new_n16819, new_n16820, new_n16821, new_n16822, new_n16823, new_n16824,
    new_n16825, new_n16826, new_n16827, new_n16828, new_n16829, new_n16830,
    new_n16831, new_n16832, new_n16833, new_n16834, new_n16835, new_n16836,
    new_n16837, new_n16838, new_n16839, new_n16840, new_n16841, new_n16842,
    new_n16843, new_n16844, new_n16845, new_n16846, new_n16847, new_n16848,
    new_n16849, new_n16850, new_n16851, new_n16852, new_n16853, new_n16854,
    new_n16855, new_n16856, new_n16857, new_n16858, new_n16859, new_n16860,
    new_n16861, new_n16862, new_n16863, new_n16864, new_n16865, new_n16866,
    new_n16867, new_n16868, new_n16869, new_n16870, new_n16871, new_n16872,
    new_n16873, new_n16874, new_n16875, new_n16876, new_n16877, new_n16878,
    new_n16879, new_n16880, new_n16881, new_n16882, new_n16883, new_n16884,
    new_n16885, new_n16886, new_n16887, new_n16888, new_n16889, new_n16890,
    new_n16891, new_n16892, new_n16893, new_n16894, new_n16895, new_n16896,
    new_n16897, new_n16898, new_n16899, new_n16900, new_n16901, new_n16902,
    new_n16903, new_n16904, new_n16905, new_n16906, new_n16907, new_n16908,
    new_n16909, new_n16910, new_n16911, new_n16912, new_n16913, new_n16914,
    new_n16915, new_n16916, new_n16917, new_n16918, new_n16919, new_n16920,
    new_n16921, new_n16922, new_n16923, new_n16924, new_n16925, new_n16926,
    new_n16927, new_n16928, new_n16929, new_n16930, new_n16931, new_n16932,
    new_n16933, new_n16934, new_n16935, new_n16936, new_n16937, new_n16938,
    new_n16939, new_n16940, new_n16941, new_n16942, new_n16943, new_n16944,
    new_n16945, new_n16946, new_n16947, new_n16948, new_n16949, new_n16950,
    new_n16951, new_n16952, new_n16953, new_n16954, new_n16955, new_n16956,
    new_n16957, new_n16958, new_n16959, new_n16960, new_n16961, new_n16962,
    new_n16963, new_n16964, new_n16965, new_n16966, new_n16967, new_n16968,
    new_n16969, new_n16970, new_n16971, new_n16972, new_n16973, new_n16974,
    new_n16975, new_n16976, new_n16977, new_n16978, new_n16979, new_n16980,
    new_n16981, new_n16982, new_n16983, new_n16984, new_n16985, new_n16986,
    new_n16987, new_n16988, new_n16989, new_n16990, new_n16991, new_n16992,
    new_n16993, new_n16994, new_n16995, new_n16996, new_n16997, new_n16998,
    new_n16999, new_n17000, new_n17001, new_n17002, new_n17003, new_n17004,
    new_n17005, new_n17006, new_n17007, new_n17008, new_n17009, new_n17010,
    new_n17011, new_n17012, new_n17013, new_n17014, new_n17015, new_n17016,
    new_n17017, new_n17018, new_n17019, new_n17020, new_n17021, new_n17022,
    new_n17023, new_n17024, new_n17025, new_n17026, new_n17027, new_n17028,
    new_n17029, new_n17030, new_n17031, new_n17032, new_n17033, new_n17034,
    new_n17035, new_n17036, new_n17037, new_n17038, new_n17039, new_n17040,
    new_n17041, new_n17042, new_n17043, new_n17044, new_n17045, new_n17046,
    new_n17047, new_n17048, new_n17049, new_n17050, new_n17051, new_n17052,
    new_n17053, new_n17054, new_n17055, new_n17056, new_n17057, new_n17058,
    new_n17059, new_n17060, new_n17061, new_n17062, new_n17063, new_n17064,
    new_n17065, new_n17066, new_n17067, new_n17068, new_n17069, new_n17070,
    new_n17071, new_n17072, new_n17073, new_n17074, new_n17075, new_n17076,
    new_n17077, new_n17078, new_n17079, new_n17080, new_n17081, new_n17082,
    new_n17083, new_n17084, new_n17085, new_n17086, new_n17087, new_n17088,
    new_n17089, new_n17090, new_n17091, new_n17092, new_n17093, new_n17094,
    new_n17095, new_n17096, new_n17097, new_n17098, new_n17099, new_n17100,
    new_n17101, new_n17102, new_n17103, new_n17104, new_n17105, new_n17106,
    new_n17107, new_n17108, new_n17109, new_n17110, new_n17111, new_n17112,
    new_n17113, new_n17114, new_n17115, new_n17116, new_n17117, new_n17118,
    new_n17119, new_n17120, new_n17121, new_n17122, new_n17123, new_n17124,
    new_n17125, new_n17126, new_n17127, new_n17128, new_n17129, new_n17130,
    new_n17131, new_n17132, new_n17133, new_n17134, new_n17135, new_n17136,
    new_n17137, new_n17138, new_n17139, new_n17140, new_n17141, new_n17142,
    new_n17143, new_n17144, new_n17145, new_n17146, new_n17147, new_n17148,
    new_n17149, new_n17150, new_n17151, new_n17152, new_n17153, new_n17154,
    new_n17155, new_n17156, new_n17157, new_n17158, new_n17159, new_n17160,
    new_n17161, new_n17162, new_n17163, new_n17164, new_n17165, new_n17166,
    new_n17167, new_n17168, new_n17169, new_n17170, new_n17171, new_n17172,
    new_n17173, new_n17174, new_n17175, new_n17176, new_n17177, new_n17178,
    new_n17179, new_n17180, new_n17181, new_n17182, new_n17183, new_n17184,
    new_n17185, new_n17186, new_n17187, new_n17188, new_n17189, new_n17190,
    new_n17191, new_n17192, new_n17193, new_n17194, new_n17195, new_n17196,
    new_n17197, new_n17198, new_n17199, new_n17200, new_n17201, new_n17202,
    new_n17203, new_n17204, new_n17205, new_n17206, new_n17207, new_n17208,
    new_n17209, new_n17210, new_n17211, new_n17212, new_n17213, new_n17214,
    new_n17215, new_n17216, new_n17217, new_n17218, new_n17219, new_n17220,
    new_n17221, new_n17222, new_n17223, new_n17224, new_n17225, new_n17226,
    new_n17227, new_n17228, new_n17229, new_n17230, new_n17231, new_n17232,
    new_n17233, new_n17234, new_n17235, new_n17236, new_n17237, new_n17238,
    new_n17239, new_n17240, new_n17241, new_n17242, new_n17243, new_n17244,
    new_n17245, new_n17246, new_n17247, new_n17248, new_n17249, new_n17250,
    new_n17251, new_n17252, new_n17253, new_n17254, new_n17255, new_n17256,
    new_n17257, new_n17258, new_n17259, new_n17260, new_n17261, new_n17262,
    new_n17263, new_n17264, new_n17265, new_n17266, new_n17267, new_n17268,
    new_n17269, new_n17270, new_n17271, new_n17272, new_n17273, new_n17274,
    new_n17275, new_n17276, new_n17277, new_n17278, new_n17279, new_n17280,
    new_n17281, new_n17282, new_n17283, new_n17284, new_n17285, new_n17286,
    new_n17287, new_n17288, new_n17289, new_n17290, new_n17291, new_n17292,
    new_n17293, new_n17294, new_n17295, new_n17296, new_n17297, new_n17298,
    new_n17299, new_n17300, new_n17301, new_n17302, new_n17303, new_n17304,
    new_n17305, new_n17306, new_n17307, new_n17308, new_n17309, new_n17310,
    new_n17311, new_n17312, new_n17313, new_n17314, new_n17315, new_n17316,
    new_n17317, new_n17318, new_n17319, new_n17320, new_n17321, new_n17322,
    new_n17323, new_n17324, new_n17325, new_n17326, new_n17327, new_n17328,
    new_n17329, new_n17330, new_n17331, new_n17332, new_n17333, new_n17334,
    new_n17335, new_n17336, new_n17337, new_n17338, new_n17339, new_n17340,
    new_n17341, new_n17342, new_n17343, new_n17344, new_n17345, new_n17346,
    new_n17347, new_n17348, new_n17349, new_n17350, new_n17351, new_n17352,
    new_n17353, new_n17354, new_n17355, new_n17356, new_n17357, new_n17358,
    new_n17359, new_n17360, new_n17361, new_n17362, new_n17363, new_n17364,
    new_n17365, new_n17366, new_n17367, new_n17368, new_n17369, new_n17370,
    new_n17371, new_n17372, new_n17373, new_n17374, new_n17375, new_n17376,
    new_n17377, new_n17378, new_n17379, new_n17380, new_n17381, new_n17382,
    new_n17383, new_n17384, new_n17385, new_n17386, new_n17387, new_n17388,
    new_n17389, new_n17390, new_n17391, new_n17392, new_n17393, new_n17394,
    new_n17395, new_n17396, new_n17397, new_n17398, new_n17399, new_n17400,
    new_n17401, new_n17402, new_n17403, new_n17404, new_n17405, new_n17406,
    new_n17407, new_n17408, new_n17409, new_n17410, new_n17411, new_n17412,
    new_n17413, new_n17414, new_n17415, new_n17416, new_n17417, new_n17418,
    new_n17419, new_n17420, new_n17421, new_n17422, new_n17423, new_n17424,
    new_n17425, new_n17426, new_n17427, new_n17428, new_n17429, new_n17430,
    new_n17431, new_n17432, new_n17433, new_n17434, new_n17435, new_n17436,
    new_n17437, new_n17438, new_n17439, new_n17440, new_n17441, new_n17442,
    new_n17443, new_n17444, new_n17445, new_n17446, new_n17447, new_n17448,
    new_n17449, new_n17450, new_n17451, new_n17452, new_n17453, new_n17454,
    new_n17455, new_n17456, new_n17457, new_n17458, new_n17459, new_n17460,
    new_n17461, new_n17462, new_n17463, new_n17464, new_n17465, new_n17466,
    new_n17467, new_n17468, new_n17469, new_n17470, new_n17471, new_n17472,
    new_n17473, new_n17474, new_n17475, new_n17476, new_n17477, new_n17478,
    new_n17479, new_n17480, new_n17481, new_n17482, new_n17483, new_n17484,
    new_n17485, new_n17486, new_n17487, new_n17488, new_n17489, new_n17490,
    new_n17491, new_n17492, new_n17493, new_n17494, new_n17495, new_n17496,
    new_n17497, new_n17498, new_n17499, new_n17500, new_n17501, new_n17502,
    new_n17503, new_n17504, new_n17505, new_n17506, new_n17507, new_n17508,
    new_n17509, new_n17510, new_n17511, new_n17512, new_n17513, new_n17514,
    new_n17515, new_n17516, new_n17517, new_n17518, new_n17519, new_n17520,
    new_n17521, new_n17522, new_n17523, new_n17524, new_n17525, new_n17526,
    new_n17527, new_n17528, new_n17529, new_n17530, new_n17531, new_n17532,
    new_n17533, new_n17534, new_n17535, new_n17536, new_n17537, new_n17538,
    new_n17539, new_n17540, new_n17541, new_n17542, new_n17543, new_n17544,
    new_n17545, new_n17546, new_n17547, new_n17548, new_n17549, new_n17550,
    new_n17551, new_n17552, new_n17553, new_n17554, new_n17555, new_n17556,
    new_n17557, new_n17558, new_n17559, new_n17560, new_n17561, new_n17562,
    new_n17563, new_n17564, new_n17565, new_n17566, new_n17567, new_n17568,
    new_n17569, new_n17570, new_n17571, new_n17572, new_n17573, new_n17574,
    new_n17575, new_n17576, new_n17577, new_n17578, new_n17579, new_n17580,
    new_n17581, new_n17582, new_n17583, new_n17584, new_n17585, new_n17586,
    new_n17587, new_n17588, new_n17589, new_n17590, new_n17591, new_n17592,
    new_n17593, new_n17594, new_n17595, new_n17596, new_n17597, new_n17598,
    new_n17599, new_n17600, new_n17601, new_n17602, new_n17603, new_n17604,
    new_n17605, new_n17606, new_n17607, new_n17608, new_n17609, new_n17610,
    new_n17611, new_n17612, new_n17613, new_n17614, new_n17615, new_n17616,
    new_n17617, new_n17618, new_n17619, new_n17620, new_n17621, new_n17622,
    new_n17623, new_n17624, new_n17625, new_n17626, new_n17627, new_n17628,
    new_n17629, new_n17630, new_n17631, new_n17632, new_n17633, new_n17634,
    new_n17635, new_n17636, new_n17637, new_n17638, new_n17639, new_n17640,
    new_n17641, new_n17642, new_n17643, new_n17644, new_n17645, new_n17646,
    new_n17647, new_n17648, new_n17649, new_n17650, new_n17651, new_n17652,
    new_n17653, new_n17654, new_n17655, new_n17656, new_n17657, new_n17658,
    new_n17659, new_n17660, new_n17661, new_n17662, new_n17663, new_n17664,
    new_n17665, new_n17666, new_n17667, new_n17668, new_n17669, new_n17670,
    new_n17671, new_n17672, new_n17673, new_n17674, new_n17675, new_n17676,
    new_n17677, new_n17678, new_n17679, new_n17680, new_n17681, new_n17682,
    new_n17683, new_n17684, new_n17685, new_n17686, new_n17687, new_n17688,
    new_n17689, new_n17690, new_n17691, new_n17692, new_n17693, new_n17694,
    new_n17695, new_n17696, new_n17697, new_n17698, new_n17699, new_n17700,
    new_n17701, new_n17702, new_n17703, new_n17704, new_n17705, new_n17706,
    new_n17707, new_n17708, new_n17709, new_n17710, new_n17711, new_n17712,
    new_n17713, new_n17714, new_n17715, new_n17716, new_n17717, new_n17718,
    new_n17719, new_n17720, new_n17721, new_n17722, new_n17723, new_n17724,
    new_n17725, new_n17726, new_n17727, new_n17728, new_n17729, new_n17730,
    new_n17731, new_n17732, new_n17733, new_n17734, new_n17735, new_n17736,
    new_n17737, new_n17738, new_n17739, new_n17740, new_n17741, new_n17742,
    new_n17743, new_n17744, new_n17745, new_n17746, new_n17747, new_n17748,
    new_n17749, new_n17750, new_n17751, new_n17752, new_n17753, new_n17754,
    new_n17755, new_n17756, new_n17757, new_n17758, new_n17759, new_n17760,
    new_n17761, new_n17762, new_n17763, new_n17764, new_n17765, new_n17766,
    new_n17767, new_n17768, new_n17769, new_n17770, new_n17771, new_n17772,
    new_n17773, new_n17774, new_n17775, new_n17776, new_n17777, new_n17778,
    new_n17779, new_n17780, new_n17781, new_n17782, new_n17783, new_n17784,
    new_n17785, new_n17786, new_n17787, new_n17788, new_n17789, new_n17790,
    new_n17791, new_n17792, new_n17793, new_n17794, new_n17795, new_n17796,
    new_n17797, new_n17798, new_n17799, new_n17800, new_n17801, new_n17802,
    new_n17803, new_n17804, new_n17805, new_n17806, new_n17807, new_n17808,
    new_n17809, new_n17810, new_n17811, new_n17812, new_n17813, new_n17814,
    new_n17815, new_n17816, new_n17817, new_n17818, new_n17819, new_n17820,
    new_n17821, new_n17822, new_n17823, new_n17824, new_n17825, new_n17826,
    new_n17827, new_n17828, new_n17829, new_n17830, new_n17831, new_n17832,
    new_n17833, new_n17834, new_n17835, new_n17836, new_n17837, new_n17838,
    new_n17839, new_n17840, new_n17841, new_n17842, new_n17843, new_n17844,
    new_n17845, new_n17846, new_n17847, new_n17848, new_n17849, new_n17850,
    new_n17851, new_n17852, new_n17853, new_n17854, new_n17855, new_n17856,
    new_n17857, new_n17858, new_n17859, new_n17860, new_n17861, new_n17862,
    new_n17863, new_n17864, new_n17865, new_n17866, new_n17867, new_n17868,
    new_n17869, new_n17870, new_n17871, new_n17872, new_n17873, new_n17874,
    new_n17875, new_n17876, new_n17877, new_n17878, new_n17879, new_n17880,
    new_n17881, new_n17882, new_n17883, new_n17884, new_n17885, new_n17886,
    new_n17887, new_n17888, new_n17889, new_n17890, new_n17891, new_n17892,
    new_n17893, new_n17894, new_n17895, new_n17896, new_n17897, new_n17898,
    new_n17899, new_n17900, new_n17901, new_n17902, new_n17903, new_n17904,
    new_n17905, new_n17906, new_n17907, new_n17908, new_n17909, new_n17910,
    new_n17911, new_n17912, new_n17913, new_n17914, new_n17915, new_n17916,
    new_n17917, new_n17918, new_n17919, new_n17920, new_n17921, new_n17922,
    new_n17923, new_n17924, new_n17925, new_n17926, new_n17927, new_n17928,
    new_n17929, new_n17930, new_n17931, new_n17932, new_n17933, new_n17934,
    new_n17935, new_n17936, new_n17937, new_n17938, new_n17939, new_n17940,
    new_n17941, new_n17942, new_n17943, new_n17944, new_n17945, new_n17946,
    new_n17947, new_n17948, new_n17949, new_n17950, new_n17951, new_n17952,
    new_n17953, new_n17954, new_n17955, new_n17956, new_n17957, new_n17958,
    new_n17959, new_n17960, new_n17961, new_n17962, new_n17963, new_n17964,
    new_n17965, new_n17966, new_n17967, new_n17968, new_n17969, new_n17970,
    new_n17971, new_n17972, new_n17973, new_n17974, new_n17975, new_n17976,
    new_n17977, new_n17978, new_n17979, new_n17980, new_n17981, new_n17982,
    new_n17983, new_n17984, new_n17985, new_n17986, new_n17987, new_n17988,
    new_n17989, new_n17990, new_n17991, new_n17992, new_n17993, new_n17994,
    new_n17995, new_n17996, new_n17997, new_n17998, new_n17999, new_n18000,
    new_n18001, new_n18002, new_n18003, new_n18004, new_n18005, new_n18006,
    new_n18007, new_n18008, new_n18009, new_n18010, new_n18011, new_n18012,
    new_n18013, new_n18014, new_n18015, new_n18016, new_n18017, new_n18018,
    new_n18019, new_n18020, new_n18021, new_n18022, new_n18023, new_n18024,
    new_n18025, new_n18026, new_n18027, new_n18028, new_n18029, new_n18030,
    new_n18031, new_n18032, new_n18033, new_n18034, new_n18035, new_n18036,
    new_n18037, new_n18038, new_n18039, new_n18040, new_n18041, new_n18042,
    new_n18043, new_n18044, new_n18045, new_n18046, new_n18047, new_n18048,
    new_n18049, new_n18050, new_n18051, new_n18052, new_n18053, new_n18054,
    new_n18055, new_n18056, new_n18057, new_n18058, new_n18059, new_n18060,
    new_n18061, new_n18062, new_n18063, new_n18064, new_n18065, new_n18066,
    new_n18067, new_n18068, new_n18069, new_n18070, new_n18071, new_n18072,
    new_n18073, new_n18074, new_n18075, new_n18076, new_n18077, new_n18078,
    new_n18079, new_n18080, new_n18081, new_n18082, new_n18083, new_n18084,
    new_n18085, new_n18086, new_n18087, new_n18088, new_n18089, new_n18090,
    new_n18091, new_n18092, new_n18093, new_n18094, new_n18095, new_n18096,
    new_n18097, new_n18098, new_n18099, new_n18100, new_n18101, new_n18102,
    new_n18103, new_n18104, new_n18105, new_n18106, new_n18107, new_n18108,
    new_n18109, new_n18110, new_n18111, new_n18112, new_n18113, new_n18114,
    new_n18115, new_n18116, new_n18117, new_n18118, new_n18119, new_n18120,
    new_n18121, new_n18122, new_n18123, new_n18124, new_n18125, new_n18126,
    new_n18127, new_n18128, new_n18129, new_n18130, new_n18131, new_n18132,
    new_n18133, new_n18134, new_n18135, new_n18136, new_n18137, new_n18138,
    new_n18139, new_n18140, new_n18141, new_n18142, new_n18143, new_n18144,
    new_n18145, new_n18146, new_n18147, new_n18148, new_n18149, new_n18150,
    new_n18151, new_n18152, new_n18153, new_n18154, new_n18155, new_n18156,
    new_n18157, new_n18158, new_n18159, new_n18160, new_n18161, new_n18162,
    new_n18163, new_n18164, new_n18165, new_n18166, new_n18167, new_n18168,
    new_n18169, new_n18170, new_n18171, new_n18172, new_n18173, new_n18174,
    new_n18175, new_n18176, new_n18177, new_n18178, new_n18179, new_n18180,
    new_n18181, new_n18182, new_n18183, new_n18184, new_n18185, new_n18186,
    new_n18187, new_n18188, new_n18189, new_n18190, new_n18191, new_n18192,
    new_n18193, new_n18194, new_n18195, new_n18196, new_n18197, new_n18198,
    new_n18199, new_n18200, new_n18201, new_n18202, new_n18203, new_n18204,
    new_n18205, new_n18206, new_n18207, new_n18208, new_n18209, new_n18210,
    new_n18211, new_n18212, new_n18213, new_n18214, new_n18215, new_n18216,
    new_n18217, new_n18218, new_n18219, new_n18220, new_n18221, new_n18222,
    new_n18223, new_n18224, new_n18225, new_n18226, new_n18227, new_n18228,
    new_n18229, new_n18230, new_n18231, new_n18232, new_n18233, new_n18234,
    new_n18235, new_n18236, new_n18237, new_n18238, new_n18239, new_n18240,
    new_n18241, new_n18242, new_n18243, new_n18244, new_n18245, new_n18246,
    new_n18247, new_n18248, new_n18249, new_n18250, new_n18251, new_n18252,
    new_n18253, new_n18254, new_n18255, new_n18256, new_n18257, new_n18258,
    new_n18259, new_n18260, new_n18261, new_n18262, new_n18263, new_n18264,
    new_n18265, new_n18266, new_n18267, new_n18268, new_n18269, new_n18270,
    new_n18271, new_n18272, new_n18273, new_n18274, new_n18275, new_n18276,
    new_n18277, new_n18278, new_n18279, new_n18280, new_n18281, new_n18282,
    new_n18283, new_n18284, new_n18285, new_n18286, new_n18287, new_n18288,
    new_n18289, new_n18290, new_n18291, new_n18292, new_n18293, new_n18294,
    new_n18295, new_n18296, new_n18297, new_n18298, new_n18299, new_n18300,
    new_n18301, new_n18302, new_n18303, new_n18304, new_n18305, new_n18306,
    new_n18307, new_n18308, new_n18309, new_n18310, new_n18311, new_n18312,
    new_n18313, new_n18314, new_n18315, new_n18316, new_n18317, new_n18318,
    new_n18319, new_n18320, new_n18321, new_n18322, new_n18323, new_n18324,
    new_n18325, new_n18326, new_n18327, new_n18328, new_n18329, new_n18330,
    new_n18331, new_n18332, new_n18333, new_n18334, new_n18335, new_n18336,
    new_n18337, new_n18338, new_n18339, new_n18340, new_n18341, new_n18342,
    new_n18343, new_n18344, new_n18345, new_n18346, new_n18347, new_n18348,
    new_n18349, new_n18350, new_n18351, new_n18352, new_n18353, new_n18354,
    new_n18355, new_n18356, new_n18357, new_n18358, new_n18359, new_n18360,
    new_n18361, new_n18362, new_n18363, new_n18364, new_n18365, new_n18366,
    new_n18367, new_n18368, new_n18369, new_n18370, new_n18371, new_n18372,
    new_n18373, new_n18374, new_n18375, new_n18376, new_n18377, new_n18378,
    new_n18379, new_n18380, new_n18381, new_n18382, new_n18383, new_n18384,
    new_n18385, new_n18386, new_n18387, new_n18388, new_n18389, new_n18390,
    new_n18391, new_n18392, new_n18393, new_n18394, new_n18395, new_n18396,
    new_n18397, new_n18398, new_n18399, new_n18400, new_n18401, new_n18402,
    new_n18403, new_n18404, new_n18405, new_n18406, new_n18407, new_n18408,
    new_n18409, new_n18410, new_n18411, new_n18412, new_n18413, new_n18414,
    new_n18415, new_n18416, new_n18417, new_n18418, new_n18419, new_n18420,
    new_n18421, new_n18422, new_n18423, new_n18424, new_n18425, new_n18426,
    new_n18427, new_n18428, new_n18429, new_n18430, new_n18431, new_n18432,
    new_n18433, new_n18434, new_n18435, new_n18436, new_n18437, new_n18438,
    new_n18439, new_n18440, new_n18441, new_n18442, new_n18443, new_n18444,
    new_n18445, new_n18446, new_n18447, new_n18448, new_n18449, new_n18450,
    new_n18451, new_n18452, new_n18453, new_n18454, new_n18455, new_n18456,
    new_n18457, new_n18458, new_n18459, new_n18460, new_n18461, new_n18462,
    new_n18463, new_n18464, new_n18465, new_n18466, new_n18467, new_n18468,
    new_n18469, new_n18470, new_n18471, new_n18472, new_n18473, new_n18474,
    new_n18475, new_n18476, new_n18477, new_n18478, new_n18479, new_n18480,
    new_n18481, new_n18482, new_n18483, new_n18484, new_n18485, new_n18486,
    new_n18487, new_n18488, new_n18489, new_n18490, new_n18491, new_n18492,
    new_n18493, new_n18494, new_n18495, new_n18496, new_n18497, new_n18498,
    new_n18499, new_n18500, new_n18501, new_n18502, new_n18503, new_n18504,
    new_n18505, new_n18506, new_n18507, new_n18508, new_n18509, new_n18510,
    new_n18511, new_n18512, new_n18513, new_n18514, new_n18515, new_n18516,
    new_n18517, new_n18518, new_n18519, new_n18520, new_n18521, new_n18522,
    new_n18523, new_n18524, new_n18525, new_n18526, new_n18527, new_n18528,
    new_n18529, new_n18530, new_n18531, new_n18532, new_n18533, new_n18534,
    new_n18535, new_n18536, new_n18537, new_n18538, new_n18539, new_n18540,
    new_n18541, new_n18542, new_n18543, new_n18544, new_n18545, new_n18546,
    new_n18547, new_n18548, new_n18549, new_n18550, new_n18551, new_n18552,
    new_n18553, new_n18554, new_n18555, new_n18556, new_n18557, new_n18558,
    new_n18559, new_n18560, new_n18561, new_n18562, new_n18563, new_n18564,
    new_n18565, new_n18566, new_n18567, new_n18568, new_n18569, new_n18570,
    new_n18571, new_n18572, new_n18573, new_n18574, new_n18575, new_n18576,
    new_n18577, new_n18578, new_n18579, new_n18580, new_n18581, new_n18582,
    new_n18583, new_n18584, new_n18585, new_n18586, new_n18587, new_n18588,
    new_n18589, new_n18590, new_n18591, new_n18592, new_n18593, new_n18594,
    new_n18595, new_n18596, new_n18597, new_n18598, new_n18599, new_n18600,
    new_n18601, new_n18602, new_n18603, new_n18604, new_n18605, new_n18606,
    new_n18607, new_n18608, new_n18609, new_n18610, new_n18611, new_n18612,
    new_n18613, new_n18614, new_n18615, new_n18616, new_n18617, new_n18618,
    new_n18619, new_n18620, new_n18621, new_n18622, new_n18623, new_n18624,
    new_n18625, new_n18626, new_n18627, new_n18628, new_n18629, new_n18630,
    new_n18631, new_n18632, new_n18633, new_n18634, new_n18635, new_n18636,
    new_n18637, new_n18638, new_n18639, new_n18640, new_n18641, new_n18642,
    new_n18643, new_n18644, new_n18645, new_n18646, new_n18647, new_n18648,
    new_n18649, new_n18650, new_n18651, new_n18652, new_n18653, new_n18654,
    new_n18655, new_n18656, new_n18657, new_n18658, new_n18659, new_n18660,
    new_n18661, new_n18662, new_n18663, new_n18664, new_n18665, new_n18666,
    new_n18667, new_n18668, new_n18669, new_n18670, new_n18671, new_n18672,
    new_n18673, new_n18674, new_n18675, new_n18676, new_n18677, new_n18678,
    new_n18679, new_n18680, new_n18681, new_n18682, new_n18683, new_n18684,
    new_n18685, new_n18686, new_n18687, new_n18688, new_n18689, new_n18690,
    new_n18691, new_n18692, new_n18693, new_n18694, new_n18695, new_n18696,
    new_n18697, new_n18698, new_n18699, new_n18700, new_n18701, new_n18702,
    new_n18703, new_n18704, new_n18705, new_n18706, new_n18707, new_n18708,
    new_n18709, new_n18710, new_n18711, new_n18712, new_n18713, new_n18714,
    new_n18715, new_n18716, new_n18717, new_n18718, new_n18719, new_n18720,
    new_n18721, new_n18722, new_n18723, new_n18724, new_n18725, new_n18726,
    new_n18727, new_n18728, new_n18729, new_n18730, new_n18731, new_n18732,
    new_n18733, new_n18734, new_n18735, new_n18736, new_n18737, new_n18738,
    new_n18739, new_n18740, new_n18741, new_n18742, new_n18743, new_n18744,
    new_n18745, new_n18746, new_n18747, new_n18748, new_n18749, new_n18750,
    new_n18751, new_n18752, new_n18753, new_n18754, new_n18755, new_n18756,
    new_n18757, new_n18758, new_n18759, new_n18760, new_n18761, new_n18762,
    new_n18763, new_n18764, new_n18765, new_n18766, new_n18767, new_n18768,
    new_n18769, new_n18770, new_n18771, new_n18772, new_n18773, new_n18774,
    new_n18775, new_n18776, new_n18777, new_n18778, new_n18779, new_n18780,
    new_n18781, new_n18782, new_n18783, new_n18784, new_n18785, new_n18786,
    new_n18787, new_n18788, new_n18789, new_n18790, new_n18791, new_n18792,
    new_n18793, new_n18794, new_n18795, new_n18796, new_n18797, new_n18798,
    new_n18799, new_n18800, new_n18801, new_n18802, new_n18803, new_n18804,
    new_n18805, new_n18806, new_n18807, new_n18808, new_n18809, new_n18810,
    new_n18811, new_n18812, new_n18813, new_n18814, new_n18815, new_n18816,
    new_n18817, new_n18818, new_n18819, new_n18820, new_n18821, new_n18822,
    new_n18823, new_n18824, new_n18825, new_n18826, new_n18827, new_n18828,
    new_n18829, new_n18830, new_n18831, new_n18832, new_n18833, new_n18834,
    new_n18835, new_n18836, new_n18837, new_n18838, new_n18839, new_n18840,
    new_n18841, new_n18842, new_n18843, new_n18844, new_n18845, new_n18846,
    new_n18847, new_n18848, new_n18849, new_n18850, new_n18851, new_n18852,
    new_n18853, new_n18854, new_n18855, new_n18856, new_n18857, new_n18858,
    new_n18859, new_n18860, new_n18861, new_n18862, new_n18863, new_n18864,
    new_n18865, new_n18866, new_n18867, new_n18868, new_n18869, new_n18870,
    new_n18871, new_n18872, new_n18873, new_n18874, new_n18875, new_n18876,
    new_n18877, new_n18878, new_n18879, new_n18880, new_n18881, new_n18882,
    new_n18883, new_n18884, new_n18885, new_n18886, new_n18887, new_n18888,
    new_n18889, new_n18890, new_n18891, new_n18892, new_n18893, new_n18894,
    new_n18895, new_n18896, new_n18897, new_n18898, new_n18899, new_n18900,
    new_n18901, new_n18902, new_n18903, new_n18904, new_n18905, new_n18906,
    new_n18907, new_n18908, new_n18909, new_n18910, new_n18911, new_n18912,
    new_n18913, new_n18914, new_n18915, new_n18916, new_n18917, new_n18918,
    new_n18919, new_n18920, new_n18921, new_n18922, new_n18923, new_n18924,
    new_n18925, new_n18926, new_n18927, new_n18928, new_n18929, new_n18930,
    new_n18931, new_n18932, new_n18933, new_n18934, new_n18935, new_n18936,
    new_n18937, new_n18938, new_n18939, new_n18940, new_n18941, new_n18942,
    new_n18943, new_n18944, new_n18945, new_n18946, new_n18947, new_n18948,
    new_n18949, new_n18950, new_n18951, new_n18952, new_n18953, new_n18954,
    new_n18955, new_n18956, new_n18957, new_n18958, new_n18959, new_n18960,
    new_n18961, new_n18962, new_n18963, new_n18964, new_n18965, new_n18966,
    new_n18967, new_n18968, new_n18969, new_n18970, new_n18971, new_n18972,
    new_n18973, new_n18974, new_n18975, new_n18976, new_n18977, new_n18978,
    new_n18979, new_n18980, new_n18981, new_n18982, new_n18983, new_n18984,
    new_n18985, new_n18986, new_n18987, new_n18988, new_n18989, new_n18990,
    new_n18991, new_n18992, new_n18993, new_n18994, new_n18995, new_n18996,
    new_n18997, new_n18998, new_n18999, new_n19000, new_n19001, new_n19002,
    new_n19003, new_n19004, new_n19005, new_n19006, new_n19007, new_n19008,
    new_n19009, new_n19010, new_n19011, new_n19012, new_n19013, new_n19014,
    new_n19015, new_n19016, new_n19017, new_n19018, new_n19019, new_n19020,
    new_n19021, new_n19022, new_n19023, new_n19024, new_n19025, new_n19026,
    new_n19027, new_n19028, new_n19029, new_n19030, new_n19031, new_n19032,
    new_n19033, new_n19034, new_n19035, new_n19036, new_n19037, new_n19038,
    new_n19039, new_n19040, new_n19041, new_n19042, new_n19043, new_n19044,
    new_n19045, new_n19046, new_n19047, new_n19048, new_n19049, new_n19050,
    new_n19051, new_n19052, new_n19053, new_n19054, new_n19055, new_n19056,
    new_n19057, new_n19058, new_n19059, new_n19060, new_n19061, new_n19062,
    new_n19063, new_n19064, new_n19065, new_n19066, new_n19067, new_n19068,
    new_n19069, new_n19070, new_n19071, new_n19072, new_n19073, new_n19074,
    new_n19075, new_n19076, new_n19077, new_n19078, new_n19079, new_n19080,
    new_n19081, new_n19082, new_n19083, new_n19084, new_n19085, new_n19086,
    new_n19087, new_n19088, new_n19089, new_n19090, new_n19091, new_n19092,
    new_n19093, new_n19094, new_n19095, new_n19096, new_n19097, new_n19098,
    new_n19099, new_n19100, new_n19101, new_n19102, new_n19103, new_n19104,
    new_n19105, new_n19106, new_n19107, new_n19108, new_n19109, new_n19110,
    new_n19111, new_n19112, new_n19113, new_n19114, new_n19115, new_n19116,
    new_n19117, new_n19118, new_n19119, new_n19120, new_n19121, new_n19122,
    new_n19123, new_n19124, new_n19125, new_n19126, new_n19127, new_n19128,
    new_n19129, new_n19130, new_n19131, new_n19132, new_n19133, new_n19134,
    new_n19135, new_n19136, new_n19137, new_n19138, new_n19139, new_n19140,
    new_n19141, new_n19142, new_n19143, new_n19144, new_n19145, new_n19146,
    new_n19147, new_n19148, new_n19149, new_n19150, new_n19151, new_n19152,
    new_n19153, new_n19154, new_n19155, new_n19156, new_n19157, new_n19158,
    new_n19159, new_n19160, new_n19161, new_n19162, new_n19163, new_n19164,
    new_n19165, new_n19166, new_n19167, new_n19168, new_n19169, new_n19170,
    new_n19171, new_n19172, new_n19173, new_n19174, new_n19175, new_n19176,
    new_n19177, new_n19178, new_n19179, new_n19180, new_n19181, new_n19182,
    new_n19183, new_n19184, new_n19185, new_n19186, new_n19187, new_n19188,
    new_n19189, new_n19190, new_n19191, new_n19192, new_n19193, new_n19194,
    new_n19195, new_n19196, new_n19197, new_n19198, new_n19199, new_n19200,
    new_n19201, new_n19202, new_n19203, new_n19204, new_n19205, new_n19206,
    new_n19207, new_n19208, new_n19209, new_n19210, new_n19211, new_n19212,
    new_n19213, new_n19214, new_n19215, new_n19216, new_n19217, new_n19218,
    new_n19219, new_n19220, new_n19221, new_n19222, new_n19223, new_n19224,
    new_n19225, new_n19226, new_n19227, new_n19228, new_n19229, new_n19230,
    new_n19231, new_n19232, new_n19233, new_n19234, new_n19235, new_n19236,
    new_n19237, new_n19238, new_n19239, new_n19240, new_n19241, new_n19242,
    new_n19243, new_n19244, new_n19245, new_n19246, new_n19247, new_n19248,
    new_n19249, new_n19250, new_n19251, new_n19252, new_n19253, new_n19254,
    new_n19255, new_n19256, new_n19257, new_n19258, new_n19259, new_n19260,
    new_n19261, new_n19262, new_n19263, new_n19264, new_n19265, new_n19266,
    new_n19267, new_n19268, new_n19269, new_n19270, new_n19271, new_n19272,
    new_n19273, new_n19274, new_n19275, new_n19276, new_n19277, new_n19278,
    new_n19279, new_n19280, new_n19281, new_n19282, new_n19283, new_n19284,
    new_n19285, new_n19286, new_n19287, new_n19288, new_n19289, new_n19290,
    new_n19291, new_n19292, new_n19293, new_n19294, new_n19295, new_n19296,
    new_n19297, new_n19298, new_n19299, new_n19300, new_n19301, new_n19302,
    new_n19303, new_n19304, new_n19305, new_n19306, new_n19307, new_n19308,
    new_n19309, new_n19310, new_n19311, new_n19312, new_n19313, new_n19314,
    new_n19315, new_n19316, new_n19317, new_n19318, new_n19319, new_n19320,
    new_n19321, new_n19322, new_n19323, new_n19324, new_n19325, new_n19326,
    new_n19327, new_n19328, new_n19329, new_n19330, new_n19331, new_n19332,
    new_n19333, new_n19334, new_n19335, new_n19336, new_n19337, new_n19338,
    new_n19339, new_n19340, new_n19341, new_n19342, new_n19343, new_n19344,
    new_n19345, new_n19346, new_n19347, new_n19348, new_n19349, new_n19350,
    new_n19351, new_n19352, new_n19353, new_n19354, new_n19355, new_n19356,
    new_n19357, new_n19358, new_n19359, new_n19360, new_n19361, new_n19362,
    new_n19363, new_n19364, new_n19365, new_n19366, new_n19367, new_n19368,
    new_n19369, new_n19370, new_n19371, new_n19372, new_n19373, new_n19374,
    new_n19375, new_n19376, new_n19377, new_n19378, new_n19379, new_n19380,
    new_n19381, new_n19382, new_n19383, new_n19384, new_n19385, new_n19386,
    new_n19387, new_n19388, new_n19389, new_n19390, new_n19391, new_n19392,
    new_n19393, new_n19394, new_n19395, new_n19396, new_n19397, new_n19398,
    new_n19399, new_n19400, new_n19401, new_n19402, new_n19403, new_n19404,
    new_n19405, new_n19406, new_n19407, new_n19408, new_n19409, new_n19410,
    new_n19411, new_n19412, new_n19413, new_n19414, new_n19415, new_n19416,
    new_n19417, new_n19418, new_n19419, new_n19420, new_n19421, new_n19422,
    new_n19423, new_n19424, new_n19425, new_n19426, new_n19427, new_n19428,
    new_n19429, new_n19430, new_n19431, new_n19432, new_n19433, new_n19434,
    new_n19435, new_n19436, new_n19437, new_n19438, new_n19439, new_n19440,
    new_n19441, new_n19442, new_n19443, new_n19444, new_n19445, new_n19446,
    new_n19447, new_n19448, new_n19449, new_n19450, new_n19451, new_n19452,
    new_n19453, new_n19454, new_n19455, new_n19456, new_n19457, new_n19458,
    new_n19459, new_n19460, new_n19461, new_n19462, new_n19463, new_n19464,
    new_n19465, new_n19466, new_n19467, new_n19468, new_n19469, new_n19470,
    new_n19471, new_n19472, new_n19473, new_n19474, new_n19475, new_n19476,
    new_n19477, new_n19478, new_n19479, new_n19480, new_n19481, new_n19482,
    new_n19483, new_n19484, new_n19485, new_n19486, new_n19487, new_n19488,
    new_n19489, new_n19490, new_n19491, new_n19492, new_n19493, new_n19494,
    new_n19495, new_n19496, new_n19497, new_n19498, new_n19499, new_n19500,
    new_n19501, new_n19502, new_n19503, new_n19504, new_n19505, new_n19506,
    new_n19507, new_n19508, new_n19509, new_n19510, new_n19511, new_n19512,
    new_n19513, new_n19514, new_n19515, new_n19516, new_n19517, new_n19518,
    new_n19519, new_n19520, new_n19521, new_n19522, new_n19523, new_n19524,
    new_n19525, new_n19526, new_n19527, new_n19528, new_n19529, new_n19530,
    new_n19531, new_n19532, new_n19533, new_n19534, new_n19535, new_n19536,
    new_n19537, new_n19538, new_n19539, new_n19540, new_n19541, new_n19542,
    new_n19543, new_n19544, new_n19545, new_n19546, new_n19547, new_n19548,
    new_n19549, new_n19550, new_n19551, new_n19552, new_n19553, new_n19554,
    new_n19555, new_n19556, new_n19557, new_n19558, new_n19559, new_n19560,
    new_n19561, new_n19562, new_n19563, new_n19564, new_n19565, new_n19566,
    new_n19567, new_n19568, new_n19569, new_n19570, new_n19571, new_n19572,
    new_n19573, new_n19574, new_n19575, new_n19576, new_n19577, new_n19578,
    new_n19579, new_n19580, new_n19581, new_n19582, new_n19583, new_n19584,
    new_n19585, new_n19586, new_n19587, new_n19588, new_n19589, new_n19590,
    new_n19591, new_n19592, new_n19593, new_n19594, new_n19595, new_n19596,
    new_n19597, new_n19598, new_n19599, new_n19600, new_n19601, new_n19602,
    new_n19603, new_n19604, new_n19605, new_n19606, new_n19607, new_n19608,
    new_n19609, new_n19610, new_n19611, new_n19612, new_n19613, new_n19614,
    new_n19615, new_n19616, new_n19617, new_n19618, new_n19619, new_n19620,
    new_n19621, new_n19622, new_n19623, new_n19624, new_n19625, new_n19626,
    new_n19627, new_n19628, new_n19629, new_n19630, new_n19631, new_n19632,
    new_n19633, new_n19634, new_n19635, new_n19636, new_n19637, new_n19638,
    new_n19639, new_n19640, new_n19641, new_n19642, new_n19643, new_n19644,
    new_n19645, new_n19646, new_n19647, new_n19648, new_n19649, new_n19650,
    new_n19651, new_n19652, new_n19653, new_n19654, new_n19655, new_n19656,
    new_n19657, new_n19658, new_n19659, new_n19660, new_n19661, new_n19662,
    new_n19663, new_n19664, new_n19665, new_n19666, new_n19667, new_n19668,
    new_n19669, new_n19670, new_n19671, new_n19672, new_n19673, new_n19674,
    new_n19675, new_n19676, new_n19677, new_n19678, new_n19679, new_n19680,
    new_n19681, new_n19682, new_n19683, new_n19684, new_n19685, new_n19686,
    new_n19687, new_n19688, new_n19689, new_n19690, new_n19691, new_n19692,
    new_n19693, new_n19694, new_n19695, new_n19696, new_n19697, new_n19698,
    new_n19699, new_n19700, new_n19701, new_n19702, new_n19703, new_n19704,
    new_n19705, new_n19706, new_n19707, new_n19708, new_n19709, new_n19710,
    new_n19711, new_n19712, new_n19713, new_n19714;
  assign new_n129 = n1 & n65;
  assign new_n130 = n1 & n66;
  assign new_n131 = n2 & n65;
  assign new_n132 = new_n131 ^ new_n130;
  assign new_n133 = n67 ^ n3;
  assign new_n134 = ~new_n133 & new_n129;
  assign new_n135 = n2 & n66;
  assign new_n136 = ~n65 & ~n67;
  assign new_n137 = new_n136 ^ n65;
  assign new_n138 = n1 & new_n137;
  assign new_n139 = new_n138 ^ new_n136;
  assign new_n140 = ~new_n135 & new_n139;
  assign new_n141 = new_n140 ^ new_n138;
  assign new_n142 = ~n1 & ~n3;
  assign new_n143 = new_n142 ^ n1;
  assign new_n144 = ~new_n143 & n65;
  assign new_n145 = new_n144 ^ n1;
  assign new_n146 = ~new_n141 & new_n145;
  assign new_n147 = new_n146 ^ new_n135;
  assign new_n148 = ~new_n134 & new_n147;
  assign new_n149 = n66 & n67;
  assign new_n150 = ~n65 & ~n66;
  assign new_n151 = new_n150 ^ n65;
  assign new_n152 = new_n151 ^ n66;
  assign new_n153 = ~n67 & new_n152;
  assign new_n154 = new_n153 ^ new_n149;
  assign new_n155 = n3 ^ n2;
  assign new_n156 = new_n154 & new_n155;
  assign new_n157 = new_n156 ^ n2;
  assign new_n158 = new_n157 ^ n68;
  assign new_n159 = ~n66 & n3;
  assign new_n160 = new_n159 ^ new_n133;
  assign new_n161 = ~n2 & new_n160;
  assign new_n162 = new_n161 ^ new_n133;
  assign new_n163 = new_n162 ^ new_n158;
  assign new_n164 = ~n1 & new_n163;
  assign new_n165 = new_n164 ^ new_n158;
  assign new_n166 = ~n66 & ~n67;
  assign new_n167 = ~n65 & new_n166;
  assign new_n168 = new_n167 ^ n65;
  assign new_n169 = n1 & n3;
  assign new_n170 = new_n169 ^ n3;
  assign new_n171 = new_n169 ^ new_n135;
  assign new_n172 = new_n171 ^ new_n169;
  assign new_n173 = new_n170 & new_n172;
  assign new_n174 = new_n173 ^ new_n169;
  assign new_n175 = ~new_n168 & new_n174;
  assign new_n176 = n4 & n65;
  assign new_n177 = new_n176 ^ n3;
  assign new_n178 = new_n177 ^ new_n175;
  assign new_n179 = new_n178 ^ new_n165;
  assign new_n180 = ~n2 & n3;
  assign new_n181 = n67 & new_n180;
  assign new_n182 = n2 & n68;
  assign new_n183 = new_n182 ^ new_n181;
  assign new_n184 = new_n183 ^ n3;
  assign new_n185 = ~n68 & ~new_n149;
  assign new_n186 = ~new_n153 & n68;
  assign new_n187 = new_n186 ^ new_n185;
  assign new_n188 = new_n155 & new_n187;
  assign new_n189 = new_n188 ^ n2;
  assign new_n190 = new_n189 ^ n69;
  assign new_n191 = new_n190 ^ new_n184;
  assign new_n192 = ~n1 & new_n191;
  assign new_n193 = new_n192 ^ new_n190;
  assign new_n194 = n3 & n4;
  assign new_n195 = new_n194 ^ n5;
  assign new_n196 = ~n65 & new_n195;
  assign new_n197 = n4 ^ n3;
  assign new_n198 = n66 ^ n4;
  assign new_n199 = ~new_n198 & new_n197;
  assign new_n200 = new_n199 ^ n3;
  assign new_n201 = new_n200 ^ n5;
  assign new_n202 = new_n201 ^ new_n196;
  assign new_n203 = new_n202 ^ new_n193;
  assign new_n204 = new_n165 & new_n178;
  assign new_n205 = new_n204 ^ new_n203;
  assign new_n206 = n6 ^ n5;
  assign new_n207 = ~new_n206 & new_n197;
  assign new_n208 = new_n207 ^ new_n197;
  assign new_n209 = ~new_n151 & new_n208;
  assign new_n210 = ~new_n197 & n6;
  assign new_n211 = new_n210 ^ new_n194;
  assign new_n212 = new_n206 & new_n211;
  assign new_n213 = n65 & new_n212;
  assign new_n214 = new_n213 ^ new_n209;
  assign new_n215 = n67 & new_n197;
  assign new_n216 = new_n215 ^ new_n214;
  assign new_n217 = ~new_n197 & n5;
  assign new_n218 = new_n217 ^ new_n194;
  assign new_n219 = n66 & new_n218;
  assign new_n220 = new_n219 ^ new_n216;
  assign new_n221 = n5 ^ n3;
  assign new_n222 = ~new_n197 & ~new_n221;
  assign new_n223 = n6 & new_n222;
  assign new_n224 = new_n223 ^ new_n210;
  assign new_n225 = new_n224 ^ n66;
  assign new_n226 = new_n225 ^ new_n224;
  assign new_n227 = new_n223 ^ n6;
  assign new_n228 = new_n227 ^ new_n224;
  assign new_n229 = ~new_n226 & new_n228;
  assign new_n230 = new_n229 ^ new_n224;
  assign new_n231 = ~n65 & new_n230;
  assign new_n232 = new_n231 ^ new_n223;
  assign new_n233 = new_n232 ^ n6;
  assign new_n234 = new_n233 ^ new_n220;
  assign new_n235 = ~new_n185 & n69;
  assign new_n236 = ~n69 & ~new_n186;
  assign new_n237 = new_n236 ^ new_n235;
  assign new_n238 = new_n155 & new_n237;
  assign new_n239 = new_n238 ^ n2;
  assign new_n240 = new_n239 ^ n70;
  assign new_n241 = n2 ^ n1;
  assign new_n242 = n69 ^ n3;
  assign new_n243 = n68 ^ n3;
  assign new_n244 = ~n68 & ~new_n243;
  assign new_n245 = new_n244 ^ new_n242;
  assign new_n246 = new_n245 ^ n68;
  assign new_n247 = ~new_n246 & new_n241;
  assign new_n248 = new_n247 ^ new_n244;
  assign new_n249 = new_n248 ^ n68;
  assign new_n250 = new_n249 ^ new_n240;
  assign new_n251 = ~n1 & ~new_n250;
  assign new_n252 = new_n251 ^ new_n240;
  assign new_n253 = new_n252 ^ new_n234;
  assign new_n254 = new_n204 ^ new_n202;
  assign new_n255 = ~new_n254 & new_n203;
  assign new_n256 = new_n255 ^ new_n193;
  assign new_n257 = new_n256 ^ new_n253;
  assign new_n258 = ~new_n220 & new_n232;
  assign new_n259 = new_n154 ^ n68;
  assign new_n260 = ~new_n259 & new_n208;
  assign new_n261 = n67 & new_n218;
  assign new_n262 = new_n261 ^ new_n260;
  assign new_n263 = n66 & new_n212;
  assign new_n264 = n68 & new_n207;
  assign new_n265 = new_n264 ^ new_n263;
  assign new_n266 = new_n265 ^ new_n262;
  assign new_n267 = new_n266 ^ n6;
  assign new_n268 = new_n267 ^ new_n258;
  assign new_n269 = n7 ^ n6;
  assign new_n270 = n65 & new_n269;
  assign new_n271 = new_n270 ^ new_n268;
  assign new_n272 = n69 & new_n180;
  assign new_n273 = n2 & n70;
  assign new_n274 = new_n273 ^ new_n272;
  assign new_n275 = new_n274 ^ n3;
  assign new_n276 = ~n70 & ~new_n235;
  assign new_n277 = ~new_n236 & n70;
  assign new_n278 = new_n277 ^ new_n276;
  assign new_n279 = new_n155 & new_n278;
  assign new_n280 = new_n279 ^ n2;
  assign new_n281 = new_n280 ^ n71;
  assign new_n282 = new_n281 ^ new_n275;
  assign new_n283 = ~n1 & new_n282;
  assign new_n284 = new_n283 ^ new_n281;
  assign new_n285 = new_n284 ^ new_n271;
  assign new_n286 = new_n256 ^ new_n252;
  assign new_n287 = ~new_n253 & new_n286;
  assign new_n288 = new_n287 ^ new_n256;
  assign new_n289 = new_n288 ^ new_n285;
  assign new_n290 = ~n6 & ~n7;
  assign new_n291 = new_n290 ^ new_n269;
  assign new_n292 = ~new_n290 & n66;
  assign new_n293 = ~n8 & n65;
  assign new_n294 = new_n293 ^ n65;
  assign new_n295 = new_n294 ^ new_n292;
  assign new_n296 = new_n291 & new_n295;
  assign new_n297 = ~new_n291 & n65;
  assign new_n298 = new_n297 ^ new_n296;
  assign new_n299 = ~new_n291 & ~new_n293;
  assign new_n300 = new_n299 ^ new_n291;
  assign new_n301 = new_n300 ^ new_n297;
  assign new_n302 = new_n301 ^ new_n298;
  assign new_n303 = n68 & new_n218;
  assign new_n304 = new_n187 ^ n69;
  assign new_n305 = ~new_n304 & new_n208;
  assign new_n306 = new_n305 ^ new_n303;
  assign new_n307 = n69 & new_n207;
  assign new_n308 = n67 & new_n212;
  assign new_n309 = new_n308 ^ new_n307;
  assign new_n310 = new_n309 ^ new_n306;
  assign new_n311 = new_n310 ^ n6;
  assign new_n312 = new_n311 ^ new_n302;
  assign new_n313 = ~new_n258 & ~new_n270;
  assign new_n314 = ~new_n313 & new_n267;
  assign new_n315 = new_n314 ^ new_n312;
  assign new_n316 = ~new_n276 & n71;
  assign new_n317 = ~n71 & ~new_n277;
  assign new_n318 = new_n317 ^ new_n316;
  assign new_n319 = new_n155 & new_n318;
  assign new_n320 = new_n319 ^ n2;
  assign new_n321 = new_n320 ^ n72;
  assign new_n322 = ~n70 & n3;
  assign new_n323 = n71 ^ n3;
  assign new_n324 = new_n323 ^ new_n322;
  assign new_n325 = n2 & new_n324;
  assign new_n326 = new_n325 ^ new_n322;
  assign new_n327 = new_n326 ^ new_n321;
  assign new_n328 = ~n1 & new_n327;
  assign new_n329 = new_n328 ^ new_n321;
  assign new_n330 = new_n329 ^ new_n315;
  assign new_n331 = new_n288 ^ new_n271;
  assign new_n332 = ~new_n285 & new_n331;
  assign new_n333 = new_n332 ^ new_n288;
  assign new_n334 = new_n333 ^ new_n330;
  assign new_n335 = new_n314 ^ new_n311;
  assign new_n336 = new_n312 & new_n335;
  assign new_n337 = new_n336 ^ new_n314;
  assign new_n338 = n69 & new_n218;
  assign new_n339 = new_n237 ^ n70;
  assign new_n340 = ~new_n339 & new_n208;
  assign new_n341 = new_n340 ^ new_n338;
  assign new_n342 = n70 & new_n207;
  assign new_n343 = n68 & new_n212;
  assign new_n344 = new_n343 ^ new_n342;
  assign new_n345 = new_n344 ^ new_n341;
  assign new_n346 = new_n345 ^ n6;
  assign new_n347 = n9 ^ n8;
  assign new_n348 = ~new_n347 & new_n269;
  assign new_n349 = new_n348 ^ new_n269;
  assign new_n350 = ~new_n151 & new_n349;
  assign new_n351 = n67 & new_n269;
  assign new_n352 = new_n351 ^ new_n350;
  assign new_n353 = n8 ^ n7;
  assign new_n354 = ~new_n269 & new_n353;
  assign new_n355 = n66 & new_n354;
  assign new_n356 = new_n355 ^ new_n352;
  assign new_n357 = new_n356 ^ new_n301;
  assign new_n358 = new_n290 & new_n293;
  assign new_n359 = new_n358 ^ new_n356;
  assign new_n360 = ~new_n270 & new_n302;
  assign new_n361 = new_n360 ^ new_n359;
  assign new_n362 = new_n361 ^ new_n357;
  assign new_n363 = ~n9 & new_n362;
  assign new_n364 = new_n363 ^ new_n361;
  assign new_n365 = new_n364 ^ new_n346;
  assign new_n366 = new_n365 ^ new_n337;
  assign new_n367 = n71 & new_n180;
  assign new_n368 = n2 & n72;
  assign new_n369 = new_n368 ^ new_n367;
  assign new_n370 = new_n369 ^ n3;
  assign new_n371 = n72 ^ n71;
  assign new_n372 = new_n318 & new_n371;
  assign new_n373 = ~new_n372 & new_n155;
  assign new_n374 = new_n373 ^ n2;
  assign new_n375 = new_n374 ^ n73;
  assign new_n376 = new_n375 ^ new_n370;
  assign new_n377 = ~n1 & new_n376;
  assign new_n378 = new_n377 ^ new_n375;
  assign new_n379 = new_n378 ^ new_n366;
  assign new_n380 = new_n333 ^ new_n315;
  assign new_n381 = ~new_n380 & new_n330;
  assign new_n382 = new_n381 ^ new_n333;
  assign new_n383 = new_n382 ^ new_n379;
  assign new_n384 = n9 & new_n361;
  assign new_n385 = ~new_n359 & new_n384;
  assign new_n386 = ~new_n259 & new_n349;
  assign new_n387 = n67 & new_n354;
  assign new_n388 = new_n387 ^ new_n386;
  assign new_n389 = ~n9 & ~new_n269;
  assign new_n390 = new_n389 ^ new_n290;
  assign new_n391 = new_n347 & new_n390;
  assign new_n392 = n66 & new_n391;
  assign new_n393 = n68 & new_n348;
  assign new_n394 = new_n393 ^ new_n392;
  assign new_n395 = new_n394 ^ new_n388;
  assign new_n396 = new_n395 ^ n9;
  assign new_n397 = n10 ^ n9;
  assign new_n398 = n65 & new_n397;
  assign new_n399 = new_n398 ^ new_n396;
  assign new_n400 = new_n399 ^ new_n385;
  assign new_n401 = n70 & new_n218;
  assign new_n402 = new_n278 ^ n71;
  assign new_n403 = ~new_n402 & new_n208;
  assign new_n404 = new_n403 ^ new_n401;
  assign new_n405 = n69 & new_n212;
  assign new_n406 = n71 & new_n207;
  assign new_n407 = new_n406 ^ new_n405;
  assign new_n408 = new_n407 ^ new_n404;
  assign new_n409 = new_n408 ^ n6;
  assign new_n410 = new_n409 ^ new_n400;
  assign new_n411 = new_n364 ^ new_n337;
  assign new_n412 = ~new_n411 & new_n365;
  assign new_n413 = new_n412 ^ new_n337;
  assign new_n414 = new_n413 ^ new_n410;
  assign new_n415 = n73 ^ n3;
  assign new_n416 = ~n72 & n3;
  assign new_n417 = new_n416 ^ new_n415;
  assign new_n418 = ~n2 & new_n417;
  assign new_n419 = new_n418 ^ new_n415;
  assign new_n420 = n73 ^ n72;
  assign new_n421 = ~n73 & n72;
  assign new_n422 = new_n421 ^ new_n420;
  assign new_n423 = ~new_n316 & new_n422;
  assign new_n424 = ~new_n317 & new_n421;
  assign new_n425 = new_n424 ^ new_n423;
  assign new_n426 = ~new_n425 & new_n155;
  assign new_n427 = new_n426 ^ n2;
  assign new_n428 = new_n427 ^ n74;
  assign new_n429 = new_n428 ^ new_n419;
  assign new_n430 = ~n1 & new_n429;
  assign new_n431 = new_n430 ^ new_n428;
  assign new_n432 = new_n431 ^ new_n414;
  assign new_n433 = new_n382 ^ new_n366;
  assign new_n434 = ~new_n433 & new_n379;
  assign new_n435 = new_n434 ^ new_n382;
  assign new_n436 = new_n435 ^ new_n432;
  assign new_n437 = ~new_n385 & ~new_n398;
  assign new_n438 = ~new_n437 & new_n396;
  assign new_n439 = n66 ^ n10;
  assign new_n440 = ~new_n439 & new_n397;
  assign new_n441 = new_n440 ^ n9;
  assign new_n442 = new_n441 ^ n11;
  assign new_n443 = ~n9 & ~n10;
  assign new_n444 = new_n443 ^ new_n397;
  assign new_n445 = new_n444 ^ n11;
  assign new_n446 = ~n65 & ~new_n445;
  assign new_n447 = new_n446 ^ new_n442;
  assign new_n448 = new_n447 ^ new_n438;
  assign new_n449 = n68 & new_n354;
  assign new_n450 = ~new_n304 & new_n349;
  assign new_n451 = new_n450 ^ new_n449;
  assign new_n452 = n69 & new_n348;
  assign new_n453 = n67 & new_n391;
  assign new_n454 = new_n453 ^ new_n452;
  assign new_n455 = new_n454 ^ new_n451;
  assign new_n456 = new_n455 ^ n9;
  assign new_n457 = new_n456 ^ new_n448;
  assign new_n458 = n71 & new_n218;
  assign new_n459 = new_n318 ^ n72;
  assign new_n460 = ~new_n459 & new_n208;
  assign new_n461 = new_n460 ^ new_n458;
  assign new_n462 = n72 & new_n207;
  assign new_n463 = n70 & new_n212;
  assign new_n464 = new_n463 ^ new_n462;
  assign new_n465 = new_n464 ^ new_n461;
  assign new_n466 = new_n465 ^ n6;
  assign new_n467 = new_n466 ^ new_n457;
  assign new_n468 = new_n413 ^ new_n400;
  assign new_n469 = ~new_n410 & new_n468;
  assign new_n470 = new_n469 ^ new_n413;
  assign new_n471 = new_n470 ^ new_n467;
  assign new_n472 = ~n74 & n73;
  assign new_n473 = ~new_n423 & new_n472;
  assign new_n474 = new_n424 ^ n73;
  assign new_n475 = n74 & new_n474;
  assign new_n476 = new_n475 ^ n74;
  assign new_n477 = new_n476 ^ new_n473;
  assign new_n478 = ~new_n477 & new_n155;
  assign new_n479 = new_n478 ^ n2;
  assign new_n480 = new_n479 ^ n75;
  assign new_n481 = n74 ^ n3;
  assign new_n482 = ~n73 & n3;
  assign new_n483 = new_n482 ^ new_n481;
  assign new_n484 = ~n2 & new_n483;
  assign new_n485 = new_n484 ^ new_n481;
  assign new_n486 = new_n485 ^ new_n480;
  assign new_n487 = ~n1 & new_n486;
  assign new_n488 = new_n487 ^ new_n480;
  assign new_n489 = new_n488 ^ new_n471;
  assign new_n490 = new_n435 ^ new_n414;
  assign new_n491 = ~new_n432 & new_n490;
  assign new_n492 = new_n491 ^ new_n435;
  assign new_n493 = new_n492 ^ new_n489;
  assign new_n494 = ~new_n398 & ~new_n447;
  assign new_n495 = n12 & new_n494;
  assign new_n496 = ~new_n444 & n11;
  assign new_n497 = new_n496 ^ new_n397;
  assign new_n498 = ~n11 & ~new_n397;
  assign new_n499 = new_n498 ^ new_n443;
  assign new_n500 = new_n499 ^ new_n497;
  assign new_n501 = ~new_n500 & n65;
  assign new_n502 = ~new_n397 & n12;
  assign new_n503 = n12 ^ n11;
  assign new_n504 = new_n503 ^ new_n498;
  assign new_n505 = new_n504 ^ new_n502;
  assign new_n506 = new_n505 ^ new_n397;
  assign new_n507 = ~new_n151 & ~new_n506;
  assign new_n508 = n67 & new_n397;
  assign new_n509 = new_n508 ^ new_n507;
  assign new_n510 = n66 & new_n499;
  assign new_n511 = new_n510 ^ new_n509;
  assign new_n512 = new_n511 ^ new_n501;
  assign new_n513 = new_n499 ^ new_n397;
  assign new_n514 = ~n12 & new_n513;
  assign new_n515 = new_n514 ^ n12;
  assign new_n516 = ~new_n515 & n65;
  assign new_n517 = new_n516 ^ n12;
  assign new_n518 = new_n517 ^ new_n512;
  assign new_n519 = new_n518 ^ new_n495;
  assign new_n520 = n69 & new_n354;
  assign new_n521 = ~new_n339 & new_n349;
  assign new_n522 = new_n521 ^ new_n520;
  assign new_n523 = n70 & new_n348;
  assign new_n524 = n68 & new_n391;
  assign new_n525 = new_n524 ^ new_n523;
  assign new_n526 = new_n525 ^ new_n522;
  assign new_n527 = new_n526 ^ n9;
  assign new_n528 = new_n527 ^ new_n519;
  assign new_n529 = new_n456 ^ new_n447;
  assign new_n530 = ~new_n529 & new_n448;
  assign new_n531 = new_n530 ^ new_n438;
  assign new_n532 = new_n531 ^ new_n528;
  assign new_n533 = n72 & new_n218;
  assign new_n534 = new_n372 ^ n73;
  assign new_n535 = new_n208 & new_n534;
  assign new_n536 = new_n535 ^ new_n533;
  assign new_n537 = n73 & new_n207;
  assign new_n538 = n71 & new_n212;
  assign new_n539 = new_n538 ^ new_n537;
  assign new_n540 = new_n539 ^ new_n536;
  assign new_n541 = new_n540 ^ n6;
  assign new_n542 = new_n541 ^ new_n532;
  assign new_n543 = new_n470 ^ new_n457;
  assign new_n544 = ~new_n467 & new_n543;
  assign new_n545 = new_n544 ^ new_n470;
  assign new_n546 = new_n545 ^ new_n542;
  assign new_n547 = n74 & new_n180;
  assign new_n548 = n2 & n75;
  assign new_n549 = new_n548 ^ new_n547;
  assign new_n550 = new_n549 ^ n3;
  assign new_n551 = new_n473 ^ n74;
  assign new_n552 = n75 & new_n551;
  assign new_n553 = ~n75 & ~new_n475;
  assign new_n554 = new_n553 ^ new_n552;
  assign new_n555 = new_n155 & new_n554;
  assign new_n556 = new_n555 ^ n2;
  assign new_n557 = new_n556 ^ n76;
  assign new_n558 = new_n557 ^ new_n550;
  assign new_n559 = ~n1 & new_n558;
  assign new_n560 = new_n559 ^ new_n557;
  assign new_n561 = new_n560 ^ new_n546;
  assign new_n562 = new_n492 ^ new_n471;
  assign new_n563 = ~new_n489 & new_n562;
  assign new_n564 = new_n563 ^ new_n492;
  assign new_n565 = new_n564 ^ new_n561;
  assign new_n566 = n70 & new_n354;
  assign new_n567 = ~new_n402 & new_n349;
  assign new_n568 = new_n567 ^ new_n566;
  assign new_n569 = n71 & new_n348;
  assign new_n570 = n69 & new_n391;
  assign new_n571 = new_n570 ^ new_n569;
  assign new_n572 = new_n571 ^ new_n568;
  assign new_n573 = new_n572 ^ n9;
  assign new_n574 = ~new_n259 & ~new_n506;
  assign new_n575 = n67 & new_n499;
  assign new_n576 = new_n575 ^ new_n574;
  assign new_n577 = ~new_n505 & n68;
  assign new_n578 = new_n502 ^ new_n444;
  assign new_n579 = ~new_n578 & new_n503;
  assign new_n580 = n66 & new_n579;
  assign new_n581 = new_n580 ^ new_n577;
  assign new_n582 = new_n581 ^ new_n576;
  assign new_n583 = new_n582 ^ n12;
  assign new_n584 = n13 ^ n12;
  assign new_n585 = n65 & new_n584;
  assign new_n586 = new_n585 ^ new_n583;
  assign new_n587 = ~new_n512 & new_n495;
  assign new_n588 = new_n587 ^ new_n586;
  assign new_n589 = new_n588 ^ new_n573;
  assign new_n590 = new_n531 ^ new_n519;
  assign new_n591 = ~new_n528 & new_n590;
  assign new_n592 = new_n591 ^ new_n531;
  assign new_n593 = new_n592 ^ new_n589;
  assign new_n594 = n73 & new_n218;
  assign new_n595 = new_n425 ^ n74;
  assign new_n596 = new_n208 & new_n595;
  assign new_n597 = new_n596 ^ new_n594;
  assign new_n598 = n74 & new_n207;
  assign new_n599 = n72 & new_n212;
  assign new_n600 = new_n599 ^ new_n598;
  assign new_n601 = new_n600 ^ new_n597;
  assign new_n602 = new_n601 ^ n6;
  assign new_n603 = new_n602 ^ new_n593;
  assign new_n604 = new_n545 ^ new_n532;
  assign new_n605 = ~new_n542 & new_n604;
  assign new_n606 = new_n605 ^ new_n545;
  assign new_n607 = new_n606 ^ new_n603;
  assign new_n608 = ~n76 & ~new_n552;
  assign new_n609 = ~new_n553 & n76;
  assign new_n610 = new_n609 ^ new_n608;
  assign new_n611 = new_n155 & new_n610;
  assign new_n612 = new_n611 ^ n2;
  assign new_n613 = new_n612 ^ n77;
  assign new_n614 = n76 ^ n3;
  assign new_n615 = ~n75 & n3;
  assign new_n616 = new_n615 ^ new_n614;
  assign new_n617 = ~n2 & new_n616;
  assign new_n618 = new_n617 ^ new_n614;
  assign new_n619 = new_n618 ^ new_n613;
  assign new_n620 = ~n1 & new_n619;
  assign new_n621 = new_n620 ^ new_n613;
  assign new_n622 = new_n621 ^ new_n607;
  assign new_n623 = new_n564 ^ new_n546;
  assign new_n624 = ~new_n561 & new_n623;
  assign new_n625 = new_n624 ^ new_n564;
  assign new_n626 = new_n625 ^ new_n622;
  assign new_n627 = ~new_n585 & ~new_n587;
  assign new_n628 = ~new_n627 & new_n583;
  assign new_n629 = n66 ^ n13;
  assign new_n630 = ~new_n629 & new_n584;
  assign new_n631 = new_n630 ^ n12;
  assign new_n632 = new_n631 ^ n14;
  assign new_n633 = n65 & new_n632;
  assign new_n634 = ~new_n151 & new_n584;
  assign new_n635 = ~new_n633 & ~new_n634;
  assign new_n636 = new_n635 ^ new_n628;
  assign new_n637 = n68 & new_n499;
  assign new_n638 = ~new_n304 & ~new_n506;
  assign new_n639 = new_n638 ^ new_n637;
  assign new_n640 = ~new_n505 & n69;
  assign new_n641 = n67 & new_n579;
  assign new_n642 = new_n641 ^ new_n640;
  assign new_n643 = new_n642 ^ new_n639;
  assign new_n644 = new_n643 ^ n12;
  assign new_n645 = new_n644 ^ new_n636;
  assign new_n646 = n71 & new_n354;
  assign new_n647 = ~new_n459 & new_n349;
  assign new_n648 = new_n647 ^ new_n646;
  assign new_n649 = n72 & new_n348;
  assign new_n650 = n70 & new_n391;
  assign new_n651 = new_n650 ^ new_n649;
  assign new_n652 = new_n651 ^ new_n648;
  assign new_n653 = new_n652 ^ n9;
  assign new_n654 = new_n653 ^ new_n645;
  assign new_n655 = new_n592 ^ new_n573;
  assign new_n656 = ~new_n589 & new_n655;
  assign new_n657 = new_n656 ^ new_n592;
  assign new_n658 = new_n657 ^ new_n654;
  assign new_n659 = n74 & new_n218;
  assign new_n660 = new_n477 ^ n75;
  assign new_n661 = new_n208 & new_n660;
  assign new_n662 = new_n661 ^ new_n659;
  assign new_n663 = n73 & new_n212;
  assign new_n664 = n75 & new_n207;
  assign new_n665 = new_n664 ^ new_n663;
  assign new_n666 = new_n665 ^ new_n662;
  assign new_n667 = new_n666 ^ n6;
  assign new_n668 = new_n667 ^ new_n658;
  assign new_n669 = new_n606 ^ new_n593;
  assign new_n670 = ~new_n603 & new_n669;
  assign new_n671 = new_n670 ^ new_n606;
  assign new_n672 = new_n671 ^ new_n668;
  assign new_n673 = n76 & new_n180;
  assign new_n674 = n2 & n77;
  assign new_n675 = new_n674 ^ new_n673;
  assign new_n676 = new_n675 ^ n3;
  assign new_n677 = ~new_n608 & n77;
  assign new_n678 = ~n77 & ~new_n609;
  assign new_n679 = new_n678 ^ new_n677;
  assign new_n680 = new_n155 & new_n679;
  assign new_n681 = new_n680 ^ n2;
  assign new_n682 = new_n681 ^ n78;
  assign new_n683 = new_n682 ^ new_n676;
  assign new_n684 = ~n1 & new_n683;
  assign new_n685 = new_n684 ^ new_n682;
  assign new_n686 = new_n685 ^ new_n672;
  assign new_n687 = new_n625 ^ new_n607;
  assign new_n688 = ~new_n622 & new_n687;
  assign new_n689 = new_n688 ^ new_n625;
  assign new_n690 = new_n689 ^ new_n686;
  assign new_n691 = n69 & new_n499;
  assign new_n692 = ~new_n339 & ~new_n506;
  assign new_n693 = new_n692 ^ new_n691;
  assign new_n694 = ~new_n505 & n70;
  assign new_n695 = n68 & new_n579;
  assign new_n696 = new_n695 ^ new_n694;
  assign new_n697 = new_n696 ^ new_n693;
  assign new_n698 = new_n697 ^ n12;
  assign new_n699 = n15 ^ n14;
  assign new_n700 = ~new_n699 & new_n584;
  assign new_n701 = new_n700 ^ new_n584;
  assign new_n702 = ~new_n151 & new_n701;
  assign new_n703 = n67 & new_n584;
  assign new_n704 = new_n703 ^ new_n702;
  assign new_n705 = ~new_n584 & n14;
  assign new_n706 = n12 & n13;
  assign new_n707 = new_n706 ^ new_n705;
  assign new_n708 = n66 & new_n707;
  assign new_n709 = new_n708 ^ new_n704;
  assign new_n710 = n14 & new_n706;
  assign new_n711 = n65 & new_n710;
  assign new_n712 = new_n711 ^ n65;
  assign new_n713 = new_n712 ^ new_n634;
  assign new_n714 = new_n713 ^ new_n711;
  assign new_n715 = n15 & new_n714;
  assign new_n716 = new_n715 ^ new_n711;
  assign new_n717 = new_n716 ^ new_n709;
  assign new_n718 = new_n717 ^ new_n698;
  assign new_n719 = new_n644 ^ new_n635;
  assign new_n720 = ~new_n636 & new_n719;
  assign new_n721 = new_n720 ^ new_n628;
  assign new_n722 = new_n721 ^ new_n718;
  assign new_n723 = n72 & new_n354;
  assign new_n724 = new_n349 & new_n534;
  assign new_n725 = new_n724 ^ new_n723;
  assign new_n726 = n73 & new_n348;
  assign new_n727 = n71 & new_n391;
  assign new_n728 = new_n727 ^ new_n726;
  assign new_n729 = new_n728 ^ new_n725;
  assign new_n730 = new_n729 ^ n9;
  assign new_n731 = new_n730 ^ new_n722;
  assign new_n732 = new_n657 ^ new_n645;
  assign new_n733 = ~new_n732 & new_n654;
  assign new_n734 = new_n733 ^ new_n657;
  assign new_n735 = new_n734 ^ new_n731;
  assign new_n736 = n75 & new_n218;
  assign new_n737 = new_n554 ^ n76;
  assign new_n738 = ~new_n737 & new_n208;
  assign new_n739 = new_n738 ^ new_n736;
  assign new_n740 = n76 & new_n207;
  assign new_n741 = n74 & new_n212;
  assign new_n742 = new_n741 ^ new_n740;
  assign new_n743 = new_n742 ^ new_n739;
  assign new_n744 = new_n743 ^ n6;
  assign new_n745 = new_n744 ^ new_n735;
  assign new_n746 = new_n671 ^ new_n658;
  assign new_n747 = ~new_n746 & new_n668;
  assign new_n748 = new_n747 ^ new_n671;
  assign new_n749 = new_n748 ^ new_n745;
  assign new_n750 = n77 & new_n180;
  assign new_n751 = n2 & n78;
  assign new_n752 = new_n751 ^ new_n750;
  assign new_n753 = new_n752 ^ n3;
  assign new_n754 = ~n78 & ~new_n677;
  assign new_n755 = ~new_n678 & n78;
  assign new_n756 = new_n755 ^ new_n754;
  assign new_n757 = new_n155 & new_n756;
  assign new_n758 = new_n757 ^ n2;
  assign new_n759 = new_n758 ^ n79;
  assign new_n760 = new_n759 ^ new_n753;
  assign new_n761 = ~n1 & new_n760;
  assign new_n762 = new_n761 ^ new_n759;
  assign new_n763 = new_n762 ^ new_n749;
  assign new_n764 = new_n689 ^ new_n672;
  assign new_n765 = ~new_n764 & new_n686;
  assign new_n766 = new_n765 ^ new_n689;
  assign new_n767 = new_n766 ^ new_n763;
  assign new_n768 = n70 & new_n499;
  assign new_n769 = ~new_n402 & ~new_n506;
  assign new_n770 = new_n769 ^ new_n768;
  assign new_n771 = ~new_n505 & n71;
  assign new_n772 = n69 & new_n579;
  assign new_n773 = new_n772 ^ new_n771;
  assign new_n774 = new_n773 ^ new_n770;
  assign new_n775 = new_n774 ^ n12;
  assign new_n776 = ~new_n713 & n15;
  assign new_n777 = ~new_n709 & new_n776;
  assign new_n778 = n16 ^ n15;
  assign new_n779 = n65 & new_n778;
  assign new_n780 = new_n779 ^ new_n777;
  assign new_n781 = ~new_n259 & new_n701;
  assign new_n782 = n67 & new_n707;
  assign new_n783 = new_n782 ^ new_n781;
  assign new_n784 = n68 & new_n700;
  assign new_n785 = ~new_n584 & n15;
  assign new_n786 = new_n785 ^ new_n706;
  assign new_n787 = new_n699 & new_n786;
  assign new_n788 = n66 & new_n787;
  assign new_n789 = new_n788 ^ new_n784;
  assign new_n790 = new_n789 ^ new_n783;
  assign new_n791 = new_n790 ^ n15;
  assign new_n792 = new_n791 ^ new_n780;
  assign new_n793 = new_n792 ^ new_n775;
  assign new_n794 = new_n721 ^ new_n698;
  assign new_n795 = ~new_n718 & new_n794;
  assign new_n796 = new_n795 ^ new_n721;
  assign new_n797 = new_n796 ^ new_n793;
  assign new_n798 = n73 & new_n354;
  assign new_n799 = new_n349 & new_n595;
  assign new_n800 = new_n799 ^ new_n798;
  assign new_n801 = n74 & new_n348;
  assign new_n802 = n72 & new_n391;
  assign new_n803 = new_n802 ^ new_n801;
  assign new_n804 = new_n803 ^ new_n800;
  assign new_n805 = new_n804 ^ n9;
  assign new_n806 = new_n805 ^ new_n797;
  assign new_n807 = new_n734 ^ new_n722;
  assign new_n808 = ~new_n731 & new_n807;
  assign new_n809 = new_n808 ^ new_n734;
  assign new_n810 = new_n809 ^ new_n806;
  assign new_n811 = n76 & new_n218;
  assign new_n812 = new_n610 ^ n77;
  assign new_n813 = ~new_n812 & new_n208;
  assign new_n814 = new_n813 ^ new_n811;
  assign new_n815 = n77 & new_n207;
  assign new_n816 = n75 & new_n212;
  assign new_n817 = new_n816 ^ new_n815;
  assign new_n818 = new_n817 ^ new_n814;
  assign new_n819 = new_n818 ^ n6;
  assign new_n820 = new_n819 ^ new_n810;
  assign new_n821 = new_n748 ^ new_n735;
  assign new_n822 = ~new_n745 & new_n821;
  assign new_n823 = new_n822 ^ new_n748;
  assign new_n824 = new_n823 ^ new_n820;
  assign new_n825 = n79 ^ n78;
  assign new_n826 = new_n756 & new_n825;
  assign new_n827 = ~new_n826 & new_n155;
  assign new_n828 = new_n827 ^ n2;
  assign new_n829 = new_n828 ^ n80;
  assign new_n830 = n79 ^ n3;
  assign new_n831 = ~n78 & n3;
  assign new_n832 = new_n831 ^ new_n830;
  assign new_n833 = ~n2 & new_n832;
  assign new_n834 = new_n833 ^ new_n830;
  assign new_n835 = new_n834 ^ new_n829;
  assign new_n836 = ~n1 & new_n835;
  assign new_n837 = new_n836 ^ new_n829;
  assign new_n838 = new_n837 ^ new_n824;
  assign new_n839 = new_n766 ^ new_n749;
  assign new_n840 = ~new_n763 & new_n839;
  assign new_n841 = new_n840 ^ new_n766;
  assign new_n842 = new_n841 ^ new_n838;
  assign new_n843 = ~n15 & ~n16;
  assign new_n844 = new_n843 ^ new_n778;
  assign new_n845 = new_n844 ^ n17;
  assign new_n846 = ~n65 & ~new_n845;
  assign new_n847 = n66 ^ n16;
  assign new_n848 = ~new_n847 & new_n778;
  assign new_n849 = new_n848 ^ n15;
  assign new_n850 = new_n849 ^ n17;
  assign new_n851 = new_n850 ^ new_n846;
  assign new_n852 = ~new_n777 & ~new_n779;
  assign new_n853 = ~new_n852 & new_n791;
  assign new_n854 = new_n853 ^ new_n851;
  assign new_n855 = n68 & new_n707;
  assign new_n856 = ~new_n304 & new_n701;
  assign new_n857 = new_n856 ^ new_n855;
  assign new_n858 = n69 & new_n700;
  assign new_n859 = n67 & new_n787;
  assign new_n860 = new_n859 ^ new_n858;
  assign new_n861 = new_n860 ^ new_n857;
  assign new_n862 = new_n861 ^ n15;
  assign new_n863 = new_n862 ^ new_n854;
  assign new_n864 = n71 & new_n499;
  assign new_n865 = ~new_n459 & ~new_n506;
  assign new_n866 = new_n865 ^ new_n864;
  assign new_n867 = ~new_n505 & n72;
  assign new_n868 = n70 & new_n579;
  assign new_n869 = new_n868 ^ new_n867;
  assign new_n870 = new_n869 ^ new_n866;
  assign new_n871 = new_n870 ^ n12;
  assign new_n872 = new_n871 ^ new_n863;
  assign new_n873 = new_n796 ^ new_n775;
  assign new_n874 = ~new_n793 & new_n873;
  assign new_n875 = new_n874 ^ new_n796;
  assign new_n876 = new_n875 ^ new_n872;
  assign new_n877 = n74 & new_n354;
  assign new_n878 = new_n349 & new_n660;
  assign new_n879 = new_n878 ^ new_n877;
  assign new_n880 = n75 & new_n348;
  assign new_n881 = n73 & new_n391;
  assign new_n882 = new_n881 ^ new_n880;
  assign new_n883 = new_n882 ^ new_n879;
  assign new_n884 = new_n883 ^ n9;
  assign new_n885 = new_n884 ^ new_n876;
  assign new_n886 = new_n809 ^ new_n797;
  assign new_n887 = ~new_n806 & new_n886;
  assign new_n888 = new_n887 ^ new_n809;
  assign new_n889 = new_n888 ^ new_n885;
  assign new_n890 = n77 & new_n218;
  assign new_n891 = new_n679 ^ n78;
  assign new_n892 = ~new_n891 & new_n208;
  assign new_n893 = new_n892 ^ new_n890;
  assign new_n894 = n78 & new_n207;
  assign new_n895 = n76 & new_n212;
  assign new_n896 = new_n895 ^ new_n894;
  assign new_n897 = new_n896 ^ new_n893;
  assign new_n898 = new_n897 ^ n6;
  assign new_n899 = new_n898 ^ new_n889;
  assign new_n900 = new_n823 ^ new_n810;
  assign new_n901 = ~new_n820 & new_n900;
  assign new_n902 = new_n901 ^ new_n823;
  assign new_n903 = new_n902 ^ new_n899;
  assign new_n904 = n79 & new_n180;
  assign new_n905 = n2 & n80;
  assign new_n906 = new_n905 ^ new_n904;
  assign new_n907 = new_n906 ^ n3;
  assign new_n908 = n80 ^ n79;
  assign new_n909 = ~n80 & new_n756;
  assign new_n910 = new_n909 ^ new_n755;
  assign new_n911 = ~new_n910 & new_n908;
  assign new_n912 = ~new_n911 & new_n155;
  assign new_n913 = new_n912 ^ n2;
  assign new_n914 = new_n913 ^ n81;
  assign new_n915 = new_n914 ^ new_n907;
  assign new_n916 = ~n1 & new_n915;
  assign new_n917 = new_n916 ^ new_n914;
  assign new_n918 = new_n917 ^ new_n903;
  assign new_n919 = new_n841 ^ new_n824;
  assign new_n920 = ~new_n838 & new_n919;
  assign new_n921 = new_n920 ^ new_n841;
  assign new_n922 = new_n921 ^ new_n918;
  assign new_n923 = n18 ^ n17;
  assign new_n924 = ~new_n923 & new_n778;
  assign new_n925 = new_n924 ^ new_n778;
  assign new_n926 = ~new_n151 & new_n925;
  assign new_n927 = n67 & new_n778;
  assign new_n928 = new_n927 ^ new_n926;
  assign new_n929 = ~new_n778 & n17;
  assign new_n930 = new_n929 ^ new_n844;
  assign new_n931 = ~new_n930 & n66;
  assign new_n932 = new_n931 ^ new_n928;
  assign new_n933 = new_n932 ^ n18;
  assign new_n934 = ~new_n778 & n18;
  assign new_n935 = new_n934 ^ new_n844;
  assign new_n936 = ~new_n935 & new_n923;
  assign new_n937 = n65 & new_n936;
  assign new_n938 = new_n937 ^ new_n933;
  assign new_n939 = ~new_n779 & ~new_n851;
  assign new_n940 = n18 & new_n939;
  assign new_n941 = new_n940 ^ new_n938;
  assign new_n942 = n69 & new_n707;
  assign new_n943 = ~new_n339 & new_n701;
  assign new_n944 = new_n943 ^ new_n942;
  assign new_n945 = n70 & new_n700;
  assign new_n946 = n68 & new_n787;
  assign new_n947 = new_n946 ^ new_n945;
  assign new_n948 = new_n947 ^ new_n944;
  assign new_n949 = new_n948 ^ n15;
  assign new_n950 = new_n949 ^ new_n941;
  assign new_n951 = new_n862 ^ new_n851;
  assign new_n952 = ~new_n951 & new_n854;
  assign new_n953 = new_n952 ^ new_n853;
  assign new_n954 = new_n953 ^ new_n950;
  assign new_n955 = n72 & new_n499;
  assign new_n956 = ~new_n506 & new_n534;
  assign new_n957 = new_n956 ^ new_n955;
  assign new_n958 = ~new_n505 & n73;
  assign new_n959 = n71 & new_n579;
  assign new_n960 = new_n959 ^ new_n958;
  assign new_n961 = new_n960 ^ new_n957;
  assign new_n962 = new_n961 ^ n12;
  assign new_n963 = new_n962 ^ new_n954;
  assign new_n964 = new_n875 ^ new_n863;
  assign new_n965 = ~new_n872 & new_n964;
  assign new_n966 = new_n965 ^ new_n875;
  assign new_n967 = new_n966 ^ new_n963;
  assign new_n968 = n75 & new_n354;
  assign new_n969 = ~new_n737 & new_n349;
  assign new_n970 = new_n969 ^ new_n968;
  assign new_n971 = n76 & new_n348;
  assign new_n972 = n74 & new_n391;
  assign new_n973 = new_n972 ^ new_n971;
  assign new_n974 = new_n973 ^ new_n970;
  assign new_n975 = new_n974 ^ n9;
  assign new_n976 = new_n975 ^ new_n967;
  assign new_n977 = new_n888 ^ new_n876;
  assign new_n978 = ~new_n885 & new_n977;
  assign new_n979 = new_n978 ^ new_n888;
  assign new_n980 = new_n979 ^ new_n976;
  assign new_n981 = n78 & new_n218;
  assign new_n982 = new_n756 ^ n79;
  assign new_n983 = ~new_n982 & new_n208;
  assign new_n984 = new_n983 ^ new_n981;
  assign new_n985 = n79 & new_n207;
  assign new_n986 = n77 & new_n212;
  assign new_n987 = new_n986 ^ new_n985;
  assign new_n988 = new_n987 ^ new_n984;
  assign new_n989 = new_n988 ^ n6;
  assign new_n990 = new_n989 ^ new_n980;
  assign new_n991 = new_n902 ^ new_n889;
  assign new_n992 = ~new_n899 & new_n991;
  assign new_n993 = new_n992 ^ new_n902;
  assign new_n994 = new_n993 ^ new_n990;
  assign new_n995 = n81 ^ n80;
  assign new_n996 = ~new_n911 & new_n995;
  assign new_n997 = ~new_n996 & new_n155;
  assign new_n998 = new_n997 ^ n2;
  assign new_n999 = new_n998 ^ n82;
  assign new_n1000 = n81 ^ n3;
  assign new_n1001 = n80 ^ n3;
  assign new_n1002 = ~n80 & ~new_n1001;
  assign new_n1003 = new_n1002 ^ new_n1000;
  assign new_n1004 = new_n1003 ^ n80;
  assign new_n1005 = ~new_n1004 & new_n241;
  assign new_n1006 = new_n1005 ^ new_n1002;
  assign new_n1007 = new_n1006 ^ n80;
  assign new_n1008 = new_n1007 ^ new_n999;
  assign new_n1009 = ~n1 & ~new_n1008;
  assign new_n1010 = new_n1009 ^ new_n999;
  assign new_n1011 = new_n1010 ^ new_n994;
  assign new_n1012 = new_n921 ^ new_n903;
  assign new_n1013 = ~new_n918 & new_n1012;
  assign new_n1014 = new_n1013 ^ new_n921;
  assign new_n1015 = new_n1014 ^ new_n1011;
  assign new_n1016 = new_n938 & new_n940;
  assign new_n1017 = ~new_n259 & new_n925;
  assign new_n1018 = ~new_n930 & n67;
  assign new_n1019 = new_n1018 ^ new_n1017;
  assign new_n1020 = n68 & new_n924;
  assign new_n1021 = n66 & new_n936;
  assign new_n1022 = new_n1021 ^ new_n1020;
  assign new_n1023 = new_n1022 ^ new_n1019;
  assign new_n1024 = new_n1023 ^ n18;
  assign new_n1025 = n19 ^ n18;
  assign new_n1026 = n65 & new_n1025;
  assign new_n1027 = new_n1026 ^ new_n1024;
  assign new_n1028 = new_n1027 ^ new_n1016;
  assign new_n1029 = n70 & new_n707;
  assign new_n1030 = ~new_n402 & new_n701;
  assign new_n1031 = new_n1030 ^ new_n1029;
  assign new_n1032 = n71 & new_n700;
  assign new_n1033 = n69 & new_n787;
  assign new_n1034 = new_n1033 ^ new_n1032;
  assign new_n1035 = new_n1034 ^ new_n1031;
  assign new_n1036 = new_n1035 ^ n15;
  assign new_n1037 = new_n1036 ^ new_n1028;
  assign new_n1038 = new_n953 ^ new_n941;
  assign new_n1039 = ~new_n950 & new_n1038;
  assign new_n1040 = new_n1039 ^ new_n953;
  assign new_n1041 = new_n1040 ^ new_n1037;
  assign new_n1042 = n73 & new_n499;
  assign new_n1043 = ~new_n506 & new_n595;
  assign new_n1044 = new_n1043 ^ new_n1042;
  assign new_n1045 = ~new_n505 & n74;
  assign new_n1046 = n72 & new_n579;
  assign new_n1047 = new_n1046 ^ new_n1045;
  assign new_n1048 = new_n1047 ^ new_n1044;
  assign new_n1049 = new_n1048 ^ n12;
  assign new_n1050 = new_n1049 ^ new_n1041;
  assign new_n1051 = new_n966 ^ new_n954;
  assign new_n1052 = ~new_n963 & new_n1051;
  assign new_n1053 = new_n1052 ^ new_n966;
  assign new_n1054 = new_n1053 ^ new_n1050;
  assign new_n1055 = n76 & new_n354;
  assign new_n1056 = ~new_n812 & new_n349;
  assign new_n1057 = new_n1056 ^ new_n1055;
  assign new_n1058 = n77 & new_n348;
  assign new_n1059 = n75 & new_n391;
  assign new_n1060 = new_n1059 ^ new_n1058;
  assign new_n1061 = new_n1060 ^ new_n1057;
  assign new_n1062 = new_n1061 ^ n9;
  assign new_n1063 = new_n1062 ^ new_n1054;
  assign new_n1064 = new_n979 ^ new_n967;
  assign new_n1065 = ~new_n976 & new_n1064;
  assign new_n1066 = new_n1065 ^ new_n979;
  assign new_n1067 = new_n1066 ^ new_n1063;
  assign new_n1068 = n79 & new_n218;
  assign new_n1069 = new_n826 ^ n80;
  assign new_n1070 = new_n208 & new_n1069;
  assign new_n1071 = new_n1070 ^ new_n1068;
  assign new_n1072 = n80 & new_n207;
  assign new_n1073 = n78 & new_n212;
  assign new_n1074 = new_n1073 ^ new_n1072;
  assign new_n1075 = new_n1074 ^ new_n1071;
  assign new_n1076 = new_n1075 ^ n6;
  assign new_n1077 = new_n1076 ^ new_n1067;
  assign new_n1078 = new_n993 ^ new_n980;
  assign new_n1079 = ~new_n990 & new_n1078;
  assign new_n1080 = new_n1079 ^ new_n993;
  assign new_n1081 = new_n1080 ^ new_n1077;
  assign new_n1082 = n82 ^ n3;
  assign new_n1083 = ~n81 & n3;
  assign new_n1084 = new_n1083 ^ new_n1082;
  assign new_n1085 = ~n2 & new_n1084;
  assign new_n1086 = new_n1085 ^ new_n1082;
  assign new_n1087 = n82 ^ n81;
  assign new_n1088 = ~new_n996 & new_n1087;
  assign new_n1089 = ~new_n1088 & new_n155;
  assign new_n1090 = new_n1089 ^ n2;
  assign new_n1091 = new_n1090 ^ n83;
  assign new_n1092 = new_n1091 ^ new_n1086;
  assign new_n1093 = ~n1 & new_n1092;
  assign new_n1094 = new_n1093 ^ new_n1091;
  assign new_n1095 = new_n1094 ^ new_n1081;
  assign new_n1096 = new_n1014 ^ new_n994;
  assign new_n1097 = ~new_n1011 & new_n1096;
  assign new_n1098 = new_n1097 ^ new_n1014;
  assign new_n1099 = new_n1098 ^ new_n1095;
  assign new_n1100 = ~new_n1016 & ~new_n1026;
  assign new_n1101 = ~new_n1100 & new_n1024;
  assign new_n1102 = ~new_n930 & n68;
  assign new_n1103 = ~new_n304 & new_n925;
  assign new_n1104 = new_n1103 ^ new_n1102;
  assign new_n1105 = n69 & new_n924;
  assign new_n1106 = n67 & new_n936;
  assign new_n1107 = new_n1106 ^ new_n1105;
  assign new_n1108 = new_n1107 ^ new_n1104;
  assign new_n1109 = new_n1108 ^ n18;
  assign new_n1110 = n66 ^ n19;
  assign new_n1111 = ~new_n1110 & new_n1025;
  assign new_n1112 = new_n1111 ^ n18;
  assign new_n1113 = new_n1112 ^ n20;
  assign new_n1114 = ~n18 & ~n19;
  assign new_n1115 = new_n1114 ^ new_n1025;
  assign new_n1116 = new_n1115 ^ n20;
  assign new_n1117 = ~n65 & ~new_n1116;
  assign new_n1118 = new_n1117 ^ new_n1113;
  assign new_n1119 = new_n1118 ^ new_n1109;
  assign new_n1120 = new_n1119 ^ new_n1101;
  assign new_n1121 = n71 & new_n707;
  assign new_n1122 = ~new_n459 & new_n701;
  assign new_n1123 = new_n1122 ^ new_n1121;
  assign new_n1124 = n72 & new_n700;
  assign new_n1125 = n70 & new_n787;
  assign new_n1126 = new_n1125 ^ new_n1124;
  assign new_n1127 = new_n1126 ^ new_n1123;
  assign new_n1128 = new_n1127 ^ n15;
  assign new_n1129 = new_n1128 ^ new_n1120;
  assign new_n1130 = new_n1040 ^ new_n1028;
  assign new_n1131 = ~new_n1037 & new_n1130;
  assign new_n1132 = new_n1131 ^ new_n1040;
  assign new_n1133 = new_n1132 ^ new_n1129;
  assign new_n1134 = n74 & new_n499;
  assign new_n1135 = ~new_n506 & new_n660;
  assign new_n1136 = new_n1135 ^ new_n1134;
  assign new_n1137 = ~new_n505 & n75;
  assign new_n1138 = n73 & new_n579;
  assign new_n1139 = new_n1138 ^ new_n1137;
  assign new_n1140 = new_n1139 ^ new_n1136;
  assign new_n1141 = new_n1140 ^ n12;
  assign new_n1142 = new_n1141 ^ new_n1133;
  assign new_n1143 = new_n1053 ^ new_n1041;
  assign new_n1144 = ~new_n1050 & new_n1143;
  assign new_n1145 = new_n1144 ^ new_n1053;
  assign new_n1146 = new_n1145 ^ new_n1142;
  assign new_n1147 = n77 & new_n354;
  assign new_n1148 = ~new_n891 & new_n349;
  assign new_n1149 = new_n1148 ^ new_n1147;
  assign new_n1150 = n78 & new_n348;
  assign new_n1151 = n76 & new_n391;
  assign new_n1152 = new_n1151 ^ new_n1150;
  assign new_n1153 = new_n1152 ^ new_n1149;
  assign new_n1154 = new_n1153 ^ n9;
  assign new_n1155 = new_n1154 ^ new_n1146;
  assign new_n1156 = new_n1066 ^ new_n1054;
  assign new_n1157 = ~new_n1063 & new_n1156;
  assign new_n1158 = new_n1157 ^ new_n1066;
  assign new_n1159 = new_n1158 ^ new_n1155;
  assign new_n1160 = n80 & new_n218;
  assign new_n1161 = new_n911 ^ n81;
  assign new_n1162 = new_n208 & new_n1161;
  assign new_n1163 = new_n1162 ^ new_n1160;
  assign new_n1164 = n79 & new_n212;
  assign new_n1165 = n81 & new_n207;
  assign new_n1166 = new_n1165 ^ new_n1164;
  assign new_n1167 = new_n1166 ^ new_n1163;
  assign new_n1168 = new_n1167 ^ n6;
  assign new_n1169 = new_n1168 ^ new_n1159;
  assign new_n1170 = new_n1080 ^ new_n1067;
  assign new_n1171 = ~new_n1077 & new_n1170;
  assign new_n1172 = new_n1171 ^ new_n1080;
  assign new_n1173 = new_n1172 ^ new_n1169;
  assign new_n1174 = n82 & new_n180;
  assign new_n1175 = n2 & n83;
  assign new_n1176 = new_n1175 ^ new_n1174;
  assign new_n1177 = new_n1176 ^ n3;
  assign new_n1178 = n83 ^ n82;
  assign new_n1179 = ~new_n1088 & new_n1178;
  assign new_n1180 = ~new_n1179 & new_n155;
  assign new_n1181 = new_n1180 ^ n2;
  assign new_n1182 = new_n1181 ^ n84;
  assign new_n1183 = new_n1182 ^ new_n1177;
  assign new_n1184 = ~n1 & new_n1183;
  assign new_n1185 = new_n1184 ^ new_n1182;
  assign new_n1186 = new_n1185 ^ new_n1173;
  assign new_n1187 = new_n1098 ^ new_n1081;
  assign new_n1188 = ~new_n1095 & new_n1187;
  assign new_n1189 = new_n1188 ^ new_n1098;
  assign new_n1190 = new_n1189 ^ new_n1186;
  assign new_n1191 = n21 ^ n20;
  assign new_n1192 = ~new_n1191 & new_n1025;
  assign new_n1193 = new_n1192 ^ new_n1025;
  assign new_n1194 = ~new_n151 & new_n1193;
  assign new_n1195 = n67 & new_n1025;
  assign new_n1196 = new_n1195 ^ new_n1194;
  assign new_n1197 = ~new_n1025 & n20;
  assign new_n1198 = new_n1197 ^ new_n1115;
  assign new_n1199 = ~new_n1198 & n66;
  assign new_n1200 = new_n1199 ^ new_n1196;
  assign new_n1201 = new_n1200 ^ n21;
  assign new_n1202 = ~new_n1025 & n21;
  assign new_n1203 = new_n1202 ^ new_n1115;
  assign new_n1204 = ~new_n1203 & new_n1191;
  assign new_n1205 = n65 & new_n1204;
  assign new_n1206 = new_n1205 ^ new_n1201;
  assign new_n1207 = ~new_n1026 & ~new_n1118;
  assign new_n1208 = n21 & new_n1207;
  assign new_n1209 = new_n1208 ^ new_n1206;
  assign new_n1210 = ~new_n930 & n69;
  assign new_n1211 = ~new_n339 & new_n925;
  assign new_n1212 = new_n1211 ^ new_n1210;
  assign new_n1213 = n70 & new_n924;
  assign new_n1214 = n68 & new_n936;
  assign new_n1215 = new_n1214 ^ new_n1213;
  assign new_n1216 = new_n1215 ^ new_n1212;
  assign new_n1217 = new_n1216 ^ n18;
  assign new_n1218 = new_n1217 ^ new_n1209;
  assign new_n1219 = new_n1109 ^ new_n1101;
  assign new_n1220 = ~new_n1119 & new_n1219;
  assign new_n1221 = new_n1220 ^ new_n1101;
  assign new_n1222 = new_n1221 ^ new_n1218;
  assign new_n1223 = n72 & new_n707;
  assign new_n1224 = new_n534 & new_n701;
  assign new_n1225 = new_n1224 ^ new_n1223;
  assign new_n1226 = n73 & new_n700;
  assign new_n1227 = n71 & new_n787;
  assign new_n1228 = new_n1227 ^ new_n1226;
  assign new_n1229 = new_n1228 ^ new_n1225;
  assign new_n1230 = new_n1229 ^ n15;
  assign new_n1231 = new_n1230 ^ new_n1222;
  assign new_n1232 = new_n1132 ^ new_n1120;
  assign new_n1233 = ~new_n1129 & new_n1232;
  assign new_n1234 = new_n1233 ^ new_n1132;
  assign new_n1235 = new_n1234 ^ new_n1231;
  assign new_n1236 = n75 & new_n499;
  assign new_n1237 = ~new_n506 & ~new_n737;
  assign new_n1238 = new_n1237 ^ new_n1236;
  assign new_n1239 = ~new_n505 & n76;
  assign new_n1240 = n74 & new_n579;
  assign new_n1241 = new_n1240 ^ new_n1239;
  assign new_n1242 = new_n1241 ^ new_n1238;
  assign new_n1243 = new_n1242 ^ n12;
  assign new_n1244 = new_n1243 ^ new_n1235;
  assign new_n1245 = new_n1145 ^ new_n1133;
  assign new_n1246 = ~new_n1142 & new_n1245;
  assign new_n1247 = new_n1246 ^ new_n1145;
  assign new_n1248 = new_n1247 ^ new_n1244;
  assign new_n1249 = n78 & new_n354;
  assign new_n1250 = ~new_n982 & new_n349;
  assign new_n1251 = new_n1250 ^ new_n1249;
  assign new_n1252 = n79 & new_n348;
  assign new_n1253 = n77 & new_n391;
  assign new_n1254 = new_n1253 ^ new_n1252;
  assign new_n1255 = new_n1254 ^ new_n1251;
  assign new_n1256 = new_n1255 ^ n9;
  assign new_n1257 = new_n1256 ^ new_n1248;
  assign new_n1258 = new_n1158 ^ new_n1146;
  assign new_n1259 = ~new_n1155 & new_n1258;
  assign new_n1260 = new_n1259 ^ new_n1158;
  assign new_n1261 = new_n1260 ^ new_n1257;
  assign new_n1262 = n81 & new_n218;
  assign new_n1263 = new_n996 ^ n82;
  assign new_n1264 = new_n208 & new_n1263;
  assign new_n1265 = new_n1264 ^ new_n1262;
  assign new_n1266 = n82 & new_n207;
  assign new_n1267 = n80 & new_n212;
  assign new_n1268 = new_n1267 ^ new_n1266;
  assign new_n1269 = new_n1268 ^ new_n1265;
  assign new_n1270 = new_n1269 ^ n6;
  assign new_n1271 = new_n1270 ^ new_n1261;
  assign new_n1272 = new_n1172 ^ new_n1159;
  assign new_n1273 = ~new_n1169 & new_n1272;
  assign new_n1274 = new_n1273 ^ new_n1172;
  assign new_n1275 = new_n1274 ^ new_n1271;
  assign new_n1276 = n84 ^ n83;
  assign new_n1277 = ~new_n1179 & new_n1276;
  assign new_n1278 = ~new_n1277 & new_n155;
  assign new_n1279 = new_n1278 ^ n2;
  assign new_n1280 = new_n1279 ^ n85;
  assign new_n1281 = n84 ^ n3;
  assign new_n1282 = n83 ^ n3;
  assign new_n1283 = ~n83 & ~new_n1282;
  assign new_n1284 = new_n1283 ^ new_n1281;
  assign new_n1285 = new_n1284 ^ n83;
  assign new_n1286 = ~new_n1285 & new_n241;
  assign new_n1287 = new_n1286 ^ new_n1283;
  assign new_n1288 = new_n1287 ^ n83;
  assign new_n1289 = new_n1288 ^ new_n1280;
  assign new_n1290 = ~n1 & ~new_n1289;
  assign new_n1291 = new_n1290 ^ new_n1280;
  assign new_n1292 = new_n1291 ^ new_n1275;
  assign new_n1293 = new_n1189 ^ new_n1173;
  assign new_n1294 = ~new_n1186 & new_n1293;
  assign new_n1295 = new_n1294 ^ new_n1189;
  assign new_n1296 = new_n1295 ^ new_n1292;
  assign new_n1297 = new_n1206 & new_n1208;
  assign new_n1298 = ~new_n259 & new_n1193;
  assign new_n1299 = ~new_n1198 & n67;
  assign new_n1300 = new_n1299 ^ new_n1298;
  assign new_n1301 = n68 & new_n1192;
  assign new_n1302 = n66 & new_n1204;
  assign new_n1303 = new_n1302 ^ new_n1301;
  assign new_n1304 = new_n1303 ^ new_n1300;
  assign new_n1305 = new_n1304 ^ n21;
  assign new_n1306 = n22 ^ n21;
  assign new_n1307 = n65 & new_n1306;
  assign new_n1308 = new_n1307 ^ new_n1305;
  assign new_n1309 = new_n1308 ^ new_n1297;
  assign new_n1310 = ~new_n930 & n70;
  assign new_n1311 = ~new_n402 & new_n925;
  assign new_n1312 = new_n1311 ^ new_n1310;
  assign new_n1313 = n71 & new_n924;
  assign new_n1314 = n69 & new_n936;
  assign new_n1315 = new_n1314 ^ new_n1313;
  assign new_n1316 = new_n1315 ^ new_n1312;
  assign new_n1317 = new_n1316 ^ n18;
  assign new_n1318 = new_n1317 ^ new_n1309;
  assign new_n1319 = new_n1221 ^ new_n1209;
  assign new_n1320 = ~new_n1218 & new_n1319;
  assign new_n1321 = new_n1320 ^ new_n1221;
  assign new_n1322 = new_n1321 ^ new_n1318;
  assign new_n1323 = n73 & new_n707;
  assign new_n1324 = new_n595 & new_n701;
  assign new_n1325 = new_n1324 ^ new_n1323;
  assign new_n1326 = n74 & new_n700;
  assign new_n1327 = n72 & new_n787;
  assign new_n1328 = new_n1327 ^ new_n1326;
  assign new_n1329 = new_n1328 ^ new_n1325;
  assign new_n1330 = new_n1329 ^ n15;
  assign new_n1331 = new_n1330 ^ new_n1322;
  assign new_n1332 = new_n1234 ^ new_n1222;
  assign new_n1333 = ~new_n1231 & new_n1332;
  assign new_n1334 = new_n1333 ^ new_n1234;
  assign new_n1335 = new_n1334 ^ new_n1331;
  assign new_n1336 = n76 & new_n499;
  assign new_n1337 = ~new_n506 & ~new_n812;
  assign new_n1338 = new_n1337 ^ new_n1336;
  assign new_n1339 = n75 & new_n579;
  assign new_n1340 = ~new_n505 & n77;
  assign new_n1341 = new_n1340 ^ new_n1339;
  assign new_n1342 = new_n1341 ^ new_n1338;
  assign new_n1343 = new_n1342 ^ n12;
  assign new_n1344 = new_n1343 ^ new_n1335;
  assign new_n1345 = new_n1247 ^ new_n1235;
  assign new_n1346 = ~new_n1244 & new_n1345;
  assign new_n1347 = new_n1346 ^ new_n1247;
  assign new_n1348 = new_n1347 ^ new_n1344;
  assign new_n1349 = n79 & new_n354;
  assign new_n1350 = new_n349 & new_n1069;
  assign new_n1351 = new_n1350 ^ new_n1349;
  assign new_n1352 = n80 & new_n348;
  assign new_n1353 = n78 & new_n391;
  assign new_n1354 = new_n1353 ^ new_n1352;
  assign new_n1355 = new_n1354 ^ new_n1351;
  assign new_n1356 = new_n1355 ^ n9;
  assign new_n1357 = new_n1356 ^ new_n1348;
  assign new_n1358 = new_n1260 ^ new_n1248;
  assign new_n1359 = ~new_n1257 & new_n1358;
  assign new_n1360 = new_n1359 ^ new_n1260;
  assign new_n1361 = new_n1360 ^ new_n1357;
  assign new_n1362 = n82 & new_n218;
  assign new_n1363 = new_n1088 ^ n83;
  assign new_n1364 = new_n208 & new_n1363;
  assign new_n1365 = new_n1364 ^ new_n1362;
  assign new_n1366 = n83 & new_n207;
  assign new_n1367 = n81 & new_n212;
  assign new_n1368 = new_n1367 ^ new_n1366;
  assign new_n1369 = new_n1368 ^ new_n1365;
  assign new_n1370 = new_n1369 ^ n6;
  assign new_n1371 = new_n1370 ^ new_n1361;
  assign new_n1372 = new_n1274 ^ new_n1261;
  assign new_n1373 = ~new_n1271 & new_n1372;
  assign new_n1374 = new_n1373 ^ new_n1274;
  assign new_n1375 = new_n1374 ^ new_n1371;
  assign new_n1376 = n85 ^ n84;
  assign new_n1377 = ~new_n1277 & new_n1376;
  assign new_n1378 = ~new_n1377 & new_n155;
  assign new_n1379 = new_n1378 ^ n2;
  assign new_n1380 = new_n1379 ^ n86;
  assign new_n1381 = ~n84 & n3;
  assign new_n1382 = n85 ^ n3;
  assign new_n1383 = new_n1382 ^ new_n1381;
  assign new_n1384 = n2 & new_n1383;
  assign new_n1385 = new_n1384 ^ new_n1381;
  assign new_n1386 = new_n1385 ^ new_n1380;
  assign new_n1387 = ~n1 & new_n1386;
  assign new_n1388 = new_n1387 ^ new_n1380;
  assign new_n1389 = new_n1388 ^ new_n1375;
  assign new_n1390 = new_n1295 ^ new_n1275;
  assign new_n1391 = ~new_n1292 & new_n1390;
  assign new_n1392 = new_n1391 ^ new_n1295;
  assign new_n1393 = new_n1392 ^ new_n1389;
  assign new_n1394 = ~new_n1297 & ~new_n1307;
  assign new_n1395 = ~new_n1394 & new_n1305;
  assign new_n1396 = ~n21 & ~n22;
  assign new_n1397 = new_n1396 ^ new_n1306;
  assign new_n1398 = new_n1397 ^ n23;
  assign new_n1399 = ~n65 & ~new_n1398;
  assign new_n1400 = n66 ^ n22;
  assign new_n1401 = ~new_n1400 & new_n1306;
  assign new_n1402 = new_n1401 ^ n21;
  assign new_n1403 = new_n1402 ^ n23;
  assign new_n1404 = new_n1403 ^ new_n1399;
  assign new_n1405 = ~new_n1198 & n68;
  assign new_n1406 = ~new_n304 & new_n1193;
  assign new_n1407 = new_n1406 ^ new_n1405;
  assign new_n1408 = n69 & new_n1192;
  assign new_n1409 = n67 & new_n1204;
  assign new_n1410 = new_n1409 ^ new_n1408;
  assign new_n1411 = new_n1410 ^ new_n1407;
  assign new_n1412 = new_n1411 ^ n21;
  assign new_n1413 = new_n1412 ^ new_n1404;
  assign new_n1414 = new_n1413 ^ new_n1395;
  assign new_n1415 = ~new_n930 & n71;
  assign new_n1416 = ~new_n459 & new_n925;
  assign new_n1417 = new_n1416 ^ new_n1415;
  assign new_n1418 = n72 & new_n924;
  assign new_n1419 = n70 & new_n936;
  assign new_n1420 = new_n1419 ^ new_n1418;
  assign new_n1421 = new_n1420 ^ new_n1417;
  assign new_n1422 = new_n1421 ^ n18;
  assign new_n1423 = new_n1422 ^ new_n1414;
  assign new_n1424 = new_n1321 ^ new_n1309;
  assign new_n1425 = ~new_n1318 & new_n1424;
  assign new_n1426 = new_n1425 ^ new_n1321;
  assign new_n1427 = new_n1426 ^ new_n1423;
  assign new_n1428 = n74 & new_n707;
  assign new_n1429 = new_n660 & new_n701;
  assign new_n1430 = new_n1429 ^ new_n1428;
  assign new_n1431 = n75 & new_n700;
  assign new_n1432 = n73 & new_n787;
  assign new_n1433 = new_n1432 ^ new_n1431;
  assign new_n1434 = new_n1433 ^ new_n1430;
  assign new_n1435 = new_n1434 ^ n15;
  assign new_n1436 = new_n1435 ^ new_n1427;
  assign new_n1437 = new_n1334 ^ new_n1322;
  assign new_n1438 = ~new_n1331 & new_n1437;
  assign new_n1439 = new_n1438 ^ new_n1334;
  assign new_n1440 = new_n1439 ^ new_n1436;
  assign new_n1441 = n77 & new_n499;
  assign new_n1442 = ~new_n506 & ~new_n891;
  assign new_n1443 = new_n1442 ^ new_n1441;
  assign new_n1444 = ~new_n505 & n78;
  assign new_n1445 = n76 & new_n579;
  assign new_n1446 = new_n1445 ^ new_n1444;
  assign new_n1447 = new_n1446 ^ new_n1443;
  assign new_n1448 = new_n1447 ^ n12;
  assign new_n1449 = new_n1448 ^ new_n1440;
  assign new_n1450 = new_n1347 ^ new_n1335;
  assign new_n1451 = ~new_n1344 & new_n1450;
  assign new_n1452 = new_n1451 ^ new_n1347;
  assign new_n1453 = new_n1452 ^ new_n1449;
  assign new_n1454 = n80 & new_n354;
  assign new_n1455 = new_n349 & new_n1161;
  assign new_n1456 = new_n1455 ^ new_n1454;
  assign new_n1457 = n81 & new_n348;
  assign new_n1458 = n79 & new_n391;
  assign new_n1459 = new_n1458 ^ new_n1457;
  assign new_n1460 = new_n1459 ^ new_n1456;
  assign new_n1461 = new_n1460 ^ n9;
  assign new_n1462 = new_n1461 ^ new_n1453;
  assign new_n1463 = new_n1360 ^ new_n1348;
  assign new_n1464 = ~new_n1357 & new_n1463;
  assign new_n1465 = new_n1464 ^ new_n1360;
  assign new_n1466 = new_n1465 ^ new_n1462;
  assign new_n1467 = n83 & new_n218;
  assign new_n1468 = new_n1179 ^ n84;
  assign new_n1469 = new_n208 & new_n1468;
  assign new_n1470 = new_n1469 ^ new_n1467;
  assign new_n1471 = n84 & new_n207;
  assign new_n1472 = n82 & new_n212;
  assign new_n1473 = new_n1472 ^ new_n1471;
  assign new_n1474 = new_n1473 ^ new_n1470;
  assign new_n1475 = new_n1474 ^ n6;
  assign new_n1476 = new_n1475 ^ new_n1466;
  assign new_n1477 = new_n1374 ^ new_n1361;
  assign new_n1478 = ~new_n1371 & new_n1477;
  assign new_n1479 = new_n1478 ^ new_n1374;
  assign new_n1480 = new_n1479 ^ new_n1476;
  assign new_n1481 = n86 ^ n85;
  assign new_n1482 = ~new_n1377 & new_n1481;
  assign new_n1483 = ~new_n1482 & new_n155;
  assign new_n1484 = new_n1483 ^ n2;
  assign new_n1485 = new_n1484 ^ n87;
  assign new_n1486 = n86 ^ n3;
  assign new_n1487 = ~n85 & n3;
  assign new_n1488 = new_n1487 ^ new_n1486;
  assign new_n1489 = ~n2 & new_n1488;
  assign new_n1490 = new_n1489 ^ new_n1486;
  assign new_n1491 = new_n1490 ^ new_n1485;
  assign new_n1492 = ~n1 & new_n1491;
  assign new_n1493 = new_n1492 ^ new_n1485;
  assign new_n1494 = new_n1493 ^ new_n1480;
  assign new_n1495 = new_n1392 ^ new_n1375;
  assign new_n1496 = ~new_n1389 & new_n1495;
  assign new_n1497 = new_n1496 ^ new_n1392;
  assign new_n1498 = new_n1497 ^ new_n1494;
  assign new_n1499 = n24 ^ n23;
  assign new_n1500 = ~new_n1499 & new_n1306;
  assign new_n1501 = new_n1500 ^ new_n1306;
  assign new_n1502 = ~new_n151 & new_n1501;
  assign new_n1503 = n67 & new_n1306;
  assign new_n1504 = new_n1503 ^ new_n1502;
  assign new_n1505 = ~new_n1306 & n23;
  assign new_n1506 = new_n1505 ^ new_n1397;
  assign new_n1507 = ~new_n1506 & n66;
  assign new_n1508 = new_n1507 ^ new_n1504;
  assign new_n1509 = new_n1508 ^ n24;
  assign new_n1510 = ~new_n1306 & n24;
  assign new_n1511 = new_n1510 ^ new_n1397;
  assign new_n1512 = ~new_n1511 & new_n1499;
  assign new_n1513 = n65 & new_n1512;
  assign new_n1514 = new_n1513 ^ new_n1509;
  assign new_n1515 = ~new_n1307 & ~new_n1404;
  assign new_n1516 = n24 & new_n1515;
  assign new_n1517 = new_n1516 ^ new_n1514;
  assign new_n1518 = ~new_n1198 & n69;
  assign new_n1519 = ~new_n339 & new_n1193;
  assign new_n1520 = new_n1519 ^ new_n1518;
  assign new_n1521 = n70 & new_n1192;
  assign new_n1522 = n68 & new_n1204;
  assign new_n1523 = new_n1522 ^ new_n1521;
  assign new_n1524 = new_n1523 ^ new_n1520;
  assign new_n1525 = new_n1524 ^ n21;
  assign new_n1526 = new_n1525 ^ new_n1517;
  assign new_n1527 = new_n1412 ^ new_n1395;
  assign new_n1528 = ~new_n1413 & new_n1527;
  assign new_n1529 = new_n1528 ^ new_n1395;
  assign new_n1530 = new_n1529 ^ new_n1526;
  assign new_n1531 = ~new_n930 & n72;
  assign new_n1532 = new_n534 & new_n925;
  assign new_n1533 = new_n1532 ^ new_n1531;
  assign new_n1534 = n73 & new_n924;
  assign new_n1535 = n71 & new_n936;
  assign new_n1536 = new_n1535 ^ new_n1534;
  assign new_n1537 = new_n1536 ^ new_n1533;
  assign new_n1538 = new_n1537 ^ n18;
  assign new_n1539 = new_n1538 ^ new_n1530;
  assign new_n1540 = new_n1426 ^ new_n1414;
  assign new_n1541 = ~new_n1423 & new_n1540;
  assign new_n1542 = new_n1541 ^ new_n1426;
  assign new_n1543 = new_n1542 ^ new_n1539;
  assign new_n1544 = n75 & new_n707;
  assign new_n1545 = ~new_n737 & new_n701;
  assign new_n1546 = new_n1545 ^ new_n1544;
  assign new_n1547 = n76 & new_n700;
  assign new_n1548 = n74 & new_n787;
  assign new_n1549 = new_n1548 ^ new_n1547;
  assign new_n1550 = new_n1549 ^ new_n1546;
  assign new_n1551 = new_n1550 ^ n15;
  assign new_n1552 = new_n1551 ^ new_n1543;
  assign new_n1553 = new_n1439 ^ new_n1427;
  assign new_n1554 = ~new_n1436 & new_n1553;
  assign new_n1555 = new_n1554 ^ new_n1439;
  assign new_n1556 = new_n1555 ^ new_n1552;
  assign new_n1557 = n78 & new_n499;
  assign new_n1558 = ~new_n506 & ~new_n982;
  assign new_n1559 = new_n1558 ^ new_n1557;
  assign new_n1560 = ~new_n505 & n79;
  assign new_n1561 = n77 & new_n579;
  assign new_n1562 = new_n1561 ^ new_n1560;
  assign new_n1563 = new_n1562 ^ new_n1559;
  assign new_n1564 = new_n1563 ^ n12;
  assign new_n1565 = new_n1564 ^ new_n1556;
  assign new_n1566 = new_n1452 ^ new_n1440;
  assign new_n1567 = ~new_n1449 & new_n1566;
  assign new_n1568 = new_n1567 ^ new_n1452;
  assign new_n1569 = new_n1568 ^ new_n1565;
  assign new_n1570 = n81 & new_n354;
  assign new_n1571 = new_n349 & new_n1263;
  assign new_n1572 = new_n1571 ^ new_n1570;
  assign new_n1573 = n82 & new_n348;
  assign new_n1574 = n80 & new_n391;
  assign new_n1575 = new_n1574 ^ new_n1573;
  assign new_n1576 = new_n1575 ^ new_n1572;
  assign new_n1577 = new_n1576 ^ n9;
  assign new_n1578 = new_n1577 ^ new_n1569;
  assign new_n1579 = new_n1465 ^ new_n1453;
  assign new_n1580 = ~new_n1462 & new_n1579;
  assign new_n1581 = new_n1580 ^ new_n1465;
  assign new_n1582 = new_n1581 ^ new_n1578;
  assign new_n1583 = n84 & new_n218;
  assign new_n1584 = new_n1277 ^ n85;
  assign new_n1585 = new_n208 & new_n1584;
  assign new_n1586 = new_n1585 ^ new_n1583;
  assign new_n1587 = n85 & new_n207;
  assign new_n1588 = n83 & new_n212;
  assign new_n1589 = new_n1588 ^ new_n1587;
  assign new_n1590 = new_n1589 ^ new_n1586;
  assign new_n1591 = new_n1590 ^ n6;
  assign new_n1592 = new_n1591 ^ new_n1582;
  assign new_n1593 = new_n1479 ^ new_n1466;
  assign new_n1594 = ~new_n1476 & new_n1593;
  assign new_n1595 = new_n1594 ^ new_n1479;
  assign new_n1596 = new_n1595 ^ new_n1592;
  assign new_n1597 = n87 ^ n3;
  assign new_n1598 = ~n86 & n3;
  assign new_n1599 = new_n1598 ^ new_n1597;
  assign new_n1600 = ~n2 & new_n1599;
  assign new_n1601 = new_n1600 ^ new_n1597;
  assign new_n1602 = n87 ^ n86;
  assign new_n1603 = ~new_n1482 & new_n1602;
  assign new_n1604 = ~new_n1603 & new_n155;
  assign new_n1605 = new_n1604 ^ n2;
  assign new_n1606 = new_n1605 ^ n88;
  assign new_n1607 = new_n1606 ^ new_n1601;
  assign new_n1608 = ~n1 & new_n1607;
  assign new_n1609 = new_n1608 ^ new_n1606;
  assign new_n1610 = new_n1609 ^ new_n1596;
  assign new_n1611 = new_n1497 ^ new_n1480;
  assign new_n1612 = ~new_n1494 & new_n1611;
  assign new_n1613 = new_n1612 ^ new_n1497;
  assign new_n1614 = new_n1613 ^ new_n1610;
  assign new_n1615 = new_n1514 & new_n1516;
  assign new_n1616 = ~new_n259 & new_n1501;
  assign new_n1617 = ~new_n1506 & n67;
  assign new_n1618 = new_n1617 ^ new_n1616;
  assign new_n1619 = n68 & new_n1500;
  assign new_n1620 = n66 & new_n1512;
  assign new_n1621 = new_n1620 ^ new_n1619;
  assign new_n1622 = new_n1621 ^ new_n1618;
  assign new_n1623 = new_n1622 ^ n24;
  assign new_n1624 = n25 ^ n24;
  assign new_n1625 = n65 & new_n1624;
  assign new_n1626 = new_n1625 ^ new_n1623;
  assign new_n1627 = new_n1626 ^ new_n1615;
  assign new_n1628 = ~new_n1198 & n70;
  assign new_n1629 = ~new_n402 & new_n1193;
  assign new_n1630 = new_n1629 ^ new_n1628;
  assign new_n1631 = n71 & new_n1192;
  assign new_n1632 = n69 & new_n1204;
  assign new_n1633 = new_n1632 ^ new_n1631;
  assign new_n1634 = new_n1633 ^ new_n1630;
  assign new_n1635 = new_n1634 ^ n21;
  assign new_n1636 = new_n1635 ^ new_n1627;
  assign new_n1637 = new_n1529 ^ new_n1517;
  assign new_n1638 = ~new_n1526 & new_n1637;
  assign new_n1639 = new_n1638 ^ new_n1529;
  assign new_n1640 = new_n1639 ^ new_n1636;
  assign new_n1641 = ~new_n930 & n73;
  assign new_n1642 = new_n595 & new_n925;
  assign new_n1643 = new_n1642 ^ new_n1641;
  assign new_n1644 = n74 & new_n924;
  assign new_n1645 = n72 & new_n936;
  assign new_n1646 = new_n1645 ^ new_n1644;
  assign new_n1647 = new_n1646 ^ new_n1643;
  assign new_n1648 = new_n1647 ^ n18;
  assign new_n1649 = new_n1648 ^ new_n1640;
  assign new_n1650 = new_n1542 ^ new_n1530;
  assign new_n1651 = ~new_n1539 & new_n1650;
  assign new_n1652 = new_n1651 ^ new_n1542;
  assign new_n1653 = new_n1652 ^ new_n1649;
  assign new_n1654 = n76 & new_n707;
  assign new_n1655 = ~new_n812 & new_n701;
  assign new_n1656 = new_n1655 ^ new_n1654;
  assign new_n1657 = n77 & new_n700;
  assign new_n1658 = n75 & new_n787;
  assign new_n1659 = new_n1658 ^ new_n1657;
  assign new_n1660 = new_n1659 ^ new_n1656;
  assign new_n1661 = new_n1660 ^ n15;
  assign new_n1662 = new_n1661 ^ new_n1653;
  assign new_n1663 = new_n1555 ^ new_n1543;
  assign new_n1664 = ~new_n1552 & new_n1663;
  assign new_n1665 = new_n1664 ^ new_n1555;
  assign new_n1666 = new_n1665 ^ new_n1662;
  assign new_n1667 = n79 & new_n499;
  assign new_n1668 = ~new_n506 & new_n1069;
  assign new_n1669 = new_n1668 ^ new_n1667;
  assign new_n1670 = ~new_n505 & n80;
  assign new_n1671 = n78 & new_n579;
  assign new_n1672 = new_n1671 ^ new_n1670;
  assign new_n1673 = new_n1672 ^ new_n1669;
  assign new_n1674 = new_n1673 ^ n12;
  assign new_n1675 = new_n1674 ^ new_n1666;
  assign new_n1676 = new_n1568 ^ new_n1556;
  assign new_n1677 = ~new_n1565 & new_n1676;
  assign new_n1678 = new_n1677 ^ new_n1568;
  assign new_n1679 = new_n1678 ^ new_n1675;
  assign new_n1680 = n82 & new_n354;
  assign new_n1681 = new_n349 & new_n1363;
  assign new_n1682 = new_n1681 ^ new_n1680;
  assign new_n1683 = n83 & new_n348;
  assign new_n1684 = n81 & new_n391;
  assign new_n1685 = new_n1684 ^ new_n1683;
  assign new_n1686 = new_n1685 ^ new_n1682;
  assign new_n1687 = new_n1686 ^ n9;
  assign new_n1688 = new_n1687 ^ new_n1679;
  assign new_n1689 = new_n1581 ^ new_n1569;
  assign new_n1690 = ~new_n1578 & new_n1689;
  assign new_n1691 = new_n1690 ^ new_n1581;
  assign new_n1692 = new_n1691 ^ new_n1688;
  assign new_n1693 = n85 & new_n218;
  assign new_n1694 = new_n1377 ^ n86;
  assign new_n1695 = new_n208 & new_n1694;
  assign new_n1696 = new_n1695 ^ new_n1693;
  assign new_n1697 = n86 & new_n207;
  assign new_n1698 = n84 & new_n212;
  assign new_n1699 = new_n1698 ^ new_n1697;
  assign new_n1700 = new_n1699 ^ new_n1696;
  assign new_n1701 = new_n1700 ^ n6;
  assign new_n1702 = new_n1701 ^ new_n1692;
  assign new_n1703 = new_n1595 ^ new_n1582;
  assign new_n1704 = ~new_n1592 & new_n1703;
  assign new_n1705 = new_n1704 ^ new_n1595;
  assign new_n1706 = new_n1705 ^ new_n1702;
  assign new_n1707 = n88 ^ n87;
  assign new_n1708 = ~new_n1603 & new_n1707;
  assign new_n1709 = ~new_n1708 & new_n155;
  assign new_n1710 = new_n1709 ^ n2;
  assign new_n1711 = new_n1710 ^ n89;
  assign new_n1712 = n88 ^ n3;
  assign new_n1713 = ~n87 & n3;
  assign new_n1714 = new_n1713 ^ new_n1712;
  assign new_n1715 = ~n2 & new_n1714;
  assign new_n1716 = new_n1715 ^ new_n1712;
  assign new_n1717 = new_n1716 ^ new_n1711;
  assign new_n1718 = ~n1 & new_n1717;
  assign new_n1719 = new_n1718 ^ new_n1711;
  assign new_n1720 = new_n1719 ^ new_n1706;
  assign new_n1721 = new_n1613 ^ new_n1596;
  assign new_n1722 = ~new_n1610 & new_n1721;
  assign new_n1723 = new_n1722 ^ new_n1613;
  assign new_n1724 = new_n1723 ^ new_n1720;
  assign new_n1725 = ~new_n1615 & ~new_n1625;
  assign new_n1726 = ~new_n1725 & new_n1623;
  assign new_n1727 = ~new_n1506 & n68;
  assign new_n1728 = ~new_n304 & new_n1501;
  assign new_n1729 = new_n1728 ^ new_n1727;
  assign new_n1730 = n69 & new_n1500;
  assign new_n1731 = n67 & new_n1512;
  assign new_n1732 = new_n1731 ^ new_n1730;
  assign new_n1733 = new_n1732 ^ new_n1729;
  assign new_n1734 = new_n1733 ^ n24;
  assign new_n1735 = n66 ^ n25;
  assign new_n1736 = ~new_n1735 & new_n1624;
  assign new_n1737 = new_n1736 ^ n24;
  assign new_n1738 = new_n1737 ^ n26;
  assign new_n1739 = n24 & n25;
  assign new_n1740 = new_n1739 ^ n26;
  assign new_n1741 = ~n65 & new_n1740;
  assign new_n1742 = new_n1741 ^ new_n1738;
  assign new_n1743 = new_n1742 ^ new_n1734;
  assign new_n1744 = new_n1743 ^ new_n1726;
  assign new_n1745 = ~new_n1198 & n71;
  assign new_n1746 = ~new_n459 & new_n1193;
  assign new_n1747 = new_n1746 ^ new_n1745;
  assign new_n1748 = n72 & new_n1192;
  assign new_n1749 = n70 & new_n1204;
  assign new_n1750 = new_n1749 ^ new_n1748;
  assign new_n1751 = new_n1750 ^ new_n1747;
  assign new_n1752 = new_n1751 ^ n21;
  assign new_n1753 = new_n1752 ^ new_n1744;
  assign new_n1754 = new_n1639 ^ new_n1627;
  assign new_n1755 = ~new_n1636 & new_n1754;
  assign new_n1756 = new_n1755 ^ new_n1639;
  assign new_n1757 = new_n1756 ^ new_n1753;
  assign new_n1758 = ~new_n930 & n74;
  assign new_n1759 = new_n660 & new_n925;
  assign new_n1760 = new_n1759 ^ new_n1758;
  assign new_n1761 = n75 & new_n924;
  assign new_n1762 = n73 & new_n936;
  assign new_n1763 = new_n1762 ^ new_n1761;
  assign new_n1764 = new_n1763 ^ new_n1760;
  assign new_n1765 = new_n1764 ^ n18;
  assign new_n1766 = new_n1765 ^ new_n1757;
  assign new_n1767 = new_n1652 ^ new_n1640;
  assign new_n1768 = ~new_n1649 & new_n1767;
  assign new_n1769 = new_n1768 ^ new_n1652;
  assign new_n1770 = new_n1769 ^ new_n1766;
  assign new_n1771 = n77 & new_n707;
  assign new_n1772 = ~new_n891 & new_n701;
  assign new_n1773 = new_n1772 ^ new_n1771;
  assign new_n1774 = n78 & new_n700;
  assign new_n1775 = n76 & new_n787;
  assign new_n1776 = new_n1775 ^ new_n1774;
  assign new_n1777 = new_n1776 ^ new_n1773;
  assign new_n1778 = new_n1777 ^ n15;
  assign new_n1779 = new_n1778 ^ new_n1770;
  assign new_n1780 = new_n1665 ^ new_n1653;
  assign new_n1781 = ~new_n1662 & new_n1780;
  assign new_n1782 = new_n1781 ^ new_n1665;
  assign new_n1783 = new_n1782 ^ new_n1779;
  assign new_n1784 = n80 & new_n499;
  assign new_n1785 = ~new_n506 & new_n1161;
  assign new_n1786 = new_n1785 ^ new_n1784;
  assign new_n1787 = ~new_n505 & n81;
  assign new_n1788 = n79 & new_n579;
  assign new_n1789 = new_n1788 ^ new_n1787;
  assign new_n1790 = new_n1789 ^ new_n1786;
  assign new_n1791 = new_n1790 ^ n12;
  assign new_n1792 = new_n1791 ^ new_n1783;
  assign new_n1793 = new_n1678 ^ new_n1666;
  assign new_n1794 = ~new_n1675 & new_n1793;
  assign new_n1795 = new_n1794 ^ new_n1678;
  assign new_n1796 = new_n1795 ^ new_n1792;
  assign new_n1797 = n83 & new_n354;
  assign new_n1798 = new_n349 & new_n1468;
  assign new_n1799 = new_n1798 ^ new_n1797;
  assign new_n1800 = n84 & new_n348;
  assign new_n1801 = n82 & new_n391;
  assign new_n1802 = new_n1801 ^ new_n1800;
  assign new_n1803 = new_n1802 ^ new_n1799;
  assign new_n1804 = new_n1803 ^ n9;
  assign new_n1805 = new_n1804 ^ new_n1796;
  assign new_n1806 = new_n1691 ^ new_n1679;
  assign new_n1807 = ~new_n1688 & new_n1806;
  assign new_n1808 = new_n1807 ^ new_n1691;
  assign new_n1809 = new_n1808 ^ new_n1805;
  assign new_n1810 = n86 & new_n218;
  assign new_n1811 = new_n1482 ^ n87;
  assign new_n1812 = new_n208 & new_n1811;
  assign new_n1813 = new_n1812 ^ new_n1810;
  assign new_n1814 = n87 & new_n207;
  assign new_n1815 = n85 & new_n212;
  assign new_n1816 = new_n1815 ^ new_n1814;
  assign new_n1817 = new_n1816 ^ new_n1813;
  assign new_n1818 = new_n1817 ^ n6;
  assign new_n1819 = new_n1818 ^ new_n1809;
  assign new_n1820 = new_n1705 ^ new_n1692;
  assign new_n1821 = ~new_n1702 & new_n1820;
  assign new_n1822 = new_n1821 ^ new_n1705;
  assign new_n1823 = new_n1822 ^ new_n1819;
  assign new_n1824 = n89 ^ n88;
  assign new_n1825 = ~new_n1708 & new_n1824;
  assign new_n1826 = ~new_n1825 & new_n155;
  assign new_n1827 = new_n1826 ^ n2;
  assign new_n1828 = new_n1827 ^ n90;
  assign new_n1829 = n89 ^ n3;
  assign new_n1830 = ~n88 & n3;
  assign new_n1831 = new_n1830 ^ new_n1829;
  assign new_n1832 = ~n2 & new_n1831;
  assign new_n1833 = new_n1832 ^ new_n1829;
  assign new_n1834 = new_n1833 ^ new_n1828;
  assign new_n1835 = ~n1 & new_n1834;
  assign new_n1836 = new_n1835 ^ new_n1828;
  assign new_n1837 = new_n1836 ^ new_n1823;
  assign new_n1838 = new_n1723 ^ new_n1706;
  assign new_n1839 = ~new_n1720 & new_n1838;
  assign new_n1840 = new_n1839 ^ new_n1723;
  assign new_n1841 = new_n1840 ^ new_n1837;
  assign new_n1842 = ~new_n930 & n75;
  assign new_n1843 = ~new_n737 & new_n925;
  assign new_n1844 = new_n1843 ^ new_n1842;
  assign new_n1845 = n76 & new_n924;
  assign new_n1846 = n74 & new_n936;
  assign new_n1847 = new_n1846 ^ new_n1845;
  assign new_n1848 = new_n1847 ^ new_n1844;
  assign new_n1849 = new_n1848 ^ n18;
  assign new_n1850 = new_n1769 ^ new_n1757;
  assign new_n1851 = ~new_n1766 & new_n1850;
  assign new_n1852 = new_n1851 ^ new_n1769;
  assign new_n1853 = new_n1852 ^ new_n1849;
  assign new_n1854 = ~new_n1506 & n69;
  assign new_n1855 = ~new_n339 & new_n1501;
  assign new_n1856 = new_n1855 ^ new_n1854;
  assign new_n1857 = n70 & new_n1500;
  assign new_n1858 = n68 & new_n1512;
  assign new_n1859 = new_n1858 ^ new_n1857;
  assign new_n1860 = new_n1859 ^ new_n1856;
  assign new_n1861 = new_n1860 ^ n24;
  assign new_n1862 = n27 ^ n26;
  assign new_n1863 = ~new_n1862 & new_n1624;
  assign new_n1864 = new_n1863 ^ new_n1624;
  assign new_n1865 = ~new_n151 & new_n1864;
  assign new_n1866 = ~new_n1624 & n27;
  assign new_n1867 = new_n1866 ^ new_n1739;
  assign new_n1868 = new_n1862 & new_n1867;
  assign new_n1869 = n65 & new_n1868;
  assign new_n1870 = new_n1869 ^ new_n1865;
  assign new_n1871 = n67 & new_n1624;
  assign new_n1872 = new_n1871 ^ new_n1870;
  assign new_n1873 = ~new_n1624 & n26;
  assign new_n1874 = new_n1873 ^ new_n1739;
  assign new_n1875 = n66 & new_n1874;
  assign new_n1876 = new_n1875 ^ new_n1872;
  assign new_n1877 = ~new_n1625 & ~new_n1742;
  assign new_n1878 = n27 & new_n1877;
  assign new_n1879 = new_n1878 ^ n27;
  assign new_n1880 = new_n1879 ^ new_n1876;
  assign new_n1881 = new_n1880 ^ new_n1861;
  assign new_n1882 = new_n1734 ^ new_n1726;
  assign new_n1883 = ~new_n1743 & new_n1882;
  assign new_n1884 = new_n1883 ^ new_n1726;
  assign new_n1885 = new_n1884 ^ new_n1881;
  assign new_n1886 = ~new_n1198 & n72;
  assign new_n1887 = new_n534 & new_n1193;
  assign new_n1888 = new_n1887 ^ new_n1886;
  assign new_n1889 = n73 & new_n1192;
  assign new_n1890 = n71 & new_n1204;
  assign new_n1891 = new_n1890 ^ new_n1889;
  assign new_n1892 = new_n1891 ^ new_n1888;
  assign new_n1893 = new_n1892 ^ n21;
  assign new_n1894 = new_n1893 ^ new_n1885;
  assign new_n1895 = new_n1756 ^ new_n1744;
  assign new_n1896 = ~new_n1753 & new_n1895;
  assign new_n1897 = new_n1896 ^ new_n1756;
  assign new_n1898 = new_n1897 ^ new_n1894;
  assign new_n1899 = new_n1898 ^ new_n1853;
  assign new_n1900 = n78 & new_n707;
  assign new_n1901 = ~new_n982 & new_n701;
  assign new_n1902 = new_n1901 ^ new_n1900;
  assign new_n1903 = n79 & new_n700;
  assign new_n1904 = n77 & new_n787;
  assign new_n1905 = new_n1904 ^ new_n1903;
  assign new_n1906 = new_n1905 ^ new_n1902;
  assign new_n1907 = new_n1906 ^ n15;
  assign new_n1908 = new_n1907 ^ new_n1899;
  assign new_n1909 = new_n1782 ^ new_n1770;
  assign new_n1910 = ~new_n1779 & new_n1909;
  assign new_n1911 = new_n1910 ^ new_n1782;
  assign new_n1912 = new_n1911 ^ new_n1908;
  assign new_n1913 = n81 & new_n499;
  assign new_n1914 = ~new_n506 & new_n1263;
  assign new_n1915 = new_n1914 ^ new_n1913;
  assign new_n1916 = ~new_n505 & n82;
  assign new_n1917 = n80 & new_n579;
  assign new_n1918 = new_n1917 ^ new_n1916;
  assign new_n1919 = new_n1918 ^ new_n1915;
  assign new_n1920 = new_n1919 ^ n12;
  assign new_n1921 = new_n1920 ^ new_n1912;
  assign new_n1922 = new_n1795 ^ new_n1783;
  assign new_n1923 = ~new_n1792 & new_n1922;
  assign new_n1924 = new_n1923 ^ new_n1795;
  assign new_n1925 = new_n1924 ^ new_n1921;
  assign new_n1926 = n84 & new_n354;
  assign new_n1927 = new_n349 & new_n1584;
  assign new_n1928 = new_n1927 ^ new_n1926;
  assign new_n1929 = n85 & new_n348;
  assign new_n1930 = n83 & new_n391;
  assign new_n1931 = new_n1930 ^ new_n1929;
  assign new_n1932 = new_n1931 ^ new_n1928;
  assign new_n1933 = new_n1932 ^ n9;
  assign new_n1934 = new_n1933 ^ new_n1925;
  assign new_n1935 = new_n1808 ^ new_n1796;
  assign new_n1936 = ~new_n1805 & new_n1935;
  assign new_n1937 = new_n1936 ^ new_n1808;
  assign new_n1938 = new_n1937 ^ new_n1934;
  assign new_n1939 = n87 & new_n218;
  assign new_n1940 = new_n1603 ^ n88;
  assign new_n1941 = new_n208 & new_n1940;
  assign new_n1942 = new_n1941 ^ new_n1939;
  assign new_n1943 = n88 & new_n207;
  assign new_n1944 = n86 & new_n212;
  assign new_n1945 = new_n1944 ^ new_n1943;
  assign new_n1946 = new_n1945 ^ new_n1942;
  assign new_n1947 = new_n1946 ^ n6;
  assign new_n1948 = new_n1947 ^ new_n1938;
  assign new_n1949 = new_n1822 ^ new_n1809;
  assign new_n1950 = ~new_n1819 & new_n1949;
  assign new_n1951 = new_n1950 ^ new_n1822;
  assign new_n1952 = new_n1951 ^ new_n1948;
  assign new_n1953 = n90 ^ n89;
  assign new_n1954 = ~new_n1825 & new_n1953;
  assign new_n1955 = ~new_n1954 & new_n155;
  assign new_n1956 = new_n1955 ^ n2;
  assign new_n1957 = new_n1956 ^ n91;
  assign new_n1958 = ~n89 & n3;
  assign new_n1959 = n90 ^ n3;
  assign new_n1960 = new_n1959 ^ new_n1958;
  assign new_n1961 = n2 & new_n1960;
  assign new_n1962 = new_n1961 ^ new_n1958;
  assign new_n1963 = new_n1962 ^ new_n1957;
  assign new_n1964 = ~n1 & new_n1963;
  assign new_n1965 = new_n1964 ^ new_n1957;
  assign new_n1966 = new_n1965 ^ new_n1952;
  assign new_n1967 = new_n1840 ^ new_n1823;
  assign new_n1968 = ~new_n1837 & new_n1967;
  assign new_n1969 = new_n1968 ^ new_n1840;
  assign new_n1970 = new_n1969 ^ new_n1966;
  assign new_n1971 = ~new_n1506 & n70;
  assign new_n1972 = ~new_n402 & new_n1501;
  assign new_n1973 = new_n1972 ^ new_n1971;
  assign new_n1974 = n71 & new_n1500;
  assign new_n1975 = n69 & new_n1512;
  assign new_n1976 = new_n1975 ^ new_n1974;
  assign new_n1977 = new_n1976 ^ new_n1973;
  assign new_n1978 = new_n1977 ^ n24;
  assign new_n1979 = ~new_n1876 & new_n1878;
  assign new_n1980 = n28 ^ n27;
  assign new_n1981 = n65 & new_n1980;
  assign new_n1982 = new_n1981 ^ new_n1979;
  assign new_n1983 = ~new_n154 & ~new_n1862;
  assign new_n1984 = new_n1983 ^ new_n259;
  assign new_n1985 = ~new_n1984 & new_n1624;
  assign new_n1986 = n67 & new_n1874;
  assign new_n1987 = n66 & new_n1868;
  assign new_n1988 = new_n1987 ^ new_n1986;
  assign new_n1989 = ~new_n1985 & ~new_n1988;
  assign new_n1990 = new_n1989 ^ n27;
  assign new_n1991 = new_n1990 ^ new_n1982;
  assign new_n1992 = new_n1991 ^ new_n1978;
  assign new_n1993 = new_n1884 ^ new_n1861;
  assign new_n1994 = ~new_n1881 & new_n1993;
  assign new_n1995 = new_n1994 ^ new_n1884;
  assign new_n1996 = new_n1995 ^ new_n1992;
  assign new_n1997 = ~new_n1198 & n73;
  assign new_n1998 = new_n595 & new_n1193;
  assign new_n1999 = new_n1998 ^ new_n1997;
  assign new_n2000 = n74 & new_n1192;
  assign new_n2001 = n72 & new_n1204;
  assign new_n2002 = new_n2001 ^ new_n2000;
  assign new_n2003 = new_n2002 ^ new_n1999;
  assign new_n2004 = new_n2003 ^ n21;
  assign new_n2005 = new_n2004 ^ new_n1996;
  assign new_n2006 = new_n1897 ^ new_n1885;
  assign new_n2007 = ~new_n1894 & new_n2006;
  assign new_n2008 = new_n2007 ^ new_n1897;
  assign new_n2009 = new_n2008 ^ new_n2005;
  assign new_n2010 = ~new_n930 & n76;
  assign new_n2011 = ~new_n812 & new_n925;
  assign new_n2012 = new_n2011 ^ new_n2010;
  assign new_n2013 = n77 & new_n924;
  assign new_n2014 = n75 & new_n936;
  assign new_n2015 = new_n2014 ^ new_n2013;
  assign new_n2016 = new_n2015 ^ new_n2012;
  assign new_n2017 = new_n2016 ^ n18;
  assign new_n2018 = new_n2017 ^ new_n2009;
  assign new_n2019 = new_n1898 ^ new_n1849;
  assign new_n2020 = ~new_n2019 & new_n1853;
  assign new_n2021 = new_n2020 ^ new_n1852;
  assign new_n2022 = new_n2021 ^ new_n2018;
  assign new_n2023 = n79 & new_n707;
  assign new_n2024 = new_n701 & new_n1069;
  assign new_n2025 = new_n2024 ^ new_n2023;
  assign new_n2026 = n80 & new_n700;
  assign new_n2027 = n78 & new_n787;
  assign new_n2028 = new_n2027 ^ new_n2026;
  assign new_n2029 = new_n2028 ^ new_n2025;
  assign new_n2030 = new_n2029 ^ n15;
  assign new_n2031 = new_n2030 ^ new_n2022;
  assign new_n2032 = new_n1911 ^ new_n1899;
  assign new_n2033 = ~new_n1908 & new_n2032;
  assign new_n2034 = new_n2033 ^ new_n1911;
  assign new_n2035 = new_n2034 ^ new_n2031;
  assign new_n2036 = n82 & new_n499;
  assign new_n2037 = ~new_n506 & new_n1363;
  assign new_n2038 = new_n2037 ^ new_n2036;
  assign new_n2039 = ~new_n505 & n83;
  assign new_n2040 = n81 & new_n579;
  assign new_n2041 = new_n2040 ^ new_n2039;
  assign new_n2042 = new_n2041 ^ new_n2038;
  assign new_n2043 = new_n2042 ^ n12;
  assign new_n2044 = new_n2043 ^ new_n2035;
  assign new_n2045 = new_n1924 ^ new_n1912;
  assign new_n2046 = ~new_n1921 & new_n2045;
  assign new_n2047 = new_n2046 ^ new_n1924;
  assign new_n2048 = new_n2047 ^ new_n2044;
  assign new_n2049 = n85 & new_n354;
  assign new_n2050 = new_n349 & new_n1694;
  assign new_n2051 = new_n2050 ^ new_n2049;
  assign new_n2052 = n86 & new_n348;
  assign new_n2053 = n84 & new_n391;
  assign new_n2054 = new_n2053 ^ new_n2052;
  assign new_n2055 = new_n2054 ^ new_n2051;
  assign new_n2056 = new_n2055 ^ n9;
  assign new_n2057 = new_n2056 ^ new_n2048;
  assign new_n2058 = new_n1937 ^ new_n1925;
  assign new_n2059 = ~new_n1934 & new_n2058;
  assign new_n2060 = new_n2059 ^ new_n1937;
  assign new_n2061 = new_n2060 ^ new_n2057;
  assign new_n2062 = n88 & new_n218;
  assign new_n2063 = new_n1708 ^ n89;
  assign new_n2064 = new_n208 & new_n2063;
  assign new_n2065 = new_n2064 ^ new_n2062;
  assign new_n2066 = n89 & new_n207;
  assign new_n2067 = n87 & new_n212;
  assign new_n2068 = new_n2067 ^ new_n2066;
  assign new_n2069 = new_n2068 ^ new_n2065;
  assign new_n2070 = new_n2069 ^ n6;
  assign new_n2071 = new_n2070 ^ new_n2061;
  assign new_n2072 = new_n1951 ^ new_n1938;
  assign new_n2073 = ~new_n1948 & new_n2072;
  assign new_n2074 = new_n2073 ^ new_n1951;
  assign new_n2075 = new_n2074 ^ new_n2071;
  assign new_n2076 = n91 ^ n90;
  assign new_n2077 = ~new_n1954 & new_n2076;
  assign new_n2078 = ~new_n2077 & new_n155;
  assign new_n2079 = new_n2078 ^ n2;
  assign new_n2080 = new_n2079 ^ n92;
  assign new_n2081 = ~n90 & n3;
  assign new_n2082 = n91 ^ n3;
  assign new_n2083 = new_n2082 ^ new_n2081;
  assign new_n2084 = n2 & new_n2083;
  assign new_n2085 = new_n2084 ^ new_n2081;
  assign new_n2086 = new_n2085 ^ new_n2080;
  assign new_n2087 = ~n1 & new_n2086;
  assign new_n2088 = new_n2087 ^ new_n2080;
  assign new_n2089 = new_n2088 ^ new_n2075;
  assign new_n2090 = new_n1969 ^ new_n1952;
  assign new_n2091 = ~new_n1966 & new_n2090;
  assign new_n2092 = new_n2091 ^ new_n1969;
  assign new_n2093 = new_n2092 ^ new_n2089;
  assign new_n2094 = ~new_n1506 & n71;
  assign new_n2095 = ~new_n459 & new_n1501;
  assign new_n2096 = new_n2095 ^ new_n2094;
  assign new_n2097 = n72 & new_n1500;
  assign new_n2098 = n70 & new_n1512;
  assign new_n2099 = new_n2098 ^ new_n2097;
  assign new_n2100 = new_n2099 ^ new_n2096;
  assign new_n2101 = new_n2100 ^ n24;
  assign new_n2102 = ~new_n1979 & ~new_n1981;
  assign new_n2103 = ~new_n1990 & ~new_n2102;
  assign new_n2104 = n27 & n28;
  assign new_n2105 = new_n2104 ^ n29;
  assign new_n2106 = ~n65 & new_n2105;
  assign new_n2107 = n66 ^ n28;
  assign new_n2108 = ~new_n2107 & new_n1980;
  assign new_n2109 = new_n2108 ^ n27;
  assign new_n2110 = new_n2109 ^ n29;
  assign new_n2111 = new_n2110 ^ new_n2106;
  assign new_n2112 = n68 & new_n1874;
  assign new_n2113 = ~new_n304 & new_n1864;
  assign new_n2114 = new_n2113 ^ new_n2112;
  assign new_n2115 = n69 & new_n1863;
  assign new_n2116 = n67 & new_n1868;
  assign new_n2117 = new_n2116 ^ new_n2115;
  assign new_n2118 = new_n2117 ^ new_n2114;
  assign new_n2119 = new_n2118 ^ n27;
  assign new_n2120 = new_n2119 ^ new_n2111;
  assign new_n2121 = new_n2120 ^ new_n2103;
  assign new_n2122 = new_n2121 ^ new_n2101;
  assign new_n2123 = new_n1995 ^ new_n1978;
  assign new_n2124 = new_n1992 & new_n2123;
  assign new_n2125 = new_n2124 ^ new_n1995;
  assign new_n2126 = new_n2125 ^ new_n2122;
  assign new_n2127 = ~new_n1198 & n74;
  assign new_n2128 = new_n660 & new_n1193;
  assign new_n2129 = new_n2128 ^ new_n2127;
  assign new_n2130 = n73 & new_n1204;
  assign new_n2131 = n75 & new_n1192;
  assign new_n2132 = new_n2131 ^ new_n2130;
  assign new_n2133 = new_n2132 ^ new_n2129;
  assign new_n2134 = new_n2133 ^ n21;
  assign new_n2135 = new_n2134 ^ new_n2126;
  assign new_n2136 = new_n2008 ^ new_n1996;
  assign new_n2137 = ~new_n2136 & new_n2005;
  assign new_n2138 = new_n2137 ^ new_n2008;
  assign new_n2139 = new_n2138 ^ new_n2135;
  assign new_n2140 = ~new_n930 & n77;
  assign new_n2141 = ~new_n891 & new_n925;
  assign new_n2142 = new_n2141 ^ new_n2140;
  assign new_n2143 = n78 & new_n924;
  assign new_n2144 = n76 & new_n936;
  assign new_n2145 = new_n2144 ^ new_n2143;
  assign new_n2146 = new_n2145 ^ new_n2142;
  assign new_n2147 = new_n2146 ^ n18;
  assign new_n2148 = new_n2147 ^ new_n2139;
  assign new_n2149 = new_n2021 ^ new_n2009;
  assign new_n2150 = ~new_n2149 & new_n2018;
  assign new_n2151 = new_n2150 ^ new_n2021;
  assign new_n2152 = new_n2151 ^ new_n2148;
  assign new_n2153 = n80 & new_n707;
  assign new_n2154 = new_n701 & new_n1161;
  assign new_n2155 = new_n2154 ^ new_n2153;
  assign new_n2156 = n81 & new_n700;
  assign new_n2157 = n79 & new_n787;
  assign new_n2158 = new_n2157 ^ new_n2156;
  assign new_n2159 = new_n2158 ^ new_n2155;
  assign new_n2160 = new_n2159 ^ n15;
  assign new_n2161 = new_n2160 ^ new_n2152;
  assign new_n2162 = new_n2034 ^ new_n2022;
  assign new_n2163 = ~new_n2162 & new_n2031;
  assign new_n2164 = new_n2163 ^ new_n2034;
  assign new_n2165 = new_n2164 ^ new_n2161;
  assign new_n2166 = n83 & new_n499;
  assign new_n2167 = ~new_n506 & new_n1468;
  assign new_n2168 = new_n2167 ^ new_n2166;
  assign new_n2169 = ~new_n505 & n84;
  assign new_n2170 = n82 & new_n579;
  assign new_n2171 = new_n2170 ^ new_n2169;
  assign new_n2172 = new_n2171 ^ new_n2168;
  assign new_n2173 = new_n2172 ^ n12;
  assign new_n2174 = new_n2173 ^ new_n2165;
  assign new_n2175 = new_n2047 ^ new_n2035;
  assign new_n2176 = ~new_n2175 & new_n2044;
  assign new_n2177 = new_n2176 ^ new_n2047;
  assign new_n2178 = new_n2177 ^ new_n2174;
  assign new_n2179 = n86 & new_n354;
  assign new_n2180 = new_n349 & new_n1811;
  assign new_n2181 = new_n2180 ^ new_n2179;
  assign new_n2182 = n87 & new_n348;
  assign new_n2183 = n85 & new_n391;
  assign new_n2184 = new_n2183 ^ new_n2182;
  assign new_n2185 = new_n2184 ^ new_n2181;
  assign new_n2186 = new_n2185 ^ n9;
  assign new_n2187 = new_n2186 ^ new_n2178;
  assign new_n2188 = new_n2060 ^ new_n2048;
  assign new_n2189 = ~new_n2188 & new_n2057;
  assign new_n2190 = new_n2189 ^ new_n2060;
  assign new_n2191 = new_n2190 ^ new_n2187;
  assign new_n2192 = n89 & new_n218;
  assign new_n2193 = new_n1825 ^ n90;
  assign new_n2194 = new_n208 & new_n2193;
  assign new_n2195 = new_n2194 ^ new_n2192;
  assign new_n2196 = n90 & new_n207;
  assign new_n2197 = n88 & new_n212;
  assign new_n2198 = new_n2197 ^ new_n2196;
  assign new_n2199 = new_n2198 ^ new_n2195;
  assign new_n2200 = new_n2199 ^ n6;
  assign new_n2201 = new_n2200 ^ new_n2191;
  assign new_n2202 = new_n2074 ^ new_n2061;
  assign new_n2203 = ~new_n2202 & new_n2071;
  assign new_n2204 = new_n2203 ^ new_n2074;
  assign new_n2205 = new_n2204 ^ new_n2201;
  assign new_n2206 = n92 ^ n91;
  assign new_n2207 = ~new_n2077 & new_n2206;
  assign new_n2208 = ~new_n2207 & new_n155;
  assign new_n2209 = new_n2208 ^ n2;
  assign new_n2210 = new_n2209 ^ n93;
  assign new_n2211 = n92 ^ n3;
  assign new_n2212 = ~n91 & ~new_n2082;
  assign new_n2213 = new_n2212 ^ new_n2211;
  assign new_n2214 = new_n2213 ^ n91;
  assign new_n2215 = ~new_n2214 & new_n241;
  assign new_n2216 = new_n2215 ^ new_n2212;
  assign new_n2217 = new_n2216 ^ n91;
  assign new_n2218 = new_n2217 ^ new_n2210;
  assign new_n2219 = ~n1 & ~new_n2218;
  assign new_n2220 = new_n2219 ^ new_n2210;
  assign new_n2221 = new_n2220 ^ new_n2205;
  assign new_n2222 = new_n2092 ^ new_n2075;
  assign new_n2223 = ~new_n2222 & new_n2089;
  assign new_n2224 = new_n2223 ^ new_n2092;
  assign new_n2225 = new_n2224 ^ new_n2221;
  assign new_n2226 = ~new_n1506 & n72;
  assign new_n2227 = new_n534 & new_n1501;
  assign new_n2228 = new_n2227 ^ new_n2226;
  assign new_n2229 = n73 & new_n1500;
  assign new_n2230 = n71 & new_n1512;
  assign new_n2231 = new_n2230 ^ new_n2229;
  assign new_n2232 = new_n2231 ^ new_n2228;
  assign new_n2233 = new_n2232 ^ n24;
  assign new_n2234 = n29 & n65;
  assign new_n2235 = new_n2234 ^ n65;
  assign new_n2236 = ~new_n2235 & n30;
  assign new_n2237 = ~new_n1981 & ~new_n2111;
  assign new_n2238 = new_n2236 & new_n2237;
  assign new_n2239 = n30 ^ n29;
  assign new_n2240 = ~new_n2239 & new_n1980;
  assign new_n2241 = new_n2240 ^ new_n1980;
  assign new_n2242 = ~new_n151 & new_n2241;
  assign new_n2243 = n67 & new_n1980;
  assign new_n2244 = new_n2243 ^ new_n2242;
  assign new_n2245 = ~new_n1980 & n29;
  assign new_n2246 = new_n2245 ^ new_n2104;
  assign new_n2247 = n66 & new_n2246;
  assign new_n2248 = new_n2247 ^ new_n2244;
  assign new_n2249 = ~new_n2248 & new_n2238;
  assign new_n2250 = new_n2248 ^ n30;
  assign new_n2251 = new_n2104 & new_n2234;
  assign new_n2252 = new_n2251 ^ new_n2237;
  assign new_n2253 = ~new_n2248 & new_n2252;
  assign new_n2254 = new_n2253 ^ new_n2237;
  assign new_n2255 = ~new_n2250 & ~new_n2254;
  assign new_n2256 = ~new_n2249 & ~new_n2255;
  assign new_n2257 = n69 & new_n1874;
  assign new_n2258 = ~new_n339 & new_n1864;
  assign new_n2259 = new_n2258 ^ new_n2257;
  assign new_n2260 = n70 & new_n1863;
  assign new_n2261 = n68 & new_n1868;
  assign new_n2262 = new_n2261 ^ new_n2260;
  assign new_n2263 = new_n2262 ^ new_n2259;
  assign new_n2264 = new_n2263 ^ n27;
  assign new_n2265 = new_n2264 ^ new_n2256;
  assign new_n2266 = new_n2119 ^ new_n2103;
  assign new_n2267 = ~new_n2120 & new_n2266;
  assign new_n2268 = new_n2267 ^ new_n2103;
  assign new_n2269 = new_n2268 ^ new_n2265;
  assign new_n2270 = new_n2269 ^ new_n2233;
  assign new_n2271 = new_n2125 ^ new_n2101;
  assign new_n2272 = ~new_n2122 & new_n2271;
  assign new_n2273 = new_n2272 ^ new_n2125;
  assign new_n2274 = new_n2273 ^ new_n2270;
  assign new_n2275 = ~new_n1198 & n75;
  assign new_n2276 = ~new_n737 & new_n1193;
  assign new_n2277 = new_n2276 ^ new_n2275;
  assign new_n2278 = n74 & new_n1204;
  assign new_n2279 = n76 & new_n1192;
  assign new_n2280 = new_n2279 ^ new_n2278;
  assign new_n2281 = new_n2280 ^ new_n2277;
  assign new_n2282 = new_n2281 ^ n21;
  assign new_n2283 = new_n2282 ^ new_n2274;
  assign new_n2284 = new_n2138 ^ new_n2126;
  assign new_n2285 = ~new_n2135 & new_n2284;
  assign new_n2286 = new_n2285 ^ new_n2138;
  assign new_n2287 = new_n2286 ^ new_n2283;
  assign new_n2288 = ~new_n930 & n78;
  assign new_n2289 = ~new_n982 & new_n925;
  assign new_n2290 = new_n2289 ^ new_n2288;
  assign new_n2291 = n79 & new_n924;
  assign new_n2292 = n77 & new_n936;
  assign new_n2293 = new_n2292 ^ new_n2291;
  assign new_n2294 = new_n2293 ^ new_n2290;
  assign new_n2295 = new_n2294 ^ n18;
  assign new_n2296 = new_n2295 ^ new_n2287;
  assign new_n2297 = new_n2151 ^ new_n2139;
  assign new_n2298 = ~new_n2148 & new_n2297;
  assign new_n2299 = new_n2298 ^ new_n2151;
  assign new_n2300 = new_n2299 ^ new_n2296;
  assign new_n2301 = n81 & new_n707;
  assign new_n2302 = new_n701 & new_n1263;
  assign new_n2303 = new_n2302 ^ new_n2301;
  assign new_n2304 = n82 & new_n700;
  assign new_n2305 = n80 & new_n787;
  assign new_n2306 = new_n2305 ^ new_n2304;
  assign new_n2307 = new_n2306 ^ new_n2303;
  assign new_n2308 = new_n2307 ^ n15;
  assign new_n2309 = new_n2308 ^ new_n2300;
  assign new_n2310 = new_n2164 ^ new_n2152;
  assign new_n2311 = ~new_n2161 & new_n2310;
  assign new_n2312 = new_n2311 ^ new_n2164;
  assign new_n2313 = new_n2312 ^ new_n2309;
  assign new_n2314 = n84 & new_n499;
  assign new_n2315 = ~new_n506 & new_n1584;
  assign new_n2316 = new_n2315 ^ new_n2314;
  assign new_n2317 = ~new_n505 & n85;
  assign new_n2318 = n83 & new_n579;
  assign new_n2319 = new_n2318 ^ new_n2317;
  assign new_n2320 = new_n2319 ^ new_n2316;
  assign new_n2321 = new_n2320 ^ n12;
  assign new_n2322 = new_n2321 ^ new_n2313;
  assign new_n2323 = new_n2177 ^ new_n2165;
  assign new_n2324 = ~new_n2174 & new_n2323;
  assign new_n2325 = new_n2324 ^ new_n2177;
  assign new_n2326 = new_n2325 ^ new_n2322;
  assign new_n2327 = n87 & new_n354;
  assign new_n2328 = new_n349 & new_n1940;
  assign new_n2329 = new_n2328 ^ new_n2327;
  assign new_n2330 = n88 & new_n348;
  assign new_n2331 = n86 & new_n391;
  assign new_n2332 = new_n2331 ^ new_n2330;
  assign new_n2333 = new_n2332 ^ new_n2329;
  assign new_n2334 = new_n2333 ^ n9;
  assign new_n2335 = new_n2334 ^ new_n2326;
  assign new_n2336 = new_n2190 ^ new_n2178;
  assign new_n2337 = ~new_n2187 & new_n2336;
  assign new_n2338 = new_n2337 ^ new_n2190;
  assign new_n2339 = new_n2338 ^ new_n2335;
  assign new_n2340 = n90 & new_n218;
  assign new_n2341 = new_n1954 ^ n91;
  assign new_n2342 = new_n208 & new_n2341;
  assign new_n2343 = new_n2342 ^ new_n2340;
  assign new_n2344 = n91 & new_n207;
  assign new_n2345 = n89 & new_n212;
  assign new_n2346 = new_n2345 ^ new_n2344;
  assign new_n2347 = new_n2346 ^ new_n2343;
  assign new_n2348 = new_n2347 ^ n6;
  assign new_n2349 = new_n2348 ^ new_n2339;
  assign new_n2350 = new_n2204 ^ new_n2191;
  assign new_n2351 = ~new_n2201 & new_n2350;
  assign new_n2352 = new_n2351 ^ new_n2204;
  assign new_n2353 = new_n2352 ^ new_n2349;
  assign new_n2354 = n93 ^ n92;
  assign new_n2355 = ~new_n2207 & new_n2354;
  assign new_n2356 = ~new_n2355 & new_n155;
  assign new_n2357 = new_n2356 ^ n2;
  assign new_n2358 = new_n2357 ^ n94;
  assign new_n2359 = n93 ^ n3;
  assign new_n2360 = ~n92 & ~new_n2211;
  assign new_n2361 = new_n2360 ^ new_n2359;
  assign new_n2362 = new_n2361 ^ n92;
  assign new_n2363 = ~new_n2362 & new_n241;
  assign new_n2364 = new_n2363 ^ new_n2360;
  assign new_n2365 = new_n2364 ^ n92;
  assign new_n2366 = new_n2365 ^ new_n2358;
  assign new_n2367 = ~n1 & ~new_n2366;
  assign new_n2368 = new_n2367 ^ new_n2358;
  assign new_n2369 = new_n2368 ^ new_n2353;
  assign new_n2370 = new_n2224 ^ new_n2205;
  assign new_n2371 = ~new_n2221 & new_n2370;
  assign new_n2372 = new_n2371 ^ new_n2224;
  assign new_n2373 = new_n2372 ^ new_n2369;
  assign new_n2374 = n70 & new_n1874;
  assign new_n2375 = ~new_n402 & new_n1864;
  assign new_n2376 = new_n2375 ^ new_n2374;
  assign new_n2377 = n71 & new_n1863;
  assign new_n2378 = n69 & new_n1868;
  assign new_n2379 = new_n2378 ^ new_n2377;
  assign new_n2380 = new_n2379 ^ new_n2376;
  assign new_n2381 = new_n2380 ^ n27;
  assign new_n2382 = n31 ^ n30;
  assign new_n2383 = n65 & new_n2382;
  assign new_n2384 = new_n2383 ^ new_n2249;
  assign new_n2385 = ~new_n259 & new_n2241;
  assign new_n2386 = n67 & new_n2246;
  assign new_n2387 = new_n2386 ^ new_n2385;
  assign new_n2388 = n68 & new_n2240;
  assign new_n2389 = ~new_n1980 & n30;
  assign new_n2390 = new_n2389 ^ new_n2104;
  assign new_n2391 = new_n2239 & new_n2390;
  assign new_n2392 = n66 & new_n2391;
  assign new_n2393 = new_n2392 ^ new_n2388;
  assign new_n2394 = new_n2393 ^ new_n2387;
  assign new_n2395 = new_n2394 ^ n30;
  assign new_n2396 = new_n2395 ^ new_n2384;
  assign new_n2397 = new_n2396 ^ new_n2381;
  assign new_n2398 = new_n2268 ^ new_n2256;
  assign new_n2399 = ~new_n2265 & new_n2398;
  assign new_n2400 = new_n2399 ^ new_n2268;
  assign new_n2401 = new_n2400 ^ new_n2397;
  assign new_n2402 = ~new_n1506 & n73;
  assign new_n2403 = new_n595 & new_n1501;
  assign new_n2404 = new_n2403 ^ new_n2402;
  assign new_n2405 = n74 & new_n1500;
  assign new_n2406 = n72 & new_n1512;
  assign new_n2407 = new_n2406 ^ new_n2405;
  assign new_n2408 = new_n2407 ^ new_n2404;
  assign new_n2409 = new_n2408 ^ n24;
  assign new_n2410 = new_n2409 ^ new_n2401;
  assign new_n2411 = new_n2273 ^ new_n2233;
  assign new_n2412 = ~new_n2270 & new_n2411;
  assign new_n2413 = new_n2412 ^ new_n2273;
  assign new_n2414 = new_n2413 ^ new_n2410;
  assign new_n2415 = ~new_n1198 & n76;
  assign new_n2416 = ~new_n812 & new_n1193;
  assign new_n2417 = new_n2416 ^ new_n2415;
  assign new_n2418 = n77 & new_n1192;
  assign new_n2419 = n75 & new_n1204;
  assign new_n2420 = new_n2419 ^ new_n2418;
  assign new_n2421 = new_n2420 ^ new_n2417;
  assign new_n2422 = new_n2421 ^ n21;
  assign new_n2423 = new_n2422 ^ new_n2414;
  assign new_n2424 = new_n2286 ^ new_n2274;
  assign new_n2425 = ~new_n2283 & new_n2424;
  assign new_n2426 = new_n2425 ^ new_n2286;
  assign new_n2427 = new_n2426 ^ new_n2423;
  assign new_n2428 = ~new_n930 & n79;
  assign new_n2429 = new_n925 & new_n1069;
  assign new_n2430 = new_n2429 ^ new_n2428;
  assign new_n2431 = n80 & new_n924;
  assign new_n2432 = n78 & new_n936;
  assign new_n2433 = new_n2432 ^ new_n2431;
  assign new_n2434 = new_n2433 ^ new_n2430;
  assign new_n2435 = new_n2434 ^ n18;
  assign new_n2436 = new_n2435 ^ new_n2427;
  assign new_n2437 = new_n2299 ^ new_n2287;
  assign new_n2438 = ~new_n2296 & new_n2437;
  assign new_n2439 = new_n2438 ^ new_n2299;
  assign new_n2440 = new_n2439 ^ new_n2436;
  assign new_n2441 = n82 & new_n707;
  assign new_n2442 = new_n701 & new_n1363;
  assign new_n2443 = new_n2442 ^ new_n2441;
  assign new_n2444 = n83 & new_n700;
  assign new_n2445 = n81 & new_n787;
  assign new_n2446 = new_n2445 ^ new_n2444;
  assign new_n2447 = new_n2446 ^ new_n2443;
  assign new_n2448 = new_n2447 ^ n15;
  assign new_n2449 = new_n2448 ^ new_n2440;
  assign new_n2450 = new_n2312 ^ new_n2300;
  assign new_n2451 = ~new_n2309 & new_n2450;
  assign new_n2452 = new_n2451 ^ new_n2312;
  assign new_n2453 = new_n2452 ^ new_n2449;
  assign new_n2454 = n85 & new_n499;
  assign new_n2455 = ~new_n506 & new_n1694;
  assign new_n2456 = new_n2455 ^ new_n2454;
  assign new_n2457 = ~new_n505 & n86;
  assign new_n2458 = n84 & new_n579;
  assign new_n2459 = new_n2458 ^ new_n2457;
  assign new_n2460 = new_n2459 ^ new_n2456;
  assign new_n2461 = new_n2460 ^ n12;
  assign new_n2462 = new_n2461 ^ new_n2453;
  assign new_n2463 = new_n2325 ^ new_n2313;
  assign new_n2464 = ~new_n2322 & new_n2463;
  assign new_n2465 = new_n2464 ^ new_n2325;
  assign new_n2466 = new_n2465 ^ new_n2462;
  assign new_n2467 = n88 & new_n354;
  assign new_n2468 = new_n349 & new_n2063;
  assign new_n2469 = new_n2468 ^ new_n2467;
  assign new_n2470 = n89 & new_n348;
  assign new_n2471 = n87 & new_n391;
  assign new_n2472 = new_n2471 ^ new_n2470;
  assign new_n2473 = new_n2472 ^ new_n2469;
  assign new_n2474 = new_n2473 ^ n9;
  assign new_n2475 = new_n2474 ^ new_n2466;
  assign new_n2476 = new_n2338 ^ new_n2326;
  assign new_n2477 = ~new_n2335 & new_n2476;
  assign new_n2478 = new_n2477 ^ new_n2338;
  assign new_n2479 = new_n2478 ^ new_n2475;
  assign new_n2480 = n91 & new_n218;
  assign new_n2481 = new_n2077 ^ n92;
  assign new_n2482 = new_n208 & new_n2481;
  assign new_n2483 = new_n2482 ^ new_n2480;
  assign new_n2484 = n92 & new_n207;
  assign new_n2485 = n90 & new_n212;
  assign new_n2486 = new_n2485 ^ new_n2484;
  assign new_n2487 = new_n2486 ^ new_n2483;
  assign new_n2488 = new_n2487 ^ n6;
  assign new_n2489 = new_n2488 ^ new_n2479;
  assign new_n2490 = new_n2352 ^ new_n2339;
  assign new_n2491 = ~new_n2349 & new_n2490;
  assign new_n2492 = new_n2491 ^ new_n2352;
  assign new_n2493 = new_n2492 ^ new_n2489;
  assign new_n2494 = n94 ^ n3;
  assign new_n2495 = ~n93 & n3;
  assign new_n2496 = new_n2495 ^ new_n2494;
  assign new_n2497 = ~n2 & new_n2496;
  assign new_n2498 = new_n2497 ^ new_n2494;
  assign new_n2499 = n94 ^ n93;
  assign new_n2500 = n94 ^ n92;
  assign new_n2501 = ~new_n2207 & ~new_n2500;
  assign new_n2502 = new_n2499 & new_n2501;
  assign new_n2503 = new_n2502 ^ new_n2499;
  assign new_n2504 = ~new_n2503 & new_n155;
  assign new_n2505 = new_n2504 ^ n2;
  assign new_n2506 = new_n2505 ^ n95;
  assign new_n2507 = new_n2506 ^ new_n2498;
  assign new_n2508 = ~n1 & new_n2507;
  assign new_n2509 = new_n2508 ^ new_n2506;
  assign new_n2510 = new_n2509 ^ new_n2493;
  assign new_n2511 = new_n2372 ^ new_n2353;
  assign new_n2512 = ~new_n2369 & new_n2511;
  assign new_n2513 = new_n2512 ^ new_n2372;
  assign new_n2514 = new_n2513 ^ new_n2510;
  assign new_n2515 = n71 & new_n1874;
  assign new_n2516 = ~new_n459 & new_n1864;
  assign new_n2517 = new_n2516 ^ new_n2515;
  assign new_n2518 = n72 & new_n1863;
  assign new_n2519 = n70 & new_n1868;
  assign new_n2520 = new_n2519 ^ new_n2518;
  assign new_n2521 = new_n2520 ^ new_n2517;
  assign new_n2522 = new_n2521 ^ n27;
  assign new_n2523 = new_n2400 ^ new_n2381;
  assign new_n2524 = ~new_n2397 & new_n2523;
  assign new_n2525 = new_n2524 ^ new_n2400;
  assign new_n2526 = new_n2525 ^ new_n2522;
  assign new_n2527 = ~new_n2249 & ~new_n2383;
  assign new_n2528 = ~new_n2527 & new_n2395;
  assign new_n2529 = n68 & new_n2246;
  assign new_n2530 = ~new_n304 & new_n2241;
  assign new_n2531 = new_n2530 ^ new_n2529;
  assign new_n2532 = n69 & new_n2240;
  assign new_n2533 = n67 & new_n2391;
  assign new_n2534 = new_n2533 ^ new_n2532;
  assign new_n2535 = new_n2534 ^ new_n2531;
  assign new_n2536 = new_n2535 ^ n30;
  assign new_n2537 = n66 ^ n31;
  assign new_n2538 = ~new_n2537 & new_n2382;
  assign new_n2539 = new_n2538 ^ n30;
  assign new_n2540 = new_n2539 ^ n32;
  assign new_n2541 = ~n30 & ~n31;
  assign new_n2542 = new_n2541 ^ new_n2382;
  assign new_n2543 = new_n2542 ^ n32;
  assign new_n2544 = ~n65 & ~new_n2543;
  assign new_n2545 = new_n2544 ^ new_n2540;
  assign new_n2546 = new_n2545 ^ new_n2536;
  assign new_n2547 = new_n2546 ^ new_n2528;
  assign new_n2548 = new_n2547 ^ new_n2526;
  assign new_n2549 = ~new_n1506 & n74;
  assign new_n2550 = new_n660 & new_n1501;
  assign new_n2551 = new_n2550 ^ new_n2549;
  assign new_n2552 = n75 & new_n1500;
  assign new_n2553 = n73 & new_n1512;
  assign new_n2554 = new_n2553 ^ new_n2552;
  assign new_n2555 = new_n2554 ^ new_n2551;
  assign new_n2556 = new_n2555 ^ n24;
  assign new_n2557 = new_n2556 ^ new_n2548;
  assign new_n2558 = new_n2413 ^ new_n2401;
  assign new_n2559 = ~new_n2410 & new_n2558;
  assign new_n2560 = new_n2559 ^ new_n2413;
  assign new_n2561 = new_n2560 ^ new_n2557;
  assign new_n2562 = ~new_n1198 & n77;
  assign new_n2563 = ~new_n891 & new_n1193;
  assign new_n2564 = new_n2563 ^ new_n2562;
  assign new_n2565 = n78 & new_n1192;
  assign new_n2566 = n76 & new_n1204;
  assign new_n2567 = new_n2566 ^ new_n2565;
  assign new_n2568 = new_n2567 ^ new_n2564;
  assign new_n2569 = new_n2568 ^ n21;
  assign new_n2570 = new_n2569 ^ new_n2561;
  assign new_n2571 = new_n2426 ^ new_n2414;
  assign new_n2572 = ~new_n2423 & new_n2571;
  assign new_n2573 = new_n2572 ^ new_n2426;
  assign new_n2574 = new_n2573 ^ new_n2570;
  assign new_n2575 = ~new_n930 & n80;
  assign new_n2576 = new_n925 & new_n1161;
  assign new_n2577 = new_n2576 ^ new_n2575;
  assign new_n2578 = n81 & new_n924;
  assign new_n2579 = n79 & new_n936;
  assign new_n2580 = new_n2579 ^ new_n2578;
  assign new_n2581 = new_n2580 ^ new_n2577;
  assign new_n2582 = new_n2581 ^ n18;
  assign new_n2583 = new_n2582 ^ new_n2574;
  assign new_n2584 = new_n2439 ^ new_n2427;
  assign new_n2585 = ~new_n2436 & new_n2584;
  assign new_n2586 = new_n2585 ^ new_n2439;
  assign new_n2587 = new_n2586 ^ new_n2583;
  assign new_n2588 = n83 & new_n707;
  assign new_n2589 = new_n701 & new_n1468;
  assign new_n2590 = new_n2589 ^ new_n2588;
  assign new_n2591 = n84 & new_n700;
  assign new_n2592 = n82 & new_n787;
  assign new_n2593 = new_n2592 ^ new_n2591;
  assign new_n2594 = new_n2593 ^ new_n2590;
  assign new_n2595 = new_n2594 ^ n15;
  assign new_n2596 = new_n2595 ^ new_n2587;
  assign new_n2597 = new_n2452 ^ new_n2440;
  assign new_n2598 = ~new_n2449 & new_n2597;
  assign new_n2599 = new_n2598 ^ new_n2452;
  assign new_n2600 = new_n2599 ^ new_n2596;
  assign new_n2601 = n86 & new_n499;
  assign new_n2602 = ~new_n506 & new_n1811;
  assign new_n2603 = new_n2602 ^ new_n2601;
  assign new_n2604 = ~new_n505 & n87;
  assign new_n2605 = n85 & new_n579;
  assign new_n2606 = new_n2605 ^ new_n2604;
  assign new_n2607 = new_n2606 ^ new_n2603;
  assign new_n2608 = new_n2607 ^ n12;
  assign new_n2609 = new_n2608 ^ new_n2600;
  assign new_n2610 = new_n2465 ^ new_n2453;
  assign new_n2611 = ~new_n2462 & new_n2610;
  assign new_n2612 = new_n2611 ^ new_n2465;
  assign new_n2613 = new_n2612 ^ new_n2609;
  assign new_n2614 = n89 & new_n354;
  assign new_n2615 = new_n349 & new_n2193;
  assign new_n2616 = new_n2615 ^ new_n2614;
  assign new_n2617 = n90 & new_n348;
  assign new_n2618 = n88 & new_n391;
  assign new_n2619 = new_n2618 ^ new_n2617;
  assign new_n2620 = new_n2619 ^ new_n2616;
  assign new_n2621 = new_n2620 ^ n9;
  assign new_n2622 = new_n2621 ^ new_n2613;
  assign new_n2623 = new_n2478 ^ new_n2466;
  assign new_n2624 = ~new_n2475 & new_n2623;
  assign new_n2625 = new_n2624 ^ new_n2478;
  assign new_n2626 = new_n2625 ^ new_n2622;
  assign new_n2627 = n92 & new_n218;
  assign new_n2628 = new_n2207 ^ n93;
  assign new_n2629 = new_n208 & new_n2628;
  assign new_n2630 = new_n2629 ^ new_n2627;
  assign new_n2631 = n93 & new_n207;
  assign new_n2632 = n91 & new_n212;
  assign new_n2633 = new_n2632 ^ new_n2631;
  assign new_n2634 = new_n2633 ^ new_n2630;
  assign new_n2635 = new_n2634 ^ n6;
  assign new_n2636 = new_n2635 ^ new_n2626;
  assign new_n2637 = new_n2492 ^ new_n2479;
  assign new_n2638 = ~new_n2489 & new_n2637;
  assign new_n2639 = new_n2638 ^ new_n2492;
  assign new_n2640 = new_n2639 ^ new_n2636;
  assign new_n2641 = n95 ^ n94;
  assign new_n2642 = ~new_n2503 & new_n2641;
  assign new_n2643 = ~new_n2642 & new_n155;
  assign new_n2644 = new_n2643 ^ n2;
  assign new_n2645 = new_n2644 ^ n96;
  assign new_n2646 = n95 ^ n3;
  assign new_n2647 = ~n94 & ~new_n2494;
  assign new_n2648 = new_n2647 ^ new_n2646;
  assign new_n2649 = new_n2648 ^ n94;
  assign new_n2650 = ~new_n2649 & new_n241;
  assign new_n2651 = new_n2650 ^ new_n2647;
  assign new_n2652 = new_n2651 ^ n94;
  assign new_n2653 = new_n2652 ^ new_n2645;
  assign new_n2654 = ~n1 & ~new_n2653;
  assign new_n2655 = new_n2654 ^ new_n2645;
  assign new_n2656 = new_n2655 ^ new_n2640;
  assign new_n2657 = new_n2513 ^ new_n2493;
  assign new_n2658 = ~new_n2510 & new_n2657;
  assign new_n2659 = new_n2658 ^ new_n2513;
  assign new_n2660 = new_n2659 ^ new_n2656;
  assign new_n2661 = n33 ^ n32;
  assign new_n2662 = ~new_n2382 & n33;
  assign new_n2663 = new_n2662 ^ new_n2542;
  assign new_n2664 = ~new_n2663 & new_n2661;
  assign new_n2665 = n65 & new_n2664;
  assign new_n2666 = ~new_n2661 & new_n2382;
  assign new_n2667 = new_n2666 ^ new_n2382;
  assign new_n2668 = ~new_n151 & new_n2667;
  assign new_n2669 = n67 & new_n2382;
  assign new_n2670 = new_n2669 ^ new_n2668;
  assign new_n2671 = ~new_n2382 & n32;
  assign new_n2672 = new_n2671 ^ new_n2542;
  assign new_n2673 = ~new_n2672 & n66;
  assign new_n2674 = new_n2673 ^ new_n2670;
  assign new_n2675 = new_n2674 ^ n33;
  assign new_n2676 = new_n2675 ^ new_n2665;
  assign new_n2677 = ~new_n2383 & ~new_n2545;
  assign new_n2678 = n33 & new_n2677;
  assign new_n2679 = new_n2678 ^ new_n2676;
  assign new_n2680 = n69 & new_n2246;
  assign new_n2681 = ~new_n339 & new_n2241;
  assign new_n2682 = new_n2681 ^ new_n2680;
  assign new_n2683 = n70 & new_n2240;
  assign new_n2684 = n68 & new_n2391;
  assign new_n2685 = new_n2684 ^ new_n2683;
  assign new_n2686 = new_n2685 ^ new_n2682;
  assign new_n2687 = new_n2686 ^ n30;
  assign new_n2688 = new_n2687 ^ new_n2679;
  assign new_n2689 = new_n2536 ^ new_n2528;
  assign new_n2690 = ~new_n2546 & new_n2689;
  assign new_n2691 = new_n2690 ^ new_n2528;
  assign new_n2692 = new_n2691 ^ new_n2688;
  assign new_n2693 = n72 & new_n1874;
  assign new_n2694 = new_n534 & new_n1864;
  assign new_n2695 = new_n2694 ^ new_n2693;
  assign new_n2696 = n73 & new_n1863;
  assign new_n2697 = n71 & new_n1868;
  assign new_n2698 = new_n2697 ^ new_n2696;
  assign new_n2699 = new_n2698 ^ new_n2695;
  assign new_n2700 = new_n2699 ^ n27;
  assign new_n2701 = new_n2700 ^ new_n2692;
  assign new_n2702 = new_n2547 ^ new_n2522;
  assign new_n2703 = ~new_n2702 & new_n2526;
  assign new_n2704 = new_n2703 ^ new_n2525;
  assign new_n2705 = new_n2704 ^ new_n2701;
  assign new_n2706 = ~new_n1506 & n75;
  assign new_n2707 = ~new_n737 & new_n1501;
  assign new_n2708 = new_n2707 ^ new_n2706;
  assign new_n2709 = n76 & new_n1500;
  assign new_n2710 = n74 & new_n1512;
  assign new_n2711 = new_n2710 ^ new_n2709;
  assign new_n2712 = new_n2711 ^ new_n2708;
  assign new_n2713 = new_n2712 ^ n24;
  assign new_n2714 = new_n2713 ^ new_n2705;
  assign new_n2715 = new_n2560 ^ new_n2548;
  assign new_n2716 = ~new_n2557 & new_n2715;
  assign new_n2717 = new_n2716 ^ new_n2560;
  assign new_n2718 = new_n2717 ^ new_n2714;
  assign new_n2719 = ~new_n1198 & n78;
  assign new_n2720 = ~new_n982 & new_n1193;
  assign new_n2721 = new_n2720 ^ new_n2719;
  assign new_n2722 = n79 & new_n1192;
  assign new_n2723 = n77 & new_n1204;
  assign new_n2724 = new_n2723 ^ new_n2722;
  assign new_n2725 = new_n2724 ^ new_n2721;
  assign new_n2726 = new_n2725 ^ n21;
  assign new_n2727 = new_n2726 ^ new_n2718;
  assign new_n2728 = new_n2573 ^ new_n2561;
  assign new_n2729 = ~new_n2570 & new_n2728;
  assign new_n2730 = new_n2729 ^ new_n2573;
  assign new_n2731 = new_n2730 ^ new_n2727;
  assign new_n2732 = ~new_n930 & n81;
  assign new_n2733 = new_n925 & new_n1263;
  assign new_n2734 = new_n2733 ^ new_n2732;
  assign new_n2735 = n82 & new_n924;
  assign new_n2736 = n80 & new_n936;
  assign new_n2737 = new_n2736 ^ new_n2735;
  assign new_n2738 = new_n2737 ^ new_n2734;
  assign new_n2739 = new_n2738 ^ n18;
  assign new_n2740 = new_n2739 ^ new_n2731;
  assign new_n2741 = new_n2586 ^ new_n2574;
  assign new_n2742 = ~new_n2583 & new_n2741;
  assign new_n2743 = new_n2742 ^ new_n2586;
  assign new_n2744 = new_n2743 ^ new_n2740;
  assign new_n2745 = n84 & new_n707;
  assign new_n2746 = new_n701 & new_n1584;
  assign new_n2747 = new_n2746 ^ new_n2745;
  assign new_n2748 = n85 & new_n700;
  assign new_n2749 = n83 & new_n787;
  assign new_n2750 = new_n2749 ^ new_n2748;
  assign new_n2751 = new_n2750 ^ new_n2747;
  assign new_n2752 = new_n2751 ^ n15;
  assign new_n2753 = new_n2752 ^ new_n2744;
  assign new_n2754 = new_n2599 ^ new_n2587;
  assign new_n2755 = ~new_n2596 & new_n2754;
  assign new_n2756 = new_n2755 ^ new_n2599;
  assign new_n2757 = new_n2756 ^ new_n2753;
  assign new_n2758 = n87 & new_n499;
  assign new_n2759 = ~new_n506 & new_n1940;
  assign new_n2760 = new_n2759 ^ new_n2758;
  assign new_n2761 = ~new_n505 & n88;
  assign new_n2762 = n86 & new_n579;
  assign new_n2763 = new_n2762 ^ new_n2761;
  assign new_n2764 = new_n2763 ^ new_n2760;
  assign new_n2765 = new_n2764 ^ n12;
  assign new_n2766 = new_n2765 ^ new_n2757;
  assign new_n2767 = new_n2612 ^ new_n2600;
  assign new_n2768 = ~new_n2609 & new_n2767;
  assign new_n2769 = new_n2768 ^ new_n2612;
  assign new_n2770 = new_n2769 ^ new_n2766;
  assign new_n2771 = n90 & new_n354;
  assign new_n2772 = new_n349 & new_n2341;
  assign new_n2773 = new_n2772 ^ new_n2771;
  assign new_n2774 = n91 & new_n348;
  assign new_n2775 = n89 & new_n391;
  assign new_n2776 = new_n2775 ^ new_n2774;
  assign new_n2777 = new_n2776 ^ new_n2773;
  assign new_n2778 = new_n2777 ^ n9;
  assign new_n2779 = new_n2778 ^ new_n2770;
  assign new_n2780 = new_n2625 ^ new_n2613;
  assign new_n2781 = ~new_n2622 & new_n2780;
  assign new_n2782 = new_n2781 ^ new_n2625;
  assign new_n2783 = new_n2782 ^ new_n2779;
  assign new_n2784 = n93 & new_n218;
  assign new_n2785 = new_n2355 ^ n94;
  assign new_n2786 = new_n208 & new_n2785;
  assign new_n2787 = new_n2786 ^ new_n2784;
  assign new_n2788 = n94 & new_n207;
  assign new_n2789 = n92 & new_n212;
  assign new_n2790 = new_n2789 ^ new_n2788;
  assign new_n2791 = new_n2790 ^ new_n2787;
  assign new_n2792 = new_n2791 ^ n6;
  assign new_n2793 = new_n2792 ^ new_n2783;
  assign new_n2794 = new_n2639 ^ new_n2626;
  assign new_n2795 = ~new_n2636 & new_n2794;
  assign new_n2796 = new_n2795 ^ new_n2639;
  assign new_n2797 = new_n2796 ^ new_n2793;
  assign new_n2798 = n96 ^ n95;
  assign new_n2799 = ~new_n2642 & new_n2798;
  assign new_n2800 = ~new_n2799 & new_n155;
  assign new_n2801 = new_n2800 ^ n2;
  assign new_n2802 = new_n2801 ^ n97;
  assign new_n2803 = n96 ^ n3;
  assign new_n2804 = ~n95 & n3;
  assign new_n2805 = new_n2804 ^ new_n2803;
  assign new_n2806 = ~n2 & new_n2805;
  assign new_n2807 = new_n2806 ^ new_n2803;
  assign new_n2808 = new_n2807 ^ new_n2802;
  assign new_n2809 = ~n1 & new_n2808;
  assign new_n2810 = new_n2809 ^ new_n2802;
  assign new_n2811 = new_n2810 ^ new_n2797;
  assign new_n2812 = new_n2659 ^ new_n2640;
  assign new_n2813 = ~new_n2656 & new_n2812;
  assign new_n2814 = new_n2813 ^ new_n2659;
  assign new_n2815 = new_n2814 ^ new_n2811;
  assign new_n2816 = new_n2676 & new_n2678;
  assign new_n2817 = ~new_n259 & new_n2667;
  assign new_n2818 = ~new_n2672 & n67;
  assign new_n2819 = new_n2818 ^ new_n2817;
  assign new_n2820 = n68 & new_n2666;
  assign new_n2821 = n66 & new_n2664;
  assign new_n2822 = new_n2821 ^ new_n2820;
  assign new_n2823 = new_n2822 ^ new_n2819;
  assign new_n2824 = new_n2823 ^ n33;
  assign new_n2825 = n34 ^ n33;
  assign new_n2826 = n65 & new_n2825;
  assign new_n2827 = new_n2826 ^ new_n2824;
  assign new_n2828 = new_n2827 ^ new_n2816;
  assign new_n2829 = n70 & new_n2246;
  assign new_n2830 = ~new_n402 & new_n2241;
  assign new_n2831 = new_n2830 ^ new_n2829;
  assign new_n2832 = n71 & new_n2240;
  assign new_n2833 = n69 & new_n2391;
  assign new_n2834 = new_n2833 ^ new_n2832;
  assign new_n2835 = new_n2834 ^ new_n2831;
  assign new_n2836 = new_n2835 ^ n30;
  assign new_n2837 = new_n2836 ^ new_n2828;
  assign new_n2838 = new_n2691 ^ new_n2679;
  assign new_n2839 = ~new_n2688 & new_n2838;
  assign new_n2840 = new_n2839 ^ new_n2691;
  assign new_n2841 = new_n2840 ^ new_n2837;
  assign new_n2842 = n73 & new_n1874;
  assign new_n2843 = new_n595 & new_n1864;
  assign new_n2844 = new_n2843 ^ new_n2842;
  assign new_n2845 = n74 & new_n1863;
  assign new_n2846 = n72 & new_n1868;
  assign new_n2847 = new_n2846 ^ new_n2845;
  assign new_n2848 = new_n2847 ^ new_n2844;
  assign new_n2849 = new_n2848 ^ n27;
  assign new_n2850 = new_n2849 ^ new_n2841;
  assign new_n2851 = new_n2704 ^ new_n2692;
  assign new_n2852 = ~new_n2701 & new_n2851;
  assign new_n2853 = new_n2852 ^ new_n2704;
  assign new_n2854 = new_n2853 ^ new_n2850;
  assign new_n2855 = ~new_n1506 & n76;
  assign new_n2856 = ~new_n812 & new_n1501;
  assign new_n2857 = new_n2856 ^ new_n2855;
  assign new_n2858 = n77 & new_n1500;
  assign new_n2859 = n75 & new_n1512;
  assign new_n2860 = new_n2859 ^ new_n2858;
  assign new_n2861 = new_n2860 ^ new_n2857;
  assign new_n2862 = new_n2861 ^ n24;
  assign new_n2863 = new_n2862 ^ new_n2854;
  assign new_n2864 = new_n2717 ^ new_n2705;
  assign new_n2865 = ~new_n2714 & new_n2864;
  assign new_n2866 = new_n2865 ^ new_n2717;
  assign new_n2867 = new_n2866 ^ new_n2863;
  assign new_n2868 = ~new_n1198 & n79;
  assign new_n2869 = new_n1069 & new_n1193;
  assign new_n2870 = new_n2869 ^ new_n2868;
  assign new_n2871 = n80 & new_n1192;
  assign new_n2872 = n78 & new_n1204;
  assign new_n2873 = new_n2872 ^ new_n2871;
  assign new_n2874 = new_n2873 ^ new_n2870;
  assign new_n2875 = new_n2874 ^ n21;
  assign new_n2876 = new_n2875 ^ new_n2867;
  assign new_n2877 = new_n2730 ^ new_n2718;
  assign new_n2878 = ~new_n2727 & new_n2877;
  assign new_n2879 = new_n2878 ^ new_n2730;
  assign new_n2880 = new_n2879 ^ new_n2876;
  assign new_n2881 = ~new_n930 & n82;
  assign new_n2882 = new_n925 & new_n1363;
  assign new_n2883 = new_n2882 ^ new_n2881;
  assign new_n2884 = n83 & new_n924;
  assign new_n2885 = n81 & new_n936;
  assign new_n2886 = new_n2885 ^ new_n2884;
  assign new_n2887 = new_n2886 ^ new_n2883;
  assign new_n2888 = new_n2887 ^ n18;
  assign new_n2889 = new_n2888 ^ new_n2880;
  assign new_n2890 = new_n2743 ^ new_n2731;
  assign new_n2891 = ~new_n2740 & new_n2890;
  assign new_n2892 = new_n2891 ^ new_n2743;
  assign new_n2893 = new_n2892 ^ new_n2889;
  assign new_n2894 = n85 & new_n707;
  assign new_n2895 = new_n701 & new_n1694;
  assign new_n2896 = new_n2895 ^ new_n2894;
  assign new_n2897 = n86 & new_n700;
  assign new_n2898 = n84 & new_n787;
  assign new_n2899 = new_n2898 ^ new_n2897;
  assign new_n2900 = new_n2899 ^ new_n2896;
  assign new_n2901 = new_n2900 ^ n15;
  assign new_n2902 = new_n2901 ^ new_n2893;
  assign new_n2903 = new_n2756 ^ new_n2744;
  assign new_n2904 = ~new_n2753 & new_n2903;
  assign new_n2905 = new_n2904 ^ new_n2756;
  assign new_n2906 = new_n2905 ^ new_n2902;
  assign new_n2907 = n88 & new_n499;
  assign new_n2908 = ~new_n506 & new_n2063;
  assign new_n2909 = new_n2908 ^ new_n2907;
  assign new_n2910 = ~new_n505 & n89;
  assign new_n2911 = n87 & new_n579;
  assign new_n2912 = new_n2911 ^ new_n2910;
  assign new_n2913 = new_n2912 ^ new_n2909;
  assign new_n2914 = new_n2913 ^ n12;
  assign new_n2915 = new_n2914 ^ new_n2906;
  assign new_n2916 = new_n2769 ^ new_n2757;
  assign new_n2917 = ~new_n2766 & new_n2916;
  assign new_n2918 = new_n2917 ^ new_n2769;
  assign new_n2919 = new_n2918 ^ new_n2915;
  assign new_n2920 = n91 & new_n354;
  assign new_n2921 = new_n349 & new_n2481;
  assign new_n2922 = new_n2921 ^ new_n2920;
  assign new_n2923 = n92 & new_n348;
  assign new_n2924 = n90 & new_n391;
  assign new_n2925 = new_n2924 ^ new_n2923;
  assign new_n2926 = new_n2925 ^ new_n2922;
  assign new_n2927 = new_n2926 ^ n9;
  assign new_n2928 = new_n2927 ^ new_n2919;
  assign new_n2929 = new_n2782 ^ new_n2770;
  assign new_n2930 = ~new_n2779 & new_n2929;
  assign new_n2931 = new_n2930 ^ new_n2782;
  assign new_n2932 = new_n2931 ^ new_n2928;
  assign new_n2933 = n94 & new_n218;
  assign new_n2934 = new_n2503 ^ n95;
  assign new_n2935 = new_n208 & new_n2934;
  assign new_n2936 = new_n2935 ^ new_n2933;
  assign new_n2937 = n95 & new_n207;
  assign new_n2938 = n93 & new_n212;
  assign new_n2939 = new_n2938 ^ new_n2937;
  assign new_n2940 = new_n2939 ^ new_n2936;
  assign new_n2941 = new_n2940 ^ n6;
  assign new_n2942 = new_n2941 ^ new_n2932;
  assign new_n2943 = new_n2796 ^ new_n2783;
  assign new_n2944 = ~new_n2793 & new_n2943;
  assign new_n2945 = new_n2944 ^ new_n2796;
  assign new_n2946 = new_n2945 ^ new_n2942;
  assign new_n2947 = n97 ^ n96;
  assign new_n2948 = n97 ^ n95;
  assign new_n2949 = ~new_n2948 & new_n2642;
  assign new_n2950 = new_n2949 ^ n95;
  assign new_n2951 = new_n2950 ^ n97;
  assign new_n2952 = new_n2947 & new_n2951;
  assign new_n2953 = ~new_n2952 & new_n155;
  assign new_n2954 = new_n2953 ^ n2;
  assign new_n2955 = new_n2954 ^ n98;
  assign new_n2956 = n97 ^ n3;
  assign new_n2957 = ~n96 & n3;
  assign new_n2958 = new_n2957 ^ new_n2956;
  assign new_n2959 = ~n2 & new_n2958;
  assign new_n2960 = new_n2959 ^ new_n2956;
  assign new_n2961 = new_n2960 ^ new_n2955;
  assign new_n2962 = ~n1 & new_n2961;
  assign new_n2963 = new_n2962 ^ new_n2955;
  assign new_n2964 = new_n2963 ^ new_n2946;
  assign new_n2965 = new_n2814 ^ new_n2797;
  assign new_n2966 = ~new_n2811 & new_n2965;
  assign new_n2967 = new_n2966 ^ new_n2814;
  assign new_n2968 = new_n2967 ^ new_n2964;
  assign new_n2969 = ~new_n2816 & ~new_n2826;
  assign new_n2970 = ~new_n2969 & new_n2824;
  assign new_n2971 = ~n33 & ~n34;
  assign new_n2972 = new_n2971 ^ new_n2825;
  assign new_n2973 = new_n2972 ^ n35;
  assign new_n2974 = ~n65 & ~new_n2973;
  assign new_n2975 = n66 ^ n34;
  assign new_n2976 = ~new_n2975 & new_n2825;
  assign new_n2977 = new_n2976 ^ n33;
  assign new_n2978 = new_n2977 ^ n35;
  assign new_n2979 = new_n2978 ^ new_n2974;
  assign new_n2980 = ~new_n2672 & n68;
  assign new_n2981 = ~new_n304 & new_n2667;
  assign new_n2982 = new_n2981 ^ new_n2980;
  assign new_n2983 = n69 & new_n2666;
  assign new_n2984 = n67 & new_n2664;
  assign new_n2985 = new_n2984 ^ new_n2983;
  assign new_n2986 = new_n2985 ^ new_n2982;
  assign new_n2987 = new_n2986 ^ n33;
  assign new_n2988 = new_n2987 ^ new_n2979;
  assign new_n2989 = new_n2988 ^ new_n2970;
  assign new_n2990 = n71 & new_n2246;
  assign new_n2991 = ~new_n459 & new_n2241;
  assign new_n2992 = new_n2991 ^ new_n2990;
  assign new_n2993 = n72 & new_n2240;
  assign new_n2994 = n70 & new_n2391;
  assign new_n2995 = new_n2994 ^ new_n2993;
  assign new_n2996 = new_n2995 ^ new_n2992;
  assign new_n2997 = new_n2996 ^ n30;
  assign new_n2998 = new_n2997 ^ new_n2989;
  assign new_n2999 = new_n2840 ^ new_n2828;
  assign new_n3000 = ~new_n2837 & new_n2999;
  assign new_n3001 = new_n3000 ^ new_n2840;
  assign new_n3002 = new_n3001 ^ new_n2998;
  assign new_n3003 = n74 & new_n1874;
  assign new_n3004 = new_n660 & new_n1864;
  assign new_n3005 = new_n3004 ^ new_n3003;
  assign new_n3006 = n75 & new_n1863;
  assign new_n3007 = n73 & new_n1868;
  assign new_n3008 = new_n3007 ^ new_n3006;
  assign new_n3009 = new_n3008 ^ new_n3005;
  assign new_n3010 = new_n3009 ^ n27;
  assign new_n3011 = new_n3010 ^ new_n3002;
  assign new_n3012 = new_n2853 ^ new_n2841;
  assign new_n3013 = ~new_n2850 & new_n3012;
  assign new_n3014 = new_n3013 ^ new_n2853;
  assign new_n3015 = new_n3014 ^ new_n3011;
  assign new_n3016 = ~new_n1506 & n77;
  assign new_n3017 = ~new_n891 & new_n1501;
  assign new_n3018 = new_n3017 ^ new_n3016;
  assign new_n3019 = n78 & new_n1500;
  assign new_n3020 = n76 & new_n1512;
  assign new_n3021 = new_n3020 ^ new_n3019;
  assign new_n3022 = new_n3021 ^ new_n3018;
  assign new_n3023 = new_n3022 ^ n24;
  assign new_n3024 = new_n3023 ^ new_n3015;
  assign new_n3025 = new_n2866 ^ new_n2854;
  assign new_n3026 = ~new_n2863 & new_n3025;
  assign new_n3027 = new_n3026 ^ new_n2866;
  assign new_n3028 = new_n3027 ^ new_n3024;
  assign new_n3029 = ~new_n1198 & n80;
  assign new_n3030 = new_n1161 & new_n1193;
  assign new_n3031 = new_n3030 ^ new_n3029;
  assign new_n3032 = n81 & new_n1192;
  assign new_n3033 = n79 & new_n1204;
  assign new_n3034 = new_n3033 ^ new_n3032;
  assign new_n3035 = new_n3034 ^ new_n3031;
  assign new_n3036 = new_n3035 ^ n21;
  assign new_n3037 = new_n3036 ^ new_n3028;
  assign new_n3038 = new_n2879 ^ new_n2867;
  assign new_n3039 = ~new_n2876 & new_n3038;
  assign new_n3040 = new_n3039 ^ new_n2879;
  assign new_n3041 = new_n3040 ^ new_n3037;
  assign new_n3042 = ~new_n930 & n83;
  assign new_n3043 = new_n925 & new_n1468;
  assign new_n3044 = new_n3043 ^ new_n3042;
  assign new_n3045 = n84 & new_n924;
  assign new_n3046 = n82 & new_n936;
  assign new_n3047 = new_n3046 ^ new_n3045;
  assign new_n3048 = new_n3047 ^ new_n3044;
  assign new_n3049 = new_n3048 ^ n18;
  assign new_n3050 = new_n3049 ^ new_n3041;
  assign new_n3051 = new_n2892 ^ new_n2880;
  assign new_n3052 = ~new_n2889 & new_n3051;
  assign new_n3053 = new_n3052 ^ new_n2892;
  assign new_n3054 = new_n3053 ^ new_n3050;
  assign new_n3055 = n86 & new_n707;
  assign new_n3056 = new_n701 & new_n1811;
  assign new_n3057 = new_n3056 ^ new_n3055;
  assign new_n3058 = n87 & new_n700;
  assign new_n3059 = n85 & new_n787;
  assign new_n3060 = new_n3059 ^ new_n3058;
  assign new_n3061 = new_n3060 ^ new_n3057;
  assign new_n3062 = new_n3061 ^ n15;
  assign new_n3063 = new_n3062 ^ new_n3054;
  assign new_n3064 = new_n2905 ^ new_n2893;
  assign new_n3065 = ~new_n2902 & new_n3064;
  assign new_n3066 = new_n3065 ^ new_n2905;
  assign new_n3067 = new_n3066 ^ new_n3063;
  assign new_n3068 = n89 & new_n499;
  assign new_n3069 = ~new_n506 & new_n2193;
  assign new_n3070 = new_n3069 ^ new_n3068;
  assign new_n3071 = ~new_n505 & n90;
  assign new_n3072 = n88 & new_n579;
  assign new_n3073 = new_n3072 ^ new_n3071;
  assign new_n3074 = new_n3073 ^ new_n3070;
  assign new_n3075 = new_n3074 ^ n12;
  assign new_n3076 = new_n3075 ^ new_n3067;
  assign new_n3077 = new_n2918 ^ new_n2906;
  assign new_n3078 = ~new_n2915 & new_n3077;
  assign new_n3079 = new_n3078 ^ new_n2918;
  assign new_n3080 = new_n3079 ^ new_n3076;
  assign new_n3081 = n92 & new_n354;
  assign new_n3082 = new_n349 & new_n2628;
  assign new_n3083 = new_n3082 ^ new_n3081;
  assign new_n3084 = n93 & new_n348;
  assign new_n3085 = n91 & new_n391;
  assign new_n3086 = new_n3085 ^ new_n3084;
  assign new_n3087 = new_n3086 ^ new_n3083;
  assign new_n3088 = new_n3087 ^ n9;
  assign new_n3089 = new_n3088 ^ new_n3080;
  assign new_n3090 = new_n2931 ^ new_n2919;
  assign new_n3091 = ~new_n2928 & new_n3090;
  assign new_n3092 = new_n3091 ^ new_n2931;
  assign new_n3093 = new_n3092 ^ new_n3089;
  assign new_n3094 = n95 & new_n218;
  assign new_n3095 = new_n2642 ^ n96;
  assign new_n3096 = new_n208 & new_n3095;
  assign new_n3097 = new_n3096 ^ new_n3094;
  assign new_n3098 = n96 & new_n207;
  assign new_n3099 = n94 & new_n212;
  assign new_n3100 = new_n3099 ^ new_n3098;
  assign new_n3101 = new_n3100 ^ new_n3097;
  assign new_n3102 = new_n3101 ^ n6;
  assign new_n3103 = new_n3102 ^ new_n3093;
  assign new_n3104 = new_n2945 ^ new_n2932;
  assign new_n3105 = ~new_n2942 & new_n3104;
  assign new_n3106 = new_n3105 ^ new_n2945;
  assign new_n3107 = new_n3106 ^ new_n3103;
  assign new_n3108 = n97 & new_n180;
  assign new_n3109 = n2 & n98;
  assign new_n3110 = new_n3109 ^ new_n3108;
  assign new_n3111 = new_n3110 ^ n3;
  assign new_n3112 = n98 ^ n97;
  assign new_n3113 = n98 ^ n95;
  assign new_n3114 = new_n3113 ^ new_n2642;
  assign new_n3115 = new_n3113 ^ new_n2947;
  assign new_n3116 = new_n3113 & new_n3115;
  assign new_n3117 = new_n3116 ^ new_n3113;
  assign new_n3118 = ~new_n3114 & new_n3117;
  assign new_n3119 = new_n3118 ^ new_n3116;
  assign new_n3120 = new_n3119 ^ new_n3113;
  assign new_n3121 = new_n3120 ^ new_n2947;
  assign new_n3122 = new_n3112 & new_n3121;
  assign new_n3123 = new_n3122 ^ n97;
  assign new_n3124 = new_n3123 ^ n98;
  assign new_n3125 = ~new_n3124 & new_n155;
  assign new_n3126 = new_n3125 ^ n2;
  assign new_n3127 = new_n3126 ^ n99;
  assign new_n3128 = new_n3127 ^ new_n3111;
  assign new_n3129 = ~n1 & new_n3128;
  assign new_n3130 = new_n3129 ^ new_n3127;
  assign new_n3131 = new_n3130 ^ new_n3107;
  assign new_n3132 = new_n2967 ^ new_n2946;
  assign new_n3133 = ~new_n2964 & new_n3132;
  assign new_n3134 = new_n3133 ^ new_n2967;
  assign new_n3135 = new_n3134 ^ new_n3131;
  assign new_n3136 = n36 ^ n35;
  assign new_n3137 = ~new_n3136 & new_n2825;
  assign new_n3138 = new_n3137 ^ new_n2825;
  assign new_n3139 = ~new_n151 & new_n3138;
  assign new_n3140 = n67 & new_n2825;
  assign new_n3141 = new_n3140 ^ new_n3139;
  assign new_n3142 = ~new_n2825 & n35;
  assign new_n3143 = new_n3142 ^ new_n2972;
  assign new_n3144 = ~new_n3143 & n66;
  assign new_n3145 = new_n3144 ^ new_n3141;
  assign new_n3146 = new_n3145 ^ n36;
  assign new_n3147 = ~new_n2825 & n36;
  assign new_n3148 = new_n3147 ^ new_n2972;
  assign new_n3149 = ~new_n3148 & new_n3136;
  assign new_n3150 = n65 & new_n3149;
  assign new_n3151 = new_n3150 ^ new_n3146;
  assign new_n3152 = ~new_n2826 & ~new_n2979;
  assign new_n3153 = n36 & new_n3152;
  assign new_n3154 = new_n3153 ^ new_n3151;
  assign new_n3155 = ~new_n2672 & n69;
  assign new_n3156 = ~new_n339 & new_n2667;
  assign new_n3157 = new_n3156 ^ new_n3155;
  assign new_n3158 = n70 & new_n2666;
  assign new_n3159 = n68 & new_n2664;
  assign new_n3160 = new_n3159 ^ new_n3158;
  assign new_n3161 = new_n3160 ^ new_n3157;
  assign new_n3162 = new_n3161 ^ n33;
  assign new_n3163 = new_n3162 ^ new_n3154;
  assign new_n3164 = new_n2987 ^ new_n2970;
  assign new_n3165 = ~new_n2988 & new_n3164;
  assign new_n3166 = new_n3165 ^ new_n2970;
  assign new_n3167 = new_n3166 ^ new_n3163;
  assign new_n3168 = n72 & new_n2246;
  assign new_n3169 = new_n534 & new_n2241;
  assign new_n3170 = new_n3169 ^ new_n3168;
  assign new_n3171 = n73 & new_n2240;
  assign new_n3172 = n71 & new_n2391;
  assign new_n3173 = new_n3172 ^ new_n3171;
  assign new_n3174 = new_n3173 ^ new_n3170;
  assign new_n3175 = new_n3174 ^ n30;
  assign new_n3176 = new_n3175 ^ new_n3167;
  assign new_n3177 = new_n3001 ^ new_n2989;
  assign new_n3178 = ~new_n2998 & new_n3177;
  assign new_n3179 = new_n3178 ^ new_n3001;
  assign new_n3180 = new_n3179 ^ new_n3176;
  assign new_n3181 = n75 & new_n1874;
  assign new_n3182 = ~new_n737 & new_n1864;
  assign new_n3183 = new_n3182 ^ new_n3181;
  assign new_n3184 = n76 & new_n1863;
  assign new_n3185 = n74 & new_n1868;
  assign new_n3186 = new_n3185 ^ new_n3184;
  assign new_n3187 = new_n3186 ^ new_n3183;
  assign new_n3188 = new_n3187 ^ n27;
  assign new_n3189 = new_n3188 ^ new_n3180;
  assign new_n3190 = new_n3014 ^ new_n3002;
  assign new_n3191 = ~new_n3011 & new_n3190;
  assign new_n3192 = new_n3191 ^ new_n3014;
  assign new_n3193 = new_n3192 ^ new_n3189;
  assign new_n3194 = ~new_n1506 & n78;
  assign new_n3195 = ~new_n982 & new_n1501;
  assign new_n3196 = new_n3195 ^ new_n3194;
  assign new_n3197 = n79 & new_n1500;
  assign new_n3198 = n77 & new_n1512;
  assign new_n3199 = new_n3198 ^ new_n3197;
  assign new_n3200 = new_n3199 ^ new_n3196;
  assign new_n3201 = new_n3200 ^ n24;
  assign new_n3202 = new_n3201 ^ new_n3193;
  assign new_n3203 = new_n3027 ^ new_n3015;
  assign new_n3204 = ~new_n3024 & new_n3203;
  assign new_n3205 = new_n3204 ^ new_n3027;
  assign new_n3206 = new_n3205 ^ new_n3202;
  assign new_n3207 = ~new_n1198 & n81;
  assign new_n3208 = new_n1193 & new_n1263;
  assign new_n3209 = new_n3208 ^ new_n3207;
  assign new_n3210 = n82 & new_n1192;
  assign new_n3211 = n80 & new_n1204;
  assign new_n3212 = new_n3211 ^ new_n3210;
  assign new_n3213 = new_n3212 ^ new_n3209;
  assign new_n3214 = new_n3213 ^ n21;
  assign new_n3215 = new_n3214 ^ new_n3206;
  assign new_n3216 = new_n3040 ^ new_n3028;
  assign new_n3217 = ~new_n3037 & new_n3216;
  assign new_n3218 = new_n3217 ^ new_n3040;
  assign new_n3219 = new_n3218 ^ new_n3215;
  assign new_n3220 = ~new_n930 & n84;
  assign new_n3221 = new_n925 & new_n1584;
  assign new_n3222 = new_n3221 ^ new_n3220;
  assign new_n3223 = n85 & new_n924;
  assign new_n3224 = n83 & new_n936;
  assign new_n3225 = new_n3224 ^ new_n3223;
  assign new_n3226 = new_n3225 ^ new_n3222;
  assign new_n3227 = new_n3226 ^ n18;
  assign new_n3228 = new_n3227 ^ new_n3219;
  assign new_n3229 = new_n3053 ^ new_n3041;
  assign new_n3230 = ~new_n3050 & new_n3229;
  assign new_n3231 = new_n3230 ^ new_n3053;
  assign new_n3232 = new_n3231 ^ new_n3228;
  assign new_n3233 = n87 & new_n707;
  assign new_n3234 = new_n701 & new_n1940;
  assign new_n3235 = new_n3234 ^ new_n3233;
  assign new_n3236 = n88 & new_n700;
  assign new_n3237 = n86 & new_n787;
  assign new_n3238 = new_n3237 ^ new_n3236;
  assign new_n3239 = new_n3238 ^ new_n3235;
  assign new_n3240 = new_n3239 ^ n15;
  assign new_n3241 = new_n3240 ^ new_n3232;
  assign new_n3242 = new_n3066 ^ new_n3054;
  assign new_n3243 = ~new_n3063 & new_n3242;
  assign new_n3244 = new_n3243 ^ new_n3066;
  assign new_n3245 = new_n3244 ^ new_n3241;
  assign new_n3246 = n90 & new_n499;
  assign new_n3247 = ~new_n506 & new_n2341;
  assign new_n3248 = new_n3247 ^ new_n3246;
  assign new_n3249 = ~new_n505 & n91;
  assign new_n3250 = n89 & new_n579;
  assign new_n3251 = new_n3250 ^ new_n3249;
  assign new_n3252 = new_n3251 ^ new_n3248;
  assign new_n3253 = new_n3252 ^ n12;
  assign new_n3254 = new_n3253 ^ new_n3245;
  assign new_n3255 = new_n3079 ^ new_n3067;
  assign new_n3256 = ~new_n3076 & new_n3255;
  assign new_n3257 = new_n3256 ^ new_n3079;
  assign new_n3258 = new_n3257 ^ new_n3254;
  assign new_n3259 = n93 & new_n354;
  assign new_n3260 = new_n349 & new_n2785;
  assign new_n3261 = new_n3260 ^ new_n3259;
  assign new_n3262 = n94 & new_n348;
  assign new_n3263 = n92 & new_n391;
  assign new_n3264 = new_n3263 ^ new_n3262;
  assign new_n3265 = new_n3264 ^ new_n3261;
  assign new_n3266 = new_n3265 ^ n9;
  assign new_n3267 = new_n3266 ^ new_n3258;
  assign new_n3268 = new_n3092 ^ new_n3080;
  assign new_n3269 = ~new_n3089 & new_n3268;
  assign new_n3270 = new_n3269 ^ new_n3092;
  assign new_n3271 = new_n3270 ^ new_n3267;
  assign new_n3272 = n96 & new_n218;
  assign new_n3273 = new_n2799 ^ n97;
  assign new_n3274 = new_n208 & new_n3273;
  assign new_n3275 = new_n3274 ^ new_n3272;
  assign new_n3276 = n97 & new_n207;
  assign new_n3277 = n95 & new_n212;
  assign new_n3278 = new_n3277 ^ new_n3276;
  assign new_n3279 = new_n3278 ^ new_n3275;
  assign new_n3280 = new_n3279 ^ n6;
  assign new_n3281 = new_n3280 ^ new_n3271;
  assign new_n3282 = new_n3106 ^ new_n3093;
  assign new_n3283 = ~new_n3103 & new_n3282;
  assign new_n3284 = new_n3283 ^ new_n3106;
  assign new_n3285 = new_n3284 ^ new_n3281;
  assign new_n3286 = n99 ^ n98;
  assign new_n3287 = ~new_n3124 & new_n3286;
  assign new_n3288 = ~new_n3287 & new_n155;
  assign new_n3289 = new_n3288 ^ n2;
  assign new_n3290 = new_n3289 ^ n100;
  assign new_n3291 = ~n98 & n3;
  assign new_n3292 = n99 ^ n3;
  assign new_n3293 = new_n3292 ^ new_n3291;
  assign new_n3294 = n2 & new_n3293;
  assign new_n3295 = new_n3294 ^ new_n3291;
  assign new_n3296 = new_n3295 ^ new_n3290;
  assign new_n3297 = ~n1 & new_n3296;
  assign new_n3298 = new_n3297 ^ new_n3290;
  assign new_n3299 = new_n3298 ^ new_n3285;
  assign new_n3300 = new_n3134 ^ new_n3107;
  assign new_n3301 = ~new_n3131 & new_n3300;
  assign new_n3302 = new_n3301 ^ new_n3134;
  assign new_n3303 = new_n3302 ^ new_n3299;
  assign new_n3304 = new_n3151 & new_n3153;
  assign new_n3305 = ~new_n259 & new_n3138;
  assign new_n3306 = ~new_n3143 & n67;
  assign new_n3307 = new_n3306 ^ new_n3305;
  assign new_n3308 = n68 & new_n3137;
  assign new_n3309 = n66 & new_n3149;
  assign new_n3310 = new_n3309 ^ new_n3308;
  assign new_n3311 = new_n3310 ^ new_n3307;
  assign new_n3312 = new_n3311 ^ n36;
  assign new_n3313 = n37 ^ n36;
  assign new_n3314 = n65 & new_n3313;
  assign new_n3315 = new_n3314 ^ new_n3312;
  assign new_n3316 = new_n3315 ^ new_n3304;
  assign new_n3317 = ~new_n2672 & n70;
  assign new_n3318 = ~new_n402 & new_n2667;
  assign new_n3319 = new_n3318 ^ new_n3317;
  assign new_n3320 = n71 & new_n2666;
  assign new_n3321 = n69 & new_n2664;
  assign new_n3322 = new_n3321 ^ new_n3320;
  assign new_n3323 = new_n3322 ^ new_n3319;
  assign new_n3324 = new_n3323 ^ n33;
  assign new_n3325 = new_n3324 ^ new_n3316;
  assign new_n3326 = new_n3166 ^ new_n3154;
  assign new_n3327 = ~new_n3163 & new_n3326;
  assign new_n3328 = new_n3327 ^ new_n3166;
  assign new_n3329 = new_n3328 ^ new_n3325;
  assign new_n3330 = n73 & new_n2246;
  assign new_n3331 = new_n595 & new_n2241;
  assign new_n3332 = new_n3331 ^ new_n3330;
  assign new_n3333 = n74 & new_n2240;
  assign new_n3334 = n72 & new_n2391;
  assign new_n3335 = new_n3334 ^ new_n3333;
  assign new_n3336 = new_n3335 ^ new_n3332;
  assign new_n3337 = new_n3336 ^ n30;
  assign new_n3338 = new_n3337 ^ new_n3329;
  assign new_n3339 = new_n3179 ^ new_n3167;
  assign new_n3340 = ~new_n3176 & new_n3339;
  assign new_n3341 = new_n3340 ^ new_n3179;
  assign new_n3342 = new_n3341 ^ new_n3338;
  assign new_n3343 = n76 & new_n1874;
  assign new_n3344 = ~new_n812 & new_n1864;
  assign new_n3345 = new_n3344 ^ new_n3343;
  assign new_n3346 = n77 & new_n1863;
  assign new_n3347 = n75 & new_n1868;
  assign new_n3348 = new_n3347 ^ new_n3346;
  assign new_n3349 = new_n3348 ^ new_n3345;
  assign new_n3350 = new_n3349 ^ n27;
  assign new_n3351 = new_n3350 ^ new_n3342;
  assign new_n3352 = new_n3192 ^ new_n3180;
  assign new_n3353 = ~new_n3189 & new_n3352;
  assign new_n3354 = new_n3353 ^ new_n3192;
  assign new_n3355 = new_n3354 ^ new_n3351;
  assign new_n3356 = ~new_n1506 & n79;
  assign new_n3357 = new_n1069 & new_n1501;
  assign new_n3358 = new_n3357 ^ new_n3356;
  assign new_n3359 = n80 & new_n1500;
  assign new_n3360 = n78 & new_n1512;
  assign new_n3361 = new_n3360 ^ new_n3359;
  assign new_n3362 = new_n3361 ^ new_n3358;
  assign new_n3363 = new_n3362 ^ n24;
  assign new_n3364 = new_n3363 ^ new_n3355;
  assign new_n3365 = new_n3205 ^ new_n3193;
  assign new_n3366 = ~new_n3202 & new_n3365;
  assign new_n3367 = new_n3366 ^ new_n3205;
  assign new_n3368 = new_n3367 ^ new_n3364;
  assign new_n3369 = ~new_n1198 & n82;
  assign new_n3370 = new_n1193 & new_n1363;
  assign new_n3371 = new_n3370 ^ new_n3369;
  assign new_n3372 = n83 & new_n1192;
  assign new_n3373 = n81 & new_n1204;
  assign new_n3374 = new_n3373 ^ new_n3372;
  assign new_n3375 = new_n3374 ^ new_n3371;
  assign new_n3376 = new_n3375 ^ n21;
  assign new_n3377 = new_n3376 ^ new_n3368;
  assign new_n3378 = new_n3218 ^ new_n3206;
  assign new_n3379 = ~new_n3215 & new_n3378;
  assign new_n3380 = new_n3379 ^ new_n3218;
  assign new_n3381 = new_n3380 ^ new_n3377;
  assign new_n3382 = ~new_n930 & n85;
  assign new_n3383 = new_n925 & new_n1694;
  assign new_n3384 = new_n3383 ^ new_n3382;
  assign new_n3385 = n86 & new_n924;
  assign new_n3386 = n84 & new_n936;
  assign new_n3387 = new_n3386 ^ new_n3385;
  assign new_n3388 = new_n3387 ^ new_n3384;
  assign new_n3389 = new_n3388 ^ n18;
  assign new_n3390 = new_n3389 ^ new_n3381;
  assign new_n3391 = new_n3231 ^ new_n3219;
  assign new_n3392 = ~new_n3228 & new_n3391;
  assign new_n3393 = new_n3392 ^ new_n3231;
  assign new_n3394 = new_n3393 ^ new_n3390;
  assign new_n3395 = n88 & new_n707;
  assign new_n3396 = new_n701 & new_n2063;
  assign new_n3397 = new_n3396 ^ new_n3395;
  assign new_n3398 = n89 & new_n700;
  assign new_n3399 = n87 & new_n787;
  assign new_n3400 = new_n3399 ^ new_n3398;
  assign new_n3401 = new_n3400 ^ new_n3397;
  assign new_n3402 = new_n3401 ^ n15;
  assign new_n3403 = new_n3402 ^ new_n3394;
  assign new_n3404 = new_n3244 ^ new_n3232;
  assign new_n3405 = ~new_n3241 & new_n3404;
  assign new_n3406 = new_n3405 ^ new_n3244;
  assign new_n3407 = new_n3406 ^ new_n3403;
  assign new_n3408 = n91 & new_n499;
  assign new_n3409 = ~new_n506 & new_n2481;
  assign new_n3410 = new_n3409 ^ new_n3408;
  assign new_n3411 = ~new_n505 & n92;
  assign new_n3412 = n90 & new_n579;
  assign new_n3413 = new_n3412 ^ new_n3411;
  assign new_n3414 = new_n3413 ^ new_n3410;
  assign new_n3415 = new_n3414 ^ n12;
  assign new_n3416 = new_n3415 ^ new_n3407;
  assign new_n3417 = new_n3257 ^ new_n3245;
  assign new_n3418 = ~new_n3254 & new_n3417;
  assign new_n3419 = new_n3418 ^ new_n3257;
  assign new_n3420 = new_n3419 ^ new_n3416;
  assign new_n3421 = n94 & new_n354;
  assign new_n3422 = new_n349 & new_n2934;
  assign new_n3423 = new_n3422 ^ new_n3421;
  assign new_n3424 = n95 & new_n348;
  assign new_n3425 = n93 & new_n391;
  assign new_n3426 = new_n3425 ^ new_n3424;
  assign new_n3427 = new_n3426 ^ new_n3423;
  assign new_n3428 = new_n3427 ^ n9;
  assign new_n3429 = new_n3428 ^ new_n3420;
  assign new_n3430 = new_n3270 ^ new_n3258;
  assign new_n3431 = ~new_n3267 & new_n3430;
  assign new_n3432 = new_n3431 ^ new_n3270;
  assign new_n3433 = new_n3432 ^ new_n3429;
  assign new_n3434 = n97 & new_n218;
  assign new_n3435 = new_n2952 ^ n98;
  assign new_n3436 = new_n208 & new_n3435;
  assign new_n3437 = new_n3436 ^ new_n3434;
  assign new_n3438 = n98 & new_n207;
  assign new_n3439 = n96 & new_n212;
  assign new_n3440 = new_n3439 ^ new_n3438;
  assign new_n3441 = new_n3440 ^ new_n3437;
  assign new_n3442 = new_n3441 ^ n6;
  assign new_n3443 = new_n3442 ^ new_n3433;
  assign new_n3444 = new_n3284 ^ new_n3271;
  assign new_n3445 = ~new_n3281 & new_n3444;
  assign new_n3446 = new_n3445 ^ new_n3284;
  assign new_n3447 = new_n3446 ^ new_n3443;
  assign new_n3448 = n99 & new_n180;
  assign new_n3449 = n2 & n100;
  assign new_n3450 = new_n3449 ^ new_n3448;
  assign new_n3451 = new_n3450 ^ n3;
  assign new_n3452 = n100 ^ n99;
  assign new_n3453 = ~new_n3287 & new_n3452;
  assign new_n3454 = ~new_n3453 & new_n155;
  assign new_n3455 = new_n3454 ^ n2;
  assign new_n3456 = new_n3455 ^ n101;
  assign new_n3457 = new_n3456 ^ new_n3451;
  assign new_n3458 = ~n1 & new_n3457;
  assign new_n3459 = new_n3458 ^ new_n3456;
  assign new_n3460 = new_n3459 ^ new_n3447;
  assign new_n3461 = new_n3302 ^ new_n3285;
  assign new_n3462 = ~new_n3299 & new_n3461;
  assign new_n3463 = new_n3462 ^ new_n3302;
  assign new_n3464 = new_n3463 ^ new_n3460;
  assign new_n3465 = ~new_n3304 & ~new_n3314;
  assign new_n3466 = ~new_n3465 & new_n3312;
  assign new_n3467 = n66 ^ n37;
  assign new_n3468 = ~new_n3467 & new_n3313;
  assign new_n3469 = new_n3468 ^ n36;
  assign new_n3470 = new_n3469 ^ n38;
  assign new_n3471 = ~n36 & ~n37;
  assign new_n3472 = new_n3471 ^ new_n3313;
  assign new_n3473 = new_n3472 ^ n38;
  assign new_n3474 = ~n65 & ~new_n3473;
  assign new_n3475 = new_n3474 ^ new_n3470;
  assign new_n3476 = new_n3475 ^ new_n3466;
  assign new_n3477 = ~new_n3143 & n68;
  assign new_n3478 = ~new_n304 & new_n3138;
  assign new_n3479 = new_n3478 ^ new_n3477;
  assign new_n3480 = n69 & new_n3137;
  assign new_n3481 = n67 & new_n3149;
  assign new_n3482 = new_n3481 ^ new_n3480;
  assign new_n3483 = new_n3482 ^ new_n3479;
  assign new_n3484 = new_n3483 ^ n36;
  assign new_n3485 = new_n3484 ^ new_n3476;
  assign new_n3486 = ~new_n2672 & n71;
  assign new_n3487 = ~new_n459 & new_n2667;
  assign new_n3488 = new_n3487 ^ new_n3486;
  assign new_n3489 = n72 & new_n2666;
  assign new_n3490 = n70 & new_n2664;
  assign new_n3491 = new_n3490 ^ new_n3489;
  assign new_n3492 = new_n3491 ^ new_n3488;
  assign new_n3493 = new_n3492 ^ n33;
  assign new_n3494 = new_n3493 ^ new_n3485;
  assign new_n3495 = new_n3328 ^ new_n3316;
  assign new_n3496 = ~new_n3325 & new_n3495;
  assign new_n3497 = new_n3496 ^ new_n3328;
  assign new_n3498 = new_n3497 ^ new_n3494;
  assign new_n3499 = n74 & new_n2246;
  assign new_n3500 = new_n660 & new_n2241;
  assign new_n3501 = new_n3500 ^ new_n3499;
  assign new_n3502 = n75 & new_n2240;
  assign new_n3503 = n73 & new_n2391;
  assign new_n3504 = new_n3503 ^ new_n3502;
  assign new_n3505 = new_n3504 ^ new_n3501;
  assign new_n3506 = new_n3505 ^ n30;
  assign new_n3507 = new_n3506 ^ new_n3498;
  assign new_n3508 = new_n3341 ^ new_n3337;
  assign new_n3509 = ~new_n3508 & new_n3338;
  assign new_n3510 = new_n3509 ^ new_n3329;
  assign new_n3511 = new_n3510 ^ new_n3507;
  assign new_n3512 = n77 & new_n1874;
  assign new_n3513 = ~new_n891 & new_n1864;
  assign new_n3514 = new_n3513 ^ new_n3512;
  assign new_n3515 = n78 & new_n1863;
  assign new_n3516 = n76 & new_n1868;
  assign new_n3517 = new_n3516 ^ new_n3515;
  assign new_n3518 = new_n3517 ^ new_n3514;
  assign new_n3519 = new_n3518 ^ n27;
  assign new_n3520 = new_n3519 ^ new_n3511;
  assign new_n3521 = new_n3354 ^ new_n3342;
  assign new_n3522 = ~new_n3351 & new_n3521;
  assign new_n3523 = new_n3522 ^ new_n3354;
  assign new_n3524 = new_n3523 ^ new_n3520;
  assign new_n3525 = ~new_n1506 & n80;
  assign new_n3526 = new_n1161 & new_n1501;
  assign new_n3527 = new_n3526 ^ new_n3525;
  assign new_n3528 = n81 & new_n1500;
  assign new_n3529 = n79 & new_n1512;
  assign new_n3530 = new_n3529 ^ new_n3528;
  assign new_n3531 = new_n3530 ^ new_n3527;
  assign new_n3532 = new_n3531 ^ n24;
  assign new_n3533 = new_n3532 ^ new_n3524;
  assign new_n3534 = new_n3367 ^ new_n3355;
  assign new_n3535 = ~new_n3364 & new_n3534;
  assign new_n3536 = new_n3535 ^ new_n3367;
  assign new_n3537 = new_n3536 ^ new_n3533;
  assign new_n3538 = ~new_n1198 & n83;
  assign new_n3539 = new_n1193 & new_n1468;
  assign new_n3540 = new_n3539 ^ new_n3538;
  assign new_n3541 = n84 & new_n1192;
  assign new_n3542 = n82 & new_n1204;
  assign new_n3543 = new_n3542 ^ new_n3541;
  assign new_n3544 = new_n3543 ^ new_n3540;
  assign new_n3545 = new_n3544 ^ n21;
  assign new_n3546 = new_n3545 ^ new_n3537;
  assign new_n3547 = new_n3380 ^ new_n3368;
  assign new_n3548 = ~new_n3377 & new_n3547;
  assign new_n3549 = new_n3548 ^ new_n3380;
  assign new_n3550 = new_n3549 ^ new_n3546;
  assign new_n3551 = ~new_n930 & n86;
  assign new_n3552 = new_n925 & new_n1811;
  assign new_n3553 = new_n3552 ^ new_n3551;
  assign new_n3554 = n87 & new_n924;
  assign new_n3555 = n85 & new_n936;
  assign new_n3556 = new_n3555 ^ new_n3554;
  assign new_n3557 = new_n3556 ^ new_n3553;
  assign new_n3558 = new_n3557 ^ n18;
  assign new_n3559 = new_n3558 ^ new_n3550;
  assign new_n3560 = new_n3393 ^ new_n3381;
  assign new_n3561 = ~new_n3390 & new_n3560;
  assign new_n3562 = new_n3561 ^ new_n3393;
  assign new_n3563 = new_n3562 ^ new_n3559;
  assign new_n3564 = n89 & new_n707;
  assign new_n3565 = new_n701 & new_n2193;
  assign new_n3566 = new_n3565 ^ new_n3564;
  assign new_n3567 = n90 & new_n700;
  assign new_n3568 = n88 & new_n787;
  assign new_n3569 = new_n3568 ^ new_n3567;
  assign new_n3570 = new_n3569 ^ new_n3566;
  assign new_n3571 = new_n3570 ^ n15;
  assign new_n3572 = new_n3571 ^ new_n3563;
  assign new_n3573 = new_n3406 ^ new_n3394;
  assign new_n3574 = ~new_n3403 & new_n3573;
  assign new_n3575 = new_n3574 ^ new_n3406;
  assign new_n3576 = new_n3575 ^ new_n3572;
  assign new_n3577 = n92 & new_n499;
  assign new_n3578 = ~new_n506 & new_n2628;
  assign new_n3579 = new_n3578 ^ new_n3577;
  assign new_n3580 = ~new_n505 & n93;
  assign new_n3581 = n91 & new_n579;
  assign new_n3582 = new_n3581 ^ new_n3580;
  assign new_n3583 = new_n3582 ^ new_n3579;
  assign new_n3584 = new_n3583 ^ n12;
  assign new_n3585 = new_n3584 ^ new_n3576;
  assign new_n3586 = new_n3419 ^ new_n3407;
  assign new_n3587 = ~new_n3416 & new_n3586;
  assign new_n3588 = new_n3587 ^ new_n3419;
  assign new_n3589 = new_n3588 ^ new_n3585;
  assign new_n3590 = n95 & new_n354;
  assign new_n3591 = new_n349 & new_n3095;
  assign new_n3592 = new_n3591 ^ new_n3590;
  assign new_n3593 = n96 & new_n348;
  assign new_n3594 = n94 & new_n391;
  assign new_n3595 = new_n3594 ^ new_n3593;
  assign new_n3596 = new_n3595 ^ new_n3592;
  assign new_n3597 = new_n3596 ^ n9;
  assign new_n3598 = new_n3597 ^ new_n3589;
  assign new_n3599 = new_n3432 ^ new_n3420;
  assign new_n3600 = ~new_n3429 & new_n3599;
  assign new_n3601 = new_n3600 ^ new_n3432;
  assign new_n3602 = new_n3601 ^ new_n3598;
  assign new_n3603 = n98 & new_n218;
  assign new_n3604 = new_n3286 ^ new_n3123;
  assign new_n3605 = new_n208 & new_n3604;
  assign new_n3606 = new_n3605 ^ new_n3603;
  assign new_n3607 = n99 & new_n207;
  assign new_n3608 = n97 & new_n212;
  assign new_n3609 = new_n3608 ^ new_n3607;
  assign new_n3610 = new_n3609 ^ new_n3606;
  assign new_n3611 = new_n3610 ^ n6;
  assign new_n3612 = new_n3611 ^ new_n3602;
  assign new_n3613 = new_n3446 ^ new_n3433;
  assign new_n3614 = ~new_n3443 & new_n3613;
  assign new_n3615 = new_n3614 ^ new_n3446;
  assign new_n3616 = new_n3615 ^ new_n3612;
  assign new_n3617 = n101 ^ n100;
  assign new_n3618 = new_n3453 & new_n3617;
  assign new_n3619 = new_n3618 ^ new_n3617;
  assign new_n3620 = ~new_n3619 & new_n155;
  assign new_n3621 = new_n3620 ^ n2;
  assign new_n3622 = new_n3621 ^ n102;
  assign new_n3623 = n101 ^ n3;
  assign new_n3624 = n100 ^ n3;
  assign new_n3625 = ~n100 & ~new_n3624;
  assign new_n3626 = new_n3625 ^ new_n3623;
  assign new_n3627 = new_n3626 ^ n100;
  assign new_n3628 = ~new_n3627 & new_n241;
  assign new_n3629 = new_n3628 ^ new_n3625;
  assign new_n3630 = new_n3629 ^ n100;
  assign new_n3631 = new_n3630 ^ new_n3622;
  assign new_n3632 = ~n1 & ~new_n3631;
  assign new_n3633 = new_n3632 ^ new_n3622;
  assign new_n3634 = new_n3633 ^ new_n3616;
  assign new_n3635 = new_n3463 ^ new_n3447;
  assign new_n3636 = ~new_n3460 & new_n3635;
  assign new_n3637 = new_n3636 ^ new_n3463;
  assign new_n3638 = new_n3637 ^ new_n3634;
  assign new_n3639 = ~new_n1506 & n81;
  assign new_n3640 = new_n1263 & new_n1501;
  assign new_n3641 = new_n3640 ^ new_n3639;
  assign new_n3642 = n82 & new_n1500;
  assign new_n3643 = n80 & new_n1512;
  assign new_n3644 = new_n3643 ^ new_n3642;
  assign new_n3645 = new_n3644 ^ new_n3641;
  assign new_n3646 = new_n3645 ^ n24;
  assign new_n3647 = new_n3536 ^ new_n3524;
  assign new_n3648 = ~new_n3533 & new_n3647;
  assign new_n3649 = new_n3648 ^ new_n3536;
  assign new_n3650 = new_n3649 ^ new_n3646;
  assign new_n3651 = n78 & new_n1874;
  assign new_n3652 = ~new_n982 & new_n1864;
  assign new_n3653 = new_n3652 ^ new_n3651;
  assign new_n3654 = n79 & new_n1863;
  assign new_n3655 = n77 & new_n1868;
  assign new_n3656 = new_n3655 ^ new_n3654;
  assign new_n3657 = new_n3656 ^ new_n3653;
  assign new_n3658 = new_n3657 ^ n27;
  assign new_n3659 = new_n3523 ^ new_n3511;
  assign new_n3660 = ~new_n3520 & new_n3659;
  assign new_n3661 = new_n3660 ^ new_n3523;
  assign new_n3662 = new_n3661 ^ new_n3658;
  assign new_n3663 = n75 & new_n2246;
  assign new_n3664 = ~new_n737 & new_n2241;
  assign new_n3665 = new_n3664 ^ new_n3663;
  assign new_n3666 = n76 & new_n2240;
  assign new_n3667 = n74 & new_n2391;
  assign new_n3668 = new_n3667 ^ new_n3666;
  assign new_n3669 = new_n3668 ^ new_n3665;
  assign new_n3670 = new_n3669 ^ n30;
  assign new_n3671 = new_n3510 ^ new_n3498;
  assign new_n3672 = ~new_n3507 & new_n3671;
  assign new_n3673 = new_n3672 ^ new_n3510;
  assign new_n3674 = new_n3673 ^ new_n3670;
  assign new_n3675 = n39 ^ n38;
  assign new_n3676 = ~new_n3675 & new_n3313;
  assign new_n3677 = new_n3676 ^ new_n3313;
  assign new_n3678 = ~new_n151 & new_n3677;
  assign new_n3679 = n67 & new_n3313;
  assign new_n3680 = new_n3679 ^ new_n3678;
  assign new_n3681 = ~new_n3313 & n38;
  assign new_n3682 = new_n3681 ^ new_n3472;
  assign new_n3683 = ~new_n3682 & n66;
  assign new_n3684 = new_n3683 ^ new_n3680;
  assign new_n3685 = new_n3684 ^ n39;
  assign new_n3686 = ~new_n3313 & n39;
  assign new_n3687 = new_n3686 ^ new_n3472;
  assign new_n3688 = ~new_n3687 & new_n3675;
  assign new_n3689 = n65 & new_n3688;
  assign new_n3690 = new_n3689 ^ new_n3685;
  assign new_n3691 = ~new_n3314 & ~new_n3475;
  assign new_n3692 = n39 & new_n3691;
  assign new_n3693 = new_n3692 ^ new_n3690;
  assign new_n3694 = ~new_n3143 & n69;
  assign new_n3695 = ~new_n339 & new_n3138;
  assign new_n3696 = new_n3695 ^ new_n3694;
  assign new_n3697 = n70 & new_n3137;
  assign new_n3698 = n68 & new_n3149;
  assign new_n3699 = new_n3698 ^ new_n3697;
  assign new_n3700 = new_n3699 ^ new_n3696;
  assign new_n3701 = new_n3700 ^ n36;
  assign new_n3702 = new_n3701 ^ new_n3693;
  assign new_n3703 = new_n3484 ^ new_n3475;
  assign new_n3704 = ~new_n3703 & new_n3476;
  assign new_n3705 = new_n3704 ^ new_n3466;
  assign new_n3706 = new_n3705 ^ new_n3702;
  assign new_n3707 = ~new_n2672 & n72;
  assign new_n3708 = new_n534 & new_n2667;
  assign new_n3709 = new_n3708 ^ new_n3707;
  assign new_n3710 = n73 & new_n2666;
  assign new_n3711 = n71 & new_n2664;
  assign new_n3712 = new_n3711 ^ new_n3710;
  assign new_n3713 = new_n3712 ^ new_n3709;
  assign new_n3714 = new_n3713 ^ n33;
  assign new_n3715 = new_n3714 ^ new_n3706;
  assign new_n3716 = new_n3497 ^ new_n3485;
  assign new_n3717 = ~new_n3494 & new_n3716;
  assign new_n3718 = new_n3717 ^ new_n3497;
  assign new_n3719 = new_n3718 ^ new_n3715;
  assign new_n3720 = new_n3719 ^ new_n3674;
  assign new_n3721 = new_n3720 ^ new_n3662;
  assign new_n3722 = new_n3721 ^ new_n3650;
  assign new_n3723 = ~new_n1198 & n84;
  assign new_n3724 = new_n1193 & new_n1584;
  assign new_n3725 = new_n3724 ^ new_n3723;
  assign new_n3726 = n85 & new_n1192;
  assign new_n3727 = n83 & new_n1204;
  assign new_n3728 = new_n3727 ^ new_n3726;
  assign new_n3729 = new_n3728 ^ new_n3725;
  assign new_n3730 = new_n3729 ^ n21;
  assign new_n3731 = new_n3730 ^ new_n3722;
  assign new_n3732 = new_n3549 ^ new_n3537;
  assign new_n3733 = ~new_n3546 & new_n3732;
  assign new_n3734 = new_n3733 ^ new_n3549;
  assign new_n3735 = new_n3734 ^ new_n3731;
  assign new_n3736 = ~new_n930 & n87;
  assign new_n3737 = new_n925 & new_n1940;
  assign new_n3738 = new_n3737 ^ new_n3736;
  assign new_n3739 = n88 & new_n924;
  assign new_n3740 = n86 & new_n936;
  assign new_n3741 = new_n3740 ^ new_n3739;
  assign new_n3742 = new_n3741 ^ new_n3738;
  assign new_n3743 = new_n3742 ^ n18;
  assign new_n3744 = new_n3743 ^ new_n3735;
  assign new_n3745 = new_n3562 ^ new_n3550;
  assign new_n3746 = ~new_n3559 & new_n3745;
  assign new_n3747 = new_n3746 ^ new_n3562;
  assign new_n3748 = new_n3747 ^ new_n3744;
  assign new_n3749 = n90 & new_n707;
  assign new_n3750 = new_n701 & new_n2341;
  assign new_n3751 = new_n3750 ^ new_n3749;
  assign new_n3752 = n91 & new_n700;
  assign new_n3753 = n89 & new_n787;
  assign new_n3754 = new_n3753 ^ new_n3752;
  assign new_n3755 = new_n3754 ^ new_n3751;
  assign new_n3756 = new_n3755 ^ n15;
  assign new_n3757 = new_n3756 ^ new_n3748;
  assign new_n3758 = new_n3575 ^ new_n3563;
  assign new_n3759 = ~new_n3572 & new_n3758;
  assign new_n3760 = new_n3759 ^ new_n3575;
  assign new_n3761 = new_n3760 ^ new_n3757;
  assign new_n3762 = n93 & new_n499;
  assign new_n3763 = ~new_n506 & new_n2785;
  assign new_n3764 = new_n3763 ^ new_n3762;
  assign new_n3765 = ~new_n505 & n94;
  assign new_n3766 = n92 & new_n579;
  assign new_n3767 = new_n3766 ^ new_n3765;
  assign new_n3768 = new_n3767 ^ new_n3764;
  assign new_n3769 = new_n3768 ^ n12;
  assign new_n3770 = new_n3769 ^ new_n3761;
  assign new_n3771 = new_n3588 ^ new_n3576;
  assign new_n3772 = ~new_n3585 & new_n3771;
  assign new_n3773 = new_n3772 ^ new_n3588;
  assign new_n3774 = new_n3773 ^ new_n3770;
  assign new_n3775 = n96 & new_n354;
  assign new_n3776 = new_n349 & new_n3273;
  assign new_n3777 = new_n3776 ^ new_n3775;
  assign new_n3778 = n97 & new_n348;
  assign new_n3779 = n95 & new_n391;
  assign new_n3780 = new_n3779 ^ new_n3778;
  assign new_n3781 = new_n3780 ^ new_n3777;
  assign new_n3782 = new_n3781 ^ n9;
  assign new_n3783 = new_n3782 ^ new_n3774;
  assign new_n3784 = new_n3601 ^ new_n3589;
  assign new_n3785 = ~new_n3598 & new_n3784;
  assign new_n3786 = new_n3785 ^ new_n3601;
  assign new_n3787 = new_n3786 ^ new_n3783;
  assign new_n3788 = n99 & new_n218;
  assign new_n3789 = new_n3287 ^ n100;
  assign new_n3790 = new_n208 & new_n3789;
  assign new_n3791 = new_n3790 ^ new_n3788;
  assign new_n3792 = n100 & new_n207;
  assign new_n3793 = n98 & new_n212;
  assign new_n3794 = new_n3793 ^ new_n3792;
  assign new_n3795 = new_n3794 ^ new_n3791;
  assign new_n3796 = new_n3795 ^ n6;
  assign new_n3797 = new_n3796 ^ new_n3787;
  assign new_n3798 = new_n3615 ^ new_n3602;
  assign new_n3799 = ~new_n3612 & new_n3798;
  assign new_n3800 = new_n3799 ^ new_n3615;
  assign new_n3801 = new_n3800 ^ new_n3797;
  assign new_n3802 = ~new_n3287 & n99;
  assign new_n3803 = new_n3802 ^ new_n3287;
  assign new_n3804 = ~n100 & ~n102;
  assign new_n3805 = n102 ^ n100;
  assign new_n3806 = new_n3805 ^ new_n3804;
  assign new_n3807 = ~new_n3806 & new_n3803;
  assign new_n3808 = ~n101 & ~new_n3807;
  assign new_n3809 = ~new_n3802 & new_n3804;
  assign new_n3810 = ~new_n3808 & ~new_n3809;
  assign new_n3811 = new_n3810 ^ n102;
  assign new_n3812 = ~new_n3811 & new_n155;
  assign new_n3813 = new_n3812 ^ n2;
  assign new_n3814 = new_n3813 ^ n103;
  assign new_n3815 = n3 & n101;
  assign new_n3816 = new_n3815 ^ n102;
  assign new_n3817 = ~n2 & new_n3816;
  assign new_n3818 = new_n3817 ^ n102;
  assign new_n3819 = new_n3818 ^ n3;
  assign new_n3820 = new_n3819 ^ new_n3814;
  assign new_n3821 = ~n1 & new_n3820;
  assign new_n3822 = new_n3821 ^ new_n3814;
  assign new_n3823 = new_n3822 ^ new_n3801;
  assign new_n3824 = new_n3637 ^ new_n3616;
  assign new_n3825 = ~new_n3634 & new_n3824;
  assign new_n3826 = new_n3825 ^ new_n3637;
  assign new_n3827 = new_n3826 ^ new_n3823;
  assign new_n3828 = new_n3690 & new_n3692;
  assign new_n3829 = ~new_n259 & new_n3677;
  assign new_n3830 = ~new_n3682 & n67;
  assign new_n3831 = new_n3830 ^ new_n3829;
  assign new_n3832 = n68 & new_n3676;
  assign new_n3833 = n66 & new_n3688;
  assign new_n3834 = new_n3833 ^ new_n3832;
  assign new_n3835 = new_n3834 ^ new_n3831;
  assign new_n3836 = new_n3835 ^ n39;
  assign new_n3837 = n40 ^ n39;
  assign new_n3838 = n65 & new_n3837;
  assign new_n3839 = new_n3838 ^ new_n3836;
  assign new_n3840 = new_n3839 ^ new_n3828;
  assign new_n3841 = ~new_n3143 & n70;
  assign new_n3842 = ~new_n402 & new_n3138;
  assign new_n3843 = new_n3842 ^ new_n3841;
  assign new_n3844 = n71 & new_n3137;
  assign new_n3845 = n69 & new_n3149;
  assign new_n3846 = new_n3845 ^ new_n3844;
  assign new_n3847 = new_n3846 ^ new_n3843;
  assign new_n3848 = new_n3847 ^ n36;
  assign new_n3849 = new_n3848 ^ new_n3840;
  assign new_n3850 = new_n3705 ^ new_n3693;
  assign new_n3851 = ~new_n3702 & new_n3850;
  assign new_n3852 = new_n3851 ^ new_n3705;
  assign new_n3853 = new_n3852 ^ new_n3849;
  assign new_n3854 = ~new_n2672 & n73;
  assign new_n3855 = new_n595 & new_n2667;
  assign new_n3856 = new_n3855 ^ new_n3854;
  assign new_n3857 = n72 & new_n2664;
  assign new_n3858 = n74 & new_n2666;
  assign new_n3859 = new_n3858 ^ new_n3857;
  assign new_n3860 = new_n3859 ^ new_n3856;
  assign new_n3861 = new_n3860 ^ n33;
  assign new_n3862 = new_n3861 ^ new_n3853;
  assign new_n3863 = new_n3718 ^ new_n3706;
  assign new_n3864 = ~new_n3715 & new_n3863;
  assign new_n3865 = new_n3864 ^ new_n3718;
  assign new_n3866 = new_n3865 ^ new_n3862;
  assign new_n3867 = n76 & new_n2246;
  assign new_n3868 = ~new_n812 & new_n2241;
  assign new_n3869 = new_n3868 ^ new_n3867;
  assign new_n3870 = n77 & new_n2240;
  assign new_n3871 = n75 & new_n2391;
  assign new_n3872 = new_n3871 ^ new_n3870;
  assign new_n3873 = new_n3872 ^ new_n3869;
  assign new_n3874 = new_n3873 ^ n30;
  assign new_n3875 = new_n3874 ^ new_n3866;
  assign new_n3876 = new_n3719 ^ new_n3670;
  assign new_n3877 = ~new_n3876 & new_n3674;
  assign new_n3878 = new_n3877 ^ new_n3673;
  assign new_n3879 = new_n3878 ^ new_n3875;
  assign new_n3880 = n79 & new_n1874;
  assign new_n3881 = new_n1069 & new_n1864;
  assign new_n3882 = new_n3881 ^ new_n3880;
  assign new_n3883 = n80 & new_n1863;
  assign new_n3884 = n78 & new_n1868;
  assign new_n3885 = new_n3884 ^ new_n3883;
  assign new_n3886 = new_n3885 ^ new_n3882;
  assign new_n3887 = new_n3886 ^ n27;
  assign new_n3888 = new_n3887 ^ new_n3879;
  assign new_n3889 = new_n3720 ^ new_n3658;
  assign new_n3890 = ~new_n3889 & new_n3662;
  assign new_n3891 = new_n3890 ^ new_n3661;
  assign new_n3892 = new_n3891 ^ new_n3888;
  assign new_n3893 = ~new_n1506 & n82;
  assign new_n3894 = new_n1363 & new_n1501;
  assign new_n3895 = new_n3894 ^ new_n3893;
  assign new_n3896 = n83 & new_n1500;
  assign new_n3897 = n81 & new_n1512;
  assign new_n3898 = new_n3897 ^ new_n3896;
  assign new_n3899 = new_n3898 ^ new_n3895;
  assign new_n3900 = new_n3899 ^ n24;
  assign new_n3901 = new_n3900 ^ new_n3892;
  assign new_n3902 = new_n3721 ^ new_n3646;
  assign new_n3903 = ~new_n3902 & new_n3650;
  assign new_n3904 = new_n3903 ^ new_n3649;
  assign new_n3905 = new_n3904 ^ new_n3901;
  assign new_n3906 = ~new_n1198 & n85;
  assign new_n3907 = new_n1193 & new_n1694;
  assign new_n3908 = new_n3907 ^ new_n3906;
  assign new_n3909 = n86 & new_n1192;
  assign new_n3910 = n84 & new_n1204;
  assign new_n3911 = new_n3910 ^ new_n3909;
  assign new_n3912 = new_n3911 ^ new_n3908;
  assign new_n3913 = new_n3912 ^ n21;
  assign new_n3914 = new_n3913 ^ new_n3905;
  assign new_n3915 = new_n3734 ^ new_n3722;
  assign new_n3916 = ~new_n3731 & new_n3915;
  assign new_n3917 = new_n3916 ^ new_n3734;
  assign new_n3918 = new_n3917 ^ new_n3914;
  assign new_n3919 = ~new_n930 & n88;
  assign new_n3920 = new_n925 & new_n2063;
  assign new_n3921 = new_n3920 ^ new_n3919;
  assign new_n3922 = n89 & new_n924;
  assign new_n3923 = n87 & new_n936;
  assign new_n3924 = new_n3923 ^ new_n3922;
  assign new_n3925 = new_n3924 ^ new_n3921;
  assign new_n3926 = new_n3925 ^ n18;
  assign new_n3927 = new_n3926 ^ new_n3918;
  assign new_n3928 = new_n3747 ^ new_n3735;
  assign new_n3929 = ~new_n3744 & new_n3928;
  assign new_n3930 = new_n3929 ^ new_n3747;
  assign new_n3931 = new_n3930 ^ new_n3927;
  assign new_n3932 = n91 & new_n707;
  assign new_n3933 = new_n701 & new_n2481;
  assign new_n3934 = new_n3933 ^ new_n3932;
  assign new_n3935 = n92 & new_n700;
  assign new_n3936 = n90 & new_n787;
  assign new_n3937 = new_n3936 ^ new_n3935;
  assign new_n3938 = new_n3937 ^ new_n3934;
  assign new_n3939 = new_n3938 ^ n15;
  assign new_n3940 = new_n3939 ^ new_n3931;
  assign new_n3941 = new_n3760 ^ new_n3748;
  assign new_n3942 = ~new_n3757 & new_n3941;
  assign new_n3943 = new_n3942 ^ new_n3760;
  assign new_n3944 = new_n3943 ^ new_n3940;
  assign new_n3945 = n94 & new_n499;
  assign new_n3946 = ~new_n506 & new_n2934;
  assign new_n3947 = new_n3946 ^ new_n3945;
  assign new_n3948 = ~new_n505 & n95;
  assign new_n3949 = n93 & new_n579;
  assign new_n3950 = new_n3949 ^ new_n3948;
  assign new_n3951 = new_n3950 ^ new_n3947;
  assign new_n3952 = new_n3951 ^ n12;
  assign new_n3953 = new_n3952 ^ new_n3944;
  assign new_n3954 = new_n3773 ^ new_n3761;
  assign new_n3955 = ~new_n3770 & new_n3954;
  assign new_n3956 = new_n3955 ^ new_n3773;
  assign new_n3957 = new_n3956 ^ new_n3953;
  assign new_n3958 = n97 & new_n354;
  assign new_n3959 = new_n349 & new_n3435;
  assign new_n3960 = new_n3959 ^ new_n3958;
  assign new_n3961 = n98 & new_n348;
  assign new_n3962 = n96 & new_n391;
  assign new_n3963 = new_n3962 ^ new_n3961;
  assign new_n3964 = new_n3963 ^ new_n3960;
  assign new_n3965 = new_n3964 ^ n9;
  assign new_n3966 = new_n3965 ^ new_n3957;
  assign new_n3967 = new_n3786 ^ new_n3774;
  assign new_n3968 = ~new_n3783 & new_n3967;
  assign new_n3969 = new_n3968 ^ new_n3786;
  assign new_n3970 = new_n3969 ^ new_n3966;
  assign new_n3971 = n100 & new_n218;
  assign new_n3972 = new_n3453 ^ n101;
  assign new_n3973 = new_n208 & new_n3972;
  assign new_n3974 = new_n3973 ^ new_n3971;
  assign new_n3975 = n101 & new_n207;
  assign new_n3976 = n99 & new_n212;
  assign new_n3977 = new_n3976 ^ new_n3975;
  assign new_n3978 = new_n3977 ^ new_n3974;
  assign new_n3979 = new_n3978 ^ n6;
  assign new_n3980 = new_n3979 ^ new_n3970;
  assign new_n3981 = new_n3800 ^ new_n3787;
  assign new_n3982 = ~new_n3797 & new_n3981;
  assign new_n3983 = new_n3982 ^ new_n3800;
  assign new_n3984 = new_n3983 ^ new_n3980;
  assign new_n3985 = n102 & new_n3810;
  assign new_n3986 = new_n3985 ^ new_n3811;
  assign new_n3987 = n103 & new_n3986;
  assign new_n3988 = ~n103 & ~new_n3985;
  assign new_n3989 = new_n3988 ^ new_n3987;
  assign new_n3990 = new_n155 & new_n3989;
  assign new_n3991 = new_n3990 ^ n2;
  assign new_n3992 = new_n3991 ^ n104;
  assign new_n3993 = n103 ^ n3;
  assign new_n3994 = ~n102 & n3;
  assign new_n3995 = new_n3994 ^ new_n3993;
  assign new_n3996 = ~n2 & new_n3995;
  assign new_n3997 = new_n3996 ^ new_n3993;
  assign new_n3998 = new_n3997 ^ new_n3992;
  assign new_n3999 = ~n1 & new_n3998;
  assign new_n4000 = new_n3999 ^ new_n3992;
  assign new_n4001 = new_n4000 ^ new_n3984;
  assign new_n4002 = new_n3826 ^ new_n3801;
  assign new_n4003 = ~new_n3823 & new_n4002;
  assign new_n4004 = new_n4003 ^ new_n3826;
  assign new_n4005 = new_n4004 ^ new_n4001;
  assign new_n4006 = ~new_n3143 & n71;
  assign new_n4007 = ~new_n459 & new_n3138;
  assign new_n4008 = new_n4007 ^ new_n4006;
  assign new_n4009 = n72 & new_n3137;
  assign new_n4010 = n70 & new_n3149;
  assign new_n4011 = new_n4010 ^ new_n4009;
  assign new_n4012 = new_n4011 ^ new_n4008;
  assign new_n4013 = new_n4012 ^ n36;
  assign new_n4014 = new_n3852 ^ new_n3840;
  assign new_n4015 = ~new_n3849 & new_n4014;
  assign new_n4016 = new_n4015 ^ new_n3852;
  assign new_n4017 = new_n4016 ^ new_n4013;
  assign new_n4018 = n66 ^ n40;
  assign new_n4019 = ~new_n4018 & new_n3837;
  assign new_n4020 = new_n4019 ^ n39;
  assign new_n4021 = new_n4020 ^ n41;
  assign new_n4022 = ~n39 & ~n40;
  assign new_n4023 = new_n4022 ^ n41;
  assign new_n4024 = ~n65 & ~new_n4023;
  assign new_n4025 = new_n4024 ^ new_n3837;
  assign new_n4026 = new_n4025 ^ new_n3838;
  assign new_n4027 = new_n4026 ^ new_n4021;
  assign new_n4028 = ~new_n3828 & ~new_n3838;
  assign new_n4029 = ~new_n4028 & new_n3836;
  assign new_n4030 = new_n4029 ^ new_n4027;
  assign new_n4031 = ~new_n3682 & n68;
  assign new_n4032 = ~new_n304 & new_n3677;
  assign new_n4033 = new_n4032 ^ new_n4031;
  assign new_n4034 = n69 & new_n3676;
  assign new_n4035 = n67 & new_n3688;
  assign new_n4036 = new_n4035 ^ new_n4034;
  assign new_n4037 = new_n4036 ^ new_n4033;
  assign new_n4038 = new_n4037 ^ n39;
  assign new_n4039 = new_n4038 ^ new_n4030;
  assign new_n4040 = new_n4039 ^ new_n4017;
  assign new_n4041 = ~new_n2672 & n74;
  assign new_n4042 = new_n660 & new_n2667;
  assign new_n4043 = new_n4042 ^ new_n4041;
  assign new_n4044 = n75 & new_n2666;
  assign new_n4045 = n73 & new_n2664;
  assign new_n4046 = new_n4045 ^ new_n4044;
  assign new_n4047 = new_n4046 ^ new_n4043;
  assign new_n4048 = new_n4047 ^ n33;
  assign new_n4049 = new_n4048 ^ new_n4040;
  assign new_n4050 = new_n3865 ^ new_n3853;
  assign new_n4051 = ~new_n3862 & new_n4050;
  assign new_n4052 = new_n4051 ^ new_n3865;
  assign new_n4053 = new_n4052 ^ new_n4049;
  assign new_n4054 = n77 & new_n2246;
  assign new_n4055 = ~new_n891 & new_n2241;
  assign new_n4056 = new_n4055 ^ new_n4054;
  assign new_n4057 = n78 & new_n2240;
  assign new_n4058 = n76 & new_n2391;
  assign new_n4059 = new_n4058 ^ new_n4057;
  assign new_n4060 = new_n4059 ^ new_n4056;
  assign new_n4061 = new_n4060 ^ n30;
  assign new_n4062 = new_n4061 ^ new_n4053;
  assign new_n4063 = new_n3878 ^ new_n3866;
  assign new_n4064 = ~new_n3875 & new_n4063;
  assign new_n4065 = new_n4064 ^ new_n3878;
  assign new_n4066 = new_n4065 ^ new_n4062;
  assign new_n4067 = n80 & new_n1874;
  assign new_n4068 = new_n1161 & new_n1864;
  assign new_n4069 = new_n4068 ^ new_n4067;
  assign new_n4070 = n79 & new_n1868;
  assign new_n4071 = n81 & new_n1863;
  assign new_n4072 = new_n4071 ^ new_n4070;
  assign new_n4073 = new_n4072 ^ new_n4069;
  assign new_n4074 = new_n4073 ^ n27;
  assign new_n4075 = new_n4074 ^ new_n4066;
  assign new_n4076 = new_n3891 ^ new_n3879;
  assign new_n4077 = ~new_n3888 & new_n4076;
  assign new_n4078 = new_n4077 ^ new_n3891;
  assign new_n4079 = new_n4078 ^ new_n4075;
  assign new_n4080 = ~new_n1506 & n83;
  assign new_n4081 = new_n1468 & new_n1501;
  assign new_n4082 = new_n4081 ^ new_n4080;
  assign new_n4083 = n84 & new_n1500;
  assign new_n4084 = n82 & new_n1512;
  assign new_n4085 = new_n4084 ^ new_n4083;
  assign new_n4086 = new_n4085 ^ new_n4082;
  assign new_n4087 = new_n4086 ^ n24;
  assign new_n4088 = new_n4087 ^ new_n4079;
  assign new_n4089 = new_n3904 ^ new_n3892;
  assign new_n4090 = ~new_n3901 & new_n4089;
  assign new_n4091 = new_n4090 ^ new_n3904;
  assign new_n4092 = new_n4091 ^ new_n4088;
  assign new_n4093 = ~new_n1198 & n86;
  assign new_n4094 = new_n1193 & new_n1811;
  assign new_n4095 = new_n4094 ^ new_n4093;
  assign new_n4096 = n87 & new_n1192;
  assign new_n4097 = n85 & new_n1204;
  assign new_n4098 = new_n4097 ^ new_n4096;
  assign new_n4099 = new_n4098 ^ new_n4095;
  assign new_n4100 = new_n4099 ^ n21;
  assign new_n4101 = new_n4100 ^ new_n4092;
  assign new_n4102 = new_n3917 ^ new_n3905;
  assign new_n4103 = ~new_n3914 & new_n4102;
  assign new_n4104 = new_n4103 ^ new_n3917;
  assign new_n4105 = new_n4104 ^ new_n4101;
  assign new_n4106 = ~new_n930 & n89;
  assign new_n4107 = new_n925 & new_n2193;
  assign new_n4108 = new_n4107 ^ new_n4106;
  assign new_n4109 = n90 & new_n924;
  assign new_n4110 = n88 & new_n936;
  assign new_n4111 = new_n4110 ^ new_n4109;
  assign new_n4112 = new_n4111 ^ new_n4108;
  assign new_n4113 = new_n4112 ^ n18;
  assign new_n4114 = new_n4113 ^ new_n4105;
  assign new_n4115 = new_n3930 ^ new_n3918;
  assign new_n4116 = ~new_n3927 & new_n4115;
  assign new_n4117 = new_n4116 ^ new_n3930;
  assign new_n4118 = new_n4117 ^ new_n4114;
  assign new_n4119 = n92 & new_n707;
  assign new_n4120 = new_n701 & new_n2628;
  assign new_n4121 = new_n4120 ^ new_n4119;
  assign new_n4122 = n93 & new_n700;
  assign new_n4123 = n91 & new_n787;
  assign new_n4124 = new_n4123 ^ new_n4122;
  assign new_n4125 = new_n4124 ^ new_n4121;
  assign new_n4126 = new_n4125 ^ n15;
  assign new_n4127 = new_n4126 ^ new_n4118;
  assign new_n4128 = new_n3943 ^ new_n3931;
  assign new_n4129 = ~new_n3940 & new_n4128;
  assign new_n4130 = new_n4129 ^ new_n3943;
  assign new_n4131 = new_n4130 ^ new_n4127;
  assign new_n4132 = n95 & new_n499;
  assign new_n4133 = ~new_n506 & new_n3095;
  assign new_n4134 = new_n4133 ^ new_n4132;
  assign new_n4135 = ~new_n505 & n96;
  assign new_n4136 = n94 & new_n579;
  assign new_n4137 = new_n4136 ^ new_n4135;
  assign new_n4138 = new_n4137 ^ new_n4134;
  assign new_n4139 = new_n4138 ^ n12;
  assign new_n4140 = new_n4139 ^ new_n4131;
  assign new_n4141 = new_n3956 ^ new_n3944;
  assign new_n4142 = ~new_n3953 & new_n4141;
  assign new_n4143 = new_n4142 ^ new_n3956;
  assign new_n4144 = new_n4143 ^ new_n4140;
  assign new_n4145 = n98 & new_n354;
  assign new_n4146 = new_n349 & new_n3604;
  assign new_n4147 = new_n4146 ^ new_n4145;
  assign new_n4148 = n99 & new_n348;
  assign new_n4149 = n97 & new_n391;
  assign new_n4150 = new_n4149 ^ new_n4148;
  assign new_n4151 = new_n4150 ^ new_n4147;
  assign new_n4152 = new_n4151 ^ n9;
  assign new_n4153 = new_n4152 ^ new_n4144;
  assign new_n4154 = new_n3969 ^ new_n3957;
  assign new_n4155 = ~new_n3966 & new_n4154;
  assign new_n4156 = new_n4155 ^ new_n3969;
  assign new_n4157 = new_n4156 ^ new_n4153;
  assign new_n4158 = n101 & new_n218;
  assign new_n4159 = new_n3619 ^ n102;
  assign new_n4160 = new_n208 & new_n4159;
  assign new_n4161 = new_n4160 ^ new_n4158;
  assign new_n4162 = n102 & new_n207;
  assign new_n4163 = n100 & new_n212;
  assign new_n4164 = new_n4163 ^ new_n4162;
  assign new_n4165 = new_n4164 ^ new_n4161;
  assign new_n4166 = new_n4165 ^ n6;
  assign new_n4167 = new_n4166 ^ new_n4157;
  assign new_n4168 = new_n3983 ^ new_n3970;
  assign new_n4169 = ~new_n3980 & new_n4168;
  assign new_n4170 = new_n4169 ^ new_n3983;
  assign new_n4171 = new_n4170 ^ new_n4167;
  assign new_n4172 = ~n104 & ~new_n3987;
  assign new_n4173 = ~new_n3988 & n104;
  assign new_n4174 = new_n4173 ^ new_n4172;
  assign new_n4175 = new_n155 & new_n4174;
  assign new_n4176 = new_n4175 ^ n2;
  assign new_n4177 = new_n4176 ^ n105;
  assign new_n4178 = n104 ^ n3;
  assign new_n4179 = ~n103 & n3;
  assign new_n4180 = new_n4179 ^ new_n4178;
  assign new_n4181 = ~n2 & new_n4180;
  assign new_n4182 = new_n4181 ^ new_n4178;
  assign new_n4183 = new_n4182 ^ new_n4177;
  assign new_n4184 = ~n1 & new_n4183;
  assign new_n4185 = new_n4184 ^ new_n4177;
  assign new_n4186 = new_n4185 ^ new_n4171;
  assign new_n4187 = new_n4004 ^ new_n3984;
  assign new_n4188 = ~new_n4001 & new_n4187;
  assign new_n4189 = new_n4188 ^ new_n4004;
  assign new_n4190 = new_n4189 ^ new_n4186;
  assign new_n4191 = ~new_n3682 & n69;
  assign new_n4192 = ~new_n339 & new_n3677;
  assign new_n4193 = new_n4192 ^ new_n4191;
  assign new_n4194 = n70 & new_n3676;
  assign new_n4195 = n68 & new_n3688;
  assign new_n4196 = new_n4195 ^ new_n4194;
  assign new_n4197 = new_n4196 ^ new_n4193;
  assign new_n4198 = new_n4197 ^ n39;
  assign new_n4199 = n42 ^ n41;
  assign new_n4200 = ~new_n4199 & new_n3837;
  assign new_n4201 = new_n4200 ^ new_n3837;
  assign new_n4202 = ~new_n151 & new_n4201;
  assign new_n4203 = ~new_n3837 & n42;
  assign new_n4204 = new_n4022 ^ new_n3837;
  assign new_n4205 = new_n4204 ^ new_n4203;
  assign new_n4206 = ~new_n4205 & new_n4199;
  assign new_n4207 = n65 & new_n4206;
  assign new_n4208 = new_n4207 ^ new_n4202;
  assign new_n4209 = n67 & new_n3837;
  assign new_n4210 = new_n4209 ^ new_n4208;
  assign new_n4211 = ~new_n3837 & n41;
  assign new_n4212 = new_n4211 ^ new_n4204;
  assign new_n4213 = ~new_n4212 & n66;
  assign new_n4214 = new_n4213 ^ new_n4210;
  assign new_n4215 = new_n4023 ^ new_n4022;
  assign new_n4216 = new_n4204 ^ new_n4022;
  assign new_n4217 = ~new_n4216 & new_n4215;
  assign new_n4218 = new_n4217 ^ new_n4022;
  assign new_n4219 = ~new_n4218 & n42;
  assign new_n4220 = ~new_n4022 & new_n3837;
  assign new_n4221 = n42 & new_n4220;
  assign new_n4222 = new_n4221 ^ new_n4219;
  assign new_n4223 = new_n4222 ^ new_n4221;
  assign new_n4224 = new_n4223 ^ new_n4222;
  assign new_n4225 = new_n4222 ^ n66;
  assign new_n4226 = new_n4225 ^ new_n4222;
  assign new_n4227 = ~new_n4226 & new_n4224;
  assign new_n4228 = new_n4227 ^ new_n4222;
  assign new_n4229 = ~n65 & new_n4228;
  assign new_n4230 = new_n4229 ^ new_n4219;
  assign new_n4231 = new_n4230 ^ new_n4214;
  assign new_n4232 = new_n4231 ^ new_n4198;
  assign new_n4233 = new_n4038 ^ new_n4027;
  assign new_n4234 = ~new_n4233 & new_n4030;
  assign new_n4235 = new_n4234 ^ new_n4029;
  assign new_n4236 = new_n4235 ^ new_n4232;
  assign new_n4237 = ~new_n3143 & n72;
  assign new_n4238 = new_n534 & new_n3138;
  assign new_n4239 = new_n4238 ^ new_n4237;
  assign new_n4240 = n71 & new_n3149;
  assign new_n4241 = n73 & new_n3137;
  assign new_n4242 = new_n4241 ^ new_n4240;
  assign new_n4243 = new_n4242 ^ new_n4239;
  assign new_n4244 = new_n4243 ^ n36;
  assign new_n4245 = new_n4244 ^ new_n4236;
  assign new_n4246 = new_n4039 ^ new_n4013;
  assign new_n4247 = ~new_n4246 & new_n4017;
  assign new_n4248 = new_n4247 ^ new_n4016;
  assign new_n4249 = new_n4248 ^ new_n4245;
  assign new_n4250 = ~new_n2672 & n75;
  assign new_n4251 = ~new_n737 & new_n2667;
  assign new_n4252 = new_n4251 ^ new_n4250;
  assign new_n4253 = n76 & new_n2666;
  assign new_n4254 = n74 & new_n2664;
  assign new_n4255 = new_n4254 ^ new_n4253;
  assign new_n4256 = new_n4255 ^ new_n4252;
  assign new_n4257 = new_n4256 ^ n33;
  assign new_n4258 = new_n4257 ^ new_n4249;
  assign new_n4259 = new_n4052 ^ new_n4040;
  assign new_n4260 = ~new_n4049 & new_n4259;
  assign new_n4261 = new_n4260 ^ new_n4052;
  assign new_n4262 = new_n4261 ^ new_n4258;
  assign new_n4263 = n78 & new_n2246;
  assign new_n4264 = ~new_n982 & new_n2241;
  assign new_n4265 = new_n4264 ^ new_n4263;
  assign new_n4266 = n79 & new_n2240;
  assign new_n4267 = n77 & new_n2391;
  assign new_n4268 = new_n4267 ^ new_n4266;
  assign new_n4269 = new_n4268 ^ new_n4265;
  assign new_n4270 = new_n4269 ^ n30;
  assign new_n4271 = new_n4270 ^ new_n4262;
  assign new_n4272 = new_n4065 ^ new_n4053;
  assign new_n4273 = ~new_n4062 & new_n4272;
  assign new_n4274 = new_n4273 ^ new_n4065;
  assign new_n4275 = new_n4274 ^ new_n4271;
  assign new_n4276 = n81 & new_n1874;
  assign new_n4277 = new_n1263 & new_n1864;
  assign new_n4278 = new_n4277 ^ new_n4276;
  assign new_n4279 = n82 & new_n1863;
  assign new_n4280 = n80 & new_n1868;
  assign new_n4281 = new_n4280 ^ new_n4279;
  assign new_n4282 = new_n4281 ^ new_n4278;
  assign new_n4283 = new_n4282 ^ n27;
  assign new_n4284 = new_n4283 ^ new_n4275;
  assign new_n4285 = new_n4078 ^ new_n4066;
  assign new_n4286 = ~new_n4075 & new_n4285;
  assign new_n4287 = new_n4286 ^ new_n4078;
  assign new_n4288 = new_n4287 ^ new_n4284;
  assign new_n4289 = ~new_n1506 & n84;
  assign new_n4290 = new_n1501 & new_n1584;
  assign new_n4291 = new_n4290 ^ new_n4289;
  assign new_n4292 = n85 & new_n1500;
  assign new_n4293 = n83 & new_n1512;
  assign new_n4294 = new_n4293 ^ new_n4292;
  assign new_n4295 = new_n4294 ^ new_n4291;
  assign new_n4296 = new_n4295 ^ n24;
  assign new_n4297 = new_n4296 ^ new_n4288;
  assign new_n4298 = new_n4091 ^ new_n4079;
  assign new_n4299 = ~new_n4088 & new_n4298;
  assign new_n4300 = new_n4299 ^ new_n4091;
  assign new_n4301 = new_n4300 ^ new_n4297;
  assign new_n4302 = ~new_n1198 & n87;
  assign new_n4303 = new_n1193 & new_n1940;
  assign new_n4304 = new_n4303 ^ new_n4302;
  assign new_n4305 = n88 & new_n1192;
  assign new_n4306 = n86 & new_n1204;
  assign new_n4307 = new_n4306 ^ new_n4305;
  assign new_n4308 = new_n4307 ^ new_n4304;
  assign new_n4309 = new_n4308 ^ n21;
  assign new_n4310 = new_n4309 ^ new_n4301;
  assign new_n4311 = new_n4104 ^ new_n4092;
  assign new_n4312 = ~new_n4101 & new_n4311;
  assign new_n4313 = new_n4312 ^ new_n4104;
  assign new_n4314 = new_n4313 ^ new_n4310;
  assign new_n4315 = ~new_n930 & n90;
  assign new_n4316 = new_n925 & new_n2341;
  assign new_n4317 = new_n4316 ^ new_n4315;
  assign new_n4318 = n91 & new_n924;
  assign new_n4319 = n89 & new_n936;
  assign new_n4320 = new_n4319 ^ new_n4318;
  assign new_n4321 = new_n4320 ^ new_n4317;
  assign new_n4322 = new_n4321 ^ n18;
  assign new_n4323 = new_n4322 ^ new_n4314;
  assign new_n4324 = new_n4117 ^ new_n4105;
  assign new_n4325 = ~new_n4114 & new_n4324;
  assign new_n4326 = new_n4325 ^ new_n4117;
  assign new_n4327 = new_n4326 ^ new_n4323;
  assign new_n4328 = n93 & new_n707;
  assign new_n4329 = new_n701 & new_n2785;
  assign new_n4330 = new_n4329 ^ new_n4328;
  assign new_n4331 = n94 & new_n700;
  assign new_n4332 = n92 & new_n787;
  assign new_n4333 = new_n4332 ^ new_n4331;
  assign new_n4334 = new_n4333 ^ new_n4330;
  assign new_n4335 = new_n4334 ^ n15;
  assign new_n4336 = new_n4335 ^ new_n4327;
  assign new_n4337 = new_n4130 ^ new_n4118;
  assign new_n4338 = ~new_n4127 & new_n4337;
  assign new_n4339 = new_n4338 ^ new_n4130;
  assign new_n4340 = new_n4339 ^ new_n4336;
  assign new_n4341 = n96 & new_n499;
  assign new_n4342 = ~new_n506 & new_n3273;
  assign new_n4343 = new_n4342 ^ new_n4341;
  assign new_n4344 = ~new_n505 & n97;
  assign new_n4345 = n95 & new_n579;
  assign new_n4346 = new_n4345 ^ new_n4344;
  assign new_n4347 = new_n4346 ^ new_n4343;
  assign new_n4348 = new_n4347 ^ n12;
  assign new_n4349 = new_n4348 ^ new_n4340;
  assign new_n4350 = new_n4143 ^ new_n4131;
  assign new_n4351 = ~new_n4140 & new_n4350;
  assign new_n4352 = new_n4351 ^ new_n4143;
  assign new_n4353 = new_n4352 ^ new_n4349;
  assign new_n4354 = n99 & new_n354;
  assign new_n4355 = new_n349 & new_n3789;
  assign new_n4356 = new_n4355 ^ new_n4354;
  assign new_n4357 = n100 & new_n348;
  assign new_n4358 = n98 & new_n391;
  assign new_n4359 = new_n4358 ^ new_n4357;
  assign new_n4360 = new_n4359 ^ new_n4356;
  assign new_n4361 = new_n4360 ^ n9;
  assign new_n4362 = new_n4361 ^ new_n4353;
  assign new_n4363 = new_n4156 ^ new_n4144;
  assign new_n4364 = ~new_n4153 & new_n4363;
  assign new_n4365 = new_n4364 ^ new_n4156;
  assign new_n4366 = new_n4365 ^ new_n4362;
  assign new_n4367 = n102 & new_n218;
  assign new_n4368 = new_n3811 ^ n103;
  assign new_n4369 = new_n208 & new_n4368;
  assign new_n4370 = new_n4369 ^ new_n4367;
  assign new_n4371 = n103 & new_n207;
  assign new_n4372 = n101 & new_n212;
  assign new_n4373 = new_n4372 ^ new_n4371;
  assign new_n4374 = new_n4373 ^ new_n4370;
  assign new_n4375 = new_n4374 ^ n6;
  assign new_n4376 = new_n4375 ^ new_n4366;
  assign new_n4377 = new_n4170 ^ new_n4157;
  assign new_n4378 = ~new_n4167 & new_n4377;
  assign new_n4379 = new_n4378 ^ new_n4170;
  assign new_n4380 = new_n4379 ^ new_n4376;
  assign new_n4381 = n104 & new_n180;
  assign new_n4382 = n2 & n105;
  assign new_n4383 = new_n4382 ^ new_n4381;
  assign new_n4384 = new_n4383 ^ n3;
  assign new_n4385 = ~n105 & ~new_n4173;
  assign new_n4386 = ~new_n4172 & n105;
  assign new_n4387 = new_n4386 ^ new_n4385;
  assign new_n4388 = new_n155 & new_n4387;
  assign new_n4389 = new_n4388 ^ n2;
  assign new_n4390 = new_n4389 ^ n106;
  assign new_n4391 = new_n4390 ^ new_n4384;
  assign new_n4392 = ~n1 & new_n4391;
  assign new_n4393 = new_n4392 ^ new_n4390;
  assign new_n4394 = new_n4393 ^ new_n4380;
  assign new_n4395 = new_n4189 ^ new_n4171;
  assign new_n4396 = ~new_n4186 & new_n4395;
  assign new_n4397 = new_n4396 ^ new_n4189;
  assign new_n4398 = new_n4397 ^ new_n4394;
  assign new_n4399 = ~new_n4214 & ~new_n4230;
  assign new_n4400 = ~new_n4399 & n42;
  assign new_n4401 = ~new_n154 & ~new_n4199;
  assign new_n4402 = new_n4401 ^ new_n259;
  assign new_n4403 = ~new_n4402 & new_n3837;
  assign new_n4404 = n66 & new_n4206;
  assign new_n4405 = ~new_n4212 & n67;
  assign new_n4406 = new_n4405 ^ new_n4404;
  assign new_n4407 = ~new_n4403 & ~new_n4406;
  assign new_n4408 = new_n4407 ^ new_n4400;
  assign new_n4409 = n43 ^ n42;
  assign new_n4410 = n65 & new_n4409;
  assign new_n4411 = new_n4410 ^ new_n4408;
  assign new_n4412 = ~new_n3682 & n70;
  assign new_n4413 = ~new_n402 & new_n3677;
  assign new_n4414 = new_n4413 ^ new_n4412;
  assign new_n4415 = n71 & new_n3676;
  assign new_n4416 = n69 & new_n3688;
  assign new_n4417 = new_n4416 ^ new_n4415;
  assign new_n4418 = new_n4417 ^ new_n4414;
  assign new_n4419 = new_n4418 ^ n39;
  assign new_n4420 = new_n4419 ^ new_n4411;
  assign new_n4421 = new_n4235 ^ new_n4198;
  assign new_n4422 = ~new_n4232 & new_n4421;
  assign new_n4423 = new_n4422 ^ new_n4235;
  assign new_n4424 = new_n4423 ^ new_n4420;
  assign new_n4425 = ~new_n3143 & n73;
  assign new_n4426 = new_n595 & new_n3138;
  assign new_n4427 = new_n4426 ^ new_n4425;
  assign new_n4428 = n74 & new_n3137;
  assign new_n4429 = n72 & new_n3149;
  assign new_n4430 = new_n4429 ^ new_n4428;
  assign new_n4431 = new_n4430 ^ new_n4427;
  assign new_n4432 = new_n4431 ^ n36;
  assign new_n4433 = new_n4432 ^ new_n4424;
  assign new_n4434 = new_n4248 ^ new_n4236;
  assign new_n4435 = ~new_n4245 & new_n4434;
  assign new_n4436 = new_n4435 ^ new_n4248;
  assign new_n4437 = new_n4436 ^ new_n4433;
  assign new_n4438 = ~new_n2672 & n76;
  assign new_n4439 = ~new_n812 & new_n2667;
  assign new_n4440 = new_n4439 ^ new_n4438;
  assign new_n4441 = n77 & new_n2666;
  assign new_n4442 = n75 & new_n2664;
  assign new_n4443 = new_n4442 ^ new_n4441;
  assign new_n4444 = new_n4443 ^ new_n4440;
  assign new_n4445 = new_n4444 ^ n33;
  assign new_n4446 = new_n4445 ^ new_n4437;
  assign new_n4447 = new_n4261 ^ new_n4249;
  assign new_n4448 = ~new_n4258 & new_n4447;
  assign new_n4449 = new_n4448 ^ new_n4261;
  assign new_n4450 = new_n4449 ^ new_n4446;
  assign new_n4451 = n79 & new_n2246;
  assign new_n4452 = new_n1069 & new_n2241;
  assign new_n4453 = new_n4452 ^ new_n4451;
  assign new_n4454 = n80 & new_n2240;
  assign new_n4455 = n78 & new_n2391;
  assign new_n4456 = new_n4455 ^ new_n4454;
  assign new_n4457 = new_n4456 ^ new_n4453;
  assign new_n4458 = new_n4457 ^ n30;
  assign new_n4459 = new_n4458 ^ new_n4450;
  assign new_n4460 = new_n4274 ^ new_n4262;
  assign new_n4461 = ~new_n4271 & new_n4460;
  assign new_n4462 = new_n4461 ^ new_n4274;
  assign new_n4463 = new_n4462 ^ new_n4459;
  assign new_n4464 = n82 & new_n1874;
  assign new_n4465 = new_n1363 & new_n1864;
  assign new_n4466 = new_n4465 ^ new_n4464;
  assign new_n4467 = n83 & new_n1863;
  assign new_n4468 = n81 & new_n1868;
  assign new_n4469 = new_n4468 ^ new_n4467;
  assign new_n4470 = new_n4469 ^ new_n4466;
  assign new_n4471 = new_n4470 ^ n27;
  assign new_n4472 = new_n4471 ^ new_n4463;
  assign new_n4473 = new_n4287 ^ new_n4275;
  assign new_n4474 = ~new_n4284 & new_n4473;
  assign new_n4475 = new_n4474 ^ new_n4287;
  assign new_n4476 = new_n4475 ^ new_n4472;
  assign new_n4477 = ~new_n1506 & n85;
  assign new_n4478 = new_n1501 & new_n1694;
  assign new_n4479 = new_n4478 ^ new_n4477;
  assign new_n4480 = n86 & new_n1500;
  assign new_n4481 = n84 & new_n1512;
  assign new_n4482 = new_n4481 ^ new_n4480;
  assign new_n4483 = new_n4482 ^ new_n4479;
  assign new_n4484 = new_n4483 ^ n24;
  assign new_n4485 = new_n4484 ^ new_n4476;
  assign new_n4486 = new_n4300 ^ new_n4288;
  assign new_n4487 = ~new_n4297 & new_n4486;
  assign new_n4488 = new_n4487 ^ new_n4300;
  assign new_n4489 = new_n4488 ^ new_n4485;
  assign new_n4490 = ~new_n1198 & n88;
  assign new_n4491 = new_n1193 & new_n2063;
  assign new_n4492 = new_n4491 ^ new_n4490;
  assign new_n4493 = n89 & new_n1192;
  assign new_n4494 = n87 & new_n1204;
  assign new_n4495 = new_n4494 ^ new_n4493;
  assign new_n4496 = new_n4495 ^ new_n4492;
  assign new_n4497 = new_n4496 ^ n21;
  assign new_n4498 = new_n4497 ^ new_n4489;
  assign new_n4499 = new_n4313 ^ new_n4301;
  assign new_n4500 = ~new_n4310 & new_n4499;
  assign new_n4501 = new_n4500 ^ new_n4313;
  assign new_n4502 = new_n4501 ^ new_n4498;
  assign new_n4503 = ~new_n930 & n91;
  assign new_n4504 = new_n925 & new_n2481;
  assign new_n4505 = new_n4504 ^ new_n4503;
  assign new_n4506 = n92 & new_n924;
  assign new_n4507 = n90 & new_n936;
  assign new_n4508 = new_n4507 ^ new_n4506;
  assign new_n4509 = new_n4508 ^ new_n4505;
  assign new_n4510 = new_n4509 ^ n18;
  assign new_n4511 = new_n4510 ^ new_n4502;
  assign new_n4512 = new_n4326 ^ new_n4314;
  assign new_n4513 = ~new_n4323 & new_n4512;
  assign new_n4514 = new_n4513 ^ new_n4326;
  assign new_n4515 = new_n4514 ^ new_n4511;
  assign new_n4516 = n94 & new_n707;
  assign new_n4517 = new_n701 & new_n2934;
  assign new_n4518 = new_n4517 ^ new_n4516;
  assign new_n4519 = n95 & new_n700;
  assign new_n4520 = n93 & new_n787;
  assign new_n4521 = new_n4520 ^ new_n4519;
  assign new_n4522 = new_n4521 ^ new_n4518;
  assign new_n4523 = new_n4522 ^ n15;
  assign new_n4524 = new_n4523 ^ new_n4515;
  assign new_n4525 = new_n4339 ^ new_n4327;
  assign new_n4526 = ~new_n4336 & new_n4525;
  assign new_n4527 = new_n4526 ^ new_n4339;
  assign new_n4528 = new_n4527 ^ new_n4524;
  assign new_n4529 = n97 & new_n499;
  assign new_n4530 = ~new_n506 & new_n3435;
  assign new_n4531 = new_n4530 ^ new_n4529;
  assign new_n4532 = ~new_n505 & n98;
  assign new_n4533 = n96 & new_n579;
  assign new_n4534 = new_n4533 ^ new_n4532;
  assign new_n4535 = new_n4534 ^ new_n4531;
  assign new_n4536 = new_n4535 ^ n12;
  assign new_n4537 = new_n4536 ^ new_n4528;
  assign new_n4538 = new_n4352 ^ new_n4340;
  assign new_n4539 = ~new_n4349 & new_n4538;
  assign new_n4540 = new_n4539 ^ new_n4352;
  assign new_n4541 = new_n4540 ^ new_n4537;
  assign new_n4542 = n100 & new_n354;
  assign new_n4543 = new_n349 & new_n3972;
  assign new_n4544 = new_n4543 ^ new_n4542;
  assign new_n4545 = n101 & new_n348;
  assign new_n4546 = n99 & new_n391;
  assign new_n4547 = new_n4546 ^ new_n4545;
  assign new_n4548 = new_n4547 ^ new_n4544;
  assign new_n4549 = new_n4548 ^ n9;
  assign new_n4550 = new_n4549 ^ new_n4541;
  assign new_n4551 = new_n4365 ^ new_n4353;
  assign new_n4552 = ~new_n4362 & new_n4551;
  assign new_n4553 = new_n4552 ^ new_n4365;
  assign new_n4554 = new_n4553 ^ new_n4550;
  assign new_n4555 = n103 & new_n218;
  assign new_n4556 = new_n3989 ^ n104;
  assign new_n4557 = ~new_n4556 & new_n208;
  assign new_n4558 = new_n4557 ^ new_n4555;
  assign new_n4559 = n104 & new_n207;
  assign new_n4560 = n102 & new_n212;
  assign new_n4561 = new_n4560 ^ new_n4559;
  assign new_n4562 = new_n4561 ^ new_n4558;
  assign new_n4563 = new_n4562 ^ n6;
  assign new_n4564 = new_n4563 ^ new_n4554;
  assign new_n4565 = new_n4379 ^ new_n4366;
  assign new_n4566 = ~new_n4376 & new_n4565;
  assign new_n4567 = new_n4566 ^ new_n4379;
  assign new_n4568 = new_n4567 ^ new_n4564;
  assign new_n4569 = n106 ^ n3;
  assign new_n4570 = ~n105 & n3;
  assign new_n4571 = new_n4570 ^ new_n4569;
  assign new_n4572 = ~n2 & new_n4571;
  assign new_n4573 = new_n4572 ^ new_n4569;
  assign new_n4574 = ~n106 & ~new_n4386;
  assign new_n4575 = ~new_n4385 & n106;
  assign new_n4576 = new_n4575 ^ new_n4574;
  assign new_n4577 = new_n155 & new_n4576;
  assign new_n4578 = new_n4577 ^ n2;
  assign new_n4579 = new_n4578 ^ n107;
  assign new_n4580 = new_n4579 ^ new_n4573;
  assign new_n4581 = ~n1 & new_n4580;
  assign new_n4582 = new_n4581 ^ new_n4579;
  assign new_n4583 = new_n4582 ^ new_n4568;
  assign new_n4584 = new_n4397 ^ new_n4380;
  assign new_n4585 = ~new_n4394 & new_n4584;
  assign new_n4586 = new_n4585 ^ new_n4397;
  assign new_n4587 = new_n4586 ^ new_n4583;
  assign new_n4588 = ~new_n4408 & ~new_n4410;
  assign new_n4589 = new_n4407 ^ n42;
  assign new_n4590 = ~new_n4588 & ~new_n4589;
  assign new_n4591 = n66 ^ n43;
  assign new_n4592 = ~new_n4591 & new_n4409;
  assign new_n4593 = new_n4592 ^ n42;
  assign new_n4594 = new_n4593 ^ n44;
  assign new_n4595 = ~n42 & ~n43;
  assign new_n4596 = new_n4595 ^ new_n4409;
  assign new_n4597 = new_n4596 ^ n44;
  assign new_n4598 = ~n65 & ~new_n4597;
  assign new_n4599 = new_n4598 ^ new_n4594;
  assign new_n4600 = new_n4599 ^ new_n4590;
  assign new_n4601 = ~new_n4212 & n68;
  assign new_n4602 = ~new_n304 & new_n4201;
  assign new_n4603 = new_n4602 ^ new_n4601;
  assign new_n4604 = n69 & new_n4200;
  assign new_n4605 = n67 & new_n4206;
  assign new_n4606 = new_n4605 ^ new_n4604;
  assign new_n4607 = new_n4606 ^ new_n4603;
  assign new_n4608 = new_n4607 ^ n42;
  assign new_n4609 = new_n4608 ^ new_n4600;
  assign new_n4610 = ~new_n3682 & n71;
  assign new_n4611 = ~new_n459 & new_n3677;
  assign new_n4612 = new_n4611 ^ new_n4610;
  assign new_n4613 = n72 & new_n3676;
  assign new_n4614 = n70 & new_n3688;
  assign new_n4615 = new_n4614 ^ new_n4613;
  assign new_n4616 = new_n4615 ^ new_n4612;
  assign new_n4617 = new_n4616 ^ n39;
  assign new_n4618 = new_n4617 ^ new_n4609;
  assign new_n4619 = new_n4423 ^ new_n4411;
  assign new_n4620 = ~new_n4619 & new_n4420;
  assign new_n4621 = new_n4620 ^ new_n4423;
  assign new_n4622 = new_n4621 ^ new_n4618;
  assign new_n4623 = ~new_n3143 & n74;
  assign new_n4624 = new_n660 & new_n3138;
  assign new_n4625 = new_n4624 ^ new_n4623;
  assign new_n4626 = n75 & new_n3137;
  assign new_n4627 = n73 & new_n3149;
  assign new_n4628 = new_n4627 ^ new_n4626;
  assign new_n4629 = new_n4628 ^ new_n4625;
  assign new_n4630 = new_n4629 ^ n36;
  assign new_n4631 = new_n4630 ^ new_n4622;
  assign new_n4632 = new_n4436 ^ new_n4424;
  assign new_n4633 = ~new_n4632 & new_n4433;
  assign new_n4634 = new_n4633 ^ new_n4436;
  assign new_n4635 = new_n4634 ^ new_n4631;
  assign new_n4636 = ~new_n2672 & n77;
  assign new_n4637 = ~new_n891 & new_n2667;
  assign new_n4638 = new_n4637 ^ new_n4636;
  assign new_n4639 = n78 & new_n2666;
  assign new_n4640 = n76 & new_n2664;
  assign new_n4641 = new_n4640 ^ new_n4639;
  assign new_n4642 = new_n4641 ^ new_n4638;
  assign new_n4643 = new_n4642 ^ n33;
  assign new_n4644 = new_n4643 ^ new_n4635;
  assign new_n4645 = new_n4449 ^ new_n4437;
  assign new_n4646 = ~new_n4645 & new_n4446;
  assign new_n4647 = new_n4646 ^ new_n4449;
  assign new_n4648 = new_n4647 ^ new_n4644;
  assign new_n4649 = n80 & new_n2246;
  assign new_n4650 = new_n1161 & new_n2241;
  assign new_n4651 = new_n4650 ^ new_n4649;
  assign new_n4652 = n81 & new_n2240;
  assign new_n4653 = n79 & new_n2391;
  assign new_n4654 = new_n4653 ^ new_n4652;
  assign new_n4655 = new_n4654 ^ new_n4651;
  assign new_n4656 = new_n4655 ^ n30;
  assign new_n4657 = new_n4656 ^ new_n4648;
  assign new_n4658 = new_n4462 ^ new_n4450;
  assign new_n4659 = ~new_n4658 & new_n4459;
  assign new_n4660 = new_n4659 ^ new_n4462;
  assign new_n4661 = new_n4660 ^ new_n4657;
  assign new_n4662 = n83 & new_n1874;
  assign new_n4663 = new_n1468 & new_n1864;
  assign new_n4664 = new_n4663 ^ new_n4662;
  assign new_n4665 = n84 & new_n1863;
  assign new_n4666 = n82 & new_n1868;
  assign new_n4667 = new_n4666 ^ new_n4665;
  assign new_n4668 = new_n4667 ^ new_n4664;
  assign new_n4669 = new_n4668 ^ n27;
  assign new_n4670 = new_n4669 ^ new_n4661;
  assign new_n4671 = new_n4475 ^ new_n4463;
  assign new_n4672 = ~new_n4671 & new_n4472;
  assign new_n4673 = new_n4672 ^ new_n4475;
  assign new_n4674 = new_n4673 ^ new_n4670;
  assign new_n4675 = ~new_n1506 & n86;
  assign new_n4676 = new_n1501 & new_n1811;
  assign new_n4677 = new_n4676 ^ new_n4675;
  assign new_n4678 = n87 & new_n1500;
  assign new_n4679 = n85 & new_n1512;
  assign new_n4680 = new_n4679 ^ new_n4678;
  assign new_n4681 = new_n4680 ^ new_n4677;
  assign new_n4682 = new_n4681 ^ n24;
  assign new_n4683 = new_n4682 ^ new_n4674;
  assign new_n4684 = new_n4488 ^ new_n4476;
  assign new_n4685 = ~new_n4684 & new_n4485;
  assign new_n4686 = new_n4685 ^ new_n4488;
  assign new_n4687 = new_n4686 ^ new_n4683;
  assign new_n4688 = ~new_n1198 & n89;
  assign new_n4689 = new_n1193 & new_n2193;
  assign new_n4690 = new_n4689 ^ new_n4688;
  assign new_n4691 = n90 & new_n1192;
  assign new_n4692 = n88 & new_n1204;
  assign new_n4693 = new_n4692 ^ new_n4691;
  assign new_n4694 = new_n4693 ^ new_n4690;
  assign new_n4695 = new_n4694 ^ n21;
  assign new_n4696 = new_n4695 ^ new_n4687;
  assign new_n4697 = new_n4501 ^ new_n4489;
  assign new_n4698 = ~new_n4697 & new_n4498;
  assign new_n4699 = new_n4698 ^ new_n4501;
  assign new_n4700 = new_n4699 ^ new_n4696;
  assign new_n4701 = ~new_n930 & n92;
  assign new_n4702 = new_n925 & new_n2628;
  assign new_n4703 = new_n4702 ^ new_n4701;
  assign new_n4704 = n93 & new_n924;
  assign new_n4705 = n91 & new_n936;
  assign new_n4706 = new_n4705 ^ new_n4704;
  assign new_n4707 = new_n4706 ^ new_n4703;
  assign new_n4708 = new_n4707 ^ n18;
  assign new_n4709 = new_n4708 ^ new_n4700;
  assign new_n4710 = new_n4514 ^ new_n4502;
  assign new_n4711 = ~new_n4710 & new_n4511;
  assign new_n4712 = new_n4711 ^ new_n4514;
  assign new_n4713 = new_n4712 ^ new_n4709;
  assign new_n4714 = n95 & new_n707;
  assign new_n4715 = new_n701 & new_n3095;
  assign new_n4716 = new_n4715 ^ new_n4714;
  assign new_n4717 = n96 & new_n700;
  assign new_n4718 = n94 & new_n787;
  assign new_n4719 = new_n4718 ^ new_n4717;
  assign new_n4720 = new_n4719 ^ new_n4716;
  assign new_n4721 = new_n4720 ^ n15;
  assign new_n4722 = new_n4721 ^ new_n4713;
  assign new_n4723 = new_n4527 ^ new_n4515;
  assign new_n4724 = ~new_n4723 & new_n4524;
  assign new_n4725 = new_n4724 ^ new_n4527;
  assign new_n4726 = new_n4725 ^ new_n4722;
  assign new_n4727 = n98 & new_n499;
  assign new_n4728 = ~new_n506 & new_n3604;
  assign new_n4729 = new_n4728 ^ new_n4727;
  assign new_n4730 = n97 & new_n579;
  assign new_n4731 = ~new_n505 & n99;
  assign new_n4732 = new_n4731 ^ new_n4730;
  assign new_n4733 = new_n4732 ^ new_n4729;
  assign new_n4734 = new_n4733 ^ n12;
  assign new_n4735 = new_n4734 ^ new_n4726;
  assign new_n4736 = new_n4540 ^ new_n4528;
  assign new_n4737 = ~new_n4736 & new_n4537;
  assign new_n4738 = new_n4737 ^ new_n4540;
  assign new_n4739 = new_n4738 ^ new_n4735;
  assign new_n4740 = n101 & new_n354;
  assign new_n4741 = new_n349 & new_n4159;
  assign new_n4742 = new_n4741 ^ new_n4740;
  assign new_n4743 = n102 & new_n348;
  assign new_n4744 = n100 & new_n391;
  assign new_n4745 = new_n4744 ^ new_n4743;
  assign new_n4746 = new_n4745 ^ new_n4742;
  assign new_n4747 = new_n4746 ^ n9;
  assign new_n4748 = new_n4747 ^ new_n4739;
  assign new_n4749 = new_n4553 ^ new_n4541;
  assign new_n4750 = ~new_n4749 & new_n4550;
  assign new_n4751 = new_n4750 ^ new_n4553;
  assign new_n4752 = new_n4751 ^ new_n4748;
  assign new_n4753 = n104 & new_n218;
  assign new_n4754 = new_n4174 ^ n105;
  assign new_n4755 = ~new_n4754 & new_n208;
  assign new_n4756 = new_n4755 ^ new_n4753;
  assign new_n4757 = n105 & new_n207;
  assign new_n4758 = n103 & new_n212;
  assign new_n4759 = new_n4758 ^ new_n4757;
  assign new_n4760 = new_n4759 ^ new_n4756;
  assign new_n4761 = new_n4760 ^ n6;
  assign new_n4762 = new_n4761 ^ new_n4752;
  assign new_n4763 = new_n4567 ^ new_n4554;
  assign new_n4764 = ~new_n4763 & new_n4564;
  assign new_n4765 = new_n4764 ^ new_n4567;
  assign new_n4766 = new_n4765 ^ new_n4762;
  assign new_n4767 = n106 & new_n180;
  assign new_n4768 = n2 & n107;
  assign new_n4769 = new_n4768 ^ new_n4767;
  assign new_n4770 = new_n4769 ^ n3;
  assign new_n4771 = ~new_n4574 & n107;
  assign new_n4772 = ~n107 & ~new_n4575;
  assign new_n4773 = new_n4772 ^ new_n4771;
  assign new_n4774 = new_n155 & new_n4773;
  assign new_n4775 = new_n4774 ^ n2;
  assign new_n4776 = new_n4775 ^ n108;
  assign new_n4777 = new_n4776 ^ new_n4770;
  assign new_n4778 = ~n1 & new_n4777;
  assign new_n4779 = new_n4778 ^ new_n4776;
  assign new_n4780 = new_n4779 ^ new_n4766;
  assign new_n4781 = new_n4586 ^ new_n4568;
  assign new_n4782 = ~new_n4781 & new_n4583;
  assign new_n4783 = new_n4782 ^ new_n4586;
  assign new_n4784 = new_n4783 ^ new_n4780;
  assign new_n4785 = ~new_n3143 & n75;
  assign new_n4786 = ~new_n737 & new_n3138;
  assign new_n4787 = new_n4786 ^ new_n4785;
  assign new_n4788 = n76 & new_n3137;
  assign new_n4789 = n74 & new_n3149;
  assign new_n4790 = new_n4789 ^ new_n4788;
  assign new_n4791 = new_n4790 ^ new_n4787;
  assign new_n4792 = new_n4791 ^ n36;
  assign new_n4793 = new_n4634 ^ new_n4622;
  assign new_n4794 = ~new_n4631 & new_n4793;
  assign new_n4795 = new_n4794 ^ new_n4634;
  assign new_n4796 = new_n4795 ^ new_n4792;
  assign new_n4797 = n45 ^ n44;
  assign new_n4798 = ~new_n4797 & new_n4409;
  assign new_n4799 = new_n4798 ^ new_n4409;
  assign new_n4800 = ~new_n151 & new_n4799;
  assign new_n4801 = n67 & new_n4409;
  assign new_n4802 = new_n4801 ^ new_n4800;
  assign new_n4803 = ~new_n4409 & n44;
  assign new_n4804 = new_n4803 ^ new_n4596;
  assign new_n4805 = ~new_n4804 & n66;
  assign new_n4806 = new_n4805 ^ new_n4802;
  assign new_n4807 = new_n4806 ^ n45;
  assign new_n4808 = ~new_n4409 & n45;
  assign new_n4809 = new_n4808 ^ new_n4596;
  assign new_n4810 = ~new_n4809 & new_n4797;
  assign new_n4811 = n65 & new_n4810;
  assign new_n4812 = new_n4811 ^ new_n4807;
  assign new_n4813 = ~new_n4410 & ~new_n4599;
  assign new_n4814 = n45 & new_n4813;
  assign new_n4815 = new_n4814 ^ new_n4812;
  assign new_n4816 = ~new_n4212 & n69;
  assign new_n4817 = ~new_n339 & new_n4201;
  assign new_n4818 = new_n4817 ^ new_n4816;
  assign new_n4819 = n70 & new_n4200;
  assign new_n4820 = n68 & new_n4206;
  assign new_n4821 = new_n4820 ^ new_n4819;
  assign new_n4822 = new_n4821 ^ new_n4818;
  assign new_n4823 = new_n4822 ^ n42;
  assign new_n4824 = new_n4823 ^ new_n4815;
  assign new_n4825 = new_n4608 ^ new_n4599;
  assign new_n4826 = ~new_n4825 & new_n4600;
  assign new_n4827 = new_n4826 ^ new_n4590;
  assign new_n4828 = new_n4827 ^ new_n4824;
  assign new_n4829 = ~new_n3682 & n72;
  assign new_n4830 = new_n534 & new_n3677;
  assign new_n4831 = new_n4830 ^ new_n4829;
  assign new_n4832 = n73 & new_n3676;
  assign new_n4833 = n71 & new_n3688;
  assign new_n4834 = new_n4833 ^ new_n4832;
  assign new_n4835 = new_n4834 ^ new_n4831;
  assign new_n4836 = new_n4835 ^ n39;
  assign new_n4837 = new_n4836 ^ new_n4828;
  assign new_n4838 = new_n4621 ^ new_n4609;
  assign new_n4839 = ~new_n4618 & new_n4838;
  assign new_n4840 = new_n4839 ^ new_n4621;
  assign new_n4841 = new_n4840 ^ new_n4837;
  assign new_n4842 = new_n4841 ^ new_n4796;
  assign new_n4843 = ~new_n2672 & n78;
  assign new_n4844 = ~new_n982 & new_n2667;
  assign new_n4845 = new_n4844 ^ new_n4843;
  assign new_n4846 = n79 & new_n2666;
  assign new_n4847 = n77 & new_n2664;
  assign new_n4848 = new_n4847 ^ new_n4846;
  assign new_n4849 = new_n4848 ^ new_n4845;
  assign new_n4850 = new_n4849 ^ n33;
  assign new_n4851 = new_n4850 ^ new_n4842;
  assign new_n4852 = new_n4647 ^ new_n4635;
  assign new_n4853 = ~new_n4644 & new_n4852;
  assign new_n4854 = new_n4853 ^ new_n4647;
  assign new_n4855 = new_n4854 ^ new_n4851;
  assign new_n4856 = n81 & new_n2246;
  assign new_n4857 = new_n1263 & new_n2241;
  assign new_n4858 = new_n4857 ^ new_n4856;
  assign new_n4859 = n82 & new_n2240;
  assign new_n4860 = n80 & new_n2391;
  assign new_n4861 = new_n4860 ^ new_n4859;
  assign new_n4862 = new_n4861 ^ new_n4858;
  assign new_n4863 = new_n4862 ^ n30;
  assign new_n4864 = new_n4863 ^ new_n4855;
  assign new_n4865 = new_n4660 ^ new_n4648;
  assign new_n4866 = ~new_n4657 & new_n4865;
  assign new_n4867 = new_n4866 ^ new_n4660;
  assign new_n4868 = new_n4867 ^ new_n4864;
  assign new_n4869 = n84 & new_n1874;
  assign new_n4870 = new_n1584 & new_n1864;
  assign new_n4871 = new_n4870 ^ new_n4869;
  assign new_n4872 = n85 & new_n1863;
  assign new_n4873 = n83 & new_n1868;
  assign new_n4874 = new_n4873 ^ new_n4872;
  assign new_n4875 = new_n4874 ^ new_n4871;
  assign new_n4876 = new_n4875 ^ n27;
  assign new_n4877 = new_n4876 ^ new_n4868;
  assign new_n4878 = new_n4673 ^ new_n4661;
  assign new_n4879 = ~new_n4670 & new_n4878;
  assign new_n4880 = new_n4879 ^ new_n4673;
  assign new_n4881 = new_n4880 ^ new_n4877;
  assign new_n4882 = ~new_n1506 & n87;
  assign new_n4883 = new_n1501 & new_n1940;
  assign new_n4884 = new_n4883 ^ new_n4882;
  assign new_n4885 = n88 & new_n1500;
  assign new_n4886 = n86 & new_n1512;
  assign new_n4887 = new_n4886 ^ new_n4885;
  assign new_n4888 = new_n4887 ^ new_n4884;
  assign new_n4889 = new_n4888 ^ n24;
  assign new_n4890 = new_n4889 ^ new_n4881;
  assign new_n4891 = new_n4686 ^ new_n4674;
  assign new_n4892 = ~new_n4683 & new_n4891;
  assign new_n4893 = new_n4892 ^ new_n4686;
  assign new_n4894 = new_n4893 ^ new_n4890;
  assign new_n4895 = ~new_n1198 & n90;
  assign new_n4896 = new_n1193 & new_n2341;
  assign new_n4897 = new_n4896 ^ new_n4895;
  assign new_n4898 = n91 & new_n1192;
  assign new_n4899 = n89 & new_n1204;
  assign new_n4900 = new_n4899 ^ new_n4898;
  assign new_n4901 = new_n4900 ^ new_n4897;
  assign new_n4902 = new_n4901 ^ n21;
  assign new_n4903 = new_n4902 ^ new_n4894;
  assign new_n4904 = new_n4699 ^ new_n4687;
  assign new_n4905 = ~new_n4696 & new_n4904;
  assign new_n4906 = new_n4905 ^ new_n4699;
  assign new_n4907 = new_n4906 ^ new_n4903;
  assign new_n4908 = ~new_n930 & n93;
  assign new_n4909 = new_n925 & new_n2785;
  assign new_n4910 = new_n4909 ^ new_n4908;
  assign new_n4911 = n94 & new_n924;
  assign new_n4912 = n92 & new_n936;
  assign new_n4913 = new_n4912 ^ new_n4911;
  assign new_n4914 = new_n4913 ^ new_n4910;
  assign new_n4915 = new_n4914 ^ n18;
  assign new_n4916 = new_n4915 ^ new_n4907;
  assign new_n4917 = new_n4712 ^ new_n4700;
  assign new_n4918 = ~new_n4709 & new_n4917;
  assign new_n4919 = new_n4918 ^ new_n4712;
  assign new_n4920 = new_n4919 ^ new_n4916;
  assign new_n4921 = n96 & new_n707;
  assign new_n4922 = new_n701 & new_n3273;
  assign new_n4923 = new_n4922 ^ new_n4921;
  assign new_n4924 = n97 & new_n700;
  assign new_n4925 = n95 & new_n787;
  assign new_n4926 = new_n4925 ^ new_n4924;
  assign new_n4927 = new_n4926 ^ new_n4923;
  assign new_n4928 = new_n4927 ^ n15;
  assign new_n4929 = new_n4928 ^ new_n4920;
  assign new_n4930 = new_n4725 ^ new_n4713;
  assign new_n4931 = ~new_n4722 & new_n4930;
  assign new_n4932 = new_n4931 ^ new_n4725;
  assign new_n4933 = new_n4932 ^ new_n4929;
  assign new_n4934 = n99 & new_n499;
  assign new_n4935 = ~new_n506 & new_n3789;
  assign new_n4936 = new_n4935 ^ new_n4934;
  assign new_n4937 = ~new_n505 & n100;
  assign new_n4938 = n98 & new_n579;
  assign new_n4939 = new_n4938 ^ new_n4937;
  assign new_n4940 = new_n4939 ^ new_n4936;
  assign new_n4941 = new_n4940 ^ n12;
  assign new_n4942 = new_n4941 ^ new_n4933;
  assign new_n4943 = new_n4738 ^ new_n4726;
  assign new_n4944 = ~new_n4735 & new_n4943;
  assign new_n4945 = new_n4944 ^ new_n4738;
  assign new_n4946 = new_n4945 ^ new_n4942;
  assign new_n4947 = n102 & new_n354;
  assign new_n4948 = new_n349 & new_n4368;
  assign new_n4949 = new_n4948 ^ new_n4947;
  assign new_n4950 = n103 & new_n348;
  assign new_n4951 = n101 & new_n391;
  assign new_n4952 = new_n4951 ^ new_n4950;
  assign new_n4953 = new_n4952 ^ new_n4949;
  assign new_n4954 = new_n4953 ^ n9;
  assign new_n4955 = new_n4954 ^ new_n4946;
  assign new_n4956 = new_n4751 ^ new_n4739;
  assign new_n4957 = ~new_n4748 & new_n4956;
  assign new_n4958 = new_n4957 ^ new_n4751;
  assign new_n4959 = new_n4958 ^ new_n4955;
  assign new_n4960 = n105 & new_n218;
  assign new_n4961 = new_n4387 ^ n106;
  assign new_n4962 = ~new_n4961 & new_n208;
  assign new_n4963 = new_n4962 ^ new_n4960;
  assign new_n4964 = n106 & new_n207;
  assign new_n4965 = n104 & new_n212;
  assign new_n4966 = new_n4965 ^ new_n4964;
  assign new_n4967 = new_n4966 ^ new_n4963;
  assign new_n4968 = new_n4967 ^ n6;
  assign new_n4969 = new_n4968 ^ new_n4959;
  assign new_n4970 = new_n4765 ^ new_n4752;
  assign new_n4971 = ~new_n4762 & new_n4970;
  assign new_n4972 = new_n4971 ^ new_n4765;
  assign new_n4973 = new_n4972 ^ new_n4969;
  assign new_n4974 = n108 ^ n107;
  assign new_n4975 = ~n108 & new_n4576;
  assign new_n4976 = new_n4975 ^ new_n4575;
  assign new_n4977 = ~new_n4976 & new_n4974;
  assign new_n4978 = ~new_n4977 & new_n155;
  assign new_n4979 = new_n4978 ^ n2;
  assign new_n4980 = new_n4979 ^ n109;
  assign new_n4981 = n108 ^ n3;
  assign new_n4982 = ~n107 & n3;
  assign new_n4983 = new_n4982 ^ new_n4981;
  assign new_n4984 = ~n2 & new_n4983;
  assign new_n4985 = new_n4984 ^ new_n4981;
  assign new_n4986 = new_n4985 ^ new_n4980;
  assign new_n4987 = ~n1 & new_n4986;
  assign new_n4988 = new_n4987 ^ new_n4980;
  assign new_n4989 = new_n4988 ^ new_n4973;
  assign new_n4990 = new_n4783 ^ new_n4766;
  assign new_n4991 = ~new_n4780 & new_n4990;
  assign new_n4992 = new_n4991 ^ new_n4783;
  assign new_n4993 = new_n4992 ^ new_n4989;
  assign new_n4994 = ~new_n3682 & n73;
  assign new_n4995 = new_n595 & new_n3677;
  assign new_n4996 = new_n4995 ^ new_n4994;
  assign new_n4997 = n74 & new_n3676;
  assign new_n4998 = n72 & new_n3688;
  assign new_n4999 = new_n4998 ^ new_n4997;
  assign new_n5000 = new_n4999 ^ new_n4996;
  assign new_n5001 = new_n5000 ^ n39;
  assign new_n5002 = new_n4840 ^ new_n4828;
  assign new_n5003 = ~new_n4837 & new_n5002;
  assign new_n5004 = new_n5003 ^ new_n4840;
  assign new_n5005 = new_n5004 ^ new_n5001;
  assign new_n5006 = new_n4812 & new_n4814;
  assign new_n5007 = ~new_n259 & new_n4799;
  assign new_n5008 = ~new_n4804 & n67;
  assign new_n5009 = new_n5008 ^ new_n5007;
  assign new_n5010 = n68 & new_n4798;
  assign new_n5011 = n66 & new_n4810;
  assign new_n5012 = new_n5011 ^ new_n5010;
  assign new_n5013 = new_n5012 ^ new_n5009;
  assign new_n5014 = new_n5013 ^ n45;
  assign new_n5015 = n46 ^ n45;
  assign new_n5016 = n65 & new_n5015;
  assign new_n5017 = new_n5016 ^ new_n5014;
  assign new_n5018 = new_n5017 ^ new_n5006;
  assign new_n5019 = ~new_n4212 & n70;
  assign new_n5020 = ~new_n402 & new_n4201;
  assign new_n5021 = new_n5020 ^ new_n5019;
  assign new_n5022 = n71 & new_n4200;
  assign new_n5023 = n69 & new_n4206;
  assign new_n5024 = new_n5023 ^ new_n5022;
  assign new_n5025 = new_n5024 ^ new_n5021;
  assign new_n5026 = new_n5025 ^ n42;
  assign new_n5027 = new_n5026 ^ new_n5018;
  assign new_n5028 = new_n4827 ^ new_n4815;
  assign new_n5029 = ~new_n4824 & new_n5028;
  assign new_n5030 = new_n5029 ^ new_n4827;
  assign new_n5031 = new_n5030 ^ new_n5027;
  assign new_n5032 = new_n5031 ^ new_n5005;
  assign new_n5033 = ~new_n3143 & n76;
  assign new_n5034 = ~new_n812 & new_n3138;
  assign new_n5035 = new_n5034 ^ new_n5033;
  assign new_n5036 = n77 & new_n3137;
  assign new_n5037 = n75 & new_n3149;
  assign new_n5038 = new_n5037 ^ new_n5036;
  assign new_n5039 = new_n5038 ^ new_n5035;
  assign new_n5040 = new_n5039 ^ n36;
  assign new_n5041 = new_n5040 ^ new_n5032;
  assign new_n5042 = new_n4841 ^ new_n4792;
  assign new_n5043 = ~new_n5042 & new_n4796;
  assign new_n5044 = new_n5043 ^ new_n4795;
  assign new_n5045 = new_n5044 ^ new_n5041;
  assign new_n5046 = ~new_n2672 & n79;
  assign new_n5047 = new_n1069 & new_n2667;
  assign new_n5048 = new_n5047 ^ new_n5046;
  assign new_n5049 = n80 & new_n2666;
  assign new_n5050 = n78 & new_n2664;
  assign new_n5051 = new_n5050 ^ new_n5049;
  assign new_n5052 = new_n5051 ^ new_n5048;
  assign new_n5053 = new_n5052 ^ n33;
  assign new_n5054 = new_n5053 ^ new_n5045;
  assign new_n5055 = new_n4854 ^ new_n4842;
  assign new_n5056 = ~new_n4851 & new_n5055;
  assign new_n5057 = new_n5056 ^ new_n4854;
  assign new_n5058 = new_n5057 ^ new_n5054;
  assign new_n5059 = n82 & new_n2246;
  assign new_n5060 = new_n1363 & new_n2241;
  assign new_n5061 = new_n5060 ^ new_n5059;
  assign new_n5062 = n83 & new_n2240;
  assign new_n5063 = n81 & new_n2391;
  assign new_n5064 = new_n5063 ^ new_n5062;
  assign new_n5065 = new_n5064 ^ new_n5061;
  assign new_n5066 = new_n5065 ^ n30;
  assign new_n5067 = new_n5066 ^ new_n5058;
  assign new_n5068 = new_n4867 ^ new_n4855;
  assign new_n5069 = ~new_n4864 & new_n5068;
  assign new_n5070 = new_n5069 ^ new_n4867;
  assign new_n5071 = new_n5070 ^ new_n5067;
  assign new_n5072 = n85 & new_n1874;
  assign new_n5073 = new_n1694 & new_n1864;
  assign new_n5074 = new_n5073 ^ new_n5072;
  assign new_n5075 = n86 & new_n1863;
  assign new_n5076 = n84 & new_n1868;
  assign new_n5077 = new_n5076 ^ new_n5075;
  assign new_n5078 = new_n5077 ^ new_n5074;
  assign new_n5079 = new_n5078 ^ n27;
  assign new_n5080 = new_n5079 ^ new_n5071;
  assign new_n5081 = new_n4880 ^ new_n4868;
  assign new_n5082 = ~new_n4877 & new_n5081;
  assign new_n5083 = new_n5082 ^ new_n4880;
  assign new_n5084 = new_n5083 ^ new_n5080;
  assign new_n5085 = ~new_n1506 & n88;
  assign new_n5086 = new_n1501 & new_n2063;
  assign new_n5087 = new_n5086 ^ new_n5085;
  assign new_n5088 = n89 & new_n1500;
  assign new_n5089 = n87 & new_n1512;
  assign new_n5090 = new_n5089 ^ new_n5088;
  assign new_n5091 = new_n5090 ^ new_n5087;
  assign new_n5092 = new_n5091 ^ n24;
  assign new_n5093 = new_n5092 ^ new_n5084;
  assign new_n5094 = new_n4893 ^ new_n4881;
  assign new_n5095 = ~new_n4890 & new_n5094;
  assign new_n5096 = new_n5095 ^ new_n4893;
  assign new_n5097 = new_n5096 ^ new_n5093;
  assign new_n5098 = ~new_n1198 & n91;
  assign new_n5099 = new_n1193 & new_n2481;
  assign new_n5100 = new_n5099 ^ new_n5098;
  assign new_n5101 = n92 & new_n1192;
  assign new_n5102 = n90 & new_n1204;
  assign new_n5103 = new_n5102 ^ new_n5101;
  assign new_n5104 = new_n5103 ^ new_n5100;
  assign new_n5105 = new_n5104 ^ n21;
  assign new_n5106 = new_n5105 ^ new_n5097;
  assign new_n5107 = new_n4906 ^ new_n4894;
  assign new_n5108 = ~new_n4903 & new_n5107;
  assign new_n5109 = new_n5108 ^ new_n4906;
  assign new_n5110 = new_n5109 ^ new_n5106;
  assign new_n5111 = ~new_n930 & n94;
  assign new_n5112 = new_n925 & new_n2934;
  assign new_n5113 = new_n5112 ^ new_n5111;
  assign new_n5114 = n95 & new_n924;
  assign new_n5115 = n93 & new_n936;
  assign new_n5116 = new_n5115 ^ new_n5114;
  assign new_n5117 = new_n5116 ^ new_n5113;
  assign new_n5118 = new_n5117 ^ n18;
  assign new_n5119 = new_n5118 ^ new_n5110;
  assign new_n5120 = new_n4919 ^ new_n4907;
  assign new_n5121 = ~new_n4916 & new_n5120;
  assign new_n5122 = new_n5121 ^ new_n4919;
  assign new_n5123 = new_n5122 ^ new_n5119;
  assign new_n5124 = n97 & new_n707;
  assign new_n5125 = new_n701 & new_n3435;
  assign new_n5126 = new_n5125 ^ new_n5124;
  assign new_n5127 = n98 & new_n700;
  assign new_n5128 = n96 & new_n787;
  assign new_n5129 = new_n5128 ^ new_n5127;
  assign new_n5130 = new_n5129 ^ new_n5126;
  assign new_n5131 = new_n5130 ^ n15;
  assign new_n5132 = new_n5131 ^ new_n5123;
  assign new_n5133 = new_n4932 ^ new_n4920;
  assign new_n5134 = ~new_n4929 & new_n5133;
  assign new_n5135 = new_n5134 ^ new_n4932;
  assign new_n5136 = new_n5135 ^ new_n5132;
  assign new_n5137 = n100 & new_n499;
  assign new_n5138 = ~new_n506 & new_n3972;
  assign new_n5139 = new_n5138 ^ new_n5137;
  assign new_n5140 = ~new_n505 & n101;
  assign new_n5141 = n99 & new_n579;
  assign new_n5142 = new_n5141 ^ new_n5140;
  assign new_n5143 = new_n5142 ^ new_n5139;
  assign new_n5144 = new_n5143 ^ n12;
  assign new_n5145 = new_n5144 ^ new_n5136;
  assign new_n5146 = new_n4945 ^ new_n4933;
  assign new_n5147 = ~new_n4942 & new_n5146;
  assign new_n5148 = new_n5147 ^ new_n4945;
  assign new_n5149 = new_n5148 ^ new_n5145;
  assign new_n5150 = n103 & new_n354;
  assign new_n5151 = ~new_n4556 & new_n349;
  assign new_n5152 = new_n5151 ^ new_n5150;
  assign new_n5153 = n104 & new_n348;
  assign new_n5154 = n102 & new_n391;
  assign new_n5155 = new_n5154 ^ new_n5153;
  assign new_n5156 = new_n5155 ^ new_n5152;
  assign new_n5157 = new_n5156 ^ n9;
  assign new_n5158 = new_n5157 ^ new_n5149;
  assign new_n5159 = new_n4958 ^ new_n4946;
  assign new_n5160 = ~new_n4955 & new_n5159;
  assign new_n5161 = new_n5160 ^ new_n4958;
  assign new_n5162 = new_n5161 ^ new_n5158;
  assign new_n5163 = n106 & new_n218;
  assign new_n5164 = new_n4576 ^ n107;
  assign new_n5165 = ~new_n5164 & new_n208;
  assign new_n5166 = new_n5165 ^ new_n5163;
  assign new_n5167 = n107 & new_n207;
  assign new_n5168 = n105 & new_n212;
  assign new_n5169 = new_n5168 ^ new_n5167;
  assign new_n5170 = new_n5169 ^ new_n5166;
  assign new_n5171 = new_n5170 ^ n6;
  assign new_n5172 = new_n5171 ^ new_n5162;
  assign new_n5173 = new_n4972 ^ new_n4959;
  assign new_n5174 = ~new_n4969 & new_n5173;
  assign new_n5175 = new_n5174 ^ new_n4972;
  assign new_n5176 = new_n5175 ^ new_n5172;
  assign new_n5177 = n109 ^ n108;
  assign new_n5178 = n109 & new_n4773;
  assign new_n5179 = new_n5178 ^ new_n4772;
  assign new_n5180 = ~new_n5179 & new_n5177;
  assign new_n5181 = ~new_n5180 & new_n155;
  assign new_n5182 = new_n5181 ^ n2;
  assign new_n5183 = new_n5182 ^ n110;
  assign new_n5184 = n109 ^ n3;
  assign new_n5185 = ~n108 & ~new_n4981;
  assign new_n5186 = new_n5185 ^ new_n5184;
  assign new_n5187 = new_n5186 ^ n108;
  assign new_n5188 = ~new_n5187 & new_n241;
  assign new_n5189 = new_n5188 ^ new_n5185;
  assign new_n5190 = new_n5189 ^ n108;
  assign new_n5191 = new_n5190 ^ new_n5183;
  assign new_n5192 = ~n1 & ~new_n5191;
  assign new_n5193 = new_n5192 ^ new_n5183;
  assign new_n5194 = new_n5193 ^ new_n5176;
  assign new_n5195 = new_n4992 ^ new_n4973;
  assign new_n5196 = ~new_n4989 & new_n5195;
  assign new_n5197 = new_n5196 ^ new_n4992;
  assign new_n5198 = new_n5197 ^ new_n5194;
  assign new_n5199 = ~new_n3143 & n77;
  assign new_n5200 = ~new_n891 & new_n3138;
  assign new_n5201 = new_n5200 ^ new_n5199;
  assign new_n5202 = n78 & new_n3137;
  assign new_n5203 = n76 & new_n3149;
  assign new_n5204 = new_n5203 ^ new_n5202;
  assign new_n5205 = new_n5204 ^ new_n5201;
  assign new_n5206 = new_n5205 ^ n36;
  assign new_n5207 = new_n5044 ^ new_n5032;
  assign new_n5208 = ~new_n5041 & new_n5207;
  assign new_n5209 = new_n5208 ^ new_n5044;
  assign new_n5210 = new_n5209 ^ new_n5206;
  assign new_n5211 = ~new_n4212 & n71;
  assign new_n5212 = ~new_n459 & new_n4201;
  assign new_n5213 = new_n5212 ^ new_n5211;
  assign new_n5214 = n72 & new_n4200;
  assign new_n5215 = n70 & new_n4206;
  assign new_n5216 = new_n5215 ^ new_n5214;
  assign new_n5217 = new_n5216 ^ new_n5213;
  assign new_n5218 = new_n5217 ^ n42;
  assign new_n5219 = new_n5030 ^ new_n5018;
  assign new_n5220 = ~new_n5027 & new_n5219;
  assign new_n5221 = new_n5220 ^ new_n5030;
  assign new_n5222 = new_n5221 ^ new_n5218;
  assign new_n5223 = ~new_n5006 & ~new_n5016;
  assign new_n5224 = ~new_n5223 & new_n5014;
  assign new_n5225 = ~n45 & ~n46;
  assign new_n5226 = new_n5225 ^ new_n5015;
  assign new_n5227 = new_n5226 ^ n47;
  assign new_n5228 = ~n65 & ~new_n5227;
  assign new_n5229 = n66 ^ n46;
  assign new_n5230 = ~new_n5229 & new_n5015;
  assign new_n5231 = new_n5230 ^ n45;
  assign new_n5232 = new_n5231 ^ n47;
  assign new_n5233 = new_n5232 ^ new_n5228;
  assign new_n5234 = ~new_n4804 & n68;
  assign new_n5235 = ~new_n304 & new_n4799;
  assign new_n5236 = new_n5235 ^ new_n5234;
  assign new_n5237 = n69 & new_n4798;
  assign new_n5238 = n67 & new_n4810;
  assign new_n5239 = new_n5238 ^ new_n5237;
  assign new_n5240 = new_n5239 ^ new_n5236;
  assign new_n5241 = new_n5240 ^ n45;
  assign new_n5242 = new_n5241 ^ new_n5233;
  assign new_n5243 = new_n5242 ^ new_n5224;
  assign new_n5244 = new_n5243 ^ new_n5222;
  assign new_n5245 = ~new_n3682 & n74;
  assign new_n5246 = new_n660 & new_n3677;
  assign new_n5247 = new_n5246 ^ new_n5245;
  assign new_n5248 = n75 & new_n3676;
  assign new_n5249 = n73 & new_n3688;
  assign new_n5250 = new_n5249 ^ new_n5248;
  assign new_n5251 = new_n5250 ^ new_n5247;
  assign new_n5252 = new_n5251 ^ n39;
  assign new_n5253 = new_n5252 ^ new_n5244;
  assign new_n5254 = new_n5031 ^ new_n5001;
  assign new_n5255 = ~new_n5254 & new_n5005;
  assign new_n5256 = new_n5255 ^ new_n5004;
  assign new_n5257 = new_n5256 ^ new_n5253;
  assign new_n5258 = new_n5257 ^ new_n5210;
  assign new_n5259 = ~new_n2672 & n80;
  assign new_n5260 = new_n1161 & new_n2667;
  assign new_n5261 = new_n5260 ^ new_n5259;
  assign new_n5262 = n81 & new_n2666;
  assign new_n5263 = n79 & new_n2664;
  assign new_n5264 = new_n5263 ^ new_n5262;
  assign new_n5265 = new_n5264 ^ new_n5261;
  assign new_n5266 = new_n5265 ^ n33;
  assign new_n5267 = new_n5266 ^ new_n5258;
  assign new_n5268 = new_n5057 ^ new_n5045;
  assign new_n5269 = ~new_n5054 & new_n5268;
  assign new_n5270 = new_n5269 ^ new_n5057;
  assign new_n5271 = new_n5270 ^ new_n5267;
  assign new_n5272 = n83 & new_n2246;
  assign new_n5273 = new_n1468 & new_n2241;
  assign new_n5274 = new_n5273 ^ new_n5272;
  assign new_n5275 = n84 & new_n2240;
  assign new_n5276 = n82 & new_n2391;
  assign new_n5277 = new_n5276 ^ new_n5275;
  assign new_n5278 = new_n5277 ^ new_n5274;
  assign new_n5279 = new_n5278 ^ n30;
  assign new_n5280 = new_n5279 ^ new_n5271;
  assign new_n5281 = new_n5070 ^ new_n5058;
  assign new_n5282 = ~new_n5067 & new_n5281;
  assign new_n5283 = new_n5282 ^ new_n5070;
  assign new_n5284 = new_n5283 ^ new_n5280;
  assign new_n5285 = n86 & new_n1874;
  assign new_n5286 = new_n1811 & new_n1864;
  assign new_n5287 = new_n5286 ^ new_n5285;
  assign new_n5288 = n87 & new_n1863;
  assign new_n5289 = n85 & new_n1868;
  assign new_n5290 = new_n5289 ^ new_n5288;
  assign new_n5291 = new_n5290 ^ new_n5287;
  assign new_n5292 = new_n5291 ^ n27;
  assign new_n5293 = new_n5292 ^ new_n5284;
  assign new_n5294 = new_n5083 ^ new_n5071;
  assign new_n5295 = ~new_n5080 & new_n5294;
  assign new_n5296 = new_n5295 ^ new_n5083;
  assign new_n5297 = new_n5296 ^ new_n5293;
  assign new_n5298 = ~new_n1506 & n89;
  assign new_n5299 = new_n1501 & new_n2193;
  assign new_n5300 = new_n5299 ^ new_n5298;
  assign new_n5301 = n90 & new_n1500;
  assign new_n5302 = n88 & new_n1512;
  assign new_n5303 = new_n5302 ^ new_n5301;
  assign new_n5304 = new_n5303 ^ new_n5300;
  assign new_n5305 = new_n5304 ^ n24;
  assign new_n5306 = new_n5305 ^ new_n5297;
  assign new_n5307 = new_n5096 ^ new_n5084;
  assign new_n5308 = ~new_n5093 & new_n5307;
  assign new_n5309 = new_n5308 ^ new_n5096;
  assign new_n5310 = new_n5309 ^ new_n5306;
  assign new_n5311 = ~new_n1198 & n92;
  assign new_n5312 = new_n1193 & new_n2628;
  assign new_n5313 = new_n5312 ^ new_n5311;
  assign new_n5314 = n93 & new_n1192;
  assign new_n5315 = n91 & new_n1204;
  assign new_n5316 = new_n5315 ^ new_n5314;
  assign new_n5317 = new_n5316 ^ new_n5313;
  assign new_n5318 = new_n5317 ^ n21;
  assign new_n5319 = new_n5318 ^ new_n5310;
  assign new_n5320 = new_n5109 ^ new_n5097;
  assign new_n5321 = ~new_n5106 & new_n5320;
  assign new_n5322 = new_n5321 ^ new_n5109;
  assign new_n5323 = new_n5322 ^ new_n5319;
  assign new_n5324 = ~new_n930 & n95;
  assign new_n5325 = new_n925 & new_n3095;
  assign new_n5326 = new_n5325 ^ new_n5324;
  assign new_n5327 = n96 & new_n924;
  assign new_n5328 = n94 & new_n936;
  assign new_n5329 = new_n5328 ^ new_n5327;
  assign new_n5330 = new_n5329 ^ new_n5326;
  assign new_n5331 = new_n5330 ^ n18;
  assign new_n5332 = new_n5331 ^ new_n5323;
  assign new_n5333 = new_n5122 ^ new_n5110;
  assign new_n5334 = ~new_n5119 & new_n5333;
  assign new_n5335 = new_n5334 ^ new_n5122;
  assign new_n5336 = new_n5335 ^ new_n5332;
  assign new_n5337 = n98 & new_n707;
  assign new_n5338 = new_n701 & new_n3604;
  assign new_n5339 = new_n5338 ^ new_n5337;
  assign new_n5340 = n99 & new_n700;
  assign new_n5341 = n97 & new_n787;
  assign new_n5342 = new_n5341 ^ new_n5340;
  assign new_n5343 = new_n5342 ^ new_n5339;
  assign new_n5344 = new_n5343 ^ n15;
  assign new_n5345 = new_n5344 ^ new_n5336;
  assign new_n5346 = new_n5135 ^ new_n5123;
  assign new_n5347 = ~new_n5132 & new_n5346;
  assign new_n5348 = new_n5347 ^ new_n5135;
  assign new_n5349 = new_n5348 ^ new_n5345;
  assign new_n5350 = n101 & new_n499;
  assign new_n5351 = ~new_n506 & new_n4159;
  assign new_n5352 = new_n5351 ^ new_n5350;
  assign new_n5353 = ~new_n505 & n102;
  assign new_n5354 = n100 & new_n579;
  assign new_n5355 = new_n5354 ^ new_n5353;
  assign new_n5356 = new_n5355 ^ new_n5352;
  assign new_n5357 = new_n5356 ^ n12;
  assign new_n5358 = new_n5357 ^ new_n5349;
  assign new_n5359 = new_n5148 ^ new_n5136;
  assign new_n5360 = ~new_n5145 & new_n5359;
  assign new_n5361 = new_n5360 ^ new_n5148;
  assign new_n5362 = new_n5361 ^ new_n5358;
  assign new_n5363 = n104 & new_n354;
  assign new_n5364 = ~new_n4754 & new_n349;
  assign new_n5365 = new_n5364 ^ new_n5363;
  assign new_n5366 = n105 & new_n348;
  assign new_n5367 = n103 & new_n391;
  assign new_n5368 = new_n5367 ^ new_n5366;
  assign new_n5369 = new_n5368 ^ new_n5365;
  assign new_n5370 = new_n5369 ^ n9;
  assign new_n5371 = new_n5370 ^ new_n5362;
  assign new_n5372 = new_n5161 ^ new_n5149;
  assign new_n5373 = ~new_n5158 & new_n5372;
  assign new_n5374 = new_n5373 ^ new_n5161;
  assign new_n5375 = new_n5374 ^ new_n5371;
  assign new_n5376 = n107 & new_n218;
  assign new_n5377 = new_n4773 ^ n108;
  assign new_n5378 = ~new_n5377 & new_n208;
  assign new_n5379 = new_n5378 ^ new_n5376;
  assign new_n5380 = n108 & new_n207;
  assign new_n5381 = n106 & new_n212;
  assign new_n5382 = new_n5381 ^ new_n5380;
  assign new_n5383 = new_n5382 ^ new_n5379;
  assign new_n5384 = new_n5383 ^ n6;
  assign new_n5385 = new_n5384 ^ new_n5375;
  assign new_n5386 = new_n5175 ^ new_n5162;
  assign new_n5387 = ~new_n5172 & new_n5386;
  assign new_n5388 = new_n5387 ^ new_n5175;
  assign new_n5389 = new_n5388 ^ new_n5385;
  assign new_n5390 = n110 ^ n109;
  assign new_n5391 = new_n5180 & new_n5390;
  assign new_n5392 = new_n5391 ^ n109;
  assign new_n5393 = new_n5392 ^ n110;
  assign new_n5394 = ~new_n5393 & new_n155;
  assign new_n5395 = new_n5394 ^ n2;
  assign new_n5396 = new_n5395 ^ n111;
  assign new_n5397 = n110 ^ n3;
  assign new_n5398 = ~n109 & ~new_n5184;
  assign new_n5399 = new_n5398 ^ new_n5397;
  assign new_n5400 = new_n5399 ^ n109;
  assign new_n5401 = ~new_n5400 & new_n241;
  assign new_n5402 = new_n5401 ^ new_n5398;
  assign new_n5403 = new_n5402 ^ n109;
  assign new_n5404 = new_n5403 ^ new_n5396;
  assign new_n5405 = ~n1 & ~new_n5404;
  assign new_n5406 = new_n5405 ^ new_n5396;
  assign new_n5407 = new_n5406 ^ new_n5389;
  assign new_n5408 = new_n5197 ^ new_n5176;
  assign new_n5409 = ~new_n5194 & new_n5408;
  assign new_n5410 = new_n5409 ^ new_n5197;
  assign new_n5411 = new_n5410 ^ new_n5407;
  assign new_n5412 = new_n5241 ^ new_n5224;
  assign new_n5413 = ~new_n5242 & new_n5412;
  assign new_n5414 = new_n5413 ^ new_n5224;
  assign new_n5415 = ~new_n5226 & n47;
  assign new_n5416 = n65 & new_n5415;
  assign new_n5417 = n48 ^ n47;
  assign new_n5418 = ~new_n5417 & new_n5015;
  assign new_n5419 = new_n5418 ^ new_n5015;
  assign new_n5420 = ~new_n151 & new_n5419;
  assign new_n5421 = n67 & new_n5015;
  assign new_n5422 = new_n5421 ^ new_n5420;
  assign new_n5423 = ~new_n5015 & n47;
  assign new_n5424 = new_n5423 ^ new_n5226;
  assign new_n5425 = ~new_n5424 & n66;
  assign new_n5426 = new_n5425 ^ new_n5422;
  assign new_n5427 = new_n5426 ^ new_n5416;
  assign new_n5428 = n48 & new_n5225;
  assign new_n5429 = ~n47 & new_n5428;
  assign new_n5430 = n65 & new_n5429;
  assign new_n5431 = new_n5430 ^ new_n5426;
  assign new_n5432 = ~new_n5016 & ~new_n5233;
  assign new_n5433 = new_n5432 ^ new_n5431;
  assign new_n5434 = new_n5433 ^ new_n5427;
  assign new_n5435 = ~n48 & ~new_n5434;
  assign new_n5436 = new_n5435 ^ new_n5433;
  assign new_n5437 = new_n5436 ^ new_n5414;
  assign new_n5438 = ~new_n4804 & n69;
  assign new_n5439 = ~new_n339 & new_n4799;
  assign new_n5440 = new_n5439 ^ new_n5438;
  assign new_n5441 = n70 & new_n4798;
  assign new_n5442 = n68 & new_n4810;
  assign new_n5443 = new_n5442 ^ new_n5441;
  assign new_n5444 = new_n5443 ^ new_n5440;
  assign new_n5445 = new_n5444 ^ n45;
  assign new_n5446 = new_n5445 ^ new_n5437;
  assign new_n5447 = new_n5243 ^ new_n5218;
  assign new_n5448 = ~new_n5447 & new_n5222;
  assign new_n5449 = new_n5448 ^ new_n5221;
  assign new_n5450 = new_n5449 ^ new_n5446;
  assign new_n5451 = ~new_n4212 & n72;
  assign new_n5452 = new_n534 & new_n4201;
  assign new_n5453 = new_n5452 ^ new_n5451;
  assign new_n5454 = n73 & new_n4200;
  assign new_n5455 = n71 & new_n4206;
  assign new_n5456 = new_n5455 ^ new_n5454;
  assign new_n5457 = new_n5456 ^ new_n5453;
  assign new_n5458 = new_n5457 ^ n42;
  assign new_n5459 = new_n5458 ^ new_n5450;
  assign new_n5460 = new_n5256 ^ new_n5244;
  assign new_n5461 = ~new_n5253 & new_n5460;
  assign new_n5462 = new_n5461 ^ new_n5256;
  assign new_n5463 = new_n5462 ^ new_n5459;
  assign new_n5464 = ~new_n3682 & n75;
  assign new_n5465 = ~new_n737 & new_n3677;
  assign new_n5466 = new_n5465 ^ new_n5464;
  assign new_n5467 = n74 & new_n3688;
  assign new_n5468 = n76 & new_n3676;
  assign new_n5469 = new_n5468 ^ new_n5467;
  assign new_n5470 = new_n5469 ^ new_n5466;
  assign new_n5471 = new_n5470 ^ n39;
  assign new_n5472 = new_n5471 ^ new_n5463;
  assign new_n5473 = ~new_n3143 & n78;
  assign new_n5474 = ~new_n982 & new_n3138;
  assign new_n5475 = new_n5474 ^ new_n5473;
  assign new_n5476 = n79 & new_n3137;
  assign new_n5477 = n77 & new_n3149;
  assign new_n5478 = new_n5477 ^ new_n5476;
  assign new_n5479 = new_n5478 ^ new_n5475;
  assign new_n5480 = new_n5479 ^ n36;
  assign new_n5481 = new_n5480 ^ new_n5472;
  assign new_n5482 = new_n5257 ^ new_n5206;
  assign new_n5483 = ~new_n5482 & new_n5210;
  assign new_n5484 = new_n5483 ^ new_n5209;
  assign new_n5485 = new_n5484 ^ new_n5481;
  assign new_n5486 = ~new_n2672 & n81;
  assign new_n5487 = new_n1263 & new_n2667;
  assign new_n5488 = new_n5487 ^ new_n5486;
  assign new_n5489 = n82 & new_n2666;
  assign new_n5490 = n80 & new_n2664;
  assign new_n5491 = new_n5490 ^ new_n5489;
  assign new_n5492 = new_n5491 ^ new_n5488;
  assign new_n5493 = new_n5492 ^ n33;
  assign new_n5494 = new_n5493 ^ new_n5485;
  assign new_n5495 = new_n5270 ^ new_n5258;
  assign new_n5496 = ~new_n5267 & new_n5495;
  assign new_n5497 = new_n5496 ^ new_n5270;
  assign new_n5498 = new_n5497 ^ new_n5494;
  assign new_n5499 = n84 & new_n2246;
  assign new_n5500 = new_n1584 & new_n2241;
  assign new_n5501 = new_n5500 ^ new_n5499;
  assign new_n5502 = n85 & new_n2240;
  assign new_n5503 = n83 & new_n2391;
  assign new_n5504 = new_n5503 ^ new_n5502;
  assign new_n5505 = new_n5504 ^ new_n5501;
  assign new_n5506 = new_n5505 ^ n30;
  assign new_n5507 = new_n5506 ^ new_n5498;
  assign new_n5508 = new_n5283 ^ new_n5271;
  assign new_n5509 = ~new_n5280 & new_n5508;
  assign new_n5510 = new_n5509 ^ new_n5283;
  assign new_n5511 = new_n5510 ^ new_n5507;
  assign new_n5512 = n87 & new_n1874;
  assign new_n5513 = new_n1864 & new_n1940;
  assign new_n5514 = new_n5513 ^ new_n5512;
  assign new_n5515 = n88 & new_n1863;
  assign new_n5516 = n86 & new_n1868;
  assign new_n5517 = new_n5516 ^ new_n5515;
  assign new_n5518 = new_n5517 ^ new_n5514;
  assign new_n5519 = new_n5518 ^ n27;
  assign new_n5520 = new_n5519 ^ new_n5511;
  assign new_n5521 = new_n5296 ^ new_n5284;
  assign new_n5522 = ~new_n5293 & new_n5521;
  assign new_n5523 = new_n5522 ^ new_n5296;
  assign new_n5524 = new_n5523 ^ new_n5520;
  assign new_n5525 = ~new_n1506 & n90;
  assign new_n5526 = new_n1501 & new_n2341;
  assign new_n5527 = new_n5526 ^ new_n5525;
  assign new_n5528 = n91 & new_n1500;
  assign new_n5529 = n89 & new_n1512;
  assign new_n5530 = new_n5529 ^ new_n5528;
  assign new_n5531 = new_n5530 ^ new_n5527;
  assign new_n5532 = new_n5531 ^ n24;
  assign new_n5533 = new_n5532 ^ new_n5524;
  assign new_n5534 = new_n5309 ^ new_n5297;
  assign new_n5535 = ~new_n5306 & new_n5534;
  assign new_n5536 = new_n5535 ^ new_n5309;
  assign new_n5537 = new_n5536 ^ new_n5533;
  assign new_n5538 = ~new_n1198 & n93;
  assign new_n5539 = new_n1193 & new_n2785;
  assign new_n5540 = new_n5539 ^ new_n5538;
  assign new_n5541 = n94 & new_n1192;
  assign new_n5542 = n92 & new_n1204;
  assign new_n5543 = new_n5542 ^ new_n5541;
  assign new_n5544 = new_n5543 ^ new_n5540;
  assign new_n5545 = new_n5544 ^ n21;
  assign new_n5546 = new_n5545 ^ new_n5537;
  assign new_n5547 = new_n5322 ^ new_n5310;
  assign new_n5548 = ~new_n5319 & new_n5547;
  assign new_n5549 = new_n5548 ^ new_n5322;
  assign new_n5550 = new_n5549 ^ new_n5546;
  assign new_n5551 = ~new_n930 & n96;
  assign new_n5552 = new_n925 & new_n3273;
  assign new_n5553 = new_n5552 ^ new_n5551;
  assign new_n5554 = n97 & new_n924;
  assign new_n5555 = n95 & new_n936;
  assign new_n5556 = new_n5555 ^ new_n5554;
  assign new_n5557 = new_n5556 ^ new_n5553;
  assign new_n5558 = new_n5557 ^ n18;
  assign new_n5559 = new_n5558 ^ new_n5550;
  assign new_n5560 = new_n5335 ^ new_n5323;
  assign new_n5561 = ~new_n5332 & new_n5560;
  assign new_n5562 = new_n5561 ^ new_n5335;
  assign new_n5563 = new_n5562 ^ new_n5559;
  assign new_n5564 = n99 & new_n707;
  assign new_n5565 = new_n701 & new_n3789;
  assign new_n5566 = new_n5565 ^ new_n5564;
  assign new_n5567 = n100 & new_n700;
  assign new_n5568 = n98 & new_n787;
  assign new_n5569 = new_n5568 ^ new_n5567;
  assign new_n5570 = new_n5569 ^ new_n5566;
  assign new_n5571 = new_n5570 ^ n15;
  assign new_n5572 = new_n5571 ^ new_n5563;
  assign new_n5573 = new_n5348 ^ new_n5336;
  assign new_n5574 = ~new_n5345 & new_n5573;
  assign new_n5575 = new_n5574 ^ new_n5348;
  assign new_n5576 = new_n5575 ^ new_n5572;
  assign new_n5577 = n102 & new_n499;
  assign new_n5578 = ~new_n506 & new_n4368;
  assign new_n5579 = new_n5578 ^ new_n5577;
  assign new_n5580 = ~new_n505 & n103;
  assign new_n5581 = n101 & new_n579;
  assign new_n5582 = new_n5581 ^ new_n5580;
  assign new_n5583 = new_n5582 ^ new_n5579;
  assign new_n5584 = new_n5583 ^ n12;
  assign new_n5585 = new_n5584 ^ new_n5576;
  assign new_n5586 = new_n5361 ^ new_n5349;
  assign new_n5587 = ~new_n5358 & new_n5586;
  assign new_n5588 = new_n5587 ^ new_n5361;
  assign new_n5589 = new_n5588 ^ new_n5585;
  assign new_n5590 = n105 & new_n354;
  assign new_n5591 = ~new_n4961 & new_n349;
  assign new_n5592 = new_n5591 ^ new_n5590;
  assign new_n5593 = n106 & new_n348;
  assign new_n5594 = n104 & new_n391;
  assign new_n5595 = new_n5594 ^ new_n5593;
  assign new_n5596 = new_n5595 ^ new_n5592;
  assign new_n5597 = new_n5596 ^ n9;
  assign new_n5598 = new_n5597 ^ new_n5589;
  assign new_n5599 = new_n5374 ^ new_n5362;
  assign new_n5600 = ~new_n5371 & new_n5599;
  assign new_n5601 = new_n5600 ^ new_n5374;
  assign new_n5602 = new_n5601 ^ new_n5598;
  assign new_n5603 = n108 & new_n218;
  assign new_n5604 = new_n4977 ^ n109;
  assign new_n5605 = new_n208 & new_n5604;
  assign new_n5606 = new_n5605 ^ new_n5603;
  assign new_n5607 = n109 & new_n207;
  assign new_n5608 = n107 & new_n212;
  assign new_n5609 = new_n5608 ^ new_n5607;
  assign new_n5610 = new_n5609 ^ new_n5606;
  assign new_n5611 = new_n5610 ^ n6;
  assign new_n5612 = new_n5611 ^ new_n5602;
  assign new_n5613 = new_n5388 ^ new_n5375;
  assign new_n5614 = ~new_n5385 & new_n5613;
  assign new_n5615 = new_n5614 ^ new_n5388;
  assign new_n5616 = new_n5615 ^ new_n5612;
  assign new_n5617 = n110 & new_n5392;
  assign new_n5618 = new_n5617 ^ new_n5393;
  assign new_n5619 = n111 & new_n5618;
  assign new_n5620 = ~n111 & ~new_n5617;
  assign new_n5621 = new_n5620 ^ new_n5619;
  assign new_n5622 = new_n155 & new_n5621;
  assign new_n5623 = new_n5622 ^ n2;
  assign new_n5624 = new_n5623 ^ n112;
  assign new_n5625 = n111 ^ n3;
  assign new_n5626 = ~n110 & n3;
  assign new_n5627 = new_n5626 ^ new_n5625;
  assign new_n5628 = ~n2 & new_n5627;
  assign new_n5629 = new_n5628 ^ new_n5625;
  assign new_n5630 = new_n5629 ^ new_n5624;
  assign new_n5631 = ~n1 & new_n5630;
  assign new_n5632 = new_n5631 ^ new_n5624;
  assign new_n5633 = new_n5632 ^ new_n5616;
  assign new_n5634 = new_n5410 ^ new_n5389;
  assign new_n5635 = ~new_n5407 & new_n5634;
  assign new_n5636 = new_n5635 ^ new_n5410;
  assign new_n5637 = new_n5636 ^ new_n5633;
  assign new_n5638 = ~new_n5431 & new_n5432;
  assign new_n5639 = n48 & new_n5638;
  assign new_n5640 = n49 ^ n48;
  assign new_n5641 = n65 & new_n5640;
  assign new_n5642 = new_n5641 ^ new_n5639;
  assign new_n5643 = ~new_n154 & new_n5417;
  assign new_n5644 = new_n5643 ^ n68;
  assign new_n5645 = new_n5015 & new_n5644;
  assign new_n5646 = ~new_n5015 & n48;
  assign new_n5647 = new_n5646 ^ new_n5226;
  assign new_n5648 = ~new_n5647 & new_n5417;
  assign new_n5649 = n66 & new_n5648;
  assign new_n5650 = ~new_n5424 & n67;
  assign new_n5651 = new_n5650 ^ new_n5649;
  assign new_n5652 = ~new_n5645 & ~new_n5651;
  assign new_n5653 = new_n5652 ^ n48;
  assign new_n5654 = new_n5653 ^ new_n5642;
  assign new_n5655 = ~new_n4804 & n70;
  assign new_n5656 = ~new_n402 & new_n4799;
  assign new_n5657 = new_n5656 ^ new_n5655;
  assign new_n5658 = n71 & new_n4798;
  assign new_n5659 = n69 & new_n4810;
  assign new_n5660 = new_n5659 ^ new_n5658;
  assign new_n5661 = new_n5660 ^ new_n5657;
  assign new_n5662 = new_n5661 ^ n45;
  assign new_n5663 = new_n5662 ^ new_n5654;
  assign new_n5664 = new_n5445 ^ new_n5436;
  assign new_n5665 = ~new_n5437 & new_n5664;
  assign new_n5666 = new_n5665 ^ new_n5414;
  assign new_n5667 = new_n5666 ^ new_n5663;
  assign new_n5668 = new_n5458 ^ new_n5446;
  assign new_n5669 = ~new_n5450 & new_n5668;
  assign new_n5670 = new_n5669 ^ new_n5449;
  assign new_n5671 = new_n5670 ^ new_n5667;
  assign new_n5672 = ~new_n4212 & n73;
  assign new_n5673 = new_n595 & new_n4201;
  assign new_n5674 = new_n5673 ^ new_n5672;
  assign new_n5675 = n74 & new_n4200;
  assign new_n5676 = n72 & new_n4206;
  assign new_n5677 = new_n5676 ^ new_n5675;
  assign new_n5678 = new_n5677 ^ new_n5674;
  assign new_n5679 = new_n5678 ^ n42;
  assign new_n5680 = new_n5679 ^ new_n5671;
  assign new_n5681 = ~new_n3682 & n76;
  assign new_n5682 = ~new_n812 & new_n3677;
  assign new_n5683 = new_n5682 ^ new_n5681;
  assign new_n5684 = n77 & new_n3676;
  assign new_n5685 = n75 & new_n3688;
  assign new_n5686 = new_n5685 ^ new_n5684;
  assign new_n5687 = new_n5686 ^ new_n5683;
  assign new_n5688 = new_n5687 ^ n39;
  assign new_n5689 = new_n5688 ^ new_n5680;
  assign new_n5690 = new_n5471 ^ new_n5459;
  assign new_n5691 = ~new_n5463 & new_n5690;
  assign new_n5692 = new_n5691 ^ new_n5462;
  assign new_n5693 = new_n5692 ^ new_n5689;
  assign new_n5694 = new_n5484 ^ new_n5472;
  assign new_n5695 = ~new_n5694 & new_n5481;
  assign new_n5696 = new_n5695 ^ new_n5484;
  assign new_n5697 = new_n5696 ^ new_n5693;
  assign new_n5698 = ~new_n3143 & n79;
  assign new_n5699 = new_n1069 & new_n3138;
  assign new_n5700 = new_n5699 ^ new_n5698;
  assign new_n5701 = n80 & new_n3137;
  assign new_n5702 = n78 & new_n3149;
  assign new_n5703 = new_n5702 ^ new_n5701;
  assign new_n5704 = new_n5703 ^ new_n5700;
  assign new_n5705 = new_n5704 ^ n36;
  assign new_n5706 = new_n5705 ^ new_n5697;
  assign new_n5707 = ~new_n2672 & n82;
  assign new_n5708 = new_n1363 & new_n2667;
  assign new_n5709 = new_n5708 ^ new_n5707;
  assign new_n5710 = n83 & new_n2666;
  assign new_n5711 = n81 & new_n2664;
  assign new_n5712 = new_n5711 ^ new_n5710;
  assign new_n5713 = new_n5712 ^ new_n5709;
  assign new_n5714 = new_n5713 ^ n33;
  assign new_n5715 = new_n5714 ^ new_n5706;
  assign new_n5716 = new_n5497 ^ new_n5485;
  assign new_n5717 = ~new_n5716 & new_n5494;
  assign new_n5718 = new_n5717 ^ new_n5497;
  assign new_n5719 = new_n5718 ^ new_n5715;
  assign new_n5720 = n85 & new_n2246;
  assign new_n5721 = new_n1694 & new_n2241;
  assign new_n5722 = new_n5721 ^ new_n5720;
  assign new_n5723 = n86 & new_n2240;
  assign new_n5724 = n84 & new_n2391;
  assign new_n5725 = new_n5724 ^ new_n5723;
  assign new_n5726 = new_n5725 ^ new_n5722;
  assign new_n5727 = new_n5726 ^ n30;
  assign new_n5728 = new_n5727 ^ new_n5719;
  assign new_n5729 = new_n5510 ^ new_n5498;
  assign new_n5730 = ~new_n5729 & new_n5507;
  assign new_n5731 = new_n5730 ^ new_n5510;
  assign new_n5732 = new_n5731 ^ new_n5728;
  assign new_n5733 = n88 & new_n1874;
  assign new_n5734 = new_n1864 & new_n2063;
  assign new_n5735 = new_n5734 ^ new_n5733;
  assign new_n5736 = n89 & new_n1863;
  assign new_n5737 = n87 & new_n1868;
  assign new_n5738 = new_n5737 ^ new_n5736;
  assign new_n5739 = new_n5738 ^ new_n5735;
  assign new_n5740 = new_n5739 ^ n27;
  assign new_n5741 = new_n5740 ^ new_n5732;
  assign new_n5742 = new_n5523 ^ new_n5511;
  assign new_n5743 = ~new_n5742 & new_n5520;
  assign new_n5744 = new_n5743 ^ new_n5523;
  assign new_n5745 = new_n5744 ^ new_n5741;
  assign new_n5746 = ~new_n1506 & n91;
  assign new_n5747 = new_n1501 & new_n2481;
  assign new_n5748 = new_n5747 ^ new_n5746;
  assign new_n5749 = n92 & new_n1500;
  assign new_n5750 = n90 & new_n1512;
  assign new_n5751 = new_n5750 ^ new_n5749;
  assign new_n5752 = new_n5751 ^ new_n5748;
  assign new_n5753 = new_n5752 ^ n24;
  assign new_n5754 = new_n5753 ^ new_n5745;
  assign new_n5755 = new_n5536 ^ new_n5524;
  assign new_n5756 = ~new_n5755 & new_n5533;
  assign new_n5757 = new_n5756 ^ new_n5536;
  assign new_n5758 = new_n5757 ^ new_n5754;
  assign new_n5759 = ~new_n1198 & n94;
  assign new_n5760 = new_n1193 & new_n2934;
  assign new_n5761 = new_n5760 ^ new_n5759;
  assign new_n5762 = n95 & new_n1192;
  assign new_n5763 = n93 & new_n1204;
  assign new_n5764 = new_n5763 ^ new_n5762;
  assign new_n5765 = new_n5764 ^ new_n5761;
  assign new_n5766 = new_n5765 ^ n21;
  assign new_n5767 = new_n5766 ^ new_n5758;
  assign new_n5768 = new_n5549 ^ new_n5537;
  assign new_n5769 = ~new_n5768 & new_n5546;
  assign new_n5770 = new_n5769 ^ new_n5549;
  assign new_n5771 = new_n5770 ^ new_n5767;
  assign new_n5772 = ~new_n930 & n97;
  assign new_n5773 = new_n925 & new_n3435;
  assign new_n5774 = new_n5773 ^ new_n5772;
  assign new_n5775 = n98 & new_n924;
  assign new_n5776 = n96 & new_n936;
  assign new_n5777 = new_n5776 ^ new_n5775;
  assign new_n5778 = new_n5777 ^ new_n5774;
  assign new_n5779 = new_n5778 ^ n18;
  assign new_n5780 = new_n5779 ^ new_n5771;
  assign new_n5781 = new_n5562 ^ new_n5550;
  assign new_n5782 = ~new_n5781 & new_n5559;
  assign new_n5783 = new_n5782 ^ new_n5562;
  assign new_n5784 = new_n5783 ^ new_n5780;
  assign new_n5785 = n100 & new_n707;
  assign new_n5786 = new_n701 & new_n3972;
  assign new_n5787 = new_n5786 ^ new_n5785;
  assign new_n5788 = n101 & new_n700;
  assign new_n5789 = n99 & new_n787;
  assign new_n5790 = new_n5789 ^ new_n5788;
  assign new_n5791 = new_n5790 ^ new_n5787;
  assign new_n5792 = new_n5791 ^ n15;
  assign new_n5793 = new_n5792 ^ new_n5784;
  assign new_n5794 = new_n5575 ^ new_n5563;
  assign new_n5795 = ~new_n5794 & new_n5572;
  assign new_n5796 = new_n5795 ^ new_n5575;
  assign new_n5797 = new_n5796 ^ new_n5793;
  assign new_n5798 = n103 & new_n499;
  assign new_n5799 = ~new_n506 & ~new_n4556;
  assign new_n5800 = new_n5799 ^ new_n5798;
  assign new_n5801 = ~new_n505 & n104;
  assign new_n5802 = n102 & new_n579;
  assign new_n5803 = new_n5802 ^ new_n5801;
  assign new_n5804 = new_n5803 ^ new_n5800;
  assign new_n5805 = new_n5804 ^ n12;
  assign new_n5806 = new_n5805 ^ new_n5797;
  assign new_n5807 = new_n5588 ^ new_n5576;
  assign new_n5808 = ~new_n5807 & new_n5585;
  assign new_n5809 = new_n5808 ^ new_n5588;
  assign new_n5810 = new_n5809 ^ new_n5806;
  assign new_n5811 = n106 & new_n354;
  assign new_n5812 = ~new_n5164 & new_n349;
  assign new_n5813 = new_n5812 ^ new_n5811;
  assign new_n5814 = n107 & new_n348;
  assign new_n5815 = n105 & new_n391;
  assign new_n5816 = new_n5815 ^ new_n5814;
  assign new_n5817 = new_n5816 ^ new_n5813;
  assign new_n5818 = new_n5817 ^ n9;
  assign new_n5819 = new_n5818 ^ new_n5810;
  assign new_n5820 = new_n5601 ^ new_n5589;
  assign new_n5821 = ~new_n5820 & new_n5598;
  assign new_n5822 = new_n5821 ^ new_n5601;
  assign new_n5823 = new_n5822 ^ new_n5819;
  assign new_n5824 = n109 & new_n218;
  assign new_n5825 = new_n5180 ^ n110;
  assign new_n5826 = new_n208 & new_n5825;
  assign new_n5827 = new_n5826 ^ new_n5824;
  assign new_n5828 = n110 & new_n207;
  assign new_n5829 = n108 & new_n212;
  assign new_n5830 = new_n5829 ^ new_n5828;
  assign new_n5831 = new_n5830 ^ new_n5827;
  assign new_n5832 = new_n5831 ^ n6;
  assign new_n5833 = new_n5832 ^ new_n5823;
  assign new_n5834 = new_n5615 ^ new_n5602;
  assign new_n5835 = ~new_n5834 & new_n5612;
  assign new_n5836 = new_n5835 ^ new_n5615;
  assign new_n5837 = new_n5836 ^ new_n5833;
  assign new_n5838 = n112 ^ n3;
  assign new_n5839 = ~n111 & n3;
  assign new_n5840 = new_n5839 ^ new_n5838;
  assign new_n5841 = ~n2 & new_n5840;
  assign new_n5842 = new_n5841 ^ new_n5838;
  assign new_n5843 = ~new_n5620 & n112;
  assign new_n5844 = ~n112 & ~new_n5619;
  assign new_n5845 = new_n5844 ^ new_n5843;
  assign new_n5846 = new_n155 & new_n5845;
  assign new_n5847 = new_n5846 ^ n2;
  assign new_n5848 = new_n5847 ^ n113;
  assign new_n5849 = new_n5848 ^ new_n5842;
  assign new_n5850 = ~n1 & new_n5849;
  assign new_n5851 = new_n5850 ^ new_n5848;
  assign new_n5852 = new_n5851 ^ new_n5837;
  assign new_n5853 = new_n5636 ^ new_n5616;
  assign new_n5854 = ~new_n5853 & new_n5633;
  assign new_n5855 = new_n5854 ^ new_n5636;
  assign new_n5856 = new_n5855 ^ new_n5852;
  assign new_n5857 = ~new_n5639 & ~new_n5641;
  assign new_n5858 = ~new_n5653 & ~new_n5857;
  assign new_n5859 = n66 ^ n49;
  assign new_n5860 = ~new_n5859 & new_n5640;
  assign new_n5861 = new_n5860 ^ n48;
  assign new_n5862 = new_n5861 ^ n50;
  assign new_n5863 = ~n48 & ~n49;
  assign new_n5864 = new_n5863 ^ new_n5640;
  assign new_n5865 = new_n5864 ^ n50;
  assign new_n5866 = ~n65 & ~new_n5865;
  assign new_n5867 = new_n5866 ^ new_n5862;
  assign new_n5868 = new_n5867 ^ new_n5858;
  assign new_n5869 = ~new_n5424 & n68;
  assign new_n5870 = ~new_n304 & new_n5419;
  assign new_n5871 = new_n5870 ^ new_n5869;
  assign new_n5872 = n69 & new_n5418;
  assign new_n5873 = n67 & new_n5648;
  assign new_n5874 = new_n5873 ^ new_n5872;
  assign new_n5875 = new_n5874 ^ new_n5871;
  assign new_n5876 = new_n5875 ^ n48;
  assign new_n5877 = new_n5876 ^ new_n5868;
  assign new_n5878 = ~new_n4804 & n71;
  assign new_n5879 = ~new_n459 & new_n4799;
  assign new_n5880 = new_n5879 ^ new_n5878;
  assign new_n5881 = n72 & new_n4798;
  assign new_n5882 = n70 & new_n4810;
  assign new_n5883 = new_n5882 ^ new_n5881;
  assign new_n5884 = new_n5883 ^ new_n5880;
  assign new_n5885 = new_n5884 ^ n45;
  assign new_n5886 = new_n5885 ^ new_n5877;
  assign new_n5887 = new_n5666 ^ new_n5654;
  assign new_n5888 = ~new_n5887 & new_n5663;
  assign new_n5889 = new_n5888 ^ new_n5666;
  assign new_n5890 = new_n5889 ^ new_n5886;
  assign new_n5891 = ~new_n4212 & n74;
  assign new_n5892 = new_n660 & new_n4201;
  assign new_n5893 = new_n5892 ^ new_n5891;
  assign new_n5894 = n75 & new_n4200;
  assign new_n5895 = n73 & new_n4206;
  assign new_n5896 = new_n5895 ^ new_n5894;
  assign new_n5897 = new_n5896 ^ new_n5893;
  assign new_n5898 = new_n5897 ^ n42;
  assign new_n5899 = new_n5898 ^ new_n5890;
  assign new_n5900 = new_n5679 ^ new_n5667;
  assign new_n5901 = ~new_n5671 & new_n5900;
  assign new_n5902 = new_n5901 ^ new_n5670;
  assign new_n5903 = new_n5902 ^ new_n5899;
  assign new_n5904 = ~new_n3682 & n77;
  assign new_n5905 = ~new_n891 & new_n3677;
  assign new_n5906 = new_n5905 ^ new_n5904;
  assign new_n5907 = n78 & new_n3676;
  assign new_n5908 = n76 & new_n3688;
  assign new_n5909 = new_n5908 ^ new_n5907;
  assign new_n5910 = new_n5909 ^ new_n5906;
  assign new_n5911 = new_n5910 ^ n39;
  assign new_n5912 = new_n5911 ^ new_n5903;
  assign new_n5913 = new_n5692 ^ new_n5680;
  assign new_n5914 = ~new_n5913 & new_n5689;
  assign new_n5915 = new_n5914 ^ new_n5692;
  assign new_n5916 = new_n5915 ^ new_n5912;
  assign new_n5917 = ~new_n3143 & n80;
  assign new_n5918 = new_n1161 & new_n3138;
  assign new_n5919 = new_n5918 ^ new_n5917;
  assign new_n5920 = n81 & new_n3137;
  assign new_n5921 = n79 & new_n3149;
  assign new_n5922 = new_n5921 ^ new_n5920;
  assign new_n5923 = new_n5922 ^ new_n5919;
  assign new_n5924 = new_n5923 ^ n36;
  assign new_n5925 = new_n5924 ^ new_n5916;
  assign new_n5926 = new_n5705 ^ new_n5693;
  assign new_n5927 = ~new_n5697 & new_n5926;
  assign new_n5928 = new_n5927 ^ new_n5696;
  assign new_n5929 = new_n5928 ^ new_n5925;
  assign new_n5930 = ~new_n2672 & n83;
  assign new_n5931 = new_n1468 & new_n2667;
  assign new_n5932 = new_n5931 ^ new_n5930;
  assign new_n5933 = n84 & new_n2666;
  assign new_n5934 = n82 & new_n2664;
  assign new_n5935 = new_n5934 ^ new_n5933;
  assign new_n5936 = new_n5935 ^ new_n5932;
  assign new_n5937 = new_n5936 ^ n33;
  assign new_n5938 = new_n5937 ^ new_n5929;
  assign new_n5939 = new_n5718 ^ new_n5706;
  assign new_n5940 = ~new_n5939 & new_n5715;
  assign new_n5941 = new_n5940 ^ new_n5718;
  assign new_n5942 = new_n5941 ^ new_n5938;
  assign new_n5943 = n86 & new_n2246;
  assign new_n5944 = new_n1811 & new_n2241;
  assign new_n5945 = new_n5944 ^ new_n5943;
  assign new_n5946 = n87 & new_n2240;
  assign new_n5947 = n85 & new_n2391;
  assign new_n5948 = new_n5947 ^ new_n5946;
  assign new_n5949 = new_n5948 ^ new_n5945;
  assign new_n5950 = new_n5949 ^ n30;
  assign new_n5951 = new_n5950 ^ new_n5942;
  assign new_n5952 = new_n5731 ^ new_n5719;
  assign new_n5953 = ~new_n5952 & new_n5728;
  assign new_n5954 = new_n5953 ^ new_n5731;
  assign new_n5955 = new_n5954 ^ new_n5951;
  assign new_n5956 = n89 & new_n1874;
  assign new_n5957 = new_n1864 & new_n2193;
  assign new_n5958 = new_n5957 ^ new_n5956;
  assign new_n5959 = n90 & new_n1863;
  assign new_n5960 = n88 & new_n1868;
  assign new_n5961 = new_n5960 ^ new_n5959;
  assign new_n5962 = new_n5961 ^ new_n5958;
  assign new_n5963 = new_n5962 ^ n27;
  assign new_n5964 = new_n5963 ^ new_n5955;
  assign new_n5965 = new_n5744 ^ new_n5732;
  assign new_n5966 = ~new_n5965 & new_n5741;
  assign new_n5967 = new_n5966 ^ new_n5744;
  assign new_n5968 = new_n5967 ^ new_n5964;
  assign new_n5969 = ~new_n1506 & n92;
  assign new_n5970 = new_n1501 & new_n2628;
  assign new_n5971 = new_n5970 ^ new_n5969;
  assign new_n5972 = n93 & new_n1500;
  assign new_n5973 = n91 & new_n1512;
  assign new_n5974 = new_n5973 ^ new_n5972;
  assign new_n5975 = new_n5974 ^ new_n5971;
  assign new_n5976 = new_n5975 ^ n24;
  assign new_n5977 = new_n5976 ^ new_n5968;
  assign new_n5978 = new_n5757 ^ new_n5745;
  assign new_n5979 = ~new_n5978 & new_n5754;
  assign new_n5980 = new_n5979 ^ new_n5757;
  assign new_n5981 = new_n5980 ^ new_n5977;
  assign new_n5982 = ~new_n1198 & n95;
  assign new_n5983 = new_n1193 & new_n3095;
  assign new_n5984 = new_n5983 ^ new_n5982;
  assign new_n5985 = n96 & new_n1192;
  assign new_n5986 = n94 & new_n1204;
  assign new_n5987 = new_n5986 ^ new_n5985;
  assign new_n5988 = new_n5987 ^ new_n5984;
  assign new_n5989 = new_n5988 ^ n21;
  assign new_n5990 = new_n5989 ^ new_n5981;
  assign new_n5991 = new_n5770 ^ new_n5758;
  assign new_n5992 = ~new_n5991 & new_n5767;
  assign new_n5993 = new_n5992 ^ new_n5770;
  assign new_n5994 = new_n5993 ^ new_n5990;
  assign new_n5995 = ~new_n930 & n98;
  assign new_n5996 = new_n925 & new_n3604;
  assign new_n5997 = new_n5996 ^ new_n5995;
  assign new_n5998 = n99 & new_n924;
  assign new_n5999 = n97 & new_n936;
  assign new_n6000 = new_n5999 ^ new_n5998;
  assign new_n6001 = new_n6000 ^ new_n5997;
  assign new_n6002 = new_n6001 ^ n18;
  assign new_n6003 = new_n6002 ^ new_n5994;
  assign new_n6004 = new_n5783 ^ new_n5771;
  assign new_n6005 = ~new_n6004 & new_n5780;
  assign new_n6006 = new_n6005 ^ new_n5783;
  assign new_n6007 = new_n6006 ^ new_n6003;
  assign new_n6008 = n101 & new_n707;
  assign new_n6009 = new_n701 & new_n4159;
  assign new_n6010 = new_n6009 ^ new_n6008;
  assign new_n6011 = n102 & new_n700;
  assign new_n6012 = n100 & new_n787;
  assign new_n6013 = new_n6012 ^ new_n6011;
  assign new_n6014 = new_n6013 ^ new_n6010;
  assign new_n6015 = new_n6014 ^ n15;
  assign new_n6016 = new_n6015 ^ new_n6007;
  assign new_n6017 = new_n5796 ^ new_n5784;
  assign new_n6018 = ~new_n6017 & new_n5793;
  assign new_n6019 = new_n6018 ^ new_n5796;
  assign new_n6020 = new_n6019 ^ new_n6016;
  assign new_n6021 = n104 & new_n499;
  assign new_n6022 = ~new_n506 & ~new_n4754;
  assign new_n6023 = new_n6022 ^ new_n6021;
  assign new_n6024 = ~new_n505 & n105;
  assign new_n6025 = n103 & new_n579;
  assign new_n6026 = new_n6025 ^ new_n6024;
  assign new_n6027 = new_n6026 ^ new_n6023;
  assign new_n6028 = new_n6027 ^ n12;
  assign new_n6029 = new_n6028 ^ new_n6020;
  assign new_n6030 = new_n5809 ^ new_n5797;
  assign new_n6031 = ~new_n6030 & new_n5806;
  assign new_n6032 = new_n6031 ^ new_n5809;
  assign new_n6033 = new_n6032 ^ new_n6029;
  assign new_n6034 = n107 & new_n354;
  assign new_n6035 = ~new_n5377 & new_n349;
  assign new_n6036 = new_n6035 ^ new_n6034;
  assign new_n6037 = n108 & new_n348;
  assign new_n6038 = n106 & new_n391;
  assign new_n6039 = new_n6038 ^ new_n6037;
  assign new_n6040 = new_n6039 ^ new_n6036;
  assign new_n6041 = new_n6040 ^ n9;
  assign new_n6042 = new_n6041 ^ new_n6033;
  assign new_n6043 = new_n5822 ^ new_n5810;
  assign new_n6044 = ~new_n6043 & new_n5819;
  assign new_n6045 = new_n6044 ^ new_n5822;
  assign new_n6046 = new_n6045 ^ new_n6042;
  assign new_n6047 = n110 & new_n218;
  assign new_n6048 = n111 ^ n110;
  assign new_n6049 = new_n6048 ^ new_n5392;
  assign new_n6050 = new_n208 & new_n6049;
  assign new_n6051 = new_n6050 ^ new_n6047;
  assign new_n6052 = n111 & new_n207;
  assign new_n6053 = n109 & new_n212;
  assign new_n6054 = new_n6053 ^ new_n6052;
  assign new_n6055 = new_n6054 ^ new_n6051;
  assign new_n6056 = new_n6055 ^ n6;
  assign new_n6057 = new_n6056 ^ new_n6046;
  assign new_n6058 = new_n5836 ^ new_n5823;
  assign new_n6059 = ~new_n6058 & new_n5833;
  assign new_n6060 = new_n6059 ^ new_n5836;
  assign new_n6061 = new_n6060 ^ new_n6057;
  assign new_n6062 = n112 & new_n180;
  assign new_n6063 = n2 & n113;
  assign new_n6064 = new_n6063 ^ new_n6062;
  assign new_n6065 = new_n6064 ^ n3;
  assign new_n6066 = ~new_n5844 & n113;
  assign new_n6067 = ~n113 & ~new_n5843;
  assign new_n6068 = new_n6067 ^ new_n6066;
  assign new_n6069 = new_n155 & new_n6068;
  assign new_n6070 = new_n6069 ^ n2;
  assign new_n6071 = new_n6070 ^ n114;
  assign new_n6072 = new_n6071 ^ new_n6065;
  assign new_n6073 = ~n1 & new_n6072;
  assign new_n6074 = new_n6073 ^ new_n6071;
  assign new_n6075 = new_n6074 ^ new_n6061;
  assign new_n6076 = new_n5855 ^ new_n5837;
  assign new_n6077 = ~new_n6076 & new_n5852;
  assign new_n6078 = new_n6077 ^ new_n5855;
  assign new_n6079 = new_n6078 ^ new_n6075;
  assign new_n6080 = ~new_n4212 & n75;
  assign new_n6081 = ~new_n737 & new_n4201;
  assign new_n6082 = new_n6081 ^ new_n6080;
  assign new_n6083 = n76 & new_n4200;
  assign new_n6084 = n74 & new_n4206;
  assign new_n6085 = new_n6084 ^ new_n6083;
  assign new_n6086 = new_n6085 ^ new_n6082;
  assign new_n6087 = new_n6086 ^ n42;
  assign new_n6088 = new_n5902 ^ new_n5890;
  assign new_n6089 = ~new_n5899 & new_n6088;
  assign new_n6090 = new_n6089 ^ new_n5902;
  assign new_n6091 = new_n6090 ^ new_n6087;
  assign new_n6092 = ~new_n5424 & n69;
  assign new_n6093 = ~new_n339 & new_n5419;
  assign new_n6094 = new_n6093 ^ new_n6092;
  assign new_n6095 = n70 & new_n5418;
  assign new_n6096 = n68 & new_n5648;
  assign new_n6097 = new_n6096 ^ new_n6095;
  assign new_n6098 = new_n6097 ^ new_n6094;
  assign new_n6099 = new_n6098 ^ n48;
  assign new_n6100 = ~new_n5641 & ~new_n5867;
  assign new_n6101 = n51 & new_n6100;
  assign new_n6102 = new_n6101 ^ new_n6099;
  assign new_n6103 = n51 ^ n50;
  assign new_n6104 = ~new_n6103 & new_n5640;
  assign new_n6105 = new_n6104 ^ new_n5640;
  assign new_n6106 = ~new_n151 & new_n6105;
  assign new_n6107 = n67 & new_n5640;
  assign new_n6108 = new_n6107 ^ new_n6106;
  assign new_n6109 = ~new_n5640 & n50;
  assign new_n6110 = new_n6109 ^ new_n5864;
  assign new_n6111 = ~new_n6110 & n66;
  assign new_n6112 = new_n6111 ^ new_n6108;
  assign new_n6113 = new_n6112 ^ n51;
  assign new_n6114 = ~new_n5864 & n50;
  assign new_n6115 = n65 & new_n6114;
  assign new_n6116 = ~new_n6113 & new_n6115;
  assign new_n6117 = new_n6116 ^ new_n6113;
  assign new_n6118 = ~n50 & new_n5863;
  assign new_n6119 = n65 & new_n6118;
  assign new_n6120 = ~new_n6119 & new_n6117;
  assign new_n6121 = new_n6120 ^ new_n6102;
  assign new_n6122 = new_n5876 ^ new_n5867;
  assign new_n6123 = ~new_n6122 & new_n5868;
  assign new_n6124 = new_n6123 ^ new_n5858;
  assign new_n6125 = new_n6124 ^ new_n6121;
  assign new_n6126 = new_n5889 ^ new_n5877;
  assign new_n6127 = ~new_n5886 & new_n6126;
  assign new_n6128 = new_n6127 ^ new_n5889;
  assign new_n6129 = new_n6128 ^ new_n6125;
  assign new_n6130 = ~new_n4804 & n72;
  assign new_n6131 = new_n534 & new_n4799;
  assign new_n6132 = new_n6131 ^ new_n6130;
  assign new_n6133 = n73 & new_n4798;
  assign new_n6134 = n71 & new_n4810;
  assign new_n6135 = new_n6134 ^ new_n6133;
  assign new_n6136 = new_n6135 ^ new_n6132;
  assign new_n6137 = new_n6136 ^ n45;
  assign new_n6138 = new_n6137 ^ new_n6129;
  assign new_n6139 = new_n6138 ^ new_n6091;
  assign new_n6140 = ~new_n3682 & n78;
  assign new_n6141 = ~new_n982 & new_n3677;
  assign new_n6142 = new_n6141 ^ new_n6140;
  assign new_n6143 = n79 & new_n3676;
  assign new_n6144 = n77 & new_n3688;
  assign new_n6145 = new_n6144 ^ new_n6143;
  assign new_n6146 = new_n6145 ^ new_n6142;
  assign new_n6147 = new_n6146 ^ n39;
  assign new_n6148 = new_n6147 ^ new_n6139;
  assign new_n6149 = new_n5915 ^ new_n5903;
  assign new_n6150 = ~new_n5912 & new_n6149;
  assign new_n6151 = new_n6150 ^ new_n5915;
  assign new_n6152 = new_n6151 ^ new_n6148;
  assign new_n6153 = ~new_n3143 & n81;
  assign new_n6154 = new_n1263 & new_n3138;
  assign new_n6155 = new_n6154 ^ new_n6153;
  assign new_n6156 = n82 & new_n3137;
  assign new_n6157 = n80 & new_n3149;
  assign new_n6158 = new_n6157 ^ new_n6156;
  assign new_n6159 = new_n6158 ^ new_n6155;
  assign new_n6160 = new_n6159 ^ n36;
  assign new_n6161 = new_n6160 ^ new_n6152;
  assign new_n6162 = new_n5928 ^ new_n5916;
  assign new_n6163 = ~new_n5925 & new_n6162;
  assign new_n6164 = new_n6163 ^ new_n5928;
  assign new_n6165 = new_n6164 ^ new_n6161;
  assign new_n6166 = ~new_n2672 & n84;
  assign new_n6167 = new_n1584 & new_n2667;
  assign new_n6168 = new_n6167 ^ new_n6166;
  assign new_n6169 = n85 & new_n2666;
  assign new_n6170 = n83 & new_n2664;
  assign new_n6171 = new_n6170 ^ new_n6169;
  assign new_n6172 = new_n6171 ^ new_n6168;
  assign new_n6173 = new_n6172 ^ n33;
  assign new_n6174 = new_n6173 ^ new_n6165;
  assign new_n6175 = new_n5941 ^ new_n5929;
  assign new_n6176 = ~new_n5938 & new_n6175;
  assign new_n6177 = new_n6176 ^ new_n5941;
  assign new_n6178 = new_n6177 ^ new_n6174;
  assign new_n6179 = n87 & new_n2246;
  assign new_n6180 = new_n1940 & new_n2241;
  assign new_n6181 = new_n6180 ^ new_n6179;
  assign new_n6182 = n88 & new_n2240;
  assign new_n6183 = n86 & new_n2391;
  assign new_n6184 = new_n6183 ^ new_n6182;
  assign new_n6185 = new_n6184 ^ new_n6181;
  assign new_n6186 = new_n6185 ^ n30;
  assign new_n6187 = new_n6186 ^ new_n6178;
  assign new_n6188 = new_n5954 ^ new_n5942;
  assign new_n6189 = ~new_n5951 & new_n6188;
  assign new_n6190 = new_n6189 ^ new_n5954;
  assign new_n6191 = new_n6190 ^ new_n6187;
  assign new_n6192 = n90 & new_n1874;
  assign new_n6193 = new_n1864 & new_n2341;
  assign new_n6194 = new_n6193 ^ new_n6192;
  assign new_n6195 = n91 & new_n1863;
  assign new_n6196 = n89 & new_n1868;
  assign new_n6197 = new_n6196 ^ new_n6195;
  assign new_n6198 = new_n6197 ^ new_n6194;
  assign new_n6199 = new_n6198 ^ n27;
  assign new_n6200 = new_n6199 ^ new_n6191;
  assign new_n6201 = new_n5967 ^ new_n5955;
  assign new_n6202 = ~new_n5964 & new_n6201;
  assign new_n6203 = new_n6202 ^ new_n5967;
  assign new_n6204 = new_n6203 ^ new_n6200;
  assign new_n6205 = ~new_n1506 & n93;
  assign new_n6206 = new_n1501 & new_n2785;
  assign new_n6207 = new_n6206 ^ new_n6205;
  assign new_n6208 = n94 & new_n1500;
  assign new_n6209 = n92 & new_n1512;
  assign new_n6210 = new_n6209 ^ new_n6208;
  assign new_n6211 = new_n6210 ^ new_n6207;
  assign new_n6212 = new_n6211 ^ n24;
  assign new_n6213 = new_n6212 ^ new_n6204;
  assign new_n6214 = new_n5980 ^ new_n5968;
  assign new_n6215 = ~new_n5977 & new_n6214;
  assign new_n6216 = new_n6215 ^ new_n5980;
  assign new_n6217 = new_n6216 ^ new_n6213;
  assign new_n6218 = ~new_n1198 & n96;
  assign new_n6219 = new_n1193 & new_n3273;
  assign new_n6220 = new_n6219 ^ new_n6218;
  assign new_n6221 = n97 & new_n1192;
  assign new_n6222 = n95 & new_n1204;
  assign new_n6223 = new_n6222 ^ new_n6221;
  assign new_n6224 = new_n6223 ^ new_n6220;
  assign new_n6225 = new_n6224 ^ n21;
  assign new_n6226 = new_n6225 ^ new_n6217;
  assign new_n6227 = new_n5993 ^ new_n5981;
  assign new_n6228 = ~new_n5990 & new_n6227;
  assign new_n6229 = new_n6228 ^ new_n5993;
  assign new_n6230 = new_n6229 ^ new_n6226;
  assign new_n6231 = ~new_n930 & n99;
  assign new_n6232 = new_n925 & new_n3789;
  assign new_n6233 = new_n6232 ^ new_n6231;
  assign new_n6234 = n100 & new_n924;
  assign new_n6235 = n98 & new_n936;
  assign new_n6236 = new_n6235 ^ new_n6234;
  assign new_n6237 = new_n6236 ^ new_n6233;
  assign new_n6238 = new_n6237 ^ n18;
  assign new_n6239 = new_n6238 ^ new_n6230;
  assign new_n6240 = new_n6006 ^ new_n5994;
  assign new_n6241 = ~new_n6003 & new_n6240;
  assign new_n6242 = new_n6241 ^ new_n6006;
  assign new_n6243 = new_n6242 ^ new_n6239;
  assign new_n6244 = n102 & new_n707;
  assign new_n6245 = new_n701 & new_n4368;
  assign new_n6246 = new_n6245 ^ new_n6244;
  assign new_n6247 = n103 & new_n700;
  assign new_n6248 = n101 & new_n787;
  assign new_n6249 = new_n6248 ^ new_n6247;
  assign new_n6250 = new_n6249 ^ new_n6246;
  assign new_n6251 = new_n6250 ^ n15;
  assign new_n6252 = new_n6251 ^ new_n6243;
  assign new_n6253 = new_n6019 ^ new_n6007;
  assign new_n6254 = ~new_n6016 & new_n6253;
  assign new_n6255 = new_n6254 ^ new_n6019;
  assign new_n6256 = new_n6255 ^ new_n6252;
  assign new_n6257 = n105 & new_n499;
  assign new_n6258 = ~new_n506 & ~new_n4961;
  assign new_n6259 = new_n6258 ^ new_n6257;
  assign new_n6260 = ~new_n505 & n106;
  assign new_n6261 = n104 & new_n579;
  assign new_n6262 = new_n6261 ^ new_n6260;
  assign new_n6263 = new_n6262 ^ new_n6259;
  assign new_n6264 = new_n6263 ^ n12;
  assign new_n6265 = new_n6264 ^ new_n6256;
  assign new_n6266 = new_n6032 ^ new_n6020;
  assign new_n6267 = ~new_n6029 & new_n6266;
  assign new_n6268 = new_n6267 ^ new_n6032;
  assign new_n6269 = new_n6268 ^ new_n6265;
  assign new_n6270 = n108 & new_n354;
  assign new_n6271 = new_n349 & new_n5604;
  assign new_n6272 = new_n6271 ^ new_n6270;
  assign new_n6273 = n109 & new_n348;
  assign new_n6274 = n107 & new_n391;
  assign new_n6275 = new_n6274 ^ new_n6273;
  assign new_n6276 = new_n6275 ^ new_n6272;
  assign new_n6277 = new_n6276 ^ n9;
  assign new_n6278 = new_n6277 ^ new_n6269;
  assign new_n6279 = new_n6045 ^ new_n6033;
  assign new_n6280 = ~new_n6042 & new_n6279;
  assign new_n6281 = new_n6280 ^ new_n6045;
  assign new_n6282 = new_n6281 ^ new_n6278;
  assign new_n6283 = n111 & new_n218;
  assign new_n6284 = new_n5621 ^ n112;
  assign new_n6285 = ~new_n6284 & new_n208;
  assign new_n6286 = new_n6285 ^ new_n6283;
  assign new_n6287 = n112 & new_n207;
  assign new_n6288 = n110 & new_n212;
  assign new_n6289 = new_n6288 ^ new_n6287;
  assign new_n6290 = new_n6289 ^ new_n6286;
  assign new_n6291 = new_n6290 ^ n6;
  assign new_n6292 = new_n6291 ^ new_n6282;
  assign new_n6293 = new_n6060 ^ new_n6046;
  assign new_n6294 = ~new_n6057 & new_n6293;
  assign new_n6295 = new_n6294 ^ new_n6060;
  assign new_n6296 = new_n6295 ^ new_n6292;
  assign new_n6297 = ~n114 & ~new_n6066;
  assign new_n6298 = ~new_n6067 & n114;
  assign new_n6299 = new_n6298 ^ new_n6297;
  assign new_n6300 = new_n155 & new_n6299;
  assign new_n6301 = new_n6300 ^ n2;
  assign new_n6302 = new_n6301 ^ n115;
  assign new_n6303 = n114 ^ n3;
  assign new_n6304 = ~n113 & n3;
  assign new_n6305 = new_n6304 ^ new_n6303;
  assign new_n6306 = ~n2 & new_n6305;
  assign new_n6307 = new_n6306 ^ new_n6303;
  assign new_n6308 = new_n6307 ^ new_n6302;
  assign new_n6309 = ~n1 & new_n6308;
  assign new_n6310 = new_n6309 ^ new_n6302;
  assign new_n6311 = new_n6310 ^ new_n6296;
  assign new_n6312 = new_n6078 ^ new_n6061;
  assign new_n6313 = ~new_n6075 & new_n6312;
  assign new_n6314 = new_n6313 ^ new_n6078;
  assign new_n6315 = new_n6314 ^ new_n6311;
  assign new_n6316 = ~new_n3682 & n79;
  assign new_n6317 = new_n1069 & new_n3677;
  assign new_n6318 = new_n6317 ^ new_n6316;
  assign new_n6319 = n80 & new_n3676;
  assign new_n6320 = n78 & new_n3688;
  assign new_n6321 = new_n6320 ^ new_n6319;
  assign new_n6322 = new_n6321 ^ new_n6318;
  assign new_n6323 = new_n6322 ^ n39;
  assign new_n6324 = new_n6151 ^ new_n6139;
  assign new_n6325 = ~new_n6148 & new_n6324;
  assign new_n6326 = new_n6325 ^ new_n6151;
  assign new_n6327 = new_n6326 ^ new_n6323;
  assign new_n6328 = new_n6125 ^ new_n6120;
  assign new_n6329 = new_n6120 ^ new_n6101;
  assign new_n6330 = ~new_n6328 & new_n6329;
  assign new_n6331 = new_n6330 ^ new_n6120;
  assign new_n6332 = ~new_n5424 & n70;
  assign new_n6333 = ~new_n402 & new_n5419;
  assign new_n6334 = new_n6333 ^ new_n6332;
  assign new_n6335 = n71 & new_n5418;
  assign new_n6336 = n69 & new_n5648;
  assign new_n6337 = new_n6336 ^ new_n6335;
  assign new_n6338 = new_n6337 ^ new_n6334;
  assign new_n6339 = new_n6338 ^ n48;
  assign new_n6340 = new_n6339 ^ new_n6331;
  assign new_n6341 = ~new_n259 & new_n6105;
  assign new_n6342 = ~new_n6110 & n67;
  assign new_n6343 = new_n6342 ^ new_n6341;
  assign new_n6344 = n68 & new_n6104;
  assign new_n6345 = ~new_n5640 & n51;
  assign new_n6346 = new_n6345 ^ new_n5864;
  assign new_n6347 = ~new_n6346 & new_n6103;
  assign new_n6348 = n66 & new_n6347;
  assign new_n6349 = new_n6348 ^ new_n6344;
  assign new_n6350 = new_n6349 ^ new_n6343;
  assign new_n6351 = new_n6350 ^ n51;
  assign new_n6352 = n52 ^ n51;
  assign new_n6353 = n65 & new_n6352;
  assign new_n6354 = new_n6353 ^ new_n6351;
  assign new_n6355 = new_n6354 ^ new_n6339;
  assign new_n6356 = new_n6355 ^ new_n6340;
  assign new_n6357 = new_n6356 ^ new_n6339;
  assign new_n6358 = new_n6099 & new_n6124;
  assign new_n6359 = new_n6358 ^ new_n6357;
  assign new_n6360 = ~new_n4804 & n73;
  assign new_n6361 = new_n595 & new_n4799;
  assign new_n6362 = new_n6361 ^ new_n6360;
  assign new_n6363 = n74 & new_n4798;
  assign new_n6364 = n72 & new_n4810;
  assign new_n6365 = new_n6364 ^ new_n6363;
  assign new_n6366 = new_n6365 ^ new_n6362;
  assign new_n6367 = new_n6366 ^ n45;
  assign new_n6368 = new_n6367 ^ new_n6359;
  assign new_n6369 = new_n6137 ^ new_n6125;
  assign new_n6370 = ~new_n6369 & new_n6129;
  assign new_n6371 = new_n6370 ^ new_n6128;
  assign new_n6372 = new_n6371 ^ new_n6368;
  assign new_n6373 = ~new_n4212 & n76;
  assign new_n6374 = ~new_n812 & new_n4201;
  assign new_n6375 = new_n6374 ^ new_n6373;
  assign new_n6376 = n77 & new_n4200;
  assign new_n6377 = n75 & new_n4206;
  assign new_n6378 = new_n6377 ^ new_n6376;
  assign new_n6379 = new_n6378 ^ new_n6375;
  assign new_n6380 = new_n6379 ^ n42;
  assign new_n6381 = new_n6380 ^ new_n6372;
  assign new_n6382 = new_n6138 ^ new_n6087;
  assign new_n6383 = ~new_n6382 & new_n6091;
  assign new_n6384 = new_n6383 ^ new_n6090;
  assign new_n6385 = new_n6384 ^ new_n6381;
  assign new_n6386 = new_n6385 ^ new_n6327;
  assign new_n6387 = ~new_n3143 & n82;
  assign new_n6388 = new_n1363 & new_n3138;
  assign new_n6389 = new_n6388 ^ new_n6387;
  assign new_n6390 = n83 & new_n3137;
  assign new_n6391 = n81 & new_n3149;
  assign new_n6392 = new_n6391 ^ new_n6390;
  assign new_n6393 = new_n6392 ^ new_n6389;
  assign new_n6394 = new_n6393 ^ n36;
  assign new_n6395 = new_n6394 ^ new_n6386;
  assign new_n6396 = new_n6164 ^ new_n6152;
  assign new_n6397 = ~new_n6161 & new_n6396;
  assign new_n6398 = new_n6397 ^ new_n6164;
  assign new_n6399 = new_n6398 ^ new_n6395;
  assign new_n6400 = ~new_n2672 & n85;
  assign new_n6401 = new_n1694 & new_n2667;
  assign new_n6402 = new_n6401 ^ new_n6400;
  assign new_n6403 = n86 & new_n2666;
  assign new_n6404 = n84 & new_n2664;
  assign new_n6405 = new_n6404 ^ new_n6403;
  assign new_n6406 = new_n6405 ^ new_n6402;
  assign new_n6407 = new_n6406 ^ n33;
  assign new_n6408 = new_n6407 ^ new_n6399;
  assign new_n6409 = new_n6177 ^ new_n6173;
  assign new_n6410 = ~new_n6409 & new_n6174;
  assign new_n6411 = new_n6410 ^ new_n6165;
  assign new_n6412 = new_n6411 ^ new_n6408;
  assign new_n6413 = n88 & new_n2246;
  assign new_n6414 = new_n2063 & new_n2241;
  assign new_n6415 = new_n6414 ^ new_n6413;
  assign new_n6416 = n89 & new_n2240;
  assign new_n6417 = n87 & new_n2391;
  assign new_n6418 = new_n6417 ^ new_n6416;
  assign new_n6419 = new_n6418 ^ new_n6415;
  assign new_n6420 = new_n6419 ^ n30;
  assign new_n6421 = new_n6420 ^ new_n6412;
  assign new_n6422 = new_n6190 ^ new_n6178;
  assign new_n6423 = ~new_n6187 & new_n6422;
  assign new_n6424 = new_n6423 ^ new_n6190;
  assign new_n6425 = new_n6424 ^ new_n6421;
  assign new_n6426 = n91 & new_n1874;
  assign new_n6427 = new_n1864 & new_n2481;
  assign new_n6428 = new_n6427 ^ new_n6426;
  assign new_n6429 = n92 & new_n1863;
  assign new_n6430 = n90 & new_n1868;
  assign new_n6431 = new_n6430 ^ new_n6429;
  assign new_n6432 = new_n6431 ^ new_n6428;
  assign new_n6433 = new_n6432 ^ n27;
  assign new_n6434 = new_n6433 ^ new_n6425;
  assign new_n6435 = new_n6203 ^ new_n6191;
  assign new_n6436 = ~new_n6200 & new_n6435;
  assign new_n6437 = new_n6436 ^ new_n6203;
  assign new_n6438 = new_n6437 ^ new_n6434;
  assign new_n6439 = ~new_n1506 & n94;
  assign new_n6440 = new_n1501 & new_n2934;
  assign new_n6441 = new_n6440 ^ new_n6439;
  assign new_n6442 = n95 & new_n1500;
  assign new_n6443 = n93 & new_n1512;
  assign new_n6444 = new_n6443 ^ new_n6442;
  assign new_n6445 = new_n6444 ^ new_n6441;
  assign new_n6446 = new_n6445 ^ n24;
  assign new_n6447 = new_n6446 ^ new_n6438;
  assign new_n6448 = new_n6216 ^ new_n6204;
  assign new_n6449 = ~new_n6213 & new_n6448;
  assign new_n6450 = new_n6449 ^ new_n6216;
  assign new_n6451 = new_n6450 ^ new_n6447;
  assign new_n6452 = ~new_n1198 & n97;
  assign new_n6453 = new_n1193 & new_n3435;
  assign new_n6454 = new_n6453 ^ new_n6452;
  assign new_n6455 = n98 & new_n1192;
  assign new_n6456 = n96 & new_n1204;
  assign new_n6457 = new_n6456 ^ new_n6455;
  assign new_n6458 = new_n6457 ^ new_n6454;
  assign new_n6459 = new_n6458 ^ n21;
  assign new_n6460 = new_n6459 ^ new_n6451;
  assign new_n6461 = new_n6229 ^ new_n6217;
  assign new_n6462 = ~new_n6226 & new_n6461;
  assign new_n6463 = new_n6462 ^ new_n6229;
  assign new_n6464 = new_n6463 ^ new_n6460;
  assign new_n6465 = ~new_n930 & n100;
  assign new_n6466 = new_n925 & new_n3972;
  assign new_n6467 = new_n6466 ^ new_n6465;
  assign new_n6468 = n101 & new_n924;
  assign new_n6469 = n99 & new_n936;
  assign new_n6470 = new_n6469 ^ new_n6468;
  assign new_n6471 = new_n6470 ^ new_n6467;
  assign new_n6472 = new_n6471 ^ n18;
  assign new_n6473 = new_n6472 ^ new_n6464;
  assign new_n6474 = new_n6242 ^ new_n6230;
  assign new_n6475 = ~new_n6239 & new_n6474;
  assign new_n6476 = new_n6475 ^ new_n6242;
  assign new_n6477 = new_n6476 ^ new_n6473;
  assign new_n6478 = n103 & new_n707;
  assign new_n6479 = ~new_n4556 & new_n701;
  assign new_n6480 = new_n6479 ^ new_n6478;
  assign new_n6481 = n104 & new_n700;
  assign new_n6482 = n102 & new_n787;
  assign new_n6483 = new_n6482 ^ new_n6481;
  assign new_n6484 = new_n6483 ^ new_n6480;
  assign new_n6485 = new_n6484 ^ n15;
  assign new_n6486 = new_n6485 ^ new_n6477;
  assign new_n6487 = new_n6255 ^ new_n6243;
  assign new_n6488 = ~new_n6252 & new_n6487;
  assign new_n6489 = new_n6488 ^ new_n6255;
  assign new_n6490 = new_n6489 ^ new_n6486;
  assign new_n6491 = n106 & new_n499;
  assign new_n6492 = ~new_n506 & ~new_n5164;
  assign new_n6493 = new_n6492 ^ new_n6491;
  assign new_n6494 = ~new_n505 & n107;
  assign new_n6495 = n105 & new_n579;
  assign new_n6496 = new_n6495 ^ new_n6494;
  assign new_n6497 = new_n6496 ^ new_n6493;
  assign new_n6498 = new_n6497 ^ n12;
  assign new_n6499 = new_n6498 ^ new_n6490;
  assign new_n6500 = new_n6268 ^ new_n6256;
  assign new_n6501 = ~new_n6265 & new_n6500;
  assign new_n6502 = new_n6501 ^ new_n6268;
  assign new_n6503 = new_n6502 ^ new_n6499;
  assign new_n6504 = n109 & new_n354;
  assign new_n6505 = new_n349 & new_n5825;
  assign new_n6506 = new_n6505 ^ new_n6504;
  assign new_n6507 = n110 & new_n348;
  assign new_n6508 = n108 & new_n391;
  assign new_n6509 = new_n6508 ^ new_n6507;
  assign new_n6510 = new_n6509 ^ new_n6506;
  assign new_n6511 = new_n6510 ^ n9;
  assign new_n6512 = new_n6511 ^ new_n6503;
  assign new_n6513 = new_n6281 ^ new_n6269;
  assign new_n6514 = ~new_n6278 & new_n6513;
  assign new_n6515 = new_n6514 ^ new_n6281;
  assign new_n6516 = new_n6515 ^ new_n6512;
  assign new_n6517 = n112 & new_n218;
  assign new_n6518 = new_n5845 ^ n113;
  assign new_n6519 = ~new_n6518 & new_n208;
  assign new_n6520 = new_n6519 ^ new_n6517;
  assign new_n6521 = n113 & new_n207;
  assign new_n6522 = n111 & new_n212;
  assign new_n6523 = new_n6522 ^ new_n6521;
  assign new_n6524 = new_n6523 ^ new_n6520;
  assign new_n6525 = new_n6524 ^ n6;
  assign new_n6526 = new_n6525 ^ new_n6516;
  assign new_n6527 = new_n6295 ^ new_n6282;
  assign new_n6528 = ~new_n6292 & new_n6527;
  assign new_n6529 = new_n6528 ^ new_n6295;
  assign new_n6530 = new_n6529 ^ new_n6526;
  assign new_n6531 = n115 ^ n3;
  assign new_n6532 = ~n114 & n3;
  assign new_n6533 = new_n6532 ^ new_n6531;
  assign new_n6534 = ~n2 & new_n6533;
  assign new_n6535 = new_n6534 ^ new_n6531;
  assign new_n6536 = ~new_n6297 & n115;
  assign new_n6537 = ~n115 & ~new_n6298;
  assign new_n6538 = new_n6537 ^ new_n6536;
  assign new_n6539 = new_n155 & new_n6538;
  assign new_n6540 = new_n6539 ^ n2;
  assign new_n6541 = new_n6540 ^ n116;
  assign new_n6542 = new_n6541 ^ new_n6535;
  assign new_n6543 = ~n1 & new_n6542;
  assign new_n6544 = new_n6543 ^ new_n6541;
  assign new_n6545 = new_n6544 ^ new_n6530;
  assign new_n6546 = new_n6314 ^ new_n6296;
  assign new_n6547 = ~new_n6311 & new_n6546;
  assign new_n6548 = new_n6547 ^ new_n6314;
  assign new_n6549 = new_n6548 ^ new_n6545;
  assign new_n6550 = ~new_n4212 & n77;
  assign new_n6551 = ~new_n891 & new_n4201;
  assign new_n6552 = new_n6551 ^ new_n6550;
  assign new_n6553 = n78 & new_n4200;
  assign new_n6554 = n76 & new_n4206;
  assign new_n6555 = new_n6554 ^ new_n6553;
  assign new_n6556 = new_n6555 ^ new_n6552;
  assign new_n6557 = new_n6556 ^ n42;
  assign new_n6558 = new_n6384 ^ new_n6372;
  assign new_n6559 = ~new_n6381 & new_n6558;
  assign new_n6560 = new_n6559 ^ new_n6384;
  assign new_n6561 = new_n6560 ^ new_n6557;
  assign new_n6562 = new_n6358 ^ new_n6339;
  assign new_n6563 = new_n6562 ^ new_n6355;
  assign new_n6564 = new_n6563 ^ new_n6339;
  assign new_n6565 = ~new_n6563 & new_n6356;
  assign new_n6566 = new_n6565 ^ new_n6356;
  assign new_n6567 = new_n6564 & new_n6566;
  assign new_n6568 = new_n6567 ^ new_n6339;
  assign new_n6569 = ~new_n6359 & ~new_n6568;
  assign new_n6570 = new_n6569 ^ new_n6565;
  assign new_n6571 = new_n6570 ^ new_n6339;
  assign new_n6572 = new_n6571 ^ new_n6358;
  assign new_n6573 = new_n6101 & new_n6120;
  assign new_n6574 = ~new_n6573 & new_n6354;
  assign new_n6575 = new_n6574 ^ new_n6572;
  assign new_n6576 = ~new_n5424 & n71;
  assign new_n6577 = ~new_n459 & new_n5419;
  assign new_n6578 = new_n6577 ^ new_n6576;
  assign new_n6579 = n72 & new_n5418;
  assign new_n6580 = n70 & new_n5648;
  assign new_n6581 = new_n6580 ^ new_n6579;
  assign new_n6582 = new_n6581 ^ new_n6578;
  assign new_n6583 = new_n6582 ^ n48;
  assign new_n6584 = new_n6583 ^ new_n6575;
  assign new_n6585 = ~n51 & ~n52;
  assign new_n6586 = new_n6585 ^ new_n6352;
  assign new_n6587 = new_n6586 ^ n53;
  assign new_n6588 = ~n65 & ~new_n6587;
  assign new_n6589 = n66 ^ n52;
  assign new_n6590 = ~new_n6589 & new_n6352;
  assign new_n6591 = new_n6590 ^ n51;
  assign new_n6592 = new_n6591 ^ n53;
  assign new_n6593 = new_n6592 ^ new_n6588;
  assign new_n6594 = ~new_n6574 & new_n6351;
  assign new_n6595 = new_n6594 ^ new_n6593;
  assign new_n6596 = ~new_n6110 & n68;
  assign new_n6597 = ~new_n304 & new_n6105;
  assign new_n6598 = new_n6597 ^ new_n6596;
  assign new_n6599 = n69 & new_n6104;
  assign new_n6600 = n67 & new_n6347;
  assign new_n6601 = new_n6600 ^ new_n6599;
  assign new_n6602 = new_n6601 ^ new_n6598;
  assign new_n6603 = new_n6602 ^ n51;
  assign new_n6604 = new_n6603 ^ new_n6595;
  assign new_n6605 = new_n6604 ^ new_n6584;
  assign new_n6606 = ~new_n4804 & n74;
  assign new_n6607 = new_n660 & new_n4799;
  assign new_n6608 = new_n6607 ^ new_n6606;
  assign new_n6609 = n75 & new_n4798;
  assign new_n6610 = n73 & new_n4810;
  assign new_n6611 = new_n6610 ^ new_n6609;
  assign new_n6612 = new_n6611 ^ new_n6608;
  assign new_n6613 = new_n6612 ^ n45;
  assign new_n6614 = new_n6613 ^ new_n6605;
  assign new_n6615 = new_n6371 ^ new_n6359;
  assign new_n6616 = ~new_n6368 & new_n6615;
  assign new_n6617 = new_n6616 ^ new_n6371;
  assign new_n6618 = new_n6617 ^ new_n6614;
  assign new_n6619 = new_n6618 ^ new_n6561;
  assign new_n6620 = ~new_n3682 & n80;
  assign new_n6621 = new_n1161 & new_n3677;
  assign new_n6622 = new_n6621 ^ new_n6620;
  assign new_n6623 = n81 & new_n3676;
  assign new_n6624 = n79 & new_n3688;
  assign new_n6625 = new_n6624 ^ new_n6623;
  assign new_n6626 = new_n6625 ^ new_n6622;
  assign new_n6627 = new_n6626 ^ n39;
  assign new_n6628 = new_n6627 ^ new_n6619;
  assign new_n6629 = new_n6385 ^ new_n6323;
  assign new_n6630 = ~new_n6629 & new_n6327;
  assign new_n6631 = new_n6630 ^ new_n6326;
  assign new_n6632 = new_n6631 ^ new_n6628;
  assign new_n6633 = ~new_n3143 & n83;
  assign new_n6634 = new_n1468 & new_n3138;
  assign new_n6635 = new_n6634 ^ new_n6633;
  assign new_n6636 = n84 & new_n3137;
  assign new_n6637 = n82 & new_n3149;
  assign new_n6638 = new_n6637 ^ new_n6636;
  assign new_n6639 = new_n6638 ^ new_n6635;
  assign new_n6640 = new_n6639 ^ n36;
  assign new_n6641 = new_n6640 ^ new_n6632;
  assign new_n6642 = new_n6398 ^ new_n6386;
  assign new_n6643 = ~new_n6395 & new_n6642;
  assign new_n6644 = new_n6643 ^ new_n6398;
  assign new_n6645 = new_n6644 ^ new_n6641;
  assign new_n6646 = ~new_n2672 & n86;
  assign new_n6647 = new_n1811 & new_n2667;
  assign new_n6648 = new_n6647 ^ new_n6646;
  assign new_n6649 = n87 & new_n2666;
  assign new_n6650 = n85 & new_n2664;
  assign new_n6651 = new_n6650 ^ new_n6649;
  assign new_n6652 = new_n6651 ^ new_n6648;
  assign new_n6653 = new_n6652 ^ n33;
  assign new_n6654 = new_n6653 ^ new_n6645;
  assign new_n6655 = new_n6411 ^ new_n6407;
  assign new_n6656 = ~new_n6655 & new_n6408;
  assign new_n6657 = new_n6656 ^ new_n6399;
  assign new_n6658 = new_n6657 ^ new_n6654;
  assign new_n6659 = n89 & new_n2246;
  assign new_n6660 = new_n2193 & new_n2241;
  assign new_n6661 = new_n6660 ^ new_n6659;
  assign new_n6662 = n90 & new_n2240;
  assign new_n6663 = n88 & new_n2391;
  assign new_n6664 = new_n6663 ^ new_n6662;
  assign new_n6665 = new_n6664 ^ new_n6661;
  assign new_n6666 = new_n6665 ^ n30;
  assign new_n6667 = new_n6666 ^ new_n6658;
  assign new_n6668 = new_n6424 ^ new_n6412;
  assign new_n6669 = ~new_n6421 & new_n6668;
  assign new_n6670 = new_n6669 ^ new_n6424;
  assign new_n6671 = new_n6670 ^ new_n6667;
  assign new_n6672 = n92 & new_n1874;
  assign new_n6673 = new_n1864 & new_n2628;
  assign new_n6674 = new_n6673 ^ new_n6672;
  assign new_n6675 = n93 & new_n1863;
  assign new_n6676 = n91 & new_n1868;
  assign new_n6677 = new_n6676 ^ new_n6675;
  assign new_n6678 = new_n6677 ^ new_n6674;
  assign new_n6679 = new_n6678 ^ n27;
  assign new_n6680 = new_n6679 ^ new_n6671;
  assign new_n6681 = new_n6437 ^ new_n6425;
  assign new_n6682 = ~new_n6434 & new_n6681;
  assign new_n6683 = new_n6682 ^ new_n6437;
  assign new_n6684 = new_n6683 ^ new_n6680;
  assign new_n6685 = ~new_n1506 & n95;
  assign new_n6686 = new_n1501 & new_n3095;
  assign new_n6687 = new_n6686 ^ new_n6685;
  assign new_n6688 = n96 & new_n1500;
  assign new_n6689 = n94 & new_n1512;
  assign new_n6690 = new_n6689 ^ new_n6688;
  assign new_n6691 = new_n6690 ^ new_n6687;
  assign new_n6692 = new_n6691 ^ n24;
  assign new_n6693 = new_n6692 ^ new_n6684;
  assign new_n6694 = new_n6450 ^ new_n6438;
  assign new_n6695 = ~new_n6447 & new_n6694;
  assign new_n6696 = new_n6695 ^ new_n6450;
  assign new_n6697 = new_n6696 ^ new_n6693;
  assign new_n6698 = ~new_n1198 & n98;
  assign new_n6699 = new_n1193 & new_n3604;
  assign new_n6700 = new_n6699 ^ new_n6698;
  assign new_n6701 = n99 & new_n1192;
  assign new_n6702 = n97 & new_n1204;
  assign new_n6703 = new_n6702 ^ new_n6701;
  assign new_n6704 = new_n6703 ^ new_n6700;
  assign new_n6705 = new_n6704 ^ n21;
  assign new_n6706 = new_n6705 ^ new_n6697;
  assign new_n6707 = new_n6463 ^ new_n6451;
  assign new_n6708 = ~new_n6460 & new_n6707;
  assign new_n6709 = new_n6708 ^ new_n6463;
  assign new_n6710 = new_n6709 ^ new_n6706;
  assign new_n6711 = ~new_n930 & n101;
  assign new_n6712 = new_n925 & new_n4159;
  assign new_n6713 = new_n6712 ^ new_n6711;
  assign new_n6714 = n102 & new_n924;
  assign new_n6715 = n100 & new_n936;
  assign new_n6716 = new_n6715 ^ new_n6714;
  assign new_n6717 = new_n6716 ^ new_n6713;
  assign new_n6718 = new_n6717 ^ n18;
  assign new_n6719 = new_n6718 ^ new_n6710;
  assign new_n6720 = new_n6476 ^ new_n6464;
  assign new_n6721 = ~new_n6473 & new_n6720;
  assign new_n6722 = new_n6721 ^ new_n6476;
  assign new_n6723 = new_n6722 ^ new_n6719;
  assign new_n6724 = n104 & new_n707;
  assign new_n6725 = ~new_n4754 & new_n701;
  assign new_n6726 = new_n6725 ^ new_n6724;
  assign new_n6727 = n105 & new_n700;
  assign new_n6728 = n103 & new_n787;
  assign new_n6729 = new_n6728 ^ new_n6727;
  assign new_n6730 = new_n6729 ^ new_n6726;
  assign new_n6731 = new_n6730 ^ n15;
  assign new_n6732 = new_n6731 ^ new_n6723;
  assign new_n6733 = new_n6489 ^ new_n6477;
  assign new_n6734 = ~new_n6486 & new_n6733;
  assign new_n6735 = new_n6734 ^ new_n6489;
  assign new_n6736 = new_n6735 ^ new_n6732;
  assign new_n6737 = n107 & new_n499;
  assign new_n6738 = ~new_n506 & ~new_n5377;
  assign new_n6739 = new_n6738 ^ new_n6737;
  assign new_n6740 = ~new_n505 & n108;
  assign new_n6741 = n106 & new_n579;
  assign new_n6742 = new_n6741 ^ new_n6740;
  assign new_n6743 = new_n6742 ^ new_n6739;
  assign new_n6744 = new_n6743 ^ n12;
  assign new_n6745 = new_n6744 ^ new_n6736;
  assign new_n6746 = new_n6502 ^ new_n6490;
  assign new_n6747 = ~new_n6499 & new_n6746;
  assign new_n6748 = new_n6747 ^ new_n6502;
  assign new_n6749 = new_n6748 ^ new_n6745;
  assign new_n6750 = n110 & new_n354;
  assign new_n6751 = new_n349 & new_n6049;
  assign new_n6752 = new_n6751 ^ new_n6750;
  assign new_n6753 = n111 & new_n348;
  assign new_n6754 = n109 & new_n391;
  assign new_n6755 = new_n6754 ^ new_n6753;
  assign new_n6756 = new_n6755 ^ new_n6752;
  assign new_n6757 = new_n6756 ^ n9;
  assign new_n6758 = new_n6757 ^ new_n6749;
  assign new_n6759 = new_n6515 ^ new_n6503;
  assign new_n6760 = ~new_n6512 & new_n6759;
  assign new_n6761 = new_n6760 ^ new_n6515;
  assign new_n6762 = new_n6761 ^ new_n6758;
  assign new_n6763 = n113 & new_n218;
  assign new_n6764 = new_n6068 ^ n114;
  assign new_n6765 = ~new_n6764 & new_n208;
  assign new_n6766 = new_n6765 ^ new_n6763;
  assign new_n6767 = n114 & new_n207;
  assign new_n6768 = n112 & new_n212;
  assign new_n6769 = new_n6768 ^ new_n6767;
  assign new_n6770 = new_n6769 ^ new_n6766;
  assign new_n6771 = new_n6770 ^ n6;
  assign new_n6772 = new_n6771 ^ new_n6762;
  assign new_n6773 = new_n6529 ^ new_n6516;
  assign new_n6774 = ~new_n6526 & new_n6773;
  assign new_n6775 = new_n6774 ^ new_n6529;
  assign new_n6776 = new_n6775 ^ new_n6772;
  assign new_n6777 = ~n116 & ~new_n6536;
  assign new_n6778 = ~new_n6537 & n116;
  assign new_n6779 = new_n6778 ^ new_n6777;
  assign new_n6780 = new_n155 & new_n6779;
  assign new_n6781 = new_n6780 ^ n2;
  assign new_n6782 = new_n6781 ^ n117;
  assign new_n6783 = n116 ^ n3;
  assign new_n6784 = ~n115 & ~new_n6531;
  assign new_n6785 = new_n6784 ^ new_n6783;
  assign new_n6786 = new_n6785 ^ n115;
  assign new_n6787 = ~new_n6786 & new_n241;
  assign new_n6788 = new_n6787 ^ new_n6784;
  assign new_n6789 = new_n6788 ^ n115;
  assign new_n6790 = new_n6789 ^ new_n6782;
  assign new_n6791 = ~n1 & ~new_n6790;
  assign new_n6792 = new_n6791 ^ new_n6782;
  assign new_n6793 = new_n6792 ^ new_n6776;
  assign new_n6794 = new_n6548 ^ new_n6530;
  assign new_n6795 = ~new_n6545 & new_n6794;
  assign new_n6796 = new_n6795 ^ new_n6548;
  assign new_n6797 = new_n6796 ^ new_n6793;
  assign new_n6798 = n54 ^ n53;
  assign new_n6799 = ~new_n6798 & new_n6352;
  assign new_n6800 = new_n6799 ^ new_n6352;
  assign new_n6801 = ~new_n151 & new_n6800;
  assign new_n6802 = n67 & new_n6352;
  assign new_n6803 = new_n6802 ^ new_n6801;
  assign new_n6804 = ~new_n6352 & n53;
  assign new_n6805 = new_n6804 ^ new_n6586;
  assign new_n6806 = ~new_n6805 & n66;
  assign new_n6807 = new_n6806 ^ new_n6803;
  assign new_n6808 = new_n6807 ^ n54;
  assign new_n6809 = ~new_n6352 & n54;
  assign new_n6810 = new_n6809 ^ new_n6586;
  assign new_n6811 = ~new_n6810 & new_n6798;
  assign new_n6812 = n65 & new_n6811;
  assign new_n6813 = new_n6812 ^ new_n6808;
  assign new_n6814 = ~new_n6353 & ~new_n6593;
  assign new_n6815 = n54 & new_n6814;
  assign new_n6816 = new_n6815 ^ new_n6813;
  assign new_n6817 = ~new_n6110 & n69;
  assign new_n6818 = ~new_n339 & new_n6105;
  assign new_n6819 = new_n6818 ^ new_n6817;
  assign new_n6820 = n70 & new_n6104;
  assign new_n6821 = n68 & new_n6347;
  assign new_n6822 = new_n6821 ^ new_n6820;
  assign new_n6823 = new_n6822 ^ new_n6819;
  assign new_n6824 = new_n6823 ^ n51;
  assign new_n6825 = new_n6824 ^ new_n6816;
  assign new_n6826 = new_n6603 ^ new_n6593;
  assign new_n6827 = ~new_n6826 & new_n6595;
  assign new_n6828 = new_n6827 ^ new_n6594;
  assign new_n6829 = new_n6828 ^ new_n6825;
  assign new_n6830 = ~new_n5424 & n72;
  assign new_n6831 = new_n534 & new_n5419;
  assign new_n6832 = new_n6831 ^ new_n6830;
  assign new_n6833 = n73 & new_n5418;
  assign new_n6834 = n71 & new_n5648;
  assign new_n6835 = new_n6834 ^ new_n6833;
  assign new_n6836 = new_n6835 ^ new_n6832;
  assign new_n6837 = new_n6836 ^ n48;
  assign new_n6838 = new_n6837 ^ new_n6829;
  assign new_n6839 = new_n6604 ^ new_n6583;
  assign new_n6840 = ~new_n6584 & ~new_n6839;
  assign new_n6841 = new_n6840 ^ new_n6575;
  assign new_n6842 = new_n6841 ^ new_n6838;
  assign new_n6843 = ~new_n4804 & n75;
  assign new_n6844 = ~new_n737 & new_n4799;
  assign new_n6845 = new_n6844 ^ new_n6843;
  assign new_n6846 = n74 & new_n4810;
  assign new_n6847 = n76 & new_n4798;
  assign new_n6848 = new_n6847 ^ new_n6846;
  assign new_n6849 = new_n6848 ^ new_n6845;
  assign new_n6850 = new_n6849 ^ n45;
  assign new_n6851 = new_n6850 ^ new_n6842;
  assign new_n6852 = new_n6617 ^ new_n6605;
  assign new_n6853 = ~new_n6852 & new_n6614;
  assign new_n6854 = new_n6853 ^ new_n6617;
  assign new_n6855 = new_n6854 ^ new_n6851;
  assign new_n6856 = ~new_n4212 & n78;
  assign new_n6857 = ~new_n982 & new_n4201;
  assign new_n6858 = new_n6857 ^ new_n6856;
  assign new_n6859 = n79 & new_n4200;
  assign new_n6860 = n77 & new_n4206;
  assign new_n6861 = new_n6860 ^ new_n6859;
  assign new_n6862 = new_n6861 ^ new_n6858;
  assign new_n6863 = new_n6862 ^ n42;
  assign new_n6864 = new_n6863 ^ new_n6855;
  assign new_n6865 = new_n6618 ^ new_n6557;
  assign new_n6866 = new_n6561 & new_n6865;
  assign new_n6867 = new_n6866 ^ new_n6560;
  assign new_n6868 = new_n6867 ^ new_n6864;
  assign new_n6869 = new_n6631 ^ new_n6619;
  assign new_n6870 = ~new_n6869 & new_n6628;
  assign new_n6871 = new_n6870 ^ new_n6631;
  assign new_n6872 = new_n6871 ^ new_n6868;
  assign new_n6873 = ~new_n3682 & n81;
  assign new_n6874 = new_n1263 & new_n3677;
  assign new_n6875 = new_n6874 ^ new_n6873;
  assign new_n6876 = n80 & new_n3688;
  assign new_n6877 = n82 & new_n3676;
  assign new_n6878 = new_n6877 ^ new_n6876;
  assign new_n6879 = new_n6878 ^ new_n6875;
  assign new_n6880 = new_n6879 ^ n39;
  assign new_n6881 = new_n6880 ^ new_n6872;
  assign new_n6882 = ~new_n3143 & n84;
  assign new_n6883 = new_n1584 & new_n3138;
  assign new_n6884 = new_n6883 ^ new_n6882;
  assign new_n6885 = n85 & new_n3137;
  assign new_n6886 = n83 & new_n3149;
  assign new_n6887 = new_n6886 ^ new_n6885;
  assign new_n6888 = new_n6887 ^ new_n6884;
  assign new_n6889 = new_n6888 ^ n36;
  assign new_n6890 = new_n6889 ^ new_n6881;
  assign new_n6891 = new_n6644 ^ new_n6632;
  assign new_n6892 = ~new_n6891 & new_n6641;
  assign new_n6893 = new_n6892 ^ new_n6644;
  assign new_n6894 = new_n6893 ^ new_n6890;
  assign new_n6895 = ~new_n2672 & n87;
  assign new_n6896 = new_n1940 & new_n2667;
  assign new_n6897 = new_n6896 ^ new_n6895;
  assign new_n6898 = n88 & new_n2666;
  assign new_n6899 = n86 & new_n2664;
  assign new_n6900 = new_n6899 ^ new_n6898;
  assign new_n6901 = new_n6900 ^ new_n6897;
  assign new_n6902 = new_n6901 ^ n33;
  assign new_n6903 = new_n6902 ^ new_n6894;
  assign new_n6904 = new_n6657 ^ new_n6653;
  assign new_n6905 = ~new_n6654 & ~new_n6904;
  assign new_n6906 = new_n6905 ^ new_n6645;
  assign new_n6907 = new_n6906 ^ new_n6903;
  assign new_n6908 = n90 & new_n2246;
  assign new_n6909 = new_n2241 & new_n2341;
  assign new_n6910 = new_n6909 ^ new_n6908;
  assign new_n6911 = n91 & new_n2240;
  assign new_n6912 = n89 & new_n2391;
  assign new_n6913 = new_n6912 ^ new_n6911;
  assign new_n6914 = new_n6913 ^ new_n6910;
  assign new_n6915 = new_n6914 ^ n30;
  assign new_n6916 = new_n6915 ^ new_n6907;
  assign new_n6917 = new_n6670 ^ new_n6658;
  assign new_n6918 = ~new_n6917 & new_n6667;
  assign new_n6919 = new_n6918 ^ new_n6670;
  assign new_n6920 = new_n6919 ^ new_n6916;
  assign new_n6921 = n93 & new_n1874;
  assign new_n6922 = new_n1864 & new_n2785;
  assign new_n6923 = new_n6922 ^ new_n6921;
  assign new_n6924 = n94 & new_n1863;
  assign new_n6925 = n92 & new_n1868;
  assign new_n6926 = new_n6925 ^ new_n6924;
  assign new_n6927 = new_n6926 ^ new_n6923;
  assign new_n6928 = new_n6927 ^ n27;
  assign new_n6929 = new_n6928 ^ new_n6920;
  assign new_n6930 = new_n6683 ^ new_n6671;
  assign new_n6931 = ~new_n6930 & new_n6680;
  assign new_n6932 = new_n6931 ^ new_n6683;
  assign new_n6933 = new_n6932 ^ new_n6929;
  assign new_n6934 = ~new_n1506 & n96;
  assign new_n6935 = new_n1501 & new_n3273;
  assign new_n6936 = new_n6935 ^ new_n6934;
  assign new_n6937 = n97 & new_n1500;
  assign new_n6938 = n95 & new_n1512;
  assign new_n6939 = new_n6938 ^ new_n6937;
  assign new_n6940 = new_n6939 ^ new_n6936;
  assign new_n6941 = new_n6940 ^ n24;
  assign new_n6942 = new_n6941 ^ new_n6933;
  assign new_n6943 = new_n6696 ^ new_n6684;
  assign new_n6944 = ~new_n6943 & new_n6693;
  assign new_n6945 = new_n6944 ^ new_n6696;
  assign new_n6946 = new_n6945 ^ new_n6942;
  assign new_n6947 = ~new_n1198 & n99;
  assign new_n6948 = new_n1193 & new_n3789;
  assign new_n6949 = new_n6948 ^ new_n6947;
  assign new_n6950 = n100 & new_n1192;
  assign new_n6951 = n98 & new_n1204;
  assign new_n6952 = new_n6951 ^ new_n6950;
  assign new_n6953 = new_n6952 ^ new_n6949;
  assign new_n6954 = new_n6953 ^ n21;
  assign new_n6955 = new_n6954 ^ new_n6946;
  assign new_n6956 = new_n6709 ^ new_n6697;
  assign new_n6957 = ~new_n6956 & new_n6706;
  assign new_n6958 = new_n6957 ^ new_n6709;
  assign new_n6959 = new_n6958 ^ new_n6955;
  assign new_n6960 = ~new_n930 & n102;
  assign new_n6961 = new_n925 & new_n4368;
  assign new_n6962 = new_n6961 ^ new_n6960;
  assign new_n6963 = n103 & new_n924;
  assign new_n6964 = n101 & new_n936;
  assign new_n6965 = new_n6964 ^ new_n6963;
  assign new_n6966 = new_n6965 ^ new_n6962;
  assign new_n6967 = new_n6966 ^ n18;
  assign new_n6968 = new_n6967 ^ new_n6959;
  assign new_n6969 = new_n6722 ^ new_n6710;
  assign new_n6970 = ~new_n6969 & new_n6719;
  assign new_n6971 = new_n6970 ^ new_n6722;
  assign new_n6972 = new_n6971 ^ new_n6968;
  assign new_n6973 = n105 & new_n707;
  assign new_n6974 = ~new_n4961 & new_n701;
  assign new_n6975 = new_n6974 ^ new_n6973;
  assign new_n6976 = n106 & new_n700;
  assign new_n6977 = n104 & new_n787;
  assign new_n6978 = new_n6977 ^ new_n6976;
  assign new_n6979 = new_n6978 ^ new_n6975;
  assign new_n6980 = new_n6979 ^ n15;
  assign new_n6981 = new_n6980 ^ new_n6972;
  assign new_n6982 = new_n6735 ^ new_n6723;
  assign new_n6983 = ~new_n6982 & new_n6732;
  assign new_n6984 = new_n6983 ^ new_n6735;
  assign new_n6985 = new_n6984 ^ new_n6981;
  assign new_n6986 = n108 & new_n499;
  assign new_n6987 = ~new_n506 & new_n5604;
  assign new_n6988 = new_n6987 ^ new_n6986;
  assign new_n6989 = ~new_n505 & n109;
  assign new_n6990 = n107 & new_n579;
  assign new_n6991 = new_n6990 ^ new_n6989;
  assign new_n6992 = new_n6991 ^ new_n6988;
  assign new_n6993 = new_n6992 ^ n12;
  assign new_n6994 = new_n6993 ^ new_n6985;
  assign new_n6995 = new_n6748 ^ new_n6736;
  assign new_n6996 = ~new_n6995 & new_n6745;
  assign new_n6997 = new_n6996 ^ new_n6748;
  assign new_n6998 = new_n6997 ^ new_n6994;
  assign new_n6999 = n111 & new_n354;
  assign new_n7000 = ~new_n6284 & new_n349;
  assign new_n7001 = new_n7000 ^ new_n6999;
  assign new_n7002 = n112 & new_n348;
  assign new_n7003 = n110 & new_n391;
  assign new_n7004 = new_n7003 ^ new_n7002;
  assign new_n7005 = new_n7004 ^ new_n7001;
  assign new_n7006 = new_n7005 ^ n9;
  assign new_n7007 = new_n7006 ^ new_n6998;
  assign new_n7008 = new_n6761 ^ new_n6749;
  assign new_n7009 = ~new_n7008 & new_n6758;
  assign new_n7010 = new_n7009 ^ new_n6761;
  assign new_n7011 = new_n7010 ^ new_n7007;
  assign new_n7012 = n114 & new_n218;
  assign new_n7013 = new_n6299 ^ n115;
  assign new_n7014 = ~new_n7013 & new_n208;
  assign new_n7015 = new_n7014 ^ new_n7012;
  assign new_n7016 = n115 & new_n207;
  assign new_n7017 = n113 & new_n212;
  assign new_n7018 = new_n7017 ^ new_n7016;
  assign new_n7019 = new_n7018 ^ new_n7015;
  assign new_n7020 = new_n7019 ^ n6;
  assign new_n7021 = new_n7020 ^ new_n7011;
  assign new_n7022 = new_n6775 ^ new_n6762;
  assign new_n7023 = ~new_n7022 & new_n6772;
  assign new_n7024 = new_n7023 ^ new_n6775;
  assign new_n7025 = new_n7024 ^ new_n7021;
  assign new_n7026 = ~new_n6777 & n117;
  assign new_n7027 = ~n117 & ~new_n6778;
  assign new_n7028 = new_n7027 ^ new_n7026;
  assign new_n7029 = new_n155 & new_n7028;
  assign new_n7030 = new_n7029 ^ n2;
  assign new_n7031 = new_n7030 ^ n118;
  assign new_n7032 = n117 ^ n3;
  assign new_n7033 = ~n116 & ~new_n6783;
  assign new_n7034 = new_n7033 ^ new_n7032;
  assign new_n7035 = new_n7034 ^ n116;
  assign new_n7036 = ~new_n7035 & new_n241;
  assign new_n7037 = new_n7036 ^ new_n7033;
  assign new_n7038 = new_n7037 ^ n116;
  assign new_n7039 = new_n7038 ^ new_n7031;
  assign new_n7040 = ~n1 & ~new_n7039;
  assign new_n7041 = new_n7040 ^ new_n7031;
  assign new_n7042 = new_n7041 ^ new_n7025;
  assign new_n7043 = new_n6796 ^ new_n6776;
  assign new_n7044 = ~new_n7043 & new_n6793;
  assign new_n7045 = new_n7044 ^ new_n6796;
  assign new_n7046 = new_n7045 ^ new_n7042;
  assign new_n7047 = new_n6997 ^ new_n6985;
  assign new_n7048 = ~new_n6994 & new_n7047;
  assign new_n7049 = new_n7048 ^ new_n6997;
  assign new_n7050 = n109 & new_n499;
  assign new_n7051 = ~new_n506 & new_n5825;
  assign new_n7052 = new_n7051 ^ new_n7050;
  assign new_n7053 = ~new_n505 & n110;
  assign new_n7054 = n108 & new_n579;
  assign new_n7055 = new_n7054 ^ new_n7053;
  assign new_n7056 = new_n7055 ^ new_n7052;
  assign new_n7057 = new_n7056 ^ n12;
  assign new_n7058 = ~new_n4212 & n79;
  assign new_n7059 = new_n1069 & new_n4201;
  assign new_n7060 = new_n7059 ^ new_n7058;
  assign new_n7061 = n80 & new_n4200;
  assign new_n7062 = n78 & new_n4206;
  assign new_n7063 = new_n7062 ^ new_n7061;
  assign new_n7064 = new_n7063 ^ new_n7060;
  assign new_n7065 = new_n7064 ^ n42;
  assign new_n7066 = new_n6867 ^ new_n6855;
  assign new_n7067 = ~new_n7066 & new_n6864;
  assign new_n7068 = new_n7067 ^ new_n6867;
  assign new_n7069 = new_n7068 ^ new_n7065;
  assign new_n7070 = new_n6813 & new_n6815;
  assign new_n7071 = ~new_n259 & new_n6800;
  assign new_n7072 = ~new_n6805 & n67;
  assign new_n7073 = new_n7072 ^ new_n7071;
  assign new_n7074 = n68 & new_n6799;
  assign new_n7075 = n66 & new_n6811;
  assign new_n7076 = new_n7075 ^ new_n7074;
  assign new_n7077 = new_n7076 ^ new_n7073;
  assign new_n7078 = new_n7077 ^ n54;
  assign new_n7079 = n55 ^ n54;
  assign new_n7080 = n65 & new_n7079;
  assign new_n7081 = new_n7080 ^ new_n7078;
  assign new_n7082 = new_n7081 ^ new_n7070;
  assign new_n7083 = ~new_n6110 & n70;
  assign new_n7084 = ~new_n402 & new_n6105;
  assign new_n7085 = new_n7084 ^ new_n7083;
  assign new_n7086 = n71 & new_n6104;
  assign new_n7087 = n69 & new_n6347;
  assign new_n7088 = new_n7087 ^ new_n7086;
  assign new_n7089 = new_n7088 ^ new_n7085;
  assign new_n7090 = new_n7089 ^ n51;
  assign new_n7091 = new_n7090 ^ new_n7082;
  assign new_n7092 = new_n6828 ^ new_n6816;
  assign new_n7093 = ~new_n6825 & new_n7092;
  assign new_n7094 = new_n7093 ^ new_n6828;
  assign new_n7095 = new_n7094 ^ new_n7091;
  assign new_n7096 = ~new_n5424 & n73;
  assign new_n7097 = new_n595 & new_n5419;
  assign new_n7098 = new_n7097 ^ new_n7096;
  assign new_n7099 = n74 & new_n5418;
  assign new_n7100 = n72 & new_n5648;
  assign new_n7101 = new_n7100 ^ new_n7099;
  assign new_n7102 = new_n7101 ^ new_n7098;
  assign new_n7103 = new_n7102 ^ n48;
  assign new_n7104 = new_n7103 ^ new_n7095;
  assign new_n7105 = new_n6841 ^ new_n6829;
  assign new_n7106 = ~new_n6838 & ~new_n7105;
  assign new_n7107 = new_n7106 ^ new_n6841;
  assign new_n7108 = new_n7107 ^ new_n7104;
  assign new_n7109 = ~new_n4804 & n76;
  assign new_n7110 = ~new_n812 & new_n4799;
  assign new_n7111 = new_n7110 ^ new_n7109;
  assign new_n7112 = n77 & new_n4798;
  assign new_n7113 = n75 & new_n4810;
  assign new_n7114 = new_n7113 ^ new_n7112;
  assign new_n7115 = new_n7114 ^ new_n7111;
  assign new_n7116 = new_n7115 ^ n45;
  assign new_n7117 = new_n7116 ^ new_n7108;
  assign new_n7118 = new_n6854 ^ new_n6842;
  assign new_n7119 = ~new_n7118 & new_n6851;
  assign new_n7120 = new_n7119 ^ new_n6854;
  assign new_n7121 = new_n7120 ^ new_n7117;
  assign new_n7122 = new_n7121 ^ new_n7069;
  assign new_n7123 = ~new_n3682 & n82;
  assign new_n7124 = new_n1363 & new_n3677;
  assign new_n7125 = new_n7124 ^ new_n7123;
  assign new_n7126 = n83 & new_n3676;
  assign new_n7127 = n81 & new_n3688;
  assign new_n7128 = new_n7127 ^ new_n7126;
  assign new_n7129 = new_n7128 ^ new_n7125;
  assign new_n7130 = new_n7129 ^ n39;
  assign new_n7131 = new_n7130 ^ new_n7122;
  assign new_n7132 = new_n6880 ^ new_n6868;
  assign new_n7133 = ~new_n6872 & new_n7132;
  assign new_n7134 = new_n7133 ^ new_n6871;
  assign new_n7135 = new_n7134 ^ new_n7131;
  assign new_n7136 = ~new_n3143 & n85;
  assign new_n7137 = new_n1694 & new_n3138;
  assign new_n7138 = new_n7137 ^ new_n7136;
  assign new_n7139 = n86 & new_n3137;
  assign new_n7140 = n84 & new_n3149;
  assign new_n7141 = new_n7140 ^ new_n7139;
  assign new_n7142 = new_n7141 ^ new_n7138;
  assign new_n7143 = new_n7142 ^ n36;
  assign new_n7144 = new_n7143 ^ new_n7135;
  assign new_n7145 = new_n6893 ^ new_n6881;
  assign new_n7146 = ~new_n7145 & new_n6890;
  assign new_n7147 = new_n7146 ^ new_n6893;
  assign new_n7148 = new_n7147 ^ new_n7144;
  assign new_n7149 = ~new_n2672 & n88;
  assign new_n7150 = new_n2063 & new_n2667;
  assign new_n7151 = new_n7150 ^ new_n7149;
  assign new_n7152 = n89 & new_n2666;
  assign new_n7153 = n87 & new_n2664;
  assign new_n7154 = new_n7153 ^ new_n7152;
  assign new_n7155 = new_n7154 ^ new_n7151;
  assign new_n7156 = new_n7155 ^ n33;
  assign new_n7157 = new_n7156 ^ new_n7148;
  assign new_n7158 = new_n6906 ^ new_n6894;
  assign new_n7159 = new_n6903 & new_n7158;
  assign new_n7160 = new_n7159 ^ new_n6906;
  assign new_n7161 = new_n7160 ^ new_n7157;
  assign new_n7162 = n91 & new_n2246;
  assign new_n7163 = new_n2241 & new_n2481;
  assign new_n7164 = new_n7163 ^ new_n7162;
  assign new_n7165 = n92 & new_n2240;
  assign new_n7166 = n90 & new_n2391;
  assign new_n7167 = new_n7166 ^ new_n7165;
  assign new_n7168 = new_n7167 ^ new_n7164;
  assign new_n7169 = new_n7168 ^ n30;
  assign new_n7170 = new_n7169 ^ new_n7161;
  assign new_n7171 = new_n6919 ^ new_n6907;
  assign new_n7172 = ~new_n6916 & new_n7171;
  assign new_n7173 = new_n7172 ^ new_n6919;
  assign new_n7174 = new_n7173 ^ new_n7170;
  assign new_n7175 = n94 & new_n1874;
  assign new_n7176 = new_n1864 & new_n2934;
  assign new_n7177 = new_n7176 ^ new_n7175;
  assign new_n7178 = n95 & new_n1863;
  assign new_n7179 = n93 & new_n1868;
  assign new_n7180 = new_n7179 ^ new_n7178;
  assign new_n7181 = new_n7180 ^ new_n7177;
  assign new_n7182 = new_n7181 ^ n27;
  assign new_n7183 = new_n7182 ^ new_n7174;
  assign new_n7184 = new_n6932 ^ new_n6920;
  assign new_n7185 = ~new_n6929 & new_n7184;
  assign new_n7186 = new_n7185 ^ new_n6932;
  assign new_n7187 = new_n7186 ^ new_n7183;
  assign new_n7188 = ~new_n1506 & n97;
  assign new_n7189 = new_n1501 & new_n3435;
  assign new_n7190 = new_n7189 ^ new_n7188;
  assign new_n7191 = n98 & new_n1500;
  assign new_n7192 = n96 & new_n1512;
  assign new_n7193 = new_n7192 ^ new_n7191;
  assign new_n7194 = new_n7193 ^ new_n7190;
  assign new_n7195 = new_n7194 ^ n24;
  assign new_n7196 = new_n7195 ^ new_n7187;
  assign new_n7197 = new_n6945 ^ new_n6933;
  assign new_n7198 = ~new_n6942 & new_n7197;
  assign new_n7199 = new_n7198 ^ new_n6945;
  assign new_n7200 = new_n7199 ^ new_n7196;
  assign new_n7201 = ~new_n1198 & n100;
  assign new_n7202 = new_n1193 & new_n3972;
  assign new_n7203 = new_n7202 ^ new_n7201;
  assign new_n7204 = n101 & new_n1192;
  assign new_n7205 = n99 & new_n1204;
  assign new_n7206 = new_n7205 ^ new_n7204;
  assign new_n7207 = new_n7206 ^ new_n7203;
  assign new_n7208 = new_n7207 ^ n21;
  assign new_n7209 = new_n7208 ^ new_n7200;
  assign new_n7210 = new_n6958 ^ new_n6946;
  assign new_n7211 = ~new_n6955 & new_n7210;
  assign new_n7212 = new_n7211 ^ new_n6958;
  assign new_n7213 = new_n7212 ^ new_n7209;
  assign new_n7214 = ~new_n930 & n103;
  assign new_n7215 = ~new_n4556 & new_n925;
  assign new_n7216 = new_n7215 ^ new_n7214;
  assign new_n7217 = n104 & new_n924;
  assign new_n7218 = n102 & new_n936;
  assign new_n7219 = new_n7218 ^ new_n7217;
  assign new_n7220 = new_n7219 ^ new_n7216;
  assign new_n7221 = new_n7220 ^ n18;
  assign new_n7222 = new_n7221 ^ new_n7213;
  assign new_n7223 = new_n6971 ^ new_n6959;
  assign new_n7224 = ~new_n6968 & new_n7223;
  assign new_n7225 = new_n7224 ^ new_n6971;
  assign new_n7226 = new_n7225 ^ new_n7222;
  assign new_n7227 = n106 & new_n707;
  assign new_n7228 = ~new_n5164 & new_n701;
  assign new_n7229 = new_n7228 ^ new_n7227;
  assign new_n7230 = n107 & new_n700;
  assign new_n7231 = n105 & new_n787;
  assign new_n7232 = new_n7231 ^ new_n7230;
  assign new_n7233 = new_n7232 ^ new_n7229;
  assign new_n7234 = new_n7233 ^ n15;
  assign new_n7235 = new_n7234 ^ new_n7226;
  assign new_n7236 = new_n6984 ^ new_n6972;
  assign new_n7237 = ~new_n6981 & new_n7236;
  assign new_n7238 = new_n7237 ^ new_n6984;
  assign new_n7239 = new_n7238 ^ new_n7235;
  assign new_n7240 = new_n7239 ^ new_n7057;
  assign new_n7241 = new_n7240 ^ new_n7049;
  assign new_n7242 = n112 & new_n354;
  assign new_n7243 = ~new_n6518 & new_n349;
  assign new_n7244 = new_n7243 ^ new_n7242;
  assign new_n7245 = n113 & new_n348;
  assign new_n7246 = n111 & new_n391;
  assign new_n7247 = new_n7246 ^ new_n7245;
  assign new_n7248 = new_n7247 ^ new_n7244;
  assign new_n7249 = new_n7248 ^ n9;
  assign new_n7250 = new_n7249 ^ new_n7241;
  assign new_n7251 = new_n7010 ^ new_n6998;
  assign new_n7252 = ~new_n7007 & new_n7251;
  assign new_n7253 = new_n7252 ^ new_n7010;
  assign new_n7254 = new_n7253 ^ new_n7250;
  assign new_n7255 = n115 & new_n218;
  assign new_n7256 = new_n6538 ^ n116;
  assign new_n7257 = ~new_n7256 & new_n208;
  assign new_n7258 = new_n7257 ^ new_n7255;
  assign new_n7259 = n116 & new_n207;
  assign new_n7260 = n114 & new_n212;
  assign new_n7261 = new_n7260 ^ new_n7259;
  assign new_n7262 = new_n7261 ^ new_n7258;
  assign new_n7263 = new_n7262 ^ n6;
  assign new_n7264 = new_n7263 ^ new_n7254;
  assign new_n7265 = new_n7024 ^ new_n7011;
  assign new_n7266 = ~new_n7021 & new_n7265;
  assign new_n7267 = new_n7266 ^ new_n7024;
  assign new_n7268 = new_n7267 ^ new_n7264;
  assign new_n7269 = n117 & new_n180;
  assign new_n7270 = n2 & n118;
  assign new_n7271 = new_n7270 ^ new_n7269;
  assign new_n7272 = new_n7271 ^ n3;
  assign new_n7273 = ~n118 & ~new_n7026;
  assign new_n7274 = ~new_n7027 & n118;
  assign new_n7275 = new_n7274 ^ new_n7273;
  assign new_n7276 = new_n155 & new_n7275;
  assign new_n7277 = new_n7276 ^ n2;
  assign new_n7278 = new_n7277 ^ n119;
  assign new_n7279 = new_n7278 ^ new_n7272;
  assign new_n7280 = ~n1 & new_n7279;
  assign new_n7281 = new_n7280 ^ new_n7278;
  assign new_n7282 = new_n7281 ^ new_n7268;
  assign new_n7283 = new_n7045 ^ new_n7025;
  assign new_n7284 = ~new_n7042 & new_n7283;
  assign new_n7285 = new_n7284 ^ new_n7045;
  assign new_n7286 = new_n7285 ^ new_n7282;
  assign new_n7287 = ~new_n4804 & n77;
  assign new_n7288 = ~new_n891 & new_n4799;
  assign new_n7289 = new_n7288 ^ new_n7287;
  assign new_n7290 = n78 & new_n4798;
  assign new_n7291 = n76 & new_n4810;
  assign new_n7292 = new_n7291 ^ new_n7290;
  assign new_n7293 = new_n7292 ^ new_n7289;
  assign new_n7294 = new_n7293 ^ n45;
  assign new_n7295 = new_n7120 ^ new_n7108;
  assign new_n7296 = ~new_n7295 & new_n7117;
  assign new_n7297 = new_n7296 ^ new_n7120;
  assign new_n7298 = new_n7297 ^ new_n7294;
  assign new_n7299 = ~new_n7070 & ~new_n7080;
  assign new_n7300 = ~new_n7299 & new_n7078;
  assign new_n7301 = ~new_n6805 & n68;
  assign new_n7302 = ~new_n304 & new_n6800;
  assign new_n7303 = new_n7302 ^ new_n7301;
  assign new_n7304 = n69 & new_n6799;
  assign new_n7305 = n67 & new_n6811;
  assign new_n7306 = new_n7305 ^ new_n7304;
  assign new_n7307 = new_n7306 ^ new_n7303;
  assign new_n7308 = new_n7307 ^ n54;
  assign new_n7309 = n66 ^ n55;
  assign new_n7310 = ~new_n7309 & new_n7079;
  assign new_n7311 = new_n7310 ^ n54;
  assign new_n7312 = new_n7311 ^ n56;
  assign new_n7313 = n54 & n55;
  assign new_n7314 = new_n7313 ^ n56;
  assign new_n7315 = ~n65 & new_n7314;
  assign new_n7316 = new_n7315 ^ new_n7312;
  assign new_n7317 = new_n7316 ^ new_n7308;
  assign new_n7318 = new_n7317 ^ new_n7300;
  assign new_n7319 = ~new_n6110 & n71;
  assign new_n7320 = ~new_n459 & new_n6105;
  assign new_n7321 = new_n7320 ^ new_n7319;
  assign new_n7322 = n72 & new_n6104;
  assign new_n7323 = n70 & new_n6347;
  assign new_n7324 = new_n7323 ^ new_n7322;
  assign new_n7325 = new_n7324 ^ new_n7321;
  assign new_n7326 = new_n7325 ^ n51;
  assign new_n7327 = new_n7326 ^ new_n7318;
  assign new_n7328 = new_n7094 ^ new_n7082;
  assign new_n7329 = ~new_n7091 & new_n7328;
  assign new_n7330 = new_n7329 ^ new_n7094;
  assign new_n7331 = new_n7330 ^ new_n7327;
  assign new_n7332 = ~new_n5424 & n74;
  assign new_n7333 = new_n660 & new_n5419;
  assign new_n7334 = new_n7333 ^ new_n7332;
  assign new_n7335 = n75 & new_n5418;
  assign new_n7336 = n73 & new_n5648;
  assign new_n7337 = new_n7336 ^ new_n7335;
  assign new_n7338 = new_n7337 ^ new_n7334;
  assign new_n7339 = new_n7338 ^ n48;
  assign new_n7340 = new_n7339 ^ new_n7331;
  assign new_n7341 = new_n7107 ^ new_n7095;
  assign new_n7342 = ~new_n7104 & ~new_n7341;
  assign new_n7343 = new_n7342 ^ new_n7107;
  assign new_n7344 = new_n7343 ^ new_n7340;
  assign new_n7345 = new_n7344 ^ new_n7298;
  assign new_n7346 = ~new_n4212 & n80;
  assign new_n7347 = new_n1161 & new_n4201;
  assign new_n7348 = new_n7347 ^ new_n7346;
  assign new_n7349 = n81 & new_n4200;
  assign new_n7350 = n79 & new_n4206;
  assign new_n7351 = new_n7350 ^ new_n7349;
  assign new_n7352 = new_n7351 ^ new_n7348;
  assign new_n7353 = new_n7352 ^ n42;
  assign new_n7354 = new_n7353 ^ new_n7345;
  assign new_n7355 = new_n7121 ^ new_n7065;
  assign new_n7356 = new_n7069 & new_n7355;
  assign new_n7357 = new_n7356 ^ new_n7068;
  assign new_n7358 = new_n7357 ^ new_n7354;
  assign new_n7359 = ~new_n3682 & n83;
  assign new_n7360 = new_n1468 & new_n3677;
  assign new_n7361 = new_n7360 ^ new_n7359;
  assign new_n7362 = n84 & new_n3676;
  assign new_n7363 = n82 & new_n3688;
  assign new_n7364 = new_n7363 ^ new_n7362;
  assign new_n7365 = new_n7364 ^ new_n7361;
  assign new_n7366 = new_n7365 ^ n39;
  assign new_n7367 = new_n7366 ^ new_n7358;
  assign new_n7368 = new_n7134 ^ new_n7122;
  assign new_n7369 = ~new_n7368 & new_n7131;
  assign new_n7370 = new_n7369 ^ new_n7134;
  assign new_n7371 = new_n7370 ^ new_n7367;
  assign new_n7372 = ~new_n3143 & n86;
  assign new_n7373 = new_n1811 & new_n3138;
  assign new_n7374 = new_n7373 ^ new_n7372;
  assign new_n7375 = n87 & new_n3137;
  assign new_n7376 = n85 & new_n3149;
  assign new_n7377 = new_n7376 ^ new_n7375;
  assign new_n7378 = new_n7377 ^ new_n7374;
  assign new_n7379 = new_n7378 ^ n36;
  assign new_n7380 = new_n7379 ^ new_n7371;
  assign new_n7381 = new_n7147 ^ new_n7135;
  assign new_n7382 = ~new_n7381 & new_n7144;
  assign new_n7383 = new_n7382 ^ new_n7147;
  assign new_n7384 = new_n7383 ^ new_n7380;
  assign new_n7385 = ~new_n2672 & n89;
  assign new_n7386 = new_n2193 & new_n2667;
  assign new_n7387 = new_n7386 ^ new_n7385;
  assign new_n7388 = n90 & new_n2666;
  assign new_n7389 = n88 & new_n2664;
  assign new_n7390 = new_n7389 ^ new_n7388;
  assign new_n7391 = new_n7390 ^ new_n7387;
  assign new_n7392 = new_n7391 ^ n33;
  assign new_n7393 = new_n7392 ^ new_n7384;
  assign new_n7394 = new_n7160 ^ new_n7148;
  assign new_n7395 = new_n7157 & new_n7394;
  assign new_n7396 = new_n7395 ^ new_n7160;
  assign new_n7397 = new_n7396 ^ new_n7393;
  assign new_n7398 = n92 & new_n2246;
  assign new_n7399 = new_n2241 & new_n2628;
  assign new_n7400 = new_n7399 ^ new_n7398;
  assign new_n7401 = n93 & new_n2240;
  assign new_n7402 = n91 & new_n2391;
  assign new_n7403 = new_n7402 ^ new_n7401;
  assign new_n7404 = new_n7403 ^ new_n7400;
  assign new_n7405 = new_n7404 ^ n30;
  assign new_n7406 = new_n7405 ^ new_n7397;
  assign new_n7407 = new_n7173 ^ new_n7161;
  assign new_n7408 = ~new_n7170 & new_n7407;
  assign new_n7409 = new_n7408 ^ new_n7173;
  assign new_n7410 = new_n7409 ^ new_n7406;
  assign new_n7411 = n95 & new_n1874;
  assign new_n7412 = new_n1864 & new_n3095;
  assign new_n7413 = new_n7412 ^ new_n7411;
  assign new_n7414 = n96 & new_n1863;
  assign new_n7415 = n94 & new_n1868;
  assign new_n7416 = new_n7415 ^ new_n7414;
  assign new_n7417 = new_n7416 ^ new_n7413;
  assign new_n7418 = new_n7417 ^ n27;
  assign new_n7419 = new_n7418 ^ new_n7410;
  assign new_n7420 = new_n7186 ^ new_n7174;
  assign new_n7421 = ~new_n7183 & new_n7420;
  assign new_n7422 = new_n7421 ^ new_n7186;
  assign new_n7423 = new_n7422 ^ new_n7419;
  assign new_n7424 = ~new_n1506 & n98;
  assign new_n7425 = new_n1501 & new_n3604;
  assign new_n7426 = new_n7425 ^ new_n7424;
  assign new_n7427 = n99 & new_n1500;
  assign new_n7428 = n97 & new_n1512;
  assign new_n7429 = new_n7428 ^ new_n7427;
  assign new_n7430 = new_n7429 ^ new_n7426;
  assign new_n7431 = new_n7430 ^ n24;
  assign new_n7432 = new_n7431 ^ new_n7423;
  assign new_n7433 = new_n7199 ^ new_n7187;
  assign new_n7434 = ~new_n7196 & new_n7433;
  assign new_n7435 = new_n7434 ^ new_n7199;
  assign new_n7436 = new_n7435 ^ new_n7432;
  assign new_n7437 = ~new_n1198 & n101;
  assign new_n7438 = new_n1193 & new_n4159;
  assign new_n7439 = new_n7438 ^ new_n7437;
  assign new_n7440 = n102 & new_n1192;
  assign new_n7441 = n100 & new_n1204;
  assign new_n7442 = new_n7441 ^ new_n7440;
  assign new_n7443 = new_n7442 ^ new_n7439;
  assign new_n7444 = new_n7443 ^ n21;
  assign new_n7445 = new_n7444 ^ new_n7436;
  assign new_n7446 = new_n7212 ^ new_n7200;
  assign new_n7447 = ~new_n7209 & new_n7446;
  assign new_n7448 = new_n7447 ^ new_n7212;
  assign new_n7449 = new_n7448 ^ new_n7445;
  assign new_n7450 = ~new_n930 & n104;
  assign new_n7451 = ~new_n4754 & new_n925;
  assign new_n7452 = new_n7451 ^ new_n7450;
  assign new_n7453 = n105 & new_n924;
  assign new_n7454 = n103 & new_n936;
  assign new_n7455 = new_n7454 ^ new_n7453;
  assign new_n7456 = new_n7455 ^ new_n7452;
  assign new_n7457 = new_n7456 ^ n18;
  assign new_n7458 = new_n7457 ^ new_n7449;
  assign new_n7459 = new_n7225 ^ new_n7213;
  assign new_n7460 = ~new_n7222 & new_n7459;
  assign new_n7461 = new_n7460 ^ new_n7225;
  assign new_n7462 = new_n7461 ^ new_n7458;
  assign new_n7463 = n107 & new_n707;
  assign new_n7464 = ~new_n5377 & new_n701;
  assign new_n7465 = new_n7464 ^ new_n7463;
  assign new_n7466 = n108 & new_n700;
  assign new_n7467 = n106 & new_n787;
  assign new_n7468 = new_n7467 ^ new_n7466;
  assign new_n7469 = new_n7468 ^ new_n7465;
  assign new_n7470 = new_n7469 ^ n15;
  assign new_n7471 = new_n7470 ^ new_n7462;
  assign new_n7472 = new_n7238 ^ new_n7226;
  assign new_n7473 = ~new_n7235 & new_n7472;
  assign new_n7474 = new_n7473 ^ new_n7238;
  assign new_n7475 = new_n7474 ^ new_n7471;
  assign new_n7476 = n110 & new_n499;
  assign new_n7477 = ~new_n506 & new_n6049;
  assign new_n7478 = new_n7477 ^ new_n7476;
  assign new_n7479 = n109 & new_n579;
  assign new_n7480 = ~new_n505 & n111;
  assign new_n7481 = new_n7480 ^ new_n7479;
  assign new_n7482 = new_n7481 ^ new_n7478;
  assign new_n7483 = new_n7482 ^ n12;
  assign new_n7484 = new_n7483 ^ new_n7475;
  assign new_n7485 = new_n7057 ^ new_n7049;
  assign new_n7486 = ~new_n7240 & new_n7485;
  assign new_n7487 = new_n7486 ^ new_n7049;
  assign new_n7488 = new_n7487 ^ new_n7484;
  assign new_n7489 = n113 & new_n354;
  assign new_n7490 = ~new_n6764 & new_n349;
  assign new_n7491 = new_n7490 ^ new_n7489;
  assign new_n7492 = n114 & new_n348;
  assign new_n7493 = n112 & new_n391;
  assign new_n7494 = new_n7493 ^ new_n7492;
  assign new_n7495 = new_n7494 ^ new_n7491;
  assign new_n7496 = new_n7495 ^ n9;
  assign new_n7497 = new_n7496 ^ new_n7488;
  assign new_n7498 = new_n7253 ^ new_n7241;
  assign new_n7499 = ~new_n7250 & new_n7498;
  assign new_n7500 = new_n7499 ^ new_n7253;
  assign new_n7501 = new_n7500 ^ new_n7497;
  assign new_n7502 = n116 & new_n218;
  assign new_n7503 = new_n6779 ^ n117;
  assign new_n7504 = ~new_n7503 & new_n208;
  assign new_n7505 = new_n7504 ^ new_n7502;
  assign new_n7506 = n117 & new_n207;
  assign new_n7507 = n115 & new_n212;
  assign new_n7508 = new_n7507 ^ new_n7506;
  assign new_n7509 = new_n7508 ^ new_n7505;
  assign new_n7510 = new_n7509 ^ n6;
  assign new_n7511 = new_n7510 ^ new_n7501;
  assign new_n7512 = new_n7267 ^ new_n7254;
  assign new_n7513 = ~new_n7264 & new_n7512;
  assign new_n7514 = new_n7513 ^ new_n7267;
  assign new_n7515 = new_n7514 ^ new_n7511;
  assign new_n7516 = n118 & new_n180;
  assign new_n7517 = n2 & n119;
  assign new_n7518 = new_n7517 ^ new_n7516;
  assign new_n7519 = new_n7518 ^ n3;
  assign new_n7520 = n119 ^ n118;
  assign new_n7521 = new_n7275 & new_n7520;
  assign new_n7522 = ~new_n7521 & new_n155;
  assign new_n7523 = new_n7522 ^ n2;
  assign new_n7524 = new_n7523 ^ n120;
  assign new_n7525 = new_n7524 ^ new_n7519;
  assign new_n7526 = ~n1 & new_n7525;
  assign new_n7527 = new_n7526 ^ new_n7524;
  assign new_n7528 = new_n7527 ^ new_n7515;
  assign new_n7529 = new_n7285 ^ new_n7268;
  assign new_n7530 = ~new_n7282 & new_n7529;
  assign new_n7531 = new_n7530 ^ new_n7285;
  assign new_n7532 = new_n7531 ^ new_n7528;
  assign new_n7533 = ~new_n6805 & n69;
  assign new_n7534 = ~new_n339 & new_n6800;
  assign new_n7535 = new_n7534 ^ new_n7533;
  assign new_n7536 = n70 & new_n6799;
  assign new_n7537 = n68 & new_n6811;
  assign new_n7538 = new_n7537 ^ new_n7536;
  assign new_n7539 = new_n7538 ^ new_n7535;
  assign new_n7540 = new_n7539 ^ n54;
  assign new_n7541 = n57 ^ n56;
  assign new_n7542 = ~new_n7541 & new_n7079;
  assign new_n7543 = new_n7542 ^ new_n7079;
  assign new_n7544 = ~new_n151 & new_n7543;
  assign new_n7545 = ~new_n7079 & n57;
  assign new_n7546 = new_n7545 ^ new_n7313;
  assign new_n7547 = new_n7541 & new_n7546;
  assign new_n7548 = n65 & new_n7547;
  assign new_n7549 = new_n7548 ^ new_n7544;
  assign new_n7550 = n67 & new_n7079;
  assign new_n7551 = new_n7550 ^ new_n7549;
  assign new_n7552 = ~new_n7079 & n56;
  assign new_n7553 = new_n7552 ^ new_n7313;
  assign new_n7554 = n66 & new_n7553;
  assign new_n7555 = new_n7554 ^ new_n7551;
  assign new_n7556 = ~new_n7080 & ~new_n7316;
  assign new_n7557 = n57 & new_n7556;
  assign new_n7558 = new_n7557 ^ n57;
  assign new_n7559 = new_n7558 ^ new_n7555;
  assign new_n7560 = new_n7559 ^ new_n7540;
  assign new_n7561 = new_n7308 ^ new_n7300;
  assign new_n7562 = ~new_n7317 & new_n7561;
  assign new_n7563 = new_n7562 ^ new_n7300;
  assign new_n7564 = new_n7563 ^ new_n7560;
  assign new_n7565 = ~new_n6110 & n72;
  assign new_n7566 = new_n534 & new_n6105;
  assign new_n7567 = new_n7566 ^ new_n7565;
  assign new_n7568 = n73 & new_n6104;
  assign new_n7569 = n71 & new_n6347;
  assign new_n7570 = new_n7569 ^ new_n7568;
  assign new_n7571 = new_n7570 ^ new_n7567;
  assign new_n7572 = new_n7571 ^ n51;
  assign new_n7573 = new_n7572 ^ new_n7564;
  assign new_n7574 = new_n7330 ^ new_n7318;
  assign new_n7575 = ~new_n7327 & new_n7574;
  assign new_n7576 = new_n7575 ^ new_n7330;
  assign new_n7577 = new_n7576 ^ new_n7573;
  assign new_n7578 = ~new_n5424 & n75;
  assign new_n7579 = ~new_n737 & new_n5419;
  assign new_n7580 = new_n7579 ^ new_n7578;
  assign new_n7581 = n76 & new_n5418;
  assign new_n7582 = n74 & new_n5648;
  assign new_n7583 = new_n7582 ^ new_n7581;
  assign new_n7584 = new_n7583 ^ new_n7580;
  assign new_n7585 = new_n7584 ^ n48;
  assign new_n7586 = new_n7585 ^ new_n7577;
  assign new_n7587 = new_n7343 ^ new_n7331;
  assign new_n7588 = ~new_n7340 & ~new_n7587;
  assign new_n7589 = new_n7588 ^ new_n7343;
  assign new_n7590 = new_n7589 ^ new_n7586;
  assign new_n7591 = ~new_n4804 & n78;
  assign new_n7592 = ~new_n982 & new_n4799;
  assign new_n7593 = new_n7592 ^ new_n7591;
  assign new_n7594 = n79 & new_n4798;
  assign new_n7595 = n77 & new_n4810;
  assign new_n7596 = new_n7595 ^ new_n7594;
  assign new_n7597 = new_n7596 ^ new_n7593;
  assign new_n7598 = new_n7597 ^ n45;
  assign new_n7599 = new_n7598 ^ new_n7590;
  assign new_n7600 = ~new_n4212 & n81;
  assign new_n7601 = new_n1263 & new_n4201;
  assign new_n7602 = new_n7601 ^ new_n7600;
  assign new_n7603 = n82 & new_n4200;
  assign new_n7604 = n80 & new_n4206;
  assign new_n7605 = new_n7604 ^ new_n7603;
  assign new_n7606 = new_n7605 ^ new_n7602;
  assign new_n7607 = new_n7606 ^ n42;
  assign new_n7608 = new_n7607 ^ new_n7599;
  assign new_n7609 = new_n7344 ^ new_n7294;
  assign new_n7610 = new_n7298 & new_n7609;
  assign new_n7611 = new_n7610 ^ new_n7297;
  assign new_n7612 = new_n7611 ^ new_n7608;
  assign new_n7613 = new_n7357 ^ new_n7345;
  assign new_n7614 = ~new_n7613 & new_n7354;
  assign new_n7615 = new_n7614 ^ new_n7357;
  assign new_n7616 = new_n7615 ^ new_n7612;
  assign new_n7617 = ~new_n3682 & n84;
  assign new_n7618 = new_n1584 & new_n3677;
  assign new_n7619 = new_n7618 ^ new_n7617;
  assign new_n7620 = n85 & new_n3676;
  assign new_n7621 = n83 & new_n3688;
  assign new_n7622 = new_n7621 ^ new_n7620;
  assign new_n7623 = new_n7622 ^ new_n7619;
  assign new_n7624 = new_n7623 ^ n39;
  assign new_n7625 = new_n7624 ^ new_n7616;
  assign new_n7626 = new_n7370 ^ new_n7358;
  assign new_n7627 = ~new_n7626 & new_n7367;
  assign new_n7628 = new_n7627 ^ new_n7370;
  assign new_n7629 = new_n7628 ^ new_n7625;
  assign new_n7630 = ~new_n3143 & n87;
  assign new_n7631 = new_n1940 & new_n3138;
  assign new_n7632 = new_n7631 ^ new_n7630;
  assign new_n7633 = n88 & new_n3137;
  assign new_n7634 = n86 & new_n3149;
  assign new_n7635 = new_n7634 ^ new_n7633;
  assign new_n7636 = new_n7635 ^ new_n7632;
  assign new_n7637 = new_n7636 ^ n36;
  assign new_n7638 = new_n7637 ^ new_n7629;
  assign new_n7639 = new_n7383 ^ new_n7371;
  assign new_n7640 = ~new_n7639 & new_n7380;
  assign new_n7641 = new_n7640 ^ new_n7383;
  assign new_n7642 = new_n7641 ^ new_n7638;
  assign new_n7643 = ~new_n2672 & n90;
  assign new_n7644 = new_n2341 & new_n2667;
  assign new_n7645 = new_n7644 ^ new_n7643;
  assign new_n7646 = n91 & new_n2666;
  assign new_n7647 = n89 & new_n2664;
  assign new_n7648 = new_n7647 ^ new_n7646;
  assign new_n7649 = new_n7648 ^ new_n7645;
  assign new_n7650 = new_n7649 ^ n33;
  assign new_n7651 = new_n7650 ^ new_n7642;
  assign new_n7652 = new_n7396 ^ new_n7384;
  assign new_n7653 = new_n7393 & new_n7652;
  assign new_n7654 = new_n7653 ^ new_n7396;
  assign new_n7655 = new_n7654 ^ new_n7651;
  assign new_n7656 = n93 & new_n2246;
  assign new_n7657 = new_n2241 & new_n2785;
  assign new_n7658 = new_n7657 ^ new_n7656;
  assign new_n7659 = n94 & new_n2240;
  assign new_n7660 = n92 & new_n2391;
  assign new_n7661 = new_n7660 ^ new_n7659;
  assign new_n7662 = new_n7661 ^ new_n7658;
  assign new_n7663 = new_n7662 ^ n30;
  assign new_n7664 = new_n7663 ^ new_n7655;
  assign new_n7665 = new_n7409 ^ new_n7397;
  assign new_n7666 = ~new_n7406 & new_n7665;
  assign new_n7667 = new_n7666 ^ new_n7409;
  assign new_n7668 = new_n7667 ^ new_n7664;
  assign new_n7669 = n96 & new_n1874;
  assign new_n7670 = new_n1864 & new_n3273;
  assign new_n7671 = new_n7670 ^ new_n7669;
  assign new_n7672 = n97 & new_n1863;
  assign new_n7673 = n95 & new_n1868;
  assign new_n7674 = new_n7673 ^ new_n7672;
  assign new_n7675 = new_n7674 ^ new_n7671;
  assign new_n7676 = new_n7675 ^ n27;
  assign new_n7677 = new_n7676 ^ new_n7668;
  assign new_n7678 = new_n7422 ^ new_n7410;
  assign new_n7679 = ~new_n7419 & new_n7678;
  assign new_n7680 = new_n7679 ^ new_n7422;
  assign new_n7681 = new_n7680 ^ new_n7677;
  assign new_n7682 = ~new_n1506 & n99;
  assign new_n7683 = new_n1501 & new_n3789;
  assign new_n7684 = new_n7683 ^ new_n7682;
  assign new_n7685 = n100 & new_n1500;
  assign new_n7686 = n98 & new_n1512;
  assign new_n7687 = new_n7686 ^ new_n7685;
  assign new_n7688 = new_n7687 ^ new_n7684;
  assign new_n7689 = new_n7688 ^ n24;
  assign new_n7690 = new_n7689 ^ new_n7681;
  assign new_n7691 = new_n7435 ^ new_n7423;
  assign new_n7692 = ~new_n7432 & new_n7691;
  assign new_n7693 = new_n7692 ^ new_n7435;
  assign new_n7694 = new_n7693 ^ new_n7690;
  assign new_n7695 = ~new_n1198 & n102;
  assign new_n7696 = new_n1193 & new_n4368;
  assign new_n7697 = new_n7696 ^ new_n7695;
  assign new_n7698 = n103 & new_n1192;
  assign new_n7699 = n101 & new_n1204;
  assign new_n7700 = new_n7699 ^ new_n7698;
  assign new_n7701 = new_n7700 ^ new_n7697;
  assign new_n7702 = new_n7701 ^ n21;
  assign new_n7703 = new_n7702 ^ new_n7694;
  assign new_n7704 = new_n7448 ^ new_n7436;
  assign new_n7705 = ~new_n7445 & new_n7704;
  assign new_n7706 = new_n7705 ^ new_n7448;
  assign new_n7707 = new_n7706 ^ new_n7703;
  assign new_n7708 = ~new_n930 & n105;
  assign new_n7709 = ~new_n4961 & new_n925;
  assign new_n7710 = new_n7709 ^ new_n7708;
  assign new_n7711 = n106 & new_n924;
  assign new_n7712 = n104 & new_n936;
  assign new_n7713 = new_n7712 ^ new_n7711;
  assign new_n7714 = new_n7713 ^ new_n7710;
  assign new_n7715 = new_n7714 ^ n18;
  assign new_n7716 = new_n7715 ^ new_n7707;
  assign new_n7717 = new_n7461 ^ new_n7449;
  assign new_n7718 = ~new_n7458 & new_n7717;
  assign new_n7719 = new_n7718 ^ new_n7461;
  assign new_n7720 = new_n7719 ^ new_n7716;
  assign new_n7721 = n108 & new_n707;
  assign new_n7722 = new_n701 & new_n5604;
  assign new_n7723 = new_n7722 ^ new_n7721;
  assign new_n7724 = n109 & new_n700;
  assign new_n7725 = n107 & new_n787;
  assign new_n7726 = new_n7725 ^ new_n7724;
  assign new_n7727 = new_n7726 ^ new_n7723;
  assign new_n7728 = new_n7727 ^ n15;
  assign new_n7729 = new_n7728 ^ new_n7720;
  assign new_n7730 = new_n7474 ^ new_n7462;
  assign new_n7731 = ~new_n7471 & new_n7730;
  assign new_n7732 = new_n7731 ^ new_n7474;
  assign new_n7733 = new_n7732 ^ new_n7729;
  assign new_n7734 = n111 & new_n499;
  assign new_n7735 = ~new_n506 & ~new_n6284;
  assign new_n7736 = new_n7735 ^ new_n7734;
  assign new_n7737 = ~new_n505 & n112;
  assign new_n7738 = n110 & new_n579;
  assign new_n7739 = new_n7738 ^ new_n7737;
  assign new_n7740 = new_n7739 ^ new_n7736;
  assign new_n7741 = new_n7740 ^ n12;
  assign new_n7742 = new_n7741 ^ new_n7733;
  assign new_n7743 = new_n7487 ^ new_n7475;
  assign new_n7744 = ~new_n7484 & new_n7743;
  assign new_n7745 = new_n7744 ^ new_n7487;
  assign new_n7746 = new_n7745 ^ new_n7742;
  assign new_n7747 = n114 & new_n354;
  assign new_n7748 = ~new_n7013 & new_n349;
  assign new_n7749 = new_n7748 ^ new_n7747;
  assign new_n7750 = n115 & new_n348;
  assign new_n7751 = n113 & new_n391;
  assign new_n7752 = new_n7751 ^ new_n7750;
  assign new_n7753 = new_n7752 ^ new_n7749;
  assign new_n7754 = new_n7753 ^ n9;
  assign new_n7755 = new_n7754 ^ new_n7746;
  assign new_n7756 = new_n7500 ^ new_n7488;
  assign new_n7757 = ~new_n7497 & new_n7756;
  assign new_n7758 = new_n7757 ^ new_n7500;
  assign new_n7759 = new_n7758 ^ new_n7755;
  assign new_n7760 = n117 & new_n218;
  assign new_n7761 = new_n7028 ^ n118;
  assign new_n7762 = ~new_n7761 & new_n208;
  assign new_n7763 = new_n7762 ^ new_n7760;
  assign new_n7764 = n118 & new_n207;
  assign new_n7765 = n116 & new_n212;
  assign new_n7766 = new_n7765 ^ new_n7764;
  assign new_n7767 = new_n7766 ^ new_n7763;
  assign new_n7768 = new_n7767 ^ n6;
  assign new_n7769 = new_n7768 ^ new_n7759;
  assign new_n7770 = new_n7514 ^ new_n7501;
  assign new_n7771 = ~new_n7511 & new_n7770;
  assign new_n7772 = new_n7771 ^ new_n7514;
  assign new_n7773 = new_n7772 ^ new_n7769;
  assign new_n7774 = n119 & new_n180;
  assign new_n7775 = n2 & n120;
  assign new_n7776 = new_n7775 ^ new_n7774;
  assign new_n7777 = new_n7776 ^ n3;
  assign new_n7778 = n120 ^ n119;
  assign new_n7779 = ~n120 & new_n7275;
  assign new_n7780 = new_n7779 ^ new_n7274;
  assign new_n7781 = ~new_n7780 & new_n7778;
  assign new_n7782 = ~new_n7781 & new_n155;
  assign new_n7783 = new_n7782 ^ n2;
  assign new_n7784 = new_n7783 ^ n121;
  assign new_n7785 = new_n7784 ^ new_n7777;
  assign new_n7786 = ~n1 & new_n7785;
  assign new_n7787 = new_n7786 ^ new_n7784;
  assign new_n7788 = new_n7787 ^ new_n7773;
  assign new_n7789 = new_n7531 ^ new_n7515;
  assign new_n7790 = ~new_n7528 & new_n7789;
  assign new_n7791 = new_n7790 ^ new_n7531;
  assign new_n7792 = new_n7791 ^ new_n7788;
  assign new_n7793 = ~new_n4804 & n79;
  assign new_n7794 = new_n1069 & new_n4799;
  assign new_n7795 = new_n7794 ^ new_n7793;
  assign new_n7796 = n80 & new_n4798;
  assign new_n7797 = n78 & new_n4810;
  assign new_n7798 = new_n7797 ^ new_n7796;
  assign new_n7799 = new_n7798 ^ new_n7795;
  assign new_n7800 = new_n7799 ^ n45;
  assign new_n7801 = new_n7611 ^ new_n7590;
  assign new_n7802 = ~new_n7801 & new_n7599;
  assign new_n7803 = new_n7802 ^ new_n7611;
  assign new_n7804 = new_n7803 ^ new_n7800;
  assign new_n7805 = ~new_n6110 & n73;
  assign new_n7806 = new_n595 & new_n6105;
  assign new_n7807 = new_n7806 ^ new_n7805;
  assign new_n7808 = n74 & new_n6104;
  assign new_n7809 = n72 & new_n6347;
  assign new_n7810 = new_n7809 ^ new_n7808;
  assign new_n7811 = new_n7810 ^ new_n7807;
  assign new_n7812 = new_n7811 ^ n51;
  assign new_n7813 = new_n7576 ^ new_n7564;
  assign new_n7814 = ~new_n7573 & new_n7813;
  assign new_n7815 = new_n7814 ^ new_n7576;
  assign new_n7816 = new_n7815 ^ new_n7812;
  assign new_n7817 = ~new_n6805 & n70;
  assign new_n7818 = ~new_n402 & new_n6800;
  assign new_n7819 = new_n7818 ^ new_n7817;
  assign new_n7820 = n71 & new_n6799;
  assign new_n7821 = n69 & new_n6811;
  assign new_n7822 = new_n7821 ^ new_n7820;
  assign new_n7823 = new_n7822 ^ new_n7819;
  assign new_n7824 = new_n7823 ^ n54;
  assign new_n7825 = new_n7563 ^ new_n7540;
  assign new_n7826 = ~new_n7560 & new_n7825;
  assign new_n7827 = new_n7826 ^ new_n7563;
  assign new_n7828 = new_n7827 ^ new_n7824;
  assign new_n7829 = ~new_n154 & new_n7541;
  assign new_n7830 = new_n7829 ^ n68;
  assign new_n7831 = new_n7079 & new_n7830;
  assign new_n7832 = n67 & new_n7553;
  assign new_n7833 = n66 & new_n7547;
  assign new_n7834 = new_n7833 ^ new_n7832;
  assign new_n7835 = ~new_n7831 & ~new_n7834;
  assign new_n7836 = new_n7835 ^ n57;
  assign new_n7837 = n58 ^ n57;
  assign new_n7838 = n65 & new_n7837;
  assign new_n7839 = new_n7838 ^ new_n7836;
  assign new_n7840 = ~new_n7555 & new_n7557;
  assign new_n7841 = ~new_n7838 & ~new_n7840;
  assign new_n7842 = new_n7841 ^ new_n7840;
  assign new_n7843 = new_n7842 ^ new_n7839;
  assign new_n7844 = new_n7843 ^ new_n7841;
  assign new_n7845 = new_n7844 ^ new_n7828;
  assign new_n7846 = new_n7845 ^ new_n7816;
  assign new_n7847 = ~new_n5424 & n76;
  assign new_n7848 = ~new_n812 & new_n5419;
  assign new_n7849 = new_n7848 ^ new_n7847;
  assign new_n7850 = n77 & new_n5418;
  assign new_n7851 = n75 & new_n5648;
  assign new_n7852 = new_n7851 ^ new_n7850;
  assign new_n7853 = new_n7852 ^ new_n7849;
  assign new_n7854 = new_n7853 ^ n48;
  assign new_n7855 = new_n7854 ^ new_n7846;
  assign new_n7856 = new_n7589 ^ new_n7577;
  assign new_n7857 = ~new_n7586 & ~new_n7856;
  assign new_n7858 = new_n7857 ^ new_n7589;
  assign new_n7859 = new_n7858 ^ new_n7855;
  assign new_n7860 = new_n7859 ^ new_n7804;
  assign new_n7861 = ~new_n4212 & n82;
  assign new_n7862 = new_n1363 & new_n4201;
  assign new_n7863 = new_n7862 ^ new_n7861;
  assign new_n7864 = n83 & new_n4200;
  assign new_n7865 = n81 & new_n4206;
  assign new_n7866 = new_n7865 ^ new_n7864;
  assign new_n7867 = new_n7866 ^ new_n7863;
  assign new_n7868 = new_n7867 ^ n42;
  assign new_n7869 = new_n7868 ^ new_n7860;
  assign new_n7870 = new_n7615 ^ new_n7607;
  assign new_n7871 = new_n7612 & new_n7870;
  assign new_n7872 = new_n7871 ^ new_n7615;
  assign new_n7873 = new_n7872 ^ new_n7869;
  assign new_n7874 = ~new_n3682 & n85;
  assign new_n7875 = new_n1694 & new_n3677;
  assign new_n7876 = new_n7875 ^ new_n7874;
  assign new_n7877 = n86 & new_n3676;
  assign new_n7878 = n84 & new_n3688;
  assign new_n7879 = new_n7878 ^ new_n7877;
  assign new_n7880 = new_n7879 ^ new_n7876;
  assign new_n7881 = new_n7880 ^ n39;
  assign new_n7882 = new_n7881 ^ new_n7873;
  assign new_n7883 = new_n7628 ^ new_n7616;
  assign new_n7884 = ~new_n7883 & new_n7625;
  assign new_n7885 = new_n7884 ^ new_n7628;
  assign new_n7886 = new_n7885 ^ new_n7882;
  assign new_n7887 = ~new_n3143 & n88;
  assign new_n7888 = new_n2063 & new_n3138;
  assign new_n7889 = new_n7888 ^ new_n7887;
  assign new_n7890 = n89 & new_n3137;
  assign new_n7891 = n87 & new_n3149;
  assign new_n7892 = new_n7891 ^ new_n7890;
  assign new_n7893 = new_n7892 ^ new_n7889;
  assign new_n7894 = new_n7893 ^ n36;
  assign new_n7895 = new_n7894 ^ new_n7886;
  assign new_n7896 = new_n7641 ^ new_n7629;
  assign new_n7897 = ~new_n7896 & new_n7638;
  assign new_n7898 = new_n7897 ^ new_n7641;
  assign new_n7899 = new_n7898 ^ new_n7895;
  assign new_n7900 = ~new_n2672 & n91;
  assign new_n7901 = new_n2481 & new_n2667;
  assign new_n7902 = new_n7901 ^ new_n7900;
  assign new_n7903 = n92 & new_n2666;
  assign new_n7904 = n90 & new_n2664;
  assign new_n7905 = new_n7904 ^ new_n7903;
  assign new_n7906 = new_n7905 ^ new_n7902;
  assign new_n7907 = new_n7906 ^ n33;
  assign new_n7908 = new_n7907 ^ new_n7899;
  assign new_n7909 = new_n7654 ^ new_n7642;
  assign new_n7910 = new_n7651 & new_n7909;
  assign new_n7911 = new_n7910 ^ new_n7654;
  assign new_n7912 = new_n7911 ^ new_n7908;
  assign new_n7913 = n94 & new_n2246;
  assign new_n7914 = new_n2241 & new_n2934;
  assign new_n7915 = new_n7914 ^ new_n7913;
  assign new_n7916 = n95 & new_n2240;
  assign new_n7917 = n93 & new_n2391;
  assign new_n7918 = new_n7917 ^ new_n7916;
  assign new_n7919 = new_n7918 ^ new_n7915;
  assign new_n7920 = new_n7919 ^ n30;
  assign new_n7921 = new_n7920 ^ new_n7912;
  assign new_n7922 = new_n7667 ^ new_n7655;
  assign new_n7923 = ~new_n7664 & new_n7922;
  assign new_n7924 = new_n7923 ^ new_n7667;
  assign new_n7925 = new_n7924 ^ new_n7921;
  assign new_n7926 = n97 & new_n1874;
  assign new_n7927 = new_n1864 & new_n3435;
  assign new_n7928 = new_n7927 ^ new_n7926;
  assign new_n7929 = n98 & new_n1863;
  assign new_n7930 = n96 & new_n1868;
  assign new_n7931 = new_n7930 ^ new_n7929;
  assign new_n7932 = new_n7931 ^ new_n7928;
  assign new_n7933 = new_n7932 ^ n27;
  assign new_n7934 = new_n7933 ^ new_n7925;
  assign new_n7935 = new_n7680 ^ new_n7668;
  assign new_n7936 = ~new_n7677 & new_n7935;
  assign new_n7937 = new_n7936 ^ new_n7680;
  assign new_n7938 = new_n7937 ^ new_n7934;
  assign new_n7939 = ~new_n1506 & n100;
  assign new_n7940 = new_n1501 & new_n3972;
  assign new_n7941 = new_n7940 ^ new_n7939;
  assign new_n7942 = n101 & new_n1500;
  assign new_n7943 = n99 & new_n1512;
  assign new_n7944 = new_n7943 ^ new_n7942;
  assign new_n7945 = new_n7944 ^ new_n7941;
  assign new_n7946 = new_n7945 ^ n24;
  assign new_n7947 = new_n7946 ^ new_n7938;
  assign new_n7948 = new_n7693 ^ new_n7681;
  assign new_n7949 = ~new_n7690 & new_n7948;
  assign new_n7950 = new_n7949 ^ new_n7693;
  assign new_n7951 = new_n7950 ^ new_n7947;
  assign new_n7952 = ~new_n1198 & n103;
  assign new_n7953 = ~new_n4556 & new_n1193;
  assign new_n7954 = new_n7953 ^ new_n7952;
  assign new_n7955 = n104 & new_n1192;
  assign new_n7956 = n102 & new_n1204;
  assign new_n7957 = new_n7956 ^ new_n7955;
  assign new_n7958 = new_n7957 ^ new_n7954;
  assign new_n7959 = new_n7958 ^ n21;
  assign new_n7960 = new_n7959 ^ new_n7951;
  assign new_n7961 = new_n7706 ^ new_n7694;
  assign new_n7962 = ~new_n7703 & new_n7961;
  assign new_n7963 = new_n7962 ^ new_n7706;
  assign new_n7964 = new_n7963 ^ new_n7960;
  assign new_n7965 = ~new_n930 & n106;
  assign new_n7966 = ~new_n5164 & new_n925;
  assign new_n7967 = new_n7966 ^ new_n7965;
  assign new_n7968 = n107 & new_n924;
  assign new_n7969 = n105 & new_n936;
  assign new_n7970 = new_n7969 ^ new_n7968;
  assign new_n7971 = new_n7970 ^ new_n7967;
  assign new_n7972 = new_n7971 ^ n18;
  assign new_n7973 = new_n7972 ^ new_n7964;
  assign new_n7974 = new_n7719 ^ new_n7707;
  assign new_n7975 = ~new_n7716 & new_n7974;
  assign new_n7976 = new_n7975 ^ new_n7719;
  assign new_n7977 = new_n7976 ^ new_n7973;
  assign new_n7978 = n109 & new_n707;
  assign new_n7979 = new_n701 & new_n5825;
  assign new_n7980 = new_n7979 ^ new_n7978;
  assign new_n7981 = n110 & new_n700;
  assign new_n7982 = n108 & new_n787;
  assign new_n7983 = new_n7982 ^ new_n7981;
  assign new_n7984 = new_n7983 ^ new_n7980;
  assign new_n7985 = new_n7984 ^ n15;
  assign new_n7986 = new_n7985 ^ new_n7977;
  assign new_n7987 = new_n7732 ^ new_n7720;
  assign new_n7988 = ~new_n7729 & new_n7987;
  assign new_n7989 = new_n7988 ^ new_n7732;
  assign new_n7990 = new_n7989 ^ new_n7986;
  assign new_n7991 = n112 & new_n499;
  assign new_n7992 = ~new_n506 & ~new_n6518;
  assign new_n7993 = new_n7992 ^ new_n7991;
  assign new_n7994 = ~new_n505 & n113;
  assign new_n7995 = n111 & new_n579;
  assign new_n7996 = new_n7995 ^ new_n7994;
  assign new_n7997 = new_n7996 ^ new_n7993;
  assign new_n7998 = new_n7997 ^ n12;
  assign new_n7999 = new_n7998 ^ new_n7990;
  assign new_n8000 = new_n7745 ^ new_n7733;
  assign new_n8001 = ~new_n7742 & new_n8000;
  assign new_n8002 = new_n8001 ^ new_n7745;
  assign new_n8003 = new_n8002 ^ new_n7999;
  assign new_n8004 = n115 & new_n354;
  assign new_n8005 = ~new_n7256 & new_n349;
  assign new_n8006 = new_n8005 ^ new_n8004;
  assign new_n8007 = n116 & new_n348;
  assign new_n8008 = n114 & new_n391;
  assign new_n8009 = new_n8008 ^ new_n8007;
  assign new_n8010 = new_n8009 ^ new_n8006;
  assign new_n8011 = new_n8010 ^ n9;
  assign new_n8012 = new_n8011 ^ new_n8003;
  assign new_n8013 = new_n7758 ^ new_n7746;
  assign new_n8014 = ~new_n7755 & new_n8013;
  assign new_n8015 = new_n8014 ^ new_n7758;
  assign new_n8016 = new_n8015 ^ new_n8012;
  assign new_n8017 = n118 & new_n218;
  assign new_n8018 = new_n7275 ^ n118;
  assign new_n8019 = new_n8018 ^ new_n7520;
  assign new_n8020 = ~new_n8019 & new_n208;
  assign new_n8021 = new_n8020 ^ new_n8017;
  assign new_n8022 = n119 & new_n207;
  assign new_n8023 = n117 & new_n212;
  assign new_n8024 = new_n8023 ^ new_n8022;
  assign new_n8025 = new_n8024 ^ new_n8021;
  assign new_n8026 = new_n8025 ^ n6;
  assign new_n8027 = new_n8026 ^ new_n8016;
  assign new_n8028 = new_n7772 ^ new_n7759;
  assign new_n8029 = ~new_n7769 & new_n8028;
  assign new_n8030 = new_n8029 ^ new_n7772;
  assign new_n8031 = new_n8030 ^ new_n8027;
  assign new_n8032 = n120 & new_n180;
  assign new_n8033 = n2 & n121;
  assign new_n8034 = new_n8033 ^ new_n8032;
  assign new_n8035 = new_n8034 ^ n3;
  assign new_n8036 = ~n119 & ~n121;
  assign new_n8037 = ~n118 & ~n120;
  assign new_n8038 = ~new_n8036 & ~new_n8037;
  assign new_n8039 = ~new_n8038 & new_n8018;
  assign new_n8040 = ~n118 & new_n8036;
  assign new_n8041 = ~n120 & n121;
  assign new_n8042 = n119 & new_n8041;
  assign new_n8043 = new_n8042 ^ n120;
  assign new_n8044 = ~new_n8040 & new_n8043;
  assign new_n8045 = ~new_n8039 & new_n8044;
  assign new_n8046 = new_n8045 ^ n121;
  assign new_n8047 = ~new_n8046 & new_n155;
  assign new_n8048 = new_n8047 ^ n2;
  assign new_n8049 = new_n8048 ^ n122;
  assign new_n8050 = new_n8049 ^ new_n8035;
  assign new_n8051 = ~n1 & new_n8050;
  assign new_n8052 = new_n8051 ^ new_n8049;
  assign new_n8053 = new_n8052 ^ new_n8031;
  assign new_n8054 = new_n7791 ^ new_n7773;
  assign new_n8055 = ~new_n7788 & new_n8054;
  assign new_n8056 = new_n8055 ^ new_n7791;
  assign new_n8057 = new_n8056 ^ new_n8053;
  assign new_n8058 = n57 & n58;
  assign new_n8059 = new_n8058 ^ n59;
  assign new_n8060 = ~n65 & new_n8059;
  assign new_n8061 = n66 ^ n58;
  assign new_n8062 = ~new_n8061 & new_n7837;
  assign new_n8063 = new_n8062 ^ n57;
  assign new_n8064 = new_n8063 ^ n59;
  assign new_n8065 = new_n8064 ^ new_n8060;
  assign new_n8066 = ~new_n7836 & ~new_n7841;
  assign new_n8067 = new_n8066 ^ new_n8065;
  assign new_n8068 = n68 & new_n7553;
  assign new_n8069 = ~new_n304 & new_n7543;
  assign new_n8070 = new_n8069 ^ new_n8068;
  assign new_n8071 = n69 & new_n7542;
  assign new_n8072 = n67 & new_n7547;
  assign new_n8073 = new_n8072 ^ new_n8071;
  assign new_n8074 = new_n8073 ^ new_n8070;
  assign new_n8075 = new_n8074 ^ n57;
  assign new_n8076 = new_n8075 ^ new_n8067;
  assign new_n8077 = ~new_n6805 & n71;
  assign new_n8078 = ~new_n459 & new_n6800;
  assign new_n8079 = new_n8078 ^ new_n8077;
  assign new_n8080 = n72 & new_n6799;
  assign new_n8081 = n70 & new_n6811;
  assign new_n8082 = new_n8081 ^ new_n8080;
  assign new_n8083 = new_n8082 ^ new_n8079;
  assign new_n8084 = new_n8083 ^ n54;
  assign new_n8085 = new_n8084 ^ new_n8076;
  assign new_n8086 = new_n7844 ^ new_n7824;
  assign new_n8087 = new_n7828 & new_n8086;
  assign new_n8088 = new_n8087 ^ new_n7827;
  assign new_n8089 = new_n8088 ^ new_n8085;
  assign new_n8090 = ~new_n6110 & n74;
  assign new_n8091 = new_n660 & new_n6105;
  assign new_n8092 = new_n8091 ^ new_n8090;
  assign new_n8093 = n75 & new_n6104;
  assign new_n8094 = n73 & new_n6347;
  assign new_n8095 = new_n8094 ^ new_n8093;
  assign new_n8096 = new_n8095 ^ new_n8092;
  assign new_n8097 = new_n8096 ^ n51;
  assign new_n8098 = new_n8097 ^ new_n8089;
  assign new_n8099 = new_n7845 ^ new_n7812;
  assign new_n8100 = new_n7816 & new_n8099;
  assign new_n8101 = new_n8100 ^ new_n7815;
  assign new_n8102 = new_n8101 ^ new_n8098;
  assign new_n8103 = ~new_n5424 & n77;
  assign new_n8104 = ~new_n891 & new_n5419;
  assign new_n8105 = new_n8104 ^ new_n8103;
  assign new_n8106 = n78 & new_n5418;
  assign new_n8107 = n76 & new_n5648;
  assign new_n8108 = new_n8107 ^ new_n8106;
  assign new_n8109 = new_n8108 ^ new_n8105;
  assign new_n8110 = new_n8109 ^ n48;
  assign new_n8111 = new_n8110 ^ new_n8102;
  assign new_n8112 = new_n7858 ^ new_n7846;
  assign new_n8113 = new_n7855 & new_n8112;
  assign new_n8114 = new_n8113 ^ new_n7858;
  assign new_n8115 = new_n8114 ^ new_n8111;
  assign new_n8116 = ~new_n4804 & n80;
  assign new_n8117 = new_n1161 & new_n4799;
  assign new_n8118 = new_n8117 ^ new_n8116;
  assign new_n8119 = n79 & new_n4810;
  assign new_n8120 = n81 & new_n4798;
  assign new_n8121 = new_n8120 ^ new_n8119;
  assign new_n8122 = new_n8121 ^ new_n8118;
  assign new_n8123 = new_n8122 ^ n45;
  assign new_n8124 = new_n8123 ^ new_n8115;
  assign new_n8125 = new_n7859 ^ new_n7800;
  assign new_n8126 = ~new_n8125 & new_n7804;
  assign new_n8127 = new_n8126 ^ new_n7803;
  assign new_n8128 = new_n8127 ^ new_n8124;
  assign new_n8129 = ~new_n4212 & n83;
  assign new_n8130 = new_n1468 & new_n4201;
  assign new_n8131 = new_n8130 ^ new_n8129;
  assign new_n8132 = n84 & new_n4200;
  assign new_n8133 = n82 & new_n4206;
  assign new_n8134 = new_n8133 ^ new_n8132;
  assign new_n8135 = new_n8134 ^ new_n8131;
  assign new_n8136 = new_n8135 ^ n42;
  assign new_n8137 = new_n8136 ^ new_n8128;
  assign new_n8138 = new_n7872 ^ new_n7860;
  assign new_n8139 = ~new_n7869 & new_n8138;
  assign new_n8140 = new_n8139 ^ new_n7872;
  assign new_n8141 = new_n8140 ^ new_n8137;
  assign new_n8142 = ~new_n3682 & n86;
  assign new_n8143 = new_n1811 & new_n3677;
  assign new_n8144 = new_n8143 ^ new_n8142;
  assign new_n8145 = n87 & new_n3676;
  assign new_n8146 = n85 & new_n3688;
  assign new_n8147 = new_n8146 ^ new_n8145;
  assign new_n8148 = new_n8147 ^ new_n8144;
  assign new_n8149 = new_n8148 ^ n39;
  assign new_n8150 = new_n8149 ^ new_n8141;
  assign new_n8151 = new_n7885 ^ new_n7873;
  assign new_n8152 = ~new_n7882 & new_n8151;
  assign new_n8153 = new_n8152 ^ new_n7885;
  assign new_n8154 = new_n8153 ^ new_n8150;
  assign new_n8155 = ~new_n3143 & n89;
  assign new_n8156 = new_n2193 & new_n3138;
  assign new_n8157 = new_n8156 ^ new_n8155;
  assign new_n8158 = n90 & new_n3137;
  assign new_n8159 = n88 & new_n3149;
  assign new_n8160 = new_n8159 ^ new_n8158;
  assign new_n8161 = new_n8160 ^ new_n8157;
  assign new_n8162 = new_n8161 ^ n36;
  assign new_n8163 = new_n8162 ^ new_n8154;
  assign new_n8164 = new_n7898 ^ new_n7886;
  assign new_n8165 = ~new_n7895 & new_n8164;
  assign new_n8166 = new_n8165 ^ new_n7898;
  assign new_n8167 = new_n8166 ^ new_n8163;
  assign new_n8168 = ~new_n2672 & n92;
  assign new_n8169 = new_n2628 & new_n2667;
  assign new_n8170 = new_n8169 ^ new_n8168;
  assign new_n8171 = n93 & new_n2666;
  assign new_n8172 = n91 & new_n2664;
  assign new_n8173 = new_n8172 ^ new_n8171;
  assign new_n8174 = new_n8173 ^ new_n8170;
  assign new_n8175 = new_n8174 ^ n33;
  assign new_n8176 = new_n8175 ^ new_n8167;
  assign new_n8177 = new_n7911 ^ new_n7899;
  assign new_n8178 = ~new_n7908 & ~new_n8177;
  assign new_n8179 = new_n8178 ^ new_n7911;
  assign new_n8180 = new_n8179 ^ new_n8176;
  assign new_n8181 = n95 & new_n2246;
  assign new_n8182 = new_n2241 & new_n3095;
  assign new_n8183 = new_n8182 ^ new_n8181;
  assign new_n8184 = n96 & new_n2240;
  assign new_n8185 = n94 & new_n2391;
  assign new_n8186 = new_n8185 ^ new_n8184;
  assign new_n8187 = new_n8186 ^ new_n8183;
  assign new_n8188 = new_n8187 ^ n30;
  assign new_n8189 = new_n8188 ^ new_n8180;
  assign new_n8190 = new_n7924 ^ new_n7912;
  assign new_n8191 = ~new_n8190 & new_n7921;
  assign new_n8192 = new_n8191 ^ new_n7924;
  assign new_n8193 = new_n8192 ^ new_n8189;
  assign new_n8194 = n98 & new_n1874;
  assign new_n8195 = new_n1864 & new_n3604;
  assign new_n8196 = new_n8195 ^ new_n8194;
  assign new_n8197 = n99 & new_n1863;
  assign new_n8198 = n97 & new_n1868;
  assign new_n8199 = new_n8198 ^ new_n8197;
  assign new_n8200 = new_n8199 ^ new_n8196;
  assign new_n8201 = new_n8200 ^ n27;
  assign new_n8202 = new_n8201 ^ new_n8193;
  assign new_n8203 = new_n7937 ^ new_n7925;
  assign new_n8204 = ~new_n8203 & new_n7934;
  assign new_n8205 = new_n8204 ^ new_n7937;
  assign new_n8206 = new_n8205 ^ new_n8202;
  assign new_n8207 = ~new_n1506 & n101;
  assign new_n8208 = new_n1501 & new_n4159;
  assign new_n8209 = new_n8208 ^ new_n8207;
  assign new_n8210 = n102 & new_n1500;
  assign new_n8211 = n100 & new_n1512;
  assign new_n8212 = new_n8211 ^ new_n8210;
  assign new_n8213 = new_n8212 ^ new_n8209;
  assign new_n8214 = new_n8213 ^ n24;
  assign new_n8215 = new_n8214 ^ new_n8206;
  assign new_n8216 = new_n7950 ^ new_n7938;
  assign new_n8217 = ~new_n8216 & new_n7947;
  assign new_n8218 = new_n8217 ^ new_n7950;
  assign new_n8219 = new_n8218 ^ new_n8215;
  assign new_n8220 = ~new_n1198 & n104;
  assign new_n8221 = ~new_n4754 & new_n1193;
  assign new_n8222 = new_n8221 ^ new_n8220;
  assign new_n8223 = n105 & new_n1192;
  assign new_n8224 = n103 & new_n1204;
  assign new_n8225 = new_n8224 ^ new_n8223;
  assign new_n8226 = new_n8225 ^ new_n8222;
  assign new_n8227 = new_n8226 ^ n21;
  assign new_n8228 = new_n8227 ^ new_n8219;
  assign new_n8229 = new_n7963 ^ new_n7951;
  assign new_n8230 = ~new_n8229 & new_n7960;
  assign new_n8231 = new_n8230 ^ new_n7963;
  assign new_n8232 = new_n8231 ^ new_n8228;
  assign new_n8233 = ~new_n930 & n107;
  assign new_n8234 = ~new_n5377 & new_n925;
  assign new_n8235 = new_n8234 ^ new_n8233;
  assign new_n8236 = n108 & new_n924;
  assign new_n8237 = n106 & new_n936;
  assign new_n8238 = new_n8237 ^ new_n8236;
  assign new_n8239 = new_n8238 ^ new_n8235;
  assign new_n8240 = new_n8239 ^ n18;
  assign new_n8241 = new_n8240 ^ new_n8232;
  assign new_n8242 = new_n7976 ^ new_n7964;
  assign new_n8243 = ~new_n8242 & new_n7973;
  assign new_n8244 = new_n8243 ^ new_n7976;
  assign new_n8245 = new_n8244 ^ new_n8241;
  assign new_n8246 = n110 & new_n707;
  assign new_n8247 = new_n701 & new_n6049;
  assign new_n8248 = new_n8247 ^ new_n8246;
  assign new_n8249 = n111 & new_n700;
  assign new_n8250 = n109 & new_n787;
  assign new_n8251 = new_n8250 ^ new_n8249;
  assign new_n8252 = new_n8251 ^ new_n8248;
  assign new_n8253 = new_n8252 ^ n15;
  assign new_n8254 = new_n8253 ^ new_n8245;
  assign new_n8255 = new_n7989 ^ new_n7977;
  assign new_n8256 = ~new_n8255 & new_n7986;
  assign new_n8257 = new_n8256 ^ new_n7989;
  assign new_n8258 = new_n8257 ^ new_n8254;
  assign new_n8259 = n113 & new_n499;
  assign new_n8260 = ~new_n506 & ~new_n6764;
  assign new_n8261 = new_n8260 ^ new_n8259;
  assign new_n8262 = ~new_n505 & n114;
  assign new_n8263 = n112 & new_n579;
  assign new_n8264 = new_n8263 ^ new_n8262;
  assign new_n8265 = new_n8264 ^ new_n8261;
  assign new_n8266 = new_n8265 ^ n12;
  assign new_n8267 = new_n8266 ^ new_n8258;
  assign new_n8268 = new_n8002 ^ new_n7990;
  assign new_n8269 = ~new_n8268 & new_n7999;
  assign new_n8270 = new_n8269 ^ new_n8002;
  assign new_n8271 = new_n8270 ^ new_n8267;
  assign new_n8272 = n116 & new_n354;
  assign new_n8273 = ~new_n7503 & new_n349;
  assign new_n8274 = new_n8273 ^ new_n8272;
  assign new_n8275 = n117 & new_n348;
  assign new_n8276 = n115 & new_n391;
  assign new_n8277 = new_n8276 ^ new_n8275;
  assign new_n8278 = new_n8277 ^ new_n8274;
  assign new_n8279 = new_n8278 ^ n9;
  assign new_n8280 = new_n8279 ^ new_n8271;
  assign new_n8281 = new_n8015 ^ new_n8003;
  assign new_n8282 = ~new_n8281 & new_n8012;
  assign new_n8283 = new_n8282 ^ new_n8015;
  assign new_n8284 = new_n8283 ^ new_n8280;
  assign new_n8285 = n119 & new_n218;
  assign new_n8286 = new_n7521 ^ n120;
  assign new_n8287 = new_n208 & new_n8286;
  assign new_n8288 = new_n8287 ^ new_n8285;
  assign new_n8289 = n120 & new_n207;
  assign new_n8290 = n118 & new_n212;
  assign new_n8291 = new_n8290 ^ new_n8289;
  assign new_n8292 = new_n8291 ^ new_n8288;
  assign new_n8293 = new_n8292 ^ n6;
  assign new_n8294 = n121 & new_n180;
  assign new_n8295 = n2 & n122;
  assign new_n8296 = new_n8295 ^ new_n8294;
  assign new_n8297 = new_n8296 ^ n3;
  assign new_n8298 = n121 & new_n8045;
  assign new_n8299 = new_n8298 ^ new_n8046;
  assign new_n8300 = n122 & new_n8299;
  assign new_n8301 = ~n122 & ~new_n8298;
  assign new_n8302 = new_n8301 ^ new_n8300;
  assign new_n8303 = new_n155 & new_n8302;
  assign new_n8304 = new_n8303 ^ n2;
  assign new_n8305 = new_n8304 ^ n123;
  assign new_n8306 = new_n8305 ^ new_n8297;
  assign new_n8307 = ~n1 & new_n8306;
  assign new_n8308 = new_n8307 ^ new_n8305;
  assign new_n8309 = new_n8308 ^ new_n8293;
  assign new_n8310 = new_n8309 ^ new_n8284;
  assign new_n8311 = new_n8030 ^ new_n8016;
  assign new_n8312 = ~new_n8311 & new_n8027;
  assign new_n8313 = new_n8312 ^ new_n8030;
  assign new_n8314 = new_n8313 ^ new_n8310;
  assign new_n8315 = new_n8056 ^ new_n8031;
  assign new_n8316 = ~new_n8315 & new_n8053;
  assign new_n8317 = new_n8316 ^ new_n8056;
  assign new_n8318 = new_n8317 ^ new_n8314;
  assign new_n8319 = ~new_n5424 & n78;
  assign new_n8320 = ~new_n982 & new_n5419;
  assign new_n8321 = new_n8320 ^ new_n8319;
  assign new_n8322 = n79 & new_n5418;
  assign new_n8323 = n77 & new_n5648;
  assign new_n8324 = new_n8323 ^ new_n8322;
  assign new_n8325 = new_n8324 ^ new_n8321;
  assign new_n8326 = new_n8325 ^ n48;
  assign new_n8327 = new_n8114 ^ new_n8102;
  assign new_n8328 = ~new_n8111 & ~new_n8327;
  assign new_n8329 = new_n8328 ^ new_n8114;
  assign new_n8330 = new_n8329 ^ new_n8326;
  assign new_n8331 = ~new_n6110 & n75;
  assign new_n8332 = ~new_n737 & new_n6105;
  assign new_n8333 = new_n8332 ^ new_n8331;
  assign new_n8334 = n76 & new_n6104;
  assign new_n8335 = n74 & new_n6347;
  assign new_n8336 = new_n8335 ^ new_n8334;
  assign new_n8337 = new_n8336 ^ new_n8333;
  assign new_n8338 = new_n8337 ^ n51;
  assign new_n8339 = new_n8101 ^ new_n8089;
  assign new_n8340 = ~new_n8098 & new_n8339;
  assign new_n8341 = new_n8340 ^ new_n8101;
  assign new_n8342 = new_n8341 ^ new_n8338;
  assign new_n8343 = n60 ^ n59;
  assign new_n8344 = ~new_n8343 & new_n7837;
  assign new_n8345 = new_n8344 ^ new_n7837;
  assign new_n8346 = ~new_n151 & new_n8345;
  assign new_n8347 = ~new_n7837 & n60;
  assign new_n8348 = new_n8347 ^ new_n8058;
  assign new_n8349 = new_n8343 & new_n8348;
  assign new_n8350 = n65 & new_n8349;
  assign new_n8351 = new_n8350 ^ new_n8346;
  assign new_n8352 = n67 & new_n7837;
  assign new_n8353 = new_n8352 ^ new_n8351;
  assign new_n8354 = ~new_n7837 & n59;
  assign new_n8355 = new_n8354 ^ new_n8058;
  assign new_n8356 = n66 & new_n8355;
  assign new_n8357 = new_n8356 ^ new_n8353;
  assign new_n8358 = ~new_n7838 & ~new_n8065;
  assign new_n8359 = n60 & new_n8358;
  assign new_n8360 = new_n8359 ^ n60;
  assign new_n8361 = new_n8360 ^ new_n8357;
  assign new_n8362 = new_n8075 ^ new_n8065;
  assign new_n8363 = ~new_n8362 & new_n8067;
  assign new_n8364 = new_n8363 ^ new_n8066;
  assign new_n8365 = new_n8364 ^ new_n8361;
  assign new_n8366 = n69 & new_n7553;
  assign new_n8367 = ~new_n339 & new_n7543;
  assign new_n8368 = new_n8367 ^ new_n8366;
  assign new_n8369 = n70 & new_n7542;
  assign new_n8370 = n68 & new_n7547;
  assign new_n8371 = new_n8370 ^ new_n8369;
  assign new_n8372 = new_n8371 ^ new_n8368;
  assign new_n8373 = new_n8372 ^ n57;
  assign new_n8374 = new_n8373 ^ new_n8365;
  assign new_n8375 = ~new_n6805 & n72;
  assign new_n8376 = new_n534 & new_n6800;
  assign new_n8377 = new_n8376 ^ new_n8375;
  assign new_n8378 = n73 & new_n6799;
  assign new_n8379 = n71 & new_n6811;
  assign new_n8380 = new_n8379 ^ new_n8378;
  assign new_n8381 = new_n8380 ^ new_n8377;
  assign new_n8382 = new_n8381 ^ n54;
  assign new_n8383 = new_n8382 ^ new_n8374;
  assign new_n8384 = new_n8088 ^ new_n8076;
  assign new_n8385 = ~new_n8085 & new_n8384;
  assign new_n8386 = new_n8385 ^ new_n8088;
  assign new_n8387 = new_n8386 ^ new_n8383;
  assign new_n8388 = new_n8387 ^ new_n8342;
  assign new_n8389 = new_n8388 ^ new_n8330;
  assign new_n8390 = ~new_n4804 & n81;
  assign new_n8391 = new_n1263 & new_n4799;
  assign new_n8392 = new_n8391 ^ new_n8390;
  assign new_n8393 = n82 & new_n4798;
  assign new_n8394 = n80 & new_n4810;
  assign new_n8395 = new_n8394 ^ new_n8393;
  assign new_n8396 = new_n8395 ^ new_n8392;
  assign new_n8397 = new_n8396 ^ n45;
  assign new_n8398 = new_n8397 ^ new_n8389;
  assign new_n8399 = new_n8127 ^ new_n8115;
  assign new_n8400 = ~new_n8399 & new_n8124;
  assign new_n8401 = new_n8400 ^ new_n8127;
  assign new_n8402 = new_n8401 ^ new_n8398;
  assign new_n8403 = ~new_n4212 & n84;
  assign new_n8404 = new_n1584 & new_n4201;
  assign new_n8405 = new_n8404 ^ new_n8403;
  assign new_n8406 = n85 & new_n4200;
  assign new_n8407 = n83 & new_n4206;
  assign new_n8408 = new_n8407 ^ new_n8406;
  assign new_n8409 = new_n8408 ^ new_n8405;
  assign new_n8410 = new_n8409 ^ n42;
  assign new_n8411 = new_n8410 ^ new_n8402;
  assign new_n8412 = new_n8140 ^ new_n8128;
  assign new_n8413 = ~new_n8412 & new_n8137;
  assign new_n8414 = new_n8413 ^ new_n8140;
  assign new_n8415 = new_n8414 ^ new_n8411;
  assign new_n8416 = ~new_n3682 & n87;
  assign new_n8417 = new_n1940 & new_n3677;
  assign new_n8418 = new_n8417 ^ new_n8416;
  assign new_n8419 = n88 & new_n3676;
  assign new_n8420 = n86 & new_n3688;
  assign new_n8421 = new_n8420 ^ new_n8419;
  assign new_n8422 = new_n8421 ^ new_n8418;
  assign new_n8423 = new_n8422 ^ n39;
  assign new_n8424 = new_n8423 ^ new_n8415;
  assign new_n8425 = new_n8153 ^ new_n8141;
  assign new_n8426 = ~new_n8425 & new_n8150;
  assign new_n8427 = new_n8426 ^ new_n8153;
  assign new_n8428 = new_n8427 ^ new_n8424;
  assign new_n8429 = ~new_n3143 & n90;
  assign new_n8430 = new_n2341 & new_n3138;
  assign new_n8431 = new_n8430 ^ new_n8429;
  assign new_n8432 = n91 & new_n3137;
  assign new_n8433 = n89 & new_n3149;
  assign new_n8434 = new_n8433 ^ new_n8432;
  assign new_n8435 = new_n8434 ^ new_n8431;
  assign new_n8436 = new_n8435 ^ n36;
  assign new_n8437 = new_n8436 ^ new_n8428;
  assign new_n8438 = new_n8166 ^ new_n8154;
  assign new_n8439 = ~new_n8438 & new_n8163;
  assign new_n8440 = new_n8439 ^ new_n8166;
  assign new_n8441 = new_n8440 ^ new_n8437;
  assign new_n8442 = ~new_n2672 & n93;
  assign new_n8443 = new_n2667 & new_n2785;
  assign new_n8444 = new_n8443 ^ new_n8442;
  assign new_n8445 = n94 & new_n2666;
  assign new_n8446 = n92 & new_n2664;
  assign new_n8447 = new_n8446 ^ new_n8445;
  assign new_n8448 = new_n8447 ^ new_n8444;
  assign new_n8449 = new_n8448 ^ n33;
  assign new_n8450 = new_n8449 ^ new_n8441;
  assign new_n8451 = new_n8179 ^ new_n8167;
  assign new_n8452 = new_n8176 & new_n8451;
  assign new_n8453 = new_n8452 ^ new_n8179;
  assign new_n8454 = new_n8453 ^ new_n8450;
  assign new_n8455 = n96 & new_n2246;
  assign new_n8456 = new_n2241 & new_n3273;
  assign new_n8457 = new_n8456 ^ new_n8455;
  assign new_n8458 = n97 & new_n2240;
  assign new_n8459 = n95 & new_n2391;
  assign new_n8460 = new_n8459 ^ new_n8458;
  assign new_n8461 = new_n8460 ^ new_n8457;
  assign new_n8462 = new_n8461 ^ n30;
  assign new_n8463 = new_n8462 ^ new_n8454;
  assign new_n8464 = new_n8192 ^ new_n8188;
  assign new_n8465 = ~new_n8464 & new_n8189;
  assign new_n8466 = new_n8465 ^ new_n8180;
  assign new_n8467 = new_n8466 ^ new_n8463;
  assign new_n8468 = n99 & new_n1874;
  assign new_n8469 = new_n1864 & new_n3789;
  assign new_n8470 = new_n8469 ^ new_n8468;
  assign new_n8471 = n100 & new_n1863;
  assign new_n8472 = n98 & new_n1868;
  assign new_n8473 = new_n8472 ^ new_n8471;
  assign new_n8474 = new_n8473 ^ new_n8470;
  assign new_n8475 = new_n8474 ^ n27;
  assign new_n8476 = new_n8475 ^ new_n8467;
  assign new_n8477 = new_n8205 ^ new_n8193;
  assign new_n8478 = ~new_n8202 & new_n8477;
  assign new_n8479 = new_n8478 ^ new_n8205;
  assign new_n8480 = new_n8479 ^ new_n8476;
  assign new_n8481 = ~new_n1506 & n102;
  assign new_n8482 = new_n1501 & new_n4368;
  assign new_n8483 = new_n8482 ^ new_n8481;
  assign new_n8484 = n103 & new_n1500;
  assign new_n8485 = n101 & new_n1512;
  assign new_n8486 = new_n8485 ^ new_n8484;
  assign new_n8487 = new_n8486 ^ new_n8483;
  assign new_n8488 = new_n8487 ^ n24;
  assign new_n8489 = new_n8488 ^ new_n8480;
  assign new_n8490 = new_n8218 ^ new_n8206;
  assign new_n8491 = ~new_n8215 & new_n8490;
  assign new_n8492 = new_n8491 ^ new_n8218;
  assign new_n8493 = new_n8492 ^ new_n8489;
  assign new_n8494 = ~new_n1198 & n105;
  assign new_n8495 = ~new_n4961 & new_n1193;
  assign new_n8496 = new_n8495 ^ new_n8494;
  assign new_n8497 = n106 & new_n1192;
  assign new_n8498 = n104 & new_n1204;
  assign new_n8499 = new_n8498 ^ new_n8497;
  assign new_n8500 = new_n8499 ^ new_n8496;
  assign new_n8501 = new_n8500 ^ n21;
  assign new_n8502 = new_n8501 ^ new_n8493;
  assign new_n8503 = new_n8231 ^ new_n8219;
  assign new_n8504 = ~new_n8228 & new_n8503;
  assign new_n8505 = new_n8504 ^ new_n8231;
  assign new_n8506 = new_n8505 ^ new_n8502;
  assign new_n8507 = ~new_n930 & n108;
  assign new_n8508 = new_n925 & new_n5604;
  assign new_n8509 = new_n8508 ^ new_n8507;
  assign new_n8510 = n109 & new_n924;
  assign new_n8511 = n107 & new_n936;
  assign new_n8512 = new_n8511 ^ new_n8510;
  assign new_n8513 = new_n8512 ^ new_n8509;
  assign new_n8514 = new_n8513 ^ n18;
  assign new_n8515 = new_n8514 ^ new_n8506;
  assign new_n8516 = new_n8244 ^ new_n8232;
  assign new_n8517 = ~new_n8241 & new_n8516;
  assign new_n8518 = new_n8517 ^ new_n8244;
  assign new_n8519 = new_n8518 ^ new_n8515;
  assign new_n8520 = n111 & new_n707;
  assign new_n8521 = ~new_n6284 & new_n701;
  assign new_n8522 = new_n8521 ^ new_n8520;
  assign new_n8523 = n112 & new_n700;
  assign new_n8524 = n110 & new_n787;
  assign new_n8525 = new_n8524 ^ new_n8523;
  assign new_n8526 = new_n8525 ^ new_n8522;
  assign new_n8527 = new_n8526 ^ n15;
  assign new_n8528 = new_n8527 ^ new_n8519;
  assign new_n8529 = new_n8257 ^ new_n8245;
  assign new_n8530 = ~new_n8254 & new_n8529;
  assign new_n8531 = new_n8530 ^ new_n8257;
  assign new_n8532 = new_n8531 ^ new_n8528;
  assign new_n8533 = n114 & new_n499;
  assign new_n8534 = ~new_n506 & ~new_n7013;
  assign new_n8535 = new_n8534 ^ new_n8533;
  assign new_n8536 = ~new_n505 & n115;
  assign new_n8537 = n113 & new_n579;
  assign new_n8538 = new_n8537 ^ new_n8536;
  assign new_n8539 = new_n8538 ^ new_n8535;
  assign new_n8540 = new_n8539 ^ n12;
  assign new_n8541 = new_n8540 ^ new_n8532;
  assign new_n8542 = new_n8270 ^ new_n8258;
  assign new_n8543 = ~new_n8267 & new_n8542;
  assign new_n8544 = new_n8543 ^ new_n8270;
  assign new_n8545 = new_n8544 ^ new_n8541;
  assign new_n8546 = n117 & new_n354;
  assign new_n8547 = ~new_n7761 & new_n349;
  assign new_n8548 = new_n8547 ^ new_n8546;
  assign new_n8549 = n118 & new_n348;
  assign new_n8550 = n116 & new_n391;
  assign new_n8551 = new_n8550 ^ new_n8549;
  assign new_n8552 = new_n8551 ^ new_n8548;
  assign new_n8553 = new_n8552 ^ n9;
  assign new_n8554 = new_n8553 ^ new_n8545;
  assign new_n8555 = new_n8283 ^ new_n8271;
  assign new_n8556 = ~new_n8280 & new_n8555;
  assign new_n8557 = new_n8556 ^ new_n8283;
  assign new_n8558 = new_n8557 ^ new_n8554;
  assign new_n8559 = n120 & new_n218;
  assign new_n8560 = new_n7781 ^ n121;
  assign new_n8561 = new_n208 & new_n8560;
  assign new_n8562 = new_n8561 ^ new_n8559;
  assign new_n8563 = n121 & new_n207;
  assign new_n8564 = n119 & new_n212;
  assign new_n8565 = new_n8564 ^ new_n8563;
  assign new_n8566 = new_n8565 ^ new_n8562;
  assign new_n8567 = new_n8566 ^ n6;
  assign new_n8568 = n122 & new_n180;
  assign new_n8569 = n2 & n123;
  assign new_n8570 = new_n8569 ^ new_n8568;
  assign new_n8571 = new_n8570 ^ n3;
  assign new_n8572 = ~new_n8301 & n123;
  assign new_n8573 = ~n123 & ~new_n8300;
  assign new_n8574 = new_n8573 ^ new_n8572;
  assign new_n8575 = new_n155 & new_n8574;
  assign new_n8576 = new_n8575 ^ n2;
  assign new_n8577 = new_n8576 ^ n124;
  assign new_n8578 = new_n8577 ^ new_n8571;
  assign new_n8579 = ~n1 & new_n8578;
  assign new_n8580 = new_n8579 ^ new_n8577;
  assign new_n8581 = new_n8580 ^ new_n8567;
  assign new_n8582 = new_n8581 ^ new_n8558;
  assign new_n8583 = new_n8293 & new_n8308;
  assign new_n8584 = new_n8583 ^ new_n8309;
  assign new_n8585 = ~new_n8284 & ~new_n8584;
  assign new_n8586 = ~new_n8313 & new_n8585;
  assign new_n8587 = new_n8284 & new_n8583;
  assign new_n8588 = new_n8313 & new_n8587;
  assign new_n8589 = new_n8588 ^ new_n8586;
  assign new_n8590 = new_n8587 ^ new_n8309;
  assign new_n8591 = new_n8590 ^ new_n8585;
  assign new_n8592 = new_n8591 ^ new_n8284;
  assign new_n8593 = ~new_n8313 & new_n8592;
  assign new_n8594 = ~new_n8585 & ~new_n8593;
  assign new_n8595 = new_n8594 ^ new_n8314;
  assign new_n8596 = new_n8595 ^ new_n8589;
  assign new_n8597 = new_n8596 ^ new_n8594;
  assign new_n8598 = new_n8317 & new_n8597;
  assign new_n8599 = new_n8598 ^ new_n8594;
  assign new_n8600 = ~new_n8589 & new_n8599;
  assign new_n8601 = new_n8600 ^ new_n8582;
  assign new_n8602 = ~new_n8586 & new_n8582;
  assign new_n8603 = ~new_n8602 & new_n8596;
  assign new_n8604 = ~new_n8603 & new_n8317;
  assign new_n8605 = new_n8582 & new_n8594;
  assign new_n8606 = ~new_n8588 & ~new_n8605;
  assign new_n8607 = ~new_n8604 & new_n8606;
  assign new_n8608 = n70 & new_n7553;
  assign new_n8609 = ~new_n402 & new_n7543;
  assign new_n8610 = new_n8609 ^ new_n8608;
  assign new_n8611 = n71 & new_n7542;
  assign new_n8612 = n69 & new_n7547;
  assign new_n8613 = new_n8612 ^ new_n8611;
  assign new_n8614 = new_n8613 ^ new_n8610;
  assign new_n8615 = new_n8614 ^ n57;
  assign new_n8616 = ~new_n154 & new_n8343;
  assign new_n8617 = new_n8616 ^ n68;
  assign new_n8618 = new_n7837 & new_n8617;
  assign new_n8619 = n66 & new_n8349;
  assign new_n8620 = n67 & new_n8355;
  assign new_n8621 = new_n8620 ^ new_n8619;
  assign new_n8622 = ~new_n8618 & ~new_n8621;
  assign new_n8623 = new_n8622 ^ n60;
  assign new_n8624 = ~new_n8357 & new_n8359;
  assign new_n8625 = n61 ^ n60;
  assign new_n8626 = n65 & new_n8625;
  assign new_n8627 = ~new_n8624 & ~new_n8626;
  assign new_n8628 = new_n8627 ^ new_n8623;
  assign new_n8629 = new_n8626 ^ new_n8624;
  assign new_n8630 = new_n8629 ^ new_n8627;
  assign new_n8631 = new_n8630 ^ new_n8628;
  assign new_n8632 = new_n8631 ^ new_n8615;
  assign new_n8633 = new_n8373 ^ new_n8361;
  assign new_n8634 = ~new_n8633 & new_n8365;
  assign new_n8635 = new_n8634 ^ new_n8364;
  assign new_n8636 = new_n8635 ^ new_n8632;
  assign new_n8637 = ~new_n6805 & n73;
  assign new_n8638 = new_n595 & new_n6800;
  assign new_n8639 = new_n8638 ^ new_n8637;
  assign new_n8640 = n74 & new_n6799;
  assign new_n8641 = n72 & new_n6811;
  assign new_n8642 = new_n8641 ^ new_n8640;
  assign new_n8643 = new_n8642 ^ new_n8639;
  assign new_n8644 = new_n8643 ^ n54;
  assign new_n8645 = new_n8644 ^ new_n8636;
  assign new_n8646 = new_n8386 ^ new_n8374;
  assign new_n8647 = ~new_n8383 & new_n8646;
  assign new_n8648 = new_n8647 ^ new_n8386;
  assign new_n8649 = new_n8648 ^ new_n8645;
  assign new_n8650 = ~new_n6110 & n76;
  assign new_n8651 = ~new_n812 & new_n6105;
  assign new_n8652 = new_n8651 ^ new_n8650;
  assign new_n8653 = n77 & new_n6104;
  assign new_n8654 = n75 & new_n6347;
  assign new_n8655 = new_n8654 ^ new_n8653;
  assign new_n8656 = new_n8655 ^ new_n8652;
  assign new_n8657 = new_n8656 ^ n51;
  assign new_n8658 = new_n8657 ^ new_n8649;
  assign new_n8659 = new_n8387 ^ new_n8338;
  assign new_n8660 = ~new_n8659 & new_n8342;
  assign new_n8661 = new_n8660 ^ new_n8341;
  assign new_n8662 = new_n8661 ^ new_n8658;
  assign new_n8663 = ~new_n5424 & n79;
  assign new_n8664 = new_n1069 & new_n5419;
  assign new_n8665 = new_n8664 ^ new_n8663;
  assign new_n8666 = n80 & new_n5418;
  assign new_n8667 = n78 & new_n5648;
  assign new_n8668 = new_n8667 ^ new_n8666;
  assign new_n8669 = new_n8668 ^ new_n8665;
  assign new_n8670 = new_n8669 ^ n48;
  assign new_n8671 = new_n8670 ^ new_n8662;
  assign new_n8672 = new_n8388 ^ new_n8326;
  assign new_n8673 = ~new_n8330 & ~new_n8672;
  assign new_n8674 = new_n8673 ^ new_n8329;
  assign new_n8675 = new_n8674 ^ new_n8671;
  assign new_n8676 = ~new_n4804 & n82;
  assign new_n8677 = new_n1363 & new_n4799;
  assign new_n8678 = new_n8677 ^ new_n8676;
  assign new_n8679 = n83 & new_n4798;
  assign new_n8680 = n81 & new_n4810;
  assign new_n8681 = new_n8680 ^ new_n8679;
  assign new_n8682 = new_n8681 ^ new_n8678;
  assign new_n8683 = new_n8682 ^ n45;
  assign new_n8684 = new_n8683 ^ new_n8675;
  assign new_n8685 = new_n8401 ^ new_n8389;
  assign new_n8686 = ~new_n8685 & new_n8398;
  assign new_n8687 = new_n8686 ^ new_n8401;
  assign new_n8688 = new_n8687 ^ new_n8684;
  assign new_n8689 = ~new_n4212 & n85;
  assign new_n8690 = new_n1694 & new_n4201;
  assign new_n8691 = new_n8690 ^ new_n8689;
  assign new_n8692 = n86 & new_n4200;
  assign new_n8693 = n84 & new_n4206;
  assign new_n8694 = new_n8693 ^ new_n8692;
  assign new_n8695 = new_n8694 ^ new_n8691;
  assign new_n8696 = new_n8695 ^ n42;
  assign new_n8697 = new_n8696 ^ new_n8688;
  assign new_n8698 = new_n8414 ^ new_n8402;
  assign new_n8699 = ~new_n8698 & new_n8411;
  assign new_n8700 = new_n8699 ^ new_n8414;
  assign new_n8701 = new_n8700 ^ new_n8697;
  assign new_n8702 = ~new_n3682 & n88;
  assign new_n8703 = new_n2063 & new_n3677;
  assign new_n8704 = new_n8703 ^ new_n8702;
  assign new_n8705 = n89 & new_n3676;
  assign new_n8706 = n87 & new_n3688;
  assign new_n8707 = new_n8706 ^ new_n8705;
  assign new_n8708 = new_n8707 ^ new_n8704;
  assign new_n8709 = new_n8708 ^ n39;
  assign new_n8710 = new_n8709 ^ new_n8701;
  assign new_n8711 = new_n8427 ^ new_n8415;
  assign new_n8712 = ~new_n8711 & new_n8424;
  assign new_n8713 = new_n8712 ^ new_n8427;
  assign new_n8714 = new_n8713 ^ new_n8710;
  assign new_n8715 = ~new_n3143 & n91;
  assign new_n8716 = new_n2481 & new_n3138;
  assign new_n8717 = new_n8716 ^ new_n8715;
  assign new_n8718 = n92 & new_n3137;
  assign new_n8719 = n90 & new_n3149;
  assign new_n8720 = new_n8719 ^ new_n8718;
  assign new_n8721 = new_n8720 ^ new_n8717;
  assign new_n8722 = new_n8721 ^ n36;
  assign new_n8723 = new_n8722 ^ new_n8714;
  assign new_n8724 = new_n8440 ^ new_n8428;
  assign new_n8725 = ~new_n8724 & new_n8437;
  assign new_n8726 = new_n8725 ^ new_n8440;
  assign new_n8727 = new_n8726 ^ new_n8723;
  assign new_n8728 = ~new_n2672 & n94;
  assign new_n8729 = new_n2667 & new_n2934;
  assign new_n8730 = new_n8729 ^ new_n8728;
  assign new_n8731 = n95 & new_n2666;
  assign new_n8732 = n93 & new_n2664;
  assign new_n8733 = new_n8732 ^ new_n8731;
  assign new_n8734 = new_n8733 ^ new_n8730;
  assign new_n8735 = new_n8734 ^ n33;
  assign new_n8736 = new_n8735 ^ new_n8727;
  assign new_n8737 = new_n8453 ^ new_n8441;
  assign new_n8738 = new_n8450 & new_n8737;
  assign new_n8739 = new_n8738 ^ new_n8453;
  assign new_n8740 = new_n8739 ^ new_n8736;
  assign new_n8741 = n97 & new_n2246;
  assign new_n8742 = new_n2241 & new_n3435;
  assign new_n8743 = new_n8742 ^ new_n8741;
  assign new_n8744 = n98 & new_n2240;
  assign new_n8745 = n96 & new_n2391;
  assign new_n8746 = new_n8745 ^ new_n8744;
  assign new_n8747 = new_n8746 ^ new_n8743;
  assign new_n8748 = new_n8747 ^ n30;
  assign new_n8749 = new_n8748 ^ new_n8740;
  assign new_n8750 = new_n8466 ^ new_n8462;
  assign new_n8751 = ~new_n8750 & new_n8463;
  assign new_n8752 = new_n8751 ^ new_n8454;
  assign new_n8753 = new_n8752 ^ new_n8749;
  assign new_n8754 = n100 & new_n1874;
  assign new_n8755 = new_n1864 & new_n3972;
  assign new_n8756 = new_n8755 ^ new_n8754;
  assign new_n8757 = n101 & new_n1863;
  assign new_n8758 = n99 & new_n1868;
  assign new_n8759 = new_n8758 ^ new_n8757;
  assign new_n8760 = new_n8759 ^ new_n8756;
  assign new_n8761 = new_n8760 ^ n27;
  assign new_n8762 = new_n8761 ^ new_n8753;
  assign new_n8763 = new_n8479 ^ new_n8467;
  assign new_n8764 = ~new_n8476 & new_n8763;
  assign new_n8765 = new_n8764 ^ new_n8479;
  assign new_n8766 = new_n8765 ^ new_n8762;
  assign new_n8767 = ~new_n1506 & n103;
  assign new_n8768 = ~new_n4556 & new_n1501;
  assign new_n8769 = new_n8768 ^ new_n8767;
  assign new_n8770 = n104 & new_n1500;
  assign new_n8771 = n102 & new_n1512;
  assign new_n8772 = new_n8771 ^ new_n8770;
  assign new_n8773 = new_n8772 ^ new_n8769;
  assign new_n8774 = new_n8773 ^ n24;
  assign new_n8775 = new_n8774 ^ new_n8766;
  assign new_n8776 = new_n8492 ^ new_n8480;
  assign new_n8777 = ~new_n8489 & new_n8776;
  assign new_n8778 = new_n8777 ^ new_n8492;
  assign new_n8779 = new_n8778 ^ new_n8775;
  assign new_n8780 = ~new_n1198 & n106;
  assign new_n8781 = ~new_n5164 & new_n1193;
  assign new_n8782 = new_n8781 ^ new_n8780;
  assign new_n8783 = n107 & new_n1192;
  assign new_n8784 = n105 & new_n1204;
  assign new_n8785 = new_n8784 ^ new_n8783;
  assign new_n8786 = new_n8785 ^ new_n8782;
  assign new_n8787 = new_n8786 ^ n21;
  assign new_n8788 = new_n8787 ^ new_n8779;
  assign new_n8789 = new_n8505 ^ new_n8493;
  assign new_n8790 = ~new_n8502 & new_n8789;
  assign new_n8791 = new_n8790 ^ new_n8505;
  assign new_n8792 = new_n8791 ^ new_n8788;
  assign new_n8793 = ~new_n930 & n109;
  assign new_n8794 = new_n925 & new_n5825;
  assign new_n8795 = new_n8794 ^ new_n8793;
  assign new_n8796 = n110 & new_n924;
  assign new_n8797 = n108 & new_n936;
  assign new_n8798 = new_n8797 ^ new_n8796;
  assign new_n8799 = new_n8798 ^ new_n8795;
  assign new_n8800 = new_n8799 ^ n18;
  assign new_n8801 = new_n8800 ^ new_n8792;
  assign new_n8802 = new_n8518 ^ new_n8506;
  assign new_n8803 = ~new_n8515 & new_n8802;
  assign new_n8804 = new_n8803 ^ new_n8518;
  assign new_n8805 = new_n8804 ^ new_n8801;
  assign new_n8806 = n112 & new_n707;
  assign new_n8807 = ~new_n6518 & new_n701;
  assign new_n8808 = new_n8807 ^ new_n8806;
  assign new_n8809 = n113 & new_n700;
  assign new_n8810 = n111 & new_n787;
  assign new_n8811 = new_n8810 ^ new_n8809;
  assign new_n8812 = new_n8811 ^ new_n8808;
  assign new_n8813 = new_n8812 ^ n15;
  assign new_n8814 = new_n8813 ^ new_n8805;
  assign new_n8815 = new_n8531 ^ new_n8519;
  assign new_n8816 = ~new_n8528 & new_n8815;
  assign new_n8817 = new_n8816 ^ new_n8531;
  assign new_n8818 = new_n8817 ^ new_n8814;
  assign new_n8819 = n115 & new_n499;
  assign new_n8820 = ~new_n506 & ~new_n7256;
  assign new_n8821 = new_n8820 ^ new_n8819;
  assign new_n8822 = ~new_n505 & n116;
  assign new_n8823 = n114 & new_n579;
  assign new_n8824 = new_n8823 ^ new_n8822;
  assign new_n8825 = new_n8824 ^ new_n8821;
  assign new_n8826 = new_n8825 ^ n12;
  assign new_n8827 = new_n8826 ^ new_n8818;
  assign new_n8828 = new_n8544 ^ new_n8532;
  assign new_n8829 = ~new_n8541 & new_n8828;
  assign new_n8830 = new_n8829 ^ new_n8544;
  assign new_n8831 = new_n8830 ^ new_n8827;
  assign new_n8832 = n118 & new_n354;
  assign new_n8833 = ~new_n8019 & new_n349;
  assign new_n8834 = new_n8833 ^ new_n8832;
  assign new_n8835 = n119 & new_n348;
  assign new_n8836 = n117 & new_n391;
  assign new_n8837 = new_n8836 ^ new_n8835;
  assign new_n8838 = new_n8837 ^ new_n8834;
  assign new_n8839 = new_n8838 ^ n9;
  assign new_n8840 = new_n8839 ^ new_n8831;
  assign new_n8841 = new_n8557 ^ new_n8545;
  assign new_n8842 = ~new_n8554 & new_n8841;
  assign new_n8843 = new_n8842 ^ new_n8557;
  assign new_n8844 = new_n8843 ^ new_n8840;
  assign new_n8845 = new_n8580 ^ new_n8558;
  assign new_n8846 = ~new_n8581 & new_n8845;
  assign new_n8847 = new_n8846 ^ new_n8558;
  assign new_n8848 = new_n8847 ^ new_n8844;
  assign new_n8849 = n121 & new_n218;
  assign new_n8850 = new_n8046 ^ n122;
  assign new_n8851 = new_n208 & new_n8850;
  assign new_n8852 = new_n8851 ^ new_n8849;
  assign new_n8853 = n122 & new_n207;
  assign new_n8854 = n120 & new_n212;
  assign new_n8855 = new_n8854 ^ new_n8853;
  assign new_n8856 = new_n8855 ^ new_n8852;
  assign new_n8857 = new_n8856 ^ n6;
  assign new_n8858 = n123 & new_n180;
  assign new_n8859 = n2 & n124;
  assign new_n8860 = new_n8859 ^ new_n8858;
  assign new_n8861 = new_n8860 ^ n3;
  assign new_n8862 = n124 ^ n123;
  assign new_n8863 = new_n8574 & new_n8862;
  assign new_n8864 = ~new_n8863 & new_n155;
  assign new_n8865 = new_n8864 ^ n2;
  assign new_n8866 = new_n8865 ^ n125;
  assign new_n8867 = new_n8866 ^ new_n8861;
  assign new_n8868 = ~n1 & new_n8867;
  assign new_n8869 = new_n8868 ^ new_n8866;
  assign new_n8870 = new_n8869 ^ new_n8857;
  assign new_n8871 = new_n8870 ^ new_n8848;
  assign new_n8872 = new_n8871 ^ new_n8607;
  assign new_n8873 = ~new_n8847 & new_n8844;
  assign new_n8874 = new_n8857 & new_n8869;
  assign new_n8875 = new_n8874 ^ new_n8870;
  assign new_n8876 = ~new_n8875 & new_n8873;
  assign new_n8877 = new_n8873 ^ new_n8848;
  assign new_n8878 = new_n8874 & new_n8877;
  assign new_n8879 = new_n8878 ^ new_n8876;
  assign new_n8880 = new_n8879 ^ new_n8871;
  assign new_n8881 = ~new_n8607 & ~new_n8880;
  assign new_n8882 = new_n8875 ^ new_n8847;
  assign new_n8883 = ~new_n8848 & new_n8882;
  assign new_n8884 = new_n8883 ^ new_n8847;
  assign new_n8885 = ~new_n8874 & ~new_n8884;
  assign new_n8886 = new_n8885 ^ new_n8881;
  assign new_n8887 = ~new_n8879 & ~new_n8886;
  assign new_n8888 = ~new_n6110 & n77;
  assign new_n8889 = ~new_n891 & new_n6105;
  assign new_n8890 = new_n8889 ^ new_n8888;
  assign new_n8891 = n78 & new_n6104;
  assign new_n8892 = n76 & new_n6347;
  assign new_n8893 = new_n8892 ^ new_n8891;
  assign new_n8894 = new_n8893 ^ new_n8890;
  assign new_n8895 = new_n8894 ^ n51;
  assign new_n8896 = new_n8661 ^ new_n8649;
  assign new_n8897 = ~new_n8896 & new_n8658;
  assign new_n8898 = new_n8897 ^ new_n8661;
  assign new_n8899 = new_n8898 ^ new_n8895;
  assign new_n8900 = n71 & new_n7553;
  assign new_n8901 = ~new_n459 & new_n7543;
  assign new_n8902 = new_n8901 ^ new_n8900;
  assign new_n8903 = n72 & new_n7542;
  assign new_n8904 = n70 & new_n7547;
  assign new_n8905 = new_n8904 ^ new_n8903;
  assign new_n8906 = new_n8905 ^ new_n8902;
  assign new_n8907 = new_n8906 ^ n57;
  assign new_n8908 = ~new_n8623 & ~new_n8627;
  assign new_n8909 = n66 ^ n61;
  assign new_n8910 = ~new_n8909 & new_n8625;
  assign new_n8911 = new_n8910 ^ n60;
  assign new_n8912 = new_n8911 ^ n62;
  assign new_n8913 = n60 & n61;
  assign new_n8914 = new_n8913 ^ n62;
  assign new_n8915 = ~n65 & new_n8914;
  assign new_n8916 = new_n8915 ^ new_n8912;
  assign new_n8917 = new_n8916 ^ new_n8908;
  assign new_n8918 = n68 & new_n8355;
  assign new_n8919 = ~new_n304 & new_n8345;
  assign new_n8920 = new_n8919 ^ new_n8918;
  assign new_n8921 = n69 & new_n8344;
  assign new_n8922 = n67 & new_n8349;
  assign new_n8923 = new_n8922 ^ new_n8921;
  assign new_n8924 = new_n8923 ^ new_n8920;
  assign new_n8925 = new_n8924 ^ n60;
  assign new_n8926 = new_n8925 ^ new_n8917;
  assign new_n8927 = new_n8926 ^ new_n8907;
  assign new_n8928 = new_n8635 ^ new_n8631;
  assign new_n8929 = ~new_n8928 & new_n8632;
  assign new_n8930 = new_n8929 ^ new_n8635;
  assign new_n8931 = new_n8930 ^ new_n8927;
  assign new_n8932 = ~new_n6805 & n74;
  assign new_n8933 = new_n660 & new_n6800;
  assign new_n8934 = new_n8933 ^ new_n8932;
  assign new_n8935 = n75 & new_n6799;
  assign new_n8936 = n73 & new_n6811;
  assign new_n8937 = new_n8936 ^ new_n8935;
  assign new_n8938 = new_n8937 ^ new_n8934;
  assign new_n8939 = new_n8938 ^ n54;
  assign new_n8940 = new_n8939 ^ new_n8931;
  assign new_n8941 = new_n8648 ^ new_n8636;
  assign new_n8942 = ~new_n8941 & new_n8645;
  assign new_n8943 = new_n8942 ^ new_n8648;
  assign new_n8944 = new_n8943 ^ new_n8940;
  assign new_n8945 = new_n8944 ^ new_n8899;
  assign new_n8946 = ~new_n5424 & n80;
  assign new_n8947 = new_n1161 & new_n5419;
  assign new_n8948 = new_n8947 ^ new_n8946;
  assign new_n8949 = n81 & new_n5418;
  assign new_n8950 = n79 & new_n5648;
  assign new_n8951 = new_n8950 ^ new_n8949;
  assign new_n8952 = new_n8951 ^ new_n8948;
  assign new_n8953 = new_n8952 ^ n48;
  assign new_n8954 = new_n8953 ^ new_n8945;
  assign new_n8955 = new_n8674 ^ new_n8662;
  assign new_n8956 = new_n8671 & new_n8955;
  assign new_n8957 = new_n8956 ^ new_n8674;
  assign new_n8958 = new_n8957 ^ new_n8954;
  assign new_n8959 = ~new_n4804 & n83;
  assign new_n8960 = new_n1468 & new_n4799;
  assign new_n8961 = new_n8960 ^ new_n8959;
  assign new_n8962 = n84 & new_n4798;
  assign new_n8963 = n82 & new_n4810;
  assign new_n8964 = new_n8963 ^ new_n8962;
  assign new_n8965 = new_n8964 ^ new_n8961;
  assign new_n8966 = new_n8965 ^ n45;
  assign new_n8967 = new_n8966 ^ new_n8958;
  assign new_n8968 = new_n8687 ^ new_n8675;
  assign new_n8969 = ~new_n8684 & new_n8968;
  assign new_n8970 = new_n8969 ^ new_n8687;
  assign new_n8971 = new_n8970 ^ new_n8967;
  assign new_n8972 = ~new_n4212 & n86;
  assign new_n8973 = new_n1811 & new_n4201;
  assign new_n8974 = new_n8973 ^ new_n8972;
  assign new_n8975 = n87 & new_n4200;
  assign new_n8976 = n85 & new_n4206;
  assign new_n8977 = new_n8976 ^ new_n8975;
  assign new_n8978 = new_n8977 ^ new_n8974;
  assign new_n8979 = new_n8978 ^ n42;
  assign new_n8980 = new_n8979 ^ new_n8971;
  assign new_n8981 = new_n8700 ^ new_n8688;
  assign new_n8982 = ~new_n8697 & new_n8981;
  assign new_n8983 = new_n8982 ^ new_n8700;
  assign new_n8984 = new_n8983 ^ new_n8980;
  assign new_n8985 = ~new_n3682 & n89;
  assign new_n8986 = new_n2193 & new_n3677;
  assign new_n8987 = new_n8986 ^ new_n8985;
  assign new_n8988 = n90 & new_n3676;
  assign new_n8989 = n88 & new_n3688;
  assign new_n8990 = new_n8989 ^ new_n8988;
  assign new_n8991 = new_n8990 ^ new_n8987;
  assign new_n8992 = new_n8991 ^ n39;
  assign new_n8993 = new_n8992 ^ new_n8984;
  assign new_n8994 = new_n8713 ^ new_n8701;
  assign new_n8995 = ~new_n8710 & new_n8994;
  assign new_n8996 = new_n8995 ^ new_n8713;
  assign new_n8997 = new_n8996 ^ new_n8993;
  assign new_n8998 = ~new_n3143 & n92;
  assign new_n8999 = new_n2628 & new_n3138;
  assign new_n9000 = new_n8999 ^ new_n8998;
  assign new_n9001 = n93 & new_n3137;
  assign new_n9002 = n91 & new_n3149;
  assign new_n9003 = new_n9002 ^ new_n9001;
  assign new_n9004 = new_n9003 ^ new_n9000;
  assign new_n9005 = new_n9004 ^ n36;
  assign new_n9006 = new_n9005 ^ new_n8997;
  assign new_n9007 = new_n8726 ^ new_n8714;
  assign new_n9008 = ~new_n8723 & new_n9007;
  assign new_n9009 = new_n9008 ^ new_n8726;
  assign new_n9010 = new_n9009 ^ new_n9006;
  assign new_n9011 = ~new_n2672 & n95;
  assign new_n9012 = new_n2667 & new_n3095;
  assign new_n9013 = new_n9012 ^ new_n9011;
  assign new_n9014 = n96 & new_n2666;
  assign new_n9015 = n94 & new_n2664;
  assign new_n9016 = new_n9015 ^ new_n9014;
  assign new_n9017 = new_n9016 ^ new_n9013;
  assign new_n9018 = new_n9017 ^ n33;
  assign new_n9019 = new_n9018 ^ new_n9010;
  assign new_n9020 = new_n8739 ^ new_n8727;
  assign new_n9021 = ~new_n8736 & ~new_n9020;
  assign new_n9022 = new_n9021 ^ new_n8739;
  assign new_n9023 = new_n9022 ^ new_n9019;
  assign new_n9024 = n98 & new_n2246;
  assign new_n9025 = new_n2241 & new_n3604;
  assign new_n9026 = new_n9025 ^ new_n9024;
  assign new_n9027 = n99 & new_n2240;
  assign new_n9028 = n97 & new_n2391;
  assign new_n9029 = new_n9028 ^ new_n9027;
  assign new_n9030 = new_n9029 ^ new_n9026;
  assign new_n9031 = new_n9030 ^ n30;
  assign new_n9032 = new_n9031 ^ new_n9023;
  assign new_n9033 = new_n8752 ^ new_n8748;
  assign new_n9034 = ~new_n8749 & ~new_n9033;
  assign new_n9035 = new_n9034 ^ new_n8740;
  assign new_n9036 = new_n9035 ^ new_n9032;
  assign new_n9037 = n101 & new_n1874;
  assign new_n9038 = new_n1864 & new_n4159;
  assign new_n9039 = new_n9038 ^ new_n9037;
  assign new_n9040 = n102 & new_n1863;
  assign new_n9041 = n100 & new_n1868;
  assign new_n9042 = new_n9041 ^ new_n9040;
  assign new_n9043 = new_n9042 ^ new_n9039;
  assign new_n9044 = new_n9043 ^ n27;
  assign new_n9045 = new_n9044 ^ new_n9036;
  assign new_n9046 = new_n8765 ^ new_n8753;
  assign new_n9047 = ~new_n9046 & new_n8762;
  assign new_n9048 = new_n9047 ^ new_n8765;
  assign new_n9049 = new_n9048 ^ new_n9045;
  assign new_n9050 = ~new_n1506 & n104;
  assign new_n9051 = ~new_n4754 & new_n1501;
  assign new_n9052 = new_n9051 ^ new_n9050;
  assign new_n9053 = n105 & new_n1500;
  assign new_n9054 = n103 & new_n1512;
  assign new_n9055 = new_n9054 ^ new_n9053;
  assign new_n9056 = new_n9055 ^ new_n9052;
  assign new_n9057 = new_n9056 ^ n24;
  assign new_n9058 = new_n9057 ^ new_n9049;
  assign new_n9059 = new_n8778 ^ new_n8766;
  assign new_n9060 = ~new_n9059 & new_n8775;
  assign new_n9061 = new_n9060 ^ new_n8778;
  assign new_n9062 = new_n9061 ^ new_n9058;
  assign new_n9063 = ~new_n1198 & n107;
  assign new_n9064 = ~new_n5377 & new_n1193;
  assign new_n9065 = new_n9064 ^ new_n9063;
  assign new_n9066 = n108 & new_n1192;
  assign new_n9067 = n106 & new_n1204;
  assign new_n9068 = new_n9067 ^ new_n9066;
  assign new_n9069 = new_n9068 ^ new_n9065;
  assign new_n9070 = new_n9069 ^ n21;
  assign new_n9071 = new_n9070 ^ new_n9062;
  assign new_n9072 = new_n8791 ^ new_n8779;
  assign new_n9073 = ~new_n9072 & new_n8788;
  assign new_n9074 = new_n9073 ^ new_n8791;
  assign new_n9075 = new_n9074 ^ new_n9071;
  assign new_n9076 = ~new_n930 & n110;
  assign new_n9077 = new_n925 & new_n6049;
  assign new_n9078 = new_n9077 ^ new_n9076;
  assign new_n9079 = n111 & new_n924;
  assign new_n9080 = n109 & new_n936;
  assign new_n9081 = new_n9080 ^ new_n9079;
  assign new_n9082 = new_n9081 ^ new_n9078;
  assign new_n9083 = new_n9082 ^ n18;
  assign new_n9084 = new_n9083 ^ new_n9075;
  assign new_n9085 = new_n8804 ^ new_n8792;
  assign new_n9086 = ~new_n9085 & new_n8801;
  assign new_n9087 = new_n9086 ^ new_n8804;
  assign new_n9088 = new_n9087 ^ new_n9084;
  assign new_n9089 = n113 & new_n707;
  assign new_n9090 = ~new_n6764 & new_n701;
  assign new_n9091 = new_n9090 ^ new_n9089;
  assign new_n9092 = n114 & new_n700;
  assign new_n9093 = n112 & new_n787;
  assign new_n9094 = new_n9093 ^ new_n9092;
  assign new_n9095 = new_n9094 ^ new_n9091;
  assign new_n9096 = new_n9095 ^ n15;
  assign new_n9097 = new_n9096 ^ new_n9088;
  assign new_n9098 = new_n8817 ^ new_n8805;
  assign new_n9099 = ~new_n9098 & new_n8814;
  assign new_n9100 = new_n9099 ^ new_n8817;
  assign new_n9101 = new_n9100 ^ new_n9097;
  assign new_n9102 = n116 & new_n499;
  assign new_n9103 = ~new_n506 & ~new_n7503;
  assign new_n9104 = new_n9103 ^ new_n9102;
  assign new_n9105 = ~new_n505 & n117;
  assign new_n9106 = n115 & new_n579;
  assign new_n9107 = new_n9106 ^ new_n9105;
  assign new_n9108 = new_n9107 ^ new_n9104;
  assign new_n9109 = new_n9108 ^ n12;
  assign new_n9110 = new_n9109 ^ new_n9101;
  assign new_n9111 = new_n8830 ^ new_n8818;
  assign new_n9112 = ~new_n9111 & new_n8827;
  assign new_n9113 = new_n9112 ^ new_n8830;
  assign new_n9114 = new_n9113 ^ new_n9110;
  assign new_n9115 = n122 & new_n218;
  assign new_n9116 = new_n8302 ^ n123;
  assign new_n9117 = ~new_n9116 & new_n208;
  assign new_n9118 = new_n9117 ^ new_n9115;
  assign new_n9119 = n123 & new_n207;
  assign new_n9120 = n121 & new_n212;
  assign new_n9121 = new_n9120 ^ new_n9119;
  assign new_n9122 = new_n9121 ^ new_n9118;
  assign new_n9123 = new_n9122 ^ n6;
  assign new_n9124 = n119 & new_n354;
  assign new_n9125 = new_n349 & new_n8286;
  assign new_n9126 = new_n9125 ^ new_n9124;
  assign new_n9127 = n120 & new_n348;
  assign new_n9128 = n118 & new_n391;
  assign new_n9129 = new_n9128 ^ new_n9127;
  assign new_n9130 = new_n9129 ^ new_n9126;
  assign new_n9131 = new_n9130 ^ n9;
  assign new_n9132 = new_n9131 ^ new_n9123;
  assign new_n9133 = n124 & new_n180;
  assign new_n9134 = n2 & n125;
  assign new_n9135 = new_n9134 ^ new_n9133;
  assign new_n9136 = new_n9135 ^ n3;
  assign new_n9137 = n125 & new_n8572;
  assign new_n9138 = ~n124 & ~new_n9137;
  assign new_n9139 = ~n125 & new_n8573;
  assign new_n9140 = ~new_n9138 & ~new_n9139;
  assign new_n9141 = new_n9140 ^ n125;
  assign new_n9142 = ~new_n9141 & new_n155;
  assign new_n9143 = new_n9142 ^ n2;
  assign new_n9144 = new_n9143 ^ n126;
  assign new_n9145 = new_n9144 ^ new_n9136;
  assign new_n9146 = ~n1 & new_n9145;
  assign new_n9147 = new_n9146 ^ new_n9144;
  assign new_n9148 = new_n9147 ^ new_n9132;
  assign new_n9149 = new_n9148 ^ new_n9114;
  assign new_n9150 = new_n8843 ^ new_n8831;
  assign new_n9151 = ~new_n9150 & new_n8840;
  assign new_n9152 = new_n9151 ^ new_n8843;
  assign new_n9153 = new_n9152 ^ new_n9149;
  assign new_n9154 = new_n9153 ^ new_n8887;
  assign new_n9155 = ~new_n8877 & new_n9153;
  assign new_n9156 = ~new_n9155 & new_n8874;
  assign new_n9157 = ~new_n9156 & new_n8607;
  assign new_n9158 = ~new_n8876 & ~new_n9153;
  assign new_n9159 = new_n8885 ^ new_n8880;
  assign new_n9160 = ~new_n9158 & new_n9159;
  assign new_n9161 = ~new_n9157 & ~new_n9160;
  assign new_n9162 = ~new_n9153 & new_n8884;
  assign new_n9163 = ~new_n9161 & ~new_n9162;
  assign new_n9164 = ~new_n6805 & n75;
  assign new_n9165 = ~new_n737 & new_n6800;
  assign new_n9166 = new_n9165 ^ new_n9164;
  assign new_n9167 = n76 & new_n6799;
  assign new_n9168 = n74 & new_n6811;
  assign new_n9169 = new_n9168 ^ new_n9167;
  assign new_n9170 = new_n9169 ^ new_n9166;
  assign new_n9171 = new_n9170 ^ n54;
  assign new_n9172 = new_n8943 ^ new_n8931;
  assign new_n9173 = ~new_n8940 & new_n9172;
  assign new_n9174 = new_n9173 ^ new_n8943;
  assign new_n9175 = new_n9174 ^ new_n9171;
  assign new_n9176 = n69 & new_n8355;
  assign new_n9177 = ~new_n339 & new_n8345;
  assign new_n9178 = new_n9177 ^ new_n9176;
  assign new_n9179 = n70 & new_n8344;
  assign new_n9180 = n68 & new_n8349;
  assign new_n9181 = new_n9180 ^ new_n9179;
  assign new_n9182 = new_n9181 ^ new_n9178;
  assign new_n9183 = n63 ^ n62;
  assign new_n9184 = ~new_n9183 & new_n8625;
  assign new_n9185 = new_n9184 ^ new_n8625;
  assign new_n9186 = ~new_n151 & new_n9185;
  assign new_n9187 = ~new_n8625 & n63;
  assign new_n9188 = new_n9187 ^ new_n8913;
  assign new_n9189 = new_n9183 & new_n9188;
  assign new_n9190 = n65 & new_n9189;
  assign new_n9191 = new_n9190 ^ new_n9186;
  assign new_n9192 = n67 & new_n8625;
  assign new_n9193 = new_n9192 ^ new_n9191;
  assign new_n9194 = ~new_n8625 & n62;
  assign new_n9195 = new_n9194 ^ new_n8913;
  assign new_n9196 = n66 & new_n9195;
  assign new_n9197 = new_n9196 ^ new_n9193;
  assign new_n9198 = ~new_n8626 & ~new_n8916;
  assign new_n9199 = n63 & new_n9198;
  assign new_n9200 = new_n9199 ^ n63;
  assign new_n9201 = new_n9200 ^ new_n9197;
  assign new_n9202 = new_n9201 ^ new_n9182;
  assign new_n9203 = new_n8916 ^ n60;
  assign new_n9204 = new_n9203 ^ new_n8924;
  assign new_n9205 = ~new_n8917 & new_n9204;
  assign new_n9206 = new_n9205 ^ new_n8924;
  assign new_n9207 = new_n9206 ^ new_n9202;
  assign new_n9208 = n72 & new_n7553;
  assign new_n9209 = new_n534 & new_n7543;
  assign new_n9210 = new_n9209 ^ new_n9208;
  assign new_n9211 = n73 & new_n7542;
  assign new_n9212 = n71 & new_n7547;
  assign new_n9213 = new_n9212 ^ new_n9211;
  assign new_n9214 = new_n9213 ^ new_n9210;
  assign new_n9215 = new_n9214 ^ n57;
  assign new_n9216 = new_n9215 ^ new_n9207;
  assign new_n9217 = new_n8930 ^ new_n8907;
  assign new_n9218 = ~new_n8927 & new_n9217;
  assign new_n9219 = new_n9218 ^ new_n8930;
  assign new_n9220 = new_n9219 ^ new_n9216;
  assign new_n9221 = new_n9220 ^ new_n9175;
  assign new_n9222 = ~new_n5424 & n81;
  assign new_n9223 = new_n1263 & new_n5419;
  assign new_n9224 = new_n9223 ^ new_n9222;
  assign new_n9225 = n82 & new_n5418;
  assign new_n9226 = n80 & new_n5648;
  assign new_n9227 = new_n9226 ^ new_n9225;
  assign new_n9228 = new_n9227 ^ new_n9224;
  assign new_n9229 = new_n9228 ^ n48;
  assign new_n9230 = ~new_n6110 & n78;
  assign new_n9231 = ~new_n982 & new_n6105;
  assign new_n9232 = new_n9231 ^ new_n9230;
  assign new_n9233 = n79 & new_n6104;
  assign new_n9234 = n77 & new_n6347;
  assign new_n9235 = new_n9234 ^ new_n9233;
  assign new_n9236 = new_n9235 ^ new_n9232;
  assign new_n9237 = new_n9236 ^ n51;
  assign new_n9238 = new_n9237 ^ new_n9229;
  assign new_n9239 = new_n9238 ^ new_n9221;
  assign new_n9240 = new_n8944 ^ new_n8895;
  assign new_n9241 = ~new_n9240 & new_n8899;
  assign new_n9242 = new_n9241 ^ new_n8898;
  assign new_n9243 = new_n9242 ^ new_n9239;
  assign new_n9244 = new_n8957 ^ new_n8945;
  assign new_n9245 = ~new_n8954 & ~new_n9244;
  assign new_n9246 = new_n9245 ^ new_n8957;
  assign new_n9247 = new_n9246 ^ new_n9243;
  assign new_n9248 = ~new_n4804 & n84;
  assign new_n9249 = new_n1584 & new_n4799;
  assign new_n9250 = new_n9249 ^ new_n9248;
  assign new_n9251 = n85 & new_n4798;
  assign new_n9252 = n83 & new_n4810;
  assign new_n9253 = new_n9252 ^ new_n9251;
  assign new_n9254 = new_n9253 ^ new_n9250;
  assign new_n9255 = new_n9254 ^ n45;
  assign new_n9256 = new_n9255 ^ new_n9247;
  assign new_n9257 = new_n8970 ^ new_n8958;
  assign new_n9258 = ~new_n9257 & new_n8967;
  assign new_n9259 = new_n9258 ^ new_n8970;
  assign new_n9260 = new_n9259 ^ new_n9256;
  assign new_n9261 = ~new_n4212 & n87;
  assign new_n9262 = new_n1940 & new_n4201;
  assign new_n9263 = new_n9262 ^ new_n9261;
  assign new_n9264 = n88 & new_n4200;
  assign new_n9265 = n86 & new_n4206;
  assign new_n9266 = new_n9265 ^ new_n9264;
  assign new_n9267 = new_n9266 ^ new_n9263;
  assign new_n9268 = new_n9267 ^ n42;
  assign new_n9269 = new_n9268 ^ new_n9260;
  assign new_n9270 = new_n8983 ^ new_n8971;
  assign new_n9271 = ~new_n9270 & new_n8980;
  assign new_n9272 = new_n9271 ^ new_n8983;
  assign new_n9273 = new_n9272 ^ new_n9269;
  assign new_n9274 = ~new_n3682 & n90;
  assign new_n9275 = new_n2341 & new_n3677;
  assign new_n9276 = new_n9275 ^ new_n9274;
  assign new_n9277 = n91 & new_n3676;
  assign new_n9278 = n89 & new_n3688;
  assign new_n9279 = new_n9278 ^ new_n9277;
  assign new_n9280 = new_n9279 ^ new_n9276;
  assign new_n9281 = new_n9280 ^ n39;
  assign new_n9282 = new_n9281 ^ new_n9273;
  assign new_n9283 = new_n8996 ^ new_n8984;
  assign new_n9284 = ~new_n9283 & new_n8993;
  assign new_n9285 = new_n9284 ^ new_n8996;
  assign new_n9286 = new_n9285 ^ new_n9282;
  assign new_n9287 = ~new_n3143 & n93;
  assign new_n9288 = new_n2785 & new_n3138;
  assign new_n9289 = new_n9288 ^ new_n9287;
  assign new_n9290 = n94 & new_n3137;
  assign new_n9291 = n92 & new_n3149;
  assign new_n9292 = new_n9291 ^ new_n9290;
  assign new_n9293 = new_n9292 ^ new_n9289;
  assign new_n9294 = new_n9293 ^ n36;
  assign new_n9295 = new_n9294 ^ new_n9286;
  assign new_n9296 = new_n9009 ^ new_n8997;
  assign new_n9297 = ~new_n9296 & new_n9006;
  assign new_n9298 = new_n9297 ^ new_n9009;
  assign new_n9299 = new_n9298 ^ new_n9295;
  assign new_n9300 = ~new_n2672 & n96;
  assign new_n9301 = new_n2667 & new_n3273;
  assign new_n9302 = new_n9301 ^ new_n9300;
  assign new_n9303 = n97 & new_n2666;
  assign new_n9304 = n95 & new_n2664;
  assign new_n9305 = new_n9304 ^ new_n9303;
  assign new_n9306 = new_n9305 ^ new_n9302;
  assign new_n9307 = new_n9306 ^ n33;
  assign new_n9308 = new_n9307 ^ new_n9299;
  assign new_n9309 = new_n9022 ^ new_n9010;
  assign new_n9310 = new_n9019 & new_n9309;
  assign new_n9311 = new_n9310 ^ new_n9022;
  assign new_n9312 = new_n9311 ^ new_n9308;
  assign new_n9313 = n99 & new_n2246;
  assign new_n9314 = new_n2241 & new_n3789;
  assign new_n9315 = new_n9314 ^ new_n9313;
  assign new_n9316 = n100 & new_n2240;
  assign new_n9317 = n98 & new_n2391;
  assign new_n9318 = new_n9317 ^ new_n9316;
  assign new_n9319 = new_n9318 ^ new_n9315;
  assign new_n9320 = new_n9319 ^ n30;
  assign new_n9321 = new_n9320 ^ new_n9312;
  assign new_n9322 = new_n9035 ^ new_n9031;
  assign new_n9323 = new_n9032 & new_n9322;
  assign new_n9324 = new_n9323 ^ new_n9023;
  assign new_n9325 = new_n9324 ^ new_n9321;
  assign new_n9326 = n102 & new_n1874;
  assign new_n9327 = new_n1864 & new_n4368;
  assign new_n9328 = new_n9327 ^ new_n9326;
  assign new_n9329 = n103 & new_n1863;
  assign new_n9330 = n101 & new_n1868;
  assign new_n9331 = new_n9330 ^ new_n9329;
  assign new_n9332 = new_n9331 ^ new_n9328;
  assign new_n9333 = new_n9332 ^ n27;
  assign new_n9334 = new_n9333 ^ new_n9325;
  assign new_n9335 = new_n9048 ^ new_n9036;
  assign new_n9336 = ~new_n9335 & new_n9045;
  assign new_n9337 = new_n9336 ^ new_n9048;
  assign new_n9338 = new_n9337 ^ new_n9334;
  assign new_n9339 = ~new_n1506 & n105;
  assign new_n9340 = ~new_n4961 & new_n1501;
  assign new_n9341 = new_n9340 ^ new_n9339;
  assign new_n9342 = n106 & new_n1500;
  assign new_n9343 = n104 & new_n1512;
  assign new_n9344 = new_n9343 ^ new_n9342;
  assign new_n9345 = new_n9344 ^ new_n9341;
  assign new_n9346 = new_n9345 ^ n24;
  assign new_n9347 = new_n9346 ^ new_n9338;
  assign new_n9348 = new_n9061 ^ new_n9049;
  assign new_n9349 = ~new_n9348 & new_n9058;
  assign new_n9350 = new_n9349 ^ new_n9061;
  assign new_n9351 = new_n9350 ^ new_n9347;
  assign new_n9352 = ~new_n1198 & n108;
  assign new_n9353 = new_n1193 & new_n5604;
  assign new_n9354 = new_n9353 ^ new_n9352;
  assign new_n9355 = n109 & new_n1192;
  assign new_n9356 = n107 & new_n1204;
  assign new_n9357 = new_n9356 ^ new_n9355;
  assign new_n9358 = new_n9357 ^ new_n9354;
  assign new_n9359 = new_n9358 ^ n21;
  assign new_n9360 = new_n9359 ^ new_n9351;
  assign new_n9361 = new_n9074 ^ new_n9062;
  assign new_n9362 = ~new_n9361 & new_n9071;
  assign new_n9363 = new_n9362 ^ new_n9074;
  assign new_n9364 = new_n9363 ^ new_n9360;
  assign new_n9365 = ~new_n930 & n111;
  assign new_n9366 = ~new_n6284 & new_n925;
  assign new_n9367 = new_n9366 ^ new_n9365;
  assign new_n9368 = n112 & new_n924;
  assign new_n9369 = n110 & new_n936;
  assign new_n9370 = new_n9369 ^ new_n9368;
  assign new_n9371 = new_n9370 ^ new_n9367;
  assign new_n9372 = new_n9371 ^ n18;
  assign new_n9373 = new_n9372 ^ new_n9364;
  assign new_n9374 = new_n9087 ^ new_n9075;
  assign new_n9375 = ~new_n9374 & new_n9084;
  assign new_n9376 = new_n9375 ^ new_n9087;
  assign new_n9377 = new_n9376 ^ new_n9373;
  assign new_n9378 = n114 & new_n707;
  assign new_n9379 = ~new_n7013 & new_n701;
  assign new_n9380 = new_n9379 ^ new_n9378;
  assign new_n9381 = n115 & new_n700;
  assign new_n9382 = n113 & new_n787;
  assign new_n9383 = new_n9382 ^ new_n9381;
  assign new_n9384 = new_n9383 ^ new_n9380;
  assign new_n9385 = new_n9384 ^ n15;
  assign new_n9386 = new_n9385 ^ new_n9377;
  assign new_n9387 = new_n9100 ^ new_n9088;
  assign new_n9388 = ~new_n9387 & new_n9097;
  assign new_n9389 = new_n9388 ^ new_n9100;
  assign new_n9390 = new_n9389 ^ new_n9386;
  assign new_n9391 = n117 & new_n499;
  assign new_n9392 = ~new_n506 & ~new_n7761;
  assign new_n9393 = new_n9392 ^ new_n9391;
  assign new_n9394 = ~new_n505 & n118;
  assign new_n9395 = n116 & new_n579;
  assign new_n9396 = new_n9395 ^ new_n9394;
  assign new_n9397 = new_n9396 ^ new_n9393;
  assign new_n9398 = new_n9397 ^ n12;
  assign new_n9399 = new_n9398 ^ new_n9390;
  assign new_n9400 = new_n9113 ^ new_n9101;
  assign new_n9401 = ~new_n9400 & new_n9110;
  assign new_n9402 = new_n9401 ^ new_n9113;
  assign new_n9403 = new_n9402 ^ new_n9399;
  assign new_n9404 = n123 & new_n218;
  assign new_n9405 = new_n8574 ^ n124;
  assign new_n9406 = ~new_n9405 & new_n208;
  assign new_n9407 = new_n9406 ^ new_n9404;
  assign new_n9408 = n124 & new_n207;
  assign new_n9409 = n122 & new_n212;
  assign new_n9410 = new_n9409 ^ new_n9408;
  assign new_n9411 = new_n9410 ^ new_n9407;
  assign new_n9412 = new_n9411 ^ n6;
  assign new_n9413 = n120 & new_n354;
  assign new_n9414 = new_n349 & new_n8560;
  assign new_n9415 = new_n9414 ^ new_n9413;
  assign new_n9416 = n121 & new_n348;
  assign new_n9417 = n119 & new_n391;
  assign new_n9418 = new_n9417 ^ new_n9416;
  assign new_n9419 = new_n9418 ^ new_n9415;
  assign new_n9420 = new_n9419 ^ n9;
  assign new_n9421 = new_n9420 ^ new_n9412;
  assign new_n9422 = new_n9421 ^ new_n9403;
  assign new_n9423 = n126 ^ n125;
  assign new_n9424 = ~n125 & n126;
  assign new_n9425 = new_n9424 ^ new_n9423;
  assign new_n9426 = ~new_n9138 & new_n9425;
  assign new_n9427 = ~new_n9140 & new_n9424;
  assign new_n9428 = new_n9427 ^ new_n9426;
  assign new_n9429 = ~new_n9428 & new_n155;
  assign new_n9430 = new_n9429 ^ n2;
  assign new_n9431 = new_n9430 ^ n127;
  assign new_n9432 = n126 ^ n3;
  assign new_n9433 = n125 ^ n3;
  assign new_n9434 = ~n125 & ~new_n9433;
  assign new_n9435 = new_n9434 ^ new_n9432;
  assign new_n9436 = new_n9435 ^ n125;
  assign new_n9437 = ~new_n9436 & new_n241;
  assign new_n9438 = new_n9437 ^ new_n9434;
  assign new_n9439 = new_n9438 ^ n125;
  assign new_n9440 = new_n9439 ^ new_n9431;
  assign new_n9441 = ~n1 & ~new_n9440;
  assign new_n9442 = new_n9441 ^ new_n9431;
  assign new_n9443 = new_n9442 ^ new_n9422;
  assign new_n9444 = new_n9131 ^ new_n9114;
  assign new_n9445 = new_n9152 ^ new_n9114;
  assign new_n9446 = ~new_n9445 & new_n9444;
  assign new_n9447 = new_n9446 ^ new_n9152;
  assign new_n9448 = new_n9447 ^ new_n9443;
  assign new_n9449 = new_n9147 ^ new_n9123;
  assign new_n9450 = new_n9444 ^ new_n9152;
  assign new_n9451 = new_n9450 ^ new_n9123;
  assign new_n9452 = new_n9449 & new_n9451;
  assign new_n9453 = new_n9452 ^ new_n9147;
  assign new_n9454 = new_n9453 ^ new_n9448;
  assign new_n9455 = new_n9454 ^ new_n9163;
  assign new_n9456 = n73 & new_n7553;
  assign new_n9457 = new_n595 & new_n7543;
  assign new_n9458 = new_n9457 ^ new_n9456;
  assign new_n9459 = n74 & new_n7542;
  assign new_n9460 = n72 & new_n7547;
  assign new_n9461 = new_n9460 ^ new_n9459;
  assign new_n9462 = new_n9461 ^ new_n9458;
  assign new_n9463 = new_n9462 ^ n57;
  assign new_n9464 = new_n9219 ^ new_n9207;
  assign new_n9465 = ~new_n9216 & new_n9464;
  assign new_n9466 = new_n9465 ^ new_n9219;
  assign new_n9467 = new_n9466 ^ new_n9463;
  assign new_n9468 = new_n9202 ^ new_n8924;
  assign new_n9469 = ~new_n9468 & new_n8925;
  assign new_n9470 = new_n8908 & new_n8916;
  assign new_n9471 = new_n9470 ^ new_n8917;
  assign new_n9472 = new_n9469 & new_n9471;
  assign new_n9473 = new_n9470 ^ new_n9201;
  assign new_n9474 = new_n9182 ^ n60;
  assign new_n9475 = new_n9474 ^ new_n9201;
  assign new_n9476 = ~new_n9475 & new_n9473;
  assign new_n9477 = new_n9476 ^ new_n9470;
  assign new_n9478 = ~new_n9472 & ~new_n9477;
  assign new_n9479 = n70 & new_n8355;
  assign new_n9480 = ~new_n402 & new_n8345;
  assign new_n9481 = new_n9480 ^ new_n9479;
  assign new_n9482 = n71 & new_n8344;
  assign new_n9483 = n69 & new_n8349;
  assign new_n9484 = new_n9483 ^ new_n9482;
  assign new_n9485 = new_n9484 ^ new_n9481;
  assign new_n9486 = new_n9485 ^ n60;
  assign new_n9487 = ~new_n154 & new_n9183;
  assign new_n9488 = new_n9487 ^ n68;
  assign new_n9489 = new_n8625 & new_n9488;
  assign new_n9490 = n67 & new_n9195;
  assign new_n9491 = n66 & new_n9189;
  assign new_n9492 = new_n9491 ^ new_n9490;
  assign new_n9493 = ~new_n9489 & ~new_n9492;
  assign new_n9494 = new_n9493 ^ n63;
  assign new_n9495 = n64 ^ n63;
  assign new_n9496 = n65 & new_n9495;
  assign new_n9497 = new_n9496 ^ new_n9494;
  assign new_n9498 = ~new_n9197 & new_n9199;
  assign new_n9499 = new_n9498 ^ new_n9497;
  assign new_n9500 = new_n9499 ^ new_n9486;
  assign new_n9501 = new_n9500 ^ new_n9478;
  assign new_n9502 = new_n9501 ^ new_n9467;
  assign new_n9503 = ~new_n6805 & n76;
  assign new_n9504 = ~new_n812 & new_n6800;
  assign new_n9505 = new_n9504 ^ new_n9503;
  assign new_n9506 = n77 & new_n6799;
  assign new_n9507 = n75 & new_n6811;
  assign new_n9508 = new_n9507 ^ new_n9506;
  assign new_n9509 = new_n9508 ^ new_n9505;
  assign new_n9510 = new_n9509 ^ n54;
  assign new_n9511 = new_n9510 ^ new_n9502;
  assign new_n9512 = new_n9220 ^ new_n9171;
  assign new_n9513 = ~new_n9512 & new_n9175;
  assign new_n9514 = new_n9513 ^ new_n9174;
  assign new_n9515 = new_n9514 ^ new_n9511;
  assign new_n9516 = new_n9242 ^ new_n9221;
  assign new_n9517 = new_n9237 ^ new_n9221;
  assign new_n9518 = ~new_n9517 & new_n9516;
  assign new_n9519 = new_n9518 ^ new_n9242;
  assign new_n9520 = new_n9519 ^ new_n9515;
  assign new_n9521 = ~new_n6110 & n79;
  assign new_n9522 = new_n1069 & new_n6105;
  assign new_n9523 = new_n9522 ^ new_n9521;
  assign new_n9524 = n80 & new_n6104;
  assign new_n9525 = n78 & new_n6347;
  assign new_n9526 = new_n9525 ^ new_n9524;
  assign new_n9527 = new_n9526 ^ new_n9523;
  assign new_n9528 = new_n9527 ^ n51;
  assign new_n9529 = new_n9528 ^ new_n9520;
  assign new_n9530 = ~new_n5424 & n82;
  assign new_n9531 = new_n1363 & new_n5419;
  assign new_n9532 = new_n9531 ^ new_n9530;
  assign new_n9533 = n83 & new_n5418;
  assign new_n9534 = n81 & new_n5648;
  assign new_n9535 = new_n9534 ^ new_n9533;
  assign new_n9536 = new_n9535 ^ new_n9532;
  assign new_n9537 = new_n9536 ^ n48;
  assign new_n9538 = new_n9537 ^ new_n9529;
  assign new_n9539 = new_n9246 ^ new_n9229;
  assign new_n9540 = ~new_n9243 & ~new_n9539;
  assign new_n9541 = new_n9540 ^ new_n9246;
  assign new_n9542 = new_n9541 ^ new_n9538;
  assign new_n9543 = ~new_n4804 & n85;
  assign new_n9544 = new_n1694 & new_n4799;
  assign new_n9545 = new_n9544 ^ new_n9543;
  assign new_n9546 = n86 & new_n4798;
  assign new_n9547 = n84 & new_n4810;
  assign new_n9548 = new_n9547 ^ new_n9546;
  assign new_n9549 = new_n9548 ^ new_n9545;
  assign new_n9550 = new_n9549 ^ n45;
  assign new_n9551 = new_n9550 ^ new_n9542;
  assign new_n9552 = new_n9259 ^ new_n9247;
  assign new_n9553 = ~new_n9552 & new_n9256;
  assign new_n9554 = new_n9553 ^ new_n9259;
  assign new_n9555 = new_n9554 ^ new_n9551;
  assign new_n9556 = ~new_n4212 & n88;
  assign new_n9557 = new_n2063 & new_n4201;
  assign new_n9558 = new_n9557 ^ new_n9556;
  assign new_n9559 = n89 & new_n4200;
  assign new_n9560 = n87 & new_n4206;
  assign new_n9561 = new_n9560 ^ new_n9559;
  assign new_n9562 = new_n9561 ^ new_n9558;
  assign new_n9563 = new_n9562 ^ n42;
  assign new_n9564 = new_n9563 ^ new_n9555;
  assign new_n9565 = new_n9272 ^ new_n9260;
  assign new_n9566 = ~new_n9565 & new_n9269;
  assign new_n9567 = new_n9566 ^ new_n9272;
  assign new_n9568 = new_n9567 ^ new_n9564;
  assign new_n9569 = ~new_n3682 & n91;
  assign new_n9570 = new_n2481 & new_n3677;
  assign new_n9571 = new_n9570 ^ new_n9569;
  assign new_n9572 = n92 & new_n3676;
  assign new_n9573 = n90 & new_n3688;
  assign new_n9574 = new_n9573 ^ new_n9572;
  assign new_n9575 = new_n9574 ^ new_n9571;
  assign new_n9576 = new_n9575 ^ n39;
  assign new_n9577 = new_n9576 ^ new_n9568;
  assign new_n9578 = new_n9285 ^ new_n9273;
  assign new_n9579 = ~new_n9578 & new_n9282;
  assign new_n9580 = new_n9579 ^ new_n9285;
  assign new_n9581 = new_n9580 ^ new_n9577;
  assign new_n9582 = ~new_n3143 & n94;
  assign new_n9583 = new_n2934 & new_n3138;
  assign new_n9584 = new_n9583 ^ new_n9582;
  assign new_n9585 = n95 & new_n3137;
  assign new_n9586 = n93 & new_n3149;
  assign new_n9587 = new_n9586 ^ new_n9585;
  assign new_n9588 = new_n9587 ^ new_n9584;
  assign new_n9589 = new_n9588 ^ n36;
  assign new_n9590 = new_n9589 ^ new_n9581;
  assign new_n9591 = new_n9298 ^ new_n9286;
  assign new_n9592 = ~new_n9591 & new_n9295;
  assign new_n9593 = new_n9592 ^ new_n9298;
  assign new_n9594 = new_n9593 ^ new_n9590;
  assign new_n9595 = ~new_n2672 & n97;
  assign new_n9596 = new_n2667 & new_n3435;
  assign new_n9597 = new_n9596 ^ new_n9595;
  assign new_n9598 = n98 & new_n2666;
  assign new_n9599 = n96 & new_n2664;
  assign new_n9600 = new_n9599 ^ new_n9598;
  assign new_n9601 = new_n9600 ^ new_n9597;
  assign new_n9602 = new_n9601 ^ n33;
  assign new_n9603 = new_n9602 ^ new_n9594;
  assign new_n9604 = new_n9311 ^ new_n9299;
  assign new_n9605 = new_n9308 & new_n9604;
  assign new_n9606 = new_n9605 ^ new_n9311;
  assign new_n9607 = new_n9606 ^ new_n9603;
  assign new_n9608 = n100 & new_n2246;
  assign new_n9609 = new_n2241 & new_n3972;
  assign new_n9610 = new_n9609 ^ new_n9608;
  assign new_n9611 = n101 & new_n2240;
  assign new_n9612 = n99 & new_n2391;
  assign new_n9613 = new_n9612 ^ new_n9611;
  assign new_n9614 = new_n9613 ^ new_n9610;
  assign new_n9615 = new_n9614 ^ n30;
  assign new_n9616 = new_n9615 ^ new_n9607;
  assign new_n9617 = new_n9324 ^ new_n9320;
  assign new_n9618 = ~new_n9617 & new_n9321;
  assign new_n9619 = new_n9618 ^ new_n9312;
  assign new_n9620 = new_n9619 ^ new_n9616;
  assign new_n9621 = n103 & new_n1874;
  assign new_n9622 = ~new_n4556 & new_n1864;
  assign new_n9623 = new_n9622 ^ new_n9621;
  assign new_n9624 = n104 & new_n1863;
  assign new_n9625 = n102 & new_n1868;
  assign new_n9626 = new_n9625 ^ new_n9624;
  assign new_n9627 = new_n9626 ^ new_n9623;
  assign new_n9628 = new_n9627 ^ n27;
  assign new_n9629 = new_n9628 ^ new_n9620;
  assign new_n9630 = new_n9337 ^ new_n9325;
  assign new_n9631 = ~new_n9334 & new_n9630;
  assign new_n9632 = new_n9631 ^ new_n9337;
  assign new_n9633 = new_n9632 ^ new_n9629;
  assign new_n9634 = ~new_n1506 & n106;
  assign new_n9635 = ~new_n5164 & new_n1501;
  assign new_n9636 = new_n9635 ^ new_n9634;
  assign new_n9637 = n107 & new_n1500;
  assign new_n9638 = n105 & new_n1512;
  assign new_n9639 = new_n9638 ^ new_n9637;
  assign new_n9640 = new_n9639 ^ new_n9636;
  assign new_n9641 = new_n9640 ^ n24;
  assign new_n9642 = new_n9641 ^ new_n9633;
  assign new_n9643 = new_n9350 ^ new_n9338;
  assign new_n9644 = ~new_n9347 & new_n9643;
  assign new_n9645 = new_n9644 ^ new_n9350;
  assign new_n9646 = new_n9645 ^ new_n9642;
  assign new_n9647 = ~new_n1198 & n109;
  assign new_n9648 = new_n1193 & new_n5825;
  assign new_n9649 = new_n9648 ^ new_n9647;
  assign new_n9650 = n110 & new_n1192;
  assign new_n9651 = n108 & new_n1204;
  assign new_n9652 = new_n9651 ^ new_n9650;
  assign new_n9653 = new_n9652 ^ new_n9649;
  assign new_n9654 = new_n9653 ^ n21;
  assign new_n9655 = new_n9654 ^ new_n9646;
  assign new_n9656 = new_n9363 ^ new_n9351;
  assign new_n9657 = ~new_n9360 & new_n9656;
  assign new_n9658 = new_n9657 ^ new_n9363;
  assign new_n9659 = new_n9658 ^ new_n9655;
  assign new_n9660 = ~new_n930 & n112;
  assign new_n9661 = ~new_n6518 & new_n925;
  assign new_n9662 = new_n9661 ^ new_n9660;
  assign new_n9663 = n113 & new_n924;
  assign new_n9664 = n111 & new_n936;
  assign new_n9665 = new_n9664 ^ new_n9663;
  assign new_n9666 = new_n9665 ^ new_n9662;
  assign new_n9667 = new_n9666 ^ n18;
  assign new_n9668 = new_n9667 ^ new_n9659;
  assign new_n9669 = new_n9376 ^ new_n9364;
  assign new_n9670 = ~new_n9373 & new_n9669;
  assign new_n9671 = new_n9670 ^ new_n9376;
  assign new_n9672 = new_n9671 ^ new_n9668;
  assign new_n9673 = n115 & new_n707;
  assign new_n9674 = ~new_n7256 & new_n701;
  assign new_n9675 = new_n9674 ^ new_n9673;
  assign new_n9676 = n116 & new_n700;
  assign new_n9677 = n114 & new_n787;
  assign new_n9678 = new_n9677 ^ new_n9676;
  assign new_n9679 = new_n9678 ^ new_n9675;
  assign new_n9680 = new_n9679 ^ n15;
  assign new_n9681 = new_n9680 ^ new_n9672;
  assign new_n9682 = new_n9389 ^ new_n9377;
  assign new_n9683 = ~new_n9386 & new_n9682;
  assign new_n9684 = new_n9683 ^ new_n9389;
  assign new_n9685 = new_n9684 ^ new_n9681;
  assign new_n9686 = n118 & new_n499;
  assign new_n9687 = ~new_n506 & ~new_n8019;
  assign new_n9688 = new_n9687 ^ new_n9686;
  assign new_n9689 = ~new_n505 & n119;
  assign new_n9690 = n117 & new_n579;
  assign new_n9691 = new_n9690 ^ new_n9689;
  assign new_n9692 = new_n9691 ^ new_n9688;
  assign new_n9693 = new_n9692 ^ n12;
  assign new_n9694 = new_n9693 ^ new_n9685;
  assign new_n9695 = new_n9402 ^ new_n9390;
  assign new_n9696 = ~new_n9399 & new_n9695;
  assign new_n9697 = new_n9696 ^ new_n9402;
  assign new_n9698 = new_n9697 ^ new_n9694;
  assign new_n9699 = n124 & new_n218;
  assign new_n9700 = new_n8863 ^ n125;
  assign new_n9701 = new_n208 & new_n9700;
  assign new_n9702 = new_n9701 ^ new_n9699;
  assign new_n9703 = n125 & new_n207;
  assign new_n9704 = n123 & new_n212;
  assign new_n9705 = new_n9704 ^ new_n9703;
  assign new_n9706 = new_n9705 ^ new_n9702;
  assign new_n9707 = new_n9706 ^ n6;
  assign new_n9708 = n121 & new_n354;
  assign new_n9709 = new_n349 & new_n8850;
  assign new_n9710 = new_n9709 ^ new_n9708;
  assign new_n9711 = n122 & new_n348;
  assign new_n9712 = n120 & new_n391;
  assign new_n9713 = new_n9712 ^ new_n9711;
  assign new_n9714 = new_n9713 ^ new_n9710;
  assign new_n9715 = new_n9714 ^ n9;
  assign new_n9716 = new_n9715 ^ new_n9707;
  assign new_n9717 = new_n9716 ^ new_n9698;
  assign new_n9718 = n127 ^ n126;
  assign new_n9719 = ~n127 & n126;
  assign new_n9720 = new_n9719 ^ new_n9718;
  assign new_n9721 = ~new_n9426 & new_n9720;
  assign new_n9722 = ~new_n9427 & new_n9719;
  assign new_n9723 = new_n9722 ^ new_n9721;
  assign new_n9724 = ~new_n9723 & new_n155;
  assign new_n9725 = new_n9724 ^ n2;
  assign new_n9726 = new_n9725 ^ n128;
  assign new_n9727 = n127 ^ n3;
  assign new_n9728 = ~n126 & n3;
  assign new_n9729 = new_n9728 ^ new_n9727;
  assign new_n9730 = ~n2 & new_n9729;
  assign new_n9731 = new_n9730 ^ new_n9727;
  assign new_n9732 = new_n9731 ^ new_n9726;
  assign new_n9733 = ~n1 & new_n9732;
  assign new_n9734 = new_n9733 ^ new_n9726;
  assign new_n9735 = new_n9734 ^ new_n9717;
  assign new_n9736 = new_n9412 ^ new_n9403;
  assign new_n9737 = ~new_n9421 & new_n9736;
  assign new_n9738 = new_n9737 ^ new_n9403;
  assign new_n9739 = new_n9738 ^ new_n9735;
  assign new_n9740 = new_n9447 ^ new_n9422;
  assign new_n9741 = ~new_n9443 & new_n9740;
  assign new_n9742 = new_n9741 ^ new_n9447;
  assign new_n9743 = new_n9742 ^ new_n9739;
  assign new_n9744 = new_n9448 ^ new_n9163;
  assign new_n9745 = ~new_n9454 & ~new_n9744;
  assign new_n9746 = new_n9745 ^ new_n9163;
  assign new_n9747 = new_n9746 ^ new_n9743;
  assign new_n9748 = ~new_n6805 & n77;
  assign new_n9749 = ~new_n891 & new_n6800;
  assign new_n9750 = new_n9749 ^ new_n9748;
  assign new_n9751 = n78 & new_n6799;
  assign new_n9752 = n76 & new_n6811;
  assign new_n9753 = new_n9752 ^ new_n9751;
  assign new_n9754 = new_n9753 ^ new_n9750;
  assign new_n9755 = new_n9754 ^ n54;
  assign new_n9756 = new_n9514 ^ new_n9502;
  assign new_n9757 = ~new_n9511 & new_n9756;
  assign new_n9758 = new_n9757 ^ new_n9514;
  assign new_n9759 = new_n9758 ^ new_n9755;
  assign new_n9760 = new_n9493 & new_n9498;
  assign new_n9761 = ~new_n9494 & new_n9496;
  assign new_n9762 = ~new_n9760 & ~new_n9761;
  assign new_n9763 = n68 & new_n9195;
  assign new_n9764 = ~new_n304 & new_n9185;
  assign new_n9765 = new_n9764 ^ new_n9763;
  assign new_n9766 = n69 & new_n9184;
  assign new_n9767 = n67 & new_n9189;
  assign new_n9768 = new_n9767 ^ new_n9766;
  assign new_n9769 = new_n9768 ^ new_n9765;
  assign new_n9770 = new_n9769 ^ n63;
  assign new_n9771 = n64 & n65;
  assign new_n9772 = new_n9771 ^ n66;
  assign new_n9773 = ~new_n9495 & new_n9772;
  assign new_n9774 = new_n9773 ^ n66;
  assign new_n9775 = new_n9774 ^ new_n9770;
  assign new_n9776 = new_n9775 ^ new_n9762;
  assign new_n9777 = n71 & new_n8355;
  assign new_n9778 = ~new_n459 & new_n8345;
  assign new_n9779 = new_n9778 ^ new_n9777;
  assign new_n9780 = n72 & new_n8344;
  assign new_n9781 = n70 & new_n8349;
  assign new_n9782 = new_n9781 ^ new_n9780;
  assign new_n9783 = new_n9782 ^ new_n9779;
  assign new_n9784 = new_n9783 ^ n60;
  assign new_n9785 = new_n9784 ^ new_n9776;
  assign new_n9786 = new_n9499 ^ new_n9478;
  assign new_n9787 = new_n9500 & new_n9786;
  assign new_n9788 = new_n9787 ^ new_n9478;
  assign new_n9789 = new_n9788 ^ new_n9785;
  assign new_n9790 = n74 & new_n7553;
  assign new_n9791 = new_n660 & new_n7543;
  assign new_n9792 = new_n9791 ^ new_n9790;
  assign new_n9793 = n75 & new_n7542;
  assign new_n9794 = n73 & new_n7547;
  assign new_n9795 = new_n9794 ^ new_n9793;
  assign new_n9796 = new_n9795 ^ new_n9792;
  assign new_n9797 = new_n9796 ^ n57;
  assign new_n9798 = new_n9797 ^ new_n9789;
  assign new_n9799 = new_n9501 ^ new_n9463;
  assign new_n9800 = ~new_n9799 & new_n9467;
  assign new_n9801 = new_n9800 ^ new_n9466;
  assign new_n9802 = new_n9801 ^ new_n9798;
  assign new_n9803 = new_n9802 ^ new_n9759;
  assign new_n9804 = ~new_n6110 & n80;
  assign new_n9805 = new_n1161 & new_n6105;
  assign new_n9806 = new_n9805 ^ new_n9804;
  assign new_n9807 = n81 & new_n6104;
  assign new_n9808 = n79 & new_n6347;
  assign new_n9809 = new_n9808 ^ new_n9807;
  assign new_n9810 = new_n9809 ^ new_n9806;
  assign new_n9811 = new_n9810 ^ n51;
  assign new_n9812 = new_n9811 ^ new_n9803;
  assign new_n9813 = new_n9528 ^ new_n9515;
  assign new_n9814 = ~new_n9813 & new_n9520;
  assign new_n9815 = new_n9814 ^ new_n9519;
  assign new_n9816 = new_n9815 ^ new_n9812;
  assign new_n9817 = ~new_n5424 & n83;
  assign new_n9818 = new_n1468 & new_n5419;
  assign new_n9819 = new_n9818 ^ new_n9817;
  assign new_n9820 = n84 & new_n5418;
  assign new_n9821 = n82 & new_n5648;
  assign new_n9822 = new_n9821 ^ new_n9820;
  assign new_n9823 = new_n9822 ^ new_n9819;
  assign new_n9824 = new_n9823 ^ n48;
  assign new_n9825 = new_n9824 ^ new_n9816;
  assign new_n9826 = new_n9541 ^ new_n9529;
  assign new_n9827 = ~new_n9538 & ~new_n9826;
  assign new_n9828 = new_n9827 ^ new_n9541;
  assign new_n9829 = new_n9828 ^ new_n9825;
  assign new_n9830 = ~new_n4804 & n86;
  assign new_n9831 = new_n1811 & new_n4799;
  assign new_n9832 = new_n9831 ^ new_n9830;
  assign new_n9833 = n85 & new_n4810;
  assign new_n9834 = n87 & new_n4798;
  assign new_n9835 = new_n9834 ^ new_n9833;
  assign new_n9836 = new_n9835 ^ new_n9832;
  assign new_n9837 = new_n9836 ^ n45;
  assign new_n9838 = new_n9837 ^ new_n9829;
  assign new_n9839 = new_n9554 ^ new_n9542;
  assign new_n9840 = ~new_n9839 & new_n9551;
  assign new_n9841 = new_n9840 ^ new_n9554;
  assign new_n9842 = new_n9841 ^ new_n9838;
  assign new_n9843 = ~new_n4212 & n89;
  assign new_n9844 = new_n2193 & new_n4201;
  assign new_n9845 = new_n9844 ^ new_n9843;
  assign new_n9846 = n90 & new_n4200;
  assign new_n9847 = n88 & new_n4206;
  assign new_n9848 = new_n9847 ^ new_n9846;
  assign new_n9849 = new_n9848 ^ new_n9845;
  assign new_n9850 = new_n9849 ^ n42;
  assign new_n9851 = new_n9850 ^ new_n9842;
  assign new_n9852 = new_n9567 ^ new_n9555;
  assign new_n9853 = ~new_n9852 & new_n9564;
  assign new_n9854 = new_n9853 ^ new_n9567;
  assign new_n9855 = new_n9854 ^ new_n9851;
  assign new_n9856 = ~new_n3682 & n92;
  assign new_n9857 = new_n2628 & new_n3677;
  assign new_n9858 = new_n9857 ^ new_n9856;
  assign new_n9859 = n93 & new_n3676;
  assign new_n9860 = n91 & new_n3688;
  assign new_n9861 = new_n9860 ^ new_n9859;
  assign new_n9862 = new_n9861 ^ new_n9858;
  assign new_n9863 = new_n9862 ^ n39;
  assign new_n9864 = new_n9863 ^ new_n9855;
  assign new_n9865 = new_n9580 ^ new_n9568;
  assign new_n9866 = ~new_n9865 & new_n9577;
  assign new_n9867 = new_n9866 ^ new_n9580;
  assign new_n9868 = new_n9867 ^ new_n9864;
  assign new_n9869 = ~new_n3143 & n95;
  assign new_n9870 = new_n3095 & new_n3138;
  assign new_n9871 = new_n9870 ^ new_n9869;
  assign new_n9872 = n96 & new_n3137;
  assign new_n9873 = n94 & new_n3149;
  assign new_n9874 = new_n9873 ^ new_n9872;
  assign new_n9875 = new_n9874 ^ new_n9871;
  assign new_n9876 = new_n9875 ^ n36;
  assign new_n9877 = new_n9876 ^ new_n9868;
  assign new_n9878 = new_n9593 ^ new_n9581;
  assign new_n9879 = ~new_n9878 & new_n9590;
  assign new_n9880 = new_n9879 ^ new_n9593;
  assign new_n9881 = new_n9880 ^ new_n9877;
  assign new_n9882 = ~new_n2672 & n98;
  assign new_n9883 = new_n2667 & new_n3604;
  assign new_n9884 = new_n9883 ^ new_n9882;
  assign new_n9885 = n99 & new_n2666;
  assign new_n9886 = n97 & new_n2664;
  assign new_n9887 = new_n9886 ^ new_n9885;
  assign new_n9888 = new_n9887 ^ new_n9884;
  assign new_n9889 = new_n9888 ^ n33;
  assign new_n9890 = new_n9889 ^ new_n9881;
  assign new_n9891 = new_n9606 ^ new_n9594;
  assign new_n9892 = new_n9603 & new_n9891;
  assign new_n9893 = new_n9892 ^ new_n9606;
  assign new_n9894 = new_n9893 ^ new_n9890;
  assign new_n9895 = n101 & new_n2246;
  assign new_n9896 = new_n2241 & new_n4159;
  assign new_n9897 = new_n9896 ^ new_n9895;
  assign new_n9898 = n102 & new_n2240;
  assign new_n9899 = n100 & new_n2391;
  assign new_n9900 = new_n9899 ^ new_n9898;
  assign new_n9901 = new_n9900 ^ new_n9897;
  assign new_n9902 = new_n9901 ^ n30;
  assign new_n9903 = new_n9902 ^ new_n9894;
  assign new_n9904 = new_n9619 ^ new_n9607;
  assign new_n9905 = ~new_n9616 & new_n9904;
  assign new_n9906 = new_n9905 ^ new_n9619;
  assign new_n9907 = new_n9906 ^ new_n9903;
  assign new_n9908 = n104 & new_n1874;
  assign new_n9909 = ~new_n4754 & new_n1864;
  assign new_n9910 = new_n9909 ^ new_n9908;
  assign new_n9911 = n105 & new_n1863;
  assign new_n9912 = n103 & new_n1868;
  assign new_n9913 = new_n9912 ^ new_n9911;
  assign new_n9914 = new_n9913 ^ new_n9910;
  assign new_n9915 = new_n9914 ^ n27;
  assign new_n9916 = new_n9915 ^ new_n9907;
  assign new_n9917 = new_n9632 ^ new_n9620;
  assign new_n9918 = ~new_n9629 & new_n9917;
  assign new_n9919 = new_n9918 ^ new_n9632;
  assign new_n9920 = new_n9919 ^ new_n9916;
  assign new_n9921 = ~new_n1506 & n107;
  assign new_n9922 = ~new_n5377 & new_n1501;
  assign new_n9923 = new_n9922 ^ new_n9921;
  assign new_n9924 = n108 & new_n1500;
  assign new_n9925 = n106 & new_n1512;
  assign new_n9926 = new_n9925 ^ new_n9924;
  assign new_n9927 = new_n9926 ^ new_n9923;
  assign new_n9928 = new_n9927 ^ n24;
  assign new_n9929 = new_n9928 ^ new_n9920;
  assign new_n9930 = new_n9645 ^ new_n9633;
  assign new_n9931 = ~new_n9642 & new_n9930;
  assign new_n9932 = new_n9931 ^ new_n9645;
  assign new_n9933 = new_n9932 ^ new_n9929;
  assign new_n9934 = ~new_n1198 & n110;
  assign new_n9935 = new_n1193 & new_n6049;
  assign new_n9936 = new_n9935 ^ new_n9934;
  assign new_n9937 = n111 & new_n1192;
  assign new_n9938 = n109 & new_n1204;
  assign new_n9939 = new_n9938 ^ new_n9937;
  assign new_n9940 = new_n9939 ^ new_n9936;
  assign new_n9941 = new_n9940 ^ n21;
  assign new_n9942 = new_n9941 ^ new_n9933;
  assign new_n9943 = new_n9658 ^ new_n9646;
  assign new_n9944 = ~new_n9655 & new_n9943;
  assign new_n9945 = new_n9944 ^ new_n9658;
  assign new_n9946 = new_n9945 ^ new_n9942;
  assign new_n9947 = ~new_n930 & n113;
  assign new_n9948 = ~new_n6764 & new_n925;
  assign new_n9949 = new_n9948 ^ new_n9947;
  assign new_n9950 = n114 & new_n924;
  assign new_n9951 = n112 & new_n936;
  assign new_n9952 = new_n9951 ^ new_n9950;
  assign new_n9953 = new_n9952 ^ new_n9949;
  assign new_n9954 = new_n9953 ^ n18;
  assign new_n9955 = new_n9954 ^ new_n9946;
  assign new_n9956 = new_n9671 ^ new_n9659;
  assign new_n9957 = ~new_n9668 & new_n9956;
  assign new_n9958 = new_n9957 ^ new_n9671;
  assign new_n9959 = new_n9958 ^ new_n9955;
  assign new_n9960 = n116 & new_n707;
  assign new_n9961 = ~new_n7503 & new_n701;
  assign new_n9962 = new_n9961 ^ new_n9960;
  assign new_n9963 = n117 & new_n700;
  assign new_n9964 = n115 & new_n787;
  assign new_n9965 = new_n9964 ^ new_n9963;
  assign new_n9966 = new_n9965 ^ new_n9962;
  assign new_n9967 = new_n9966 ^ n15;
  assign new_n9968 = new_n9967 ^ new_n9959;
  assign new_n9969 = new_n9684 ^ new_n9672;
  assign new_n9970 = ~new_n9681 & new_n9969;
  assign new_n9971 = new_n9970 ^ new_n9684;
  assign new_n9972 = new_n9971 ^ new_n9968;
  assign new_n9973 = n119 & new_n499;
  assign new_n9974 = ~new_n506 & new_n8286;
  assign new_n9975 = new_n9974 ^ new_n9973;
  assign new_n9976 = ~new_n505 & n120;
  assign new_n9977 = n118 & new_n579;
  assign new_n9978 = new_n9977 ^ new_n9976;
  assign new_n9979 = new_n9978 ^ new_n9975;
  assign new_n9980 = new_n9979 ^ n12;
  assign new_n9981 = new_n9980 ^ new_n9972;
  assign new_n9982 = new_n9697 ^ new_n9685;
  assign new_n9983 = ~new_n9694 & new_n9982;
  assign new_n9984 = new_n9983 ^ new_n9697;
  assign new_n9985 = new_n9984 ^ new_n9981;
  assign new_n9986 = n125 & new_n218;
  assign new_n9987 = new_n9423 ^ new_n9140;
  assign new_n9988 = new_n208 & new_n9987;
  assign new_n9989 = new_n9988 ^ new_n9986;
  assign new_n9990 = n126 & new_n207;
  assign new_n9991 = n124 & new_n212;
  assign new_n9992 = new_n9991 ^ new_n9990;
  assign new_n9993 = new_n9992 ^ new_n9989;
  assign new_n9994 = new_n9993 ^ n6;
  assign new_n9995 = n122 & new_n354;
  assign new_n9996 = ~new_n9116 & new_n349;
  assign new_n9997 = new_n9996 ^ new_n9995;
  assign new_n9998 = n123 & new_n348;
  assign new_n9999 = n121 & new_n391;
  assign new_n10000 = new_n9999 ^ new_n9998;
  assign new_n10001 = new_n10000 ^ new_n9997;
  assign new_n10002 = new_n10001 ^ n9;
  assign new_n10003 = new_n10002 ^ new_n9994;
  assign new_n10004 = new_n10003 ^ new_n9985;
  assign new_n10005 = ~n127 & n128;
  assign new_n10006 = n128 ^ n127;
  assign new_n10007 = new_n10006 ^ new_n10005;
  assign new_n10008 = ~new_n9721 & new_n10007;
  assign new_n10009 = ~new_n9722 & new_n10005;
  assign new_n10010 = new_n10009 ^ new_n10008;
  assign new_n10011 = ~new_n10010 & new_n155;
  assign new_n10012 = new_n10011 ^ n2;
  assign new_n10013 = ~n3 & ~new_n10006;
  assign new_n10014 = new_n10013 ^ n127;
  assign new_n10015 = ~new_n10014 & new_n155;
  assign new_n10016 = new_n10015 ^ new_n10012;
  assign new_n10017 = ~n1 & new_n10016;
  assign new_n10018 = new_n10017 ^ new_n10012;
  assign new_n10019 = n2 & n3;
  assign new_n10020 = new_n10019 ^ n127;
  assign new_n10021 = new_n10020 ^ new_n10019;
  assign new_n10022 = new_n10019 ^ n3;
  assign new_n10023 = ~new_n10021 & new_n10022;
  assign new_n10024 = new_n10023 ^ new_n10019;
  assign new_n10025 = ~n128 & new_n10024;
  assign new_n10026 = ~new_n10018 & ~new_n10025;
  assign new_n10027 = new_n10026 ^ new_n10004;
  assign new_n10028 = new_n9707 ^ new_n9698;
  assign new_n10029 = ~new_n9716 & new_n10028;
  assign new_n10030 = new_n10029 ^ new_n9698;
  assign new_n10031 = new_n10030 ^ new_n10027;
  assign new_n10032 = new_n9738 ^ new_n9734;
  assign new_n10033 = ~new_n10032 & new_n9735;
  assign new_n10034 = new_n10033 ^ new_n9717;
  assign new_n10035 = new_n10034 ^ new_n10031;
  assign new_n10036 = new_n9746 ^ new_n9742;
  assign new_n10037 = ~new_n9743 & ~new_n10036;
  assign new_n10038 = new_n10037 ^ new_n9746;
  assign new_n10039 = new_n10038 ^ new_n10035;
  assign new_n10040 = new_n9994 ^ new_n9985;
  assign new_n10041 = ~new_n10003 & new_n10040;
  assign new_n10042 = new_n10041 ^ new_n9985;
  assign new_n10043 = ~n3 & new_n155;
  assign new_n10044 = ~n1 & new_n10043;
  assign new_n10045 = new_n10044 ^ new_n155;
  assign new_n10046 = n3 & new_n155;
  assign new_n10047 = ~n1 & new_n10046;
  assign new_n10048 = new_n10047 ^ new_n155;
  assign new_n10049 = new_n10048 ^ new_n155;
  assign new_n10050 = new_n10049 ^ new_n10045;
  assign new_n10051 = new_n10045 ^ new_n10009;
  assign new_n10052 = new_n10051 ^ new_n10045;
  assign new_n10053 = new_n10050 & new_n10052;
  assign new_n10054 = new_n10053 ^ new_n10045;
  assign new_n10055 = n128 & new_n10054;
  assign new_n10056 = new_n10055 ^ new_n155;
  assign new_n10057 = new_n10056 ^ new_n155;
  assign new_n10058 = new_n10057 ^ n3;
  assign new_n10059 = new_n10058 ^ new_n10042;
  assign new_n10060 = ~new_n6805 & n78;
  assign new_n10061 = ~new_n982 & new_n6800;
  assign new_n10062 = new_n10061 ^ new_n10060;
  assign new_n10063 = n79 & new_n6799;
  assign new_n10064 = n77 & new_n6811;
  assign new_n10065 = new_n10064 ^ new_n10063;
  assign new_n10066 = new_n10065 ^ new_n10062;
  assign new_n10067 = new_n10066 ^ n54;
  assign new_n10068 = new_n9802 ^ new_n9755;
  assign new_n10069 = ~new_n10068 & new_n9759;
  assign new_n10070 = new_n10069 ^ new_n9758;
  assign new_n10071 = new_n10070 ^ new_n10067;
  assign new_n10072 = n75 & new_n7553;
  assign new_n10073 = ~new_n737 & new_n7543;
  assign new_n10074 = new_n10073 ^ new_n10072;
  assign new_n10075 = n76 & new_n7542;
  assign new_n10076 = n74 & new_n7547;
  assign new_n10077 = new_n10076 ^ new_n10075;
  assign new_n10078 = new_n10077 ^ new_n10074;
  assign new_n10079 = new_n10078 ^ n57;
  assign new_n10080 = new_n9801 ^ new_n9789;
  assign new_n10081 = ~new_n9798 & new_n10080;
  assign new_n10082 = new_n10081 ^ new_n9801;
  assign new_n10083 = new_n10082 ^ new_n10079;
  assign new_n10084 = n64 & n66;
  assign new_n10085 = new_n10084 ^ n67;
  assign new_n10086 = ~new_n9495 & new_n10085;
  assign new_n10087 = new_n10086 ^ n67;
  assign new_n10088 = new_n9770 ^ new_n9762;
  assign new_n10089 = ~new_n9775 & ~new_n10088;
  assign new_n10090 = new_n10089 ^ new_n9762;
  assign new_n10091 = new_n10090 ^ new_n10087;
  assign new_n10092 = n69 & new_n9195;
  assign new_n10093 = ~new_n339 & new_n9185;
  assign new_n10094 = new_n10093 ^ new_n10092;
  assign new_n10095 = n70 & new_n9184;
  assign new_n10096 = n68 & new_n9189;
  assign new_n10097 = new_n10096 ^ new_n10095;
  assign new_n10098 = new_n10097 ^ new_n10094;
  assign new_n10099 = new_n10098 ^ n63;
  assign new_n10100 = new_n10099 ^ new_n10091;
  assign new_n10101 = n72 & new_n8355;
  assign new_n10102 = new_n534 & new_n8345;
  assign new_n10103 = new_n10102 ^ new_n10101;
  assign new_n10104 = n73 & new_n8344;
  assign new_n10105 = n71 & new_n8349;
  assign new_n10106 = new_n10105 ^ new_n10104;
  assign new_n10107 = new_n10106 ^ new_n10103;
  assign new_n10108 = new_n10107 ^ n60;
  assign new_n10109 = new_n10108 ^ new_n10100;
  assign new_n10110 = new_n9788 ^ new_n9776;
  assign new_n10111 = new_n9785 & new_n10110;
  assign new_n10112 = new_n10111 ^ new_n9788;
  assign new_n10113 = new_n10112 ^ new_n10109;
  assign new_n10114 = new_n10113 ^ new_n10083;
  assign new_n10115 = new_n10114 ^ new_n10071;
  assign new_n10116 = ~new_n6110 & n81;
  assign new_n10117 = new_n1263 & new_n6105;
  assign new_n10118 = new_n10117 ^ new_n10116;
  assign new_n10119 = n82 & new_n6104;
  assign new_n10120 = n80 & new_n6347;
  assign new_n10121 = new_n10120 ^ new_n10119;
  assign new_n10122 = new_n10121 ^ new_n10118;
  assign new_n10123 = new_n10122 ^ n51;
  assign new_n10124 = new_n10123 ^ new_n10115;
  assign new_n10125 = new_n9815 ^ new_n9803;
  assign new_n10126 = ~new_n9812 & new_n10125;
  assign new_n10127 = new_n10126 ^ new_n9815;
  assign new_n10128 = new_n10127 ^ new_n10124;
  assign new_n10129 = ~new_n5424 & n84;
  assign new_n10130 = new_n1584 & new_n5419;
  assign new_n10131 = new_n10130 ^ new_n10129;
  assign new_n10132 = n85 & new_n5418;
  assign new_n10133 = n83 & new_n5648;
  assign new_n10134 = new_n10133 ^ new_n10132;
  assign new_n10135 = new_n10134 ^ new_n10131;
  assign new_n10136 = new_n10135 ^ n48;
  assign new_n10137 = new_n10136 ^ new_n10128;
  assign new_n10138 = new_n9828 ^ new_n9816;
  assign new_n10139 = ~new_n9825 & ~new_n10138;
  assign new_n10140 = new_n10139 ^ new_n9828;
  assign new_n10141 = new_n10140 ^ new_n10137;
  assign new_n10142 = ~new_n4804 & n87;
  assign new_n10143 = new_n1940 & new_n4799;
  assign new_n10144 = new_n10143 ^ new_n10142;
  assign new_n10145 = n88 & new_n4798;
  assign new_n10146 = n86 & new_n4810;
  assign new_n10147 = new_n10146 ^ new_n10145;
  assign new_n10148 = new_n10147 ^ new_n10144;
  assign new_n10149 = new_n10148 ^ n45;
  assign new_n10150 = new_n10149 ^ new_n10141;
  assign new_n10151 = new_n9841 ^ new_n9829;
  assign new_n10152 = ~new_n10151 & new_n9838;
  assign new_n10153 = new_n10152 ^ new_n9841;
  assign new_n10154 = new_n10153 ^ new_n10150;
  assign new_n10155 = ~new_n4212 & n90;
  assign new_n10156 = new_n2341 & new_n4201;
  assign new_n10157 = new_n10156 ^ new_n10155;
  assign new_n10158 = n91 & new_n4200;
  assign new_n10159 = n89 & new_n4206;
  assign new_n10160 = new_n10159 ^ new_n10158;
  assign new_n10161 = new_n10160 ^ new_n10157;
  assign new_n10162 = new_n10161 ^ n42;
  assign new_n10163 = new_n10162 ^ new_n10154;
  assign new_n10164 = new_n9854 ^ new_n9842;
  assign new_n10165 = ~new_n10164 & new_n9851;
  assign new_n10166 = new_n10165 ^ new_n9854;
  assign new_n10167 = new_n10166 ^ new_n10163;
  assign new_n10168 = ~new_n3682 & n93;
  assign new_n10169 = new_n2785 & new_n3677;
  assign new_n10170 = new_n10169 ^ new_n10168;
  assign new_n10171 = n94 & new_n3676;
  assign new_n10172 = n92 & new_n3688;
  assign new_n10173 = new_n10172 ^ new_n10171;
  assign new_n10174 = new_n10173 ^ new_n10170;
  assign new_n10175 = new_n10174 ^ n39;
  assign new_n10176 = new_n10175 ^ new_n10167;
  assign new_n10177 = new_n9867 ^ new_n9855;
  assign new_n10178 = ~new_n10177 & new_n9864;
  assign new_n10179 = new_n10178 ^ new_n9867;
  assign new_n10180 = new_n10179 ^ new_n10176;
  assign new_n10181 = ~new_n3143 & n96;
  assign new_n10182 = new_n3138 & new_n3273;
  assign new_n10183 = new_n10182 ^ new_n10181;
  assign new_n10184 = n97 & new_n3137;
  assign new_n10185 = n95 & new_n3149;
  assign new_n10186 = new_n10185 ^ new_n10184;
  assign new_n10187 = new_n10186 ^ new_n10183;
  assign new_n10188 = new_n10187 ^ n36;
  assign new_n10189 = new_n10188 ^ new_n10180;
  assign new_n10190 = new_n9880 ^ new_n9868;
  assign new_n10191 = ~new_n10190 & new_n9877;
  assign new_n10192 = new_n10191 ^ new_n9880;
  assign new_n10193 = new_n10192 ^ new_n10189;
  assign new_n10194 = ~new_n2672 & n99;
  assign new_n10195 = new_n2667 & new_n3789;
  assign new_n10196 = new_n10195 ^ new_n10194;
  assign new_n10197 = n100 & new_n2666;
  assign new_n10198 = n98 & new_n2664;
  assign new_n10199 = new_n10198 ^ new_n10197;
  assign new_n10200 = new_n10199 ^ new_n10196;
  assign new_n10201 = new_n10200 ^ n33;
  assign new_n10202 = new_n10201 ^ new_n10193;
  assign new_n10203 = new_n9893 ^ new_n9881;
  assign new_n10204 = new_n9890 & new_n10203;
  assign new_n10205 = new_n10204 ^ new_n9893;
  assign new_n10206 = new_n10205 ^ new_n10202;
  assign new_n10207 = n102 & new_n2246;
  assign new_n10208 = new_n2241 & new_n4368;
  assign new_n10209 = new_n10208 ^ new_n10207;
  assign new_n10210 = n103 & new_n2240;
  assign new_n10211 = n101 & new_n2391;
  assign new_n10212 = new_n10211 ^ new_n10210;
  assign new_n10213 = new_n10212 ^ new_n10209;
  assign new_n10214 = new_n10213 ^ n30;
  assign new_n10215 = new_n10214 ^ new_n10206;
  assign new_n10216 = new_n9906 ^ new_n9894;
  assign new_n10217 = ~new_n9903 & new_n10216;
  assign new_n10218 = new_n10217 ^ new_n9906;
  assign new_n10219 = new_n10218 ^ new_n10215;
  assign new_n10220 = n105 & new_n1874;
  assign new_n10221 = ~new_n4961 & new_n1864;
  assign new_n10222 = new_n10221 ^ new_n10220;
  assign new_n10223 = n106 & new_n1863;
  assign new_n10224 = n104 & new_n1868;
  assign new_n10225 = new_n10224 ^ new_n10223;
  assign new_n10226 = new_n10225 ^ new_n10222;
  assign new_n10227 = new_n10226 ^ n27;
  assign new_n10228 = new_n10227 ^ new_n10219;
  assign new_n10229 = new_n9919 ^ new_n9907;
  assign new_n10230 = ~new_n9916 & new_n10229;
  assign new_n10231 = new_n10230 ^ new_n9919;
  assign new_n10232 = new_n10231 ^ new_n10228;
  assign new_n10233 = ~new_n1506 & n108;
  assign new_n10234 = new_n1501 & new_n5604;
  assign new_n10235 = new_n10234 ^ new_n10233;
  assign new_n10236 = n109 & new_n1500;
  assign new_n10237 = n107 & new_n1512;
  assign new_n10238 = new_n10237 ^ new_n10236;
  assign new_n10239 = new_n10238 ^ new_n10235;
  assign new_n10240 = new_n10239 ^ n24;
  assign new_n10241 = new_n10240 ^ new_n10232;
  assign new_n10242 = new_n9932 ^ new_n9920;
  assign new_n10243 = ~new_n9929 & new_n10242;
  assign new_n10244 = new_n10243 ^ new_n9932;
  assign new_n10245 = new_n10244 ^ new_n10241;
  assign new_n10246 = ~new_n1198 & n111;
  assign new_n10247 = ~new_n6284 & new_n1193;
  assign new_n10248 = new_n10247 ^ new_n10246;
  assign new_n10249 = n112 & new_n1192;
  assign new_n10250 = n110 & new_n1204;
  assign new_n10251 = new_n10250 ^ new_n10249;
  assign new_n10252 = new_n10251 ^ new_n10248;
  assign new_n10253 = new_n10252 ^ n21;
  assign new_n10254 = new_n10253 ^ new_n10245;
  assign new_n10255 = new_n9945 ^ new_n9933;
  assign new_n10256 = ~new_n9942 & new_n10255;
  assign new_n10257 = new_n10256 ^ new_n9945;
  assign new_n10258 = new_n10257 ^ new_n10254;
  assign new_n10259 = ~new_n930 & n114;
  assign new_n10260 = ~new_n7013 & new_n925;
  assign new_n10261 = new_n10260 ^ new_n10259;
  assign new_n10262 = n115 & new_n924;
  assign new_n10263 = n113 & new_n936;
  assign new_n10264 = new_n10263 ^ new_n10262;
  assign new_n10265 = new_n10264 ^ new_n10261;
  assign new_n10266 = new_n10265 ^ n18;
  assign new_n10267 = new_n10266 ^ new_n10258;
  assign new_n10268 = new_n9958 ^ new_n9946;
  assign new_n10269 = ~new_n9955 & new_n10268;
  assign new_n10270 = new_n10269 ^ new_n9958;
  assign new_n10271 = new_n10270 ^ new_n10267;
  assign new_n10272 = n117 & new_n707;
  assign new_n10273 = ~new_n7761 & new_n701;
  assign new_n10274 = new_n10273 ^ new_n10272;
  assign new_n10275 = n118 & new_n700;
  assign new_n10276 = n116 & new_n787;
  assign new_n10277 = new_n10276 ^ new_n10275;
  assign new_n10278 = new_n10277 ^ new_n10274;
  assign new_n10279 = new_n10278 ^ n15;
  assign new_n10280 = new_n10279 ^ new_n10271;
  assign new_n10281 = new_n9971 ^ new_n9959;
  assign new_n10282 = ~new_n9968 & new_n10281;
  assign new_n10283 = new_n10282 ^ new_n9971;
  assign new_n10284 = new_n10283 ^ new_n10280;
  assign new_n10285 = n123 & new_n354;
  assign new_n10286 = ~new_n9405 & new_n349;
  assign new_n10287 = new_n10286 ^ new_n10285;
  assign new_n10288 = n124 & new_n348;
  assign new_n10289 = n122 & new_n391;
  assign new_n10290 = new_n10289 ^ new_n10288;
  assign new_n10291 = new_n10290 ^ new_n10287;
  assign new_n10292 = new_n10291 ^ n9;
  assign new_n10293 = n120 & new_n499;
  assign new_n10294 = ~new_n506 & new_n8560;
  assign new_n10295 = new_n10294 ^ new_n10293;
  assign new_n10296 = ~new_n505 & n121;
  assign new_n10297 = n119 & new_n579;
  assign new_n10298 = new_n10297 ^ new_n10296;
  assign new_n10299 = new_n10298 ^ new_n10295;
  assign new_n10300 = new_n10299 ^ n12;
  assign new_n10301 = new_n10300 ^ new_n10292;
  assign new_n10302 = new_n10301 ^ new_n10284;
  assign new_n10303 = n126 & new_n218;
  assign new_n10304 = new_n9428 ^ n127;
  assign new_n10305 = new_n208 & new_n10304;
  assign new_n10306 = new_n10305 ^ new_n10303;
  assign new_n10307 = n127 & new_n207;
  assign new_n10308 = n125 & new_n212;
  assign new_n10309 = new_n10308 ^ new_n10307;
  assign new_n10310 = new_n10309 ^ new_n10306;
  assign new_n10311 = new_n10310 ^ n6;
  assign new_n10312 = new_n10311 ^ new_n10302;
  assign new_n10313 = new_n9984 ^ new_n9972;
  assign new_n10314 = ~new_n9981 & new_n10313;
  assign new_n10315 = new_n10314 ^ new_n9984;
  assign new_n10316 = new_n10315 ^ new_n10312;
  assign new_n10317 = new_n10316 ^ new_n10059;
  assign new_n10318 = new_n10030 ^ new_n10026;
  assign new_n10319 = ~new_n10027 & new_n10318;
  assign new_n10320 = new_n10319 ^ new_n10004;
  assign new_n10321 = new_n10320 ^ new_n10317;
  assign new_n10322 = new_n10038 ^ new_n10031;
  assign new_n10323 = new_n10035 & new_n10322;
  assign new_n10324 = new_n10323 ^ new_n10038;
  assign new_n10325 = new_n10324 ^ new_n10321;
  assign new_n10326 = n73 & new_n8355;
  assign new_n10327 = new_n595 & new_n8345;
  assign new_n10328 = new_n10327 ^ new_n10326;
  assign new_n10329 = n74 & new_n8344;
  assign new_n10330 = n72 & new_n8349;
  assign new_n10331 = new_n10330 ^ new_n10329;
  assign new_n10332 = new_n10331 ^ new_n10328;
  assign new_n10333 = new_n10332 ^ n60;
  assign new_n10334 = n70 & new_n9195;
  assign new_n10335 = ~new_n402 & new_n9185;
  assign new_n10336 = new_n10335 ^ new_n10334;
  assign new_n10337 = n71 & new_n9184;
  assign new_n10338 = n69 & new_n9189;
  assign new_n10339 = new_n10338 ^ new_n10337;
  assign new_n10340 = new_n10339 ^ new_n10336;
  assign new_n10341 = n64 & n68;
  assign new_n10342 = n68 ^ n67;
  assign new_n10343 = ~n64 & new_n10342;
  assign new_n10344 = new_n10343 ^ n67;
  assign new_n10345 = new_n10344 ^ new_n10341;
  assign new_n10346 = ~n63 & ~new_n10345;
  assign new_n10347 = new_n10346 ^ new_n10344;
  assign new_n10348 = new_n10347 ^ n3;
  assign new_n10349 = new_n10348 ^ new_n10340;
  assign new_n10350 = new_n10349 ^ new_n10333;
  assign new_n10351 = new_n10099 ^ new_n10087;
  assign new_n10352 = ~new_n10091 & ~new_n10351;
  assign new_n10353 = new_n10352 ^ new_n10090;
  assign new_n10354 = new_n10353 ^ new_n10350;
  assign new_n10355 = n76 & new_n7553;
  assign new_n10356 = ~new_n812 & new_n7543;
  assign new_n10357 = new_n10356 ^ new_n10355;
  assign new_n10358 = n77 & new_n7542;
  assign new_n10359 = n75 & new_n7547;
  assign new_n10360 = new_n10359 ^ new_n10358;
  assign new_n10361 = new_n10360 ^ new_n10357;
  assign new_n10362 = new_n10361 ^ n57;
  assign new_n10363 = new_n10362 ^ new_n10354;
  assign new_n10364 = new_n10112 ^ new_n10100;
  assign new_n10365 = new_n10109 & new_n10364;
  assign new_n10366 = new_n10365 ^ new_n10112;
  assign new_n10367 = new_n10366 ^ new_n10363;
  assign new_n10368 = ~new_n6805 & n79;
  assign new_n10369 = new_n1069 & new_n6800;
  assign new_n10370 = new_n10369 ^ new_n10368;
  assign new_n10371 = n80 & new_n6799;
  assign new_n10372 = n78 & new_n6811;
  assign new_n10373 = new_n10372 ^ new_n10371;
  assign new_n10374 = new_n10373 ^ new_n10370;
  assign new_n10375 = new_n10374 ^ n54;
  assign new_n10376 = new_n10375 ^ new_n10367;
  assign new_n10377 = new_n10113 ^ new_n10079;
  assign new_n10378 = ~new_n10377 & new_n10083;
  assign new_n10379 = new_n10378 ^ new_n10082;
  assign new_n10380 = new_n10379 ^ new_n10376;
  assign new_n10381 = ~new_n6110 & n82;
  assign new_n10382 = new_n1363 & new_n6105;
  assign new_n10383 = new_n10382 ^ new_n10381;
  assign new_n10384 = n83 & new_n6104;
  assign new_n10385 = n81 & new_n6347;
  assign new_n10386 = new_n10385 ^ new_n10384;
  assign new_n10387 = new_n10386 ^ new_n10383;
  assign new_n10388 = new_n10387 ^ n51;
  assign new_n10389 = new_n10388 ^ new_n10380;
  assign new_n10390 = new_n10114 ^ new_n10067;
  assign new_n10391 = ~new_n10390 & new_n10071;
  assign new_n10392 = new_n10391 ^ new_n10070;
  assign new_n10393 = new_n10392 ^ new_n10389;
  assign new_n10394 = ~new_n5424 & n85;
  assign new_n10395 = new_n1694 & new_n5419;
  assign new_n10396 = new_n10395 ^ new_n10394;
  assign new_n10397 = n86 & new_n5418;
  assign new_n10398 = n84 & new_n5648;
  assign new_n10399 = new_n10398 ^ new_n10397;
  assign new_n10400 = new_n10399 ^ new_n10396;
  assign new_n10401 = new_n10400 ^ n48;
  assign new_n10402 = new_n10401 ^ new_n10393;
  assign new_n10403 = new_n10127 ^ new_n10115;
  assign new_n10404 = ~new_n10124 & new_n10403;
  assign new_n10405 = new_n10404 ^ new_n10127;
  assign new_n10406 = new_n10405 ^ new_n10402;
  assign new_n10407 = ~new_n4804 & n88;
  assign new_n10408 = new_n2063 & new_n4799;
  assign new_n10409 = new_n10408 ^ new_n10407;
  assign new_n10410 = n89 & new_n4798;
  assign new_n10411 = n87 & new_n4810;
  assign new_n10412 = new_n10411 ^ new_n10410;
  assign new_n10413 = new_n10412 ^ new_n10409;
  assign new_n10414 = new_n10413 ^ n45;
  assign new_n10415 = new_n10414 ^ new_n10406;
  assign new_n10416 = new_n10140 ^ new_n10128;
  assign new_n10417 = ~new_n10137 & ~new_n10416;
  assign new_n10418 = new_n10417 ^ new_n10140;
  assign new_n10419 = new_n10418 ^ new_n10415;
  assign new_n10420 = ~new_n4212 & n91;
  assign new_n10421 = new_n2481 & new_n4201;
  assign new_n10422 = new_n10421 ^ new_n10420;
  assign new_n10423 = n92 & new_n4200;
  assign new_n10424 = n90 & new_n4206;
  assign new_n10425 = new_n10424 ^ new_n10423;
  assign new_n10426 = new_n10425 ^ new_n10422;
  assign new_n10427 = new_n10426 ^ n42;
  assign new_n10428 = new_n10427 ^ new_n10419;
  assign new_n10429 = new_n10153 ^ new_n10141;
  assign new_n10430 = ~new_n10429 & new_n10150;
  assign new_n10431 = new_n10430 ^ new_n10153;
  assign new_n10432 = new_n10431 ^ new_n10428;
  assign new_n10433 = ~new_n3682 & n94;
  assign new_n10434 = new_n2934 & new_n3677;
  assign new_n10435 = new_n10434 ^ new_n10433;
  assign new_n10436 = n95 & new_n3676;
  assign new_n10437 = n93 & new_n3688;
  assign new_n10438 = new_n10437 ^ new_n10436;
  assign new_n10439 = new_n10438 ^ new_n10435;
  assign new_n10440 = new_n10439 ^ n39;
  assign new_n10441 = new_n10440 ^ new_n10432;
  assign new_n10442 = new_n10166 ^ new_n10154;
  assign new_n10443 = ~new_n10442 & new_n10163;
  assign new_n10444 = new_n10443 ^ new_n10166;
  assign new_n10445 = new_n10444 ^ new_n10441;
  assign new_n10446 = ~new_n3143 & n97;
  assign new_n10447 = new_n3138 & new_n3435;
  assign new_n10448 = new_n10447 ^ new_n10446;
  assign new_n10449 = n98 & new_n3137;
  assign new_n10450 = n96 & new_n3149;
  assign new_n10451 = new_n10450 ^ new_n10449;
  assign new_n10452 = new_n10451 ^ new_n10448;
  assign new_n10453 = new_n10452 ^ n36;
  assign new_n10454 = new_n10453 ^ new_n10445;
  assign new_n10455 = new_n10179 ^ new_n10167;
  assign new_n10456 = ~new_n10455 & new_n10176;
  assign new_n10457 = new_n10456 ^ new_n10179;
  assign new_n10458 = new_n10457 ^ new_n10454;
  assign new_n10459 = ~new_n2672 & n100;
  assign new_n10460 = new_n2667 & new_n3972;
  assign new_n10461 = new_n10460 ^ new_n10459;
  assign new_n10462 = n101 & new_n2666;
  assign new_n10463 = n99 & new_n2664;
  assign new_n10464 = new_n10463 ^ new_n10462;
  assign new_n10465 = new_n10464 ^ new_n10461;
  assign new_n10466 = new_n10465 ^ n33;
  assign new_n10467 = new_n10466 ^ new_n10458;
  assign new_n10468 = new_n10192 ^ new_n10180;
  assign new_n10469 = ~new_n10468 & new_n10189;
  assign new_n10470 = new_n10469 ^ new_n10192;
  assign new_n10471 = new_n10470 ^ new_n10467;
  assign new_n10472 = n103 & new_n2246;
  assign new_n10473 = ~new_n4556 & new_n2241;
  assign new_n10474 = new_n10473 ^ new_n10472;
  assign new_n10475 = n104 & new_n2240;
  assign new_n10476 = n102 & new_n2391;
  assign new_n10477 = new_n10476 ^ new_n10475;
  assign new_n10478 = new_n10477 ^ new_n10474;
  assign new_n10479 = new_n10478 ^ n30;
  assign new_n10480 = new_n10479 ^ new_n10471;
  assign new_n10481 = new_n10205 ^ new_n10193;
  assign new_n10482 = new_n10202 & new_n10481;
  assign new_n10483 = new_n10482 ^ new_n10205;
  assign new_n10484 = new_n10483 ^ new_n10480;
  assign new_n10485 = n106 & new_n1874;
  assign new_n10486 = ~new_n5164 & new_n1864;
  assign new_n10487 = new_n10486 ^ new_n10485;
  assign new_n10488 = n107 & new_n1863;
  assign new_n10489 = n105 & new_n1868;
  assign new_n10490 = new_n10489 ^ new_n10488;
  assign new_n10491 = new_n10490 ^ new_n10487;
  assign new_n10492 = new_n10491 ^ n27;
  assign new_n10493 = new_n10492 ^ new_n10484;
  assign new_n10494 = new_n10218 ^ new_n10206;
  assign new_n10495 = ~new_n10215 & new_n10494;
  assign new_n10496 = new_n10495 ^ new_n10218;
  assign new_n10497 = new_n10496 ^ new_n10493;
  assign new_n10498 = ~new_n1506 & n109;
  assign new_n10499 = new_n1501 & new_n5825;
  assign new_n10500 = new_n10499 ^ new_n10498;
  assign new_n10501 = n110 & new_n1500;
  assign new_n10502 = n108 & new_n1512;
  assign new_n10503 = new_n10502 ^ new_n10501;
  assign new_n10504 = new_n10503 ^ new_n10500;
  assign new_n10505 = new_n10504 ^ n24;
  assign new_n10506 = new_n10505 ^ new_n10497;
  assign new_n10507 = new_n10231 ^ new_n10219;
  assign new_n10508 = ~new_n10228 & new_n10507;
  assign new_n10509 = new_n10508 ^ new_n10231;
  assign new_n10510 = new_n10509 ^ new_n10506;
  assign new_n10511 = ~new_n1198 & n112;
  assign new_n10512 = ~new_n6518 & new_n1193;
  assign new_n10513 = new_n10512 ^ new_n10511;
  assign new_n10514 = n113 & new_n1192;
  assign new_n10515 = n111 & new_n1204;
  assign new_n10516 = new_n10515 ^ new_n10514;
  assign new_n10517 = new_n10516 ^ new_n10513;
  assign new_n10518 = new_n10517 ^ n21;
  assign new_n10519 = new_n10518 ^ new_n10510;
  assign new_n10520 = new_n10244 ^ new_n10232;
  assign new_n10521 = ~new_n10241 & new_n10520;
  assign new_n10522 = new_n10521 ^ new_n10244;
  assign new_n10523 = new_n10522 ^ new_n10519;
  assign new_n10524 = ~new_n930 & n115;
  assign new_n10525 = ~new_n7256 & new_n925;
  assign new_n10526 = new_n10525 ^ new_n10524;
  assign new_n10527 = n116 & new_n924;
  assign new_n10528 = n114 & new_n936;
  assign new_n10529 = new_n10528 ^ new_n10527;
  assign new_n10530 = new_n10529 ^ new_n10526;
  assign new_n10531 = new_n10530 ^ n18;
  assign new_n10532 = new_n10531 ^ new_n10523;
  assign new_n10533 = new_n10257 ^ new_n10245;
  assign new_n10534 = ~new_n10254 & new_n10533;
  assign new_n10535 = new_n10534 ^ new_n10257;
  assign new_n10536 = new_n10535 ^ new_n10532;
  assign new_n10537 = n118 & new_n707;
  assign new_n10538 = ~new_n8019 & new_n701;
  assign new_n10539 = new_n10538 ^ new_n10537;
  assign new_n10540 = n119 & new_n700;
  assign new_n10541 = n117 & new_n787;
  assign new_n10542 = new_n10541 ^ new_n10540;
  assign new_n10543 = new_n10542 ^ new_n10539;
  assign new_n10544 = new_n10543 ^ n15;
  assign new_n10545 = new_n10544 ^ new_n10536;
  assign new_n10546 = new_n10270 ^ new_n10258;
  assign new_n10547 = ~new_n10267 & new_n10546;
  assign new_n10548 = new_n10547 ^ new_n10270;
  assign new_n10549 = new_n10548 ^ new_n10545;
  assign new_n10550 = n121 & new_n499;
  assign new_n10551 = ~new_n506 & new_n8850;
  assign new_n10552 = new_n10551 ^ new_n10550;
  assign new_n10553 = ~new_n505 & n122;
  assign new_n10554 = n120 & new_n579;
  assign new_n10555 = new_n10554 ^ new_n10553;
  assign new_n10556 = new_n10555 ^ new_n10552;
  assign new_n10557 = new_n10556 ^ n12;
  assign new_n10558 = new_n10557 ^ new_n10549;
  assign new_n10559 = new_n10283 ^ new_n10271;
  assign new_n10560 = ~new_n10280 & new_n10559;
  assign new_n10561 = new_n10560 ^ new_n10283;
  assign new_n10562 = new_n10561 ^ new_n10558;
  assign new_n10563 = new_n10292 ^ new_n10284;
  assign new_n10564 = ~new_n10301 & new_n10563;
  assign new_n10565 = new_n10564 ^ new_n10284;
  assign new_n10566 = new_n10565 ^ new_n10562;
  assign new_n10567 = n124 & new_n354;
  assign new_n10568 = new_n349 & new_n9700;
  assign new_n10569 = new_n10568 ^ new_n10567;
  assign new_n10570 = n125 & new_n348;
  assign new_n10571 = n123 & new_n391;
  assign new_n10572 = new_n10571 ^ new_n10570;
  assign new_n10573 = new_n10572 ^ new_n10569;
  assign new_n10574 = new_n10573 ^ n9;
  assign new_n10575 = new_n10574 ^ new_n10566;
  assign new_n10576 = new_n10315 ^ new_n10302;
  assign new_n10577 = ~new_n10312 & new_n10576;
  assign new_n10578 = new_n10577 ^ new_n10315;
  assign new_n10579 = new_n10578 ^ new_n10575;
  assign new_n10580 = n127 & new_n218;
  assign new_n10581 = new_n9723 ^ n128;
  assign new_n10582 = new_n208 & new_n10581;
  assign new_n10583 = new_n10582 ^ new_n10580;
  assign new_n10584 = n128 & new_n207;
  assign new_n10585 = n126 & new_n212;
  assign new_n10586 = new_n10585 ^ new_n10584;
  assign new_n10587 = new_n10586 ^ new_n10583;
  assign new_n10588 = new_n10587 ^ n6;
  assign new_n10589 = new_n10588 ^ new_n10579;
  assign new_n10590 = new_n10316 ^ new_n10058;
  assign new_n10591 = ~new_n10590 & new_n10059;
  assign new_n10592 = new_n10591 ^ new_n10042;
  assign new_n10593 = new_n10592 ^ new_n10589;
  assign new_n10594 = new_n10324 ^ new_n10317;
  assign new_n10595 = ~new_n10321 & ~new_n10594;
  assign new_n10596 = new_n10595 ^ new_n10324;
  assign new_n10597 = new_n10596 ^ new_n10593;
  assign new_n10598 = ~new_n6110 & n83;
  assign new_n10599 = new_n1468 & new_n6105;
  assign new_n10600 = new_n10599 ^ new_n10598;
  assign new_n10601 = n84 & new_n6104;
  assign new_n10602 = n82 & new_n6347;
  assign new_n10603 = new_n10602 ^ new_n10601;
  assign new_n10604 = new_n10603 ^ new_n10600;
  assign new_n10605 = new_n10604 ^ n51;
  assign new_n10606 = new_n10379 ^ new_n10367;
  assign new_n10607 = ~new_n10606 & new_n10376;
  assign new_n10608 = new_n10607 ^ new_n10379;
  assign new_n10609 = new_n10608 ^ new_n10605;
  assign new_n10610 = ~new_n6805 & n80;
  assign new_n10611 = new_n1161 & new_n6800;
  assign new_n10612 = new_n10611 ^ new_n10610;
  assign new_n10613 = n79 & new_n6811;
  assign new_n10614 = n81 & new_n6799;
  assign new_n10615 = new_n10614 ^ new_n10613;
  assign new_n10616 = new_n10615 ^ new_n10612;
  assign new_n10617 = new_n10616 ^ n54;
  assign new_n10618 = n77 & new_n7553;
  assign new_n10619 = ~new_n891 & new_n7543;
  assign new_n10620 = new_n10619 ^ new_n10618;
  assign new_n10621 = n78 & new_n7542;
  assign new_n10622 = n76 & new_n7547;
  assign new_n10623 = new_n10622 ^ new_n10621;
  assign new_n10624 = new_n10623 ^ new_n10620;
  assign new_n10625 = new_n10624 ^ n57;
  assign new_n10626 = n71 & new_n9195;
  assign new_n10627 = ~new_n459 & new_n9185;
  assign new_n10628 = new_n10627 ^ new_n10626;
  assign new_n10629 = n72 & new_n9184;
  assign new_n10630 = n70 & new_n9189;
  assign new_n10631 = new_n10630 ^ new_n10629;
  assign new_n10632 = new_n10631 ^ new_n10628;
  assign new_n10633 = n64 & n69;
  assign new_n10634 = new_n10633 ^ n69;
  assign new_n10635 = new_n10634 ^ new_n10341;
  assign new_n10636 = new_n10635 ^ new_n10633;
  assign new_n10637 = ~n63 & ~new_n10636;
  assign new_n10638 = new_n10637 ^ new_n10635;
  assign new_n10639 = new_n10638 ^ n3;
  assign new_n10640 = new_n10639 ^ new_n10632;
  assign new_n10641 = new_n10340 ^ n3;
  assign new_n10642 = new_n10344 ^ n3;
  assign new_n10643 = ~new_n10641 & new_n10642;
  assign new_n10644 = new_n10643 ^ n3;
  assign new_n10645 = new_n10341 ^ n3;
  assign new_n10646 = new_n10641 & new_n10645;
  assign new_n10647 = new_n10646 ^ n3;
  assign new_n10648 = new_n10647 ^ new_n10644;
  assign new_n10649 = ~n63 & new_n10648;
  assign new_n10650 = new_n10649 ^ new_n10644;
  assign new_n10651 = new_n10650 ^ new_n10640;
  assign new_n10652 = n74 & new_n8355;
  assign new_n10653 = new_n660 & new_n8345;
  assign new_n10654 = new_n10653 ^ new_n10652;
  assign new_n10655 = n75 & new_n8344;
  assign new_n10656 = n73 & new_n8349;
  assign new_n10657 = new_n10656 ^ new_n10655;
  assign new_n10658 = new_n10657 ^ new_n10654;
  assign new_n10659 = new_n10658 ^ n60;
  assign new_n10660 = new_n10659 ^ new_n10651;
  assign new_n10661 = new_n10660 ^ new_n10625;
  assign new_n10662 = new_n10353 ^ new_n10333;
  assign new_n10663 = ~new_n10662 & new_n10350;
  assign new_n10664 = new_n10663 ^ new_n10353;
  assign new_n10665 = new_n10664 ^ new_n10661;
  assign new_n10666 = new_n10665 ^ new_n10617;
  assign new_n10667 = new_n10366 ^ new_n10354;
  assign new_n10668 = ~new_n10363 & ~new_n10667;
  assign new_n10669 = new_n10668 ^ new_n10366;
  assign new_n10670 = new_n10669 ^ new_n10666;
  assign new_n10671 = new_n10670 ^ new_n10609;
  assign new_n10672 = ~new_n5424 & n86;
  assign new_n10673 = new_n1811 & new_n5419;
  assign new_n10674 = new_n10673 ^ new_n10672;
  assign new_n10675 = n87 & new_n5418;
  assign new_n10676 = n85 & new_n5648;
  assign new_n10677 = new_n10676 ^ new_n10675;
  assign new_n10678 = new_n10677 ^ new_n10674;
  assign new_n10679 = new_n10678 ^ n48;
  assign new_n10680 = new_n10679 ^ new_n10671;
  assign new_n10681 = new_n10392 ^ new_n10380;
  assign new_n10682 = ~new_n10681 & new_n10389;
  assign new_n10683 = new_n10682 ^ new_n10392;
  assign new_n10684 = new_n10683 ^ new_n10680;
  assign new_n10685 = ~new_n4804 & n89;
  assign new_n10686 = new_n2193 & new_n4799;
  assign new_n10687 = new_n10686 ^ new_n10685;
  assign new_n10688 = n90 & new_n4798;
  assign new_n10689 = n88 & new_n4810;
  assign new_n10690 = new_n10689 ^ new_n10688;
  assign new_n10691 = new_n10690 ^ new_n10687;
  assign new_n10692 = new_n10691 ^ n45;
  assign new_n10693 = new_n10692 ^ new_n10684;
  assign new_n10694 = new_n10405 ^ new_n10393;
  assign new_n10695 = ~new_n10694 & new_n10402;
  assign new_n10696 = new_n10695 ^ new_n10405;
  assign new_n10697 = new_n10696 ^ new_n10693;
  assign new_n10698 = ~new_n4212 & n92;
  assign new_n10699 = new_n2628 & new_n4201;
  assign new_n10700 = new_n10699 ^ new_n10698;
  assign new_n10701 = n93 & new_n4200;
  assign new_n10702 = n91 & new_n4206;
  assign new_n10703 = new_n10702 ^ new_n10701;
  assign new_n10704 = new_n10703 ^ new_n10700;
  assign new_n10705 = new_n10704 ^ n42;
  assign new_n10706 = new_n10705 ^ new_n10697;
  assign new_n10707 = new_n10418 ^ new_n10406;
  assign new_n10708 = new_n10415 & new_n10707;
  assign new_n10709 = new_n10708 ^ new_n10418;
  assign new_n10710 = new_n10709 ^ new_n10706;
  assign new_n10711 = ~new_n3682 & n95;
  assign new_n10712 = new_n3095 & new_n3677;
  assign new_n10713 = new_n10712 ^ new_n10711;
  assign new_n10714 = n96 & new_n3676;
  assign new_n10715 = n94 & new_n3688;
  assign new_n10716 = new_n10715 ^ new_n10714;
  assign new_n10717 = new_n10716 ^ new_n10713;
  assign new_n10718 = new_n10717 ^ n39;
  assign new_n10719 = new_n10718 ^ new_n10710;
  assign new_n10720 = new_n10431 ^ new_n10419;
  assign new_n10721 = ~new_n10428 & new_n10720;
  assign new_n10722 = new_n10721 ^ new_n10431;
  assign new_n10723 = new_n10722 ^ new_n10719;
  assign new_n10724 = ~new_n3143 & n98;
  assign new_n10725 = new_n3138 & new_n3604;
  assign new_n10726 = new_n10725 ^ new_n10724;
  assign new_n10727 = n99 & new_n3137;
  assign new_n10728 = n97 & new_n3149;
  assign new_n10729 = new_n10728 ^ new_n10727;
  assign new_n10730 = new_n10729 ^ new_n10726;
  assign new_n10731 = new_n10730 ^ n36;
  assign new_n10732 = new_n10731 ^ new_n10723;
  assign new_n10733 = new_n10444 ^ new_n10432;
  assign new_n10734 = ~new_n10441 & new_n10733;
  assign new_n10735 = new_n10734 ^ new_n10444;
  assign new_n10736 = new_n10735 ^ new_n10732;
  assign new_n10737 = ~new_n2672 & n101;
  assign new_n10738 = new_n2667 & new_n4159;
  assign new_n10739 = new_n10738 ^ new_n10737;
  assign new_n10740 = n102 & new_n2666;
  assign new_n10741 = n100 & new_n2664;
  assign new_n10742 = new_n10741 ^ new_n10740;
  assign new_n10743 = new_n10742 ^ new_n10739;
  assign new_n10744 = new_n10743 ^ n33;
  assign new_n10745 = new_n10744 ^ new_n10736;
  assign new_n10746 = new_n10457 ^ new_n10445;
  assign new_n10747 = ~new_n10454 & new_n10746;
  assign new_n10748 = new_n10747 ^ new_n10457;
  assign new_n10749 = new_n10748 ^ new_n10745;
  assign new_n10750 = n104 & new_n2246;
  assign new_n10751 = ~new_n4754 & new_n2241;
  assign new_n10752 = new_n10751 ^ new_n10750;
  assign new_n10753 = n105 & new_n2240;
  assign new_n10754 = n103 & new_n2391;
  assign new_n10755 = new_n10754 ^ new_n10753;
  assign new_n10756 = new_n10755 ^ new_n10752;
  assign new_n10757 = new_n10756 ^ n30;
  assign new_n10758 = new_n10757 ^ new_n10749;
  assign new_n10759 = new_n10470 ^ new_n10458;
  assign new_n10760 = ~new_n10467 & new_n10759;
  assign new_n10761 = new_n10760 ^ new_n10470;
  assign new_n10762 = new_n10761 ^ new_n10758;
  assign new_n10763 = n107 & new_n1874;
  assign new_n10764 = ~new_n5377 & new_n1864;
  assign new_n10765 = new_n10764 ^ new_n10763;
  assign new_n10766 = n108 & new_n1863;
  assign new_n10767 = n106 & new_n1868;
  assign new_n10768 = new_n10767 ^ new_n10766;
  assign new_n10769 = new_n10768 ^ new_n10765;
  assign new_n10770 = new_n10769 ^ n27;
  assign new_n10771 = new_n10770 ^ new_n10762;
  assign new_n10772 = new_n10483 ^ new_n10471;
  assign new_n10773 = ~new_n10480 & ~new_n10772;
  assign new_n10774 = new_n10773 ^ new_n10483;
  assign new_n10775 = new_n10774 ^ new_n10771;
  assign new_n10776 = ~new_n1506 & n110;
  assign new_n10777 = new_n1501 & new_n6049;
  assign new_n10778 = new_n10777 ^ new_n10776;
  assign new_n10779 = n111 & new_n1500;
  assign new_n10780 = n109 & new_n1512;
  assign new_n10781 = new_n10780 ^ new_n10779;
  assign new_n10782 = new_n10781 ^ new_n10778;
  assign new_n10783 = new_n10782 ^ n24;
  assign new_n10784 = new_n10783 ^ new_n10775;
  assign new_n10785 = new_n10496 ^ new_n10484;
  assign new_n10786 = ~new_n10785 & new_n10493;
  assign new_n10787 = new_n10786 ^ new_n10496;
  assign new_n10788 = new_n10787 ^ new_n10784;
  assign new_n10789 = ~new_n1198 & n113;
  assign new_n10790 = ~new_n6764 & new_n1193;
  assign new_n10791 = new_n10790 ^ new_n10789;
  assign new_n10792 = n114 & new_n1192;
  assign new_n10793 = n112 & new_n1204;
  assign new_n10794 = new_n10793 ^ new_n10792;
  assign new_n10795 = new_n10794 ^ new_n10791;
  assign new_n10796 = new_n10795 ^ n21;
  assign new_n10797 = new_n10796 ^ new_n10788;
  assign new_n10798 = new_n10509 ^ new_n10497;
  assign new_n10799 = ~new_n10798 & new_n10506;
  assign new_n10800 = new_n10799 ^ new_n10509;
  assign new_n10801 = new_n10800 ^ new_n10797;
  assign new_n10802 = ~new_n930 & n116;
  assign new_n10803 = ~new_n7503 & new_n925;
  assign new_n10804 = new_n10803 ^ new_n10802;
  assign new_n10805 = n117 & new_n924;
  assign new_n10806 = n115 & new_n936;
  assign new_n10807 = new_n10806 ^ new_n10805;
  assign new_n10808 = new_n10807 ^ new_n10804;
  assign new_n10809 = new_n10808 ^ n18;
  assign new_n10810 = new_n10809 ^ new_n10801;
  assign new_n10811 = new_n10522 ^ new_n10510;
  assign new_n10812 = ~new_n10811 & new_n10519;
  assign new_n10813 = new_n10812 ^ new_n10522;
  assign new_n10814 = new_n10813 ^ new_n10810;
  assign new_n10815 = n119 & new_n707;
  assign new_n10816 = new_n701 & new_n8286;
  assign new_n10817 = new_n10816 ^ new_n10815;
  assign new_n10818 = n120 & new_n700;
  assign new_n10819 = n118 & new_n787;
  assign new_n10820 = new_n10819 ^ new_n10818;
  assign new_n10821 = new_n10820 ^ new_n10817;
  assign new_n10822 = new_n10821 ^ n15;
  assign new_n10823 = new_n10822 ^ new_n10814;
  assign new_n10824 = new_n10535 ^ new_n10523;
  assign new_n10825 = ~new_n10824 & new_n10532;
  assign new_n10826 = new_n10825 ^ new_n10535;
  assign new_n10827 = new_n10826 ^ new_n10823;
  assign new_n10828 = n122 & new_n499;
  assign new_n10829 = ~new_n506 & ~new_n9116;
  assign new_n10830 = new_n10829 ^ new_n10828;
  assign new_n10831 = ~new_n505 & n123;
  assign new_n10832 = n121 & new_n579;
  assign new_n10833 = new_n10832 ^ new_n10831;
  assign new_n10834 = new_n10833 ^ new_n10830;
  assign new_n10835 = new_n10834 ^ n12;
  assign new_n10836 = new_n10835 ^ new_n10827;
  assign new_n10837 = new_n10548 ^ new_n10536;
  assign new_n10838 = ~new_n10837 & new_n10545;
  assign new_n10839 = new_n10838 ^ new_n10548;
  assign new_n10840 = new_n10839 ^ new_n10836;
  assign new_n10841 = n125 & new_n354;
  assign new_n10842 = new_n349 & new_n9987;
  assign new_n10843 = new_n10842 ^ new_n10841;
  assign new_n10844 = n126 & new_n348;
  assign new_n10845 = n124 & new_n391;
  assign new_n10846 = new_n10845 ^ new_n10844;
  assign new_n10847 = new_n10846 ^ new_n10843;
  assign new_n10848 = new_n10847 ^ n9;
  assign new_n10849 = new_n10848 ^ new_n10840;
  assign new_n10850 = new_n10561 ^ new_n10549;
  assign new_n10851 = ~new_n10850 & new_n10558;
  assign new_n10852 = new_n10851 ^ new_n10561;
  assign new_n10853 = new_n10852 ^ new_n10849;
  assign new_n10854 = n127 & new_n212;
  assign new_n10855 = new_n208 & new_n10010;
  assign new_n10856 = new_n10855 ^ new_n10854;
  assign new_n10857 = n128 & new_n218;
  assign new_n10858 = new_n10857 ^ new_n10856;
  assign new_n10859 = new_n10858 ^ n6;
  assign new_n10860 = new_n10859 ^ new_n10853;
  assign new_n10861 = new_n10574 ^ new_n10562;
  assign new_n10862 = ~new_n10566 & new_n10861;
  assign new_n10863 = new_n10862 ^ new_n10565;
  assign new_n10864 = new_n10863 ^ new_n10860;
  assign new_n10865 = new_n10588 ^ new_n10575;
  assign new_n10866 = ~new_n10579 & new_n10865;
  assign new_n10867 = new_n10866 ^ new_n10578;
  assign new_n10868 = new_n10867 ^ new_n10864;
  assign new_n10869 = new_n10596 ^ new_n10589;
  assign new_n10870 = new_n10593 & new_n10869;
  assign new_n10871 = new_n10870 ^ new_n10596;
  assign new_n10872 = new_n10871 ^ new_n10868;
  assign new_n10873 = ~new_n6110 & n84;
  assign new_n10874 = new_n1584 & new_n6105;
  assign new_n10875 = new_n10874 ^ new_n10873;
  assign new_n10876 = n85 & new_n6104;
  assign new_n10877 = n83 & new_n6347;
  assign new_n10878 = new_n10877 ^ new_n10876;
  assign new_n10879 = new_n10878 ^ new_n10875;
  assign new_n10880 = new_n10879 ^ n51;
  assign new_n10881 = ~new_n6805 & n81;
  assign new_n10882 = new_n1263 & new_n6800;
  assign new_n10883 = new_n10882 ^ new_n10881;
  assign new_n10884 = n82 & new_n6799;
  assign new_n10885 = n80 & new_n6811;
  assign new_n10886 = new_n10885 ^ new_n10884;
  assign new_n10887 = new_n10886 ^ new_n10883;
  assign new_n10888 = new_n10887 ^ n54;
  assign new_n10889 = n78 & new_n7553;
  assign new_n10890 = ~new_n982 & new_n7543;
  assign new_n10891 = new_n10890 ^ new_n10889;
  assign new_n10892 = n79 & new_n7542;
  assign new_n10893 = n77 & new_n7547;
  assign new_n10894 = new_n10893 ^ new_n10892;
  assign new_n10895 = new_n10894 ^ new_n10891;
  assign new_n10896 = new_n10895 ^ n57;
  assign new_n10897 = new_n10659 ^ new_n10640;
  assign new_n10898 = ~new_n10651 & new_n10897;
  assign new_n10899 = new_n10898 ^ new_n10650;
  assign new_n10900 = new_n10899 ^ new_n10896;
  assign new_n10901 = n75 & new_n8355;
  assign new_n10902 = ~new_n737 & new_n8345;
  assign new_n10903 = new_n10902 ^ new_n10901;
  assign new_n10904 = n76 & new_n8344;
  assign new_n10905 = n74 & new_n8349;
  assign new_n10906 = new_n10905 ^ new_n10904;
  assign new_n10907 = new_n10906 ^ new_n10903;
  assign new_n10908 = new_n10907 ^ n60;
  assign new_n10909 = new_n10632 ^ n3;
  assign new_n10910 = new_n10635 ^ n3;
  assign new_n10911 = ~new_n10909 & new_n10910;
  assign new_n10912 = new_n10911 ^ n3;
  assign new_n10913 = new_n10633 ^ n3;
  assign new_n10914 = new_n10909 & new_n10913;
  assign new_n10915 = new_n10914 ^ n3;
  assign new_n10916 = new_n10915 ^ new_n10912;
  assign new_n10917 = ~n63 & new_n10916;
  assign new_n10918 = new_n10917 ^ new_n10912;
  assign new_n10919 = new_n10918 ^ new_n10908;
  assign new_n10920 = n72 & new_n9195;
  assign new_n10921 = new_n534 & new_n9185;
  assign new_n10922 = new_n10921 ^ new_n10920;
  assign new_n10923 = n73 & new_n9184;
  assign new_n10924 = n71 & new_n9189;
  assign new_n10925 = new_n10924 ^ new_n10923;
  assign new_n10926 = new_n10925 ^ new_n10922;
  assign new_n10927 = n64 & n70;
  assign new_n10928 = new_n10927 ^ n70;
  assign new_n10929 = new_n10928 ^ new_n10634;
  assign new_n10930 = new_n10929 ^ n69;
  assign new_n10931 = new_n10930 ^ new_n10927;
  assign new_n10932 = ~n63 & ~new_n10931;
  assign new_n10933 = new_n10932 ^ new_n10930;
  assign new_n10934 = new_n10933 ^ n3;
  assign new_n10935 = new_n10934 ^ new_n10926;
  assign new_n10936 = new_n10935 ^ new_n10919;
  assign new_n10937 = new_n10936 ^ new_n10900;
  assign new_n10938 = new_n10937 ^ new_n10888;
  assign new_n10939 = new_n10664 ^ new_n10660;
  assign new_n10940 = ~new_n10661 & ~new_n10939;
  assign new_n10941 = new_n10940 ^ new_n10625;
  assign new_n10942 = new_n10941 ^ new_n10938;
  assign new_n10943 = new_n10942 ^ new_n10880;
  assign new_n10944 = new_n10669 ^ new_n10617;
  assign new_n10945 = ~new_n10666 & ~new_n10944;
  assign new_n10946 = new_n10945 ^ new_n10669;
  assign new_n10947 = new_n10946 ^ new_n10943;
  assign new_n10948 = new_n10670 ^ new_n10605;
  assign new_n10949 = new_n10609 & new_n10948;
  assign new_n10950 = new_n10949 ^ new_n10608;
  assign new_n10951 = new_n10950 ^ new_n10947;
  assign new_n10952 = ~new_n5424 & n87;
  assign new_n10953 = new_n1940 & new_n5419;
  assign new_n10954 = new_n10953 ^ new_n10952;
  assign new_n10955 = n88 & new_n5418;
  assign new_n10956 = n86 & new_n5648;
  assign new_n10957 = new_n10956 ^ new_n10955;
  assign new_n10958 = new_n10957 ^ new_n10954;
  assign new_n10959 = new_n10958 ^ n48;
  assign new_n10960 = new_n10959 ^ new_n10951;
  assign new_n10961 = ~new_n4804 & n90;
  assign new_n10962 = new_n2341 & new_n4799;
  assign new_n10963 = new_n10962 ^ new_n10961;
  assign new_n10964 = n91 & new_n4798;
  assign new_n10965 = n89 & new_n4810;
  assign new_n10966 = new_n10965 ^ new_n10964;
  assign new_n10967 = new_n10966 ^ new_n10963;
  assign new_n10968 = new_n10967 ^ n45;
  assign new_n10969 = new_n10968 ^ new_n10960;
  assign new_n10970 = new_n10683 ^ new_n10671;
  assign new_n10971 = ~new_n10970 & new_n10680;
  assign new_n10972 = new_n10971 ^ new_n10683;
  assign new_n10973 = new_n10972 ^ new_n10969;
  assign new_n10974 = ~new_n4212 & n93;
  assign new_n10975 = new_n2785 & new_n4201;
  assign new_n10976 = new_n10975 ^ new_n10974;
  assign new_n10977 = n94 & new_n4200;
  assign new_n10978 = n92 & new_n4206;
  assign new_n10979 = new_n10978 ^ new_n10977;
  assign new_n10980 = new_n10979 ^ new_n10976;
  assign new_n10981 = new_n10980 ^ n42;
  assign new_n10982 = new_n10981 ^ new_n10973;
  assign new_n10983 = new_n10696 ^ new_n10684;
  assign new_n10984 = ~new_n10983 & new_n10693;
  assign new_n10985 = new_n10984 ^ new_n10696;
  assign new_n10986 = new_n10985 ^ new_n10982;
  assign new_n10987 = ~new_n3682 & n96;
  assign new_n10988 = new_n3273 & new_n3677;
  assign new_n10989 = new_n10988 ^ new_n10987;
  assign new_n10990 = n97 & new_n3676;
  assign new_n10991 = n95 & new_n3688;
  assign new_n10992 = new_n10991 ^ new_n10990;
  assign new_n10993 = new_n10992 ^ new_n10989;
  assign new_n10994 = new_n10993 ^ n39;
  assign new_n10995 = new_n10994 ^ new_n10986;
  assign new_n10996 = new_n10709 ^ new_n10697;
  assign new_n10997 = new_n10706 & new_n10996;
  assign new_n10998 = new_n10997 ^ new_n10709;
  assign new_n10999 = new_n10998 ^ new_n10995;
  assign new_n11000 = ~new_n3143 & n99;
  assign new_n11001 = new_n3138 & new_n3789;
  assign new_n11002 = new_n11001 ^ new_n11000;
  assign new_n11003 = n100 & new_n3137;
  assign new_n11004 = n98 & new_n3149;
  assign new_n11005 = new_n11004 ^ new_n11003;
  assign new_n11006 = new_n11005 ^ new_n11002;
  assign new_n11007 = new_n11006 ^ n36;
  assign new_n11008 = new_n11007 ^ new_n10999;
  assign new_n11009 = new_n10722 ^ new_n10710;
  assign new_n11010 = ~new_n10719 & new_n11009;
  assign new_n11011 = new_n11010 ^ new_n10722;
  assign new_n11012 = new_n11011 ^ new_n11008;
  assign new_n11013 = ~new_n2672 & n102;
  assign new_n11014 = new_n2667 & new_n4368;
  assign new_n11015 = new_n11014 ^ new_n11013;
  assign new_n11016 = n103 & new_n2666;
  assign new_n11017 = n101 & new_n2664;
  assign new_n11018 = new_n11017 ^ new_n11016;
  assign new_n11019 = new_n11018 ^ new_n11015;
  assign new_n11020 = new_n11019 ^ n33;
  assign new_n11021 = new_n11020 ^ new_n11012;
  assign new_n11022 = new_n10735 ^ new_n10723;
  assign new_n11023 = ~new_n10732 & new_n11022;
  assign new_n11024 = new_n11023 ^ new_n10735;
  assign new_n11025 = new_n11024 ^ new_n11021;
  assign new_n11026 = n105 & new_n2246;
  assign new_n11027 = ~new_n4961 & new_n2241;
  assign new_n11028 = new_n11027 ^ new_n11026;
  assign new_n11029 = n106 & new_n2240;
  assign new_n11030 = n104 & new_n2391;
  assign new_n11031 = new_n11030 ^ new_n11029;
  assign new_n11032 = new_n11031 ^ new_n11028;
  assign new_n11033 = new_n11032 ^ n30;
  assign new_n11034 = new_n11033 ^ new_n11025;
  assign new_n11035 = new_n10748 ^ new_n10736;
  assign new_n11036 = ~new_n10745 & new_n11035;
  assign new_n11037 = new_n11036 ^ new_n10748;
  assign new_n11038 = new_n11037 ^ new_n11034;
  assign new_n11039 = n108 & new_n1874;
  assign new_n11040 = new_n1864 & new_n5604;
  assign new_n11041 = new_n11040 ^ new_n11039;
  assign new_n11042 = n109 & new_n1863;
  assign new_n11043 = n107 & new_n1868;
  assign new_n11044 = new_n11043 ^ new_n11042;
  assign new_n11045 = new_n11044 ^ new_n11041;
  assign new_n11046 = new_n11045 ^ n27;
  assign new_n11047 = new_n11046 ^ new_n11038;
  assign new_n11048 = new_n10761 ^ new_n10749;
  assign new_n11049 = ~new_n10758 & new_n11048;
  assign new_n11050 = new_n11049 ^ new_n10761;
  assign new_n11051 = new_n11050 ^ new_n11047;
  assign new_n11052 = ~new_n1506 & n111;
  assign new_n11053 = ~new_n6284 & new_n1501;
  assign new_n11054 = new_n11053 ^ new_n11052;
  assign new_n11055 = n112 & new_n1500;
  assign new_n11056 = n110 & new_n1512;
  assign new_n11057 = new_n11056 ^ new_n11055;
  assign new_n11058 = new_n11057 ^ new_n11054;
  assign new_n11059 = new_n11058 ^ n24;
  assign new_n11060 = new_n11059 ^ new_n11051;
  assign new_n11061 = new_n10774 ^ new_n10762;
  assign new_n11062 = ~new_n10771 & ~new_n11061;
  assign new_n11063 = new_n11062 ^ new_n10774;
  assign new_n11064 = new_n11063 ^ new_n11060;
  assign new_n11065 = ~new_n1198 & n114;
  assign new_n11066 = ~new_n7013 & new_n1193;
  assign new_n11067 = new_n11066 ^ new_n11065;
  assign new_n11068 = n115 & new_n1192;
  assign new_n11069 = n113 & new_n1204;
  assign new_n11070 = new_n11069 ^ new_n11068;
  assign new_n11071 = new_n11070 ^ new_n11067;
  assign new_n11072 = new_n11071 ^ n21;
  assign new_n11073 = new_n11072 ^ new_n11064;
  assign new_n11074 = new_n10787 ^ new_n10775;
  assign new_n11075 = ~new_n11074 & new_n10784;
  assign new_n11076 = new_n11075 ^ new_n10787;
  assign new_n11077 = new_n11076 ^ new_n11073;
  assign new_n11078 = ~new_n930 & n117;
  assign new_n11079 = ~new_n7761 & new_n925;
  assign new_n11080 = new_n11079 ^ new_n11078;
  assign new_n11081 = n118 & new_n924;
  assign new_n11082 = n116 & new_n936;
  assign new_n11083 = new_n11082 ^ new_n11081;
  assign new_n11084 = new_n11083 ^ new_n11080;
  assign new_n11085 = new_n11084 ^ n18;
  assign new_n11086 = new_n11085 ^ new_n11077;
  assign new_n11087 = new_n10800 ^ new_n10788;
  assign new_n11088 = ~new_n11087 & new_n10797;
  assign new_n11089 = new_n11088 ^ new_n10800;
  assign new_n11090 = new_n11089 ^ new_n11086;
  assign new_n11091 = n120 & new_n707;
  assign new_n11092 = new_n701 & new_n8560;
  assign new_n11093 = new_n11092 ^ new_n11091;
  assign new_n11094 = n121 & new_n700;
  assign new_n11095 = n119 & new_n787;
  assign new_n11096 = new_n11095 ^ new_n11094;
  assign new_n11097 = new_n11096 ^ new_n11093;
  assign new_n11098 = new_n11097 ^ n15;
  assign new_n11099 = new_n11098 ^ new_n11090;
  assign new_n11100 = new_n10813 ^ new_n10801;
  assign new_n11101 = ~new_n11100 & new_n10810;
  assign new_n11102 = new_n11101 ^ new_n10813;
  assign new_n11103 = new_n11102 ^ new_n11099;
  assign new_n11104 = n123 & new_n499;
  assign new_n11105 = ~new_n506 & ~new_n9405;
  assign new_n11106 = new_n11105 ^ new_n11104;
  assign new_n11107 = ~new_n505 & n124;
  assign new_n11108 = n122 & new_n579;
  assign new_n11109 = new_n11108 ^ new_n11107;
  assign new_n11110 = new_n11109 ^ new_n11106;
  assign new_n11111 = new_n11110 ^ n12;
  assign new_n11112 = new_n11111 ^ new_n11103;
  assign new_n11113 = new_n10826 ^ new_n10814;
  assign new_n11114 = ~new_n11113 & new_n10823;
  assign new_n11115 = new_n11114 ^ new_n10826;
  assign new_n11116 = new_n11115 ^ new_n11112;
  assign new_n11117 = n126 & new_n354;
  assign new_n11118 = new_n349 & new_n10304;
  assign new_n11119 = new_n11118 ^ new_n11117;
  assign new_n11120 = n127 & new_n348;
  assign new_n11121 = n125 & new_n391;
  assign new_n11122 = new_n11121 ^ new_n11120;
  assign new_n11123 = new_n11122 ^ new_n11119;
  assign new_n11124 = new_n11123 ^ n9;
  assign new_n11125 = new_n11124 ^ new_n11116;
  assign new_n11126 = new_n10839 ^ new_n10827;
  assign new_n11127 = ~new_n11126 & new_n10836;
  assign new_n11128 = new_n11127 ^ new_n10839;
  assign new_n11129 = new_n11128 ^ new_n11125;
  assign new_n11130 = n128 & new_n211;
  assign new_n11131 = ~n6 & ~new_n11130;
  assign new_n11132 = new_n11131 ^ n5;
  assign new_n11133 = new_n10009 ^ n128;
  assign new_n11134 = new_n197 & new_n11133;
  assign new_n11135 = new_n11134 ^ new_n11130;
  assign new_n11136 = ~new_n11132 & ~new_n11135;
  assign new_n11137 = new_n11136 ^ n5;
  assign new_n11138 = new_n11137 ^ new_n11129;
  assign new_n11139 = new_n10852 ^ new_n10840;
  assign new_n11140 = ~new_n11139 & new_n10849;
  assign new_n11141 = new_n11140 ^ new_n10852;
  assign new_n11142 = new_n11141 ^ new_n11138;
  assign new_n11143 = new_n10863 ^ new_n10853;
  assign new_n11144 = ~new_n11143 & new_n10860;
  assign new_n11145 = new_n11144 ^ new_n10863;
  assign new_n11146 = new_n11145 ^ new_n11142;
  assign new_n11147 = new_n10871 ^ new_n10867;
  assign new_n11148 = ~new_n11147 & new_n10868;
  assign new_n11149 = new_n11148 ^ new_n10871;
  assign new_n11150 = new_n11149 ^ new_n11146;
  assign new_n11151 = new_n11129 & new_n11145;
  assign new_n11152 = new_n11145 ^ new_n11129;
  assign new_n11153 = new_n11152 ^ new_n11151;
  assign new_n11154 = new_n11153 ^ new_n11149;
  assign new_n11155 = ~new_n11149 & new_n11153;
  assign new_n11156 = new_n11155 ^ new_n11154;
  assign new_n11157 = new_n11142 & new_n11156;
  assign new_n11158 = new_n11141 ^ new_n11137;
  assign new_n11159 = new_n11137 & new_n11141;
  assign new_n11160 = new_n11159 ^ new_n11158;
  assign new_n11161 = new_n11153 & new_n11159;
  assign new_n11162 = new_n11161 ^ new_n11149;
  assign new_n11163 = new_n11161 ^ new_n11151;
  assign new_n11164 = new_n11162 & new_n11163;
  assign new_n11165 = new_n11164 ^ new_n11155;
  assign new_n11166 = new_n11164 ^ new_n11151;
  assign new_n11167 = new_n11166 ^ new_n11165;
  assign new_n11168 = ~new_n11160 & ~new_n11167;
  assign new_n11169 = new_n11168 ^ new_n11166;
  assign new_n11170 = new_n11169 ^ new_n11157;
  assign new_n11171 = n79 & new_n7553;
  assign new_n11172 = new_n1069 & new_n7543;
  assign new_n11173 = new_n11172 ^ new_n11171;
  assign new_n11174 = n80 & new_n7542;
  assign new_n11175 = n78 & new_n7547;
  assign new_n11176 = new_n11175 ^ new_n11174;
  assign new_n11177 = new_n11176 ^ new_n11173;
  assign new_n11178 = new_n11177 ^ n57;
  assign new_n11179 = new_n10936 ^ new_n10899;
  assign new_n11180 = new_n10900 & new_n11179;
  assign new_n11181 = new_n11180 ^ new_n10896;
  assign new_n11182 = new_n11181 ^ new_n11178;
  assign new_n11183 = n6 ^ n3;
  assign new_n11184 = new_n10927 ^ n71;
  assign new_n11185 = ~new_n9495 & new_n11184;
  assign new_n11186 = new_n11185 ^ n71;
  assign new_n11187 = new_n11186 ^ new_n11183;
  assign new_n11188 = new_n10926 ^ n3;
  assign new_n11189 = new_n10930 ^ n3;
  assign new_n11190 = ~new_n11188 & new_n11189;
  assign new_n11191 = new_n11190 ^ n3;
  assign new_n11192 = new_n10927 ^ n3;
  assign new_n11193 = new_n11188 & new_n11192;
  assign new_n11194 = new_n11193 ^ n3;
  assign new_n11195 = new_n11194 ^ new_n11191;
  assign new_n11196 = ~n63 & new_n11195;
  assign new_n11197 = new_n11196 ^ new_n11191;
  assign new_n11198 = new_n11197 ^ new_n11187;
  assign new_n11199 = n73 & new_n9195;
  assign new_n11200 = new_n595 & new_n9185;
  assign new_n11201 = new_n11200 ^ new_n11199;
  assign new_n11202 = n74 & new_n9184;
  assign new_n11203 = n72 & new_n9189;
  assign new_n11204 = new_n11203 ^ new_n11202;
  assign new_n11205 = new_n11204 ^ new_n11201;
  assign new_n11206 = new_n11205 ^ n63;
  assign new_n11207 = new_n11206 ^ new_n11198;
  assign new_n11208 = n76 & new_n8355;
  assign new_n11209 = ~new_n812 & new_n8345;
  assign new_n11210 = new_n11209 ^ new_n11208;
  assign new_n11211 = n77 & new_n8344;
  assign new_n11212 = n75 & new_n8349;
  assign new_n11213 = new_n11212 ^ new_n11211;
  assign new_n11214 = new_n11213 ^ new_n11210;
  assign new_n11215 = new_n11214 ^ n60;
  assign new_n11216 = new_n11215 ^ new_n11207;
  assign new_n11217 = new_n10935 ^ new_n10918;
  assign new_n11218 = new_n10919 & new_n11217;
  assign new_n11219 = new_n11218 ^ new_n10908;
  assign new_n11220 = new_n11219 ^ new_n11216;
  assign new_n11221 = new_n11220 ^ new_n11182;
  assign new_n11222 = ~new_n6805 & n82;
  assign new_n11223 = new_n1363 & new_n6800;
  assign new_n11224 = new_n11223 ^ new_n11222;
  assign new_n11225 = n83 & new_n6799;
  assign new_n11226 = n81 & new_n6811;
  assign new_n11227 = new_n11226 ^ new_n11225;
  assign new_n11228 = new_n11227 ^ new_n11224;
  assign new_n11229 = new_n11228 ^ n54;
  assign new_n11230 = new_n11229 ^ new_n11221;
  assign new_n11231 = new_n10941 ^ new_n10937;
  assign new_n11232 = ~new_n10938 & new_n11231;
  assign new_n11233 = new_n11232 ^ new_n10888;
  assign new_n11234 = new_n11233 ^ new_n11230;
  assign new_n11235 = ~new_n6110 & n85;
  assign new_n11236 = new_n1694 & new_n6105;
  assign new_n11237 = new_n11236 ^ new_n11235;
  assign new_n11238 = n86 & new_n6104;
  assign new_n11239 = n84 & new_n6347;
  assign new_n11240 = new_n11239 ^ new_n11238;
  assign new_n11241 = new_n11240 ^ new_n11237;
  assign new_n11242 = new_n11241 ^ n51;
  assign new_n11243 = new_n11242 ^ new_n11234;
  assign new_n11244 = new_n10946 ^ new_n10880;
  assign new_n11245 = ~new_n11244 & new_n10943;
  assign new_n11246 = new_n11245 ^ new_n10946;
  assign new_n11247 = new_n11246 ^ new_n11243;
  assign new_n11248 = new_n10959 ^ new_n10947;
  assign new_n11249 = ~new_n11248 & new_n10951;
  assign new_n11250 = new_n11249 ^ new_n10950;
  assign new_n11251 = new_n11250 ^ new_n11247;
  assign new_n11252 = ~new_n5424 & n88;
  assign new_n11253 = new_n2063 & new_n5419;
  assign new_n11254 = new_n11253 ^ new_n11252;
  assign new_n11255 = n89 & new_n5418;
  assign new_n11256 = n87 & new_n5648;
  assign new_n11257 = new_n11256 ^ new_n11255;
  assign new_n11258 = new_n11257 ^ new_n11254;
  assign new_n11259 = new_n11258 ^ n48;
  assign new_n11260 = new_n11259 ^ new_n11251;
  assign new_n11261 = ~new_n4804 & n91;
  assign new_n11262 = new_n2481 & new_n4799;
  assign new_n11263 = new_n11262 ^ new_n11261;
  assign new_n11264 = n92 & new_n4798;
  assign new_n11265 = n90 & new_n4810;
  assign new_n11266 = new_n11265 ^ new_n11264;
  assign new_n11267 = new_n11266 ^ new_n11263;
  assign new_n11268 = new_n11267 ^ n45;
  assign new_n11269 = new_n11268 ^ new_n11260;
  assign new_n11270 = new_n10972 ^ new_n10960;
  assign new_n11271 = ~new_n10969 & new_n11270;
  assign new_n11272 = new_n11271 ^ new_n10972;
  assign new_n11273 = new_n11272 ^ new_n11269;
  assign new_n11274 = ~new_n4212 & n94;
  assign new_n11275 = new_n2934 & new_n4201;
  assign new_n11276 = new_n11275 ^ new_n11274;
  assign new_n11277 = n95 & new_n4200;
  assign new_n11278 = n93 & new_n4206;
  assign new_n11279 = new_n11278 ^ new_n11277;
  assign new_n11280 = new_n11279 ^ new_n11276;
  assign new_n11281 = new_n11280 ^ n42;
  assign new_n11282 = new_n11281 ^ new_n11273;
  assign new_n11283 = new_n10985 ^ new_n10973;
  assign new_n11284 = ~new_n10982 & new_n11283;
  assign new_n11285 = new_n11284 ^ new_n10985;
  assign new_n11286 = new_n11285 ^ new_n11282;
  assign new_n11287 = ~new_n3682 & n97;
  assign new_n11288 = new_n3435 & new_n3677;
  assign new_n11289 = new_n11288 ^ new_n11287;
  assign new_n11290 = n98 & new_n3676;
  assign new_n11291 = n96 & new_n3688;
  assign new_n11292 = new_n11291 ^ new_n11290;
  assign new_n11293 = new_n11292 ^ new_n11289;
  assign new_n11294 = new_n11293 ^ n39;
  assign new_n11295 = new_n11294 ^ new_n11286;
  assign new_n11296 = new_n10998 ^ new_n10986;
  assign new_n11297 = ~new_n10995 & ~new_n11296;
  assign new_n11298 = new_n11297 ^ new_n10998;
  assign new_n11299 = new_n11298 ^ new_n11295;
  assign new_n11300 = ~new_n3143 & n100;
  assign new_n11301 = new_n3138 & new_n3972;
  assign new_n11302 = new_n11301 ^ new_n11300;
  assign new_n11303 = n101 & new_n3137;
  assign new_n11304 = n99 & new_n3149;
  assign new_n11305 = new_n11304 ^ new_n11303;
  assign new_n11306 = new_n11305 ^ new_n11302;
  assign new_n11307 = new_n11306 ^ n36;
  assign new_n11308 = new_n11307 ^ new_n11299;
  assign new_n11309 = new_n11011 ^ new_n10999;
  assign new_n11310 = ~new_n11309 & new_n11008;
  assign new_n11311 = new_n11310 ^ new_n11011;
  assign new_n11312 = new_n11311 ^ new_n11308;
  assign new_n11313 = ~new_n2672 & n103;
  assign new_n11314 = ~new_n4556 & new_n2667;
  assign new_n11315 = new_n11314 ^ new_n11313;
  assign new_n11316 = n104 & new_n2666;
  assign new_n11317 = n102 & new_n2664;
  assign new_n11318 = new_n11317 ^ new_n11316;
  assign new_n11319 = new_n11318 ^ new_n11315;
  assign new_n11320 = new_n11319 ^ n33;
  assign new_n11321 = new_n11320 ^ new_n11312;
  assign new_n11322 = new_n11024 ^ new_n11012;
  assign new_n11323 = ~new_n11322 & new_n11021;
  assign new_n11324 = new_n11323 ^ new_n11024;
  assign new_n11325 = new_n11324 ^ new_n11321;
  assign new_n11326 = n106 & new_n2246;
  assign new_n11327 = ~new_n5164 & new_n2241;
  assign new_n11328 = new_n11327 ^ new_n11326;
  assign new_n11329 = n107 & new_n2240;
  assign new_n11330 = n105 & new_n2391;
  assign new_n11331 = new_n11330 ^ new_n11329;
  assign new_n11332 = new_n11331 ^ new_n11328;
  assign new_n11333 = new_n11332 ^ n30;
  assign new_n11334 = new_n11333 ^ new_n11325;
  assign new_n11335 = new_n11037 ^ new_n11025;
  assign new_n11336 = ~new_n11335 & new_n11034;
  assign new_n11337 = new_n11336 ^ new_n11037;
  assign new_n11338 = new_n11337 ^ new_n11334;
  assign new_n11339 = n109 & new_n1874;
  assign new_n11340 = new_n1864 & new_n5825;
  assign new_n11341 = new_n11340 ^ new_n11339;
  assign new_n11342 = n110 & new_n1863;
  assign new_n11343 = n108 & new_n1868;
  assign new_n11344 = new_n11343 ^ new_n11342;
  assign new_n11345 = new_n11344 ^ new_n11341;
  assign new_n11346 = new_n11345 ^ n27;
  assign new_n11347 = new_n11346 ^ new_n11338;
  assign new_n11348 = new_n11050 ^ new_n11038;
  assign new_n11349 = ~new_n11348 & new_n11047;
  assign new_n11350 = new_n11349 ^ new_n11050;
  assign new_n11351 = new_n11350 ^ new_n11347;
  assign new_n11352 = ~new_n1506 & n112;
  assign new_n11353 = ~new_n6518 & new_n1501;
  assign new_n11354 = new_n11353 ^ new_n11352;
  assign new_n11355 = n113 & new_n1500;
  assign new_n11356 = n111 & new_n1512;
  assign new_n11357 = new_n11356 ^ new_n11355;
  assign new_n11358 = new_n11357 ^ new_n11354;
  assign new_n11359 = new_n11358 ^ n24;
  assign new_n11360 = new_n11359 ^ new_n11351;
  assign new_n11361 = new_n11063 ^ new_n11051;
  assign new_n11362 = new_n11060 & new_n11361;
  assign new_n11363 = new_n11362 ^ new_n11063;
  assign new_n11364 = new_n11363 ^ new_n11360;
  assign new_n11365 = ~new_n1198 & n115;
  assign new_n11366 = ~new_n7256 & new_n1193;
  assign new_n11367 = new_n11366 ^ new_n11365;
  assign new_n11368 = n116 & new_n1192;
  assign new_n11369 = n114 & new_n1204;
  assign new_n11370 = new_n11369 ^ new_n11368;
  assign new_n11371 = new_n11370 ^ new_n11367;
  assign new_n11372 = new_n11371 ^ n21;
  assign new_n11373 = new_n11372 ^ new_n11364;
  assign new_n11374 = new_n11076 ^ new_n11064;
  assign new_n11375 = ~new_n11073 & new_n11374;
  assign new_n11376 = new_n11375 ^ new_n11076;
  assign new_n11377 = new_n11376 ^ new_n11373;
  assign new_n11378 = ~new_n930 & n118;
  assign new_n11379 = ~new_n8019 & new_n925;
  assign new_n11380 = new_n11379 ^ new_n11378;
  assign new_n11381 = n119 & new_n924;
  assign new_n11382 = n117 & new_n936;
  assign new_n11383 = new_n11382 ^ new_n11381;
  assign new_n11384 = new_n11383 ^ new_n11380;
  assign new_n11385 = new_n11384 ^ n18;
  assign new_n11386 = new_n11385 ^ new_n11377;
  assign new_n11387 = new_n11089 ^ new_n11077;
  assign new_n11388 = ~new_n11086 & new_n11387;
  assign new_n11389 = new_n11388 ^ new_n11089;
  assign new_n11390 = new_n11389 ^ new_n11386;
  assign new_n11391 = n121 & new_n707;
  assign new_n11392 = new_n701 & new_n8850;
  assign new_n11393 = new_n11392 ^ new_n11391;
  assign new_n11394 = n122 & new_n700;
  assign new_n11395 = n120 & new_n787;
  assign new_n11396 = new_n11395 ^ new_n11394;
  assign new_n11397 = new_n11396 ^ new_n11393;
  assign new_n11398 = new_n11397 ^ n15;
  assign new_n11399 = new_n11398 ^ new_n11390;
  assign new_n11400 = new_n11102 ^ new_n11090;
  assign new_n11401 = ~new_n11099 & new_n11400;
  assign new_n11402 = new_n11401 ^ new_n11102;
  assign new_n11403 = new_n11402 ^ new_n11399;
  assign new_n11404 = n124 & new_n499;
  assign new_n11405 = ~new_n506 & new_n9700;
  assign new_n11406 = new_n11405 ^ new_n11404;
  assign new_n11407 = ~new_n505 & n125;
  assign new_n11408 = n123 & new_n579;
  assign new_n11409 = new_n11408 ^ new_n11407;
  assign new_n11410 = new_n11409 ^ new_n11406;
  assign new_n11411 = new_n11410 ^ n12;
  assign new_n11412 = new_n11411 ^ new_n11403;
  assign new_n11413 = new_n11115 ^ new_n11103;
  assign new_n11414 = ~new_n11112 & new_n11413;
  assign new_n11415 = new_n11414 ^ new_n11115;
  assign new_n11416 = new_n11415 ^ new_n11412;
  assign new_n11417 = n127 & new_n354;
  assign new_n11418 = new_n349 & new_n10581;
  assign new_n11419 = new_n11418 ^ new_n11417;
  assign new_n11420 = n128 & new_n348;
  assign new_n11421 = n126 & new_n391;
  assign new_n11422 = new_n11421 ^ new_n11420;
  assign new_n11423 = new_n11422 ^ new_n11419;
  assign new_n11424 = new_n11423 ^ n9;
  assign new_n11425 = new_n11424 ^ new_n11416;
  assign new_n11426 = new_n11128 ^ new_n11116;
  assign new_n11427 = ~new_n11125 & new_n11426;
  assign new_n11428 = new_n11427 ^ new_n11128;
  assign new_n11429 = new_n11428 ^ new_n11425;
  assign new_n11430 = new_n11429 ^ new_n11170;
  assign new_n11431 = ~new_n11429 & new_n11153;
  assign new_n11432 = ~new_n11431 & new_n11149;
  assign new_n11433 = ~new_n11151 & new_n11160;
  assign new_n11434 = new_n11429 & new_n11433;
  assign new_n11435 = new_n11434 ^ new_n11160;
  assign new_n11436 = ~new_n11432 & new_n11435;
  assign new_n11437 = ~new_n11429 & new_n11159;
  assign new_n11438 = ~new_n11436 & ~new_n11437;
  assign new_n11439 = ~new_n11151 & new_n11149;
  assign new_n11440 = ~new_n11161 & ~new_n11431;
  assign new_n11441 = ~new_n11439 & ~new_n11440;
  assign new_n11442 = ~new_n11441 & new_n11438;
  assign new_n11443 = ~new_n4804 & n92;
  assign new_n11444 = new_n2628 & new_n4799;
  assign new_n11445 = new_n11444 ^ new_n11443;
  assign new_n11446 = n93 & new_n4798;
  assign new_n11447 = n91 & new_n4810;
  assign new_n11448 = new_n11447 ^ new_n11446;
  assign new_n11449 = new_n11448 ^ new_n11445;
  assign new_n11450 = new_n11449 ^ n45;
  assign new_n11451 = ~new_n5424 & n89;
  assign new_n11452 = new_n2193 & new_n5419;
  assign new_n11453 = new_n11452 ^ new_n11451;
  assign new_n11454 = n90 & new_n5418;
  assign new_n11455 = n88 & new_n5648;
  assign new_n11456 = new_n11455 ^ new_n11454;
  assign new_n11457 = new_n11456 ^ new_n11453;
  assign new_n11458 = new_n11457 ^ n48;
  assign new_n11459 = ~new_n6110 & n86;
  assign new_n11460 = new_n1811 & new_n6105;
  assign new_n11461 = new_n11460 ^ new_n11459;
  assign new_n11462 = n87 & new_n6104;
  assign new_n11463 = n85 & new_n6347;
  assign new_n11464 = new_n11463 ^ new_n11462;
  assign new_n11465 = new_n11464 ^ new_n11461;
  assign new_n11466 = new_n11465 ^ n51;
  assign new_n11467 = ~new_n6805 & n83;
  assign new_n11468 = new_n1468 & new_n6800;
  assign new_n11469 = new_n11468 ^ new_n11467;
  assign new_n11470 = n84 & new_n6799;
  assign new_n11471 = n82 & new_n6811;
  assign new_n11472 = new_n11471 ^ new_n11470;
  assign new_n11473 = new_n11472 ^ new_n11469;
  assign new_n11474 = new_n11473 ^ n54;
  assign new_n11475 = n77 & new_n8355;
  assign new_n11476 = ~new_n891 & new_n8345;
  assign new_n11477 = new_n11476 ^ new_n11475;
  assign new_n11478 = n78 & new_n8344;
  assign new_n11479 = n76 & new_n8349;
  assign new_n11480 = new_n11479 ^ new_n11478;
  assign new_n11481 = new_n11480 ^ new_n11477;
  assign new_n11482 = new_n11481 ^ n60;
  assign new_n11483 = n74 & new_n9195;
  assign new_n11484 = new_n660 & new_n9185;
  assign new_n11485 = new_n11484 ^ new_n11483;
  assign new_n11486 = n75 & new_n9184;
  assign new_n11487 = n73 & new_n9189;
  assign new_n11488 = new_n11487 ^ new_n11486;
  assign new_n11489 = new_n11488 ^ new_n11485;
  assign new_n11490 = new_n11489 ^ n63;
  assign new_n11491 = ~n64 & n63;
  assign new_n11492 = new_n11491 ^ n63;
  assign new_n11493 = n71 & new_n11492;
  assign new_n11494 = n72 & new_n9495;
  assign new_n11495 = new_n11494 ^ new_n11493;
  assign new_n11496 = new_n11186 ^ n6;
  assign new_n11497 = new_n11183 & new_n11496;
  assign new_n11498 = new_n11497 ^ n3;
  assign new_n11499 = new_n11498 ^ new_n11495;
  assign new_n11500 = new_n11499 ^ new_n11490;
  assign new_n11501 = new_n11500 ^ new_n11482;
  assign new_n11502 = new_n11206 ^ new_n11187;
  assign new_n11503 = ~new_n11502 & new_n11198;
  assign new_n11504 = new_n11503 ^ new_n11197;
  assign new_n11505 = new_n11504 ^ new_n11501;
  assign new_n11506 = n80 & new_n7553;
  assign new_n11507 = new_n1161 & new_n7543;
  assign new_n11508 = new_n11507 ^ new_n11506;
  assign new_n11509 = n81 & new_n7542;
  assign new_n11510 = n79 & new_n7547;
  assign new_n11511 = new_n11510 ^ new_n11509;
  assign new_n11512 = new_n11511 ^ new_n11508;
  assign new_n11513 = new_n11512 ^ n57;
  assign new_n11514 = new_n11513 ^ new_n11505;
  assign new_n11515 = new_n11219 ^ new_n11207;
  assign new_n11516 = ~new_n11216 & new_n11515;
  assign new_n11517 = new_n11516 ^ new_n11219;
  assign new_n11518 = new_n11517 ^ new_n11514;
  assign new_n11519 = new_n11518 ^ new_n11474;
  assign new_n11520 = new_n11220 ^ new_n11178;
  assign new_n11521 = ~new_n11520 & new_n11182;
  assign new_n11522 = new_n11521 ^ new_n11181;
  assign new_n11523 = new_n11522 ^ new_n11519;
  assign new_n11524 = new_n11523 ^ new_n11466;
  assign new_n11525 = new_n11233 ^ new_n11229;
  assign new_n11526 = ~new_n11525 & new_n11230;
  assign new_n11527 = new_n11526 ^ new_n11221;
  assign new_n11528 = new_n11527 ^ new_n11524;
  assign new_n11529 = new_n11528 ^ new_n11458;
  assign new_n11530 = new_n11246 ^ new_n11234;
  assign new_n11531 = ~new_n11243 & ~new_n11530;
  assign new_n11532 = new_n11531 ^ new_n11246;
  assign new_n11533 = new_n11532 ^ new_n11529;
  assign new_n11534 = new_n11533 ^ new_n11450;
  assign new_n11535 = new_n11259 ^ new_n11247;
  assign new_n11536 = ~new_n11251 & new_n11535;
  assign new_n11537 = new_n11536 ^ new_n11250;
  assign new_n11538 = new_n11537 ^ new_n11534;
  assign new_n11539 = ~new_n4212 & n95;
  assign new_n11540 = new_n3095 & new_n4201;
  assign new_n11541 = new_n11540 ^ new_n11539;
  assign new_n11542 = n96 & new_n4200;
  assign new_n11543 = n94 & new_n4206;
  assign new_n11544 = new_n11543 ^ new_n11542;
  assign new_n11545 = new_n11544 ^ new_n11541;
  assign new_n11546 = new_n11545 ^ n42;
  assign new_n11547 = new_n11546 ^ new_n11538;
  assign new_n11548 = new_n11272 ^ new_n11260;
  assign new_n11549 = ~new_n11548 & new_n11269;
  assign new_n11550 = new_n11549 ^ new_n11272;
  assign new_n11551 = new_n11550 ^ new_n11547;
  assign new_n11552 = ~new_n3682 & n98;
  assign new_n11553 = new_n3604 & new_n3677;
  assign new_n11554 = new_n11553 ^ new_n11552;
  assign new_n11555 = n99 & new_n3676;
  assign new_n11556 = n97 & new_n3688;
  assign new_n11557 = new_n11556 ^ new_n11555;
  assign new_n11558 = new_n11557 ^ new_n11554;
  assign new_n11559 = new_n11558 ^ n39;
  assign new_n11560 = new_n11559 ^ new_n11551;
  assign new_n11561 = new_n11285 ^ new_n11273;
  assign new_n11562 = ~new_n11561 & new_n11282;
  assign new_n11563 = new_n11562 ^ new_n11285;
  assign new_n11564 = new_n11563 ^ new_n11560;
  assign new_n11565 = ~new_n3143 & n101;
  assign new_n11566 = new_n3138 & new_n4159;
  assign new_n11567 = new_n11566 ^ new_n11565;
  assign new_n11568 = n102 & new_n3137;
  assign new_n11569 = n100 & new_n3149;
  assign new_n11570 = new_n11569 ^ new_n11568;
  assign new_n11571 = new_n11570 ^ new_n11567;
  assign new_n11572 = new_n11571 ^ n36;
  assign new_n11573 = new_n11572 ^ new_n11564;
  assign new_n11574 = new_n11298 ^ new_n11286;
  assign new_n11575 = new_n11295 & new_n11574;
  assign new_n11576 = new_n11575 ^ new_n11298;
  assign new_n11577 = new_n11576 ^ new_n11573;
  assign new_n11578 = ~new_n2672 & n104;
  assign new_n11579 = ~new_n4754 & new_n2667;
  assign new_n11580 = new_n11579 ^ new_n11578;
  assign new_n11581 = n105 & new_n2666;
  assign new_n11582 = n103 & new_n2664;
  assign new_n11583 = new_n11582 ^ new_n11581;
  assign new_n11584 = new_n11583 ^ new_n11580;
  assign new_n11585 = new_n11584 ^ n33;
  assign new_n11586 = new_n11585 ^ new_n11577;
  assign new_n11587 = new_n11311 ^ new_n11299;
  assign new_n11588 = ~new_n11308 & new_n11587;
  assign new_n11589 = new_n11588 ^ new_n11311;
  assign new_n11590 = new_n11589 ^ new_n11586;
  assign new_n11591 = n107 & new_n2246;
  assign new_n11592 = ~new_n5377 & new_n2241;
  assign new_n11593 = new_n11592 ^ new_n11591;
  assign new_n11594 = n108 & new_n2240;
  assign new_n11595 = n106 & new_n2391;
  assign new_n11596 = new_n11595 ^ new_n11594;
  assign new_n11597 = new_n11596 ^ new_n11593;
  assign new_n11598 = new_n11597 ^ n30;
  assign new_n11599 = new_n11598 ^ new_n11590;
  assign new_n11600 = new_n11324 ^ new_n11312;
  assign new_n11601 = ~new_n11321 & new_n11600;
  assign new_n11602 = new_n11601 ^ new_n11324;
  assign new_n11603 = new_n11602 ^ new_n11599;
  assign new_n11604 = n110 & new_n1874;
  assign new_n11605 = new_n1864 & new_n6049;
  assign new_n11606 = new_n11605 ^ new_n11604;
  assign new_n11607 = n111 & new_n1863;
  assign new_n11608 = n109 & new_n1868;
  assign new_n11609 = new_n11608 ^ new_n11607;
  assign new_n11610 = new_n11609 ^ new_n11606;
  assign new_n11611 = new_n11610 ^ n27;
  assign new_n11612 = new_n11611 ^ new_n11603;
  assign new_n11613 = new_n11337 ^ new_n11325;
  assign new_n11614 = ~new_n11334 & new_n11613;
  assign new_n11615 = new_n11614 ^ new_n11337;
  assign new_n11616 = new_n11615 ^ new_n11612;
  assign new_n11617 = ~new_n1506 & n113;
  assign new_n11618 = ~new_n6764 & new_n1501;
  assign new_n11619 = new_n11618 ^ new_n11617;
  assign new_n11620 = n114 & new_n1500;
  assign new_n11621 = n112 & new_n1512;
  assign new_n11622 = new_n11621 ^ new_n11620;
  assign new_n11623 = new_n11622 ^ new_n11619;
  assign new_n11624 = new_n11623 ^ n24;
  assign new_n11625 = new_n11624 ^ new_n11616;
  assign new_n11626 = new_n11350 ^ new_n11338;
  assign new_n11627 = ~new_n11347 & new_n11626;
  assign new_n11628 = new_n11627 ^ new_n11350;
  assign new_n11629 = new_n11628 ^ new_n11625;
  assign new_n11630 = ~new_n1198 & n116;
  assign new_n11631 = ~new_n7503 & new_n1193;
  assign new_n11632 = new_n11631 ^ new_n11630;
  assign new_n11633 = n117 & new_n1192;
  assign new_n11634 = n115 & new_n1204;
  assign new_n11635 = new_n11634 ^ new_n11633;
  assign new_n11636 = new_n11635 ^ new_n11632;
  assign new_n11637 = new_n11636 ^ n21;
  assign new_n11638 = new_n11637 ^ new_n11629;
  assign new_n11639 = new_n11363 ^ new_n11351;
  assign new_n11640 = ~new_n11360 & ~new_n11639;
  assign new_n11641 = new_n11640 ^ new_n11363;
  assign new_n11642 = new_n11641 ^ new_n11638;
  assign new_n11643 = ~new_n930 & n119;
  assign new_n11644 = new_n925 & new_n8286;
  assign new_n11645 = new_n11644 ^ new_n11643;
  assign new_n11646 = n120 & new_n924;
  assign new_n11647 = n118 & new_n936;
  assign new_n11648 = new_n11647 ^ new_n11646;
  assign new_n11649 = new_n11648 ^ new_n11645;
  assign new_n11650 = new_n11649 ^ n18;
  assign new_n11651 = new_n11650 ^ new_n11642;
  assign new_n11652 = new_n11376 ^ new_n11364;
  assign new_n11653 = ~new_n11652 & new_n11373;
  assign new_n11654 = new_n11653 ^ new_n11376;
  assign new_n11655 = new_n11654 ^ new_n11651;
  assign new_n11656 = n122 & new_n707;
  assign new_n11657 = ~new_n9116 & new_n701;
  assign new_n11658 = new_n11657 ^ new_n11656;
  assign new_n11659 = n123 & new_n700;
  assign new_n11660 = n121 & new_n787;
  assign new_n11661 = new_n11660 ^ new_n11659;
  assign new_n11662 = new_n11661 ^ new_n11658;
  assign new_n11663 = new_n11662 ^ n15;
  assign new_n11664 = new_n11663 ^ new_n11655;
  assign new_n11665 = new_n11389 ^ new_n11377;
  assign new_n11666 = ~new_n11665 & new_n11386;
  assign new_n11667 = new_n11666 ^ new_n11389;
  assign new_n11668 = new_n11667 ^ new_n11664;
  assign new_n11669 = n125 & new_n499;
  assign new_n11670 = ~new_n506 & new_n9987;
  assign new_n11671 = new_n11670 ^ new_n11669;
  assign new_n11672 = ~new_n505 & n126;
  assign new_n11673 = n124 & new_n579;
  assign new_n11674 = new_n11673 ^ new_n11672;
  assign new_n11675 = new_n11674 ^ new_n11671;
  assign new_n11676 = new_n11675 ^ n12;
  assign new_n11677 = new_n11676 ^ new_n11668;
  assign new_n11678 = new_n11402 ^ new_n11390;
  assign new_n11679 = ~new_n11678 & new_n11399;
  assign new_n11680 = new_n11679 ^ new_n11402;
  assign new_n11681 = new_n11680 ^ new_n11677;
  assign new_n11682 = n127 & new_n391;
  assign new_n11683 = new_n349 & new_n10010;
  assign new_n11684 = new_n11683 ^ new_n11682;
  assign new_n11685 = n128 & new_n354;
  assign new_n11686 = new_n11685 ^ new_n11684;
  assign new_n11687 = new_n11686 ^ n9;
  assign new_n11688 = new_n11687 ^ new_n11681;
  assign new_n11689 = new_n11415 ^ new_n11403;
  assign new_n11690 = ~new_n11689 & new_n11412;
  assign new_n11691 = new_n11690 ^ new_n11415;
  assign new_n11692 = new_n11691 ^ new_n11688;
  assign new_n11693 = new_n11428 ^ new_n11416;
  assign new_n11694 = ~new_n11693 & new_n11425;
  assign new_n11695 = new_n11694 ^ new_n11428;
  assign new_n11696 = new_n11695 ^ new_n11692;
  assign new_n11697 = new_n11696 ^ new_n11442;
  assign new_n11698 = new_n290 ^ n9;
  assign new_n11699 = new_n291 ^ new_n290;
  assign new_n11700 = new_n347 ^ new_n291;
  assign new_n11701 = new_n291 & new_n11700;
  assign new_n11702 = new_n11701 ^ new_n291;
  assign new_n11703 = ~new_n11699 & new_n11702;
  assign new_n11704 = new_n11703 ^ new_n11701;
  assign new_n11705 = new_n11704 ^ new_n291;
  assign new_n11706 = new_n11705 ^ new_n347;
  assign new_n11707 = ~new_n11698 & new_n11706;
  assign new_n11708 = new_n11707 ^ n9;
  assign new_n11709 = new_n11708 ^ n9;
  assign new_n11710 = new_n11698 & new_n11706;
  assign new_n11711 = new_n11710 ^ n8;
  assign new_n11712 = new_n11711 ^ n9;
  assign new_n11713 = new_n11712 ^ new_n11709;
  assign new_n11714 = new_n11712 ^ new_n10009;
  assign new_n11715 = new_n11714 ^ new_n11712;
  assign new_n11716 = new_n11713 & new_n11715;
  assign new_n11717 = new_n11716 ^ new_n11712;
  assign new_n11718 = n128 & new_n11717;
  assign new_n11719 = new_n11718 ^ n9;
  assign new_n11720 = ~new_n4212 & n96;
  assign new_n11721 = new_n3273 & new_n4201;
  assign new_n11722 = new_n11721 ^ new_n11720;
  assign new_n11723 = n97 & new_n4200;
  assign new_n11724 = n95 & new_n4206;
  assign new_n11725 = new_n11724 ^ new_n11723;
  assign new_n11726 = new_n11725 ^ new_n11722;
  assign new_n11727 = new_n11726 ^ n42;
  assign new_n11728 = ~new_n4804 & n93;
  assign new_n11729 = new_n2785 & new_n4799;
  assign new_n11730 = new_n11729 ^ new_n11728;
  assign new_n11731 = n94 & new_n4798;
  assign new_n11732 = n92 & new_n4810;
  assign new_n11733 = new_n11732 ^ new_n11731;
  assign new_n11734 = new_n11733 ^ new_n11730;
  assign new_n11735 = new_n11734 ^ n45;
  assign new_n11736 = ~new_n5424 & n90;
  assign new_n11737 = new_n2341 & new_n5419;
  assign new_n11738 = new_n11737 ^ new_n11736;
  assign new_n11739 = n91 & new_n5418;
  assign new_n11740 = n89 & new_n5648;
  assign new_n11741 = new_n11740 ^ new_n11739;
  assign new_n11742 = new_n11741 ^ new_n11738;
  assign new_n11743 = new_n11742 ^ n48;
  assign new_n11744 = new_n11527 ^ new_n11466;
  assign new_n11745 = ~new_n11524 & new_n11744;
  assign new_n11746 = new_n11745 ^ new_n11527;
  assign new_n11747 = new_n11746 ^ new_n11743;
  assign new_n11748 = ~new_n6110 & n87;
  assign new_n11749 = new_n1940 & new_n6105;
  assign new_n11750 = new_n11749 ^ new_n11748;
  assign new_n11751 = n88 & new_n6104;
  assign new_n11752 = n86 & new_n6347;
  assign new_n11753 = new_n11752 ^ new_n11751;
  assign new_n11754 = new_n11753 ^ new_n11750;
  assign new_n11755 = new_n11754 ^ n51;
  assign new_n11756 = ~new_n6805 & n84;
  assign new_n11757 = new_n1584 & new_n6800;
  assign new_n11758 = new_n11757 ^ new_n11756;
  assign new_n11759 = n85 & new_n6799;
  assign new_n11760 = n83 & new_n6811;
  assign new_n11761 = new_n11760 ^ new_n11759;
  assign new_n11762 = new_n11761 ^ new_n11758;
  assign new_n11763 = new_n11762 ^ n54;
  assign new_n11764 = n78 & new_n8355;
  assign new_n11765 = ~new_n982 & new_n8345;
  assign new_n11766 = new_n11765 ^ new_n11764;
  assign new_n11767 = n79 & new_n8344;
  assign new_n11768 = n77 & new_n8349;
  assign new_n11769 = new_n11768 ^ new_n11767;
  assign new_n11770 = new_n11769 ^ new_n11766;
  assign new_n11771 = new_n11770 ^ n60;
  assign new_n11772 = n75 & new_n9195;
  assign new_n11773 = ~new_n737 & new_n9185;
  assign new_n11774 = new_n11773 ^ new_n11772;
  assign new_n11775 = n76 & new_n9184;
  assign new_n11776 = n74 & new_n9189;
  assign new_n11777 = new_n11776 ^ new_n11775;
  assign new_n11778 = new_n11777 ^ new_n11774;
  assign new_n11779 = new_n11778 ^ n63;
  assign new_n11780 = new_n11779 ^ new_n11771;
  assign new_n11781 = new_n11498 ^ new_n11490;
  assign new_n11782 = ~new_n11499 & ~new_n11781;
  assign new_n11783 = new_n11782 ^ new_n11490;
  assign new_n11784 = ~n73 & new_n9495;
  assign new_n11785 = new_n11784 ^ new_n11493;
  assign new_n11786 = n72 & new_n11785;
  assign new_n11787 = new_n11786 ^ new_n11493;
  assign new_n11788 = new_n9495 ^ n72;
  assign new_n11789 = new_n11491 ^ n64;
  assign new_n11790 = new_n11789 ^ n71;
  assign new_n11791 = new_n11790 ^ new_n11785;
  assign new_n11792 = new_n11791 ^ n71;
  assign new_n11793 = new_n11788 & new_n11792;
  assign new_n11794 = new_n11793 ^ new_n420;
  assign new_n11795 = new_n11794 ^ new_n11787;
  assign new_n11796 = new_n11795 ^ new_n420;
  assign new_n11797 = new_n11796 ^ new_n11783;
  assign new_n11798 = new_n11797 ^ new_n11780;
  assign new_n11799 = n81 & new_n7553;
  assign new_n11800 = new_n1263 & new_n7543;
  assign new_n11801 = new_n11800 ^ new_n11799;
  assign new_n11802 = n82 & new_n7542;
  assign new_n11803 = n80 & new_n7547;
  assign new_n11804 = new_n11803 ^ new_n11802;
  assign new_n11805 = new_n11804 ^ new_n11801;
  assign new_n11806 = new_n11805 ^ n57;
  assign new_n11807 = new_n11806 ^ new_n11798;
  assign new_n11808 = new_n11504 ^ new_n11482;
  assign new_n11809 = ~new_n11501 & new_n11808;
  assign new_n11810 = new_n11809 ^ new_n11504;
  assign new_n11811 = new_n11810 ^ new_n11807;
  assign new_n11812 = new_n11811 ^ new_n11763;
  assign new_n11813 = new_n11517 ^ new_n11505;
  assign new_n11814 = ~new_n11514 & new_n11813;
  assign new_n11815 = new_n11814 ^ new_n11517;
  assign new_n11816 = new_n11815 ^ new_n11812;
  assign new_n11817 = new_n11816 ^ new_n11755;
  assign new_n11818 = new_n11522 ^ new_n11474;
  assign new_n11819 = ~new_n11519 & new_n11818;
  assign new_n11820 = new_n11819 ^ new_n11522;
  assign new_n11821 = new_n11820 ^ new_n11817;
  assign new_n11822 = new_n11821 ^ new_n11747;
  assign new_n11823 = new_n11822 ^ new_n11735;
  assign new_n11824 = new_n11532 ^ new_n11528;
  assign new_n11825 = new_n11529 & new_n11824;
  assign new_n11826 = new_n11825 ^ new_n11458;
  assign new_n11827 = new_n11826 ^ new_n11823;
  assign new_n11828 = new_n11827 ^ new_n11727;
  assign new_n11829 = new_n11537 ^ new_n11450;
  assign new_n11830 = new_n11534 & new_n11829;
  assign new_n11831 = new_n11830 ^ new_n11537;
  assign new_n11832 = new_n11831 ^ new_n11828;
  assign new_n11833 = ~new_n3682 & n99;
  assign new_n11834 = new_n3677 & new_n3789;
  assign new_n11835 = new_n11834 ^ new_n11833;
  assign new_n11836 = n100 & new_n3676;
  assign new_n11837 = n98 & new_n3688;
  assign new_n11838 = new_n11837 ^ new_n11836;
  assign new_n11839 = new_n11838 ^ new_n11835;
  assign new_n11840 = new_n11839 ^ n39;
  assign new_n11841 = new_n11840 ^ new_n11832;
  assign new_n11842 = new_n11550 ^ new_n11538;
  assign new_n11843 = ~new_n11842 & new_n11547;
  assign new_n11844 = new_n11843 ^ new_n11550;
  assign new_n11845 = new_n11844 ^ new_n11841;
  assign new_n11846 = ~new_n3143 & n102;
  assign new_n11847 = new_n3138 & new_n4368;
  assign new_n11848 = new_n11847 ^ new_n11846;
  assign new_n11849 = n103 & new_n3137;
  assign new_n11850 = n101 & new_n3149;
  assign new_n11851 = new_n11850 ^ new_n11849;
  assign new_n11852 = new_n11851 ^ new_n11848;
  assign new_n11853 = new_n11852 ^ n36;
  assign new_n11854 = new_n11853 ^ new_n11845;
  assign new_n11855 = new_n11563 ^ new_n11551;
  assign new_n11856 = ~new_n11855 & new_n11560;
  assign new_n11857 = new_n11856 ^ new_n11563;
  assign new_n11858 = new_n11857 ^ new_n11854;
  assign new_n11859 = ~new_n2672 & n105;
  assign new_n11860 = ~new_n4961 & new_n2667;
  assign new_n11861 = new_n11860 ^ new_n11859;
  assign new_n11862 = n106 & new_n2666;
  assign new_n11863 = n104 & new_n2664;
  assign new_n11864 = new_n11863 ^ new_n11862;
  assign new_n11865 = new_n11864 ^ new_n11861;
  assign new_n11866 = new_n11865 ^ n33;
  assign new_n11867 = new_n11866 ^ new_n11858;
  assign new_n11868 = new_n11576 ^ new_n11564;
  assign new_n11869 = new_n11573 & new_n11868;
  assign new_n11870 = new_n11869 ^ new_n11576;
  assign new_n11871 = new_n11870 ^ new_n11867;
  assign new_n11872 = n108 & new_n2246;
  assign new_n11873 = new_n2241 & new_n5604;
  assign new_n11874 = new_n11873 ^ new_n11872;
  assign new_n11875 = n109 & new_n2240;
  assign new_n11876 = n107 & new_n2391;
  assign new_n11877 = new_n11876 ^ new_n11875;
  assign new_n11878 = new_n11877 ^ new_n11874;
  assign new_n11879 = new_n11878 ^ n30;
  assign new_n11880 = new_n11879 ^ new_n11871;
  assign new_n11881 = new_n11589 ^ new_n11577;
  assign new_n11882 = ~new_n11586 & new_n11881;
  assign new_n11883 = new_n11882 ^ new_n11589;
  assign new_n11884 = new_n11883 ^ new_n11880;
  assign new_n11885 = n111 & new_n1874;
  assign new_n11886 = ~new_n6284 & new_n1864;
  assign new_n11887 = new_n11886 ^ new_n11885;
  assign new_n11888 = n112 & new_n1863;
  assign new_n11889 = n110 & new_n1868;
  assign new_n11890 = new_n11889 ^ new_n11888;
  assign new_n11891 = new_n11890 ^ new_n11887;
  assign new_n11892 = new_n11891 ^ n27;
  assign new_n11893 = new_n11892 ^ new_n11884;
  assign new_n11894 = new_n11602 ^ new_n11590;
  assign new_n11895 = ~new_n11599 & new_n11894;
  assign new_n11896 = new_n11895 ^ new_n11602;
  assign new_n11897 = new_n11896 ^ new_n11893;
  assign new_n11898 = ~new_n1506 & n114;
  assign new_n11899 = ~new_n7013 & new_n1501;
  assign new_n11900 = new_n11899 ^ new_n11898;
  assign new_n11901 = n115 & new_n1500;
  assign new_n11902 = n113 & new_n1512;
  assign new_n11903 = new_n11902 ^ new_n11901;
  assign new_n11904 = new_n11903 ^ new_n11900;
  assign new_n11905 = new_n11904 ^ n24;
  assign new_n11906 = new_n11905 ^ new_n11897;
  assign new_n11907 = new_n11615 ^ new_n11603;
  assign new_n11908 = ~new_n11612 & new_n11907;
  assign new_n11909 = new_n11908 ^ new_n11615;
  assign new_n11910 = new_n11909 ^ new_n11906;
  assign new_n11911 = ~new_n1198 & n117;
  assign new_n11912 = ~new_n7761 & new_n1193;
  assign new_n11913 = new_n11912 ^ new_n11911;
  assign new_n11914 = n118 & new_n1192;
  assign new_n11915 = n116 & new_n1204;
  assign new_n11916 = new_n11915 ^ new_n11914;
  assign new_n11917 = new_n11916 ^ new_n11913;
  assign new_n11918 = new_n11917 ^ n21;
  assign new_n11919 = new_n11918 ^ new_n11910;
  assign new_n11920 = new_n11628 ^ new_n11616;
  assign new_n11921 = ~new_n11625 & new_n11920;
  assign new_n11922 = new_n11921 ^ new_n11628;
  assign new_n11923 = new_n11922 ^ new_n11919;
  assign new_n11924 = ~new_n930 & n120;
  assign new_n11925 = new_n925 & new_n8560;
  assign new_n11926 = new_n11925 ^ new_n11924;
  assign new_n11927 = n121 & new_n924;
  assign new_n11928 = n119 & new_n936;
  assign new_n11929 = new_n11928 ^ new_n11927;
  assign new_n11930 = new_n11929 ^ new_n11926;
  assign new_n11931 = new_n11930 ^ n18;
  assign new_n11932 = new_n11931 ^ new_n11923;
  assign new_n11933 = new_n11641 ^ new_n11629;
  assign new_n11934 = ~new_n11638 & ~new_n11933;
  assign new_n11935 = new_n11934 ^ new_n11641;
  assign new_n11936 = new_n11935 ^ new_n11932;
  assign new_n11937 = n123 & new_n707;
  assign new_n11938 = ~new_n9405 & new_n701;
  assign new_n11939 = new_n11938 ^ new_n11937;
  assign new_n11940 = n124 & new_n700;
  assign new_n11941 = n122 & new_n787;
  assign new_n11942 = new_n11941 ^ new_n11940;
  assign new_n11943 = new_n11942 ^ new_n11939;
  assign new_n11944 = new_n11943 ^ n15;
  assign new_n11945 = new_n11944 ^ new_n11936;
  assign new_n11946 = new_n11654 ^ new_n11642;
  assign new_n11947 = ~new_n11946 & new_n11651;
  assign new_n11948 = new_n11947 ^ new_n11654;
  assign new_n11949 = new_n11948 ^ new_n11945;
  assign new_n11950 = n126 & new_n499;
  assign new_n11951 = ~new_n506 & new_n10304;
  assign new_n11952 = new_n11951 ^ new_n11950;
  assign new_n11953 = ~new_n505 & n127;
  assign new_n11954 = n125 & new_n579;
  assign new_n11955 = new_n11954 ^ new_n11953;
  assign new_n11956 = new_n11955 ^ new_n11952;
  assign new_n11957 = new_n11956 ^ n12;
  assign new_n11958 = new_n11957 ^ new_n11949;
  assign new_n11959 = new_n11667 ^ new_n11663;
  assign new_n11960 = ~new_n11664 & ~new_n11959;
  assign new_n11961 = new_n11960 ^ new_n11655;
  assign new_n11962 = new_n11961 ^ new_n11958;
  assign new_n11963 = new_n11962 ^ new_n11719;
  assign new_n11964 = new_n11680 ^ new_n11668;
  assign new_n11965 = ~new_n11964 & new_n11677;
  assign new_n11966 = new_n11965 ^ new_n11680;
  assign new_n11967 = new_n11966 ^ new_n11963;
  assign new_n11968 = new_n11691 ^ new_n11681;
  assign new_n11969 = ~new_n11968 & new_n11688;
  assign new_n11970 = new_n11969 ^ new_n11691;
  assign new_n11971 = new_n11970 ^ new_n11967;
  assign new_n11972 = new_n11695 ^ new_n11442;
  assign new_n11973 = ~new_n11972 & new_n11696;
  assign new_n11974 = new_n11973 ^ new_n11442;
  assign new_n11975 = new_n11974 ^ new_n11971;
  assign new_n11976 = ~new_n4212 & n97;
  assign new_n11977 = new_n3435 & new_n4201;
  assign new_n11978 = new_n11977 ^ new_n11976;
  assign new_n11979 = n98 & new_n4200;
  assign new_n11980 = n96 & new_n4206;
  assign new_n11981 = new_n11980 ^ new_n11979;
  assign new_n11982 = new_n11981 ^ new_n11978;
  assign new_n11983 = new_n11982 ^ n42;
  assign new_n11984 = ~new_n5424 & n91;
  assign new_n11985 = new_n2481 & new_n5419;
  assign new_n11986 = new_n11985 ^ new_n11984;
  assign new_n11987 = n92 & new_n5418;
  assign new_n11988 = n90 & new_n5648;
  assign new_n11989 = new_n11988 ^ new_n11987;
  assign new_n11990 = new_n11989 ^ new_n11986;
  assign new_n11991 = new_n11990 ^ n48;
  assign new_n11992 = ~new_n6110 & n88;
  assign new_n11993 = new_n2063 & new_n6105;
  assign new_n11994 = new_n11993 ^ new_n11992;
  assign new_n11995 = n89 & new_n6104;
  assign new_n11996 = n87 & new_n6347;
  assign new_n11997 = new_n11996 ^ new_n11995;
  assign new_n11998 = new_n11997 ^ new_n11994;
  assign new_n11999 = new_n11998 ^ n51;
  assign new_n12000 = n79 & new_n8355;
  assign new_n12001 = new_n1069 & new_n8345;
  assign new_n12002 = new_n12001 ^ new_n12000;
  assign new_n12003 = n80 & new_n8344;
  assign new_n12004 = n78 & new_n8349;
  assign new_n12005 = new_n12004 ^ new_n12003;
  assign new_n12006 = new_n12005 ^ new_n12002;
  assign new_n12007 = new_n12006 ^ n60;
  assign new_n12008 = new_n11797 ^ new_n11779;
  assign new_n12009 = new_n11780 & new_n12008;
  assign new_n12010 = new_n12009 ^ new_n11771;
  assign new_n12011 = new_n12010 ^ new_n12007;
  assign new_n12012 = ~new_n11783 & ~new_n11787;
  assign new_n12013 = ~new_n11793 & ~new_n12012;
  assign new_n12014 = n76 & new_n9195;
  assign new_n12015 = ~new_n812 & new_n9185;
  assign new_n12016 = new_n12015 ^ new_n12014;
  assign new_n12017 = n77 & new_n9184;
  assign new_n12018 = n75 & new_n9189;
  assign new_n12019 = new_n12018 ^ new_n12017;
  assign new_n12020 = new_n12019 ^ new_n12016;
  assign new_n12021 = new_n12020 ^ n63;
  assign new_n12022 = n74 ^ n72;
  assign new_n12023 = ~new_n11492 & new_n12022;
  assign new_n12024 = new_n12023 ^ n72;
  assign new_n12025 = new_n12024 ^ n73;
  assign new_n12026 = new_n11789 & new_n12025;
  assign new_n12027 = new_n12026 ^ n9;
  assign new_n12028 = new_n12027 ^ new_n12021;
  assign new_n12029 = new_n12028 ^ new_n12013;
  assign new_n12030 = new_n12029 ^ new_n12011;
  assign new_n12031 = n82 & new_n7553;
  assign new_n12032 = new_n1363 & new_n7543;
  assign new_n12033 = new_n12032 ^ new_n12031;
  assign new_n12034 = n83 & new_n7542;
  assign new_n12035 = n81 & new_n7547;
  assign new_n12036 = new_n12035 ^ new_n12034;
  assign new_n12037 = new_n12036 ^ new_n12033;
  assign new_n12038 = new_n12037 ^ n57;
  assign new_n12039 = new_n12038 ^ new_n12030;
  assign new_n12040 = new_n11810 ^ new_n11806;
  assign new_n12041 = ~new_n11807 & ~new_n12040;
  assign new_n12042 = new_n12041 ^ new_n11798;
  assign new_n12043 = new_n12042 ^ new_n12039;
  assign new_n12044 = ~new_n6805 & n85;
  assign new_n12045 = new_n1694 & new_n6800;
  assign new_n12046 = new_n12045 ^ new_n12044;
  assign new_n12047 = n86 & new_n6799;
  assign new_n12048 = n84 & new_n6811;
  assign new_n12049 = new_n12048 ^ new_n12047;
  assign new_n12050 = new_n12049 ^ new_n12046;
  assign new_n12051 = new_n12050 ^ n54;
  assign new_n12052 = new_n12051 ^ new_n12043;
  assign new_n12053 = new_n11815 ^ new_n11811;
  assign new_n12054 = ~new_n11812 & new_n12053;
  assign new_n12055 = new_n12054 ^ new_n11763;
  assign new_n12056 = new_n12055 ^ new_n12052;
  assign new_n12057 = new_n12056 ^ new_n11999;
  assign new_n12058 = new_n11820 ^ new_n11816;
  assign new_n12059 = ~new_n11817 & new_n12058;
  assign new_n12060 = new_n12059 ^ new_n11755;
  assign new_n12061 = new_n12060 ^ new_n12057;
  assign new_n12062 = new_n12061 ^ new_n11991;
  assign new_n12063 = new_n11821 ^ new_n11746;
  assign new_n12064 = new_n11747 & new_n12063;
  assign new_n12065 = new_n12064 ^ new_n11743;
  assign new_n12066 = new_n12065 ^ new_n12062;
  assign new_n12067 = new_n11826 ^ new_n11822;
  assign new_n12068 = ~new_n11823 & new_n12067;
  assign new_n12069 = new_n12068 ^ new_n11735;
  assign new_n12070 = new_n12069 ^ new_n12066;
  assign new_n12071 = ~new_n4804 & n94;
  assign new_n12072 = new_n2934 & new_n4799;
  assign new_n12073 = new_n12072 ^ new_n12071;
  assign new_n12074 = n95 & new_n4798;
  assign new_n12075 = n93 & new_n4810;
  assign new_n12076 = new_n12075 ^ new_n12074;
  assign new_n12077 = new_n12076 ^ new_n12073;
  assign new_n12078 = new_n12077 ^ n45;
  assign new_n12079 = new_n12078 ^ new_n12070;
  assign new_n12080 = new_n12079 ^ new_n11983;
  assign new_n12081 = new_n11831 ^ new_n11727;
  assign new_n12082 = new_n11828 & new_n12081;
  assign new_n12083 = new_n12082 ^ new_n11831;
  assign new_n12084 = new_n12083 ^ new_n12080;
  assign new_n12085 = ~new_n3682 & n100;
  assign new_n12086 = new_n3677 & new_n3972;
  assign new_n12087 = new_n12086 ^ new_n12085;
  assign new_n12088 = n101 & new_n3676;
  assign new_n12089 = n99 & new_n3688;
  assign new_n12090 = new_n12089 ^ new_n12088;
  assign new_n12091 = new_n12090 ^ new_n12087;
  assign new_n12092 = new_n12091 ^ n39;
  assign new_n12093 = new_n12092 ^ new_n12084;
  assign new_n12094 = new_n11844 ^ new_n11832;
  assign new_n12095 = ~new_n12094 & new_n11841;
  assign new_n12096 = new_n12095 ^ new_n11844;
  assign new_n12097 = new_n12096 ^ new_n12093;
  assign new_n12098 = ~new_n3143 & n103;
  assign new_n12099 = ~new_n4556 & new_n3138;
  assign new_n12100 = new_n12099 ^ new_n12098;
  assign new_n12101 = n104 & new_n3137;
  assign new_n12102 = n102 & new_n3149;
  assign new_n12103 = new_n12102 ^ new_n12101;
  assign new_n12104 = new_n12103 ^ new_n12100;
  assign new_n12105 = new_n12104 ^ n36;
  assign new_n12106 = new_n12105 ^ new_n12097;
  assign new_n12107 = new_n11857 ^ new_n11845;
  assign new_n12108 = ~new_n12107 & new_n11854;
  assign new_n12109 = new_n12108 ^ new_n11857;
  assign new_n12110 = new_n12109 ^ new_n12106;
  assign new_n12111 = ~new_n2672 & n106;
  assign new_n12112 = ~new_n5164 & new_n2667;
  assign new_n12113 = new_n12112 ^ new_n12111;
  assign new_n12114 = n107 & new_n2666;
  assign new_n12115 = n105 & new_n2664;
  assign new_n12116 = new_n12115 ^ new_n12114;
  assign new_n12117 = new_n12116 ^ new_n12113;
  assign new_n12118 = new_n12117 ^ n33;
  assign new_n12119 = new_n12118 ^ new_n12110;
  assign new_n12120 = new_n11870 ^ new_n11858;
  assign new_n12121 = new_n11867 & new_n12120;
  assign new_n12122 = new_n12121 ^ new_n11870;
  assign new_n12123 = new_n12122 ^ new_n12119;
  assign new_n12124 = n109 & new_n2246;
  assign new_n12125 = new_n2241 & new_n5825;
  assign new_n12126 = new_n12125 ^ new_n12124;
  assign new_n12127 = n110 & new_n2240;
  assign new_n12128 = n108 & new_n2391;
  assign new_n12129 = new_n12128 ^ new_n12127;
  assign new_n12130 = new_n12129 ^ new_n12126;
  assign new_n12131 = new_n12130 ^ n30;
  assign new_n12132 = new_n12131 ^ new_n12123;
  assign new_n12133 = new_n11883 ^ new_n11871;
  assign new_n12134 = ~new_n11880 & new_n12133;
  assign new_n12135 = new_n12134 ^ new_n11883;
  assign new_n12136 = new_n12135 ^ new_n12132;
  assign new_n12137 = n112 & new_n1874;
  assign new_n12138 = ~new_n6518 & new_n1864;
  assign new_n12139 = new_n12138 ^ new_n12137;
  assign new_n12140 = n113 & new_n1863;
  assign new_n12141 = n111 & new_n1868;
  assign new_n12142 = new_n12141 ^ new_n12140;
  assign new_n12143 = new_n12142 ^ new_n12139;
  assign new_n12144 = new_n12143 ^ n27;
  assign new_n12145 = new_n12144 ^ new_n12136;
  assign new_n12146 = new_n11896 ^ new_n11884;
  assign new_n12147 = ~new_n11893 & new_n12146;
  assign new_n12148 = new_n12147 ^ new_n11896;
  assign new_n12149 = new_n12148 ^ new_n12145;
  assign new_n12150 = ~new_n1506 & n115;
  assign new_n12151 = ~new_n7256 & new_n1501;
  assign new_n12152 = new_n12151 ^ new_n12150;
  assign new_n12153 = n116 & new_n1500;
  assign new_n12154 = n114 & new_n1512;
  assign new_n12155 = new_n12154 ^ new_n12153;
  assign new_n12156 = new_n12155 ^ new_n12152;
  assign new_n12157 = new_n12156 ^ n24;
  assign new_n12158 = new_n12157 ^ new_n12149;
  assign new_n12159 = new_n11909 ^ new_n11897;
  assign new_n12160 = ~new_n11906 & new_n12159;
  assign new_n12161 = new_n12160 ^ new_n11909;
  assign new_n12162 = new_n12161 ^ new_n12158;
  assign new_n12163 = ~new_n1198 & n118;
  assign new_n12164 = ~new_n8019 & new_n1193;
  assign new_n12165 = new_n12164 ^ new_n12163;
  assign new_n12166 = n119 & new_n1192;
  assign new_n12167 = n117 & new_n1204;
  assign new_n12168 = new_n12167 ^ new_n12166;
  assign new_n12169 = new_n12168 ^ new_n12165;
  assign new_n12170 = new_n12169 ^ n21;
  assign new_n12171 = new_n12170 ^ new_n12162;
  assign new_n12172 = new_n11922 ^ new_n11910;
  assign new_n12173 = ~new_n11919 & new_n12172;
  assign new_n12174 = new_n12173 ^ new_n11922;
  assign new_n12175 = new_n12174 ^ new_n12171;
  assign new_n12176 = ~new_n930 & n121;
  assign new_n12177 = new_n925 & new_n8850;
  assign new_n12178 = new_n12177 ^ new_n12176;
  assign new_n12179 = n122 & new_n924;
  assign new_n12180 = n120 & new_n936;
  assign new_n12181 = new_n12180 ^ new_n12179;
  assign new_n12182 = new_n12181 ^ new_n12178;
  assign new_n12183 = new_n12182 ^ n18;
  assign new_n12184 = new_n12183 ^ new_n12175;
  assign new_n12185 = new_n11935 ^ new_n11923;
  assign new_n12186 = ~new_n11932 & ~new_n12185;
  assign new_n12187 = new_n12186 ^ new_n11935;
  assign new_n12188 = new_n12187 ^ new_n12184;
  assign new_n12189 = n124 & new_n707;
  assign new_n12190 = new_n701 & new_n9700;
  assign new_n12191 = new_n12190 ^ new_n12189;
  assign new_n12192 = n125 & new_n700;
  assign new_n12193 = n123 & new_n787;
  assign new_n12194 = new_n12193 ^ new_n12192;
  assign new_n12195 = new_n12194 ^ new_n12191;
  assign new_n12196 = new_n12195 ^ n15;
  assign new_n12197 = new_n12196 ^ new_n12188;
  assign new_n12198 = new_n11948 ^ new_n11936;
  assign new_n12199 = ~new_n12198 & new_n11945;
  assign new_n12200 = new_n12199 ^ new_n11948;
  assign new_n12201 = new_n12200 ^ new_n12197;
  assign new_n12202 = n127 & new_n499;
  assign new_n12203 = ~new_n506 & new_n10581;
  assign new_n12204 = new_n12203 ^ new_n12202;
  assign new_n12205 = ~new_n505 & n128;
  assign new_n12206 = n126 & new_n579;
  assign new_n12207 = new_n12206 ^ new_n12205;
  assign new_n12208 = new_n12207 ^ new_n12204;
  assign new_n12209 = new_n12208 ^ n12;
  assign new_n12210 = new_n12209 ^ new_n12201;
  assign new_n12211 = new_n11961 ^ new_n11949;
  assign new_n12212 = new_n11958 & new_n12211;
  assign new_n12213 = new_n12212 ^ new_n11961;
  assign new_n12214 = new_n12213 ^ new_n12210;
  assign new_n12215 = ~new_n11719 & ~new_n11962;
  assign new_n12216 = new_n12215 ^ new_n11963;
  assign new_n12217 = ~new_n12216 & new_n11966;
  assign new_n12218 = new_n12217 ^ new_n11963;
  assign new_n12219 = new_n11966 ^ new_n11962;
  assign new_n12220 = ~new_n11963 & new_n12219;
  assign new_n12221 = new_n12220 ^ new_n12218;
  assign new_n12222 = new_n12221 ^ new_n12217;
  assign new_n12223 = new_n11974 ^ new_n11970;
  assign new_n12224 = new_n12220 ^ new_n11966;
  assign new_n12225 = new_n12224 ^ new_n11970;
  assign new_n12226 = new_n12225 ^ new_n12221;
  assign new_n12227 = new_n12226 ^ new_n12217;
  assign new_n12228 = new_n12223 & new_n12227;
  assign new_n12229 = new_n12228 ^ new_n12222;
  assign new_n12230 = new_n12229 ^ new_n12214;
  assign new_n12231 = ~new_n12217 & new_n12214;
  assign new_n12232 = ~new_n12231 & new_n12221;
  assign new_n12233 = new_n11970 & new_n12232;
  assign new_n12234 = new_n12232 ^ new_n11970;
  assign new_n12235 = new_n12234 ^ new_n12233;
  assign new_n12236 = ~new_n12214 & new_n12224;
  assign new_n12237 = new_n12224 ^ new_n12214;
  assign new_n12238 = new_n12237 ^ new_n12236;
  assign new_n12239 = ~new_n12238 & new_n12235;
  assign new_n12240 = ~new_n11974 & new_n12239;
  assign new_n12241 = ~new_n12233 & ~new_n12236;
  assign new_n12242 = ~new_n12240 & new_n12241;
  assign new_n12243 = ~new_n3682 & n101;
  assign new_n12244 = new_n3677 & new_n4159;
  assign new_n12245 = new_n12244 ^ new_n12243;
  assign new_n12246 = n102 & new_n3676;
  assign new_n12247 = n100 & new_n3688;
  assign new_n12248 = new_n12247 ^ new_n12246;
  assign new_n12249 = new_n12248 ^ new_n12245;
  assign new_n12250 = new_n12249 ^ n39;
  assign new_n12251 = ~new_n4212 & n98;
  assign new_n12252 = new_n3604 & new_n4201;
  assign new_n12253 = new_n12252 ^ new_n12251;
  assign new_n12254 = n99 & new_n4200;
  assign new_n12255 = n97 & new_n4206;
  assign new_n12256 = new_n12255 ^ new_n12254;
  assign new_n12257 = new_n12256 ^ new_n12253;
  assign new_n12258 = new_n12257 ^ n42;
  assign new_n12259 = ~new_n4804 & n95;
  assign new_n12260 = new_n3095 & new_n4799;
  assign new_n12261 = new_n12260 ^ new_n12259;
  assign new_n12262 = n96 & new_n4798;
  assign new_n12263 = n94 & new_n4810;
  assign new_n12264 = new_n12263 ^ new_n12262;
  assign new_n12265 = new_n12264 ^ new_n12261;
  assign new_n12266 = new_n12265 ^ n45;
  assign new_n12267 = ~new_n5424 & n92;
  assign new_n12268 = new_n2628 & new_n5419;
  assign new_n12269 = new_n12268 ^ new_n12267;
  assign new_n12270 = n93 & new_n5418;
  assign new_n12271 = n91 & new_n5648;
  assign new_n12272 = new_n12271 ^ new_n12270;
  assign new_n12273 = new_n12272 ^ new_n12269;
  assign new_n12274 = new_n12273 ^ n48;
  assign new_n12275 = ~new_n6110 & n89;
  assign new_n12276 = new_n2193 & new_n6105;
  assign new_n12277 = new_n12276 ^ new_n12275;
  assign new_n12278 = n90 & new_n6104;
  assign new_n12279 = n88 & new_n6347;
  assign new_n12280 = new_n12279 ^ new_n12278;
  assign new_n12281 = new_n12280 ^ new_n12277;
  assign new_n12282 = new_n12281 ^ n51;
  assign new_n12283 = ~new_n6805 & n86;
  assign new_n12284 = new_n1811 & new_n6800;
  assign new_n12285 = new_n12284 ^ new_n12283;
  assign new_n12286 = n87 & new_n6799;
  assign new_n12287 = n85 & new_n6811;
  assign new_n12288 = new_n12287 ^ new_n12286;
  assign new_n12289 = new_n12288 ^ new_n12285;
  assign new_n12290 = new_n12289 ^ n54;
  assign new_n12291 = new_n12042 ^ new_n12038;
  assign new_n12292 = ~new_n12039 & new_n12291;
  assign new_n12293 = new_n12292 ^ new_n12030;
  assign new_n12294 = new_n12293 ^ new_n12290;
  assign new_n12295 = n83 & new_n7553;
  assign new_n12296 = new_n1468 & new_n7543;
  assign new_n12297 = new_n12296 ^ new_n12295;
  assign new_n12298 = n84 & new_n7542;
  assign new_n12299 = n82 & new_n7547;
  assign new_n12300 = new_n12299 ^ new_n12298;
  assign new_n12301 = new_n12300 ^ new_n12297;
  assign new_n12302 = new_n12301 ^ n57;
  assign new_n12303 = n80 & new_n8355;
  assign new_n12304 = new_n1161 & new_n8345;
  assign new_n12305 = new_n12304 ^ new_n12303;
  assign new_n12306 = n81 & new_n8344;
  assign new_n12307 = n79 & new_n8349;
  assign new_n12308 = new_n12307 ^ new_n12306;
  assign new_n12309 = new_n12308 ^ new_n12305;
  assign new_n12310 = new_n12309 ^ n60;
  assign new_n12311 = n77 & new_n9195;
  assign new_n12312 = ~new_n891 & new_n9185;
  assign new_n12313 = new_n12312 ^ new_n12311;
  assign new_n12314 = n78 & new_n9184;
  assign new_n12315 = n76 & new_n9189;
  assign new_n12316 = new_n12315 ^ new_n12314;
  assign new_n12317 = new_n12316 ^ new_n12313;
  assign new_n12318 = new_n12317 ^ n63;
  assign new_n12319 = n74 & new_n11492;
  assign new_n12320 = n75 & new_n9495;
  assign new_n12321 = new_n12320 ^ new_n12319;
  assign new_n12322 = n73 ^ n9;
  assign new_n12323 = ~new_n12322 & new_n12025;
  assign new_n12324 = new_n12323 ^ n73;
  assign new_n12325 = new_n11789 & new_n12324;
  assign new_n12326 = new_n12325 ^ new_n12321;
  assign new_n12327 = new_n12326 ^ new_n12318;
  assign new_n12328 = new_n12327 ^ new_n12310;
  assign new_n12329 = new_n12021 ^ new_n12013;
  assign new_n12330 = new_n12028 & new_n12329;
  assign new_n12331 = new_n12330 ^ new_n12013;
  assign new_n12332 = new_n12331 ^ new_n12328;
  assign new_n12333 = new_n12332 ^ new_n12302;
  assign new_n12334 = new_n12029 ^ new_n12007;
  assign new_n12335 = new_n12011 & new_n12334;
  assign new_n12336 = new_n12335 ^ new_n12010;
  assign new_n12337 = new_n12336 ^ new_n12333;
  assign new_n12338 = new_n12337 ^ new_n12294;
  assign new_n12339 = new_n12338 ^ new_n12282;
  assign new_n12340 = new_n12055 ^ new_n12043;
  assign new_n12341 = ~new_n12052 & new_n12340;
  assign new_n12342 = new_n12341 ^ new_n12055;
  assign new_n12343 = new_n12342 ^ new_n12339;
  assign new_n12344 = new_n12343 ^ new_n12274;
  assign new_n12345 = new_n12060 ^ new_n11999;
  assign new_n12346 = ~new_n12057 & new_n12345;
  assign new_n12347 = new_n12346 ^ new_n12060;
  assign new_n12348 = new_n12347 ^ new_n12344;
  assign new_n12349 = new_n12348 ^ new_n12266;
  assign new_n12350 = new_n12065 ^ new_n11991;
  assign new_n12351 = ~new_n12062 & new_n12350;
  assign new_n12352 = new_n12351 ^ new_n12065;
  assign new_n12353 = new_n12352 ^ new_n12349;
  assign new_n12354 = new_n12353 ^ new_n12258;
  assign new_n12355 = new_n12078 ^ new_n12066;
  assign new_n12356 = ~new_n12355 & new_n12070;
  assign new_n12357 = new_n12356 ^ new_n12069;
  assign new_n12358 = new_n12357 ^ new_n12354;
  assign new_n12359 = new_n12358 ^ new_n12250;
  assign new_n12360 = new_n12083 ^ new_n11983;
  assign new_n12361 = ~new_n12080 & new_n12360;
  assign new_n12362 = new_n12361 ^ new_n12083;
  assign new_n12363 = new_n12362 ^ new_n12359;
  assign new_n12364 = ~new_n3143 & n104;
  assign new_n12365 = ~new_n4754 & new_n3138;
  assign new_n12366 = new_n12365 ^ new_n12364;
  assign new_n12367 = n105 & new_n3137;
  assign new_n12368 = n103 & new_n3149;
  assign new_n12369 = new_n12368 ^ new_n12367;
  assign new_n12370 = new_n12369 ^ new_n12366;
  assign new_n12371 = new_n12370 ^ n36;
  assign new_n12372 = new_n12371 ^ new_n12363;
  assign new_n12373 = new_n12096 ^ new_n12084;
  assign new_n12374 = ~new_n12093 & new_n12373;
  assign new_n12375 = new_n12374 ^ new_n12096;
  assign new_n12376 = new_n12375 ^ new_n12372;
  assign new_n12377 = ~new_n2672 & n107;
  assign new_n12378 = ~new_n5377 & new_n2667;
  assign new_n12379 = new_n12378 ^ new_n12377;
  assign new_n12380 = n108 & new_n2666;
  assign new_n12381 = n106 & new_n2664;
  assign new_n12382 = new_n12381 ^ new_n12380;
  assign new_n12383 = new_n12382 ^ new_n12379;
  assign new_n12384 = new_n12383 ^ n33;
  assign new_n12385 = new_n12384 ^ new_n12376;
  assign new_n12386 = new_n12109 ^ new_n12097;
  assign new_n12387 = ~new_n12106 & new_n12386;
  assign new_n12388 = new_n12387 ^ new_n12109;
  assign new_n12389 = new_n12388 ^ new_n12385;
  assign new_n12390 = n110 & new_n2246;
  assign new_n12391 = new_n2241 & new_n6049;
  assign new_n12392 = new_n12391 ^ new_n12390;
  assign new_n12393 = n111 & new_n2240;
  assign new_n12394 = n109 & new_n2391;
  assign new_n12395 = new_n12394 ^ new_n12393;
  assign new_n12396 = new_n12395 ^ new_n12392;
  assign new_n12397 = new_n12396 ^ n30;
  assign new_n12398 = new_n12397 ^ new_n12389;
  assign new_n12399 = new_n12122 ^ new_n12110;
  assign new_n12400 = ~new_n12119 & ~new_n12399;
  assign new_n12401 = new_n12400 ^ new_n12122;
  assign new_n12402 = new_n12401 ^ new_n12398;
  assign new_n12403 = n113 & new_n1874;
  assign new_n12404 = ~new_n6764 & new_n1864;
  assign new_n12405 = new_n12404 ^ new_n12403;
  assign new_n12406 = n114 & new_n1863;
  assign new_n12407 = n112 & new_n1868;
  assign new_n12408 = new_n12407 ^ new_n12406;
  assign new_n12409 = new_n12408 ^ new_n12405;
  assign new_n12410 = new_n12409 ^ n27;
  assign new_n12411 = new_n12410 ^ new_n12402;
  assign new_n12412 = new_n12135 ^ new_n12123;
  assign new_n12413 = ~new_n12412 & new_n12132;
  assign new_n12414 = new_n12413 ^ new_n12135;
  assign new_n12415 = new_n12414 ^ new_n12411;
  assign new_n12416 = ~new_n1506 & n116;
  assign new_n12417 = ~new_n7503 & new_n1501;
  assign new_n12418 = new_n12417 ^ new_n12416;
  assign new_n12419 = n117 & new_n1500;
  assign new_n12420 = n115 & new_n1512;
  assign new_n12421 = new_n12420 ^ new_n12419;
  assign new_n12422 = new_n12421 ^ new_n12418;
  assign new_n12423 = new_n12422 ^ n24;
  assign new_n12424 = new_n12423 ^ new_n12415;
  assign new_n12425 = new_n12148 ^ new_n12136;
  assign new_n12426 = ~new_n12425 & new_n12145;
  assign new_n12427 = new_n12426 ^ new_n12148;
  assign new_n12428 = new_n12427 ^ new_n12424;
  assign new_n12429 = ~new_n1198 & n119;
  assign new_n12430 = new_n1193 & new_n8286;
  assign new_n12431 = new_n12430 ^ new_n12429;
  assign new_n12432 = n120 & new_n1192;
  assign new_n12433 = n118 & new_n1204;
  assign new_n12434 = new_n12433 ^ new_n12432;
  assign new_n12435 = new_n12434 ^ new_n12431;
  assign new_n12436 = new_n12435 ^ n21;
  assign new_n12437 = new_n12436 ^ new_n12428;
  assign new_n12438 = new_n12161 ^ new_n12149;
  assign new_n12439 = ~new_n12438 & new_n12158;
  assign new_n12440 = new_n12439 ^ new_n12161;
  assign new_n12441 = new_n12440 ^ new_n12437;
  assign new_n12442 = ~new_n930 & n122;
  assign new_n12443 = ~new_n9116 & new_n925;
  assign new_n12444 = new_n12443 ^ new_n12442;
  assign new_n12445 = n123 & new_n924;
  assign new_n12446 = n121 & new_n936;
  assign new_n12447 = new_n12446 ^ new_n12445;
  assign new_n12448 = new_n12447 ^ new_n12444;
  assign new_n12449 = new_n12448 ^ n18;
  assign new_n12450 = new_n12449 ^ new_n12441;
  assign new_n12451 = new_n12174 ^ new_n12162;
  assign new_n12452 = ~new_n12451 & new_n12171;
  assign new_n12453 = new_n12452 ^ new_n12174;
  assign new_n12454 = new_n12453 ^ new_n12450;
  assign new_n12455 = n125 & new_n707;
  assign new_n12456 = new_n701 & new_n9987;
  assign new_n12457 = new_n12456 ^ new_n12455;
  assign new_n12458 = n126 & new_n700;
  assign new_n12459 = n124 & new_n787;
  assign new_n12460 = new_n12459 ^ new_n12458;
  assign new_n12461 = new_n12460 ^ new_n12457;
  assign new_n12462 = new_n12461 ^ n15;
  assign new_n12463 = new_n12462 ^ new_n12454;
  assign new_n12464 = new_n12187 ^ new_n12175;
  assign new_n12465 = new_n12184 & new_n12464;
  assign new_n12466 = new_n12465 ^ new_n12187;
  assign new_n12467 = new_n12466 ^ new_n12463;
  assign new_n12468 = n127 & new_n579;
  assign new_n12469 = ~new_n506 & new_n10010;
  assign new_n12470 = new_n12469 ^ new_n12468;
  assign new_n12471 = n128 & new_n499;
  assign new_n12472 = new_n12471 ^ new_n12470;
  assign new_n12473 = new_n12472 ^ n12;
  assign new_n12474 = new_n12473 ^ new_n12467;
  assign new_n12475 = new_n12200 ^ new_n12188;
  assign new_n12476 = ~new_n12197 & new_n12475;
  assign new_n12477 = new_n12476 ^ new_n12200;
  assign new_n12478 = new_n12477 ^ new_n12474;
  assign new_n12479 = new_n12213 ^ new_n12209;
  assign new_n12480 = new_n12210 & new_n12479;
  assign new_n12481 = new_n12480 ^ new_n12201;
  assign new_n12482 = new_n12481 ^ new_n12478;
  assign new_n12483 = new_n12482 ^ new_n12242;
  assign new_n12484 = new_n443 ^ n12;
  assign new_n12485 = new_n444 ^ new_n443;
  assign new_n12486 = new_n503 ^ new_n444;
  assign new_n12487 = new_n444 & new_n12486;
  assign new_n12488 = new_n12487 ^ new_n444;
  assign new_n12489 = ~new_n12485 & new_n12488;
  assign new_n12490 = new_n12489 ^ new_n12487;
  assign new_n12491 = new_n12490 ^ new_n444;
  assign new_n12492 = new_n12491 ^ new_n503;
  assign new_n12493 = ~new_n12484 & new_n12492;
  assign new_n12494 = new_n12493 ^ n12;
  assign new_n12495 = new_n12494 ^ n12;
  assign new_n12496 = new_n12484 & new_n12492;
  assign new_n12497 = new_n12496 ^ n11;
  assign new_n12498 = new_n12497 ^ n12;
  assign new_n12499 = new_n12498 ^ new_n12495;
  assign new_n12500 = new_n12498 ^ new_n10009;
  assign new_n12501 = new_n12500 ^ new_n12498;
  assign new_n12502 = new_n12499 & new_n12501;
  assign new_n12503 = new_n12502 ^ new_n12498;
  assign new_n12504 = n128 & new_n12503;
  assign new_n12505 = new_n12504 ^ n12;
  assign new_n12506 = ~new_n3143 & n105;
  assign new_n12507 = ~new_n4961 & new_n3138;
  assign new_n12508 = new_n12507 ^ new_n12506;
  assign new_n12509 = n106 & new_n3137;
  assign new_n12510 = n104 & new_n3149;
  assign new_n12511 = new_n12510 ^ new_n12509;
  assign new_n12512 = new_n12511 ^ new_n12508;
  assign new_n12513 = new_n12512 ^ n36;
  assign new_n12514 = ~new_n3682 & n102;
  assign new_n12515 = new_n3677 & new_n4368;
  assign new_n12516 = new_n12515 ^ new_n12514;
  assign new_n12517 = n103 & new_n3676;
  assign new_n12518 = n101 & new_n3688;
  assign new_n12519 = new_n12518 ^ new_n12517;
  assign new_n12520 = new_n12519 ^ new_n12516;
  assign new_n12521 = new_n12520 ^ n39;
  assign new_n12522 = ~new_n4212 & n99;
  assign new_n12523 = new_n3789 & new_n4201;
  assign new_n12524 = new_n12523 ^ new_n12522;
  assign new_n12525 = n100 & new_n4200;
  assign new_n12526 = n98 & new_n4206;
  assign new_n12527 = new_n12526 ^ new_n12525;
  assign new_n12528 = new_n12527 ^ new_n12524;
  assign new_n12529 = new_n12528 ^ n42;
  assign new_n12530 = ~new_n4804 & n96;
  assign new_n12531 = new_n3273 & new_n4799;
  assign new_n12532 = new_n12531 ^ new_n12530;
  assign new_n12533 = n97 & new_n4798;
  assign new_n12534 = n95 & new_n4810;
  assign new_n12535 = new_n12534 ^ new_n12533;
  assign new_n12536 = new_n12535 ^ new_n12532;
  assign new_n12537 = new_n12536 ^ n45;
  assign new_n12538 = ~new_n5424 & n93;
  assign new_n12539 = new_n2785 & new_n5419;
  assign new_n12540 = new_n12539 ^ new_n12538;
  assign new_n12541 = n94 & new_n5418;
  assign new_n12542 = n92 & new_n5648;
  assign new_n12543 = new_n12542 ^ new_n12541;
  assign new_n12544 = new_n12543 ^ new_n12540;
  assign new_n12545 = new_n12544 ^ n48;
  assign new_n12546 = ~new_n6110 & n90;
  assign new_n12547 = new_n2341 & new_n6105;
  assign new_n12548 = new_n12547 ^ new_n12546;
  assign new_n12549 = n91 & new_n6104;
  assign new_n12550 = n89 & new_n6347;
  assign new_n12551 = new_n12550 ^ new_n12549;
  assign new_n12552 = new_n12551 ^ new_n12548;
  assign new_n12553 = new_n12552 ^ n51;
  assign new_n12554 = new_n12337 ^ new_n12290;
  assign new_n12555 = ~new_n12294 & new_n12554;
  assign new_n12556 = new_n12555 ^ new_n12293;
  assign new_n12557 = new_n12556 ^ new_n12553;
  assign new_n12558 = ~new_n6805 & n87;
  assign new_n12559 = new_n1940 & new_n6800;
  assign new_n12560 = new_n12559 ^ new_n12558;
  assign new_n12561 = n88 & new_n6799;
  assign new_n12562 = n86 & new_n6811;
  assign new_n12563 = new_n12562 ^ new_n12561;
  assign new_n12564 = new_n12563 ^ new_n12560;
  assign new_n12565 = new_n12564 ^ n54;
  assign new_n12566 = n84 & new_n7553;
  assign new_n12567 = new_n1584 & new_n7543;
  assign new_n12568 = new_n12567 ^ new_n12566;
  assign new_n12569 = n85 & new_n7542;
  assign new_n12570 = n83 & new_n7547;
  assign new_n12571 = new_n12570 ^ new_n12569;
  assign new_n12572 = new_n12571 ^ new_n12568;
  assign new_n12573 = new_n12572 ^ n57;
  assign new_n12574 = n75 ^ n74;
  assign new_n12575 = ~n75 & n76;
  assign new_n12576 = new_n12575 ^ new_n12574;
  assign new_n12577 = new_n12576 ^ new_n12575;
  assign new_n12578 = n64 & new_n12577;
  assign new_n12579 = new_n12578 ^ new_n12575;
  assign new_n12580 = ~new_n9495 & new_n12579;
  assign new_n12581 = new_n12580 ^ new_n12575;
  assign new_n12582 = ~n76 & new_n12320;
  assign new_n12583 = new_n12582 ^ new_n12581;
  assign new_n12584 = new_n12325 ^ new_n12318;
  assign new_n12585 = new_n12326 & new_n12584;
  assign new_n12586 = new_n12585 ^ new_n12318;
  assign new_n12587 = new_n12586 ^ new_n12583;
  assign new_n12588 = n78 & new_n9195;
  assign new_n12589 = ~new_n982 & new_n9185;
  assign new_n12590 = new_n12589 ^ new_n12588;
  assign new_n12591 = n79 & new_n9184;
  assign new_n12592 = n77 & new_n9189;
  assign new_n12593 = new_n12592 ^ new_n12591;
  assign new_n12594 = new_n12593 ^ new_n12590;
  assign new_n12595 = new_n12594 ^ n63;
  assign new_n12596 = new_n12595 ^ new_n12587;
  assign new_n12597 = n81 & new_n8355;
  assign new_n12598 = new_n1263 & new_n8345;
  assign new_n12599 = new_n12598 ^ new_n12597;
  assign new_n12600 = n82 & new_n8344;
  assign new_n12601 = n80 & new_n8349;
  assign new_n12602 = new_n12601 ^ new_n12600;
  assign new_n12603 = new_n12602 ^ new_n12599;
  assign new_n12604 = new_n12603 ^ n60;
  assign new_n12605 = new_n12604 ^ new_n12596;
  assign new_n12606 = new_n12605 ^ new_n12573;
  assign new_n12607 = new_n12331 ^ new_n12310;
  assign new_n12608 = new_n12328 & new_n12607;
  assign new_n12609 = new_n12608 ^ new_n12331;
  assign new_n12610 = new_n12609 ^ new_n12606;
  assign new_n12611 = new_n12610 ^ new_n12565;
  assign new_n12612 = new_n12336 ^ new_n12302;
  assign new_n12613 = new_n12333 & new_n12612;
  assign new_n12614 = new_n12613 ^ new_n12336;
  assign new_n12615 = new_n12614 ^ new_n12611;
  assign new_n12616 = new_n12615 ^ new_n12557;
  assign new_n12617 = new_n12616 ^ new_n12545;
  assign new_n12618 = new_n12342 ^ new_n12338;
  assign new_n12619 = ~new_n12618 & new_n12339;
  assign new_n12620 = new_n12619 ^ new_n12282;
  assign new_n12621 = new_n12620 ^ new_n12617;
  assign new_n12622 = new_n12621 ^ new_n12537;
  assign new_n12623 = new_n12347 ^ new_n12343;
  assign new_n12624 = ~new_n12623 & new_n12344;
  assign new_n12625 = new_n12624 ^ new_n12274;
  assign new_n12626 = new_n12625 ^ new_n12622;
  assign new_n12627 = new_n12352 ^ new_n12348;
  assign new_n12628 = ~new_n12627 & new_n12349;
  assign new_n12629 = new_n12628 ^ new_n12266;
  assign new_n12630 = new_n12629 ^ new_n12626;
  assign new_n12631 = new_n12630 ^ new_n12529;
  assign new_n12632 = new_n12357 ^ new_n12353;
  assign new_n12633 = ~new_n12632 & new_n12354;
  assign new_n12634 = new_n12633 ^ new_n12258;
  assign new_n12635 = new_n12634 ^ new_n12631;
  assign new_n12636 = new_n12635 ^ new_n12521;
  assign new_n12637 = new_n12636 ^ new_n12513;
  assign new_n12638 = new_n12362 ^ new_n12250;
  assign new_n12639 = ~new_n12359 & new_n12638;
  assign new_n12640 = new_n12639 ^ new_n12362;
  assign new_n12641 = new_n12640 ^ new_n12637;
  assign new_n12642 = ~new_n2672 & n108;
  assign new_n12643 = new_n2667 & new_n5604;
  assign new_n12644 = new_n12643 ^ new_n12642;
  assign new_n12645 = n109 & new_n2666;
  assign new_n12646 = n107 & new_n2664;
  assign new_n12647 = new_n12646 ^ new_n12645;
  assign new_n12648 = new_n12647 ^ new_n12644;
  assign new_n12649 = new_n12648 ^ n33;
  assign new_n12650 = new_n12649 ^ new_n12641;
  assign new_n12651 = new_n12375 ^ new_n12363;
  assign new_n12652 = ~new_n12372 & new_n12651;
  assign new_n12653 = new_n12652 ^ new_n12375;
  assign new_n12654 = new_n12653 ^ new_n12650;
  assign new_n12655 = n111 & new_n2246;
  assign new_n12656 = ~new_n6284 & new_n2241;
  assign new_n12657 = new_n12656 ^ new_n12655;
  assign new_n12658 = n112 & new_n2240;
  assign new_n12659 = n110 & new_n2391;
  assign new_n12660 = new_n12659 ^ new_n12658;
  assign new_n12661 = new_n12660 ^ new_n12657;
  assign new_n12662 = new_n12661 ^ n30;
  assign new_n12663 = new_n12662 ^ new_n12654;
  assign new_n12664 = new_n12388 ^ new_n12376;
  assign new_n12665 = ~new_n12385 & new_n12664;
  assign new_n12666 = new_n12665 ^ new_n12388;
  assign new_n12667 = new_n12666 ^ new_n12663;
  assign new_n12668 = n114 & new_n1874;
  assign new_n12669 = ~new_n7013 & new_n1864;
  assign new_n12670 = new_n12669 ^ new_n12668;
  assign new_n12671 = n115 & new_n1863;
  assign new_n12672 = n113 & new_n1868;
  assign new_n12673 = new_n12672 ^ new_n12671;
  assign new_n12674 = new_n12673 ^ new_n12670;
  assign new_n12675 = new_n12674 ^ n27;
  assign new_n12676 = new_n12675 ^ new_n12667;
  assign new_n12677 = new_n12401 ^ new_n12389;
  assign new_n12678 = ~new_n12398 & ~new_n12677;
  assign new_n12679 = new_n12678 ^ new_n12401;
  assign new_n12680 = new_n12679 ^ new_n12676;
  assign new_n12681 = ~new_n1506 & n117;
  assign new_n12682 = ~new_n7761 & new_n1501;
  assign new_n12683 = new_n12682 ^ new_n12681;
  assign new_n12684 = n118 & new_n1500;
  assign new_n12685 = n116 & new_n1512;
  assign new_n12686 = new_n12685 ^ new_n12684;
  assign new_n12687 = new_n12686 ^ new_n12683;
  assign new_n12688 = new_n12687 ^ n24;
  assign new_n12689 = new_n12688 ^ new_n12680;
  assign new_n12690 = new_n12414 ^ new_n12402;
  assign new_n12691 = ~new_n12690 & new_n12411;
  assign new_n12692 = new_n12691 ^ new_n12414;
  assign new_n12693 = new_n12692 ^ new_n12689;
  assign new_n12694 = ~new_n1198 & n120;
  assign new_n12695 = new_n1193 & new_n8560;
  assign new_n12696 = new_n12695 ^ new_n12694;
  assign new_n12697 = n121 & new_n1192;
  assign new_n12698 = n119 & new_n1204;
  assign new_n12699 = new_n12698 ^ new_n12697;
  assign new_n12700 = new_n12699 ^ new_n12696;
  assign new_n12701 = new_n12700 ^ n21;
  assign new_n12702 = new_n12701 ^ new_n12693;
  assign new_n12703 = new_n12427 ^ new_n12415;
  assign new_n12704 = ~new_n12703 & new_n12424;
  assign new_n12705 = new_n12704 ^ new_n12427;
  assign new_n12706 = new_n12705 ^ new_n12702;
  assign new_n12707 = ~new_n930 & n123;
  assign new_n12708 = ~new_n9405 & new_n925;
  assign new_n12709 = new_n12708 ^ new_n12707;
  assign new_n12710 = n124 & new_n924;
  assign new_n12711 = n122 & new_n936;
  assign new_n12712 = new_n12711 ^ new_n12710;
  assign new_n12713 = new_n12712 ^ new_n12709;
  assign new_n12714 = new_n12713 ^ n18;
  assign new_n12715 = new_n12714 ^ new_n12706;
  assign new_n12716 = new_n12440 ^ new_n12428;
  assign new_n12717 = ~new_n12716 & new_n12437;
  assign new_n12718 = new_n12717 ^ new_n12440;
  assign new_n12719 = new_n12718 ^ new_n12715;
  assign new_n12720 = n126 & new_n707;
  assign new_n12721 = new_n701 & new_n10304;
  assign new_n12722 = new_n12721 ^ new_n12720;
  assign new_n12723 = n127 & new_n700;
  assign new_n12724 = n125 & new_n787;
  assign new_n12725 = new_n12724 ^ new_n12723;
  assign new_n12726 = new_n12725 ^ new_n12722;
  assign new_n12727 = new_n12726 ^ n15;
  assign new_n12728 = new_n12727 ^ new_n12719;
  assign new_n12729 = new_n12453 ^ new_n12441;
  assign new_n12730 = ~new_n12729 & new_n12450;
  assign new_n12731 = new_n12730 ^ new_n12453;
  assign new_n12732 = new_n12731 ^ new_n12728;
  assign new_n12733 = new_n12732 ^ new_n12505;
  assign new_n12734 = new_n12466 ^ new_n12454;
  assign new_n12735 = new_n12463 & new_n12734;
  assign new_n12736 = new_n12735 ^ new_n12466;
  assign new_n12737 = new_n12736 ^ new_n12733;
  assign new_n12738 = new_n12477 ^ new_n12467;
  assign new_n12739 = ~new_n12474 & new_n12738;
  assign new_n12740 = new_n12739 ^ new_n12477;
  assign new_n12741 = new_n12740 ^ new_n12737;
  assign new_n12742 = new_n12481 ^ new_n12242;
  assign new_n12743 = ~new_n12482 & ~new_n12742;
  assign new_n12744 = new_n12743 ^ new_n12242;
  assign new_n12745 = new_n12744 ^ new_n12741;
  assign new_n12746 = ~new_n3143 & n106;
  assign new_n12747 = ~new_n5164 & new_n3138;
  assign new_n12748 = new_n12747 ^ new_n12746;
  assign new_n12749 = n107 & new_n3137;
  assign new_n12750 = n105 & new_n3149;
  assign new_n12751 = new_n12750 ^ new_n12749;
  assign new_n12752 = new_n12751 ^ new_n12748;
  assign new_n12753 = new_n12752 ^ n36;
  assign new_n12754 = ~new_n4212 & n100;
  assign new_n12755 = new_n3972 & new_n4201;
  assign new_n12756 = new_n12755 ^ new_n12754;
  assign new_n12757 = n101 & new_n4200;
  assign new_n12758 = n99 & new_n4206;
  assign new_n12759 = new_n12758 ^ new_n12757;
  assign new_n12760 = new_n12759 ^ new_n12756;
  assign new_n12761 = new_n12760 ^ n42;
  assign new_n12762 = ~new_n4804 & n97;
  assign new_n12763 = new_n3435 & new_n4799;
  assign new_n12764 = new_n12763 ^ new_n12762;
  assign new_n12765 = n98 & new_n4798;
  assign new_n12766 = n96 & new_n4810;
  assign new_n12767 = new_n12766 ^ new_n12765;
  assign new_n12768 = new_n12767 ^ new_n12764;
  assign new_n12769 = new_n12768 ^ n45;
  assign new_n12770 = ~new_n5424 & n94;
  assign new_n12771 = new_n2934 & new_n5419;
  assign new_n12772 = new_n12771 ^ new_n12770;
  assign new_n12773 = n95 & new_n5418;
  assign new_n12774 = n93 & new_n5648;
  assign new_n12775 = new_n12774 ^ new_n12773;
  assign new_n12776 = new_n12775 ^ new_n12772;
  assign new_n12777 = new_n12776 ^ n48;
  assign new_n12778 = new_n12620 ^ new_n12616;
  assign new_n12779 = ~new_n12778 & new_n12617;
  assign new_n12780 = new_n12779 ^ new_n12545;
  assign new_n12781 = new_n12780 ^ new_n12777;
  assign new_n12782 = ~new_n6110 & n91;
  assign new_n12783 = new_n2481 & new_n6105;
  assign new_n12784 = new_n12783 ^ new_n12782;
  assign new_n12785 = n92 & new_n6104;
  assign new_n12786 = n90 & new_n6347;
  assign new_n12787 = new_n12786 ^ new_n12785;
  assign new_n12788 = new_n12787 ^ new_n12784;
  assign new_n12789 = new_n12788 ^ n51;
  assign new_n12790 = ~new_n6805 & n88;
  assign new_n12791 = new_n2063 & new_n6800;
  assign new_n12792 = new_n12791 ^ new_n12790;
  assign new_n12793 = n89 & new_n6799;
  assign new_n12794 = n87 & new_n6811;
  assign new_n12795 = new_n12794 ^ new_n12793;
  assign new_n12796 = new_n12795 ^ new_n12792;
  assign new_n12797 = new_n12796 ^ n54;
  assign new_n12798 = ~new_n12581 & ~new_n12586;
  assign new_n12799 = ~n75 & new_n12319;
  assign new_n12800 = new_n12799 ^ new_n12582;
  assign new_n12801 = ~new_n12798 & ~new_n12800;
  assign new_n12802 = n79 & new_n9195;
  assign new_n12803 = new_n1069 & new_n9185;
  assign new_n12804 = new_n12803 ^ new_n12802;
  assign new_n12805 = n80 & new_n9184;
  assign new_n12806 = n78 & new_n9189;
  assign new_n12807 = new_n12806 ^ new_n12805;
  assign new_n12808 = new_n12807 ^ new_n12804;
  assign new_n12809 = new_n12808 ^ n63;
  assign new_n12810 = n64 & n76;
  assign new_n12811 = new_n12810 ^ n77;
  assign new_n12812 = ~new_n9495 & new_n12811;
  assign new_n12813 = new_n12812 ^ n77;
  assign new_n12814 = new_n12813 ^ new_n12321;
  assign new_n12815 = new_n12814 ^ n12;
  assign new_n12816 = new_n12815 ^ new_n12809;
  assign new_n12817 = new_n12816 ^ new_n12801;
  assign new_n12818 = n82 & new_n8355;
  assign new_n12819 = new_n1363 & new_n8345;
  assign new_n12820 = new_n12819 ^ new_n12818;
  assign new_n12821 = n83 & new_n8344;
  assign new_n12822 = n81 & new_n8349;
  assign new_n12823 = new_n12822 ^ new_n12821;
  assign new_n12824 = new_n12823 ^ new_n12820;
  assign new_n12825 = new_n12824 ^ n60;
  assign new_n12826 = new_n12825 ^ new_n12817;
  assign new_n12827 = new_n12604 ^ new_n12595;
  assign new_n12828 = ~new_n12596 & ~new_n12827;
  assign new_n12829 = new_n12828 ^ new_n12587;
  assign new_n12830 = new_n12829 ^ new_n12826;
  assign new_n12831 = n85 & new_n7553;
  assign new_n12832 = new_n1694 & new_n7543;
  assign new_n12833 = new_n12832 ^ new_n12831;
  assign new_n12834 = n86 & new_n7542;
  assign new_n12835 = n84 & new_n7547;
  assign new_n12836 = new_n12835 ^ new_n12834;
  assign new_n12837 = new_n12836 ^ new_n12833;
  assign new_n12838 = new_n12837 ^ n57;
  assign new_n12839 = new_n12838 ^ new_n12830;
  assign new_n12840 = new_n12609 ^ new_n12605;
  assign new_n12841 = ~new_n12606 & new_n12840;
  assign new_n12842 = new_n12841 ^ new_n12573;
  assign new_n12843 = new_n12842 ^ new_n12839;
  assign new_n12844 = new_n12843 ^ new_n12797;
  assign new_n12845 = new_n12614 ^ new_n12610;
  assign new_n12846 = ~new_n12611 & new_n12845;
  assign new_n12847 = new_n12846 ^ new_n12565;
  assign new_n12848 = new_n12847 ^ new_n12844;
  assign new_n12849 = new_n12848 ^ new_n12789;
  assign new_n12850 = new_n12615 ^ new_n12556;
  assign new_n12851 = ~new_n12557 & ~new_n12850;
  assign new_n12852 = new_n12851 ^ new_n12553;
  assign new_n12853 = new_n12852 ^ new_n12849;
  assign new_n12854 = new_n12853 ^ new_n12781;
  assign new_n12855 = new_n12854 ^ new_n12769;
  assign new_n12856 = new_n12625 ^ new_n12621;
  assign new_n12857 = ~new_n12856 & new_n12622;
  assign new_n12858 = new_n12857 ^ new_n12537;
  assign new_n12859 = new_n12858 ^ new_n12855;
  assign new_n12860 = new_n12859 ^ new_n12761;
  assign new_n12861 = new_n12626 ^ new_n12529;
  assign new_n12862 = ~new_n12630 & new_n12861;
  assign new_n12863 = new_n12862 ^ new_n12529;
  assign new_n12864 = new_n12863 ^ new_n12860;
  assign new_n12865 = new_n12634 ^ new_n12521;
  assign new_n12866 = ~new_n12635 & new_n12865;
  assign new_n12867 = new_n12866 ^ new_n12521;
  assign new_n12868 = new_n12867 ^ new_n12864;
  assign new_n12869 = ~new_n3682 & n103;
  assign new_n12870 = ~new_n4556 & new_n3677;
  assign new_n12871 = new_n12870 ^ new_n12869;
  assign new_n12872 = n104 & new_n3676;
  assign new_n12873 = n102 & new_n3688;
  assign new_n12874 = new_n12873 ^ new_n12872;
  assign new_n12875 = new_n12874 ^ new_n12871;
  assign new_n12876 = new_n12875 ^ n39;
  assign new_n12877 = new_n12876 ^ new_n12868;
  assign new_n12878 = new_n12877 ^ new_n12753;
  assign new_n12879 = new_n12640 ^ new_n12513;
  assign new_n12880 = ~new_n12637 & new_n12879;
  assign new_n12881 = new_n12880 ^ new_n12640;
  assign new_n12882 = new_n12881 ^ new_n12878;
  assign new_n12883 = ~new_n2672 & n109;
  assign new_n12884 = new_n2667 & new_n5825;
  assign new_n12885 = new_n12884 ^ new_n12883;
  assign new_n12886 = n110 & new_n2666;
  assign new_n12887 = n108 & new_n2664;
  assign new_n12888 = new_n12887 ^ new_n12886;
  assign new_n12889 = new_n12888 ^ new_n12885;
  assign new_n12890 = new_n12889 ^ n33;
  assign new_n12891 = new_n12890 ^ new_n12882;
  assign new_n12892 = new_n12653 ^ new_n12641;
  assign new_n12893 = ~new_n12650 & new_n12892;
  assign new_n12894 = new_n12893 ^ new_n12653;
  assign new_n12895 = new_n12894 ^ new_n12891;
  assign new_n12896 = n112 & new_n2246;
  assign new_n12897 = ~new_n6518 & new_n2241;
  assign new_n12898 = new_n12897 ^ new_n12896;
  assign new_n12899 = n113 & new_n2240;
  assign new_n12900 = n111 & new_n2391;
  assign new_n12901 = new_n12900 ^ new_n12899;
  assign new_n12902 = new_n12901 ^ new_n12898;
  assign new_n12903 = new_n12902 ^ n30;
  assign new_n12904 = new_n12903 ^ new_n12895;
  assign new_n12905 = new_n12666 ^ new_n12654;
  assign new_n12906 = ~new_n12663 & new_n12905;
  assign new_n12907 = new_n12906 ^ new_n12666;
  assign new_n12908 = new_n12907 ^ new_n12904;
  assign new_n12909 = n115 & new_n1874;
  assign new_n12910 = ~new_n7256 & new_n1864;
  assign new_n12911 = new_n12910 ^ new_n12909;
  assign new_n12912 = n116 & new_n1863;
  assign new_n12913 = n114 & new_n1868;
  assign new_n12914 = new_n12913 ^ new_n12912;
  assign new_n12915 = new_n12914 ^ new_n12911;
  assign new_n12916 = new_n12915 ^ n27;
  assign new_n12917 = new_n12916 ^ new_n12908;
  assign new_n12918 = new_n12679 ^ new_n12667;
  assign new_n12919 = ~new_n12676 & ~new_n12918;
  assign new_n12920 = new_n12919 ^ new_n12679;
  assign new_n12921 = new_n12920 ^ new_n12917;
  assign new_n12922 = ~new_n1506 & n118;
  assign new_n12923 = ~new_n8019 & new_n1501;
  assign new_n12924 = new_n12923 ^ new_n12922;
  assign new_n12925 = n119 & new_n1500;
  assign new_n12926 = n117 & new_n1512;
  assign new_n12927 = new_n12926 ^ new_n12925;
  assign new_n12928 = new_n12927 ^ new_n12924;
  assign new_n12929 = new_n12928 ^ n24;
  assign new_n12930 = new_n12929 ^ new_n12921;
  assign new_n12931 = new_n12692 ^ new_n12680;
  assign new_n12932 = ~new_n12931 & new_n12689;
  assign new_n12933 = new_n12932 ^ new_n12692;
  assign new_n12934 = new_n12933 ^ new_n12930;
  assign new_n12935 = ~new_n1198 & n121;
  assign new_n12936 = new_n1193 & new_n8850;
  assign new_n12937 = new_n12936 ^ new_n12935;
  assign new_n12938 = n122 & new_n1192;
  assign new_n12939 = n120 & new_n1204;
  assign new_n12940 = new_n12939 ^ new_n12938;
  assign new_n12941 = new_n12940 ^ new_n12937;
  assign new_n12942 = new_n12941 ^ n21;
  assign new_n12943 = new_n12942 ^ new_n12934;
  assign new_n12944 = new_n12705 ^ new_n12693;
  assign new_n12945 = ~new_n12944 & new_n12702;
  assign new_n12946 = new_n12945 ^ new_n12705;
  assign new_n12947 = new_n12946 ^ new_n12943;
  assign new_n12948 = ~new_n930 & n124;
  assign new_n12949 = new_n925 & new_n9700;
  assign new_n12950 = new_n12949 ^ new_n12948;
  assign new_n12951 = n125 & new_n924;
  assign new_n12952 = n123 & new_n936;
  assign new_n12953 = new_n12952 ^ new_n12951;
  assign new_n12954 = new_n12953 ^ new_n12950;
  assign new_n12955 = new_n12954 ^ n18;
  assign new_n12956 = new_n12955 ^ new_n12947;
  assign new_n12957 = new_n12718 ^ new_n12706;
  assign new_n12958 = ~new_n12957 & new_n12715;
  assign new_n12959 = new_n12958 ^ new_n12718;
  assign new_n12960 = new_n12959 ^ new_n12956;
  assign new_n12961 = n127 & new_n707;
  assign new_n12962 = new_n701 & new_n10581;
  assign new_n12963 = new_n12962 ^ new_n12961;
  assign new_n12964 = n128 & new_n700;
  assign new_n12965 = n126 & new_n787;
  assign new_n12966 = new_n12965 ^ new_n12964;
  assign new_n12967 = new_n12966 ^ new_n12963;
  assign new_n12968 = new_n12967 ^ n15;
  assign new_n12969 = new_n12968 ^ new_n12960;
  assign new_n12970 = new_n12731 ^ new_n12719;
  assign new_n12971 = ~new_n12970 & new_n12728;
  assign new_n12972 = new_n12971 ^ new_n12731;
  assign new_n12973 = new_n12972 ^ new_n12969;
  assign new_n12974 = new_n12736 ^ new_n12732;
  assign new_n12975 = new_n12733 & new_n12974;
  assign new_n12976 = new_n12975 ^ new_n12736;
  assign new_n12977 = new_n12976 ^ new_n12973;
  assign new_n12978 = new_n12744 ^ new_n12740;
  assign new_n12979 = ~new_n12741 & ~new_n12978;
  assign new_n12980 = new_n12979 ^ new_n12744;
  assign new_n12981 = new_n12980 ^ new_n12977;
  assign new_n12982 = ~new_n2672 & n110;
  assign new_n12983 = new_n2667 & new_n6049;
  assign new_n12984 = new_n12983 ^ new_n12982;
  assign new_n12985 = n111 & new_n2666;
  assign new_n12986 = n109 & new_n2664;
  assign new_n12987 = new_n12986 ^ new_n12985;
  assign new_n12988 = new_n12987 ^ new_n12984;
  assign new_n12989 = new_n12988 ^ n33;
  assign new_n12990 = ~new_n3143 & n107;
  assign new_n12991 = ~new_n5377 & new_n3138;
  assign new_n12992 = new_n12991 ^ new_n12990;
  assign new_n12993 = n108 & new_n3137;
  assign new_n12994 = n106 & new_n3149;
  assign new_n12995 = new_n12994 ^ new_n12993;
  assign new_n12996 = new_n12995 ^ new_n12992;
  assign new_n12997 = new_n12996 ^ n36;
  assign new_n12998 = ~new_n3682 & n104;
  assign new_n12999 = ~new_n4754 & new_n3677;
  assign new_n13000 = new_n12999 ^ new_n12998;
  assign new_n13001 = n105 & new_n3676;
  assign new_n13002 = n103 & new_n3688;
  assign new_n13003 = new_n13002 ^ new_n13001;
  assign new_n13004 = new_n13003 ^ new_n13000;
  assign new_n13005 = new_n13004 ^ n39;
  assign new_n13006 = ~new_n4212 & n101;
  assign new_n13007 = new_n4159 & new_n4201;
  assign new_n13008 = new_n13007 ^ new_n13006;
  assign new_n13009 = n102 & new_n4200;
  assign new_n13010 = n100 & new_n4206;
  assign new_n13011 = new_n13010 ^ new_n13009;
  assign new_n13012 = new_n13011 ^ new_n13008;
  assign new_n13013 = new_n13012 ^ n42;
  assign new_n13014 = ~new_n4804 & n98;
  assign new_n13015 = new_n3604 & new_n4799;
  assign new_n13016 = new_n13015 ^ new_n13014;
  assign new_n13017 = n99 & new_n4798;
  assign new_n13018 = n97 & new_n4810;
  assign new_n13019 = new_n13018 ^ new_n13017;
  assign new_n13020 = new_n13019 ^ new_n13016;
  assign new_n13021 = new_n13020 ^ n45;
  assign new_n13022 = ~new_n5424 & n95;
  assign new_n13023 = new_n3095 & new_n5419;
  assign new_n13024 = new_n13023 ^ new_n13022;
  assign new_n13025 = n96 & new_n5418;
  assign new_n13026 = n94 & new_n5648;
  assign new_n13027 = new_n13026 ^ new_n13025;
  assign new_n13028 = new_n13027 ^ new_n13024;
  assign new_n13029 = new_n13028 ^ n48;
  assign new_n13030 = ~new_n6110 & n92;
  assign new_n13031 = new_n2628 & new_n6105;
  assign new_n13032 = new_n13031 ^ new_n13030;
  assign new_n13033 = n93 & new_n6104;
  assign new_n13034 = n91 & new_n6347;
  assign new_n13035 = new_n13034 ^ new_n13033;
  assign new_n13036 = new_n13035 ^ new_n13032;
  assign new_n13037 = new_n13036 ^ n51;
  assign new_n13038 = ~new_n6805 & n89;
  assign new_n13039 = new_n2193 & new_n6800;
  assign new_n13040 = new_n13039 ^ new_n13038;
  assign new_n13041 = n90 & new_n6799;
  assign new_n13042 = n88 & new_n6811;
  assign new_n13043 = new_n13042 ^ new_n13041;
  assign new_n13044 = new_n13043 ^ new_n13040;
  assign new_n13045 = new_n13044 ^ n54;
  assign new_n13046 = n86 & new_n7553;
  assign new_n13047 = new_n1811 & new_n7543;
  assign new_n13048 = new_n13047 ^ new_n13046;
  assign new_n13049 = n87 & new_n7542;
  assign new_n13050 = n85 & new_n7547;
  assign new_n13051 = new_n13050 ^ new_n13049;
  assign new_n13052 = new_n13051 ^ new_n13048;
  assign new_n13053 = new_n13052 ^ n57;
  assign new_n13054 = new_n12829 ^ new_n12817;
  assign new_n13055 = new_n12826 & new_n13054;
  assign new_n13056 = new_n13055 ^ new_n12829;
  assign new_n13057 = new_n13056 ^ new_n13053;
  assign new_n13058 = n83 & new_n8355;
  assign new_n13059 = new_n1468 & new_n8345;
  assign new_n13060 = new_n13059 ^ new_n13058;
  assign new_n13061 = n84 & new_n8344;
  assign new_n13062 = n82 & new_n8349;
  assign new_n13063 = new_n13062 ^ new_n13061;
  assign new_n13064 = new_n13063 ^ new_n13060;
  assign new_n13065 = new_n13064 ^ n60;
  assign new_n13066 = n80 & new_n9195;
  assign new_n13067 = new_n1161 & new_n9185;
  assign new_n13068 = new_n13067 ^ new_n13066;
  assign new_n13069 = n81 & new_n9184;
  assign new_n13070 = n79 & new_n9189;
  assign new_n13071 = new_n13070 ^ new_n13069;
  assign new_n13072 = new_n13071 ^ new_n13068;
  assign new_n13073 = new_n13072 ^ n63;
  assign new_n13074 = n64 & n77;
  assign new_n13075 = new_n13074 ^ n78;
  assign new_n13076 = ~new_n9495 & new_n13075;
  assign new_n13077 = new_n13076 ^ n78;
  assign new_n13078 = new_n12321 ^ n12;
  assign new_n13079 = ~new_n12814 & ~new_n13078;
  assign new_n13080 = new_n13079 ^ n12;
  assign new_n13081 = new_n13080 ^ new_n13077;
  assign new_n13082 = new_n13081 ^ new_n13073;
  assign new_n13083 = new_n13082 ^ new_n13065;
  assign new_n13084 = new_n12809 ^ new_n12801;
  assign new_n13085 = new_n12816 & new_n13084;
  assign new_n13086 = new_n13085 ^ new_n12801;
  assign new_n13087 = new_n13086 ^ new_n13083;
  assign new_n13088 = new_n13087 ^ new_n13057;
  assign new_n13089 = new_n13088 ^ new_n13045;
  assign new_n13090 = new_n12842 ^ new_n12830;
  assign new_n13091 = ~new_n12839 & new_n13090;
  assign new_n13092 = new_n13091 ^ new_n12842;
  assign new_n13093 = new_n13092 ^ new_n13089;
  assign new_n13094 = new_n13093 ^ new_n13037;
  assign new_n13095 = new_n12847 ^ new_n12797;
  assign new_n13096 = ~new_n12844 & new_n13095;
  assign new_n13097 = new_n13096 ^ new_n12847;
  assign new_n13098 = new_n13097 ^ new_n13094;
  assign new_n13099 = new_n13098 ^ new_n13029;
  assign new_n13100 = new_n12852 ^ new_n12789;
  assign new_n13101 = ~new_n12849 & new_n13100;
  assign new_n13102 = new_n13101 ^ new_n12852;
  assign new_n13103 = new_n13102 ^ new_n13099;
  assign new_n13104 = new_n13103 ^ new_n13021;
  assign new_n13105 = new_n12853 ^ new_n12777;
  assign new_n13106 = ~new_n13105 & new_n12781;
  assign new_n13107 = new_n13106 ^ new_n12780;
  assign new_n13108 = new_n13107 ^ new_n13104;
  assign new_n13109 = new_n12858 ^ new_n12769;
  assign new_n13110 = ~new_n12855 & new_n13109;
  assign new_n13111 = new_n13110 ^ new_n12858;
  assign new_n13112 = new_n13111 ^ new_n13108;
  assign new_n13113 = new_n13112 ^ new_n13013;
  assign new_n13114 = new_n12863 ^ new_n12761;
  assign new_n13115 = ~new_n12860 & new_n13114;
  assign new_n13116 = new_n13115 ^ new_n12863;
  assign new_n13117 = new_n13116 ^ new_n13113;
  assign new_n13118 = new_n13117 ^ new_n13005;
  assign new_n13119 = new_n12876 ^ new_n12864;
  assign new_n13120 = ~new_n13119 & new_n12868;
  assign new_n13121 = new_n13120 ^ new_n12867;
  assign new_n13122 = new_n13121 ^ new_n13118;
  assign new_n13123 = new_n13122 ^ new_n12997;
  assign new_n13124 = new_n13123 ^ new_n12989;
  assign new_n13125 = new_n12881 ^ new_n12753;
  assign new_n13126 = ~new_n12878 & new_n13125;
  assign new_n13127 = new_n13126 ^ new_n12881;
  assign new_n13128 = new_n13127 ^ new_n13124;
  assign new_n13129 = new_n12894 ^ new_n12882;
  assign new_n13130 = ~new_n12891 & new_n13129;
  assign new_n13131 = new_n13130 ^ new_n12894;
  assign new_n13132 = new_n13131 ^ new_n13128;
  assign new_n13133 = n113 & new_n2246;
  assign new_n13134 = ~new_n6764 & new_n2241;
  assign new_n13135 = new_n13134 ^ new_n13133;
  assign new_n13136 = n114 & new_n2240;
  assign new_n13137 = n112 & new_n2391;
  assign new_n13138 = new_n13137 ^ new_n13136;
  assign new_n13139 = new_n13138 ^ new_n13135;
  assign new_n13140 = new_n13139 ^ n30;
  assign new_n13141 = new_n13140 ^ new_n13132;
  assign new_n13142 = n116 & new_n1874;
  assign new_n13143 = ~new_n7503 & new_n1864;
  assign new_n13144 = new_n13143 ^ new_n13142;
  assign new_n13145 = n117 & new_n1863;
  assign new_n13146 = n115 & new_n1868;
  assign new_n13147 = new_n13146 ^ new_n13145;
  assign new_n13148 = new_n13147 ^ new_n13144;
  assign new_n13149 = new_n13148 ^ n27;
  assign new_n13150 = new_n13149 ^ new_n13141;
  assign new_n13151 = new_n12907 ^ new_n12895;
  assign new_n13152 = ~new_n12904 & new_n13151;
  assign new_n13153 = new_n13152 ^ new_n12907;
  assign new_n13154 = new_n13153 ^ new_n13150;
  assign new_n13155 = ~new_n1506 & n119;
  assign new_n13156 = new_n1501 & new_n8286;
  assign new_n13157 = new_n13156 ^ new_n13155;
  assign new_n13158 = n120 & new_n1500;
  assign new_n13159 = n118 & new_n1512;
  assign new_n13160 = new_n13159 ^ new_n13158;
  assign new_n13161 = new_n13160 ^ new_n13157;
  assign new_n13162 = new_n13161 ^ n24;
  assign new_n13163 = new_n13162 ^ new_n13154;
  assign new_n13164 = new_n12920 ^ new_n12908;
  assign new_n13165 = ~new_n12917 & ~new_n13164;
  assign new_n13166 = new_n13165 ^ new_n12920;
  assign new_n13167 = new_n13166 ^ new_n13163;
  assign new_n13168 = ~new_n1198 & n122;
  assign new_n13169 = ~new_n9116 & new_n1193;
  assign new_n13170 = new_n13169 ^ new_n13168;
  assign new_n13171 = n123 & new_n1192;
  assign new_n13172 = n121 & new_n1204;
  assign new_n13173 = new_n13172 ^ new_n13171;
  assign new_n13174 = new_n13173 ^ new_n13170;
  assign new_n13175 = new_n13174 ^ n21;
  assign new_n13176 = new_n13175 ^ new_n13167;
  assign new_n13177 = new_n12933 ^ new_n12921;
  assign new_n13178 = ~new_n13177 & new_n12930;
  assign new_n13179 = new_n13178 ^ new_n12933;
  assign new_n13180 = new_n13179 ^ new_n13176;
  assign new_n13181 = ~new_n930 & n125;
  assign new_n13182 = new_n925 & new_n9987;
  assign new_n13183 = new_n13182 ^ new_n13181;
  assign new_n13184 = n126 & new_n924;
  assign new_n13185 = n124 & new_n936;
  assign new_n13186 = new_n13185 ^ new_n13184;
  assign new_n13187 = new_n13186 ^ new_n13183;
  assign new_n13188 = new_n13187 ^ n18;
  assign new_n13189 = new_n13188 ^ new_n13180;
  assign new_n13190 = new_n12946 ^ new_n12934;
  assign new_n13191 = ~new_n13190 & new_n12943;
  assign new_n13192 = new_n13191 ^ new_n12946;
  assign new_n13193 = new_n13192 ^ new_n13189;
  assign new_n13194 = n127 & new_n787;
  assign new_n13195 = new_n701 & new_n10010;
  assign new_n13196 = new_n13195 ^ new_n13194;
  assign new_n13197 = n128 & new_n707;
  assign new_n13198 = new_n13197 ^ new_n13196;
  assign new_n13199 = new_n13198 ^ n15;
  assign new_n13200 = new_n13199 ^ new_n13193;
  assign new_n13201 = new_n12959 ^ new_n12947;
  assign new_n13202 = ~new_n13201 & new_n12956;
  assign new_n13203 = new_n13202 ^ new_n12959;
  assign new_n13204 = new_n13203 ^ new_n13200;
  assign new_n13205 = new_n12972 ^ new_n12960;
  assign new_n13206 = ~new_n13205 & new_n12969;
  assign new_n13207 = new_n13206 ^ new_n12972;
  assign new_n13208 = new_n13207 ^ new_n13204;
  assign new_n13209 = new_n12980 ^ new_n12976;
  assign new_n13210 = ~new_n12977 & new_n13209;
  assign new_n13211 = new_n13210 ^ new_n12980;
  assign new_n13212 = new_n13211 ^ new_n13208;
  assign new_n13213 = ~new_n2672 & n111;
  assign new_n13214 = ~new_n6284 & new_n2667;
  assign new_n13215 = new_n13214 ^ new_n13213;
  assign new_n13216 = n112 & new_n2666;
  assign new_n13217 = n110 & new_n2664;
  assign new_n13218 = new_n13217 ^ new_n13216;
  assign new_n13219 = new_n13218 ^ new_n13215;
  assign new_n13220 = new_n13219 ^ n33;
  assign new_n13221 = ~new_n3143 & n108;
  assign new_n13222 = new_n3138 & new_n5604;
  assign new_n13223 = new_n13222 ^ new_n13221;
  assign new_n13224 = n109 & new_n3137;
  assign new_n13225 = n107 & new_n3149;
  assign new_n13226 = new_n13225 ^ new_n13224;
  assign new_n13227 = new_n13226 ^ new_n13223;
  assign new_n13228 = new_n13227 ^ n36;
  assign new_n13229 = ~new_n3682 & n105;
  assign new_n13230 = ~new_n4961 & new_n3677;
  assign new_n13231 = new_n13230 ^ new_n13229;
  assign new_n13232 = n106 & new_n3676;
  assign new_n13233 = n104 & new_n3688;
  assign new_n13234 = new_n13233 ^ new_n13232;
  assign new_n13235 = new_n13234 ^ new_n13231;
  assign new_n13236 = new_n13235 ^ n39;
  assign new_n13237 = ~new_n4212 & n102;
  assign new_n13238 = new_n4201 & new_n4368;
  assign new_n13239 = new_n13238 ^ new_n13237;
  assign new_n13240 = n103 & new_n4200;
  assign new_n13241 = n101 & new_n4206;
  assign new_n13242 = new_n13241 ^ new_n13240;
  assign new_n13243 = new_n13242 ^ new_n13239;
  assign new_n13244 = new_n13243 ^ n42;
  assign new_n13245 = ~new_n4804 & n99;
  assign new_n13246 = new_n3789 & new_n4799;
  assign new_n13247 = new_n13246 ^ new_n13245;
  assign new_n13248 = n100 & new_n4798;
  assign new_n13249 = n98 & new_n4810;
  assign new_n13250 = new_n13249 ^ new_n13248;
  assign new_n13251 = new_n13250 ^ new_n13247;
  assign new_n13252 = new_n13251 ^ n45;
  assign new_n13253 = ~new_n5424 & n96;
  assign new_n13254 = new_n3273 & new_n5419;
  assign new_n13255 = new_n13254 ^ new_n13253;
  assign new_n13256 = n97 & new_n5418;
  assign new_n13257 = n95 & new_n5648;
  assign new_n13258 = new_n13257 ^ new_n13256;
  assign new_n13259 = new_n13258 ^ new_n13255;
  assign new_n13260 = new_n13259 ^ n48;
  assign new_n13261 = ~new_n6110 & n93;
  assign new_n13262 = new_n2785 & new_n6105;
  assign new_n13263 = new_n13262 ^ new_n13261;
  assign new_n13264 = n94 & new_n6104;
  assign new_n13265 = n92 & new_n6347;
  assign new_n13266 = new_n13265 ^ new_n13264;
  assign new_n13267 = new_n13266 ^ new_n13263;
  assign new_n13268 = new_n13267 ^ n51;
  assign new_n13269 = ~new_n6805 & n90;
  assign new_n13270 = new_n2341 & new_n6800;
  assign new_n13271 = new_n13270 ^ new_n13269;
  assign new_n13272 = n91 & new_n6799;
  assign new_n13273 = n89 & new_n6811;
  assign new_n13274 = new_n13273 ^ new_n13272;
  assign new_n13275 = new_n13274 ^ new_n13271;
  assign new_n13276 = new_n13275 ^ n54;
  assign new_n13277 = new_n13087 ^ new_n13053;
  assign new_n13278 = ~new_n13057 & ~new_n13277;
  assign new_n13279 = new_n13278 ^ new_n13056;
  assign new_n13280 = new_n13279 ^ new_n13276;
  assign new_n13281 = n87 & new_n7553;
  assign new_n13282 = new_n1940 & new_n7543;
  assign new_n13283 = new_n13282 ^ new_n13281;
  assign new_n13284 = n88 & new_n7542;
  assign new_n13285 = n86 & new_n7547;
  assign new_n13286 = new_n13285 ^ new_n13284;
  assign new_n13287 = new_n13286 ^ new_n13283;
  assign new_n13288 = new_n13287 ^ n57;
  assign new_n13289 = n84 & new_n8355;
  assign new_n13290 = new_n1584 & new_n8345;
  assign new_n13291 = new_n13290 ^ new_n13289;
  assign new_n13292 = n85 & new_n8344;
  assign new_n13293 = n83 & new_n8349;
  assign new_n13294 = new_n13293 ^ new_n13292;
  assign new_n13295 = new_n13294 ^ new_n13291;
  assign new_n13296 = new_n13295 ^ n60;
  assign new_n13297 = n81 & new_n9195;
  assign new_n13298 = new_n1263 & new_n9185;
  assign new_n13299 = new_n13298 ^ new_n13297;
  assign new_n13300 = n82 & new_n9184;
  assign new_n13301 = n80 & new_n9189;
  assign new_n13302 = new_n13301 ^ new_n13300;
  assign new_n13303 = new_n13302 ^ new_n13299;
  assign new_n13304 = new_n825 ^ n63;
  assign new_n13305 = n64 & n79;
  assign new_n13306 = new_n13305 ^ new_n13075;
  assign new_n13307 = n64 & new_n825;
  assign new_n13308 = new_n13307 ^ n79;
  assign new_n13309 = new_n13308 ^ new_n13306;
  assign new_n13310 = ~new_n9495 & new_n13309;
  assign new_n13311 = new_n13310 ^ new_n13304;
  assign new_n13312 = new_n13311 ^ new_n13303;
  assign new_n13313 = new_n13080 ^ new_n13073;
  assign new_n13314 = ~new_n13081 & ~new_n13313;
  assign new_n13315 = new_n13314 ^ new_n13073;
  assign new_n13316 = new_n13315 ^ new_n13312;
  assign new_n13317 = new_n13316 ^ new_n13296;
  assign new_n13318 = new_n13317 ^ new_n13288;
  assign new_n13319 = new_n13086 ^ new_n13065;
  assign new_n13320 = ~new_n13083 & new_n13319;
  assign new_n13321 = new_n13320 ^ new_n13086;
  assign new_n13322 = new_n13321 ^ new_n13318;
  assign new_n13323 = new_n13322 ^ new_n13280;
  assign new_n13324 = new_n13323 ^ new_n13268;
  assign new_n13325 = new_n13092 ^ new_n13088;
  assign new_n13326 = ~new_n13089 & new_n13325;
  assign new_n13327 = new_n13326 ^ new_n13045;
  assign new_n13328 = new_n13327 ^ new_n13324;
  assign new_n13329 = new_n13328 ^ new_n13260;
  assign new_n13330 = new_n13097 ^ new_n13093;
  assign new_n13331 = ~new_n13094 & new_n13330;
  assign new_n13332 = new_n13331 ^ new_n13037;
  assign new_n13333 = new_n13332 ^ new_n13329;
  assign new_n13334 = new_n13333 ^ new_n13252;
  assign new_n13335 = new_n13102 ^ new_n13098;
  assign new_n13336 = ~new_n13099 & new_n13335;
  assign new_n13337 = new_n13336 ^ new_n13029;
  assign new_n13338 = new_n13337 ^ new_n13334;
  assign new_n13339 = new_n13107 ^ new_n13103;
  assign new_n13340 = ~new_n13104 & new_n13339;
  assign new_n13341 = new_n13340 ^ new_n13021;
  assign new_n13342 = new_n13341 ^ new_n13338;
  assign new_n13343 = new_n13342 ^ new_n13244;
  assign new_n13344 = new_n13111 ^ new_n13013;
  assign new_n13345 = new_n13112 & new_n13344;
  assign new_n13346 = new_n13345 ^ new_n13013;
  assign new_n13347 = new_n13346 ^ new_n13343;
  assign new_n13348 = new_n13347 ^ new_n13236;
  assign new_n13349 = new_n13116 ^ new_n13005;
  assign new_n13350 = new_n13117 & new_n13349;
  assign new_n13351 = new_n13350 ^ new_n13005;
  assign new_n13352 = new_n13351 ^ new_n13348;
  assign new_n13353 = new_n13352 ^ new_n13228;
  assign new_n13354 = new_n13121 ^ new_n12997;
  assign new_n13355 = new_n13122 & new_n13354;
  assign new_n13356 = new_n13355 ^ new_n12997;
  assign new_n13357 = new_n13356 ^ new_n13353;
  assign new_n13358 = new_n13357 ^ new_n13220;
  assign new_n13359 = new_n13127 ^ new_n12989;
  assign new_n13360 = new_n13124 & new_n13359;
  assign new_n13361 = new_n13360 ^ new_n13127;
  assign new_n13362 = new_n13361 ^ new_n13358;
  assign new_n13363 = n114 & new_n2246;
  assign new_n13364 = ~new_n7013 & new_n2241;
  assign new_n13365 = new_n13364 ^ new_n13363;
  assign new_n13366 = n115 & new_n2240;
  assign new_n13367 = n113 & new_n2391;
  assign new_n13368 = new_n13367 ^ new_n13366;
  assign new_n13369 = new_n13368 ^ new_n13365;
  assign new_n13370 = new_n13369 ^ n30;
  assign new_n13371 = new_n13370 ^ new_n13362;
  assign new_n13372 = new_n13140 ^ new_n13128;
  assign new_n13373 = ~new_n13132 & new_n13372;
  assign new_n13374 = new_n13373 ^ new_n13131;
  assign new_n13375 = new_n13374 ^ new_n13371;
  assign new_n13376 = n117 & new_n1874;
  assign new_n13377 = ~new_n7761 & new_n1864;
  assign new_n13378 = new_n13377 ^ new_n13376;
  assign new_n13379 = n118 & new_n1863;
  assign new_n13380 = n116 & new_n1868;
  assign new_n13381 = new_n13380 ^ new_n13379;
  assign new_n13382 = new_n13381 ^ new_n13378;
  assign new_n13383 = new_n13382 ^ n27;
  assign new_n13384 = new_n13383 ^ new_n13375;
  assign new_n13385 = ~new_n1506 & n120;
  assign new_n13386 = new_n1501 & new_n8560;
  assign new_n13387 = new_n13386 ^ new_n13385;
  assign new_n13388 = n121 & new_n1500;
  assign new_n13389 = n119 & new_n1512;
  assign new_n13390 = new_n13389 ^ new_n13388;
  assign new_n13391 = new_n13390 ^ new_n13387;
  assign new_n13392 = new_n13391 ^ n24;
  assign new_n13393 = new_n13392 ^ new_n13384;
  assign new_n13394 = new_n13153 ^ new_n13141;
  assign new_n13395 = ~new_n13394 & new_n13150;
  assign new_n13396 = new_n13395 ^ new_n13153;
  assign new_n13397 = new_n13396 ^ new_n13393;
  assign new_n13398 = new_n13166 ^ new_n13154;
  assign new_n13399 = new_n13163 & new_n13398;
  assign new_n13400 = new_n13399 ^ new_n13166;
  assign new_n13401 = new_n13400 ^ new_n13397;
  assign new_n13402 = ~new_n1198 & n123;
  assign new_n13403 = ~new_n9405 & new_n1193;
  assign new_n13404 = new_n13403 ^ new_n13402;
  assign new_n13405 = n124 & new_n1192;
  assign new_n13406 = n122 & new_n1204;
  assign new_n13407 = new_n13406 ^ new_n13405;
  assign new_n13408 = new_n13407 ^ new_n13404;
  assign new_n13409 = new_n13408 ^ n21;
  assign new_n13410 = new_n13409 ^ new_n13401;
  assign new_n13411 = new_n13179 ^ new_n13167;
  assign new_n13412 = ~new_n13176 & new_n13411;
  assign new_n13413 = new_n13412 ^ new_n13179;
  assign new_n13414 = new_n13413 ^ new_n13410;
  assign new_n13415 = ~new_n930 & n126;
  assign new_n13416 = new_n925 & new_n10304;
  assign new_n13417 = new_n13416 ^ new_n13415;
  assign new_n13418 = n127 & new_n924;
  assign new_n13419 = n125 & new_n936;
  assign new_n13420 = new_n13419 ^ new_n13418;
  assign new_n13421 = new_n13420 ^ new_n13417;
  assign new_n13422 = new_n13421 ^ n18;
  assign new_n13423 = new_n13422 ^ new_n13414;
  assign new_n13424 = n128 & new_n786;
  assign new_n13425 = ~n15 & ~new_n13424;
  assign new_n13426 = new_n13425 ^ n14;
  assign new_n13427 = new_n584 & new_n11133;
  assign new_n13428 = new_n13427 ^ new_n13424;
  assign new_n13429 = ~new_n13426 & ~new_n13428;
  assign new_n13430 = new_n13429 ^ n14;
  assign new_n13431 = new_n13430 ^ new_n13423;
  assign new_n13432 = new_n13192 ^ new_n13180;
  assign new_n13433 = ~new_n13189 & new_n13432;
  assign new_n13434 = new_n13433 ^ new_n13192;
  assign new_n13435 = new_n13434 ^ new_n13431;
  assign new_n13436 = new_n13203 ^ new_n13193;
  assign new_n13437 = ~new_n13200 & new_n13436;
  assign new_n13438 = new_n13437 ^ new_n13203;
  assign new_n13439 = new_n13438 ^ new_n13435;
  assign new_n13440 = new_n13211 ^ new_n13207;
  assign new_n13441 = ~new_n13208 & ~new_n13440;
  assign new_n13442 = new_n13441 ^ new_n13211;
  assign new_n13443 = new_n13442 ^ new_n13439;
  assign new_n13444 = new_n13442 ^ new_n13434;
  assign new_n13445 = new_n13444 ^ new_n13438;
  assign new_n13446 = ~new_n13439 & new_n13445;
  assign new_n13447 = new_n13434 & new_n13438;
  assign new_n13448 = ~new_n13430 & new_n13423;
  assign new_n13449 = new_n13448 ^ new_n13447;
  assign new_n13450 = new_n13449 ^ new_n13446;
  assign new_n13451 = n118 & new_n1874;
  assign new_n13452 = ~new_n8019 & new_n1864;
  assign new_n13453 = new_n13452 ^ new_n13451;
  assign new_n13454 = n119 & new_n1863;
  assign new_n13455 = n117 & new_n1868;
  assign new_n13456 = new_n13455 ^ new_n13454;
  assign new_n13457 = new_n13456 ^ new_n13453;
  assign new_n13458 = new_n13457 ^ n27;
  assign new_n13459 = n115 & new_n2246;
  assign new_n13460 = ~new_n7256 & new_n2241;
  assign new_n13461 = new_n13460 ^ new_n13459;
  assign new_n13462 = n116 & new_n2240;
  assign new_n13463 = n114 & new_n2391;
  assign new_n13464 = new_n13463 ^ new_n13462;
  assign new_n13465 = new_n13464 ^ new_n13461;
  assign new_n13466 = new_n13465 ^ n30;
  assign new_n13467 = ~new_n2672 & n112;
  assign new_n13468 = ~new_n6518 & new_n2667;
  assign new_n13469 = new_n13468 ^ new_n13467;
  assign new_n13470 = n113 & new_n2666;
  assign new_n13471 = n111 & new_n2664;
  assign new_n13472 = new_n13471 ^ new_n13470;
  assign new_n13473 = new_n13472 ^ new_n13469;
  assign new_n13474 = new_n13473 ^ n33;
  assign new_n13475 = ~new_n3143 & n109;
  assign new_n13476 = new_n3138 & new_n5825;
  assign new_n13477 = new_n13476 ^ new_n13475;
  assign new_n13478 = n110 & new_n3137;
  assign new_n13479 = n108 & new_n3149;
  assign new_n13480 = new_n13479 ^ new_n13478;
  assign new_n13481 = new_n13480 ^ new_n13477;
  assign new_n13482 = new_n13481 ^ n36;
  assign new_n13483 = ~new_n3682 & n106;
  assign new_n13484 = ~new_n5164 & new_n3677;
  assign new_n13485 = new_n13484 ^ new_n13483;
  assign new_n13486 = n107 & new_n3676;
  assign new_n13487 = n105 & new_n3688;
  assign new_n13488 = new_n13487 ^ new_n13486;
  assign new_n13489 = new_n13488 ^ new_n13485;
  assign new_n13490 = new_n13489 ^ n39;
  assign new_n13491 = ~new_n4212 & n103;
  assign new_n13492 = ~new_n4556 & new_n4201;
  assign new_n13493 = new_n13492 ^ new_n13491;
  assign new_n13494 = n104 & new_n4200;
  assign new_n13495 = n102 & new_n4206;
  assign new_n13496 = new_n13495 ^ new_n13494;
  assign new_n13497 = new_n13496 ^ new_n13493;
  assign new_n13498 = new_n13497 ^ n42;
  assign new_n13499 = ~new_n4804 & n100;
  assign new_n13500 = new_n3972 & new_n4799;
  assign new_n13501 = new_n13500 ^ new_n13499;
  assign new_n13502 = n101 & new_n4798;
  assign new_n13503 = n99 & new_n4810;
  assign new_n13504 = new_n13503 ^ new_n13502;
  assign new_n13505 = new_n13504 ^ new_n13501;
  assign new_n13506 = new_n13505 ^ n45;
  assign new_n13507 = ~new_n5424 & n97;
  assign new_n13508 = new_n3435 & new_n5419;
  assign new_n13509 = new_n13508 ^ new_n13507;
  assign new_n13510 = n98 & new_n5418;
  assign new_n13511 = n96 & new_n5648;
  assign new_n13512 = new_n13511 ^ new_n13510;
  assign new_n13513 = new_n13512 ^ new_n13509;
  assign new_n13514 = new_n13513 ^ n48;
  assign new_n13515 = ~new_n6110 & n94;
  assign new_n13516 = new_n2934 & new_n6105;
  assign new_n13517 = new_n13516 ^ new_n13515;
  assign new_n13518 = n95 & new_n6104;
  assign new_n13519 = n93 & new_n6347;
  assign new_n13520 = new_n13519 ^ new_n13518;
  assign new_n13521 = new_n13520 ^ new_n13517;
  assign new_n13522 = new_n13521 ^ n51;
  assign new_n13523 = ~new_n6805 & n91;
  assign new_n13524 = new_n2481 & new_n6800;
  assign new_n13525 = new_n13524 ^ new_n13523;
  assign new_n13526 = n92 & new_n6799;
  assign new_n13527 = n90 & new_n6811;
  assign new_n13528 = new_n13527 ^ new_n13526;
  assign new_n13529 = new_n13528 ^ new_n13525;
  assign new_n13530 = new_n13529 ^ n54;
  assign new_n13531 = n88 & new_n7553;
  assign new_n13532 = new_n2063 & new_n7543;
  assign new_n13533 = new_n13532 ^ new_n13531;
  assign new_n13534 = n89 & new_n7542;
  assign new_n13535 = n87 & new_n7547;
  assign new_n13536 = new_n13535 ^ new_n13534;
  assign new_n13537 = new_n13536 ^ new_n13533;
  assign new_n13538 = new_n13537 ^ n57;
  assign new_n13539 = n85 & new_n8355;
  assign new_n13540 = new_n1694 & new_n8345;
  assign new_n13541 = new_n13540 ^ new_n13539;
  assign new_n13542 = n86 & new_n8344;
  assign new_n13543 = n84 & new_n8349;
  assign new_n13544 = new_n13543 ^ new_n13542;
  assign new_n13545 = new_n13544 ^ new_n13541;
  assign new_n13546 = new_n13545 ^ n60;
  assign new_n13547 = n82 & new_n9195;
  assign new_n13548 = new_n1363 & new_n9185;
  assign new_n13549 = new_n13548 ^ new_n13547;
  assign new_n13550 = n83 & new_n9184;
  assign new_n13551 = n81 & new_n9189;
  assign new_n13552 = new_n13551 ^ new_n13550;
  assign new_n13553 = new_n13552 ^ new_n13549;
  assign new_n13554 = new_n13553 ^ n63;
  assign new_n13555 = new_n13305 ^ n80;
  assign new_n13556 = ~new_n9495 & new_n13555;
  assign new_n13557 = new_n13556 ^ n80;
  assign new_n13558 = new_n13557 ^ n15;
  assign new_n13559 = new_n13558 ^ new_n13077;
  assign new_n13560 = new_n13559 ^ new_n13554;
  assign new_n13561 = new_n13303 ^ n64;
  assign new_n13562 = new_n13303 ^ n63;
  assign new_n13563 = new_n13562 ^ new_n13561;
  assign new_n13564 = ~n77 & n78;
  assign new_n13565 = ~n78 & n77;
  assign new_n13566 = new_n13565 ^ new_n13564;
  assign new_n13567 = new_n13565 ^ new_n13561;
  assign new_n13568 = new_n13567 ^ new_n13565;
  assign new_n13569 = ~new_n13568 & new_n13566;
  assign new_n13570 = new_n13569 ^ new_n13565;
  assign new_n13571 = ~new_n13563 & new_n13570;
  assign new_n13572 = ~new_n13303 & new_n13571;
  assign new_n13573 = ~n79 & n78;
  assign new_n13574 = ~new_n13561 & new_n13573;
  assign new_n13575 = ~n78 & n79;
  assign new_n13576 = new_n13575 ^ new_n13564;
  assign new_n13577 = ~new_n13561 & new_n13576;
  assign new_n13578 = new_n13577 ^ new_n13575;
  assign new_n13579 = new_n13578 ^ new_n13574;
  assign new_n13580 = ~new_n13562 & ~new_n13579;
  assign new_n13581 = new_n13580 ^ new_n13574;
  assign new_n13582 = new_n13581 ^ new_n13572;
  assign new_n13583 = new_n13582 ^ new_n13560;
  assign new_n13584 = new_n13583 ^ new_n13546;
  assign new_n13585 = new_n13315 ^ new_n13296;
  assign new_n13586 = new_n13316 & new_n13585;
  assign new_n13587 = new_n13586 ^ new_n13296;
  assign new_n13588 = new_n13587 ^ new_n13584;
  assign new_n13589 = new_n13588 ^ new_n13538;
  assign new_n13590 = new_n13321 ^ new_n13317;
  assign new_n13591 = ~new_n13318 & new_n13590;
  assign new_n13592 = new_n13591 ^ new_n13288;
  assign new_n13593 = new_n13592 ^ new_n13589;
  assign new_n13594 = new_n13593 ^ new_n13530;
  assign new_n13595 = new_n13322 ^ new_n13279;
  assign new_n13596 = ~new_n13280 & ~new_n13595;
  assign new_n13597 = new_n13596 ^ new_n13276;
  assign new_n13598 = new_n13597 ^ new_n13594;
  assign new_n13599 = new_n13598 ^ new_n13522;
  assign new_n13600 = new_n13327 ^ new_n13323;
  assign new_n13601 = ~new_n13600 & new_n13324;
  assign new_n13602 = new_n13601 ^ new_n13268;
  assign new_n13603 = new_n13602 ^ new_n13599;
  assign new_n13604 = new_n13603 ^ new_n13514;
  assign new_n13605 = new_n13332 ^ new_n13328;
  assign new_n13606 = ~new_n13605 & new_n13329;
  assign new_n13607 = new_n13606 ^ new_n13260;
  assign new_n13608 = new_n13607 ^ new_n13604;
  assign new_n13609 = new_n13608 ^ new_n13506;
  assign new_n13610 = new_n13337 ^ new_n13333;
  assign new_n13611 = ~new_n13610 & new_n13334;
  assign new_n13612 = new_n13611 ^ new_n13252;
  assign new_n13613 = new_n13612 ^ new_n13609;
  assign new_n13614 = new_n13613 ^ new_n13498;
  assign new_n13615 = new_n13338 ^ new_n13244;
  assign new_n13616 = ~new_n13342 & new_n13615;
  assign new_n13617 = new_n13616 ^ new_n13244;
  assign new_n13618 = new_n13617 ^ new_n13614;
  assign new_n13619 = new_n13618 ^ new_n13490;
  assign new_n13620 = new_n13343 ^ new_n13236;
  assign new_n13621 = ~new_n13347 & new_n13620;
  assign new_n13622 = new_n13621 ^ new_n13236;
  assign new_n13623 = new_n13622 ^ new_n13619;
  assign new_n13624 = new_n13623 ^ new_n13482;
  assign new_n13625 = new_n13348 ^ new_n13228;
  assign new_n13626 = ~new_n13352 & new_n13625;
  assign new_n13627 = new_n13626 ^ new_n13228;
  assign new_n13628 = new_n13627 ^ new_n13624;
  assign new_n13629 = new_n13628 ^ new_n13474;
  assign new_n13630 = new_n13356 ^ new_n13220;
  assign new_n13631 = ~new_n13357 & new_n13630;
  assign new_n13632 = new_n13631 ^ new_n13220;
  assign new_n13633 = new_n13632 ^ new_n13629;
  assign new_n13634 = new_n13633 ^ new_n13466;
  assign new_n13635 = new_n13370 ^ new_n13358;
  assign new_n13636 = ~new_n13635 & new_n13362;
  assign new_n13637 = new_n13636 ^ new_n13361;
  assign new_n13638 = new_n13637 ^ new_n13634;
  assign new_n13639 = new_n13638 ^ new_n13458;
  assign new_n13640 = new_n13383 ^ new_n13371;
  assign new_n13641 = ~new_n13640 & new_n13375;
  assign new_n13642 = new_n13641 ^ new_n13374;
  assign new_n13643 = new_n13642 ^ new_n13639;
  assign new_n13644 = ~new_n1506 & n121;
  assign new_n13645 = new_n1501 & new_n8850;
  assign new_n13646 = new_n13645 ^ new_n13644;
  assign new_n13647 = n122 & new_n1500;
  assign new_n13648 = n120 & new_n1512;
  assign new_n13649 = new_n13648 ^ new_n13647;
  assign new_n13650 = new_n13649 ^ new_n13646;
  assign new_n13651 = new_n13650 ^ n24;
  assign new_n13652 = new_n13651 ^ new_n13643;
  assign new_n13653 = new_n13396 ^ new_n13384;
  assign new_n13654 = ~new_n13393 & new_n13653;
  assign new_n13655 = new_n13654 ^ new_n13396;
  assign new_n13656 = new_n13655 ^ new_n13652;
  assign new_n13657 = ~new_n1198 & n124;
  assign new_n13658 = new_n1193 & new_n9700;
  assign new_n13659 = new_n13658 ^ new_n13657;
  assign new_n13660 = n125 & new_n1192;
  assign new_n13661 = n123 & new_n1204;
  assign new_n13662 = new_n13661 ^ new_n13660;
  assign new_n13663 = new_n13662 ^ new_n13659;
  assign new_n13664 = new_n13663 ^ n21;
  assign new_n13665 = new_n13664 ^ new_n13656;
  assign new_n13666 = new_n13409 ^ new_n13397;
  assign new_n13667 = ~new_n13401 & ~new_n13666;
  assign new_n13668 = new_n13667 ^ new_n13400;
  assign new_n13669 = new_n13668 ^ new_n13665;
  assign new_n13670 = ~new_n930 & n127;
  assign new_n13671 = new_n925 & new_n10581;
  assign new_n13672 = new_n13671 ^ new_n13670;
  assign new_n13673 = n128 & new_n924;
  assign new_n13674 = n126 & new_n936;
  assign new_n13675 = new_n13674 ^ new_n13673;
  assign new_n13676 = new_n13675 ^ new_n13672;
  assign new_n13677 = new_n13676 ^ n18;
  assign new_n13678 = new_n13677 ^ new_n13669;
  assign new_n13679 = new_n13422 ^ new_n13410;
  assign new_n13680 = ~new_n13414 & new_n13679;
  assign new_n13681 = new_n13680 ^ new_n13413;
  assign new_n13682 = new_n13681 ^ new_n13678;
  assign new_n13683 = new_n13682 ^ new_n13450;
  assign new_n13684 = ~new_n13448 & new_n13447;
  assign new_n13685 = ~new_n13684 & new_n13682;
  assign new_n13686 = ~new_n13442 & ~new_n13685;
  assign new_n13687 = new_n13448 ^ new_n13431;
  assign new_n13688 = new_n13438 ^ new_n13434;
  assign new_n13689 = new_n13688 ^ new_n13447;
  assign new_n13690 = ~new_n13682 & new_n13689;
  assign new_n13691 = ~new_n13687 & ~new_n13690;
  assign new_n13692 = ~new_n13686 & new_n13691;
  assign new_n13693 = ~new_n13448 & ~new_n13682;
  assign new_n13694 = new_n13442 ^ new_n13438;
  assign new_n13695 = ~new_n13694 & new_n13688;
  assign new_n13696 = new_n13695 ^ new_n13438;
  assign new_n13697 = ~new_n13693 & ~new_n13696;
  assign new_n13698 = ~new_n13692 & ~new_n13697;
  assign new_n13699 = n119 & new_n1874;
  assign new_n13700 = new_n1864 & new_n8286;
  assign new_n13701 = new_n13700 ^ new_n13699;
  assign new_n13702 = n120 & new_n1863;
  assign new_n13703 = n118 & new_n1868;
  assign new_n13704 = new_n13703 ^ new_n13702;
  assign new_n13705 = new_n13704 ^ new_n13701;
  assign new_n13706 = new_n13705 ^ n27;
  assign new_n13707 = n116 & new_n2246;
  assign new_n13708 = ~new_n7503 & new_n2241;
  assign new_n13709 = new_n13708 ^ new_n13707;
  assign new_n13710 = n117 & new_n2240;
  assign new_n13711 = n115 & new_n2391;
  assign new_n13712 = new_n13711 ^ new_n13710;
  assign new_n13713 = new_n13712 ^ new_n13709;
  assign new_n13714 = new_n13713 ^ n30;
  assign new_n13715 = ~new_n2672 & n113;
  assign new_n13716 = ~new_n6764 & new_n2667;
  assign new_n13717 = new_n13716 ^ new_n13715;
  assign new_n13718 = n114 & new_n2666;
  assign new_n13719 = n112 & new_n2664;
  assign new_n13720 = new_n13719 ^ new_n13718;
  assign new_n13721 = new_n13720 ^ new_n13717;
  assign new_n13722 = new_n13721 ^ n33;
  assign new_n13723 = ~new_n3143 & n110;
  assign new_n13724 = new_n3138 & new_n6049;
  assign new_n13725 = new_n13724 ^ new_n13723;
  assign new_n13726 = n111 & new_n3137;
  assign new_n13727 = n109 & new_n3149;
  assign new_n13728 = new_n13727 ^ new_n13726;
  assign new_n13729 = new_n13728 ^ new_n13725;
  assign new_n13730 = new_n13729 ^ n36;
  assign new_n13731 = new_n13622 ^ new_n13490;
  assign new_n13732 = ~new_n13619 & new_n13731;
  assign new_n13733 = new_n13732 ^ new_n13622;
  assign new_n13734 = new_n13733 ^ new_n13730;
  assign new_n13735 = ~new_n3682 & n107;
  assign new_n13736 = ~new_n5377 & new_n3677;
  assign new_n13737 = new_n13736 ^ new_n13735;
  assign new_n13738 = n108 & new_n3676;
  assign new_n13739 = n106 & new_n3688;
  assign new_n13740 = new_n13739 ^ new_n13738;
  assign new_n13741 = new_n13740 ^ new_n13737;
  assign new_n13742 = new_n13741 ^ n39;
  assign new_n13743 = ~new_n4212 & n104;
  assign new_n13744 = ~new_n4754 & new_n4201;
  assign new_n13745 = new_n13744 ^ new_n13743;
  assign new_n13746 = n105 & new_n4200;
  assign new_n13747 = n103 & new_n4206;
  assign new_n13748 = new_n13747 ^ new_n13746;
  assign new_n13749 = new_n13748 ^ new_n13745;
  assign new_n13750 = new_n13749 ^ n42;
  assign new_n13751 = ~new_n4804 & n101;
  assign new_n13752 = new_n4159 & new_n4799;
  assign new_n13753 = new_n13752 ^ new_n13751;
  assign new_n13754 = n102 & new_n4798;
  assign new_n13755 = n100 & new_n4810;
  assign new_n13756 = new_n13755 ^ new_n13754;
  assign new_n13757 = new_n13756 ^ new_n13753;
  assign new_n13758 = new_n13757 ^ n45;
  assign new_n13759 = new_n13607 ^ new_n13514;
  assign new_n13760 = ~new_n13604 & new_n13759;
  assign new_n13761 = new_n13760 ^ new_n13607;
  assign new_n13762 = new_n13761 ^ new_n13758;
  assign new_n13763 = ~new_n5424 & n98;
  assign new_n13764 = new_n3604 & new_n5419;
  assign new_n13765 = new_n13764 ^ new_n13763;
  assign new_n13766 = n99 & new_n5418;
  assign new_n13767 = n97 & new_n5648;
  assign new_n13768 = new_n13767 ^ new_n13766;
  assign new_n13769 = new_n13768 ^ new_n13765;
  assign new_n13770 = new_n13769 ^ n48;
  assign new_n13771 = ~new_n6110 & n95;
  assign new_n13772 = new_n3095 & new_n6105;
  assign new_n13773 = new_n13772 ^ new_n13771;
  assign new_n13774 = n96 & new_n6104;
  assign new_n13775 = n94 & new_n6347;
  assign new_n13776 = new_n13775 ^ new_n13774;
  assign new_n13777 = new_n13776 ^ new_n13773;
  assign new_n13778 = new_n13777 ^ n51;
  assign new_n13779 = ~new_n6805 & n92;
  assign new_n13780 = new_n2628 & new_n6800;
  assign new_n13781 = new_n13780 ^ new_n13779;
  assign new_n13782 = n93 & new_n6799;
  assign new_n13783 = n91 & new_n6811;
  assign new_n13784 = new_n13783 ^ new_n13782;
  assign new_n13785 = new_n13784 ^ new_n13781;
  assign new_n13786 = new_n13785 ^ n54;
  assign new_n13787 = new_n13592 ^ new_n13538;
  assign new_n13788 = ~new_n13589 & new_n13787;
  assign new_n13789 = new_n13788 ^ new_n13592;
  assign new_n13790 = new_n13789 ^ new_n13786;
  assign new_n13791 = n89 & new_n7553;
  assign new_n13792 = new_n2193 & new_n7543;
  assign new_n13793 = new_n13792 ^ new_n13791;
  assign new_n13794 = n90 & new_n7542;
  assign new_n13795 = n88 & new_n7547;
  assign new_n13796 = new_n13795 ^ new_n13794;
  assign new_n13797 = new_n13796 ^ new_n13793;
  assign new_n13798 = new_n13797 ^ n57;
  assign new_n13799 = new_n13587 ^ new_n13546;
  assign new_n13800 = ~new_n13584 & new_n13799;
  assign new_n13801 = new_n13800 ^ new_n13587;
  assign new_n13802 = new_n13801 ^ new_n13798;
  assign new_n13803 = n86 & new_n8355;
  assign new_n13804 = new_n1811 & new_n8345;
  assign new_n13805 = new_n13804 ^ new_n13803;
  assign new_n13806 = n87 & new_n8344;
  assign new_n13807 = n85 & new_n8349;
  assign new_n13808 = new_n13807 ^ new_n13806;
  assign new_n13809 = new_n13808 ^ new_n13805;
  assign new_n13810 = new_n13809 ^ n60;
  assign new_n13811 = n83 & new_n9195;
  assign new_n13812 = new_n1468 & new_n9185;
  assign new_n13813 = new_n13812 ^ new_n13811;
  assign new_n13814 = n84 & new_n9184;
  assign new_n13815 = n82 & new_n9189;
  assign new_n13816 = new_n13815 ^ new_n13814;
  assign new_n13817 = new_n13816 ^ new_n13813;
  assign new_n13818 = new_n13077 ^ n15;
  assign new_n13819 = new_n13557 ^ new_n13077;
  assign new_n13820 = ~new_n13818 & ~new_n13819;
  assign new_n13821 = new_n13820 ^ n15;
  assign new_n13822 = n64 & n81;
  assign new_n13823 = ~n64 & new_n995;
  assign new_n13824 = new_n13823 ^ n80;
  assign new_n13825 = new_n13824 ^ new_n13822;
  assign new_n13826 = ~n63 & ~new_n13825;
  assign new_n13827 = new_n13826 ^ new_n13824;
  assign new_n13828 = new_n13827 ^ new_n13821;
  assign new_n13829 = new_n13828 ^ new_n13817;
  assign new_n13830 = new_n13829 ^ new_n13810;
  assign new_n13831 = new_n13582 ^ new_n13554;
  assign new_n13832 = ~new_n13831 & new_n13560;
  assign new_n13833 = new_n13832 ^ new_n13582;
  assign new_n13834 = new_n13833 ^ new_n13830;
  assign new_n13835 = new_n13834 ^ new_n13802;
  assign new_n13836 = new_n13835 ^ new_n13790;
  assign new_n13837 = new_n13836 ^ new_n13778;
  assign new_n13838 = new_n13597 ^ new_n13530;
  assign new_n13839 = ~new_n13594 & new_n13838;
  assign new_n13840 = new_n13839 ^ new_n13597;
  assign new_n13841 = new_n13840 ^ new_n13837;
  assign new_n13842 = new_n13841 ^ new_n13770;
  assign new_n13843 = new_n13602 ^ new_n13522;
  assign new_n13844 = ~new_n13599 & new_n13843;
  assign new_n13845 = new_n13844 ^ new_n13602;
  assign new_n13846 = new_n13845 ^ new_n13842;
  assign new_n13847 = new_n13846 ^ new_n13762;
  assign new_n13848 = new_n13612 ^ new_n13506;
  assign new_n13849 = ~new_n13609 & new_n13848;
  assign new_n13850 = new_n13849 ^ new_n13612;
  assign new_n13851 = new_n13850 ^ new_n13847;
  assign new_n13852 = new_n13851 ^ new_n13750;
  assign new_n13853 = new_n13617 ^ new_n13613;
  assign new_n13854 = ~new_n13853 & new_n13614;
  assign new_n13855 = new_n13854 ^ new_n13498;
  assign new_n13856 = new_n13855 ^ new_n13852;
  assign new_n13857 = new_n13856 ^ new_n13742;
  assign new_n13858 = new_n13857 ^ new_n13734;
  assign new_n13859 = new_n13627 ^ new_n13482;
  assign new_n13860 = ~new_n13624 & new_n13859;
  assign new_n13861 = new_n13860 ^ new_n13627;
  assign new_n13862 = new_n13861 ^ new_n13858;
  assign new_n13863 = new_n13862 ^ new_n13722;
  assign new_n13864 = new_n13632 ^ new_n13474;
  assign new_n13865 = ~new_n13629 & new_n13864;
  assign new_n13866 = new_n13865 ^ new_n13632;
  assign new_n13867 = new_n13866 ^ new_n13863;
  assign new_n13868 = new_n13867 ^ new_n13714;
  assign new_n13869 = new_n13868 ^ new_n13706;
  assign new_n13870 = new_n13637 ^ new_n13466;
  assign new_n13871 = ~new_n13634 & new_n13870;
  assign new_n13872 = new_n13871 ^ new_n13637;
  assign new_n13873 = new_n13872 ^ new_n13869;
  assign new_n13874 = new_n13642 ^ new_n13458;
  assign new_n13875 = ~new_n13639 & new_n13874;
  assign new_n13876 = new_n13875 ^ new_n13642;
  assign new_n13877 = new_n13876 ^ new_n13873;
  assign new_n13878 = ~new_n1506 & n122;
  assign new_n13879 = ~new_n9116 & new_n1501;
  assign new_n13880 = new_n13879 ^ new_n13878;
  assign new_n13881 = n123 & new_n1500;
  assign new_n13882 = n121 & new_n1512;
  assign new_n13883 = new_n13882 ^ new_n13881;
  assign new_n13884 = new_n13883 ^ new_n13880;
  assign new_n13885 = new_n13884 ^ n24;
  assign new_n13886 = new_n13885 ^ new_n13877;
  assign new_n13887 = new_n13655 ^ new_n13643;
  assign new_n13888 = ~new_n13652 & new_n13887;
  assign new_n13889 = new_n13888 ^ new_n13655;
  assign new_n13890 = new_n13889 ^ new_n13886;
  assign new_n13891 = ~new_n1198 & n125;
  assign new_n13892 = new_n1193 & new_n9987;
  assign new_n13893 = new_n13892 ^ new_n13891;
  assign new_n13894 = n126 & new_n1192;
  assign new_n13895 = n124 & new_n1204;
  assign new_n13896 = new_n13895 ^ new_n13894;
  assign new_n13897 = new_n13896 ^ new_n13893;
  assign new_n13898 = new_n13897 ^ n21;
  assign new_n13899 = new_n13898 ^ new_n13890;
  assign new_n13900 = new_n13668 ^ new_n13656;
  assign new_n13901 = ~new_n13665 & ~new_n13900;
  assign new_n13902 = new_n13901 ^ new_n13668;
  assign new_n13903 = new_n13902 ^ new_n13899;
  assign new_n13904 = n127 & new_n936;
  assign new_n13905 = new_n925 & new_n10010;
  assign new_n13906 = new_n13905 ^ new_n13904;
  assign new_n13907 = ~new_n930 & n128;
  assign new_n13908 = new_n13907 ^ new_n13906;
  assign new_n13909 = new_n13908 ^ n18;
  assign new_n13910 = new_n13909 ^ new_n13903;
  assign new_n13911 = new_n13681 ^ new_n13669;
  assign new_n13912 = ~new_n13911 & new_n13678;
  assign new_n13913 = new_n13912 ^ new_n13681;
  assign new_n13914 = new_n13913 ^ new_n13910;
  assign new_n13915 = new_n13914 ^ new_n13698;
  assign new_n13916 = new_n13899 & new_n13909;
  assign new_n13917 = new_n13909 ^ new_n13899;
  assign new_n13918 = new_n13917 ^ new_n13916;
  assign new_n13919 = new_n13913 ^ new_n13902;
  assign new_n13920 = ~new_n13902 & new_n13913;
  assign new_n13921 = new_n13920 ^ new_n13919;
  assign new_n13922 = ~new_n13918 & ~new_n13921;
  assign new_n13923 = new_n13916 ^ new_n13698;
  assign new_n13924 = new_n13921 ^ new_n13916;
  assign new_n13925 = ~new_n13923 & ~new_n13924;
  assign new_n13926 = new_n13925 ^ new_n13922;
  assign new_n13927 = ~new_n13920 & new_n13916;
  assign new_n13928 = new_n13918 ^ new_n13698;
  assign new_n13929 = new_n13920 ^ new_n13918;
  assign new_n13930 = ~new_n13928 & new_n13929;
  assign new_n13931 = new_n13930 ^ new_n13927;
  assign new_n13932 = new_n13931 ^ new_n13926;
  assign new_n13933 = ~new_n1198 & n126;
  assign new_n13934 = new_n1193 & new_n10304;
  assign new_n13935 = new_n13934 ^ new_n13933;
  assign new_n13936 = n127 & new_n1192;
  assign new_n13937 = n125 & new_n1204;
  assign new_n13938 = new_n13937 ^ new_n13936;
  assign new_n13939 = new_n13938 ^ new_n13935;
  assign new_n13940 = new_n13939 ^ n21;
  assign new_n13941 = ~new_n1506 & n123;
  assign new_n13942 = ~new_n9405 & new_n1501;
  assign new_n13943 = new_n13942 ^ new_n13941;
  assign new_n13944 = n124 & new_n1500;
  assign new_n13945 = n122 & new_n1512;
  assign new_n13946 = new_n13945 ^ new_n13944;
  assign new_n13947 = new_n13946 ^ new_n13943;
  assign new_n13948 = new_n13947 ^ n24;
  assign new_n13949 = n120 & new_n1874;
  assign new_n13950 = new_n1864 & new_n8560;
  assign new_n13951 = new_n13950 ^ new_n13949;
  assign new_n13952 = n121 & new_n1863;
  assign new_n13953 = n119 & new_n1868;
  assign new_n13954 = new_n13953 ^ new_n13952;
  assign new_n13955 = new_n13954 ^ new_n13951;
  assign new_n13956 = new_n13955 ^ n27;
  assign new_n13957 = n117 & new_n2246;
  assign new_n13958 = ~new_n7761 & new_n2241;
  assign new_n13959 = new_n13958 ^ new_n13957;
  assign new_n13960 = n118 & new_n2240;
  assign new_n13961 = n116 & new_n2391;
  assign new_n13962 = new_n13961 ^ new_n13960;
  assign new_n13963 = new_n13962 ^ new_n13959;
  assign new_n13964 = new_n13963 ^ n30;
  assign new_n13965 = ~new_n2672 & n114;
  assign new_n13966 = ~new_n7013 & new_n2667;
  assign new_n13967 = new_n13966 ^ new_n13965;
  assign new_n13968 = n115 & new_n2666;
  assign new_n13969 = n113 & new_n2664;
  assign new_n13970 = new_n13969 ^ new_n13968;
  assign new_n13971 = new_n13970 ^ new_n13967;
  assign new_n13972 = new_n13971 ^ n33;
  assign new_n13973 = ~new_n3143 & n111;
  assign new_n13974 = ~new_n6284 & new_n3138;
  assign new_n13975 = new_n13974 ^ new_n13973;
  assign new_n13976 = n112 & new_n3137;
  assign new_n13977 = n110 & new_n3149;
  assign new_n13978 = new_n13977 ^ new_n13976;
  assign new_n13979 = new_n13978 ^ new_n13975;
  assign new_n13980 = new_n13979 ^ n36;
  assign new_n13981 = ~new_n3682 & n108;
  assign new_n13982 = new_n3677 & new_n5604;
  assign new_n13983 = new_n13982 ^ new_n13981;
  assign new_n13984 = n109 & new_n3676;
  assign new_n13985 = n107 & new_n3688;
  assign new_n13986 = new_n13985 ^ new_n13984;
  assign new_n13987 = new_n13986 ^ new_n13983;
  assign new_n13988 = new_n13987 ^ n39;
  assign new_n13989 = ~new_n4212 & n105;
  assign new_n13990 = ~new_n4961 & new_n4201;
  assign new_n13991 = new_n13990 ^ new_n13989;
  assign new_n13992 = n106 & new_n4200;
  assign new_n13993 = n104 & new_n4206;
  assign new_n13994 = new_n13993 ^ new_n13992;
  assign new_n13995 = new_n13994 ^ new_n13991;
  assign new_n13996 = new_n13995 ^ n42;
  assign new_n13997 = ~new_n4804 & n102;
  assign new_n13998 = new_n4368 & new_n4799;
  assign new_n13999 = new_n13998 ^ new_n13997;
  assign new_n14000 = n103 & new_n4798;
  assign new_n14001 = n101 & new_n4810;
  assign new_n14002 = new_n14001 ^ new_n14000;
  assign new_n14003 = new_n14002 ^ new_n13999;
  assign new_n14004 = new_n14003 ^ n45;
  assign new_n14005 = ~new_n5424 & n99;
  assign new_n14006 = new_n3789 & new_n5419;
  assign new_n14007 = new_n14006 ^ new_n14005;
  assign new_n14008 = n100 & new_n5418;
  assign new_n14009 = n98 & new_n5648;
  assign new_n14010 = new_n14009 ^ new_n14008;
  assign new_n14011 = new_n14010 ^ new_n14007;
  assign new_n14012 = new_n14011 ^ n48;
  assign new_n14013 = new_n13840 ^ new_n13836;
  assign new_n14014 = ~new_n14013 & new_n13837;
  assign new_n14015 = new_n14014 ^ new_n13778;
  assign new_n14016 = new_n14015 ^ new_n14012;
  assign new_n14017 = ~new_n6110 & n96;
  assign new_n14018 = new_n3273 & new_n6105;
  assign new_n14019 = new_n14018 ^ new_n14017;
  assign new_n14020 = n97 & new_n6104;
  assign new_n14021 = n95 & new_n6347;
  assign new_n14022 = new_n14021 ^ new_n14020;
  assign new_n14023 = new_n14022 ^ new_n14019;
  assign new_n14024 = new_n14023 ^ n51;
  assign new_n14025 = ~new_n6805 & n93;
  assign new_n14026 = new_n2785 & new_n6800;
  assign new_n14027 = new_n14026 ^ new_n14025;
  assign new_n14028 = n94 & new_n6799;
  assign new_n14029 = n92 & new_n6811;
  assign new_n14030 = new_n14029 ^ new_n14028;
  assign new_n14031 = new_n14030 ^ new_n14027;
  assign new_n14032 = new_n14031 ^ n54;
  assign new_n14033 = n90 & new_n7553;
  assign new_n14034 = new_n2341 & new_n7543;
  assign new_n14035 = new_n14034 ^ new_n14033;
  assign new_n14036 = n91 & new_n7542;
  assign new_n14037 = n89 & new_n7547;
  assign new_n14038 = new_n14037 ^ new_n14036;
  assign new_n14039 = new_n14038 ^ new_n14035;
  assign new_n14040 = new_n14039 ^ n57;
  assign new_n14041 = n87 & new_n8355;
  assign new_n14042 = new_n1940 & new_n8345;
  assign new_n14043 = new_n14042 ^ new_n14041;
  assign new_n14044 = n88 & new_n8344;
  assign new_n14045 = n86 & new_n8349;
  assign new_n14046 = new_n14045 ^ new_n14044;
  assign new_n14047 = new_n14046 ^ new_n14043;
  assign new_n14048 = new_n14047 ^ n60;
  assign new_n14049 = n84 & new_n9195;
  assign new_n14050 = new_n1584 & new_n9185;
  assign new_n14051 = new_n14050 ^ new_n14049;
  assign new_n14052 = n85 & new_n9184;
  assign new_n14053 = n83 & new_n9189;
  assign new_n14054 = new_n14053 ^ new_n14052;
  assign new_n14055 = new_n14054 ^ new_n14051;
  assign new_n14056 = new_n1087 ^ n63;
  assign new_n14057 = new_n13824 ^ n81;
  assign new_n14058 = new_n14057 ^ new_n1087;
  assign new_n14059 = ~new_n9495 & new_n14058;
  assign new_n14060 = new_n14059 ^ new_n14056;
  assign new_n14061 = new_n14060 ^ new_n14055;
  assign new_n14062 = new_n13821 ^ new_n13817;
  assign new_n14063 = new_n13822 ^ new_n13817;
  assign new_n14064 = ~new_n14062 & ~new_n14063;
  assign new_n14065 = new_n14064 ^ new_n13817;
  assign new_n14066 = new_n13824 ^ new_n13817;
  assign new_n14067 = new_n14062 & new_n14066;
  assign new_n14068 = new_n14067 ^ new_n13817;
  assign new_n14069 = new_n14068 ^ new_n14065;
  assign new_n14070 = ~new_n14069 & n63;
  assign new_n14071 = new_n14070 ^ new_n14065;
  assign new_n14072 = new_n14071 ^ new_n14061;
  assign new_n14073 = new_n14072 ^ new_n14048;
  assign new_n14074 = new_n13833 ^ new_n13829;
  assign new_n14075 = ~new_n13830 & ~new_n14074;
  assign new_n14076 = new_n14075 ^ new_n13810;
  assign new_n14077 = new_n14076 ^ new_n14073;
  assign new_n14078 = new_n14077 ^ new_n14040;
  assign new_n14079 = new_n14078 ^ new_n14032;
  assign new_n14080 = new_n13834 ^ new_n13801;
  assign new_n14081 = ~new_n14080 & new_n13802;
  assign new_n14082 = new_n14081 ^ new_n13798;
  assign new_n14083 = new_n14082 ^ new_n14079;
  assign new_n14084 = new_n14083 ^ new_n14024;
  assign new_n14085 = new_n13835 ^ new_n13786;
  assign new_n14086 = ~new_n14085 & new_n13790;
  assign new_n14087 = new_n14086 ^ new_n13789;
  assign new_n14088 = new_n14087 ^ new_n14084;
  assign new_n14089 = new_n14088 ^ new_n14016;
  assign new_n14090 = new_n14089 ^ new_n14004;
  assign new_n14091 = new_n13845 ^ new_n13841;
  assign new_n14092 = ~new_n14091 & new_n13842;
  assign new_n14093 = new_n14092 ^ new_n13770;
  assign new_n14094 = new_n14093 ^ new_n14090;
  assign new_n14095 = new_n13846 ^ new_n13761;
  assign new_n14096 = ~new_n14095 & new_n13762;
  assign new_n14097 = new_n14096 ^ new_n13758;
  assign new_n14098 = new_n14097 ^ new_n14094;
  assign new_n14099 = new_n14098 ^ new_n13996;
  assign new_n14100 = new_n13850 ^ new_n13750;
  assign new_n14101 = ~new_n13851 & new_n14100;
  assign new_n14102 = new_n14101 ^ new_n13750;
  assign new_n14103 = new_n14102 ^ new_n14099;
  assign new_n14104 = new_n14103 ^ new_n13988;
  assign new_n14105 = new_n13855 ^ new_n13742;
  assign new_n14106 = ~new_n13856 & new_n14105;
  assign new_n14107 = new_n14106 ^ new_n13742;
  assign new_n14108 = new_n14107 ^ new_n14104;
  assign new_n14109 = new_n14108 ^ new_n13980;
  assign new_n14110 = new_n13857 ^ new_n13730;
  assign new_n14111 = ~new_n14110 & new_n13734;
  assign new_n14112 = new_n14111 ^ new_n13733;
  assign new_n14113 = new_n14112 ^ new_n14109;
  assign new_n14114 = new_n14113 ^ new_n13972;
  assign new_n14115 = new_n13858 ^ new_n13722;
  assign new_n14116 = ~new_n13862 & new_n14115;
  assign new_n14117 = new_n14116 ^ new_n13722;
  assign new_n14118 = new_n14117 ^ new_n14114;
  assign new_n14119 = new_n14118 ^ new_n13964;
  assign new_n14120 = new_n13866 ^ new_n13714;
  assign new_n14121 = ~new_n13867 & new_n14120;
  assign new_n14122 = new_n14121 ^ new_n13714;
  assign new_n14123 = new_n14122 ^ new_n14119;
  assign new_n14124 = new_n14123 ^ new_n13956;
  assign new_n14125 = new_n13872 ^ new_n13706;
  assign new_n14126 = ~new_n13869 & new_n14125;
  assign new_n14127 = new_n14126 ^ new_n13872;
  assign new_n14128 = new_n14127 ^ new_n14124;
  assign new_n14129 = new_n14128 ^ new_n13948;
  assign new_n14130 = new_n13885 ^ new_n13873;
  assign new_n14131 = ~new_n14130 & new_n13877;
  assign new_n14132 = new_n14131 ^ new_n13876;
  assign new_n14133 = new_n14132 ^ new_n14129;
  assign new_n14134 = new_n14133 ^ new_n13940;
  assign new_n14135 = ~new_n935 & n128;
  assign new_n14136 = ~n18 & ~new_n14135;
  assign new_n14137 = new_n14136 ^ n17;
  assign new_n14138 = new_n778 & new_n11133;
  assign new_n14139 = new_n14138 ^ new_n14135;
  assign new_n14140 = ~new_n14137 & ~new_n14139;
  assign new_n14141 = new_n14140 ^ n17;
  assign new_n14142 = new_n14141 ^ new_n14134;
  assign new_n14143 = new_n13898 ^ new_n13886;
  assign new_n14144 = ~new_n14143 & new_n13890;
  assign new_n14145 = new_n14144 ^ new_n13889;
  assign new_n14146 = new_n14145 ^ new_n14142;
  assign new_n14147 = new_n14146 ^ new_n13932;
  assign new_n14148 = ~new_n13918 & ~new_n13920;
  assign new_n14149 = ~new_n14146 & ~new_n14148;
  assign new_n14150 = ~new_n13698 & ~new_n14149;
  assign new_n14151 = ~new_n13916 & new_n14146;
  assign new_n14152 = ~new_n13921 & ~new_n14151;
  assign new_n14153 = ~new_n14150 & new_n14152;
  assign new_n14154 = ~new_n13920 & new_n14146;
  assign new_n14155 = new_n13899 ^ new_n13698;
  assign new_n14156 = new_n13917 & new_n14155;
  assign new_n14157 = new_n14156 ^ new_n13899;
  assign new_n14158 = ~new_n14154 & new_n14157;
  assign new_n14159 = ~new_n14153 & ~new_n14158;
  assign new_n14160 = ~new_n1198 & n127;
  assign new_n14161 = new_n1193 & new_n10581;
  assign new_n14162 = new_n14161 ^ new_n14160;
  assign new_n14163 = n128 & new_n1192;
  assign new_n14164 = n126 & new_n1204;
  assign new_n14165 = new_n14164 ^ new_n14163;
  assign new_n14166 = new_n14165 ^ new_n14162;
  assign new_n14167 = new_n14166 ^ n21;
  assign new_n14168 = ~new_n1506 & n124;
  assign new_n14169 = new_n1501 & new_n9700;
  assign new_n14170 = new_n14169 ^ new_n14168;
  assign new_n14171 = n125 & new_n1500;
  assign new_n14172 = n123 & new_n1512;
  assign new_n14173 = new_n14172 ^ new_n14171;
  assign new_n14174 = new_n14173 ^ new_n14170;
  assign new_n14175 = new_n14174 ^ n24;
  assign new_n14176 = n118 & new_n2246;
  assign new_n14177 = ~new_n8019 & new_n2241;
  assign new_n14178 = new_n14177 ^ new_n14176;
  assign new_n14179 = n119 & new_n2240;
  assign new_n14180 = n117 & new_n2391;
  assign new_n14181 = new_n14180 ^ new_n14179;
  assign new_n14182 = new_n14181 ^ new_n14178;
  assign new_n14183 = new_n14182 ^ n30;
  assign new_n14184 = ~new_n2672 & n115;
  assign new_n14185 = ~new_n7256 & new_n2667;
  assign new_n14186 = new_n14185 ^ new_n14184;
  assign new_n14187 = n116 & new_n2666;
  assign new_n14188 = n114 & new_n2664;
  assign new_n14189 = new_n14188 ^ new_n14187;
  assign new_n14190 = new_n14189 ^ new_n14186;
  assign new_n14191 = new_n14190 ^ n33;
  assign new_n14192 = ~new_n3143 & n112;
  assign new_n14193 = ~new_n6518 & new_n3138;
  assign new_n14194 = new_n14193 ^ new_n14192;
  assign new_n14195 = n113 & new_n3137;
  assign new_n14196 = n111 & new_n3149;
  assign new_n14197 = new_n14196 ^ new_n14195;
  assign new_n14198 = new_n14197 ^ new_n14194;
  assign new_n14199 = new_n14198 ^ n36;
  assign new_n14200 = ~new_n3682 & n109;
  assign new_n14201 = new_n3677 & new_n5825;
  assign new_n14202 = new_n14201 ^ new_n14200;
  assign new_n14203 = n110 & new_n3676;
  assign new_n14204 = n108 & new_n3688;
  assign new_n14205 = new_n14204 ^ new_n14203;
  assign new_n14206 = new_n14205 ^ new_n14202;
  assign new_n14207 = new_n14206 ^ n39;
  assign new_n14208 = ~new_n4212 & n106;
  assign new_n14209 = ~new_n5164 & new_n4201;
  assign new_n14210 = new_n14209 ^ new_n14208;
  assign new_n14211 = n107 & new_n4200;
  assign new_n14212 = n105 & new_n4206;
  assign new_n14213 = new_n14212 ^ new_n14211;
  assign new_n14214 = new_n14213 ^ new_n14210;
  assign new_n14215 = new_n14214 ^ n42;
  assign new_n14216 = ~new_n4804 & n103;
  assign new_n14217 = ~new_n4556 & new_n4799;
  assign new_n14218 = new_n14217 ^ new_n14216;
  assign new_n14219 = n104 & new_n4798;
  assign new_n14220 = n102 & new_n4810;
  assign new_n14221 = new_n14220 ^ new_n14219;
  assign new_n14222 = new_n14221 ^ new_n14218;
  assign new_n14223 = new_n14222 ^ n45;
  assign new_n14224 = ~new_n5424 & n100;
  assign new_n14225 = new_n3972 & new_n5419;
  assign new_n14226 = new_n14225 ^ new_n14224;
  assign new_n14227 = n101 & new_n5418;
  assign new_n14228 = n99 & new_n5648;
  assign new_n14229 = new_n14228 ^ new_n14227;
  assign new_n14230 = new_n14229 ^ new_n14226;
  assign new_n14231 = new_n14230 ^ n48;
  assign new_n14232 = ~new_n6110 & n97;
  assign new_n14233 = new_n3435 & new_n6105;
  assign new_n14234 = new_n14233 ^ new_n14232;
  assign new_n14235 = n98 & new_n6104;
  assign new_n14236 = n96 & new_n6347;
  assign new_n14237 = new_n14236 ^ new_n14235;
  assign new_n14238 = new_n14237 ^ new_n14234;
  assign new_n14239 = new_n14238 ^ n51;
  assign new_n14240 = ~new_n6805 & n94;
  assign new_n14241 = new_n2934 & new_n6800;
  assign new_n14242 = new_n14241 ^ new_n14240;
  assign new_n14243 = n95 & new_n6799;
  assign new_n14244 = n93 & new_n6811;
  assign new_n14245 = new_n14244 ^ new_n14243;
  assign new_n14246 = new_n14245 ^ new_n14242;
  assign new_n14247 = new_n14246 ^ n54;
  assign new_n14248 = n88 & new_n8355;
  assign new_n14249 = new_n2063 & new_n8345;
  assign new_n14250 = new_n14249 ^ new_n14248;
  assign new_n14251 = n89 & new_n8344;
  assign new_n14252 = n87 & new_n8349;
  assign new_n14253 = new_n14252 ^ new_n14251;
  assign new_n14254 = new_n14253 ^ new_n14250;
  assign new_n14255 = new_n14254 ^ n60;
  assign new_n14256 = new_n14071 ^ new_n14048;
  assign new_n14257 = new_n14072 & new_n14256;
  assign new_n14258 = new_n14257 ^ new_n14048;
  assign new_n14259 = new_n14258 ^ new_n14255;
  assign new_n14260 = new_n14055 ^ n82;
  assign new_n14261 = ~new_n1087 & ~new_n14055;
  assign new_n14262 = new_n14055 ^ new_n1087;
  assign new_n14263 = new_n14262 ^ new_n14261;
  assign new_n14264 = ~n64 & new_n1087;
  assign new_n14265 = new_n14264 ^ new_n14263;
  assign new_n14266 = ~new_n14260 & ~new_n14265;
  assign new_n14267 = new_n995 & new_n14055;
  assign new_n14268 = n81 & new_n995;
  assign new_n14269 = new_n14268 ^ new_n14267;
  assign new_n14270 = new_n14269 ^ new_n1087;
  assign new_n14271 = new_n14261 ^ new_n11491;
  assign new_n14272 = new_n14270 & new_n14271;
  assign new_n14273 = n81 & new_n1087;
  assign new_n14274 = ~new_n14055 & ~new_n14273;
  assign new_n14275 = new_n14274 ^ n63;
  assign new_n14276 = new_n14267 ^ new_n14263;
  assign new_n14277 = new_n14273 ^ new_n14268;
  assign new_n14278 = new_n14277 ^ new_n14276;
  assign new_n14279 = new_n14275 & new_n14278;
  assign new_n14280 = new_n14279 ^ new_n14272;
  assign new_n14281 = new_n14280 ^ new_n14266;
  assign new_n14282 = n85 & new_n9195;
  assign new_n14283 = new_n1694 & new_n9185;
  assign new_n14284 = new_n14283 ^ new_n14282;
  assign new_n14285 = n86 & new_n9184;
  assign new_n14286 = n84 & new_n9189;
  assign new_n14287 = new_n14286 ^ new_n14285;
  assign new_n14288 = new_n14287 ^ new_n14284;
  assign new_n14289 = new_n14288 ^ n63;
  assign new_n14290 = new_n14264 ^ new_n1087;
  assign new_n14291 = new_n14290 ^ new_n1178;
  assign new_n14292 = ~new_n9495 & new_n14291;
  assign new_n14293 = new_n14292 ^ new_n1178;
  assign new_n14294 = new_n14293 ^ n18;
  assign new_n14295 = new_n14294 ^ new_n14289;
  assign new_n14296 = new_n14295 ^ new_n14281;
  assign new_n14297 = new_n14296 ^ new_n14259;
  assign new_n14298 = n91 & new_n7553;
  assign new_n14299 = new_n2481 & new_n7543;
  assign new_n14300 = new_n14299 ^ new_n14298;
  assign new_n14301 = n92 & new_n7542;
  assign new_n14302 = n90 & new_n7547;
  assign new_n14303 = new_n14302 ^ new_n14301;
  assign new_n14304 = new_n14303 ^ new_n14300;
  assign new_n14305 = new_n14304 ^ n57;
  assign new_n14306 = new_n14305 ^ new_n14297;
  assign new_n14307 = new_n14076 ^ new_n14040;
  assign new_n14308 = new_n14077 & new_n14307;
  assign new_n14309 = new_n14308 ^ new_n14040;
  assign new_n14310 = new_n14309 ^ new_n14306;
  assign new_n14311 = new_n14310 ^ new_n14247;
  assign new_n14312 = new_n14082 ^ new_n14078;
  assign new_n14313 = ~new_n14079 & new_n14312;
  assign new_n14314 = new_n14313 ^ new_n14032;
  assign new_n14315 = new_n14314 ^ new_n14311;
  assign new_n14316 = new_n14315 ^ new_n14239;
  assign new_n14317 = new_n14087 ^ new_n14083;
  assign new_n14318 = ~new_n14084 & new_n14317;
  assign new_n14319 = new_n14318 ^ new_n14024;
  assign new_n14320 = new_n14319 ^ new_n14316;
  assign new_n14321 = new_n14320 ^ new_n14231;
  assign new_n14322 = new_n14088 ^ new_n14015;
  assign new_n14323 = new_n14016 & new_n14322;
  assign new_n14324 = new_n14323 ^ new_n14012;
  assign new_n14325 = new_n14324 ^ new_n14321;
  assign new_n14326 = new_n14325 ^ new_n14223;
  assign new_n14327 = new_n14093 ^ new_n14089;
  assign new_n14328 = ~new_n14090 & new_n14327;
  assign new_n14329 = new_n14328 ^ new_n14004;
  assign new_n14330 = new_n14329 ^ new_n14326;
  assign new_n14331 = new_n14330 ^ new_n14215;
  assign new_n14332 = new_n14097 ^ new_n13996;
  assign new_n14333 = new_n14098 & new_n14332;
  assign new_n14334 = new_n14333 ^ new_n13996;
  assign new_n14335 = new_n14334 ^ new_n14331;
  assign new_n14336 = new_n14335 ^ new_n14207;
  assign new_n14337 = new_n14099 ^ new_n13988;
  assign new_n14338 = ~new_n14337 & new_n14103;
  assign new_n14339 = new_n14338 ^ new_n13988;
  assign new_n14340 = new_n14339 ^ new_n14336;
  assign new_n14341 = new_n14340 ^ new_n14199;
  assign new_n14342 = new_n14107 ^ new_n13980;
  assign new_n14343 = new_n14108 & new_n14342;
  assign new_n14344 = new_n14343 ^ new_n13980;
  assign new_n14345 = new_n14344 ^ new_n14341;
  assign new_n14346 = new_n14345 ^ new_n14191;
  assign new_n14347 = new_n14109 ^ new_n13972;
  assign new_n14348 = ~new_n14347 & new_n14113;
  assign new_n14349 = new_n14348 ^ new_n13972;
  assign new_n14350 = new_n14349 ^ new_n14346;
  assign new_n14351 = new_n14350 ^ new_n14183;
  assign new_n14352 = new_n14114 ^ new_n13964;
  assign new_n14353 = ~new_n14352 & new_n14118;
  assign new_n14354 = new_n14353 ^ new_n13964;
  assign new_n14355 = new_n14354 ^ new_n14351;
  assign new_n14356 = new_n14119 ^ new_n13956;
  assign new_n14357 = ~new_n14356 & new_n14123;
  assign new_n14358 = new_n14357 ^ new_n13956;
  assign new_n14359 = new_n14358 ^ new_n14355;
  assign new_n14360 = n121 & new_n1874;
  assign new_n14361 = new_n1864 & new_n8850;
  assign new_n14362 = new_n14361 ^ new_n14360;
  assign new_n14363 = n122 & new_n1863;
  assign new_n14364 = n120 & new_n1868;
  assign new_n14365 = new_n14364 ^ new_n14363;
  assign new_n14366 = new_n14365 ^ new_n14362;
  assign new_n14367 = new_n14366 ^ n27;
  assign new_n14368 = new_n14367 ^ new_n14359;
  assign new_n14369 = new_n14368 ^ new_n14175;
  assign new_n14370 = new_n14127 ^ new_n13948;
  assign new_n14371 = new_n14128 & new_n14370;
  assign new_n14372 = new_n14371 ^ new_n13948;
  assign new_n14373 = new_n14372 ^ new_n14369;
  assign new_n14374 = new_n14373 ^ new_n14167;
  assign new_n14375 = new_n14132 ^ new_n13940;
  assign new_n14376 = new_n14133 & new_n14375;
  assign new_n14377 = new_n14376 ^ new_n13940;
  assign new_n14378 = new_n14377 ^ new_n14374;
  assign new_n14379 = new_n14145 ^ new_n14141;
  assign new_n14380 = new_n14142 & new_n14379;
  assign new_n14381 = new_n14380 ^ new_n14145;
  assign new_n14382 = new_n14381 ^ new_n14378;
  assign new_n14383 = new_n14382 ^ new_n14159;
  assign new_n14384 = new_n14374 ^ new_n14159;
  assign new_n14385 = new_n14381 ^ new_n14377;
  assign new_n14386 = new_n14385 ^ new_n14159;
  assign new_n14387 = ~new_n14384 & new_n14386;
  assign new_n14388 = new_n14377 & new_n14381;
  assign new_n14389 = new_n14388 ^ new_n14387;
  assign new_n14390 = ~new_n14167 & ~new_n14373;
  assign new_n14391 = new_n14390 ^ new_n14389;
  assign new_n14392 = ~new_n1506 & n125;
  assign new_n14393 = new_n1501 & new_n9987;
  assign new_n14394 = new_n14393 ^ new_n14392;
  assign new_n14395 = n126 & new_n1500;
  assign new_n14396 = n124 & new_n1512;
  assign new_n14397 = new_n14396 ^ new_n14395;
  assign new_n14398 = new_n14397 ^ new_n14394;
  assign new_n14399 = new_n14398 ^ n24;
  assign new_n14400 = n122 & new_n1874;
  assign new_n14401 = ~new_n9116 & new_n1864;
  assign new_n14402 = new_n14401 ^ new_n14400;
  assign new_n14403 = n123 & new_n1863;
  assign new_n14404 = n121 & new_n1868;
  assign new_n14405 = new_n14404 ^ new_n14403;
  assign new_n14406 = new_n14405 ^ new_n14402;
  assign new_n14407 = new_n14406 ^ n27;
  assign new_n14408 = n119 & new_n2246;
  assign new_n14409 = new_n2241 & new_n8286;
  assign new_n14410 = new_n14409 ^ new_n14408;
  assign new_n14411 = n120 & new_n2240;
  assign new_n14412 = n118 & new_n2391;
  assign new_n14413 = new_n14412 ^ new_n14411;
  assign new_n14414 = new_n14413 ^ new_n14410;
  assign new_n14415 = new_n14414 ^ n30;
  assign new_n14416 = ~new_n2672 & n116;
  assign new_n14417 = ~new_n7503 & new_n2667;
  assign new_n14418 = new_n14417 ^ new_n14416;
  assign new_n14419 = n117 & new_n2666;
  assign new_n14420 = n115 & new_n2664;
  assign new_n14421 = new_n14420 ^ new_n14419;
  assign new_n14422 = new_n14421 ^ new_n14418;
  assign new_n14423 = new_n14422 ^ n33;
  assign new_n14424 = ~new_n3143 & n113;
  assign new_n14425 = ~new_n6764 & new_n3138;
  assign new_n14426 = new_n14425 ^ new_n14424;
  assign new_n14427 = n114 & new_n3137;
  assign new_n14428 = n112 & new_n3149;
  assign new_n14429 = new_n14428 ^ new_n14427;
  assign new_n14430 = new_n14429 ^ new_n14426;
  assign new_n14431 = new_n14430 ^ n36;
  assign new_n14432 = ~new_n5424 & n101;
  assign new_n14433 = new_n4159 & new_n5419;
  assign new_n14434 = new_n14433 ^ new_n14432;
  assign new_n14435 = n102 & new_n5418;
  assign new_n14436 = n100 & new_n5648;
  assign new_n14437 = new_n14436 ^ new_n14435;
  assign new_n14438 = new_n14437 ^ new_n14434;
  assign new_n14439 = new_n14438 ^ n48;
  assign new_n14440 = ~new_n6110 & n98;
  assign new_n14441 = new_n3604 & new_n6105;
  assign new_n14442 = new_n14441 ^ new_n14440;
  assign new_n14443 = n99 & new_n6104;
  assign new_n14444 = n97 & new_n6347;
  assign new_n14445 = new_n14444 ^ new_n14443;
  assign new_n14446 = new_n14445 ^ new_n14442;
  assign new_n14447 = new_n14446 ^ n51;
  assign new_n14448 = ~new_n6805 & n95;
  assign new_n14449 = new_n3095 & new_n6800;
  assign new_n14450 = new_n14449 ^ new_n14448;
  assign new_n14451 = n96 & new_n6799;
  assign new_n14452 = n94 & new_n6811;
  assign new_n14453 = new_n14452 ^ new_n14451;
  assign new_n14454 = new_n14453 ^ new_n14450;
  assign new_n14455 = new_n14454 ^ n54;
  assign new_n14456 = n92 & new_n7553;
  assign new_n14457 = new_n2628 & new_n7543;
  assign new_n14458 = new_n14457 ^ new_n14456;
  assign new_n14459 = n93 & new_n7542;
  assign new_n14460 = n91 & new_n7547;
  assign new_n14461 = new_n14460 ^ new_n14459;
  assign new_n14462 = new_n14461 ^ new_n14458;
  assign new_n14463 = new_n14462 ^ n57;
  assign new_n14464 = new_n14296 ^ new_n14255;
  assign new_n14465 = ~new_n14464 & new_n14259;
  assign new_n14466 = new_n14465 ^ new_n14258;
  assign new_n14467 = new_n14466 ^ new_n14463;
  assign new_n14468 = n89 & new_n8355;
  assign new_n14469 = new_n2193 & new_n8345;
  assign new_n14470 = new_n14469 ^ new_n14468;
  assign new_n14471 = n88 & new_n8349;
  assign new_n14472 = n90 & new_n8344;
  assign new_n14473 = new_n14472 ^ new_n14471;
  assign new_n14474 = new_n14473 ^ new_n14470;
  assign new_n14475 = new_n14474 ^ n60;
  assign new_n14476 = n86 & new_n9195;
  assign new_n14477 = new_n1811 & new_n9185;
  assign new_n14478 = new_n14477 ^ new_n14476;
  assign new_n14479 = n87 & new_n9184;
  assign new_n14480 = n85 & new_n9189;
  assign new_n14481 = new_n14480 ^ new_n14479;
  assign new_n14482 = new_n14481 ^ new_n14478;
  assign new_n14483 = new_n14482 ^ n63;
  assign new_n14484 = n83 & new_n11492;
  assign new_n14485 = n84 & new_n9495;
  assign new_n14486 = new_n14485 ^ new_n14484;
  assign new_n14487 = n82 ^ n18;
  assign new_n14488 = n83 ^ n81;
  assign new_n14489 = new_n11492 & new_n14488;
  assign new_n14490 = new_n14489 ^ n83;
  assign new_n14491 = new_n14490 ^ n82;
  assign new_n14492 = ~new_n14487 & new_n14491;
  assign new_n14493 = new_n14492 ^ n82;
  assign new_n14494 = new_n11789 & new_n14493;
  assign new_n14495 = new_n14494 ^ new_n14486;
  assign new_n14496 = new_n14495 ^ new_n14483;
  assign new_n14497 = new_n14496 ^ new_n14475;
  assign new_n14498 = new_n14289 ^ new_n14281;
  assign new_n14499 = ~new_n14498 & new_n14295;
  assign new_n14500 = new_n14499 ^ new_n14281;
  assign new_n14501 = new_n14500 ^ new_n14497;
  assign new_n14502 = new_n14501 ^ new_n14467;
  assign new_n14503 = new_n14309 ^ new_n14305;
  assign new_n14504 = ~new_n14503 & new_n14306;
  assign new_n14505 = new_n14504 ^ new_n14297;
  assign new_n14506 = new_n14505 ^ new_n14502;
  assign new_n14507 = new_n14506 ^ new_n14455;
  assign new_n14508 = new_n14314 ^ new_n14247;
  assign new_n14509 = ~new_n14311 & new_n14508;
  assign new_n14510 = new_n14509 ^ new_n14314;
  assign new_n14511 = new_n14510 ^ new_n14507;
  assign new_n14512 = new_n14511 ^ new_n14447;
  assign new_n14513 = new_n14319 ^ new_n14239;
  assign new_n14514 = ~new_n14316 & new_n14513;
  assign new_n14515 = new_n14514 ^ new_n14319;
  assign new_n14516 = new_n14515 ^ new_n14512;
  assign new_n14517 = new_n14516 ^ new_n14439;
  assign new_n14518 = new_n14324 ^ new_n14231;
  assign new_n14519 = ~new_n14321 & new_n14518;
  assign new_n14520 = new_n14519 ^ new_n14324;
  assign new_n14521 = new_n14520 ^ new_n14517;
  assign new_n14522 = ~new_n4804 & n104;
  assign new_n14523 = ~new_n4754 & new_n4799;
  assign new_n14524 = new_n14523 ^ new_n14522;
  assign new_n14525 = n105 & new_n4798;
  assign new_n14526 = n103 & new_n4810;
  assign new_n14527 = new_n14526 ^ new_n14525;
  assign new_n14528 = new_n14527 ^ new_n14524;
  assign new_n14529 = new_n14528 ^ n45;
  assign new_n14530 = new_n14529 ^ new_n14521;
  assign new_n14531 = new_n14329 ^ new_n14223;
  assign new_n14532 = ~new_n14326 & new_n14531;
  assign new_n14533 = new_n14532 ^ new_n14329;
  assign new_n14534 = new_n14533 ^ new_n14530;
  assign new_n14535 = ~new_n4212 & n107;
  assign new_n14536 = ~new_n5377 & new_n4201;
  assign new_n14537 = new_n14536 ^ new_n14535;
  assign new_n14538 = n108 & new_n4200;
  assign new_n14539 = n106 & new_n4206;
  assign new_n14540 = new_n14539 ^ new_n14538;
  assign new_n14541 = new_n14540 ^ new_n14537;
  assign new_n14542 = new_n14541 ^ n42;
  assign new_n14543 = new_n14542 ^ new_n14534;
  assign new_n14544 = new_n14334 ^ new_n14215;
  assign new_n14545 = ~new_n14331 & new_n14544;
  assign new_n14546 = new_n14545 ^ new_n14334;
  assign new_n14547 = new_n14546 ^ new_n14543;
  assign new_n14548 = ~new_n3682 & n110;
  assign new_n14549 = new_n3677 & new_n6049;
  assign new_n14550 = new_n14549 ^ new_n14548;
  assign new_n14551 = n111 & new_n3676;
  assign new_n14552 = n109 & new_n3688;
  assign new_n14553 = new_n14552 ^ new_n14551;
  assign new_n14554 = new_n14553 ^ new_n14550;
  assign new_n14555 = new_n14554 ^ n39;
  assign new_n14556 = new_n14555 ^ new_n14547;
  assign new_n14557 = new_n14339 ^ new_n14207;
  assign new_n14558 = ~new_n14336 & new_n14557;
  assign new_n14559 = new_n14558 ^ new_n14339;
  assign new_n14560 = new_n14559 ^ new_n14556;
  assign new_n14561 = new_n14560 ^ new_n14431;
  assign new_n14562 = new_n14344 ^ new_n14340;
  assign new_n14563 = ~new_n14562 & new_n14341;
  assign new_n14564 = new_n14563 ^ new_n14199;
  assign new_n14565 = new_n14564 ^ new_n14561;
  assign new_n14566 = new_n14565 ^ new_n14423;
  assign new_n14567 = new_n14566 ^ new_n14415;
  assign new_n14568 = new_n14349 ^ new_n14191;
  assign new_n14569 = ~new_n14346 & new_n14568;
  assign new_n14570 = new_n14569 ^ new_n14349;
  assign new_n14571 = new_n14570 ^ new_n14567;
  assign new_n14572 = new_n14354 ^ new_n14183;
  assign new_n14573 = ~new_n14351 & new_n14572;
  assign new_n14574 = new_n14573 ^ new_n14354;
  assign new_n14575 = new_n14574 ^ new_n14571;
  assign new_n14576 = new_n14575 ^ new_n14407;
  assign new_n14577 = new_n14367 ^ new_n14355;
  assign new_n14578 = ~new_n14577 & new_n14359;
  assign new_n14579 = new_n14578 ^ new_n14358;
  assign new_n14580 = new_n14579 ^ new_n14576;
  assign new_n14581 = new_n14580 ^ new_n14399;
  assign new_n14582 = new_n14372 ^ new_n14175;
  assign new_n14583 = ~new_n14369 & new_n14582;
  assign new_n14584 = new_n14583 ^ new_n14372;
  assign new_n14585 = new_n14584 ^ new_n14581;
  assign new_n14586 = n127 & new_n1204;
  assign new_n14587 = new_n1193 & new_n10010;
  assign new_n14588 = new_n14587 ^ new_n14586;
  assign new_n14589 = ~new_n1198 & n128;
  assign new_n14590 = new_n14589 ^ new_n14588;
  assign new_n14591 = new_n14590 ^ n21;
  assign new_n14592 = new_n14591 ^ new_n14585;
  assign new_n14593 = new_n14592 ^ new_n14391;
  assign new_n14594 = new_n14388 ^ new_n14385;
  assign new_n14595 = new_n14390 ^ new_n14374;
  assign new_n14596 = ~new_n14595 & new_n14594;
  assign new_n14597 = ~new_n14592 & ~new_n14596;
  assign new_n14598 = ~new_n14159 & ~new_n14597;
  assign new_n14599 = ~new_n14390 & new_n14592;
  assign new_n14600 = ~new_n14388 & ~new_n14599;
  assign new_n14601 = ~new_n14598 & new_n14600;
  assign new_n14602 = new_n14592 & new_n14594;
  assign new_n14603 = new_n14167 ^ new_n14159;
  assign new_n14604 = ~new_n14603 & new_n14374;
  assign new_n14605 = new_n14604 ^ new_n14167;
  assign new_n14606 = ~new_n14602 & ~new_n14605;
  assign new_n14607 = ~new_n14601 & ~new_n14606;
  assign new_n14608 = ~new_n1506 & n126;
  assign new_n14609 = new_n1501 & new_n10304;
  assign new_n14610 = new_n14609 ^ new_n14608;
  assign new_n14611 = n127 & new_n1500;
  assign new_n14612 = n125 & new_n1512;
  assign new_n14613 = new_n14612 ^ new_n14611;
  assign new_n14614 = new_n14613 ^ new_n14610;
  assign new_n14615 = new_n14614 ^ n24;
  assign new_n14616 = n123 & new_n1874;
  assign new_n14617 = ~new_n9405 & new_n1864;
  assign new_n14618 = new_n14617 ^ new_n14616;
  assign new_n14619 = n124 & new_n1863;
  assign new_n14620 = n122 & new_n1868;
  assign new_n14621 = new_n14620 ^ new_n14619;
  assign new_n14622 = new_n14621 ^ new_n14618;
  assign new_n14623 = new_n14622 ^ n27;
  assign new_n14624 = n120 & new_n2246;
  assign new_n14625 = new_n2241 & new_n8560;
  assign new_n14626 = new_n14625 ^ new_n14624;
  assign new_n14627 = n121 & new_n2240;
  assign new_n14628 = n119 & new_n2391;
  assign new_n14629 = new_n14628 ^ new_n14627;
  assign new_n14630 = new_n14629 ^ new_n14626;
  assign new_n14631 = new_n14630 ^ n30;
  assign new_n14632 = ~new_n2672 & n117;
  assign new_n14633 = ~new_n7761 & new_n2667;
  assign new_n14634 = new_n14633 ^ new_n14632;
  assign new_n14635 = n118 & new_n2666;
  assign new_n14636 = n116 & new_n2664;
  assign new_n14637 = new_n14636 ^ new_n14635;
  assign new_n14638 = new_n14637 ^ new_n14634;
  assign new_n14639 = new_n14638 ^ n33;
  assign new_n14640 = ~new_n3143 & n114;
  assign new_n14641 = ~new_n7013 & new_n3138;
  assign new_n14642 = new_n14641 ^ new_n14640;
  assign new_n14643 = n115 & new_n3137;
  assign new_n14644 = n113 & new_n3149;
  assign new_n14645 = new_n14644 ^ new_n14643;
  assign new_n14646 = new_n14645 ^ new_n14642;
  assign new_n14647 = new_n14646 ^ n36;
  assign new_n14648 = ~new_n3682 & n111;
  assign new_n14649 = ~new_n6284 & new_n3677;
  assign new_n14650 = new_n14649 ^ new_n14648;
  assign new_n14651 = n112 & new_n3676;
  assign new_n14652 = n110 & new_n3688;
  assign new_n14653 = new_n14652 ^ new_n14651;
  assign new_n14654 = new_n14653 ^ new_n14650;
  assign new_n14655 = new_n14654 ^ n39;
  assign new_n14656 = ~new_n4212 & n108;
  assign new_n14657 = new_n4201 & new_n5604;
  assign new_n14658 = new_n14657 ^ new_n14656;
  assign new_n14659 = n109 & new_n4200;
  assign new_n14660 = n107 & new_n4206;
  assign new_n14661 = new_n14660 ^ new_n14659;
  assign new_n14662 = new_n14661 ^ new_n14658;
  assign new_n14663 = new_n14662 ^ n42;
  assign new_n14664 = ~new_n4804 & n105;
  assign new_n14665 = ~new_n4961 & new_n4799;
  assign new_n14666 = new_n14665 ^ new_n14664;
  assign new_n14667 = n106 & new_n4798;
  assign new_n14668 = n104 & new_n4810;
  assign new_n14669 = new_n14668 ^ new_n14667;
  assign new_n14670 = new_n14669 ^ new_n14666;
  assign new_n14671 = new_n14670 ^ n45;
  assign new_n14672 = ~new_n6110 & n99;
  assign new_n14673 = new_n3789 & new_n6105;
  assign new_n14674 = new_n14673 ^ new_n14672;
  assign new_n14675 = n100 & new_n6104;
  assign new_n14676 = n98 & new_n6347;
  assign new_n14677 = new_n14676 ^ new_n14675;
  assign new_n14678 = new_n14677 ^ new_n14674;
  assign new_n14679 = new_n14678 ^ n51;
  assign new_n14680 = new_n14505 ^ new_n14455;
  assign new_n14681 = ~new_n14506 & new_n14680;
  assign new_n14682 = new_n14681 ^ new_n14455;
  assign new_n14683 = new_n14682 ^ new_n14679;
  assign new_n14684 = ~new_n6805 & n96;
  assign new_n14685 = new_n3273 & new_n6800;
  assign new_n14686 = new_n14685 ^ new_n14684;
  assign new_n14687 = n97 & new_n6799;
  assign new_n14688 = n95 & new_n6811;
  assign new_n14689 = new_n14688 ^ new_n14687;
  assign new_n14690 = new_n14689 ^ new_n14686;
  assign new_n14691 = new_n14690 ^ n54;
  assign new_n14692 = n93 & new_n7553;
  assign new_n14693 = new_n2785 & new_n7543;
  assign new_n14694 = new_n14693 ^ new_n14692;
  assign new_n14695 = n94 & new_n7542;
  assign new_n14696 = n92 & new_n7547;
  assign new_n14697 = new_n14696 ^ new_n14695;
  assign new_n14698 = new_n14697 ^ new_n14694;
  assign new_n14699 = new_n14698 ^ n57;
  assign new_n14700 = new_n14500 ^ new_n14496;
  assign new_n14701 = ~new_n14497 & ~new_n14700;
  assign new_n14702 = new_n14701 ^ new_n14475;
  assign new_n14703 = new_n14702 ^ new_n14699;
  assign new_n14704 = n90 & new_n8355;
  assign new_n14705 = new_n2341 & new_n8345;
  assign new_n14706 = new_n14705 ^ new_n14704;
  assign new_n14707 = n91 & new_n8344;
  assign new_n14708 = n89 & new_n8349;
  assign new_n14709 = new_n14708 ^ new_n14707;
  assign new_n14710 = new_n14709 ^ new_n14706;
  assign new_n14711 = new_n14710 ^ n60;
  assign new_n14712 = n87 & new_n9195;
  assign new_n14713 = new_n1940 & new_n9185;
  assign new_n14714 = new_n14713 ^ new_n14712;
  assign new_n14715 = n88 & new_n9184;
  assign new_n14716 = n86 & new_n9189;
  assign new_n14717 = new_n14716 ^ new_n14715;
  assign new_n14718 = new_n14717 ^ new_n14714;
  assign new_n14719 = new_n14718 ^ n63;
  assign new_n14720 = n84 & new_n11789;
  assign new_n14721 = ~n85 & new_n9495;
  assign new_n14722 = new_n14721 ^ new_n14484;
  assign new_n14723 = new_n14722 ^ new_n9495;
  assign new_n14724 = new_n14723 ^ new_n14720;
  assign new_n14725 = new_n14724 ^ new_n14719;
  assign new_n14726 = new_n14494 ^ new_n14483;
  assign new_n14727 = new_n14495 & new_n14726;
  assign new_n14728 = new_n14727 ^ new_n14483;
  assign new_n14729 = new_n14728 ^ new_n14725;
  assign new_n14730 = new_n14729 ^ new_n14711;
  assign new_n14731 = new_n14730 ^ new_n14703;
  assign new_n14732 = new_n14731 ^ new_n14691;
  assign new_n14733 = new_n14501 ^ new_n14463;
  assign new_n14734 = ~new_n14733 & new_n14467;
  assign new_n14735 = new_n14734 ^ new_n14466;
  assign new_n14736 = new_n14735 ^ new_n14732;
  assign new_n14737 = new_n14736 ^ new_n14683;
  assign new_n14738 = new_n14510 ^ new_n14447;
  assign new_n14739 = ~new_n14511 & new_n14738;
  assign new_n14740 = new_n14739 ^ new_n14447;
  assign new_n14741 = new_n14740 ^ new_n14737;
  assign new_n14742 = ~new_n5424 & n102;
  assign new_n14743 = new_n4368 & new_n5419;
  assign new_n14744 = new_n14743 ^ new_n14742;
  assign new_n14745 = n103 & new_n5418;
  assign new_n14746 = n101 & new_n5648;
  assign new_n14747 = new_n14746 ^ new_n14745;
  assign new_n14748 = new_n14747 ^ new_n14744;
  assign new_n14749 = new_n14748 ^ n48;
  assign new_n14750 = new_n14749 ^ new_n14741;
  assign new_n14751 = new_n14515 ^ new_n14439;
  assign new_n14752 = ~new_n14516 & new_n14751;
  assign new_n14753 = new_n14752 ^ new_n14439;
  assign new_n14754 = new_n14753 ^ new_n14750;
  assign new_n14755 = new_n14754 ^ new_n14671;
  assign new_n14756 = new_n14529 ^ new_n14517;
  assign new_n14757 = ~new_n14756 & new_n14521;
  assign new_n14758 = new_n14757 ^ new_n14520;
  assign new_n14759 = new_n14758 ^ new_n14755;
  assign new_n14760 = new_n14759 ^ new_n14663;
  assign new_n14761 = new_n14542 ^ new_n14530;
  assign new_n14762 = ~new_n14761 & new_n14534;
  assign new_n14763 = new_n14762 ^ new_n14533;
  assign new_n14764 = new_n14763 ^ new_n14760;
  assign new_n14765 = new_n14764 ^ new_n14655;
  assign new_n14766 = new_n14555 ^ new_n14543;
  assign new_n14767 = ~new_n14766 & new_n14547;
  assign new_n14768 = new_n14767 ^ new_n14546;
  assign new_n14769 = new_n14768 ^ new_n14765;
  assign new_n14770 = new_n14769 ^ new_n14647;
  assign new_n14771 = new_n14556 ^ new_n14431;
  assign new_n14772 = ~new_n14560 & new_n14771;
  assign new_n14773 = new_n14772 ^ new_n14431;
  assign new_n14774 = new_n14773 ^ new_n14770;
  assign new_n14775 = new_n14774 ^ new_n14639;
  assign new_n14776 = new_n14564 ^ new_n14423;
  assign new_n14777 = ~new_n14565 & new_n14776;
  assign new_n14778 = new_n14777 ^ new_n14423;
  assign new_n14779 = new_n14778 ^ new_n14775;
  assign new_n14780 = new_n14779 ^ new_n14631;
  assign new_n14781 = new_n14570 ^ new_n14566;
  assign new_n14782 = ~new_n14781 & new_n14567;
  assign new_n14783 = new_n14782 ^ new_n14415;
  assign new_n14784 = new_n14783 ^ new_n14780;
  assign new_n14785 = new_n14784 ^ new_n14623;
  assign new_n14786 = new_n14574 ^ new_n14407;
  assign new_n14787 = ~new_n14575 & new_n14786;
  assign new_n14788 = new_n14787 ^ new_n14407;
  assign new_n14789 = new_n14788 ^ new_n14785;
  assign new_n14790 = new_n14789 ^ new_n14615;
  assign new_n14791 = new_n14591 ^ new_n14581;
  assign new_n14792 = ~new_n14791 & new_n14585;
  assign new_n14793 = new_n14792 ^ new_n14584;
  assign new_n14794 = new_n14793 ^ new_n14790;
  assign new_n14795 = ~new_n1203 & n128;
  assign new_n14796 = ~n21 & ~new_n14795;
  assign new_n14797 = new_n14796 ^ n20;
  assign new_n14798 = new_n1025 & new_n11133;
  assign new_n14799 = new_n14798 ^ new_n14795;
  assign new_n14800 = ~new_n14797 & ~new_n14799;
  assign new_n14801 = new_n14800 ^ n20;
  assign new_n14802 = new_n14576 ^ new_n14399;
  assign new_n14803 = ~new_n14580 & new_n14802;
  assign new_n14804 = new_n14803 ^ new_n14399;
  assign new_n14805 = new_n14804 ^ new_n14801;
  assign new_n14806 = new_n14805 ^ new_n14794;
  assign new_n14807 = new_n14806 ^ new_n14607;
  assign new_n14808 = ~new_n14793 & new_n14790;
  assign new_n14809 = new_n14808 ^ new_n14794;
  assign new_n14810 = ~new_n14801 & ~new_n14804;
  assign new_n14811 = new_n14810 ^ new_n14805;
  assign new_n14812 = new_n14809 & new_n14811;
  assign new_n14813 = new_n14808 ^ new_n14607;
  assign new_n14814 = new_n14811 ^ new_n14808;
  assign new_n14815 = new_n14813 & new_n14814;
  assign new_n14816 = new_n14815 ^ new_n14812;
  assign new_n14817 = ~new_n14810 & new_n14808;
  assign new_n14818 = new_n14809 ^ new_n14607;
  assign new_n14819 = new_n14810 ^ new_n14809;
  assign new_n14820 = ~new_n14818 & ~new_n14819;
  assign new_n14821 = new_n14820 ^ new_n14817;
  assign new_n14822 = new_n14821 ^ new_n14816;
  assign new_n14823 = ~new_n1506 & n127;
  assign new_n14824 = new_n1501 & new_n10581;
  assign new_n14825 = new_n14824 ^ new_n14823;
  assign new_n14826 = n128 & new_n1500;
  assign new_n14827 = n126 & new_n1512;
  assign new_n14828 = new_n14827 ^ new_n14826;
  assign new_n14829 = new_n14828 ^ new_n14825;
  assign new_n14830 = new_n14829 ^ n24;
  assign new_n14831 = n124 & new_n1874;
  assign new_n14832 = new_n1864 & new_n9700;
  assign new_n14833 = new_n14832 ^ new_n14831;
  assign new_n14834 = n125 & new_n1863;
  assign new_n14835 = n123 & new_n1868;
  assign new_n14836 = new_n14835 ^ new_n14834;
  assign new_n14837 = new_n14836 ^ new_n14833;
  assign new_n14838 = new_n14837 ^ n27;
  assign new_n14839 = ~new_n2672 & n118;
  assign new_n14840 = ~new_n8019 & new_n2667;
  assign new_n14841 = new_n14840 ^ new_n14839;
  assign new_n14842 = n119 & new_n2666;
  assign new_n14843 = n117 & new_n2664;
  assign new_n14844 = new_n14843 ^ new_n14842;
  assign new_n14845 = new_n14844 ^ new_n14841;
  assign new_n14846 = new_n14845 ^ n33;
  assign new_n14847 = ~new_n3143 & n115;
  assign new_n14848 = ~new_n7256 & new_n3138;
  assign new_n14849 = new_n14848 ^ new_n14847;
  assign new_n14850 = n116 & new_n3137;
  assign new_n14851 = n114 & new_n3149;
  assign new_n14852 = new_n14851 ^ new_n14850;
  assign new_n14853 = new_n14852 ^ new_n14849;
  assign new_n14854 = new_n14853 ^ n36;
  assign new_n14855 = ~new_n3682 & n112;
  assign new_n14856 = ~new_n6518 & new_n3677;
  assign new_n14857 = new_n14856 ^ new_n14855;
  assign new_n14858 = n113 & new_n3676;
  assign new_n14859 = n111 & new_n3688;
  assign new_n14860 = new_n14859 ^ new_n14858;
  assign new_n14861 = new_n14860 ^ new_n14857;
  assign new_n14862 = new_n14861 ^ n39;
  assign new_n14863 = ~new_n4212 & n109;
  assign new_n14864 = new_n4201 & new_n5825;
  assign new_n14865 = new_n14864 ^ new_n14863;
  assign new_n14866 = n110 & new_n4200;
  assign new_n14867 = n108 & new_n4206;
  assign new_n14868 = new_n14867 ^ new_n14866;
  assign new_n14869 = new_n14868 ^ new_n14865;
  assign new_n14870 = new_n14869 ^ n42;
  assign new_n14871 = ~new_n4804 & n106;
  assign new_n14872 = ~new_n5164 & new_n4799;
  assign new_n14873 = new_n14872 ^ new_n14871;
  assign new_n14874 = n107 & new_n4798;
  assign new_n14875 = n105 & new_n4810;
  assign new_n14876 = new_n14875 ^ new_n14874;
  assign new_n14877 = new_n14876 ^ new_n14873;
  assign new_n14878 = new_n14877 ^ n45;
  assign new_n14879 = ~new_n6110 & n100;
  assign new_n14880 = new_n3972 & new_n6105;
  assign new_n14881 = new_n14880 ^ new_n14879;
  assign new_n14882 = n101 & new_n6104;
  assign new_n14883 = n99 & new_n6347;
  assign new_n14884 = new_n14883 ^ new_n14882;
  assign new_n14885 = new_n14884 ^ new_n14881;
  assign new_n14886 = new_n14885 ^ n51;
  assign new_n14887 = new_n14736 ^ new_n14682;
  assign new_n14888 = new_n14683 & new_n14887;
  assign new_n14889 = new_n14888 ^ new_n14679;
  assign new_n14890 = new_n14889 ^ new_n14886;
  assign new_n14891 = ~new_n6805 & n97;
  assign new_n14892 = new_n3435 & new_n6800;
  assign new_n14893 = new_n14892 ^ new_n14891;
  assign new_n14894 = n98 & new_n6799;
  assign new_n14895 = n96 & new_n6811;
  assign new_n14896 = new_n14895 ^ new_n14894;
  assign new_n14897 = new_n14896 ^ new_n14893;
  assign new_n14898 = new_n14897 ^ n54;
  assign new_n14899 = n94 & new_n7553;
  assign new_n14900 = new_n2934 & new_n7543;
  assign new_n14901 = new_n14900 ^ new_n14899;
  assign new_n14902 = n95 & new_n7542;
  assign new_n14903 = n93 & new_n7547;
  assign new_n14904 = new_n14903 ^ new_n14902;
  assign new_n14905 = new_n14904 ^ new_n14901;
  assign new_n14906 = new_n14905 ^ n57;
  assign new_n14907 = n91 & new_n8355;
  assign new_n14908 = new_n2481 & new_n8345;
  assign new_n14909 = new_n14908 ^ new_n14907;
  assign new_n14910 = n92 & new_n8344;
  assign new_n14911 = n90 & new_n8349;
  assign new_n14912 = new_n14911 ^ new_n14910;
  assign new_n14913 = new_n14912 ^ new_n14909;
  assign new_n14914 = new_n14913 ^ n60;
  assign new_n14915 = new_n14728 ^ new_n14711;
  assign new_n14916 = new_n14729 & new_n14915;
  assign new_n14917 = new_n14916 ^ new_n14711;
  assign new_n14918 = new_n14917 ^ new_n14914;
  assign new_n14919 = n88 & new_n9195;
  assign new_n14920 = new_n2063 & new_n9185;
  assign new_n14921 = new_n14920 ^ new_n14919;
  assign new_n14922 = n89 & new_n9184;
  assign new_n14923 = n87 & new_n9189;
  assign new_n14924 = new_n14923 ^ new_n14922;
  assign new_n14925 = new_n14924 ^ new_n14921;
  assign new_n14926 = new_n14925 ^ n63;
  assign new_n14927 = n86 & new_n11492;
  assign new_n14928 = new_n14927 ^ new_n14485;
  assign new_n14929 = new_n14928 ^ new_n14720;
  assign new_n14930 = new_n14929 ^ n86;
  assign new_n14931 = new_n14930 ^ n85;
  assign new_n14932 = new_n11789 & new_n14931;
  assign new_n14933 = new_n14932 ^ n21;
  assign new_n14934 = new_n14933 ^ new_n14926;
  assign new_n14935 = n84 & new_n14722;
  assign new_n14936 = new_n14935 ^ new_n14484;
  assign new_n14937 = ~new_n14724 & new_n14719;
  assign new_n14938 = new_n14937 ^ new_n14936;
  assign new_n14939 = new_n14938 ^ new_n14934;
  assign new_n14940 = new_n14939 ^ new_n14918;
  assign new_n14941 = new_n14940 ^ new_n14906;
  assign new_n14942 = new_n14730 ^ new_n14702;
  assign new_n14943 = new_n14703 & new_n14942;
  assign new_n14944 = new_n14943 ^ new_n14699;
  assign new_n14945 = new_n14944 ^ new_n14941;
  assign new_n14946 = new_n14945 ^ new_n14898;
  assign new_n14947 = new_n14735 ^ new_n14731;
  assign new_n14948 = ~new_n14732 & new_n14947;
  assign new_n14949 = new_n14948 ^ new_n14691;
  assign new_n14950 = new_n14949 ^ new_n14946;
  assign new_n14951 = new_n14950 ^ new_n14890;
  assign new_n14952 = new_n14749 ^ new_n14740;
  assign new_n14953 = ~new_n14741 & ~new_n14952;
  assign new_n14954 = new_n14953 ^ new_n14737;
  assign new_n14955 = new_n14954 ^ new_n14951;
  assign new_n14956 = ~new_n5424 & n103;
  assign new_n14957 = ~new_n4556 & new_n5419;
  assign new_n14958 = new_n14957 ^ new_n14956;
  assign new_n14959 = n104 & new_n5418;
  assign new_n14960 = n102 & new_n5648;
  assign new_n14961 = new_n14960 ^ new_n14959;
  assign new_n14962 = new_n14961 ^ new_n14958;
  assign new_n14963 = new_n14962 ^ n48;
  assign new_n14964 = new_n14963 ^ new_n14955;
  assign new_n14965 = new_n14964 ^ new_n14878;
  assign new_n14966 = new_n14750 ^ new_n14671;
  assign new_n14967 = ~new_n14966 & new_n14754;
  assign new_n14968 = new_n14967 ^ new_n14671;
  assign new_n14969 = new_n14968 ^ new_n14965;
  assign new_n14970 = new_n14969 ^ new_n14870;
  assign new_n14971 = new_n14758 ^ new_n14663;
  assign new_n14972 = new_n14759 & new_n14971;
  assign new_n14973 = new_n14972 ^ new_n14663;
  assign new_n14974 = new_n14973 ^ new_n14970;
  assign new_n14975 = new_n14974 ^ new_n14862;
  assign new_n14976 = new_n14763 ^ new_n14655;
  assign new_n14977 = new_n14764 & new_n14976;
  assign new_n14978 = new_n14977 ^ new_n14655;
  assign new_n14979 = new_n14978 ^ new_n14975;
  assign new_n14980 = new_n14979 ^ new_n14854;
  assign new_n14981 = new_n14765 ^ new_n14647;
  assign new_n14982 = ~new_n14981 & new_n14769;
  assign new_n14983 = new_n14982 ^ new_n14647;
  assign new_n14984 = new_n14983 ^ new_n14980;
  assign new_n14985 = new_n14984 ^ new_n14846;
  assign new_n14986 = new_n14770 ^ new_n14639;
  assign new_n14987 = ~new_n14986 & new_n14774;
  assign new_n14988 = new_n14987 ^ new_n14639;
  assign new_n14989 = new_n14988 ^ new_n14985;
  assign new_n14990 = new_n14775 ^ new_n14631;
  assign new_n14991 = ~new_n14990 & new_n14779;
  assign new_n14992 = new_n14991 ^ new_n14631;
  assign new_n14993 = new_n14992 ^ new_n14989;
  assign new_n14994 = n121 & new_n2246;
  assign new_n14995 = new_n2241 & new_n8850;
  assign new_n14996 = new_n14995 ^ new_n14994;
  assign new_n14997 = n122 & new_n2240;
  assign new_n14998 = n120 & new_n2391;
  assign new_n14999 = new_n14998 ^ new_n14997;
  assign new_n15000 = new_n14999 ^ new_n14996;
  assign new_n15001 = new_n15000 ^ n30;
  assign new_n15002 = new_n15001 ^ new_n14993;
  assign new_n15003 = new_n15002 ^ new_n14838;
  assign new_n15004 = new_n14783 ^ new_n14623;
  assign new_n15005 = new_n14784 & new_n15004;
  assign new_n15006 = new_n15005 ^ new_n14623;
  assign new_n15007 = new_n15006 ^ new_n15003;
  assign new_n15008 = new_n15007 ^ new_n14830;
  assign new_n15009 = new_n14785 ^ new_n14615;
  assign new_n15010 = ~new_n15009 & new_n14789;
  assign new_n15011 = new_n15010 ^ new_n14615;
  assign new_n15012 = new_n15011 ^ new_n15008;
  assign new_n15013 = new_n15012 ^ new_n14822;
  assign new_n15014 = ~new_n14808 & new_n15012;
  assign new_n15015 = ~new_n15014 & new_n14811;
  assign new_n15016 = ~new_n14810 & new_n15012;
  assign new_n15017 = ~new_n14809 & ~new_n15016;
  assign new_n15018 = ~new_n15015 & ~new_n15017;
  assign new_n15019 = ~new_n14607 & ~new_n15018;
  assign new_n15020 = new_n14811 ^ new_n14790;
  assign new_n15021 = ~new_n14794 & ~new_n15020;
  assign new_n15022 = new_n15021 ^ new_n14793;
  assign new_n15023 = ~new_n15012 & ~new_n15022;
  assign new_n15024 = new_n14810 & new_n15015;
  assign new_n15025 = ~new_n15023 & ~new_n15024;
  assign new_n15026 = ~new_n15019 & new_n15025;
  assign new_n15027 = n125 & new_n1874;
  assign new_n15028 = new_n1864 & new_n9987;
  assign new_n15029 = new_n15028 ^ new_n15027;
  assign new_n15030 = n126 & new_n1863;
  assign new_n15031 = n124 & new_n1868;
  assign new_n15032 = new_n15031 ^ new_n15030;
  assign new_n15033 = new_n15032 ^ new_n15029;
  assign new_n15034 = new_n15033 ^ n27;
  assign new_n15035 = n122 & new_n2246;
  assign new_n15036 = ~new_n9116 & new_n2241;
  assign new_n15037 = new_n15036 ^ new_n15035;
  assign new_n15038 = n123 & new_n2240;
  assign new_n15039 = n121 & new_n2391;
  assign new_n15040 = new_n15039 ^ new_n15038;
  assign new_n15041 = new_n15040 ^ new_n15037;
  assign new_n15042 = new_n15041 ^ n30;
  assign new_n15043 = ~new_n3143 & n116;
  assign new_n15044 = ~new_n7503 & new_n3138;
  assign new_n15045 = new_n15044 ^ new_n15043;
  assign new_n15046 = n117 & new_n3137;
  assign new_n15047 = n115 & new_n3149;
  assign new_n15048 = new_n15047 ^ new_n15046;
  assign new_n15049 = new_n15048 ^ new_n15045;
  assign new_n15050 = new_n15049 ^ n36;
  assign new_n15051 = ~new_n3682 & n113;
  assign new_n15052 = ~new_n6764 & new_n3677;
  assign new_n15053 = new_n15052 ^ new_n15051;
  assign new_n15054 = n114 & new_n3676;
  assign new_n15055 = n112 & new_n3688;
  assign new_n15056 = new_n15055 ^ new_n15054;
  assign new_n15057 = new_n15056 ^ new_n15053;
  assign new_n15058 = new_n15057 ^ n39;
  assign new_n15059 = ~new_n4212 & n110;
  assign new_n15060 = new_n4201 & new_n6049;
  assign new_n15061 = new_n15060 ^ new_n15059;
  assign new_n15062 = n111 & new_n4200;
  assign new_n15063 = n109 & new_n4206;
  assign new_n15064 = new_n15063 ^ new_n15062;
  assign new_n15065 = new_n15064 ^ new_n15061;
  assign new_n15066 = new_n15065 ^ n42;
  assign new_n15067 = ~new_n4804 & n107;
  assign new_n15068 = ~new_n5377 & new_n4799;
  assign new_n15069 = new_n15068 ^ new_n15067;
  assign new_n15070 = n108 & new_n4798;
  assign new_n15071 = n106 & new_n4810;
  assign new_n15072 = new_n15071 ^ new_n15070;
  assign new_n15073 = new_n15072 ^ new_n15069;
  assign new_n15074 = new_n15073 ^ n45;
  assign new_n15075 = ~new_n5424 & n104;
  assign new_n15076 = ~new_n4754 & new_n5419;
  assign new_n15077 = new_n15076 ^ new_n15075;
  assign new_n15078 = n105 & new_n5418;
  assign new_n15079 = n103 & new_n5648;
  assign new_n15080 = new_n15079 ^ new_n15078;
  assign new_n15081 = new_n15080 ^ new_n15077;
  assign new_n15082 = new_n15081 ^ n48;
  assign new_n15083 = new_n14950 ^ new_n14886;
  assign new_n15084 = new_n14890 & new_n15083;
  assign new_n15085 = new_n15084 ^ new_n14889;
  assign new_n15086 = new_n15085 ^ new_n15082;
  assign new_n15087 = ~new_n6110 & n101;
  assign new_n15088 = new_n4159 & new_n6105;
  assign new_n15089 = new_n15088 ^ new_n15087;
  assign new_n15090 = n102 & new_n6104;
  assign new_n15091 = n100 & new_n6347;
  assign new_n15092 = new_n15091 ^ new_n15090;
  assign new_n15093 = new_n15092 ^ new_n15089;
  assign new_n15094 = new_n15093 ^ n51;
  assign new_n15095 = ~new_n6805 & n98;
  assign new_n15096 = new_n3604 & new_n6800;
  assign new_n15097 = new_n15096 ^ new_n15095;
  assign new_n15098 = n99 & new_n6799;
  assign new_n15099 = n97 & new_n6811;
  assign new_n15100 = new_n15099 ^ new_n15098;
  assign new_n15101 = new_n15100 ^ new_n15097;
  assign new_n15102 = new_n15101 ^ n54;
  assign new_n15103 = n95 & new_n7553;
  assign new_n15104 = new_n3095 & new_n7543;
  assign new_n15105 = new_n15104 ^ new_n15103;
  assign new_n15106 = n96 & new_n7542;
  assign new_n15107 = n94 & new_n7547;
  assign new_n15108 = new_n15107 ^ new_n15106;
  assign new_n15109 = new_n15108 ^ new_n15105;
  assign new_n15110 = new_n15109 ^ n57;
  assign new_n15111 = n92 & new_n8355;
  assign new_n15112 = new_n2628 & new_n8345;
  assign new_n15113 = new_n15112 ^ new_n15111;
  assign new_n15114 = n93 & new_n8344;
  assign new_n15115 = n91 & new_n8349;
  assign new_n15116 = new_n15115 ^ new_n15114;
  assign new_n15117 = new_n15116 ^ new_n15113;
  assign new_n15118 = new_n15117 ^ n60;
  assign new_n15119 = n87 & new_n9495;
  assign new_n15120 = new_n15119 ^ new_n14927;
  assign new_n15121 = n89 & new_n9195;
  assign new_n15122 = new_n2193 & new_n9185;
  assign new_n15123 = new_n15122 ^ new_n15121;
  assign new_n15124 = n90 & new_n9184;
  assign new_n15125 = n88 & new_n9189;
  assign new_n15126 = new_n15125 ^ new_n15124;
  assign new_n15127 = new_n15126 ^ new_n15123;
  assign new_n15128 = new_n15127 ^ n63;
  assign new_n15129 = n85 ^ n21;
  assign new_n15130 = ~new_n15129 & new_n14931;
  assign new_n15131 = new_n15130 ^ n85;
  assign new_n15132 = new_n11789 & new_n15131;
  assign new_n15133 = new_n15132 ^ new_n15128;
  assign new_n15134 = new_n15133 ^ new_n15120;
  assign new_n15135 = new_n15134 ^ new_n15118;
  assign new_n15136 = new_n14938 ^ new_n14926;
  assign new_n15137 = new_n14934 & new_n15136;
  assign new_n15138 = new_n15137 ^ new_n14938;
  assign new_n15139 = new_n15138 ^ new_n15135;
  assign new_n15140 = new_n15139 ^ new_n15110;
  assign new_n15141 = new_n14939 ^ new_n14914;
  assign new_n15142 = new_n14918 & new_n15141;
  assign new_n15143 = new_n15142 ^ new_n14917;
  assign new_n15144 = new_n15143 ^ new_n15140;
  assign new_n15145 = new_n15144 ^ new_n15102;
  assign new_n15146 = new_n14944 ^ new_n14906;
  assign new_n15147 = new_n14941 & new_n15146;
  assign new_n15148 = new_n15147 ^ new_n14944;
  assign new_n15149 = new_n15148 ^ new_n15145;
  assign new_n15150 = new_n15149 ^ new_n15094;
  assign new_n15151 = new_n14949 ^ new_n14898;
  assign new_n15152 = new_n14946 & new_n15151;
  assign new_n15153 = new_n15152 ^ new_n14949;
  assign new_n15154 = new_n15153 ^ new_n15150;
  assign new_n15155 = new_n15154 ^ new_n15086;
  assign new_n15156 = new_n14963 ^ new_n14951;
  assign new_n15157 = new_n14955 & new_n15156;
  assign new_n15158 = new_n15157 ^ new_n14954;
  assign new_n15159 = new_n15158 ^ new_n15155;
  assign new_n15160 = new_n15159 ^ new_n15074;
  assign new_n15161 = new_n15160 ^ new_n15066;
  assign new_n15162 = new_n14968 ^ new_n14878;
  assign new_n15163 = ~new_n14965 & new_n15162;
  assign new_n15164 = new_n15163 ^ new_n14968;
  assign new_n15165 = new_n15164 ^ new_n15161;
  assign new_n15166 = new_n14973 ^ new_n14969;
  assign new_n15167 = ~new_n15166 & new_n14970;
  assign new_n15168 = new_n15167 ^ new_n14870;
  assign new_n15169 = new_n15168 ^ new_n15165;
  assign new_n15170 = new_n15169 ^ new_n15058;
  assign new_n15171 = new_n14978 ^ new_n14974;
  assign new_n15172 = ~new_n15171 & new_n14975;
  assign new_n15173 = new_n15172 ^ new_n14862;
  assign new_n15174 = new_n15173 ^ new_n15170;
  assign new_n15175 = new_n15174 ^ new_n15050;
  assign new_n15176 = new_n14983 ^ new_n14854;
  assign new_n15177 = ~new_n14980 & new_n15176;
  assign new_n15178 = new_n15177 ^ new_n14983;
  assign new_n15179 = new_n15178 ^ new_n15175;
  assign new_n15180 = ~new_n2672 & n119;
  assign new_n15181 = new_n2667 & new_n8286;
  assign new_n15182 = new_n15181 ^ new_n15180;
  assign new_n15183 = n120 & new_n2666;
  assign new_n15184 = n118 & new_n2664;
  assign new_n15185 = new_n15184 ^ new_n15183;
  assign new_n15186 = new_n15185 ^ new_n15182;
  assign new_n15187 = new_n15186 ^ n33;
  assign new_n15188 = new_n15187 ^ new_n15179;
  assign new_n15189 = new_n14988 ^ new_n14846;
  assign new_n15190 = ~new_n14985 & new_n15189;
  assign new_n15191 = new_n15190 ^ new_n14988;
  assign new_n15192 = new_n15191 ^ new_n15188;
  assign new_n15193 = new_n15192 ^ new_n15042;
  assign new_n15194 = new_n15001 ^ new_n14989;
  assign new_n15195 = ~new_n15194 & new_n14993;
  assign new_n15196 = new_n15195 ^ new_n14992;
  assign new_n15197 = new_n15196 ^ new_n15193;
  assign new_n15198 = new_n15197 ^ new_n15034;
  assign new_n15199 = new_n15006 ^ new_n14838;
  assign new_n15200 = ~new_n15003 & new_n15199;
  assign new_n15201 = new_n15200 ^ new_n15006;
  assign new_n15202 = new_n15201 ^ new_n15198;
  assign new_n15203 = n127 & new_n1512;
  assign new_n15204 = new_n1501 & new_n10010;
  assign new_n15205 = new_n15204 ^ new_n15203;
  assign new_n15206 = ~new_n1506 & n128;
  assign new_n15207 = new_n15206 ^ new_n15205;
  assign new_n15208 = new_n15207 ^ n24;
  assign new_n15209 = new_n15208 ^ new_n15202;
  assign new_n15210 = new_n15011 ^ new_n15007;
  assign new_n15211 = ~new_n15210 & new_n15008;
  assign new_n15212 = new_n15211 ^ new_n14830;
  assign new_n15213 = new_n15212 ^ new_n15209;
  assign new_n15214 = new_n15213 ^ new_n15026;
  assign new_n15215 = n126 & new_n1874;
  assign new_n15216 = new_n1864 & new_n10304;
  assign new_n15217 = new_n15216 ^ new_n15215;
  assign new_n15218 = n127 & new_n1863;
  assign new_n15219 = n125 & new_n1868;
  assign new_n15220 = new_n15219 ^ new_n15218;
  assign new_n15221 = new_n15220 ^ new_n15217;
  assign new_n15222 = new_n15221 ^ n27;
  assign new_n15223 = n123 & new_n2246;
  assign new_n15224 = ~new_n9405 & new_n2241;
  assign new_n15225 = new_n15224 ^ new_n15223;
  assign new_n15226 = n124 & new_n2240;
  assign new_n15227 = n122 & new_n2391;
  assign new_n15228 = new_n15227 ^ new_n15226;
  assign new_n15229 = new_n15228 ^ new_n15225;
  assign new_n15230 = new_n15229 ^ n30;
  assign new_n15231 = ~new_n2672 & n120;
  assign new_n15232 = new_n2667 & new_n8560;
  assign new_n15233 = new_n15232 ^ new_n15231;
  assign new_n15234 = n121 & new_n2666;
  assign new_n15235 = n119 & new_n2664;
  assign new_n15236 = new_n15235 ^ new_n15234;
  assign new_n15237 = new_n15236 ^ new_n15233;
  assign new_n15238 = new_n15237 ^ n33;
  assign new_n15239 = ~new_n3143 & n117;
  assign new_n15240 = ~new_n7761 & new_n3138;
  assign new_n15241 = new_n15240 ^ new_n15239;
  assign new_n15242 = n118 & new_n3137;
  assign new_n15243 = n116 & new_n3149;
  assign new_n15244 = new_n15243 ^ new_n15242;
  assign new_n15245 = new_n15244 ^ new_n15241;
  assign new_n15246 = new_n15245 ^ n36;
  assign new_n15247 = ~new_n3682 & n114;
  assign new_n15248 = ~new_n7013 & new_n3677;
  assign new_n15249 = new_n15248 ^ new_n15247;
  assign new_n15250 = n115 & new_n3676;
  assign new_n15251 = n113 & new_n3688;
  assign new_n15252 = new_n15251 ^ new_n15250;
  assign new_n15253 = new_n15252 ^ new_n15249;
  assign new_n15254 = new_n15253 ^ n39;
  assign new_n15255 = ~new_n4212 & n111;
  assign new_n15256 = ~new_n6284 & new_n4201;
  assign new_n15257 = new_n15256 ^ new_n15255;
  assign new_n15258 = n112 & new_n4200;
  assign new_n15259 = n110 & new_n4206;
  assign new_n15260 = new_n15259 ^ new_n15258;
  assign new_n15261 = new_n15260 ^ new_n15257;
  assign new_n15262 = new_n15261 ^ n42;
  assign new_n15263 = ~new_n5424 & n105;
  assign new_n15264 = ~new_n4961 & new_n5419;
  assign new_n15265 = new_n15264 ^ new_n15263;
  assign new_n15266 = n106 & new_n5418;
  assign new_n15267 = n104 & new_n5648;
  assign new_n15268 = new_n15267 ^ new_n15266;
  assign new_n15269 = new_n15268 ^ new_n15265;
  assign new_n15270 = new_n15269 ^ n48;
  assign new_n15271 = new_n15153 ^ new_n15149;
  assign new_n15272 = ~new_n15150 & new_n15271;
  assign new_n15273 = new_n15272 ^ new_n15094;
  assign new_n15274 = new_n15273 ^ new_n15270;
  assign new_n15275 = ~new_n6110 & n102;
  assign new_n15276 = new_n4368 & new_n6105;
  assign new_n15277 = new_n15276 ^ new_n15275;
  assign new_n15278 = n103 & new_n6104;
  assign new_n15279 = n101 & new_n6347;
  assign new_n15280 = new_n15279 ^ new_n15278;
  assign new_n15281 = new_n15280 ^ new_n15277;
  assign new_n15282 = new_n15281 ^ n51;
  assign new_n15283 = new_n15148 ^ new_n15144;
  assign new_n15284 = ~new_n15145 & new_n15283;
  assign new_n15285 = new_n15284 ^ new_n15102;
  assign new_n15286 = new_n15285 ^ new_n15282;
  assign new_n15287 = ~new_n6805 & n99;
  assign new_n15288 = new_n3789 & new_n6800;
  assign new_n15289 = new_n15288 ^ new_n15287;
  assign new_n15290 = n100 & new_n6799;
  assign new_n15291 = n98 & new_n6811;
  assign new_n15292 = new_n15291 ^ new_n15290;
  assign new_n15293 = new_n15292 ^ new_n15289;
  assign new_n15294 = new_n15293 ^ n54;
  assign new_n15295 = new_n15143 ^ new_n15139;
  assign new_n15296 = ~new_n15140 & new_n15295;
  assign new_n15297 = new_n15296 ^ new_n15110;
  assign new_n15298 = new_n15297 ^ new_n15294;
  assign new_n15299 = n96 & new_n7553;
  assign new_n15300 = new_n3273 & new_n7543;
  assign new_n15301 = new_n15300 ^ new_n15299;
  assign new_n15302 = n97 & new_n7542;
  assign new_n15303 = n95 & new_n7547;
  assign new_n15304 = new_n15303 ^ new_n15302;
  assign new_n15305 = new_n15304 ^ new_n15301;
  assign new_n15306 = new_n15305 ^ n57;
  assign new_n15307 = new_n15138 ^ new_n15134;
  assign new_n15308 = ~new_n15135 & new_n15307;
  assign new_n15309 = new_n15308 ^ new_n15118;
  assign new_n15310 = new_n15309 ^ new_n15306;
  assign new_n15311 = n93 & new_n8355;
  assign new_n15312 = new_n2785 & new_n8345;
  assign new_n15313 = new_n15312 ^ new_n15311;
  assign new_n15314 = n94 & new_n8344;
  assign new_n15315 = n92 & new_n8349;
  assign new_n15316 = new_n15315 ^ new_n15314;
  assign new_n15317 = new_n15316 ^ new_n15313;
  assign new_n15318 = new_n15317 ^ n60;
  assign new_n15319 = new_n15132 ^ new_n15120;
  assign new_n15320 = new_n15133 & new_n15319;
  assign new_n15321 = new_n15320 ^ new_n15128;
  assign new_n15322 = new_n15321 ^ new_n15318;
  assign new_n15323 = n90 & new_n9195;
  assign new_n15324 = new_n2341 & new_n9185;
  assign new_n15325 = new_n15324 ^ new_n15323;
  assign new_n15326 = n91 & new_n9184;
  assign new_n15327 = n89 & new_n9189;
  assign new_n15328 = new_n15327 ^ new_n15326;
  assign new_n15329 = new_n15328 ^ new_n15325;
  assign new_n15330 = new_n15329 ^ n63;
  assign new_n15331 = n64 & new_n1602;
  assign new_n15332 = new_n15331 ^ new_n1707;
  assign new_n15333 = ~new_n9495 & new_n15332;
  assign new_n15334 = new_n15333 ^ new_n1707;
  assign new_n15335 = new_n15334 ^ new_n15330;
  assign new_n15336 = new_n15335 ^ new_n15322;
  assign new_n15337 = new_n15336 ^ new_n15310;
  assign new_n15338 = new_n15337 ^ new_n15298;
  assign new_n15339 = new_n15338 ^ new_n15286;
  assign new_n15340 = new_n15339 ^ new_n15274;
  assign new_n15341 = new_n15154 ^ new_n15085;
  assign new_n15342 = new_n15086 & new_n15341;
  assign new_n15343 = new_n15342 ^ new_n15082;
  assign new_n15344 = new_n15343 ^ new_n15340;
  assign new_n15345 = ~new_n4804 & n108;
  assign new_n15346 = new_n4799 & new_n5604;
  assign new_n15347 = new_n15346 ^ new_n15345;
  assign new_n15348 = n109 & new_n4798;
  assign new_n15349 = n107 & new_n4810;
  assign new_n15350 = new_n15349 ^ new_n15348;
  assign new_n15351 = new_n15350 ^ new_n15347;
  assign new_n15352 = new_n15351 ^ n45;
  assign new_n15353 = new_n15352 ^ new_n15344;
  assign new_n15354 = new_n15155 ^ new_n15074;
  assign new_n15355 = ~new_n15159 & ~new_n15354;
  assign new_n15356 = new_n15355 ^ new_n15074;
  assign new_n15357 = new_n15356 ^ new_n15353;
  assign new_n15358 = new_n15357 ^ new_n15262;
  assign new_n15359 = new_n15164 ^ new_n15066;
  assign new_n15360 = ~new_n15161 & new_n15359;
  assign new_n15361 = new_n15360 ^ new_n15164;
  assign new_n15362 = new_n15361 ^ new_n15358;
  assign new_n15363 = new_n15362 ^ new_n15254;
  assign new_n15364 = new_n15168 ^ new_n15058;
  assign new_n15365 = ~new_n15169 & new_n15364;
  assign new_n15366 = new_n15365 ^ new_n15058;
  assign new_n15367 = new_n15366 ^ new_n15363;
  assign new_n15368 = new_n15367 ^ new_n15246;
  assign new_n15369 = new_n15173 ^ new_n15050;
  assign new_n15370 = ~new_n15174 & new_n15369;
  assign new_n15371 = new_n15370 ^ new_n15050;
  assign new_n15372 = new_n15371 ^ new_n15368;
  assign new_n15373 = new_n15372 ^ new_n15238;
  assign new_n15374 = new_n15187 ^ new_n15175;
  assign new_n15375 = ~new_n15374 & new_n15179;
  assign new_n15376 = new_n15375 ^ new_n15178;
  assign new_n15377 = new_n15376 ^ new_n15373;
  assign new_n15378 = new_n15377 ^ new_n15230;
  assign new_n15379 = new_n15191 ^ new_n15042;
  assign new_n15380 = ~new_n15192 & new_n15379;
  assign new_n15381 = new_n15380 ^ new_n15042;
  assign new_n15382 = new_n15381 ^ new_n15378;
  assign new_n15383 = new_n15382 ^ new_n15222;
  assign new_n15384 = new_n15193 ^ new_n15034;
  assign new_n15385 = ~new_n15197 & new_n15384;
  assign new_n15386 = new_n15385 ^ new_n15034;
  assign new_n15387 = new_n15386 ^ new_n15383;
  assign new_n15388 = ~new_n1511 & n128;
  assign new_n15389 = ~n24 & ~new_n15388;
  assign new_n15390 = new_n15389 ^ n23;
  assign new_n15391 = new_n1306 & new_n11133;
  assign new_n15392 = new_n15391 ^ new_n15388;
  assign new_n15393 = ~new_n15390 & ~new_n15392;
  assign new_n15394 = new_n15393 ^ n23;
  assign new_n15395 = new_n15394 ^ new_n15387;
  assign new_n15396 = new_n15208 ^ new_n15198;
  assign new_n15397 = ~new_n15396 & new_n15202;
  assign new_n15398 = new_n15397 ^ new_n15201;
  assign new_n15399 = new_n15398 ^ new_n15395;
  assign new_n15400 = new_n15212 ^ new_n15026;
  assign new_n15401 = ~new_n15213 & new_n15400;
  assign new_n15402 = new_n15401 ^ new_n15026;
  assign new_n15403 = new_n15402 ^ new_n15399;
  assign new_n15404 = new_n15402 ^ new_n15398;
  assign new_n15405 = new_n15399 & new_n15404;
  assign new_n15406 = new_n15405 ^ new_n15402;
  assign new_n15407 = n127 & new_n1874;
  assign new_n15408 = new_n1864 & new_n10581;
  assign new_n15409 = new_n15408 ^ new_n15407;
  assign new_n15410 = n128 & new_n1863;
  assign new_n15411 = n126 & new_n1868;
  assign new_n15412 = new_n15411 ^ new_n15410;
  assign new_n15413 = new_n15412 ^ new_n15409;
  assign new_n15414 = new_n15413 ^ n27;
  assign new_n15415 = n124 & new_n2246;
  assign new_n15416 = new_n2241 & new_n9700;
  assign new_n15417 = new_n15416 ^ new_n15415;
  assign new_n15418 = n125 & new_n2240;
  assign new_n15419 = n123 & new_n2391;
  assign new_n15420 = new_n15419 ^ new_n15418;
  assign new_n15421 = new_n15420 ^ new_n15417;
  assign new_n15422 = new_n15421 ^ n30;
  assign new_n15423 = ~new_n3143 & n118;
  assign new_n15424 = ~new_n8019 & new_n3138;
  assign new_n15425 = new_n15424 ^ new_n15423;
  assign new_n15426 = n119 & new_n3137;
  assign new_n15427 = n117 & new_n3149;
  assign new_n15428 = new_n15427 ^ new_n15426;
  assign new_n15429 = new_n15428 ^ new_n15425;
  assign new_n15430 = new_n15429 ^ n36;
  assign new_n15431 = ~new_n3682 & n115;
  assign new_n15432 = ~new_n7256 & new_n3677;
  assign new_n15433 = new_n15432 ^ new_n15431;
  assign new_n15434 = n116 & new_n3676;
  assign new_n15435 = n114 & new_n3688;
  assign new_n15436 = new_n15435 ^ new_n15434;
  assign new_n15437 = new_n15436 ^ new_n15433;
  assign new_n15438 = new_n15437 ^ n39;
  assign new_n15439 = ~new_n4212 & n112;
  assign new_n15440 = ~new_n6518 & new_n4201;
  assign new_n15441 = new_n15440 ^ new_n15439;
  assign new_n15442 = n113 & new_n4200;
  assign new_n15443 = n111 & new_n4206;
  assign new_n15444 = new_n15443 ^ new_n15442;
  assign new_n15445 = new_n15444 ^ new_n15441;
  assign new_n15446 = new_n15445 ^ n42;
  assign new_n15447 = ~new_n6110 & n103;
  assign new_n15448 = ~new_n4556 & new_n6105;
  assign new_n15449 = new_n15448 ^ new_n15447;
  assign new_n15450 = n104 & new_n6104;
  assign new_n15451 = n102 & new_n6347;
  assign new_n15452 = new_n15451 ^ new_n15450;
  assign new_n15453 = new_n15452 ^ new_n15449;
  assign new_n15454 = new_n15453 ^ n51;
  assign new_n15455 = new_n15338 ^ new_n15285;
  assign new_n15456 = new_n15286 & new_n15455;
  assign new_n15457 = new_n15456 ^ new_n15282;
  assign new_n15458 = new_n15457 ^ new_n15454;
  assign new_n15459 = ~new_n6805 & n100;
  assign new_n15460 = new_n3972 & new_n6800;
  assign new_n15461 = new_n15460 ^ new_n15459;
  assign new_n15462 = n101 & new_n6799;
  assign new_n15463 = n99 & new_n6811;
  assign new_n15464 = new_n15463 ^ new_n15462;
  assign new_n15465 = new_n15464 ^ new_n15461;
  assign new_n15466 = new_n15465 ^ n54;
  assign new_n15467 = new_n15337 ^ new_n15297;
  assign new_n15468 = new_n15298 & new_n15467;
  assign new_n15469 = new_n15468 ^ new_n15294;
  assign new_n15470 = new_n15469 ^ new_n15466;
  assign new_n15471 = n94 & new_n8355;
  assign new_n15472 = new_n2934 & new_n8345;
  assign new_n15473 = new_n15472 ^ new_n15471;
  assign new_n15474 = n95 & new_n8344;
  assign new_n15475 = n93 & new_n8349;
  assign new_n15476 = new_n15475 ^ new_n15474;
  assign new_n15477 = new_n15476 ^ new_n15473;
  assign new_n15478 = new_n15477 ^ n60;
  assign new_n15479 = new_n15335 ^ new_n15321;
  assign new_n15480 = new_n15322 & new_n15479;
  assign new_n15481 = new_n15480 ^ new_n15318;
  assign new_n15482 = new_n15481 ^ new_n15478;
  assign new_n15483 = new_n15330 ^ n87;
  assign new_n15484 = new_n15483 ^ new_n9495;
  assign new_n15485 = ~new_n15334 & ~new_n15484;
  assign new_n15486 = new_n9495 ^ n87;
  assign new_n15487 = new_n15486 ^ new_n15485;
  assign new_n15488 = n91 & new_n9195;
  assign new_n15489 = new_n2481 & new_n9185;
  assign new_n15490 = new_n15489 ^ new_n15488;
  assign new_n15491 = n92 & new_n9184;
  assign new_n15492 = n90 & new_n9189;
  assign new_n15493 = new_n15492 ^ new_n15491;
  assign new_n15494 = new_n15493 ^ new_n15490;
  assign new_n15495 = new_n15494 ^ n63;
  assign new_n15496 = n89 ^ n87;
  assign new_n15497 = new_n11492 & new_n15496;
  assign new_n15498 = new_n15497 ^ n89;
  assign new_n15499 = new_n15498 ^ n88;
  assign new_n15500 = new_n11789 & new_n15499;
  assign new_n15501 = new_n15500 ^ n24;
  assign new_n15502 = new_n15501 ^ new_n15495;
  assign new_n15503 = new_n15502 ^ new_n15487;
  assign new_n15504 = new_n15503 ^ new_n15482;
  assign new_n15505 = n97 & new_n7553;
  assign new_n15506 = new_n3435 & new_n7543;
  assign new_n15507 = new_n15506 ^ new_n15505;
  assign new_n15508 = n98 & new_n7542;
  assign new_n15509 = n96 & new_n7547;
  assign new_n15510 = new_n15509 ^ new_n15508;
  assign new_n15511 = new_n15510 ^ new_n15507;
  assign new_n15512 = new_n15511 ^ n57;
  assign new_n15513 = new_n15512 ^ new_n15504;
  assign new_n15514 = new_n15336 ^ new_n15309;
  assign new_n15515 = new_n15310 & new_n15514;
  assign new_n15516 = new_n15515 ^ new_n15306;
  assign new_n15517 = new_n15516 ^ new_n15513;
  assign new_n15518 = new_n15517 ^ new_n15470;
  assign new_n15519 = new_n15518 ^ new_n15458;
  assign new_n15520 = new_n15339 ^ new_n15273;
  assign new_n15521 = new_n15274 & new_n15520;
  assign new_n15522 = new_n15521 ^ new_n15270;
  assign new_n15523 = new_n15522 ^ new_n15519;
  assign new_n15524 = ~new_n5424 & n106;
  assign new_n15525 = ~new_n5164 & new_n5419;
  assign new_n15526 = new_n15525 ^ new_n15524;
  assign new_n15527 = n107 & new_n5418;
  assign new_n15528 = n105 & new_n5648;
  assign new_n15529 = new_n15528 ^ new_n15527;
  assign new_n15530 = new_n15529 ^ new_n15526;
  assign new_n15531 = new_n15530 ^ n48;
  assign new_n15532 = new_n15531 ^ new_n15523;
  assign new_n15533 = ~new_n4804 & n109;
  assign new_n15534 = new_n4799 & new_n5825;
  assign new_n15535 = new_n15534 ^ new_n15533;
  assign new_n15536 = n110 & new_n4798;
  assign new_n15537 = n108 & new_n4810;
  assign new_n15538 = new_n15537 ^ new_n15536;
  assign new_n15539 = new_n15538 ^ new_n15535;
  assign new_n15540 = new_n15539 ^ n45;
  assign new_n15541 = new_n15540 ^ new_n15532;
  assign new_n15542 = new_n15352 ^ new_n15340;
  assign new_n15543 = ~new_n15344 & new_n15542;
  assign new_n15544 = new_n15543 ^ new_n15343;
  assign new_n15545 = new_n15544 ^ new_n15541;
  assign new_n15546 = new_n15545 ^ new_n15446;
  assign new_n15547 = new_n15356 ^ new_n15262;
  assign new_n15548 = new_n15357 & new_n15547;
  assign new_n15549 = new_n15548 ^ new_n15262;
  assign new_n15550 = new_n15549 ^ new_n15546;
  assign new_n15551 = new_n15550 ^ new_n15438;
  assign new_n15552 = new_n15361 ^ new_n15254;
  assign new_n15553 = new_n15362 & new_n15552;
  assign new_n15554 = new_n15553 ^ new_n15254;
  assign new_n15555 = new_n15554 ^ new_n15551;
  assign new_n15556 = new_n15555 ^ new_n15430;
  assign new_n15557 = new_n15363 ^ new_n15246;
  assign new_n15558 = ~new_n15557 & new_n15367;
  assign new_n15559 = new_n15558 ^ new_n15246;
  assign new_n15560 = new_n15559 ^ new_n15556;
  assign new_n15561 = new_n15371 ^ new_n15238;
  assign new_n15562 = new_n15372 & new_n15561;
  assign new_n15563 = new_n15562 ^ new_n15238;
  assign new_n15564 = new_n15563 ^ new_n15560;
  assign new_n15565 = ~new_n2672 & n121;
  assign new_n15566 = new_n2667 & new_n8850;
  assign new_n15567 = new_n15566 ^ new_n15565;
  assign new_n15568 = n122 & new_n2666;
  assign new_n15569 = n120 & new_n2664;
  assign new_n15570 = new_n15569 ^ new_n15568;
  assign new_n15571 = new_n15570 ^ new_n15567;
  assign new_n15572 = new_n15571 ^ n33;
  assign new_n15573 = new_n15572 ^ new_n15564;
  assign new_n15574 = new_n15573 ^ new_n15422;
  assign new_n15575 = new_n15376 ^ new_n15230;
  assign new_n15576 = new_n15377 & new_n15575;
  assign new_n15577 = new_n15576 ^ new_n15230;
  assign new_n15578 = new_n15577 ^ new_n15574;
  assign new_n15579 = new_n15578 ^ new_n15414;
  assign new_n15580 = new_n15378 ^ new_n15222;
  assign new_n15581 = ~new_n15580 & new_n15382;
  assign new_n15582 = new_n15581 ^ new_n15222;
  assign new_n15583 = new_n15582 ^ new_n15579;
  assign new_n15584 = new_n15394 ^ new_n15383;
  assign new_n15585 = ~new_n15584 & new_n15387;
  assign new_n15586 = new_n15585 ^ new_n15394;
  assign new_n15587 = new_n15586 ^ new_n15583;
  assign new_n15588 = new_n15587 ^ new_n15406;
  assign new_n15589 = new_n15406 & new_n15587;
  assign new_n15590 = new_n15587 ^ new_n15578;
  assign new_n15591 = new_n15583 & new_n15590;
  assign new_n15592 = new_n15591 ^ new_n15589;
  assign new_n15593 = new_n15414 & new_n15582;
  assign new_n15594 = new_n15582 ^ new_n15414;
  assign new_n15595 = new_n15594 ^ new_n15593;
  assign new_n15596 = new_n15595 ^ new_n15592;
  assign new_n15597 = n125 & new_n2246;
  assign new_n15598 = new_n2241 & new_n9987;
  assign new_n15599 = new_n15598 ^ new_n15597;
  assign new_n15600 = n126 & new_n2240;
  assign new_n15601 = n124 & new_n2391;
  assign new_n15602 = new_n15601 ^ new_n15600;
  assign new_n15603 = new_n15602 ^ new_n15599;
  assign new_n15604 = new_n15603 ^ n30;
  assign new_n15605 = ~new_n2672 & n122;
  assign new_n15606 = ~new_n9116 & new_n2667;
  assign new_n15607 = new_n15606 ^ new_n15605;
  assign new_n15608 = n123 & new_n2666;
  assign new_n15609 = n121 & new_n2664;
  assign new_n15610 = new_n15609 ^ new_n15608;
  assign new_n15611 = new_n15610 ^ new_n15607;
  assign new_n15612 = new_n15611 ^ n33;
  assign new_n15613 = ~new_n3143 & n119;
  assign new_n15614 = new_n3138 & new_n8286;
  assign new_n15615 = new_n15614 ^ new_n15613;
  assign new_n15616 = n120 & new_n3137;
  assign new_n15617 = n118 & new_n3149;
  assign new_n15618 = new_n15617 ^ new_n15616;
  assign new_n15619 = new_n15618 ^ new_n15615;
  assign new_n15620 = new_n15619 ^ n36;
  assign new_n15621 = new_n15554 ^ new_n15438;
  assign new_n15622 = ~new_n15551 & new_n15621;
  assign new_n15623 = new_n15622 ^ new_n15554;
  assign new_n15624 = new_n15623 ^ new_n15620;
  assign new_n15625 = ~new_n3682 & n116;
  assign new_n15626 = ~new_n7503 & new_n3677;
  assign new_n15627 = new_n15626 ^ new_n15625;
  assign new_n15628 = n117 & new_n3676;
  assign new_n15629 = n115 & new_n3688;
  assign new_n15630 = new_n15629 ^ new_n15628;
  assign new_n15631 = new_n15630 ^ new_n15627;
  assign new_n15632 = new_n15631 ^ n39;
  assign new_n15633 = ~new_n4212 & n113;
  assign new_n15634 = ~new_n6764 & new_n4201;
  assign new_n15635 = new_n15634 ^ new_n15633;
  assign new_n15636 = n114 & new_n4200;
  assign new_n15637 = n112 & new_n4206;
  assign new_n15638 = new_n15637 ^ new_n15636;
  assign new_n15639 = new_n15638 ^ new_n15635;
  assign new_n15640 = new_n15639 ^ n42;
  assign new_n15641 = ~new_n4804 & n110;
  assign new_n15642 = new_n4799 & new_n6049;
  assign new_n15643 = new_n15642 ^ new_n15641;
  assign new_n15644 = n111 & new_n4798;
  assign new_n15645 = n109 & new_n4810;
  assign new_n15646 = new_n15645 ^ new_n15644;
  assign new_n15647 = new_n15646 ^ new_n15643;
  assign new_n15648 = new_n15647 ^ n45;
  assign new_n15649 = ~new_n6110 & n104;
  assign new_n15650 = ~new_n4754 & new_n6105;
  assign new_n15651 = new_n15650 ^ new_n15649;
  assign new_n15652 = n105 & new_n6104;
  assign new_n15653 = n103 & new_n6347;
  assign new_n15654 = new_n15653 ^ new_n15652;
  assign new_n15655 = new_n15654 ^ new_n15651;
  assign new_n15656 = new_n15655 ^ n51;
  assign new_n15657 = new_n15517 ^ new_n15466;
  assign new_n15658 = ~new_n15657 & new_n15470;
  assign new_n15659 = new_n15658 ^ new_n15469;
  assign new_n15660 = new_n15659 ^ new_n15656;
  assign new_n15661 = ~new_n6805 & n101;
  assign new_n15662 = new_n4159 & new_n6800;
  assign new_n15663 = new_n15662 ^ new_n15661;
  assign new_n15664 = n102 & new_n6799;
  assign new_n15665 = n100 & new_n6811;
  assign new_n15666 = new_n15665 ^ new_n15664;
  assign new_n15667 = new_n15666 ^ new_n15663;
  assign new_n15668 = new_n15667 ^ n54;
  assign new_n15669 = new_n15516 ^ new_n15504;
  assign new_n15670 = ~new_n15513 & new_n15669;
  assign new_n15671 = new_n15670 ^ new_n15516;
  assign new_n15672 = new_n15671 ^ new_n15668;
  assign new_n15673 = n98 & new_n7553;
  assign new_n15674 = new_n3604 & new_n7543;
  assign new_n15675 = new_n15674 ^ new_n15673;
  assign new_n15676 = n99 & new_n7542;
  assign new_n15677 = n97 & new_n7547;
  assign new_n15678 = new_n15677 ^ new_n15676;
  assign new_n15679 = new_n15678 ^ new_n15675;
  assign new_n15680 = new_n15679 ^ n57;
  assign new_n15681 = n95 & new_n8355;
  assign new_n15682 = new_n3095 & new_n8345;
  assign new_n15683 = new_n15682 ^ new_n15681;
  assign new_n15684 = n96 & new_n8344;
  assign new_n15685 = n94 & new_n8349;
  assign new_n15686 = new_n15685 ^ new_n15684;
  assign new_n15687 = new_n15686 ^ new_n15683;
  assign new_n15688 = new_n15687 ^ n60;
  assign new_n15689 = n92 & new_n9195;
  assign new_n15690 = new_n2628 & new_n9185;
  assign new_n15691 = new_n15690 ^ new_n15689;
  assign new_n15692 = n93 & new_n9184;
  assign new_n15693 = n91 & new_n9189;
  assign new_n15694 = new_n15693 ^ new_n15692;
  assign new_n15695 = new_n15694 ^ new_n15691;
  assign new_n15696 = new_n15695 ^ n63;
  assign new_n15697 = n89 & new_n11492;
  assign new_n15698 = n90 & new_n9495;
  assign new_n15699 = new_n15698 ^ new_n15697;
  assign new_n15700 = n88 ^ n24;
  assign new_n15701 = ~new_n15700 & new_n15499;
  assign new_n15702 = new_n15701 ^ n88;
  assign new_n15703 = new_n11789 & new_n15702;
  assign new_n15704 = new_n15703 ^ new_n15699;
  assign new_n15705 = new_n15704 ^ new_n15696;
  assign new_n15706 = new_n15705 ^ new_n15688;
  assign new_n15707 = new_n15495 ^ new_n15487;
  assign new_n15708 = ~new_n15707 & new_n15502;
  assign new_n15709 = new_n15708 ^ new_n15487;
  assign new_n15710 = new_n15709 ^ new_n15706;
  assign new_n15711 = new_n15710 ^ new_n15680;
  assign new_n15712 = new_n15503 ^ new_n15478;
  assign new_n15713 = ~new_n15712 & new_n15482;
  assign new_n15714 = new_n15713 ^ new_n15481;
  assign new_n15715 = new_n15714 ^ new_n15711;
  assign new_n15716 = new_n15715 ^ new_n15672;
  assign new_n15717 = new_n15716 ^ new_n15660;
  assign new_n15718 = new_n15518 ^ new_n15454;
  assign new_n15719 = ~new_n15718 & new_n15458;
  assign new_n15720 = new_n15719 ^ new_n15457;
  assign new_n15721 = new_n15720 ^ new_n15717;
  assign new_n15722 = ~new_n5424 & n107;
  assign new_n15723 = ~new_n5377 & new_n5419;
  assign new_n15724 = new_n15723 ^ new_n15722;
  assign new_n15725 = n108 & new_n5418;
  assign new_n15726 = n106 & new_n5648;
  assign new_n15727 = new_n15726 ^ new_n15725;
  assign new_n15728 = new_n15727 ^ new_n15724;
  assign new_n15729 = new_n15728 ^ n48;
  assign new_n15730 = new_n15729 ^ new_n15721;
  assign new_n15731 = new_n15730 ^ new_n15648;
  assign new_n15732 = new_n15531 ^ new_n15519;
  assign new_n15733 = ~new_n15732 & new_n15523;
  assign new_n15734 = new_n15733 ^ new_n15522;
  assign new_n15735 = new_n15734 ^ new_n15731;
  assign new_n15736 = new_n15544 ^ new_n15540;
  assign new_n15737 = ~new_n15736 & new_n15541;
  assign new_n15738 = new_n15737 ^ new_n15532;
  assign new_n15739 = new_n15738 ^ new_n15735;
  assign new_n15740 = new_n15739 ^ new_n15640;
  assign new_n15741 = new_n15549 ^ new_n15545;
  assign new_n15742 = ~new_n15741 & new_n15546;
  assign new_n15743 = new_n15742 ^ new_n15446;
  assign new_n15744 = new_n15743 ^ new_n15740;
  assign new_n15745 = new_n15744 ^ new_n15632;
  assign new_n15746 = new_n15745 ^ new_n15624;
  assign new_n15747 = new_n15559 ^ new_n15430;
  assign new_n15748 = ~new_n15556 & new_n15747;
  assign new_n15749 = new_n15748 ^ new_n15559;
  assign new_n15750 = new_n15749 ^ new_n15746;
  assign new_n15751 = new_n15750 ^ new_n15612;
  assign new_n15752 = new_n15572 ^ new_n15560;
  assign new_n15753 = ~new_n15752 & new_n15564;
  assign new_n15754 = new_n15753 ^ new_n15563;
  assign new_n15755 = new_n15754 ^ new_n15751;
  assign new_n15756 = new_n15755 ^ new_n15604;
  assign new_n15757 = new_n15577 ^ new_n15422;
  assign new_n15758 = ~new_n15574 & new_n15757;
  assign new_n15759 = new_n15758 ^ new_n15577;
  assign new_n15760 = new_n15759 ^ new_n15756;
  assign new_n15761 = n127 & new_n1868;
  assign new_n15762 = new_n1864 & new_n10010;
  assign new_n15763 = new_n15762 ^ new_n15761;
  assign new_n15764 = n128 & new_n1874;
  assign new_n15765 = new_n15764 ^ new_n15763;
  assign new_n15766 = new_n15765 ^ n27;
  assign new_n15767 = new_n15766 ^ new_n15760;
  assign new_n15768 = new_n15767 ^ new_n15596;
  assign new_n15769 = ~new_n15593 & ~new_n15767;
  assign new_n15770 = new_n15586 ^ new_n15578;
  assign new_n15771 = new_n15578 ^ new_n15406;
  assign new_n15772 = ~new_n15771 & new_n15770;
  assign new_n15773 = new_n15772 ^ new_n15586;
  assign new_n15774 = ~new_n15769 & new_n15773;
  assign new_n15775 = ~new_n15578 & ~new_n15586;
  assign new_n15776 = new_n15775 ^ new_n15770;
  assign new_n15777 = ~new_n15767 & new_n15776;
  assign new_n15778 = ~new_n15777 & new_n15595;
  assign new_n15779 = new_n15406 & new_n15778;
  assign new_n15780 = new_n15775 ^ new_n15582;
  assign new_n15781 = ~new_n15780 & new_n15594;
  assign new_n15782 = new_n15781 ^ new_n15582;
  assign new_n15783 = new_n15767 & new_n15782;
  assign new_n15784 = ~new_n15779 & ~new_n15783;
  assign new_n15785 = ~new_n15774 & new_n15784;
  assign new_n15786 = n126 & new_n2246;
  assign new_n15787 = new_n2241 & new_n10304;
  assign new_n15788 = new_n15787 ^ new_n15786;
  assign new_n15789 = n127 & new_n2240;
  assign new_n15790 = n125 & new_n2391;
  assign new_n15791 = new_n15790 ^ new_n15789;
  assign new_n15792 = new_n15791 ^ new_n15788;
  assign new_n15793 = new_n15792 ^ n30;
  assign new_n15794 = ~new_n2672 & n123;
  assign new_n15795 = ~new_n9405 & new_n2667;
  assign new_n15796 = new_n15795 ^ new_n15794;
  assign new_n15797 = n124 & new_n2666;
  assign new_n15798 = n122 & new_n2664;
  assign new_n15799 = new_n15798 ^ new_n15797;
  assign new_n15800 = new_n15799 ^ new_n15796;
  assign new_n15801 = new_n15800 ^ n33;
  assign new_n15802 = ~new_n3682 & n117;
  assign new_n15803 = ~new_n7761 & new_n3677;
  assign new_n15804 = new_n15803 ^ new_n15802;
  assign new_n15805 = n118 & new_n3676;
  assign new_n15806 = n116 & new_n3688;
  assign new_n15807 = new_n15806 ^ new_n15805;
  assign new_n15808 = new_n15807 ^ new_n15804;
  assign new_n15809 = new_n15808 ^ n39;
  assign new_n15810 = ~new_n4212 & n114;
  assign new_n15811 = ~new_n7013 & new_n4201;
  assign new_n15812 = new_n15811 ^ new_n15810;
  assign new_n15813 = n115 & new_n4200;
  assign new_n15814 = n113 & new_n4206;
  assign new_n15815 = new_n15814 ^ new_n15813;
  assign new_n15816 = new_n15815 ^ new_n15812;
  assign new_n15817 = new_n15816 ^ n42;
  assign new_n15818 = ~new_n4804 & n111;
  assign new_n15819 = ~new_n6284 & new_n4799;
  assign new_n15820 = new_n15819 ^ new_n15818;
  assign new_n15821 = n112 & new_n4798;
  assign new_n15822 = n110 & new_n4810;
  assign new_n15823 = new_n15822 ^ new_n15821;
  assign new_n15824 = new_n15823 ^ new_n15820;
  assign new_n15825 = new_n15824 ^ n45;
  assign new_n15826 = ~new_n5424 & n108;
  assign new_n15827 = new_n5419 & new_n5604;
  assign new_n15828 = new_n15827 ^ new_n15826;
  assign new_n15829 = n109 & new_n5418;
  assign new_n15830 = n107 & new_n5648;
  assign new_n15831 = new_n15830 ^ new_n15829;
  assign new_n15832 = new_n15831 ^ new_n15828;
  assign new_n15833 = new_n15832 ^ n48;
  assign new_n15834 = ~new_n6110 & n105;
  assign new_n15835 = ~new_n4961 & new_n6105;
  assign new_n15836 = new_n15835 ^ new_n15834;
  assign new_n15837 = n106 & new_n6104;
  assign new_n15838 = n104 & new_n6347;
  assign new_n15839 = new_n15838 ^ new_n15837;
  assign new_n15840 = new_n15839 ^ new_n15836;
  assign new_n15841 = new_n15840 ^ n51;
  assign new_n15842 = ~new_n6805 & n102;
  assign new_n15843 = new_n4368 & new_n6800;
  assign new_n15844 = new_n15843 ^ new_n15842;
  assign new_n15845 = n103 & new_n6799;
  assign new_n15846 = n101 & new_n6811;
  assign new_n15847 = new_n15846 ^ new_n15845;
  assign new_n15848 = new_n15847 ^ new_n15844;
  assign new_n15849 = new_n15848 ^ n54;
  assign new_n15850 = n99 & new_n7553;
  assign new_n15851 = new_n3789 & new_n7543;
  assign new_n15852 = new_n15851 ^ new_n15850;
  assign new_n15853 = n100 & new_n7542;
  assign new_n15854 = n98 & new_n7547;
  assign new_n15855 = new_n15854 ^ new_n15853;
  assign new_n15856 = new_n15855 ^ new_n15852;
  assign new_n15857 = new_n15856 ^ n57;
  assign new_n15858 = n96 & new_n8355;
  assign new_n15859 = new_n3273 & new_n8345;
  assign new_n15860 = new_n15859 ^ new_n15858;
  assign new_n15861 = n97 & new_n8344;
  assign new_n15862 = n95 & new_n8349;
  assign new_n15863 = new_n15862 ^ new_n15861;
  assign new_n15864 = new_n15863 ^ new_n15860;
  assign new_n15865 = new_n15864 ^ n60;
  assign new_n15866 = n93 & new_n9195;
  assign new_n15867 = new_n2785 & new_n9185;
  assign new_n15868 = new_n15867 ^ new_n15866;
  assign new_n15869 = n94 & new_n9184;
  assign new_n15870 = n92 & new_n9189;
  assign new_n15871 = new_n15870 ^ new_n15869;
  assign new_n15872 = new_n15871 ^ new_n15868;
  assign new_n15873 = new_n15872 ^ n63;
  assign new_n15874 = n90 & new_n11789;
  assign new_n15875 = ~n91 & new_n9495;
  assign new_n15876 = new_n15875 ^ new_n15697;
  assign new_n15877 = new_n15876 ^ new_n9495;
  assign new_n15878 = new_n15877 ^ new_n15874;
  assign new_n15879 = new_n15878 ^ new_n15873;
  assign new_n15880 = new_n15703 ^ new_n15696;
  assign new_n15881 = new_n15704 & new_n15880;
  assign new_n15882 = new_n15881 ^ new_n15696;
  assign new_n15883 = new_n15882 ^ new_n15879;
  assign new_n15884 = new_n15883 ^ new_n15865;
  assign new_n15885 = new_n15884 ^ new_n15857;
  assign new_n15886 = new_n15709 ^ new_n15705;
  assign new_n15887 = ~new_n15706 & ~new_n15886;
  assign new_n15888 = new_n15887 ^ new_n15688;
  assign new_n15889 = new_n15888 ^ new_n15885;
  assign new_n15890 = new_n15889 ^ new_n15849;
  assign new_n15891 = new_n15714 ^ new_n15710;
  assign new_n15892 = ~new_n15891 & new_n15711;
  assign new_n15893 = new_n15892 ^ new_n15680;
  assign new_n15894 = new_n15893 ^ new_n15890;
  assign new_n15895 = new_n15715 ^ new_n15671;
  assign new_n15896 = ~new_n15895 & new_n15672;
  assign new_n15897 = new_n15896 ^ new_n15668;
  assign new_n15898 = new_n15897 ^ new_n15894;
  assign new_n15899 = new_n15898 ^ new_n15841;
  assign new_n15900 = new_n15899 ^ new_n15833;
  assign new_n15901 = new_n15716 ^ new_n15659;
  assign new_n15902 = ~new_n15901 & new_n15660;
  assign new_n15903 = new_n15902 ^ new_n15656;
  assign new_n15904 = new_n15903 ^ new_n15900;
  assign new_n15905 = new_n15729 ^ new_n15717;
  assign new_n15906 = ~new_n15905 & new_n15721;
  assign new_n15907 = new_n15906 ^ new_n15720;
  assign new_n15908 = new_n15907 ^ new_n15904;
  assign new_n15909 = new_n15908 ^ new_n15825;
  assign new_n15910 = new_n15734 ^ new_n15648;
  assign new_n15911 = ~new_n15731 & new_n15910;
  assign new_n15912 = new_n15911 ^ new_n15734;
  assign new_n15913 = new_n15912 ^ new_n15909;
  assign new_n15914 = new_n15913 ^ new_n15817;
  assign new_n15915 = new_n15738 ^ new_n15640;
  assign new_n15916 = ~new_n15739 & new_n15915;
  assign new_n15917 = new_n15916 ^ new_n15640;
  assign new_n15918 = new_n15917 ^ new_n15914;
  assign new_n15919 = new_n15918 ^ new_n15809;
  assign new_n15920 = new_n15743 ^ new_n15632;
  assign new_n15921 = ~new_n15744 & new_n15920;
  assign new_n15922 = new_n15921 ^ new_n15632;
  assign new_n15923 = new_n15922 ^ new_n15919;
  assign new_n15924 = ~new_n3143 & n120;
  assign new_n15925 = new_n3138 & new_n8560;
  assign new_n15926 = new_n15925 ^ new_n15924;
  assign new_n15927 = n121 & new_n3137;
  assign new_n15928 = n119 & new_n3149;
  assign new_n15929 = new_n15928 ^ new_n15927;
  assign new_n15930 = new_n15929 ^ new_n15926;
  assign new_n15931 = new_n15930 ^ n36;
  assign new_n15932 = new_n15931 ^ new_n15923;
  assign new_n15933 = new_n15745 ^ new_n15620;
  assign new_n15934 = ~new_n15933 & new_n15624;
  assign new_n15935 = new_n15934 ^ new_n15623;
  assign new_n15936 = new_n15935 ^ new_n15932;
  assign new_n15937 = new_n15936 ^ new_n15801;
  assign new_n15938 = new_n15749 ^ new_n15612;
  assign new_n15939 = ~new_n15750 & new_n15938;
  assign new_n15940 = new_n15939 ^ new_n15612;
  assign new_n15941 = new_n15940 ^ new_n15937;
  assign new_n15942 = new_n15941 ^ new_n15793;
  assign new_n15943 = n128 & new_n1868;
  assign new_n15944 = new_n1864 & new_n11133;
  assign new_n15945 = new_n15944 ^ new_n15943;
  assign new_n15946 = new_n15945 ^ n27;
  assign new_n15947 = new_n15946 ^ new_n15942;
  assign new_n15948 = new_n15751 ^ new_n15604;
  assign new_n15949 = ~new_n15755 & new_n15948;
  assign new_n15950 = new_n15949 ^ new_n15604;
  assign new_n15951 = new_n15950 ^ new_n15947;
  assign new_n15952 = new_n15766 ^ new_n15756;
  assign new_n15953 = ~new_n15952 & new_n15760;
  assign new_n15954 = new_n15953 ^ new_n15759;
  assign new_n15955 = new_n15954 ^ new_n15951;
  assign new_n15956 = new_n15955 ^ new_n15785;
  assign new_n15957 = ~new_n15950 & ~new_n15954;
  assign new_n15958 = new_n15954 ^ new_n15950;
  assign new_n15959 = new_n15958 ^ new_n15957;
  assign new_n15960 = ~new_n15947 & ~new_n15959;
  assign new_n15961 = new_n15957 ^ new_n15785;
  assign new_n15962 = ~new_n15946 & new_n15942;
  assign new_n15963 = new_n15962 ^ new_n15947;
  assign new_n15964 = new_n15963 ^ new_n15957;
  assign new_n15965 = new_n15964 ^ new_n15962;
  assign new_n15966 = ~new_n15965 & new_n15961;
  assign new_n15967 = new_n15966 ^ new_n15963;
  assign new_n15968 = new_n15785 & new_n15959;
  assign new_n15969 = new_n15968 ^ new_n15967;
  assign new_n15970 = new_n15969 ^ new_n15960;
  assign new_n15971 = n127 & new_n2246;
  assign new_n15972 = new_n2241 & new_n10581;
  assign new_n15973 = new_n15972 ^ new_n15971;
  assign new_n15974 = n128 & new_n2240;
  assign new_n15975 = n126 & new_n2391;
  assign new_n15976 = new_n15975 ^ new_n15974;
  assign new_n15977 = new_n15976 ^ new_n15973;
  assign new_n15978 = new_n15977 ^ n30;
  assign new_n15979 = ~new_n2672 & n124;
  assign new_n15980 = new_n2667 & new_n9700;
  assign new_n15981 = new_n15980 ^ new_n15979;
  assign new_n15982 = n125 & new_n2666;
  assign new_n15983 = n123 & new_n2664;
  assign new_n15984 = new_n15983 ^ new_n15982;
  assign new_n15985 = new_n15984 ^ new_n15981;
  assign new_n15986 = new_n15985 ^ n33;
  assign new_n15987 = ~new_n3682 & n118;
  assign new_n15988 = ~new_n8019 & new_n3677;
  assign new_n15989 = new_n15988 ^ new_n15987;
  assign new_n15990 = n119 & new_n3676;
  assign new_n15991 = n117 & new_n3688;
  assign new_n15992 = new_n15991 ^ new_n15990;
  assign new_n15993 = new_n15992 ^ new_n15989;
  assign new_n15994 = new_n15993 ^ n39;
  assign new_n15995 = ~new_n4212 & n115;
  assign new_n15996 = ~new_n7256 & new_n4201;
  assign new_n15997 = new_n15996 ^ new_n15995;
  assign new_n15998 = n116 & new_n4200;
  assign new_n15999 = n114 & new_n4206;
  assign new_n16000 = new_n15999 ^ new_n15998;
  assign new_n16001 = new_n16000 ^ new_n15997;
  assign new_n16002 = new_n16001 ^ n42;
  assign new_n16003 = ~new_n4804 & n112;
  assign new_n16004 = ~new_n6518 & new_n4799;
  assign new_n16005 = new_n16004 ^ new_n16003;
  assign new_n16006 = n113 & new_n4798;
  assign new_n16007 = n111 & new_n4810;
  assign new_n16008 = new_n16007 ^ new_n16006;
  assign new_n16009 = new_n16008 ^ new_n16005;
  assign new_n16010 = new_n16009 ^ n45;
  assign new_n16011 = ~new_n6110 & n106;
  assign new_n16012 = ~new_n5164 & new_n6105;
  assign new_n16013 = new_n16012 ^ new_n16011;
  assign new_n16014 = n107 & new_n6104;
  assign new_n16015 = n105 & new_n6347;
  assign new_n16016 = new_n16015 ^ new_n16014;
  assign new_n16017 = new_n16016 ^ new_n16013;
  assign new_n16018 = new_n16017 ^ n51;
  assign new_n16019 = new_n15894 ^ new_n15841;
  assign new_n16020 = ~new_n16019 & new_n15898;
  assign new_n16021 = new_n16020 ^ new_n15841;
  assign new_n16022 = new_n16021 ^ new_n16018;
  assign new_n16023 = ~new_n6805 & n103;
  assign new_n16024 = ~new_n4556 & new_n6800;
  assign new_n16025 = new_n16024 ^ new_n16023;
  assign new_n16026 = n104 & new_n6799;
  assign new_n16027 = n102 & new_n6811;
  assign new_n16028 = new_n16027 ^ new_n16026;
  assign new_n16029 = new_n16028 ^ new_n16025;
  assign new_n16030 = new_n16029 ^ n54;
  assign new_n16031 = new_n15893 ^ new_n15889;
  assign new_n16032 = ~new_n15890 & new_n16031;
  assign new_n16033 = new_n16032 ^ new_n15849;
  assign new_n16034 = new_n16033 ^ new_n16030;
  assign new_n16035 = n100 & new_n7553;
  assign new_n16036 = new_n3972 & new_n7543;
  assign new_n16037 = new_n16036 ^ new_n16035;
  assign new_n16038 = n101 & new_n7542;
  assign new_n16039 = n99 & new_n7547;
  assign new_n16040 = new_n16039 ^ new_n16038;
  assign new_n16041 = new_n16040 ^ new_n16037;
  assign new_n16042 = new_n16041 ^ n57;
  assign new_n16043 = n97 & new_n8355;
  assign new_n16044 = new_n3435 & new_n8345;
  assign new_n16045 = new_n16044 ^ new_n16043;
  assign new_n16046 = n98 & new_n8344;
  assign new_n16047 = n96 & new_n8349;
  assign new_n16048 = new_n16047 ^ new_n16046;
  assign new_n16049 = new_n16048 ^ new_n16045;
  assign new_n16050 = new_n16049 ^ n60;
  assign new_n16051 = n92 ^ n90;
  assign new_n16052 = ~new_n11492 & new_n16051;
  assign new_n16053 = new_n16052 ^ n90;
  assign new_n16054 = new_n16053 ^ n91;
  assign new_n16055 = new_n11789 & new_n16054;
  assign new_n16056 = new_n16055 ^ n27;
  assign new_n16057 = n90 & new_n15876;
  assign new_n16058 = new_n16057 ^ new_n15697;
  assign new_n16059 = ~new_n15878 & new_n15873;
  assign new_n16060 = new_n16059 ^ new_n16058;
  assign new_n16061 = new_n16060 ^ new_n16056;
  assign new_n16062 = n94 & new_n9195;
  assign new_n16063 = new_n2934 & new_n9185;
  assign new_n16064 = new_n16063 ^ new_n16062;
  assign new_n16065 = n95 & new_n9184;
  assign new_n16066 = n93 & new_n9189;
  assign new_n16067 = new_n16066 ^ new_n16065;
  assign new_n16068 = new_n16067 ^ new_n16064;
  assign new_n16069 = new_n16068 ^ n63;
  assign new_n16070 = new_n16069 ^ new_n16061;
  assign new_n16071 = new_n16070 ^ new_n16050;
  assign new_n16072 = new_n15882 ^ new_n15865;
  assign new_n16073 = new_n15883 & new_n16072;
  assign new_n16074 = new_n16073 ^ new_n15865;
  assign new_n16075 = new_n16074 ^ new_n16071;
  assign new_n16076 = new_n16075 ^ new_n16042;
  assign new_n16077 = new_n15888 ^ new_n15884;
  assign new_n16078 = ~new_n15885 & new_n16077;
  assign new_n16079 = new_n16078 ^ new_n15857;
  assign new_n16080 = new_n16079 ^ new_n16076;
  assign new_n16081 = new_n16080 ^ new_n16034;
  assign new_n16082 = new_n16081 ^ new_n16022;
  assign new_n16083 = ~new_n5424 & n109;
  assign new_n16084 = new_n5419 & new_n5825;
  assign new_n16085 = new_n16084 ^ new_n16083;
  assign new_n16086 = n110 & new_n5418;
  assign new_n16087 = n108 & new_n5648;
  assign new_n16088 = new_n16087 ^ new_n16086;
  assign new_n16089 = new_n16088 ^ new_n16085;
  assign new_n16090 = new_n16089 ^ n48;
  assign new_n16091 = new_n16090 ^ new_n16082;
  assign new_n16092 = new_n15903 ^ new_n15899;
  assign new_n16093 = ~new_n15900 & new_n16092;
  assign new_n16094 = new_n16093 ^ new_n15833;
  assign new_n16095 = new_n16094 ^ new_n16091;
  assign new_n16096 = new_n16095 ^ new_n16010;
  assign new_n16097 = new_n15907 ^ new_n15825;
  assign new_n16098 = new_n15908 & new_n16097;
  assign new_n16099 = new_n16098 ^ new_n15825;
  assign new_n16100 = new_n16099 ^ new_n16096;
  assign new_n16101 = new_n16100 ^ new_n16002;
  assign new_n16102 = new_n15909 ^ new_n15817;
  assign new_n16103 = ~new_n16102 & new_n15913;
  assign new_n16104 = new_n16103 ^ new_n15817;
  assign new_n16105 = new_n16104 ^ new_n16101;
  assign new_n16106 = new_n16105 ^ new_n15994;
  assign new_n16107 = new_n15914 ^ new_n15809;
  assign new_n16108 = ~new_n16107 & new_n15918;
  assign new_n16109 = new_n16108 ^ new_n15809;
  assign new_n16110 = new_n16109 ^ new_n16106;
  assign new_n16111 = new_n15931 ^ new_n15922;
  assign new_n16112 = ~new_n15923 & ~new_n16111;
  assign new_n16113 = new_n16112 ^ new_n15919;
  assign new_n16114 = new_n16113 ^ new_n16110;
  assign new_n16115 = ~new_n3143 & n121;
  assign new_n16116 = new_n3138 & new_n8850;
  assign new_n16117 = new_n16116 ^ new_n16115;
  assign new_n16118 = n122 & new_n3137;
  assign new_n16119 = n120 & new_n3149;
  assign new_n16120 = new_n16119 ^ new_n16118;
  assign new_n16121 = new_n16120 ^ new_n16117;
  assign new_n16122 = new_n16121 ^ n36;
  assign new_n16123 = new_n16122 ^ new_n16114;
  assign new_n16124 = new_n16123 ^ new_n15986;
  assign new_n16125 = new_n15935 ^ new_n15801;
  assign new_n16126 = new_n15936 & new_n16125;
  assign new_n16127 = new_n16126 ^ new_n15801;
  assign new_n16128 = new_n16127 ^ new_n16124;
  assign new_n16129 = new_n16128 ^ new_n15978;
  assign new_n16130 = new_n15940 ^ new_n15793;
  assign new_n16131 = new_n15941 & new_n16130;
  assign new_n16132 = new_n16131 ^ new_n15793;
  assign new_n16133 = new_n16132 ^ new_n16129;
  assign new_n16134 = new_n16133 ^ new_n15970;
  assign new_n16135 = ~new_n15963 & ~new_n16133;
  assign new_n16136 = ~new_n15957 & ~new_n16135;
  assign new_n16137 = ~new_n15968 & new_n16136;
  assign new_n16138 = ~new_n16133 & new_n15959;
  assign new_n16139 = ~new_n15962 & ~new_n16138;
  assign new_n16140 = ~new_n15785 & new_n16139;
  assign new_n16141 = new_n15957 ^ new_n15946;
  assign new_n16142 = ~new_n15947 & new_n16141;
  assign new_n16143 = new_n16142 ^ new_n15942;
  assign new_n16144 = ~new_n16143 & new_n16133;
  assign new_n16145 = ~new_n16140 & ~new_n16144;
  assign new_n16146 = ~new_n16137 & new_n16145;
  assign new_n16147 = ~new_n2672 & n125;
  assign new_n16148 = new_n2667 & new_n9987;
  assign new_n16149 = new_n16148 ^ new_n16147;
  assign new_n16150 = n126 & new_n2666;
  assign new_n16151 = n124 & new_n2664;
  assign new_n16152 = new_n16151 ^ new_n16150;
  assign new_n16153 = new_n16152 ^ new_n16149;
  assign new_n16154 = new_n16153 ^ n33;
  assign new_n16155 = ~new_n3143 & n122;
  assign new_n16156 = ~new_n9116 & new_n3138;
  assign new_n16157 = new_n16156 ^ new_n16155;
  assign new_n16158 = n123 & new_n3137;
  assign new_n16159 = n121 & new_n3149;
  assign new_n16160 = new_n16159 ^ new_n16158;
  assign new_n16161 = new_n16160 ^ new_n16157;
  assign new_n16162 = new_n16161 ^ n36;
  assign new_n16163 = ~new_n3682 & n119;
  assign new_n16164 = new_n3677 & new_n8286;
  assign new_n16165 = new_n16164 ^ new_n16163;
  assign new_n16166 = n120 & new_n3676;
  assign new_n16167 = n118 & new_n3688;
  assign new_n16168 = new_n16167 ^ new_n16166;
  assign new_n16169 = new_n16168 ^ new_n16165;
  assign new_n16170 = new_n16169 ^ n39;
  assign new_n16171 = ~new_n4212 & n116;
  assign new_n16172 = ~new_n7503 & new_n4201;
  assign new_n16173 = new_n16172 ^ new_n16171;
  assign new_n16174 = n117 & new_n4200;
  assign new_n16175 = n115 & new_n4206;
  assign new_n16176 = new_n16175 ^ new_n16174;
  assign new_n16177 = new_n16176 ^ new_n16173;
  assign new_n16178 = new_n16177 ^ n42;
  assign new_n16179 = ~new_n6805 & n104;
  assign new_n16180 = ~new_n4754 & new_n6800;
  assign new_n16181 = new_n16180 ^ new_n16179;
  assign new_n16182 = n105 & new_n6799;
  assign new_n16183 = n103 & new_n6811;
  assign new_n16184 = new_n16183 ^ new_n16182;
  assign new_n16185 = new_n16184 ^ new_n16181;
  assign new_n16186 = new_n16185 ^ n54;
  assign new_n16187 = n101 & new_n7553;
  assign new_n16188 = new_n4159 & new_n7543;
  assign new_n16189 = new_n16188 ^ new_n16187;
  assign new_n16190 = n102 & new_n7542;
  assign new_n16191 = n100 & new_n7547;
  assign new_n16192 = new_n16191 ^ new_n16190;
  assign new_n16193 = new_n16192 ^ new_n16189;
  assign new_n16194 = new_n16193 ^ n57;
  assign new_n16195 = new_n16074 ^ new_n16070;
  assign new_n16196 = ~new_n16071 & new_n16195;
  assign new_n16197 = new_n16196 ^ new_n16050;
  assign new_n16198 = new_n16197 ^ new_n16194;
  assign new_n16199 = n98 & new_n8355;
  assign new_n16200 = new_n3604 & new_n8345;
  assign new_n16201 = new_n16200 ^ new_n16199;
  assign new_n16202 = n99 & new_n8344;
  assign new_n16203 = n97 & new_n8349;
  assign new_n16204 = new_n16203 ^ new_n16202;
  assign new_n16205 = new_n16204 ^ new_n16201;
  assign new_n16206 = new_n16205 ^ n60;
  assign new_n16207 = n95 & new_n9195;
  assign new_n16208 = new_n3095 & new_n9185;
  assign new_n16209 = new_n16208 ^ new_n16207;
  assign new_n16210 = n96 & new_n9184;
  assign new_n16211 = n94 & new_n9189;
  assign new_n16212 = new_n16211 ^ new_n16210;
  assign new_n16213 = new_n16212 ^ new_n16209;
  assign new_n16214 = new_n16213 ^ n63;
  assign new_n16215 = n64 & n92;
  assign new_n16216 = new_n16215 ^ n93;
  assign new_n16217 = ~new_n9495 & new_n16216;
  assign new_n16218 = new_n16217 ^ n93;
  assign new_n16219 = n91 ^ n27;
  assign new_n16220 = ~new_n16219 & new_n16054;
  assign new_n16221 = new_n16220 ^ n91;
  assign new_n16222 = new_n11789 & new_n16221;
  assign new_n16223 = new_n16222 ^ new_n16218;
  assign new_n16224 = new_n16223 ^ new_n16214;
  assign new_n16225 = new_n16224 ^ new_n16206;
  assign new_n16226 = new_n16069 ^ new_n16056;
  assign new_n16227 = ~new_n16061 & new_n16226;
  assign new_n16228 = new_n16227 ^ new_n16060;
  assign new_n16229 = new_n16228 ^ new_n16225;
  assign new_n16230 = new_n16229 ^ new_n16198;
  assign new_n16231 = new_n16230 ^ new_n16186;
  assign new_n16232 = new_n16079 ^ new_n16042;
  assign new_n16233 = new_n16076 & new_n16232;
  assign new_n16234 = new_n16233 ^ new_n16079;
  assign new_n16235 = new_n16234 ^ new_n16231;
  assign new_n16236 = new_n16080 ^ new_n16030;
  assign new_n16237 = new_n16034 & new_n16236;
  assign new_n16238 = new_n16237 ^ new_n16033;
  assign new_n16239 = new_n16238 ^ new_n16235;
  assign new_n16240 = ~new_n6110 & n107;
  assign new_n16241 = ~new_n5377 & new_n6105;
  assign new_n16242 = new_n16241 ^ new_n16240;
  assign new_n16243 = n108 & new_n6104;
  assign new_n16244 = n106 & new_n6347;
  assign new_n16245 = new_n16244 ^ new_n16243;
  assign new_n16246 = new_n16245 ^ new_n16242;
  assign new_n16247 = new_n16246 ^ n51;
  assign new_n16248 = new_n16247 ^ new_n16239;
  assign new_n16249 = new_n16081 ^ new_n16018;
  assign new_n16250 = new_n16022 & new_n16249;
  assign new_n16251 = new_n16250 ^ new_n16021;
  assign new_n16252 = new_n16251 ^ new_n16248;
  assign new_n16253 = ~new_n5424 & n110;
  assign new_n16254 = new_n5419 & new_n6049;
  assign new_n16255 = new_n16254 ^ new_n16253;
  assign new_n16256 = n111 & new_n5418;
  assign new_n16257 = n109 & new_n5648;
  assign new_n16258 = new_n16257 ^ new_n16256;
  assign new_n16259 = new_n16258 ^ new_n16255;
  assign new_n16260 = new_n16259 ^ n48;
  assign new_n16261 = new_n16260 ^ new_n16252;
  assign new_n16262 = new_n16094 ^ new_n16090;
  assign new_n16263 = ~new_n16091 & ~new_n16262;
  assign new_n16264 = new_n16263 ^ new_n16082;
  assign new_n16265 = new_n16264 ^ new_n16261;
  assign new_n16266 = ~new_n4804 & n113;
  assign new_n16267 = ~new_n6764 & new_n4799;
  assign new_n16268 = new_n16267 ^ new_n16266;
  assign new_n16269 = n114 & new_n4798;
  assign new_n16270 = n112 & new_n4810;
  assign new_n16271 = new_n16270 ^ new_n16269;
  assign new_n16272 = new_n16271 ^ new_n16268;
  assign new_n16273 = new_n16272 ^ n45;
  assign new_n16274 = new_n16273 ^ new_n16265;
  assign new_n16275 = new_n16099 ^ new_n16095;
  assign new_n16276 = ~new_n16096 & new_n16275;
  assign new_n16277 = new_n16276 ^ new_n16010;
  assign new_n16278 = new_n16277 ^ new_n16274;
  assign new_n16279 = new_n16278 ^ new_n16178;
  assign new_n16280 = new_n16104 ^ new_n16100;
  assign new_n16281 = ~new_n16101 & new_n16280;
  assign new_n16282 = new_n16281 ^ new_n16002;
  assign new_n16283 = new_n16282 ^ new_n16279;
  assign new_n16284 = new_n16283 ^ new_n16170;
  assign new_n16285 = new_n16109 ^ new_n16105;
  assign new_n16286 = ~new_n16106 & new_n16285;
  assign new_n16287 = new_n16286 ^ new_n15994;
  assign new_n16288 = new_n16287 ^ new_n16284;
  assign new_n16289 = new_n16288 ^ new_n16162;
  assign new_n16290 = new_n16122 ^ new_n16110;
  assign new_n16291 = new_n16114 & new_n16290;
  assign new_n16292 = new_n16291 ^ new_n16113;
  assign new_n16293 = new_n16292 ^ new_n16289;
  assign new_n16294 = new_n16293 ^ new_n16154;
  assign new_n16295 = new_n16127 ^ new_n15986;
  assign new_n16296 = ~new_n16124 & new_n16295;
  assign new_n16297 = new_n16296 ^ new_n16127;
  assign new_n16298 = new_n16297 ^ new_n16294;
  assign new_n16299 = n127 & new_n2391;
  assign new_n16300 = new_n2241 & new_n10010;
  assign new_n16301 = new_n16300 ^ new_n16299;
  assign new_n16302 = n128 & new_n2246;
  assign new_n16303 = new_n16302 ^ new_n16301;
  assign new_n16304 = new_n16303 ^ n30;
  assign new_n16305 = new_n16304 ^ new_n16298;
  assign new_n16306 = new_n16132 ^ new_n15978;
  assign new_n16307 = ~new_n16129 & new_n16306;
  assign new_n16308 = new_n16307 ^ new_n16132;
  assign new_n16309 = new_n16308 ^ new_n16305;
  assign new_n16310 = new_n16309 ^ new_n16146;
  assign new_n16311 = ~new_n2672 & n126;
  assign new_n16312 = new_n2667 & new_n10304;
  assign new_n16313 = new_n16312 ^ new_n16311;
  assign new_n16314 = n127 & new_n2666;
  assign new_n16315 = n125 & new_n2664;
  assign new_n16316 = new_n16315 ^ new_n16314;
  assign new_n16317 = new_n16316 ^ new_n16313;
  assign new_n16318 = new_n16317 ^ n33;
  assign new_n16319 = ~new_n3143 & n123;
  assign new_n16320 = ~new_n9405 & new_n3138;
  assign new_n16321 = new_n16320 ^ new_n16319;
  assign new_n16322 = n124 & new_n3137;
  assign new_n16323 = n122 & new_n3149;
  assign new_n16324 = new_n16323 ^ new_n16322;
  assign new_n16325 = new_n16324 ^ new_n16321;
  assign new_n16326 = new_n16325 ^ n36;
  assign new_n16327 = ~new_n3682 & n120;
  assign new_n16328 = new_n3677 & new_n8560;
  assign new_n16329 = new_n16328 ^ new_n16327;
  assign new_n16330 = n121 & new_n3676;
  assign new_n16331 = n119 & new_n3688;
  assign new_n16332 = new_n16331 ^ new_n16330;
  assign new_n16333 = new_n16332 ^ new_n16329;
  assign new_n16334 = new_n16333 ^ n39;
  assign new_n16335 = ~new_n4212 & n117;
  assign new_n16336 = ~new_n7761 & new_n4201;
  assign new_n16337 = new_n16336 ^ new_n16335;
  assign new_n16338 = n118 & new_n4200;
  assign new_n16339 = n116 & new_n4206;
  assign new_n16340 = new_n16339 ^ new_n16338;
  assign new_n16341 = new_n16340 ^ new_n16337;
  assign new_n16342 = new_n16341 ^ n42;
  assign new_n16343 = ~new_n5424 & n111;
  assign new_n16344 = ~new_n6284 & new_n5419;
  assign new_n16345 = new_n16344 ^ new_n16343;
  assign new_n16346 = n112 & new_n5418;
  assign new_n16347 = n110 & new_n5648;
  assign new_n16348 = new_n16347 ^ new_n16346;
  assign new_n16349 = new_n16348 ^ new_n16345;
  assign new_n16350 = new_n16349 ^ n48;
  assign new_n16351 = ~new_n6110 & n108;
  assign new_n16352 = new_n5604 & new_n6105;
  assign new_n16353 = new_n16352 ^ new_n16351;
  assign new_n16354 = n109 & new_n6104;
  assign new_n16355 = n107 & new_n6347;
  assign new_n16356 = new_n16355 ^ new_n16354;
  assign new_n16357 = new_n16356 ^ new_n16353;
  assign new_n16358 = new_n16357 ^ n51;
  assign new_n16359 = new_n16234 ^ new_n16230;
  assign new_n16360 = ~new_n16231 & new_n16359;
  assign new_n16361 = new_n16360 ^ new_n16186;
  assign new_n16362 = new_n16361 ^ new_n16358;
  assign new_n16363 = ~new_n6805 & n105;
  assign new_n16364 = ~new_n4961 & new_n6800;
  assign new_n16365 = new_n16364 ^ new_n16363;
  assign new_n16366 = n106 & new_n6799;
  assign new_n16367 = n104 & new_n6811;
  assign new_n16368 = new_n16367 ^ new_n16366;
  assign new_n16369 = new_n16368 ^ new_n16365;
  assign new_n16370 = new_n16369 ^ n54;
  assign new_n16371 = new_n16229 ^ new_n16197;
  assign new_n16372 = new_n16198 & new_n16371;
  assign new_n16373 = new_n16372 ^ new_n16194;
  assign new_n16374 = new_n16373 ^ new_n16370;
  assign new_n16375 = n102 & new_n7553;
  assign new_n16376 = new_n4368 & new_n7543;
  assign new_n16377 = new_n16376 ^ new_n16375;
  assign new_n16378 = n103 & new_n7542;
  assign new_n16379 = n101 & new_n7547;
  assign new_n16380 = new_n16379 ^ new_n16378;
  assign new_n16381 = new_n16380 ^ new_n16377;
  assign new_n16382 = new_n16381 ^ n57;
  assign new_n16383 = new_n16228 ^ new_n16224;
  assign new_n16384 = ~new_n16225 & new_n16383;
  assign new_n16385 = new_n16384 ^ new_n16206;
  assign new_n16386 = new_n16385 ^ new_n16382;
  assign new_n16387 = n99 & new_n8355;
  assign new_n16388 = new_n3789 & new_n8345;
  assign new_n16389 = new_n16388 ^ new_n16387;
  assign new_n16390 = n100 & new_n8344;
  assign new_n16391 = n98 & new_n8349;
  assign new_n16392 = new_n16391 ^ new_n16390;
  assign new_n16393 = new_n16392 ^ new_n16389;
  assign new_n16394 = new_n16393 ^ n60;
  assign new_n16395 = new_n16222 ^ new_n16214;
  assign new_n16396 = new_n16223 & new_n16395;
  assign new_n16397 = new_n16396 ^ new_n16214;
  assign new_n16398 = new_n2499 ^ new_n2354;
  assign new_n16399 = new_n16398 ^ n64;
  assign new_n16400 = new_n16399 ^ new_n16398;
  assign new_n16401 = new_n16398 ^ new_n2499;
  assign new_n16402 = ~new_n16400 & new_n16401;
  assign new_n16403 = new_n16402 ^ new_n16398;
  assign new_n16404 = ~new_n9495 & new_n16403;
  assign new_n16405 = new_n16404 ^ new_n2499;
  assign new_n16406 = new_n16405 ^ new_n16397;
  assign new_n16407 = n96 & new_n9195;
  assign new_n16408 = new_n3273 & new_n9185;
  assign new_n16409 = new_n16408 ^ new_n16407;
  assign new_n16410 = n97 & new_n9184;
  assign new_n16411 = n95 & new_n9189;
  assign new_n16412 = new_n16411 ^ new_n16410;
  assign new_n16413 = new_n16412 ^ new_n16409;
  assign new_n16414 = new_n16413 ^ n63;
  assign new_n16415 = new_n16414 ^ new_n16406;
  assign new_n16416 = new_n16415 ^ new_n16394;
  assign new_n16417 = new_n16416 ^ new_n16386;
  assign new_n16418 = new_n16417 ^ new_n16374;
  assign new_n16419 = new_n16418 ^ new_n16362;
  assign new_n16420 = new_n16247 ^ new_n16235;
  assign new_n16421 = ~new_n16239 & new_n16420;
  assign new_n16422 = new_n16421 ^ new_n16238;
  assign new_n16423 = new_n16422 ^ new_n16419;
  assign new_n16424 = new_n16423 ^ new_n16350;
  assign new_n16425 = new_n16260 ^ new_n16248;
  assign new_n16426 = ~new_n16252 & new_n16425;
  assign new_n16427 = new_n16426 ^ new_n16251;
  assign new_n16428 = new_n16427 ^ new_n16424;
  assign new_n16429 = ~new_n4804 & n114;
  assign new_n16430 = ~new_n7013 & new_n4799;
  assign new_n16431 = new_n16430 ^ new_n16429;
  assign new_n16432 = n115 & new_n4798;
  assign new_n16433 = n113 & new_n4810;
  assign new_n16434 = new_n16433 ^ new_n16432;
  assign new_n16435 = new_n16434 ^ new_n16431;
  assign new_n16436 = new_n16435 ^ n45;
  assign new_n16437 = new_n16436 ^ new_n16428;
  assign new_n16438 = new_n16273 ^ new_n16261;
  assign new_n16439 = new_n16265 & new_n16438;
  assign new_n16440 = new_n16439 ^ new_n16264;
  assign new_n16441 = new_n16440 ^ new_n16437;
  assign new_n16442 = new_n16441 ^ new_n16342;
  assign new_n16443 = new_n16277 ^ new_n16178;
  assign new_n16444 = ~new_n16278 & new_n16443;
  assign new_n16445 = new_n16444 ^ new_n16178;
  assign new_n16446 = new_n16445 ^ new_n16442;
  assign new_n16447 = new_n16446 ^ new_n16334;
  assign new_n16448 = new_n16282 ^ new_n16170;
  assign new_n16449 = ~new_n16283 & new_n16448;
  assign new_n16450 = new_n16449 ^ new_n16170;
  assign new_n16451 = new_n16450 ^ new_n16447;
  assign new_n16452 = new_n16451 ^ new_n16326;
  assign new_n16453 = new_n16287 ^ new_n16162;
  assign new_n16454 = ~new_n16288 & new_n16453;
  assign new_n16455 = new_n16454 ^ new_n16162;
  assign new_n16456 = new_n16455 ^ new_n16452;
  assign new_n16457 = new_n16456 ^ new_n16318;
  assign new_n16458 = new_n16289 ^ new_n16154;
  assign new_n16459 = new_n16293 & new_n16458;
  assign new_n16460 = new_n16459 ^ new_n16154;
  assign new_n16461 = new_n16460 ^ new_n16457;
  assign new_n16462 = n128 & new_n2390;
  assign new_n16463 = ~n30 & ~new_n16462;
  assign new_n16464 = new_n16463 ^ n29;
  assign new_n16465 = new_n1980 & new_n11133;
  assign new_n16466 = new_n16465 ^ new_n16462;
  assign new_n16467 = ~new_n16464 & ~new_n16466;
  assign new_n16468 = new_n16467 ^ n29;
  assign new_n16469 = new_n16468 ^ new_n16461;
  assign new_n16470 = new_n16304 ^ new_n16294;
  assign new_n16471 = ~new_n16298 & new_n16470;
  assign new_n16472 = new_n16471 ^ new_n16297;
  assign new_n16473 = new_n16472 ^ new_n16469;
  assign new_n16474 = new_n16308 ^ new_n16146;
  assign new_n16475 = ~new_n16474 & new_n16309;
  assign new_n16476 = new_n16475 ^ new_n16146;
  assign new_n16477 = new_n16476 ^ new_n16473;
  assign new_n16478 = new_n16468 ^ new_n16457;
  assign new_n16479 = ~new_n16461 & new_n16478;
  assign new_n16480 = new_n16479 ^ new_n16468;
  assign new_n16481 = new_n16452 ^ new_n16318;
  assign new_n16482 = ~new_n16456 & new_n16481;
  assign new_n16483 = new_n16482 ^ new_n16318;
  assign new_n16484 = new_n16483 ^ new_n16480;
  assign new_n16485 = ~new_n2672 & n127;
  assign new_n16486 = new_n2667 & new_n10581;
  assign new_n16487 = new_n16486 ^ new_n16485;
  assign new_n16488 = n128 & new_n2666;
  assign new_n16489 = n126 & new_n2664;
  assign new_n16490 = new_n16489 ^ new_n16488;
  assign new_n16491 = new_n16490 ^ new_n16487;
  assign new_n16492 = new_n16491 ^ n33;
  assign new_n16493 = ~new_n3143 & n124;
  assign new_n16494 = new_n3138 & new_n9700;
  assign new_n16495 = new_n16494 ^ new_n16493;
  assign new_n16496 = n125 & new_n3137;
  assign new_n16497 = n123 & new_n3149;
  assign new_n16498 = new_n16497 ^ new_n16496;
  assign new_n16499 = new_n16498 ^ new_n16495;
  assign new_n16500 = new_n16499 ^ n36;
  assign new_n16501 = ~new_n4212 & n118;
  assign new_n16502 = ~new_n8019 & new_n4201;
  assign new_n16503 = new_n16502 ^ new_n16501;
  assign new_n16504 = n119 & new_n4200;
  assign new_n16505 = n117 & new_n4206;
  assign new_n16506 = new_n16505 ^ new_n16504;
  assign new_n16507 = new_n16506 ^ new_n16503;
  assign new_n16508 = new_n16507 ^ n42;
  assign new_n16509 = ~new_n4804 & n115;
  assign new_n16510 = ~new_n7256 & new_n4799;
  assign new_n16511 = new_n16510 ^ new_n16509;
  assign new_n16512 = n116 & new_n4798;
  assign new_n16513 = n114 & new_n4810;
  assign new_n16514 = new_n16513 ^ new_n16512;
  assign new_n16515 = new_n16514 ^ new_n16511;
  assign new_n16516 = new_n16515 ^ n45;
  assign new_n16517 = ~new_n5424 & n112;
  assign new_n16518 = ~new_n6518 & new_n5419;
  assign new_n16519 = new_n16518 ^ new_n16517;
  assign new_n16520 = n113 & new_n5418;
  assign new_n16521 = n111 & new_n5648;
  assign new_n16522 = new_n16521 ^ new_n16520;
  assign new_n16523 = new_n16522 ^ new_n16519;
  assign new_n16524 = new_n16523 ^ n48;
  assign new_n16525 = ~new_n6110 & n109;
  assign new_n16526 = new_n5825 & new_n6105;
  assign new_n16527 = new_n16526 ^ new_n16525;
  assign new_n16528 = n110 & new_n6104;
  assign new_n16529 = n108 & new_n6347;
  assign new_n16530 = new_n16529 ^ new_n16528;
  assign new_n16531 = new_n16530 ^ new_n16527;
  assign new_n16532 = new_n16531 ^ n51;
  assign new_n16533 = new_n16418 ^ new_n16361;
  assign new_n16534 = new_n16362 & new_n16533;
  assign new_n16535 = new_n16534 ^ new_n16358;
  assign new_n16536 = new_n16535 ^ new_n16532;
  assign new_n16537 = ~new_n6805 & n106;
  assign new_n16538 = ~new_n5164 & new_n6800;
  assign new_n16539 = new_n16538 ^ new_n16537;
  assign new_n16540 = n107 & new_n6799;
  assign new_n16541 = n105 & new_n6811;
  assign new_n16542 = new_n16541 ^ new_n16540;
  assign new_n16543 = new_n16542 ^ new_n16539;
  assign new_n16544 = new_n16543 ^ n54;
  assign new_n16545 = new_n16417 ^ new_n16373;
  assign new_n16546 = new_n16374 & new_n16545;
  assign new_n16547 = new_n16546 ^ new_n16370;
  assign new_n16548 = new_n16547 ^ new_n16544;
  assign new_n16549 = n103 & new_n7553;
  assign new_n16550 = ~new_n4556 & new_n7543;
  assign new_n16551 = new_n16550 ^ new_n16549;
  assign new_n16552 = n104 & new_n7542;
  assign new_n16553 = n102 & new_n7547;
  assign new_n16554 = new_n16553 ^ new_n16552;
  assign new_n16555 = new_n16554 ^ new_n16551;
  assign new_n16556 = new_n16555 ^ n57;
  assign new_n16557 = new_n16416 ^ new_n16385;
  assign new_n16558 = new_n16386 & new_n16557;
  assign new_n16559 = new_n16558 ^ new_n16382;
  assign new_n16560 = new_n16559 ^ new_n16556;
  assign new_n16561 = n100 & new_n8355;
  assign new_n16562 = new_n3972 & new_n8345;
  assign new_n16563 = new_n16562 ^ new_n16561;
  assign new_n16564 = n101 & new_n8344;
  assign new_n16565 = n99 & new_n8349;
  assign new_n16566 = new_n16565 ^ new_n16564;
  assign new_n16567 = new_n16566 ^ new_n16563;
  assign new_n16568 = new_n16567 ^ n60;
  assign new_n16569 = new_n16406 ^ new_n16394;
  assign new_n16570 = ~new_n16569 & new_n16415;
  assign new_n16571 = new_n16570 ^ new_n16394;
  assign new_n16572 = new_n16571 ^ new_n16568;
  assign new_n16573 = n97 & new_n9195;
  assign new_n16574 = new_n3435 & new_n9185;
  assign new_n16575 = new_n16574 ^ new_n16573;
  assign new_n16576 = n98 & new_n9184;
  assign new_n16577 = n96 & new_n9189;
  assign new_n16578 = new_n16577 ^ new_n16576;
  assign new_n16579 = new_n16578 ^ new_n16575;
  assign new_n16580 = new_n16579 ^ n63;
  assign new_n16581 = n95 ^ n93;
  assign new_n16582 = new_n11492 & new_n16581;
  assign new_n16583 = new_n16582 ^ n95;
  assign new_n16584 = new_n16583 ^ n94;
  assign new_n16585 = new_n11789 & new_n16584;
  assign new_n16586 = new_n16585 ^ n30;
  assign new_n16587 = new_n16586 ^ new_n16580;
  assign new_n16588 = ~n93 & n94;
  assign new_n16589 = ~n92 & n93;
  assign new_n16590 = n64 & new_n16589;
  assign new_n16591 = new_n16590 ^ new_n16588;
  assign new_n16592 = ~new_n9495 & new_n16591;
  assign new_n16593 = new_n16592 ^ new_n16588;
  assign new_n16594 = ~new_n16397 & ~new_n16405;
  assign new_n16595 = new_n16594 ^ new_n16593;
  assign new_n16596 = new_n16595 ^ new_n16587;
  assign new_n16597 = new_n16596 ^ new_n16572;
  assign new_n16598 = new_n16597 ^ new_n16560;
  assign new_n16599 = new_n16598 ^ new_n16548;
  assign new_n16600 = new_n16599 ^ new_n16536;
  assign new_n16601 = new_n16600 ^ new_n16524;
  assign new_n16602 = new_n16422 ^ new_n16350;
  assign new_n16603 = new_n16423 & new_n16602;
  assign new_n16604 = new_n16603 ^ new_n16350;
  assign new_n16605 = new_n16604 ^ new_n16601;
  assign new_n16606 = new_n16605 ^ new_n16516;
  assign new_n16607 = new_n16436 ^ new_n16424;
  assign new_n16608 = ~new_n16428 & new_n16607;
  assign new_n16609 = new_n16608 ^ new_n16427;
  assign new_n16610 = new_n16609 ^ new_n16606;
  assign new_n16611 = new_n16610 ^ new_n16508;
  assign new_n16612 = new_n16437 ^ new_n16342;
  assign new_n16613 = ~new_n16441 & ~new_n16612;
  assign new_n16614 = new_n16613 ^ new_n16342;
  assign new_n16615 = new_n16614 ^ new_n16611;
  assign new_n16616 = new_n16442 ^ new_n16334;
  assign new_n16617 = ~new_n16446 & new_n16616;
  assign new_n16618 = new_n16617 ^ new_n16334;
  assign new_n16619 = new_n16618 ^ new_n16615;
  assign new_n16620 = ~new_n3682 & n121;
  assign new_n16621 = new_n3677 & new_n8850;
  assign new_n16622 = new_n16621 ^ new_n16620;
  assign new_n16623 = n122 & new_n3676;
  assign new_n16624 = n120 & new_n3688;
  assign new_n16625 = new_n16624 ^ new_n16623;
  assign new_n16626 = new_n16625 ^ new_n16622;
  assign new_n16627 = new_n16626 ^ n39;
  assign new_n16628 = new_n16627 ^ new_n16619;
  assign new_n16629 = new_n16628 ^ new_n16500;
  assign new_n16630 = new_n16450 ^ new_n16326;
  assign new_n16631 = ~new_n16451 & new_n16630;
  assign new_n16632 = new_n16631 ^ new_n16326;
  assign new_n16633 = new_n16632 ^ new_n16629;
  assign new_n16634 = new_n16633 ^ new_n16492;
  assign new_n16635 = new_n16634 ^ new_n16484;
  assign new_n16636 = new_n16476 ^ new_n16472;
  assign new_n16637 = ~new_n16473 & ~new_n16636;
  assign new_n16638 = new_n16637 ^ new_n16476;
  assign new_n16639 = new_n16638 ^ new_n16635;
  assign new_n16640 = new_n16638 ^ new_n16484;
  assign new_n16641 = new_n16635 & new_n16640;
  assign new_n16642 = ~new_n16480 & ~new_n16483;
  assign new_n16643 = new_n16642 ^ new_n16484;
  assign new_n16644 = new_n16643 ^ new_n16641;
  assign new_n16645 = new_n16492 & new_n16633;
  assign new_n16646 = new_n16645 ^ new_n16634;
  assign new_n16647 = new_n16646 ^ new_n16644;
  assign new_n16648 = ~new_n3143 & n125;
  assign new_n16649 = new_n3138 & new_n9987;
  assign new_n16650 = new_n16649 ^ new_n16648;
  assign new_n16651 = n126 & new_n3137;
  assign new_n16652 = n124 & new_n3149;
  assign new_n16653 = new_n16652 ^ new_n16651;
  assign new_n16654 = new_n16653 ^ new_n16650;
  assign new_n16655 = new_n16654 ^ n36;
  assign new_n16656 = ~new_n3682 & n122;
  assign new_n16657 = ~new_n9116 & new_n3677;
  assign new_n16658 = new_n16657 ^ new_n16656;
  assign new_n16659 = n123 & new_n3676;
  assign new_n16660 = n121 & new_n3688;
  assign new_n16661 = new_n16660 ^ new_n16659;
  assign new_n16662 = new_n16661 ^ new_n16658;
  assign new_n16663 = new_n16662 ^ n39;
  assign new_n16664 = ~new_n4804 & n116;
  assign new_n16665 = ~new_n7503 & new_n4799;
  assign new_n16666 = new_n16665 ^ new_n16664;
  assign new_n16667 = n117 & new_n4798;
  assign new_n16668 = n115 & new_n4810;
  assign new_n16669 = new_n16668 ^ new_n16667;
  assign new_n16670 = new_n16669 ^ new_n16666;
  assign new_n16671 = new_n16670 ^ n45;
  assign new_n16672 = ~new_n5424 & n113;
  assign new_n16673 = ~new_n6764 & new_n5419;
  assign new_n16674 = new_n16673 ^ new_n16672;
  assign new_n16675 = n114 & new_n5418;
  assign new_n16676 = n112 & new_n5648;
  assign new_n16677 = new_n16676 ^ new_n16675;
  assign new_n16678 = new_n16677 ^ new_n16674;
  assign new_n16679 = new_n16678 ^ n48;
  assign new_n16680 = ~new_n6110 & n110;
  assign new_n16681 = new_n6049 & new_n6105;
  assign new_n16682 = new_n16681 ^ new_n16680;
  assign new_n16683 = n111 & new_n6104;
  assign new_n16684 = n109 & new_n6347;
  assign new_n16685 = new_n16684 ^ new_n16683;
  assign new_n16686 = new_n16685 ^ new_n16682;
  assign new_n16687 = new_n16686 ^ n51;
  assign new_n16688 = new_n16598 ^ new_n16544;
  assign new_n16689 = ~new_n16688 & new_n16548;
  assign new_n16690 = new_n16689 ^ new_n16547;
  assign new_n16691 = new_n16690 ^ new_n16687;
  assign new_n16692 = ~new_n6805 & n107;
  assign new_n16693 = ~new_n5377 & new_n6800;
  assign new_n16694 = new_n16693 ^ new_n16692;
  assign new_n16695 = n108 & new_n6799;
  assign new_n16696 = n106 & new_n6811;
  assign new_n16697 = new_n16696 ^ new_n16695;
  assign new_n16698 = new_n16697 ^ new_n16694;
  assign new_n16699 = new_n16698 ^ n54;
  assign new_n16700 = new_n16597 ^ new_n16556;
  assign new_n16701 = ~new_n16700 & new_n16560;
  assign new_n16702 = new_n16701 ^ new_n16559;
  assign new_n16703 = new_n16702 ^ new_n16699;
  assign new_n16704 = n104 & new_n7553;
  assign new_n16705 = ~new_n4754 & new_n7543;
  assign new_n16706 = new_n16705 ^ new_n16704;
  assign new_n16707 = n105 & new_n7542;
  assign new_n16708 = n103 & new_n7547;
  assign new_n16709 = new_n16708 ^ new_n16707;
  assign new_n16710 = new_n16709 ^ new_n16706;
  assign new_n16711 = new_n16710 ^ n57;
  assign new_n16712 = n101 & new_n8355;
  assign new_n16713 = new_n4159 & new_n8345;
  assign new_n16714 = new_n16713 ^ new_n16712;
  assign new_n16715 = n102 & new_n8344;
  assign new_n16716 = n100 & new_n8349;
  assign new_n16717 = new_n16716 ^ new_n16715;
  assign new_n16718 = new_n16717 ^ new_n16714;
  assign new_n16719 = new_n16718 ^ n60;
  assign new_n16720 = n96 & new_n9495;
  assign new_n16721 = n95 & new_n11492;
  assign new_n16722 = new_n16721 ^ new_n16720;
  assign new_n16723 = n98 & new_n9195;
  assign new_n16724 = new_n3604 & new_n9185;
  assign new_n16725 = new_n16724 ^ new_n16723;
  assign new_n16726 = n99 & new_n9184;
  assign new_n16727 = n97 & new_n9189;
  assign new_n16728 = new_n16727 ^ new_n16726;
  assign new_n16729 = new_n16728 ^ new_n16725;
  assign new_n16730 = new_n16729 ^ n63;
  assign new_n16731 = n94 ^ n30;
  assign new_n16732 = ~new_n16731 & new_n16584;
  assign new_n16733 = new_n16732 ^ n94;
  assign new_n16734 = new_n11789 & new_n16733;
  assign new_n16735 = new_n16734 ^ new_n16730;
  assign new_n16736 = new_n16735 ^ new_n16722;
  assign new_n16737 = new_n16736 ^ new_n16719;
  assign new_n16738 = new_n16595 ^ new_n16580;
  assign new_n16739 = ~new_n16738 & new_n16587;
  assign new_n16740 = new_n16739 ^ new_n16595;
  assign new_n16741 = new_n16740 ^ new_n16737;
  assign new_n16742 = new_n16741 ^ new_n16711;
  assign new_n16743 = new_n16596 ^ new_n16568;
  assign new_n16744 = ~new_n16743 & new_n16572;
  assign new_n16745 = new_n16744 ^ new_n16571;
  assign new_n16746 = new_n16745 ^ new_n16742;
  assign new_n16747 = new_n16746 ^ new_n16703;
  assign new_n16748 = new_n16747 ^ new_n16691;
  assign new_n16749 = new_n16599 ^ new_n16532;
  assign new_n16750 = ~new_n16749 & new_n16536;
  assign new_n16751 = new_n16750 ^ new_n16535;
  assign new_n16752 = new_n16751 ^ new_n16748;
  assign new_n16753 = new_n16752 ^ new_n16679;
  assign new_n16754 = new_n16604 ^ new_n16524;
  assign new_n16755 = ~new_n16601 & new_n16754;
  assign new_n16756 = new_n16755 ^ new_n16604;
  assign new_n16757 = new_n16756 ^ new_n16753;
  assign new_n16758 = new_n16757 ^ new_n16671;
  assign new_n16759 = new_n16609 ^ new_n16516;
  assign new_n16760 = ~new_n16606 & new_n16759;
  assign new_n16761 = new_n16760 ^ new_n16609;
  assign new_n16762 = new_n16761 ^ new_n16758;
  assign new_n16763 = ~new_n4212 & n119;
  assign new_n16764 = new_n4201 & new_n8286;
  assign new_n16765 = new_n16764 ^ new_n16763;
  assign new_n16766 = n120 & new_n4200;
  assign new_n16767 = n118 & new_n4206;
  assign new_n16768 = new_n16767 ^ new_n16766;
  assign new_n16769 = new_n16768 ^ new_n16765;
  assign new_n16770 = new_n16769 ^ n42;
  assign new_n16771 = new_n16770 ^ new_n16762;
  assign new_n16772 = new_n16614 ^ new_n16508;
  assign new_n16773 = ~new_n16611 & new_n16772;
  assign new_n16774 = new_n16773 ^ new_n16614;
  assign new_n16775 = new_n16774 ^ new_n16771;
  assign new_n16776 = new_n16775 ^ new_n16663;
  assign new_n16777 = new_n16627 ^ new_n16615;
  assign new_n16778 = ~new_n16777 & new_n16619;
  assign new_n16779 = new_n16778 ^ new_n16618;
  assign new_n16780 = new_n16779 ^ new_n16776;
  assign new_n16781 = new_n16780 ^ new_n16655;
  assign new_n16782 = new_n16632 ^ new_n16500;
  assign new_n16783 = ~new_n16629 & new_n16782;
  assign new_n16784 = new_n16783 ^ new_n16632;
  assign new_n16785 = new_n16784 ^ new_n16781;
  assign new_n16786 = n127 & new_n2664;
  assign new_n16787 = new_n2667 & new_n10010;
  assign new_n16788 = new_n16787 ^ new_n16786;
  assign new_n16789 = ~new_n2672 & n128;
  assign new_n16790 = new_n16789 ^ new_n16788;
  assign new_n16791 = new_n16790 ^ n33;
  assign new_n16792 = new_n16791 ^ new_n16785;
  assign new_n16793 = new_n16792 ^ new_n16647;
  assign new_n16794 = ~new_n16792 & new_n16643;
  assign new_n16795 = ~new_n16794 & new_n16646;
  assign new_n16796 = ~new_n16645 & ~new_n16792;
  assign new_n16797 = ~new_n16642 & ~new_n16796;
  assign new_n16798 = ~new_n16795 & ~new_n16797;
  assign new_n16799 = ~new_n16638 & ~new_n16798;
  assign new_n16800 = new_n16792 ^ new_n16645;
  assign new_n16801 = new_n16646 ^ new_n16483;
  assign new_n16802 = new_n16484 & new_n16801;
  assign new_n16803 = new_n16802 ^ new_n16483;
  assign new_n16804 = new_n16803 ^ new_n16643;
  assign new_n16805 = new_n16792 & new_n16804;
  assign new_n16806 = new_n16805 ^ new_n16643;
  assign new_n16807 = new_n16800 & new_n16806;
  assign new_n16808 = new_n16807 ^ new_n16645;
  assign new_n16809 = ~new_n16799 & ~new_n16808;
  assign new_n16810 = new_n2541 ^ n33;
  assign new_n16811 = new_n2542 ^ new_n2541;
  assign new_n16812 = new_n2661 ^ new_n2542;
  assign new_n16813 = new_n2542 & new_n16812;
  assign new_n16814 = new_n16813 ^ new_n2542;
  assign new_n16815 = ~new_n16811 & new_n16814;
  assign new_n16816 = new_n16815 ^ new_n16813;
  assign new_n16817 = new_n16816 ^ new_n2542;
  assign new_n16818 = new_n16817 ^ new_n2661;
  assign new_n16819 = ~new_n16810 & new_n16818;
  assign new_n16820 = new_n16819 ^ n33;
  assign new_n16821 = new_n16820 ^ n33;
  assign new_n16822 = new_n16810 & new_n16818;
  assign new_n16823 = new_n16822 ^ n32;
  assign new_n16824 = new_n16823 ^ n33;
  assign new_n16825 = new_n16824 ^ new_n16821;
  assign new_n16826 = new_n16824 ^ new_n10009;
  assign new_n16827 = new_n16826 ^ new_n16824;
  assign new_n16828 = new_n16825 & new_n16827;
  assign new_n16829 = new_n16828 ^ new_n16824;
  assign new_n16830 = n128 & new_n16829;
  assign new_n16831 = new_n16830 ^ n33;
  assign new_n16832 = ~new_n3143 & n126;
  assign new_n16833 = new_n3138 & new_n10304;
  assign new_n16834 = new_n16833 ^ new_n16832;
  assign new_n16835 = n127 & new_n3137;
  assign new_n16836 = n125 & new_n3149;
  assign new_n16837 = new_n16836 ^ new_n16835;
  assign new_n16838 = new_n16837 ^ new_n16834;
  assign new_n16839 = new_n16838 ^ n36;
  assign new_n16840 = ~new_n3682 & n123;
  assign new_n16841 = ~new_n9405 & new_n3677;
  assign new_n16842 = new_n16841 ^ new_n16840;
  assign new_n16843 = n124 & new_n3676;
  assign new_n16844 = n122 & new_n3688;
  assign new_n16845 = new_n16844 ^ new_n16843;
  assign new_n16846 = new_n16845 ^ new_n16842;
  assign new_n16847 = new_n16846 ^ n39;
  assign new_n16848 = ~new_n4212 & n120;
  assign new_n16849 = new_n4201 & new_n8560;
  assign new_n16850 = new_n16849 ^ new_n16848;
  assign new_n16851 = n121 & new_n4200;
  assign new_n16852 = n119 & new_n4206;
  assign new_n16853 = new_n16852 ^ new_n16851;
  assign new_n16854 = new_n16853 ^ new_n16850;
  assign new_n16855 = new_n16854 ^ n42;
  assign new_n16856 = ~new_n4804 & n117;
  assign new_n16857 = ~new_n7761 & new_n4799;
  assign new_n16858 = new_n16857 ^ new_n16856;
  assign new_n16859 = n118 & new_n4798;
  assign new_n16860 = n116 & new_n4810;
  assign new_n16861 = new_n16860 ^ new_n16859;
  assign new_n16862 = new_n16861 ^ new_n16858;
  assign new_n16863 = new_n16862 ^ n45;
  assign new_n16864 = ~new_n5424 & n114;
  assign new_n16865 = ~new_n7013 & new_n5419;
  assign new_n16866 = new_n16865 ^ new_n16864;
  assign new_n16867 = n115 & new_n5418;
  assign new_n16868 = n113 & new_n5648;
  assign new_n16869 = new_n16868 ^ new_n16867;
  assign new_n16870 = new_n16869 ^ new_n16866;
  assign new_n16871 = new_n16870 ^ n48;
  assign new_n16872 = ~new_n6110 & n111;
  assign new_n16873 = ~new_n6284 & new_n6105;
  assign new_n16874 = new_n16873 ^ new_n16872;
  assign new_n16875 = n112 & new_n6104;
  assign new_n16876 = n110 & new_n6347;
  assign new_n16877 = new_n16876 ^ new_n16875;
  assign new_n16878 = new_n16877 ^ new_n16874;
  assign new_n16879 = new_n16878 ^ n51;
  assign new_n16880 = ~new_n6805 & n108;
  assign new_n16881 = new_n5604 & new_n6800;
  assign new_n16882 = new_n16881 ^ new_n16880;
  assign new_n16883 = n109 & new_n6799;
  assign new_n16884 = n107 & new_n6811;
  assign new_n16885 = new_n16884 ^ new_n16883;
  assign new_n16886 = new_n16885 ^ new_n16882;
  assign new_n16887 = new_n16886 ^ n54;
  assign new_n16888 = new_n16745 ^ new_n16741;
  assign new_n16889 = ~new_n16888 & new_n16742;
  assign new_n16890 = new_n16889 ^ new_n16711;
  assign new_n16891 = new_n16890 ^ new_n16887;
  assign new_n16892 = n105 & new_n7553;
  assign new_n16893 = ~new_n4961 & new_n7543;
  assign new_n16894 = new_n16893 ^ new_n16892;
  assign new_n16895 = n106 & new_n7542;
  assign new_n16896 = n104 & new_n7547;
  assign new_n16897 = new_n16896 ^ new_n16895;
  assign new_n16898 = new_n16897 ^ new_n16894;
  assign new_n16899 = new_n16898 ^ n57;
  assign new_n16900 = new_n16740 ^ new_n16736;
  assign new_n16901 = ~new_n16737 & ~new_n16900;
  assign new_n16902 = new_n16901 ^ new_n16719;
  assign new_n16903 = new_n16902 ^ new_n16899;
  assign new_n16904 = ~n97 & new_n9495;
  assign new_n16905 = new_n16904 ^ new_n16721;
  assign new_n16906 = n96 & new_n16905;
  assign new_n16907 = new_n16906 ^ new_n16721;
  assign new_n16908 = new_n9495 ^ n96;
  assign new_n16909 = new_n11789 ^ n95;
  assign new_n16910 = new_n16909 ^ new_n16905;
  assign new_n16911 = new_n16910 ^ n95;
  assign new_n16912 = new_n16908 & new_n16911;
  assign new_n16913 = new_n16912 ^ new_n2947;
  assign new_n16914 = new_n16913 ^ new_n16907;
  assign new_n16915 = new_n16914 ^ new_n2947;
  assign new_n16916 = new_n16734 ^ new_n16722;
  assign new_n16917 = new_n16735 & new_n16916;
  assign new_n16918 = new_n16917 ^ new_n16730;
  assign new_n16919 = new_n16918 ^ new_n16915;
  assign new_n16920 = n99 & new_n9195;
  assign new_n16921 = new_n3789 & new_n9185;
  assign new_n16922 = new_n16921 ^ new_n16920;
  assign new_n16923 = n100 & new_n9184;
  assign new_n16924 = n98 & new_n9189;
  assign new_n16925 = new_n16924 ^ new_n16923;
  assign new_n16926 = new_n16925 ^ new_n16922;
  assign new_n16927 = new_n16926 ^ n63;
  assign new_n16928 = new_n16927 ^ new_n16919;
  assign new_n16929 = n102 & new_n8355;
  assign new_n16930 = new_n4368 & new_n8345;
  assign new_n16931 = new_n16930 ^ new_n16929;
  assign new_n16932 = n103 & new_n8344;
  assign new_n16933 = n101 & new_n8349;
  assign new_n16934 = new_n16933 ^ new_n16932;
  assign new_n16935 = new_n16934 ^ new_n16931;
  assign new_n16936 = new_n16935 ^ n60;
  assign new_n16937 = new_n16936 ^ new_n16928;
  assign new_n16938 = new_n16937 ^ new_n16903;
  assign new_n16939 = new_n16938 ^ new_n16891;
  assign new_n16940 = new_n16746 ^ new_n16699;
  assign new_n16941 = ~new_n16940 & new_n16703;
  assign new_n16942 = new_n16941 ^ new_n16702;
  assign new_n16943 = new_n16942 ^ new_n16939;
  assign new_n16944 = new_n16943 ^ new_n16879;
  assign new_n16945 = new_n16747 ^ new_n16687;
  assign new_n16946 = ~new_n16945 & new_n16691;
  assign new_n16947 = new_n16946 ^ new_n16690;
  assign new_n16948 = new_n16947 ^ new_n16944;
  assign new_n16949 = new_n16948 ^ new_n16871;
  assign new_n16950 = new_n16748 ^ new_n16679;
  assign new_n16951 = ~new_n16752 & new_n16950;
  assign new_n16952 = new_n16951 ^ new_n16679;
  assign new_n16953 = new_n16952 ^ new_n16949;
  assign new_n16954 = new_n16953 ^ new_n16863;
  assign new_n16955 = new_n16756 ^ new_n16671;
  assign new_n16956 = ~new_n16757 & new_n16955;
  assign new_n16957 = new_n16956 ^ new_n16671;
  assign new_n16958 = new_n16957 ^ new_n16954;
  assign new_n16959 = new_n16958 ^ new_n16855;
  assign new_n16960 = new_n16770 ^ new_n16758;
  assign new_n16961 = ~new_n16960 & new_n16762;
  assign new_n16962 = new_n16961 ^ new_n16761;
  assign new_n16963 = new_n16962 ^ new_n16959;
  assign new_n16964 = new_n16963 ^ new_n16847;
  assign new_n16965 = new_n16774 ^ new_n16663;
  assign new_n16966 = ~new_n16775 & new_n16965;
  assign new_n16967 = new_n16966 ^ new_n16663;
  assign new_n16968 = new_n16967 ^ new_n16964;
  assign new_n16969 = new_n16968 ^ new_n16839;
  assign new_n16970 = new_n16969 ^ new_n16831;
  assign new_n16971 = new_n16779 ^ new_n16655;
  assign new_n16972 = ~new_n16780 & new_n16971;
  assign new_n16973 = new_n16972 ^ new_n16655;
  assign new_n16974 = new_n16973 ^ new_n16970;
  assign new_n16975 = new_n16791 ^ new_n16781;
  assign new_n16976 = ~new_n16975 & new_n16785;
  assign new_n16977 = new_n16976 ^ new_n16784;
  assign new_n16978 = new_n16977 ^ new_n16974;
  assign new_n16979 = new_n16978 ^ new_n16809;
  assign new_n16980 = ~new_n3143 & n127;
  assign new_n16981 = new_n3138 & new_n10581;
  assign new_n16982 = new_n16981 ^ new_n16980;
  assign new_n16983 = n128 & new_n3137;
  assign new_n16984 = n126 & new_n3149;
  assign new_n16985 = new_n16984 ^ new_n16983;
  assign new_n16986 = new_n16985 ^ new_n16982;
  assign new_n16987 = new_n16986 ^ n36;
  assign new_n16988 = ~new_n3682 & n124;
  assign new_n16989 = new_n3677 & new_n9700;
  assign new_n16990 = new_n16989 ^ new_n16988;
  assign new_n16991 = n125 & new_n3676;
  assign new_n16992 = n123 & new_n3688;
  assign new_n16993 = new_n16992 ^ new_n16991;
  assign new_n16994 = new_n16993 ^ new_n16990;
  assign new_n16995 = new_n16994 ^ n39;
  assign new_n16996 = ~new_n6110 & n112;
  assign new_n16997 = ~new_n6518 & new_n6105;
  assign new_n16998 = new_n16997 ^ new_n16996;
  assign new_n16999 = n113 & new_n6104;
  assign new_n17000 = n111 & new_n6347;
  assign new_n17001 = new_n17000 ^ new_n16999;
  assign new_n17002 = new_n17001 ^ new_n16998;
  assign new_n17003 = new_n17002 ^ n51;
  assign new_n17004 = new_n16942 ^ new_n16879;
  assign new_n17005 = new_n16943 & new_n17004;
  assign new_n17006 = new_n17005 ^ new_n16879;
  assign new_n17007 = new_n17006 ^ new_n17003;
  assign new_n17008 = ~new_n6805 & n109;
  assign new_n17009 = new_n5825 & new_n6800;
  assign new_n17010 = new_n17009 ^ new_n17008;
  assign new_n17011 = n110 & new_n6799;
  assign new_n17012 = n108 & new_n6811;
  assign new_n17013 = new_n17012 ^ new_n17011;
  assign new_n17014 = new_n17013 ^ new_n17010;
  assign new_n17015 = new_n17014 ^ n54;
  assign new_n17016 = new_n16938 ^ new_n16887;
  assign new_n17017 = new_n16891 & new_n17016;
  assign new_n17018 = new_n17017 ^ new_n16890;
  assign new_n17019 = new_n17018 ^ new_n17015;
  assign new_n17020 = n106 & new_n7553;
  assign new_n17021 = ~new_n5164 & new_n7543;
  assign new_n17022 = new_n17021 ^ new_n17020;
  assign new_n17023 = n107 & new_n7542;
  assign new_n17024 = n105 & new_n7547;
  assign new_n17025 = new_n17024 ^ new_n17023;
  assign new_n17026 = new_n17025 ^ new_n17022;
  assign new_n17027 = new_n17026 ^ n57;
  assign new_n17028 = new_n16937 ^ new_n16902;
  assign new_n17029 = new_n16903 & new_n17028;
  assign new_n17030 = new_n17029 ^ new_n16899;
  assign new_n17031 = new_n17030 ^ new_n17027;
  assign new_n17032 = n103 & new_n8355;
  assign new_n17033 = ~new_n4556 & new_n8345;
  assign new_n17034 = new_n17033 ^ new_n17032;
  assign new_n17035 = n104 & new_n8344;
  assign new_n17036 = n102 & new_n8349;
  assign new_n17037 = new_n17036 ^ new_n17035;
  assign new_n17038 = new_n17037 ^ new_n17034;
  assign new_n17039 = new_n17038 ^ n60;
  assign new_n17040 = new_n16936 ^ new_n16927;
  assign new_n17041 = ~new_n16928 & ~new_n17040;
  assign new_n17042 = new_n17041 ^ new_n16919;
  assign new_n17043 = new_n17042 ^ new_n17039;
  assign new_n17044 = ~new_n16907 & ~new_n16918;
  assign new_n17045 = ~new_n16912 & ~new_n17044;
  assign new_n17046 = n100 & new_n9195;
  assign new_n17047 = new_n3972 & new_n9185;
  assign new_n17048 = new_n17047 ^ new_n17046;
  assign new_n17049 = n101 & new_n9184;
  assign new_n17050 = n99 & new_n9189;
  assign new_n17051 = new_n17050 ^ new_n17049;
  assign new_n17052 = new_n17051 ^ new_n17048;
  assign new_n17053 = new_n17052 ^ n63;
  assign new_n17054 = n98 ^ n96;
  assign new_n17055 = ~new_n11492 & new_n17054;
  assign new_n17056 = new_n17055 ^ n96;
  assign new_n17057 = new_n17056 ^ n97;
  assign new_n17058 = new_n11789 & new_n17057;
  assign new_n17059 = new_n17058 ^ n33;
  assign new_n17060 = new_n17059 ^ new_n17053;
  assign new_n17061 = new_n17060 ^ new_n17045;
  assign new_n17062 = new_n17061 ^ new_n17043;
  assign new_n17063 = new_n17062 ^ new_n17031;
  assign new_n17064 = new_n17063 ^ new_n17019;
  assign new_n17065 = new_n17064 ^ new_n17007;
  assign new_n17066 = ~new_n5424 & n115;
  assign new_n17067 = ~new_n7256 & new_n5419;
  assign new_n17068 = new_n17067 ^ new_n17066;
  assign new_n17069 = n116 & new_n5418;
  assign new_n17070 = n114 & new_n5648;
  assign new_n17071 = new_n17070 ^ new_n17069;
  assign new_n17072 = new_n17071 ^ new_n17068;
  assign new_n17073 = new_n17072 ^ n48;
  assign new_n17074 = new_n17073 ^ new_n17065;
  assign new_n17075 = new_n16947 ^ new_n16871;
  assign new_n17076 = new_n16948 & new_n17075;
  assign new_n17077 = new_n17076 ^ new_n16871;
  assign new_n17078 = new_n17077 ^ new_n17074;
  assign new_n17079 = new_n16949 ^ new_n16863;
  assign new_n17080 = ~new_n17079 & new_n16953;
  assign new_n17081 = new_n17080 ^ new_n16863;
  assign new_n17082 = new_n17081 ^ new_n17078;
  assign new_n17083 = ~new_n4804 & n118;
  assign new_n17084 = ~new_n8019 & new_n4799;
  assign new_n17085 = new_n17084 ^ new_n17083;
  assign new_n17086 = n119 & new_n4798;
  assign new_n17087 = n117 & new_n4810;
  assign new_n17088 = new_n17087 ^ new_n17086;
  assign new_n17089 = new_n17088 ^ new_n17085;
  assign new_n17090 = new_n17089 ^ n45;
  assign new_n17091 = new_n17090 ^ new_n17082;
  assign new_n17092 = new_n16954 ^ new_n16855;
  assign new_n17093 = ~new_n17092 & new_n16958;
  assign new_n17094 = new_n17093 ^ new_n16855;
  assign new_n17095 = new_n17094 ^ new_n17091;
  assign new_n17096 = ~new_n4212 & n121;
  assign new_n17097 = new_n4201 & new_n8850;
  assign new_n17098 = new_n17097 ^ new_n17096;
  assign new_n17099 = n122 & new_n4200;
  assign new_n17100 = n120 & new_n4206;
  assign new_n17101 = new_n17100 ^ new_n17099;
  assign new_n17102 = new_n17101 ^ new_n17098;
  assign new_n17103 = new_n17102 ^ n42;
  assign new_n17104 = new_n17103 ^ new_n17095;
  assign new_n17105 = new_n17104 ^ new_n16995;
  assign new_n17106 = new_n16962 ^ new_n16847;
  assign new_n17107 = new_n16963 & new_n17106;
  assign new_n17108 = new_n17107 ^ new_n16847;
  assign new_n17109 = new_n17108 ^ new_n17105;
  assign new_n17110 = new_n17109 ^ new_n16987;
  assign new_n17111 = new_n16964 ^ new_n16839;
  assign new_n17112 = ~new_n17111 & new_n16968;
  assign new_n17113 = new_n17112 ^ new_n16839;
  assign new_n17114 = new_n17113 ^ new_n17110;
  assign new_n17115 = new_n16973 ^ new_n16969;
  assign new_n17116 = ~new_n16970 & new_n17115;
  assign new_n17117 = new_n17116 ^ new_n16831;
  assign new_n17118 = new_n17117 ^ new_n17114;
  assign new_n17119 = new_n16977 ^ new_n16809;
  assign new_n17120 = ~new_n17119 & new_n16978;
  assign new_n17121 = new_n17120 ^ new_n16809;
  assign new_n17122 = new_n17121 ^ new_n17118;
  assign new_n17123 = ~new_n3682 & n125;
  assign new_n17124 = new_n3677 & new_n9987;
  assign new_n17125 = new_n17124 ^ new_n17123;
  assign new_n17126 = n126 & new_n3676;
  assign new_n17127 = n124 & new_n3688;
  assign new_n17128 = new_n17127 ^ new_n17126;
  assign new_n17129 = new_n17128 ^ new_n17125;
  assign new_n17130 = new_n17129 ^ n39;
  assign new_n17131 = ~new_n4212 & n122;
  assign new_n17132 = ~new_n9116 & new_n4201;
  assign new_n17133 = new_n17132 ^ new_n17131;
  assign new_n17134 = n123 & new_n4200;
  assign new_n17135 = n121 & new_n4206;
  assign new_n17136 = new_n17135 ^ new_n17134;
  assign new_n17137 = new_n17136 ^ new_n17133;
  assign new_n17138 = new_n17137 ^ n42;
  assign new_n17139 = ~new_n5424 & n116;
  assign new_n17140 = ~new_n7503 & new_n5419;
  assign new_n17141 = new_n17140 ^ new_n17139;
  assign new_n17142 = n117 & new_n5418;
  assign new_n17143 = n115 & new_n5648;
  assign new_n17144 = new_n17143 ^ new_n17142;
  assign new_n17145 = new_n17144 ^ new_n17141;
  assign new_n17146 = new_n17145 ^ n48;
  assign new_n17147 = ~new_n6110 & n113;
  assign new_n17148 = ~new_n6764 & new_n6105;
  assign new_n17149 = new_n17148 ^ new_n17147;
  assign new_n17150 = n114 & new_n6104;
  assign new_n17151 = n112 & new_n6347;
  assign new_n17152 = new_n17151 ^ new_n17150;
  assign new_n17153 = new_n17152 ^ new_n17149;
  assign new_n17154 = new_n17153 ^ n51;
  assign new_n17155 = new_n17063 ^ new_n17015;
  assign new_n17156 = ~new_n17155 & new_n17019;
  assign new_n17157 = new_n17156 ^ new_n17018;
  assign new_n17158 = new_n17157 ^ new_n17154;
  assign new_n17159 = ~new_n6805 & n110;
  assign new_n17160 = new_n6049 & new_n6800;
  assign new_n17161 = new_n17160 ^ new_n17159;
  assign new_n17162 = n111 & new_n6799;
  assign new_n17163 = n109 & new_n6811;
  assign new_n17164 = new_n17163 ^ new_n17162;
  assign new_n17165 = new_n17164 ^ new_n17161;
  assign new_n17166 = new_n17165 ^ n54;
  assign new_n17167 = new_n17062 ^ new_n17027;
  assign new_n17168 = ~new_n17167 & new_n17031;
  assign new_n17169 = new_n17168 ^ new_n17030;
  assign new_n17170 = new_n17169 ^ new_n17166;
  assign new_n17171 = n107 & new_n7553;
  assign new_n17172 = ~new_n5377 & new_n7543;
  assign new_n17173 = new_n17172 ^ new_n17171;
  assign new_n17174 = n108 & new_n7542;
  assign new_n17175 = n106 & new_n7547;
  assign new_n17176 = new_n17175 ^ new_n17174;
  assign new_n17177 = new_n17176 ^ new_n17173;
  assign new_n17178 = new_n17177 ^ n57;
  assign new_n17179 = new_n17061 ^ new_n17042;
  assign new_n17180 = ~new_n17043 & ~new_n17179;
  assign new_n17181 = new_n17180 ^ new_n17039;
  assign new_n17182 = new_n17181 ^ new_n17178;
  assign new_n17183 = n104 & new_n8355;
  assign new_n17184 = ~new_n4754 & new_n8345;
  assign new_n17185 = new_n17184 ^ new_n17183;
  assign new_n17186 = n105 & new_n8344;
  assign new_n17187 = n103 & new_n8349;
  assign new_n17188 = new_n17187 ^ new_n17186;
  assign new_n17189 = new_n17188 ^ new_n17185;
  assign new_n17190 = new_n17189 ^ n60;
  assign new_n17191 = n98 & new_n11492;
  assign new_n17192 = n99 & new_n9495;
  assign new_n17193 = new_n17192 ^ new_n17191;
  assign new_n17194 = n101 & new_n9195;
  assign new_n17195 = new_n4159 & new_n9185;
  assign new_n17196 = new_n17195 ^ new_n17194;
  assign new_n17197 = n102 & new_n9184;
  assign new_n17198 = n100 & new_n9189;
  assign new_n17199 = new_n17198 ^ new_n17197;
  assign new_n17200 = new_n17199 ^ new_n17196;
  assign new_n17201 = new_n17200 ^ n63;
  assign new_n17202 = n97 ^ n33;
  assign new_n17203 = ~new_n17202 & new_n17057;
  assign new_n17204 = new_n17203 ^ n97;
  assign new_n17205 = new_n11789 & new_n17204;
  assign new_n17206 = new_n17205 ^ new_n17201;
  assign new_n17207 = new_n17206 ^ new_n17193;
  assign new_n17208 = new_n17207 ^ new_n17190;
  assign new_n17209 = new_n17053 ^ new_n17045;
  assign new_n17210 = new_n17060 & new_n17209;
  assign new_n17211 = new_n17210 ^ new_n17045;
  assign new_n17212 = new_n17211 ^ new_n17208;
  assign new_n17213 = new_n17212 ^ new_n17182;
  assign new_n17214 = new_n17213 ^ new_n17170;
  assign new_n17215 = new_n17214 ^ new_n17158;
  assign new_n17216 = new_n17215 ^ new_n17146;
  assign new_n17217 = new_n17064 ^ new_n17003;
  assign new_n17218 = ~new_n17217 & new_n17007;
  assign new_n17219 = new_n17218 ^ new_n17006;
  assign new_n17220 = new_n17219 ^ new_n17216;
  assign new_n17221 = new_n17077 ^ new_n17073;
  assign new_n17222 = ~new_n17221 & new_n17074;
  assign new_n17223 = new_n17222 ^ new_n17065;
  assign new_n17224 = new_n17223 ^ new_n17220;
  assign new_n17225 = ~new_n4804 & n119;
  assign new_n17226 = new_n4799 & new_n8286;
  assign new_n17227 = new_n17226 ^ new_n17225;
  assign new_n17228 = n120 & new_n4798;
  assign new_n17229 = n118 & new_n4810;
  assign new_n17230 = new_n17229 ^ new_n17228;
  assign new_n17231 = new_n17230 ^ new_n17227;
  assign new_n17232 = new_n17231 ^ n45;
  assign new_n17233 = new_n17232 ^ new_n17224;
  assign new_n17234 = new_n17090 ^ new_n17078;
  assign new_n17235 = ~new_n17234 & new_n17082;
  assign new_n17236 = new_n17235 ^ new_n17081;
  assign new_n17237 = new_n17236 ^ new_n17233;
  assign new_n17238 = new_n17237 ^ new_n17138;
  assign new_n17239 = new_n17103 ^ new_n17091;
  assign new_n17240 = ~new_n17239 & new_n17095;
  assign new_n17241 = new_n17240 ^ new_n17094;
  assign new_n17242 = new_n17241 ^ new_n17238;
  assign new_n17243 = new_n17242 ^ new_n17130;
  assign new_n17244 = n127 & new_n3149;
  assign new_n17245 = new_n3138 & new_n10010;
  assign new_n17246 = new_n17245 ^ new_n17244;
  assign new_n17247 = ~new_n3143 & n128;
  assign new_n17248 = new_n17247 ^ new_n17246;
  assign new_n17249 = new_n17248 ^ n36;
  assign new_n17250 = new_n17249 ^ new_n17243;
  assign new_n17251 = ~new_n17243 & new_n17249;
  assign new_n17252 = new_n17251 ^ new_n17250;
  assign new_n17253 = new_n17108 ^ new_n16995;
  assign new_n17254 = ~new_n17105 & new_n17253;
  assign new_n17255 = new_n17254 ^ new_n17108;
  assign new_n17256 = new_n17113 ^ new_n17109;
  assign new_n17257 = ~new_n17256 & new_n17110;
  assign new_n17258 = new_n17257 ^ new_n16987;
  assign new_n17259 = new_n17258 ^ new_n17255;
  assign new_n17260 = ~new_n17255 & ~new_n17258;
  assign new_n17261 = new_n17260 ^ new_n17259;
  assign new_n17262 = new_n17261 ^ new_n17252;
  assign new_n17263 = new_n17260 ^ new_n17251;
  assign new_n17264 = new_n17263 ^ new_n17262;
  assign new_n17265 = new_n17121 ^ new_n17117;
  assign new_n17266 = ~new_n17118 & ~new_n17265;
  assign new_n17267 = new_n17266 ^ new_n17121;
  assign new_n17268 = new_n17267 ^ new_n17264;
  assign new_n17269 = new_n17267 ^ new_n17255;
  assign new_n17270 = new_n17269 ^ new_n17258;
  assign new_n17271 = ~new_n17264 & ~new_n17270;
  assign new_n17272 = new_n17271 ^ new_n17263;
  assign new_n17273 = ~new_n3682 & n126;
  assign new_n17274 = new_n3677 & new_n10304;
  assign new_n17275 = new_n17274 ^ new_n17273;
  assign new_n17276 = n127 & new_n3676;
  assign new_n17277 = n125 & new_n3688;
  assign new_n17278 = new_n17277 ^ new_n17276;
  assign new_n17279 = new_n17278 ^ new_n17275;
  assign new_n17280 = new_n17279 ^ n39;
  assign new_n17281 = ~new_n4212 & n123;
  assign new_n17282 = ~new_n9405 & new_n4201;
  assign new_n17283 = new_n17282 ^ new_n17281;
  assign new_n17284 = n124 & new_n4200;
  assign new_n17285 = n122 & new_n4206;
  assign new_n17286 = new_n17285 ^ new_n17284;
  assign new_n17287 = new_n17286 ^ new_n17283;
  assign new_n17288 = new_n17287 ^ n42;
  assign new_n17289 = ~new_n5424 & n117;
  assign new_n17290 = ~new_n7761 & new_n5419;
  assign new_n17291 = new_n17290 ^ new_n17289;
  assign new_n17292 = n118 & new_n5418;
  assign new_n17293 = n116 & new_n5648;
  assign new_n17294 = new_n17293 ^ new_n17292;
  assign new_n17295 = new_n17294 ^ new_n17291;
  assign new_n17296 = new_n17295 ^ n48;
  assign new_n17297 = ~new_n6110 & n114;
  assign new_n17298 = ~new_n7013 & new_n6105;
  assign new_n17299 = new_n17298 ^ new_n17297;
  assign new_n17300 = n115 & new_n6104;
  assign new_n17301 = n113 & new_n6347;
  assign new_n17302 = new_n17301 ^ new_n17300;
  assign new_n17303 = new_n17302 ^ new_n17299;
  assign new_n17304 = new_n17303 ^ n51;
  assign new_n17305 = new_n17213 ^ new_n17166;
  assign new_n17306 = new_n17170 & new_n17305;
  assign new_n17307 = new_n17306 ^ new_n17169;
  assign new_n17308 = new_n17307 ^ new_n17304;
  assign new_n17309 = ~new_n6805 & n111;
  assign new_n17310 = ~new_n6284 & new_n6800;
  assign new_n17311 = new_n17310 ^ new_n17309;
  assign new_n17312 = n112 & new_n6799;
  assign new_n17313 = n110 & new_n6811;
  assign new_n17314 = new_n17313 ^ new_n17312;
  assign new_n17315 = new_n17314 ^ new_n17311;
  assign new_n17316 = new_n17315 ^ n54;
  assign new_n17317 = new_n17212 ^ new_n17181;
  assign new_n17318 = new_n17182 & new_n17317;
  assign new_n17319 = new_n17318 ^ new_n17178;
  assign new_n17320 = new_n17319 ^ new_n17316;
  assign new_n17321 = n108 & new_n7553;
  assign new_n17322 = new_n5604 & new_n7543;
  assign new_n17323 = new_n17322 ^ new_n17321;
  assign new_n17324 = n109 & new_n7542;
  assign new_n17325 = n107 & new_n7547;
  assign new_n17326 = new_n17325 ^ new_n17324;
  assign new_n17327 = new_n17326 ^ new_n17323;
  assign new_n17328 = new_n17327 ^ n57;
  assign new_n17329 = new_n17211 ^ new_n17207;
  assign new_n17330 = ~new_n17208 & new_n17329;
  assign new_n17331 = new_n17330 ^ new_n17190;
  assign new_n17332 = new_n17331 ^ new_n17328;
  assign new_n17333 = n105 & new_n8355;
  assign new_n17334 = ~new_n4961 & new_n8345;
  assign new_n17335 = new_n17334 ^ new_n17333;
  assign new_n17336 = n106 & new_n8344;
  assign new_n17337 = n104 & new_n8349;
  assign new_n17338 = new_n17337 ^ new_n17336;
  assign new_n17339 = new_n17338 ^ new_n17335;
  assign new_n17340 = new_n17339 ^ n60;
  assign new_n17341 = new_n17205 ^ new_n17193;
  assign new_n17342 = new_n17206 & new_n17341;
  assign new_n17343 = new_n17342 ^ new_n17201;
  assign new_n17344 = ~n100 & new_n9495;
  assign new_n17345 = new_n17344 ^ new_n17191;
  assign new_n17346 = n99 & new_n17345;
  assign new_n17347 = new_n17346 ^ new_n17191;
  assign new_n17348 = new_n9495 ^ n99;
  assign new_n17349 = new_n11789 ^ n98;
  assign new_n17350 = new_n17349 ^ new_n17345;
  assign new_n17351 = new_n17350 ^ n98;
  assign new_n17352 = new_n17348 & new_n17351;
  assign new_n17353 = new_n17352 ^ new_n3452;
  assign new_n17354 = new_n17353 ^ new_n17347;
  assign new_n17355 = new_n17354 ^ new_n3452;
  assign new_n17356 = new_n17355 ^ new_n17343;
  assign new_n17357 = n102 & new_n9195;
  assign new_n17358 = new_n4368 & new_n9185;
  assign new_n17359 = new_n17358 ^ new_n17357;
  assign new_n17360 = n103 & new_n9184;
  assign new_n17361 = n101 & new_n9189;
  assign new_n17362 = new_n17361 ^ new_n17360;
  assign new_n17363 = new_n17362 ^ new_n17359;
  assign new_n17364 = new_n17363 ^ n63;
  assign new_n17365 = new_n17364 ^ new_n17356;
  assign new_n17366 = new_n17365 ^ new_n17340;
  assign new_n17367 = new_n17366 ^ new_n17332;
  assign new_n17368 = new_n17367 ^ new_n17320;
  assign new_n17369 = new_n17368 ^ new_n17308;
  assign new_n17370 = new_n17214 ^ new_n17157;
  assign new_n17371 = new_n17158 & new_n17370;
  assign new_n17372 = new_n17371 ^ new_n17154;
  assign new_n17373 = new_n17372 ^ new_n17369;
  assign new_n17374 = new_n17373 ^ new_n17296;
  assign new_n17375 = new_n17219 ^ new_n17146;
  assign new_n17376 = new_n17216 & new_n17375;
  assign new_n17377 = new_n17376 ^ new_n17219;
  assign new_n17378 = new_n17377 ^ new_n17374;
  assign new_n17379 = ~new_n4804 & n120;
  assign new_n17380 = new_n4799 & new_n8560;
  assign new_n17381 = new_n17380 ^ new_n17379;
  assign new_n17382 = n121 & new_n4798;
  assign new_n17383 = n119 & new_n4810;
  assign new_n17384 = new_n17383 ^ new_n17382;
  assign new_n17385 = new_n17384 ^ new_n17381;
  assign new_n17386 = new_n17385 ^ n45;
  assign new_n17387 = new_n17386 ^ new_n17378;
  assign new_n17388 = new_n17232 ^ new_n17220;
  assign new_n17389 = ~new_n17224 & new_n17388;
  assign new_n17390 = new_n17389 ^ new_n17223;
  assign new_n17391 = new_n17390 ^ new_n17387;
  assign new_n17392 = new_n17391 ^ new_n17288;
  assign new_n17393 = new_n17236 ^ new_n17138;
  assign new_n17394 = new_n17237 & new_n17393;
  assign new_n17395 = new_n17394 ^ new_n17138;
  assign new_n17396 = new_n17395 ^ new_n17392;
  assign new_n17397 = new_n17396 ^ new_n17280;
  assign new_n17398 = new_n17238 ^ new_n17130;
  assign new_n17399 = ~new_n17398 & new_n17242;
  assign new_n17400 = new_n17399 ^ new_n17130;
  assign new_n17401 = new_n17400 ^ new_n17397;
  assign new_n17402 = ~new_n3148 & n128;
  assign new_n17403 = ~n36 & ~new_n17402;
  assign new_n17404 = new_n17403 ^ n35;
  assign new_n17405 = new_n2825 & new_n11133;
  assign new_n17406 = new_n17405 ^ new_n17402;
  assign new_n17407 = ~new_n17404 & ~new_n17406;
  assign new_n17408 = new_n17407 ^ n35;
  assign new_n17409 = new_n17408 ^ new_n17401;
  assign new_n17410 = new_n17409 ^ new_n17272;
  assign new_n17411 = ~new_n17260 & ~new_n17409;
  assign new_n17412 = ~new_n17251 & ~new_n17411;
  assign new_n17413 = ~new_n17252 & ~new_n17409;
  assign new_n17414 = ~new_n17413 & new_n17261;
  assign new_n17415 = ~new_n17412 & ~new_n17414;
  assign new_n17416 = ~new_n17415 & new_n17267;
  assign new_n17417 = new_n17261 ^ new_n17243;
  assign new_n17418 = ~new_n17250 & ~new_n17417;
  assign new_n17419 = new_n17418 ^ new_n17249;
  assign new_n17420 = ~new_n17419 & new_n17409;
  assign new_n17421 = new_n17260 & new_n17414;
  assign new_n17422 = ~new_n17420 & ~new_n17421;
  assign new_n17423 = ~new_n17416 & new_n17422;
  assign new_n17424 = ~new_n3682 & n127;
  assign new_n17425 = new_n3677 & new_n10581;
  assign new_n17426 = new_n17425 ^ new_n17424;
  assign new_n17427 = n128 & new_n3676;
  assign new_n17428 = n126 & new_n3688;
  assign new_n17429 = new_n17428 ^ new_n17427;
  assign new_n17430 = new_n17429 ^ new_n17426;
  assign new_n17431 = new_n17430 ^ n39;
  assign new_n17432 = ~new_n4212 & n124;
  assign new_n17433 = new_n4201 & new_n9700;
  assign new_n17434 = new_n17433 ^ new_n17432;
  assign new_n17435 = n125 & new_n4200;
  assign new_n17436 = n123 & new_n4206;
  assign new_n17437 = new_n17436 ^ new_n17435;
  assign new_n17438 = new_n17437 ^ new_n17434;
  assign new_n17439 = new_n17438 ^ n42;
  assign new_n17440 = ~new_n4804 & n121;
  assign new_n17441 = new_n4799 & new_n8850;
  assign new_n17442 = new_n17441 ^ new_n17440;
  assign new_n17443 = n122 & new_n4798;
  assign new_n17444 = n120 & new_n4810;
  assign new_n17445 = new_n17444 ^ new_n17443;
  assign new_n17446 = new_n17445 ^ new_n17442;
  assign new_n17447 = new_n17446 ^ n45;
  assign new_n17448 = ~new_n6805 & n112;
  assign new_n17449 = ~new_n6518 & new_n6800;
  assign new_n17450 = new_n17449 ^ new_n17448;
  assign new_n17451 = n113 & new_n6799;
  assign new_n17452 = n111 & new_n6811;
  assign new_n17453 = new_n17452 ^ new_n17451;
  assign new_n17454 = new_n17453 ^ new_n17450;
  assign new_n17455 = new_n17454 ^ n54;
  assign new_n17456 = n109 & new_n7553;
  assign new_n17457 = new_n5825 & new_n7543;
  assign new_n17458 = new_n17457 ^ new_n17456;
  assign new_n17459 = n110 & new_n7542;
  assign new_n17460 = n108 & new_n7547;
  assign new_n17461 = new_n17460 ^ new_n17459;
  assign new_n17462 = new_n17461 ^ new_n17458;
  assign new_n17463 = new_n17462 ^ n57;
  assign new_n17464 = new_n17366 ^ new_n17328;
  assign new_n17465 = new_n17332 & new_n17464;
  assign new_n17466 = new_n17465 ^ new_n17331;
  assign new_n17467 = new_n17466 ^ new_n17463;
  assign new_n17468 = n106 & new_n8355;
  assign new_n17469 = ~new_n5164 & new_n8345;
  assign new_n17470 = new_n17469 ^ new_n17468;
  assign new_n17471 = n107 & new_n8344;
  assign new_n17472 = n105 & new_n8349;
  assign new_n17473 = new_n17472 ^ new_n17471;
  assign new_n17474 = new_n17473 ^ new_n17470;
  assign new_n17475 = new_n17474 ^ n60;
  assign new_n17476 = new_n17356 ^ new_n17340;
  assign new_n17477 = ~new_n17476 & new_n17365;
  assign new_n17478 = new_n17477 ^ new_n17340;
  assign new_n17479 = new_n17478 ^ new_n17475;
  assign new_n17480 = ~new_n17343 & ~new_n17347;
  assign new_n17481 = ~new_n17352 & ~new_n17480;
  assign new_n17482 = n103 & new_n9195;
  assign new_n17483 = ~new_n4556 & new_n9185;
  assign new_n17484 = new_n17483 ^ new_n17482;
  assign new_n17485 = n104 & new_n9184;
  assign new_n17486 = n102 & new_n9189;
  assign new_n17487 = new_n17486 ^ new_n17485;
  assign new_n17488 = new_n17487 ^ new_n17484;
  assign new_n17489 = new_n17488 ^ n63;
  assign new_n17490 = n101 ^ n99;
  assign new_n17491 = ~new_n11492 & new_n17490;
  assign new_n17492 = new_n17491 ^ n99;
  assign new_n17493 = new_n17492 ^ n100;
  assign new_n17494 = new_n11789 & new_n17493;
  assign new_n17495 = new_n17494 ^ n36;
  assign new_n17496 = new_n17495 ^ new_n17489;
  assign new_n17497 = new_n17496 ^ new_n17481;
  assign new_n17498 = new_n17497 ^ new_n17479;
  assign new_n17499 = new_n17498 ^ new_n17467;
  assign new_n17500 = new_n17499 ^ new_n17455;
  assign new_n17501 = new_n17367 ^ new_n17319;
  assign new_n17502 = new_n17320 & new_n17501;
  assign new_n17503 = new_n17502 ^ new_n17316;
  assign new_n17504 = new_n17503 ^ new_n17500;
  assign new_n17505 = new_n17368 ^ new_n17307;
  assign new_n17506 = new_n17308 & new_n17505;
  assign new_n17507 = new_n17506 ^ new_n17304;
  assign new_n17508 = new_n17507 ^ new_n17504;
  assign new_n17509 = ~new_n6110 & n115;
  assign new_n17510 = ~new_n7256 & new_n6105;
  assign new_n17511 = new_n17510 ^ new_n17509;
  assign new_n17512 = n116 & new_n6104;
  assign new_n17513 = n114 & new_n6347;
  assign new_n17514 = new_n17513 ^ new_n17512;
  assign new_n17515 = new_n17514 ^ new_n17511;
  assign new_n17516 = new_n17515 ^ n51;
  assign new_n17517 = new_n17516 ^ new_n17508;
  assign new_n17518 = ~new_n5424 & n118;
  assign new_n17519 = ~new_n8019 & new_n5419;
  assign new_n17520 = new_n17519 ^ new_n17518;
  assign new_n17521 = n119 & new_n5418;
  assign new_n17522 = n117 & new_n5648;
  assign new_n17523 = new_n17522 ^ new_n17521;
  assign new_n17524 = new_n17523 ^ new_n17520;
  assign new_n17525 = new_n17524 ^ n48;
  assign new_n17526 = new_n17525 ^ new_n17517;
  assign new_n17527 = new_n17369 ^ new_n17296;
  assign new_n17528 = ~new_n17527 & new_n17373;
  assign new_n17529 = new_n17528 ^ new_n17296;
  assign new_n17530 = new_n17529 ^ new_n17526;
  assign new_n17531 = new_n17530 ^ new_n17447;
  assign new_n17532 = new_n17386 ^ new_n17374;
  assign new_n17533 = ~new_n17378 & new_n17532;
  assign new_n17534 = new_n17533 ^ new_n17377;
  assign new_n17535 = new_n17534 ^ new_n17531;
  assign new_n17536 = new_n17535 ^ new_n17439;
  assign new_n17537 = new_n17390 ^ new_n17288;
  assign new_n17538 = new_n17391 & new_n17537;
  assign new_n17539 = new_n17538 ^ new_n17288;
  assign new_n17540 = new_n17539 ^ new_n17536;
  assign new_n17541 = new_n17540 ^ new_n17431;
  assign new_n17542 = new_n17392 ^ new_n17280;
  assign new_n17543 = ~new_n17542 & new_n17396;
  assign new_n17544 = new_n17543 ^ new_n17280;
  assign new_n17545 = new_n17544 ^ new_n17541;
  assign new_n17546 = new_n17408 ^ new_n17397;
  assign new_n17547 = ~new_n17546 & new_n17401;
  assign new_n17548 = new_n17547 ^ new_n17408;
  assign new_n17549 = new_n17548 ^ new_n17545;
  assign new_n17550 = new_n17549 ^ new_n17423;
  assign new_n17551 = ~new_n4212 & n125;
  assign new_n17552 = new_n4201 & new_n9987;
  assign new_n17553 = new_n17552 ^ new_n17551;
  assign new_n17554 = n126 & new_n4200;
  assign new_n17555 = n124 & new_n4206;
  assign new_n17556 = new_n17555 ^ new_n17554;
  assign new_n17557 = new_n17556 ^ new_n17553;
  assign new_n17558 = new_n17557 ^ n42;
  assign new_n17559 = ~new_n4804 & n122;
  assign new_n17560 = ~new_n9116 & new_n4799;
  assign new_n17561 = new_n17560 ^ new_n17559;
  assign new_n17562 = n123 & new_n4798;
  assign new_n17563 = n121 & new_n4810;
  assign new_n17564 = new_n17563 ^ new_n17562;
  assign new_n17565 = new_n17564 ^ new_n17561;
  assign new_n17566 = new_n17565 ^ n45;
  assign new_n17567 = ~new_n6110 & n116;
  assign new_n17568 = ~new_n7503 & new_n6105;
  assign new_n17569 = new_n17568 ^ new_n17567;
  assign new_n17570 = n117 & new_n6104;
  assign new_n17571 = n115 & new_n6347;
  assign new_n17572 = new_n17571 ^ new_n17570;
  assign new_n17573 = new_n17572 ^ new_n17569;
  assign new_n17574 = new_n17573 ^ n51;
  assign new_n17575 = new_n17503 ^ new_n17455;
  assign new_n17576 = new_n17500 & new_n17575;
  assign new_n17577 = new_n17576 ^ new_n17503;
  assign new_n17578 = new_n17577 ^ new_n17574;
  assign new_n17579 = ~new_n6805 & n113;
  assign new_n17580 = ~new_n6764 & new_n6800;
  assign new_n17581 = new_n17580 ^ new_n17579;
  assign new_n17582 = n114 & new_n6799;
  assign new_n17583 = n112 & new_n6811;
  assign new_n17584 = new_n17583 ^ new_n17582;
  assign new_n17585 = new_n17584 ^ new_n17581;
  assign new_n17586 = new_n17585 ^ n54;
  assign new_n17587 = new_n17498 ^ new_n17463;
  assign new_n17588 = new_n17467 & new_n17587;
  assign new_n17589 = new_n17588 ^ new_n17466;
  assign new_n17590 = new_n17589 ^ new_n17586;
  assign new_n17591 = n110 & new_n7553;
  assign new_n17592 = new_n6049 & new_n7543;
  assign new_n17593 = new_n17592 ^ new_n17591;
  assign new_n17594 = n111 & new_n7542;
  assign new_n17595 = n109 & new_n7547;
  assign new_n17596 = new_n17595 ^ new_n17594;
  assign new_n17597 = new_n17596 ^ new_n17593;
  assign new_n17598 = new_n17597 ^ n57;
  assign new_n17599 = new_n17497 ^ new_n17475;
  assign new_n17600 = new_n17479 & new_n17599;
  assign new_n17601 = new_n17600 ^ new_n17478;
  assign new_n17602 = new_n17601 ^ new_n17598;
  assign new_n17603 = n107 & new_n8355;
  assign new_n17604 = ~new_n5377 & new_n8345;
  assign new_n17605 = new_n17604 ^ new_n17603;
  assign new_n17606 = n108 & new_n8344;
  assign new_n17607 = n106 & new_n8349;
  assign new_n17608 = new_n17607 ^ new_n17606;
  assign new_n17609 = new_n17608 ^ new_n17605;
  assign new_n17610 = new_n17609 ^ n60;
  assign new_n17611 = new_n17489 ^ new_n17481;
  assign new_n17612 = new_n17496 & new_n17611;
  assign new_n17613 = new_n17612 ^ new_n17481;
  assign new_n17614 = new_n17613 ^ new_n17610;
  assign new_n17615 = n104 & new_n9195;
  assign new_n17616 = ~new_n4754 & new_n9185;
  assign new_n17617 = new_n17616 ^ new_n17615;
  assign new_n17618 = n105 & new_n9184;
  assign new_n17619 = n103 & new_n9189;
  assign new_n17620 = new_n17619 ^ new_n17618;
  assign new_n17621 = new_n17620 ^ new_n17617;
  assign new_n17622 = new_n17621 ^ n63;
  assign new_n17623 = n101 & new_n11492;
  assign new_n17624 = n102 & new_n9495;
  assign new_n17625 = new_n17624 ^ new_n17623;
  assign new_n17626 = n100 ^ n36;
  assign new_n17627 = ~new_n17626 & new_n17493;
  assign new_n17628 = new_n17627 ^ n100;
  assign new_n17629 = new_n11789 & new_n17628;
  assign new_n17630 = new_n17629 ^ new_n17625;
  assign new_n17631 = new_n17630 ^ new_n17622;
  assign new_n17632 = new_n17631 ^ new_n17614;
  assign new_n17633 = new_n17632 ^ new_n17602;
  assign new_n17634 = new_n17633 ^ new_n17590;
  assign new_n17635 = new_n17634 ^ new_n17578;
  assign new_n17636 = new_n17516 ^ new_n17504;
  assign new_n17637 = ~new_n17508 & new_n17636;
  assign new_n17638 = new_n17637 ^ new_n17507;
  assign new_n17639 = new_n17638 ^ new_n17635;
  assign new_n17640 = ~new_n5424 & n119;
  assign new_n17641 = new_n5419 & new_n8286;
  assign new_n17642 = new_n17641 ^ new_n17640;
  assign new_n17643 = n120 & new_n5418;
  assign new_n17644 = n118 & new_n5648;
  assign new_n17645 = new_n17644 ^ new_n17643;
  assign new_n17646 = new_n17645 ^ new_n17642;
  assign new_n17647 = new_n17646 ^ n48;
  assign new_n17648 = new_n17647 ^ new_n17639;
  assign new_n17649 = new_n17529 ^ new_n17525;
  assign new_n17650 = ~new_n17526 & ~new_n17649;
  assign new_n17651 = new_n17650 ^ new_n17517;
  assign new_n17652 = new_n17651 ^ new_n17648;
  assign new_n17653 = new_n17652 ^ new_n17566;
  assign new_n17654 = new_n17534 ^ new_n17447;
  assign new_n17655 = new_n17531 & new_n17654;
  assign new_n17656 = new_n17655 ^ new_n17534;
  assign new_n17657 = new_n17656 ^ new_n17653;
  assign new_n17658 = new_n17657 ^ new_n17558;
  assign new_n17659 = new_n17539 ^ new_n17439;
  assign new_n17660 = new_n17536 & new_n17659;
  assign new_n17661 = new_n17660 ^ new_n17539;
  assign new_n17662 = new_n17661 ^ new_n17658;
  assign new_n17663 = n127 & new_n3688;
  assign new_n17664 = new_n3677 & new_n10010;
  assign new_n17665 = new_n17664 ^ new_n17663;
  assign new_n17666 = ~new_n3682 & n128;
  assign new_n17667 = new_n17666 ^ new_n17665;
  assign new_n17668 = new_n17667 ^ n39;
  assign new_n17669 = new_n17668 ^ new_n17662;
  assign new_n17670 = new_n17544 ^ new_n17431;
  assign new_n17671 = new_n17541 & new_n17670;
  assign new_n17672 = new_n17671 ^ new_n17544;
  assign new_n17673 = new_n17672 ^ new_n17669;
  assign new_n17674 = new_n17548 ^ new_n17423;
  assign new_n17675 = new_n17549 & new_n17674;
  assign new_n17676 = new_n17675 ^ new_n17423;
  assign new_n17677 = new_n17676 ^ new_n17673;
  assign new_n17678 = ~new_n4212 & n126;
  assign new_n17679 = new_n4201 & new_n10304;
  assign new_n17680 = new_n17679 ^ new_n17678;
  assign new_n17681 = n127 & new_n4200;
  assign new_n17682 = n125 & new_n4206;
  assign new_n17683 = new_n17682 ^ new_n17681;
  assign new_n17684 = new_n17683 ^ new_n17680;
  assign new_n17685 = new_n17684 ^ n42;
  assign new_n17686 = ~new_n4804 & n123;
  assign new_n17687 = ~new_n9405 & new_n4799;
  assign new_n17688 = new_n17687 ^ new_n17686;
  assign new_n17689 = n124 & new_n4798;
  assign new_n17690 = n122 & new_n4810;
  assign new_n17691 = new_n17690 ^ new_n17689;
  assign new_n17692 = new_n17691 ^ new_n17688;
  assign new_n17693 = new_n17692 ^ n45;
  assign new_n17694 = ~new_n6110 & n117;
  assign new_n17695 = ~new_n7761 & new_n6105;
  assign new_n17696 = new_n17695 ^ new_n17694;
  assign new_n17697 = n118 & new_n6104;
  assign new_n17698 = n116 & new_n6347;
  assign new_n17699 = new_n17698 ^ new_n17697;
  assign new_n17700 = new_n17699 ^ new_n17696;
  assign new_n17701 = new_n17700 ^ n51;
  assign new_n17702 = ~new_n6805 & n114;
  assign new_n17703 = ~new_n7013 & new_n6800;
  assign new_n17704 = new_n17703 ^ new_n17702;
  assign new_n17705 = n115 & new_n6799;
  assign new_n17706 = n113 & new_n6811;
  assign new_n17707 = new_n17706 ^ new_n17705;
  assign new_n17708 = new_n17707 ^ new_n17704;
  assign new_n17709 = new_n17708 ^ n54;
  assign new_n17710 = n111 & new_n7553;
  assign new_n17711 = ~new_n6284 & new_n7543;
  assign new_n17712 = new_n17711 ^ new_n17710;
  assign new_n17713 = n112 & new_n7542;
  assign new_n17714 = n110 & new_n7547;
  assign new_n17715 = new_n17714 ^ new_n17713;
  assign new_n17716 = new_n17715 ^ new_n17712;
  assign new_n17717 = new_n17716 ^ n57;
  assign new_n17718 = new_n17631 ^ new_n17610;
  assign new_n17719 = new_n17614 & new_n17718;
  assign new_n17720 = new_n17719 ^ new_n17613;
  assign new_n17721 = new_n17720 ^ new_n17717;
  assign new_n17722 = n108 & new_n8355;
  assign new_n17723 = new_n5604 & new_n8345;
  assign new_n17724 = new_n17723 ^ new_n17722;
  assign new_n17725 = n109 & new_n8344;
  assign new_n17726 = n107 & new_n8349;
  assign new_n17727 = new_n17726 ^ new_n17725;
  assign new_n17728 = new_n17727 ^ new_n17724;
  assign new_n17729 = new_n17728 ^ n60;
  assign new_n17730 = new_n17629 ^ new_n17622;
  assign new_n17731 = new_n17630 & new_n17730;
  assign new_n17732 = new_n17731 ^ new_n17622;
  assign new_n17733 = n103 ^ n102;
  assign new_n17734 = n102 ^ n101;
  assign new_n17735 = new_n17734 ^ new_n17733;
  assign new_n17736 = new_n17735 ^ new_n17734;
  assign new_n17737 = new_n17736 ^ new_n17735;
  assign new_n17738 = new_n17735 ^ n63;
  assign new_n17739 = new_n17738 ^ new_n17735;
  assign new_n17740 = ~new_n17739 & new_n17737;
  assign new_n17741 = new_n17740 ^ new_n17735;
  assign new_n17742 = ~new_n9495 & new_n17741;
  assign new_n17743 = new_n17742 ^ new_n17733;
  assign new_n17744 = new_n17743 ^ new_n17732;
  assign new_n17745 = new_n17744 ^ new_n17729;
  assign new_n17746 = n105 & new_n9195;
  assign new_n17747 = ~new_n4961 & new_n9185;
  assign new_n17748 = new_n17747 ^ new_n17746;
  assign new_n17749 = n106 & new_n9184;
  assign new_n17750 = n104 & new_n9189;
  assign new_n17751 = new_n17750 ^ new_n17749;
  assign new_n17752 = new_n17751 ^ new_n17748;
  assign new_n17753 = new_n17752 ^ n63;
  assign new_n17754 = new_n17753 ^ new_n17745;
  assign new_n17755 = new_n17754 ^ new_n17721;
  assign new_n17756 = new_n17632 ^ new_n17598;
  assign new_n17757 = new_n17602 & new_n17756;
  assign new_n17758 = new_n17757 ^ new_n17601;
  assign new_n17759 = new_n17758 ^ new_n17755;
  assign new_n17760 = new_n17759 ^ new_n17709;
  assign new_n17761 = new_n17760 ^ new_n17701;
  assign new_n17762 = new_n17633 ^ new_n17589;
  assign new_n17763 = new_n17590 & new_n17762;
  assign new_n17764 = new_n17763 ^ new_n17586;
  assign new_n17765 = new_n17764 ^ new_n17761;
  assign new_n17766 = new_n17634 ^ new_n17577;
  assign new_n17767 = new_n17578 & new_n17766;
  assign new_n17768 = new_n17767 ^ new_n17574;
  assign new_n17769 = new_n17768 ^ new_n17765;
  assign new_n17770 = ~new_n5424 & n120;
  assign new_n17771 = new_n5419 & new_n8560;
  assign new_n17772 = new_n17771 ^ new_n17770;
  assign new_n17773 = n121 & new_n5418;
  assign new_n17774 = n119 & new_n5648;
  assign new_n17775 = new_n17774 ^ new_n17773;
  assign new_n17776 = new_n17775 ^ new_n17772;
  assign new_n17777 = new_n17776 ^ n48;
  assign new_n17778 = new_n17777 ^ new_n17769;
  assign new_n17779 = new_n17647 ^ new_n17635;
  assign new_n17780 = ~new_n17639 & new_n17779;
  assign new_n17781 = new_n17780 ^ new_n17638;
  assign new_n17782 = new_n17781 ^ new_n17778;
  assign new_n17783 = new_n17782 ^ new_n17693;
  assign new_n17784 = new_n17651 ^ new_n17566;
  assign new_n17785 = ~new_n17652 & ~new_n17784;
  assign new_n17786 = new_n17785 ^ new_n17566;
  assign new_n17787 = new_n17786 ^ new_n17783;
  assign new_n17788 = new_n17787 ^ new_n17685;
  assign new_n17789 = new_n17656 ^ new_n17558;
  assign new_n17790 = ~new_n17657 & new_n17789;
  assign new_n17791 = new_n17790 ^ new_n17558;
  assign new_n17792 = new_n17791 ^ new_n17788;
  assign new_n17793 = ~new_n3687 & n128;
  assign new_n17794 = ~n39 & ~new_n17793;
  assign new_n17795 = new_n17794 ^ n38;
  assign new_n17796 = new_n3313 & new_n11133;
  assign new_n17797 = new_n17796 ^ new_n17793;
  assign new_n17798 = ~new_n17795 & ~new_n17797;
  assign new_n17799 = new_n17798 ^ n38;
  assign new_n17800 = new_n17799 ^ new_n17792;
  assign new_n17801 = new_n17668 ^ new_n17658;
  assign new_n17802 = ~new_n17801 & new_n17662;
  assign new_n17803 = new_n17802 ^ new_n17661;
  assign new_n17804 = new_n17803 ^ new_n17800;
  assign new_n17805 = new_n17676 ^ new_n17672;
  assign new_n17806 = ~new_n17673 & new_n17805;
  assign new_n17807 = new_n17806 ^ new_n17676;
  assign new_n17808 = new_n17807 ^ new_n17804;
  assign new_n17809 = new_n17807 ^ new_n17803;
  assign new_n17810 = new_n17804 & new_n17809;
  assign new_n17811 = new_n17810 ^ new_n17807;
  assign new_n17812 = ~new_n6110 & n118;
  assign new_n17813 = ~new_n8019 & new_n6105;
  assign new_n17814 = new_n17813 ^ new_n17812;
  assign new_n17815 = n119 & new_n6104;
  assign new_n17816 = n117 & new_n6347;
  assign new_n17817 = new_n17816 ^ new_n17815;
  assign new_n17818 = new_n17817 ^ new_n17814;
  assign new_n17819 = new_n17818 ^ n51;
  assign new_n17820 = new_n17764 ^ new_n17760;
  assign new_n17821 = ~new_n17761 & new_n17820;
  assign new_n17822 = new_n17821 ^ new_n17701;
  assign new_n17823 = new_n17822 ^ new_n17819;
  assign new_n17824 = ~new_n6805 & n115;
  assign new_n17825 = ~new_n7256 & new_n6800;
  assign new_n17826 = new_n17825 ^ new_n17824;
  assign new_n17827 = n116 & new_n6799;
  assign new_n17828 = n114 & new_n6811;
  assign new_n17829 = new_n17828 ^ new_n17827;
  assign new_n17830 = new_n17829 ^ new_n17826;
  assign new_n17831 = new_n17830 ^ n54;
  assign new_n17832 = new_n17758 ^ new_n17709;
  assign new_n17833 = new_n17759 & new_n17832;
  assign new_n17834 = new_n17833 ^ new_n17709;
  assign new_n17835 = new_n17834 ^ new_n17831;
  assign new_n17836 = n112 & new_n7553;
  assign new_n17837 = ~new_n6518 & new_n7543;
  assign new_n17838 = new_n17837 ^ new_n17836;
  assign new_n17839 = n113 & new_n7542;
  assign new_n17840 = n111 & new_n7547;
  assign new_n17841 = new_n17840 ^ new_n17839;
  assign new_n17842 = new_n17841 ^ new_n17838;
  assign new_n17843 = new_n17842 ^ n57;
  assign new_n17844 = new_n17754 ^ new_n17720;
  assign new_n17845 = new_n17721 & new_n17844;
  assign new_n17846 = new_n17845 ^ new_n17717;
  assign new_n17847 = new_n17846 ^ new_n17843;
  assign new_n17848 = n109 & new_n8355;
  assign new_n17849 = new_n5825 & new_n8345;
  assign new_n17850 = new_n17849 ^ new_n17848;
  assign new_n17851 = n110 & new_n8344;
  assign new_n17852 = n108 & new_n8349;
  assign new_n17853 = new_n17852 ^ new_n17851;
  assign new_n17854 = new_n17853 ^ new_n17850;
  assign new_n17855 = new_n17854 ^ n60;
  assign new_n17856 = new_n17753 ^ new_n17744;
  assign new_n17857 = ~new_n17745 & new_n17856;
  assign new_n17858 = new_n17857 ^ new_n17729;
  assign new_n17859 = new_n17858 ^ new_n17855;
  assign new_n17860 = n106 & new_n9195;
  assign new_n17861 = ~new_n5164 & new_n9185;
  assign new_n17862 = new_n17861 ^ new_n17860;
  assign new_n17863 = n107 & new_n9184;
  assign new_n17864 = n105 & new_n9189;
  assign new_n17865 = new_n17864 ^ new_n17863;
  assign new_n17866 = new_n17865 ^ new_n17862;
  assign new_n17867 = new_n17866 ^ n63;
  assign new_n17868 = n64 & n103;
  assign new_n17869 = new_n17868 ^ n104;
  assign new_n17870 = ~new_n9495 & new_n17869;
  assign new_n17871 = new_n17870 ^ n104;
  assign new_n17872 = new_n17871 ^ new_n17625;
  assign new_n17873 = new_n17872 ^ n39;
  assign new_n17874 = new_n17873 ^ new_n17867;
  assign new_n17875 = ~n103 & new_n9495;
  assign new_n17876 = new_n17875 ^ new_n17623;
  assign new_n17877 = n102 & new_n17876;
  assign new_n17878 = new_n17877 ^ new_n17623;
  assign new_n17879 = ~new_n17732 & ~new_n17743;
  assign new_n17880 = new_n17879 ^ new_n17878;
  assign new_n17881 = new_n17880 ^ new_n17874;
  assign new_n17882 = new_n17881 ^ new_n17859;
  assign new_n17883 = new_n17882 ^ new_n17847;
  assign new_n17884 = new_n17883 ^ new_n17835;
  assign new_n17885 = new_n17884 ^ new_n17823;
  assign new_n17886 = ~new_n5424 & n121;
  assign new_n17887 = new_n5419 & new_n8850;
  assign new_n17888 = new_n17887 ^ new_n17886;
  assign new_n17889 = n122 & new_n5418;
  assign new_n17890 = n120 & new_n5648;
  assign new_n17891 = new_n17890 ^ new_n17889;
  assign new_n17892 = new_n17891 ^ new_n17888;
  assign new_n17893 = new_n17892 ^ n48;
  assign new_n17894 = new_n17893 ^ new_n17885;
  assign new_n17895 = new_n17777 ^ new_n17768;
  assign new_n17896 = ~new_n17769 & ~new_n17895;
  assign new_n17897 = new_n17896 ^ new_n17765;
  assign new_n17898 = new_n17897 ^ new_n17894;
  assign new_n17899 = new_n17781 ^ new_n17693;
  assign new_n17900 = new_n17782 & new_n17899;
  assign new_n17901 = new_n17900 ^ new_n17693;
  assign new_n17902 = new_n17901 ^ new_n17898;
  assign new_n17903 = ~new_n4804 & n124;
  assign new_n17904 = new_n4799 & new_n9700;
  assign new_n17905 = new_n17904 ^ new_n17903;
  assign new_n17906 = n125 & new_n4798;
  assign new_n17907 = n123 & new_n4810;
  assign new_n17908 = new_n17907 ^ new_n17906;
  assign new_n17909 = new_n17908 ^ new_n17905;
  assign new_n17910 = new_n17909 ^ n45;
  assign new_n17911 = new_n17910 ^ new_n17902;
  assign new_n17912 = new_n17799 ^ new_n17788;
  assign new_n17913 = ~new_n17912 & new_n17792;
  assign new_n17914 = new_n17913 ^ new_n17799;
  assign new_n17915 = new_n17914 ^ new_n17911;
  assign new_n17916 = ~new_n4212 & n127;
  assign new_n17917 = new_n4201 & new_n10581;
  assign new_n17918 = new_n17917 ^ new_n17916;
  assign new_n17919 = n128 & new_n4200;
  assign new_n17920 = n126 & new_n4206;
  assign new_n17921 = new_n17920 ^ new_n17919;
  assign new_n17922 = new_n17921 ^ new_n17918;
  assign new_n17923 = new_n17922 ^ n42;
  assign new_n17924 = new_n17786 ^ new_n17685;
  assign new_n17925 = new_n17787 & new_n17924;
  assign new_n17926 = new_n17925 ^ new_n17685;
  assign new_n17927 = new_n17926 ^ new_n17923;
  assign new_n17928 = new_n17927 ^ new_n17915;
  assign new_n17929 = new_n17928 ^ new_n17811;
  assign new_n17930 = new_n17923 & new_n17926;
  assign new_n17931 = new_n17930 ^ new_n17927;
  assign new_n17932 = ~new_n17931 & new_n17811;
  assign new_n17933 = new_n17931 ^ new_n17911;
  assign new_n17934 = ~new_n17915 & new_n17933;
  assign new_n17935 = new_n17934 ^ new_n17914;
  assign new_n17936 = ~new_n17914 & new_n17911;
  assign new_n17937 = new_n17936 ^ new_n17935;
  assign new_n17938 = new_n17937 ^ new_n17932;
  assign new_n17939 = new_n17930 ^ new_n17915;
  assign new_n17940 = new_n17930 ^ new_n17811;
  assign new_n17941 = ~new_n17940 & new_n17939;
  assign new_n17942 = new_n17941 ^ new_n17938;
  assign new_n17943 = new_n17936 ^ new_n17915;
  assign new_n17944 = new_n17943 ^ new_n17942;
  assign new_n17945 = ~new_n4804 & n125;
  assign new_n17946 = new_n4799 & new_n9987;
  assign new_n17947 = new_n17946 ^ new_n17945;
  assign new_n17948 = n126 & new_n4798;
  assign new_n17949 = n124 & new_n4810;
  assign new_n17950 = new_n17949 ^ new_n17948;
  assign new_n17951 = new_n17950 ^ new_n17947;
  assign new_n17952 = new_n17951 ^ n45;
  assign new_n17953 = ~new_n5424 & n122;
  assign new_n17954 = ~new_n9116 & new_n5419;
  assign new_n17955 = new_n17954 ^ new_n17953;
  assign new_n17956 = n123 & new_n5418;
  assign new_n17957 = n121 & new_n5648;
  assign new_n17958 = new_n17957 ^ new_n17956;
  assign new_n17959 = new_n17958 ^ new_n17955;
  assign new_n17960 = new_n17959 ^ n48;
  assign new_n17961 = ~new_n6110 & n119;
  assign new_n17962 = new_n6105 & new_n8286;
  assign new_n17963 = new_n17962 ^ new_n17961;
  assign new_n17964 = n120 & new_n6104;
  assign new_n17965 = n118 & new_n6347;
  assign new_n17966 = new_n17965 ^ new_n17964;
  assign new_n17967 = new_n17966 ^ new_n17963;
  assign new_n17968 = new_n17967 ^ n51;
  assign new_n17969 = ~new_n6805 & n116;
  assign new_n17970 = ~new_n7503 & new_n6800;
  assign new_n17971 = new_n17970 ^ new_n17969;
  assign new_n17972 = n117 & new_n6799;
  assign new_n17973 = n115 & new_n6811;
  assign new_n17974 = new_n17973 ^ new_n17972;
  assign new_n17975 = new_n17974 ^ new_n17971;
  assign new_n17976 = new_n17975 ^ n54;
  assign new_n17977 = new_n17882 ^ new_n17843;
  assign new_n17978 = ~new_n17977 & new_n17847;
  assign new_n17979 = new_n17978 ^ new_n17846;
  assign new_n17980 = new_n17979 ^ new_n17976;
  assign new_n17981 = n113 & new_n7553;
  assign new_n17982 = ~new_n6764 & new_n7543;
  assign new_n17983 = new_n17982 ^ new_n17981;
  assign new_n17984 = n114 & new_n7542;
  assign new_n17985 = n112 & new_n7547;
  assign new_n17986 = new_n17985 ^ new_n17984;
  assign new_n17987 = new_n17986 ^ new_n17983;
  assign new_n17988 = new_n17987 ^ n57;
  assign new_n17989 = new_n17881 ^ new_n17855;
  assign new_n17990 = ~new_n17989 & new_n17859;
  assign new_n17991 = new_n17990 ^ new_n17858;
  assign new_n17992 = new_n17991 ^ new_n17988;
  assign new_n17993 = n110 & new_n8355;
  assign new_n17994 = new_n6049 & new_n8345;
  assign new_n17995 = new_n17994 ^ new_n17993;
  assign new_n17996 = n111 & new_n8344;
  assign new_n17997 = n109 & new_n8349;
  assign new_n17998 = new_n17997 ^ new_n17996;
  assign new_n17999 = new_n17998 ^ new_n17995;
  assign new_n18000 = new_n17999 ^ n60;
  assign new_n18001 = n107 & new_n9195;
  assign new_n18002 = ~new_n5377 & new_n9185;
  assign new_n18003 = new_n18002 ^ new_n18001;
  assign new_n18004 = n108 & new_n9184;
  assign new_n18005 = n106 & new_n9189;
  assign new_n18006 = new_n18005 ^ new_n18004;
  assign new_n18007 = new_n18006 ^ new_n18003;
  assign new_n18008 = new_n18007 ^ n63;
  assign new_n18009 = new_n17625 ^ n39;
  assign new_n18010 = ~new_n17872 & ~new_n18009;
  assign new_n18011 = new_n18010 ^ n39;
  assign new_n18012 = n64 & n104;
  assign new_n18013 = new_n18012 ^ n105;
  assign new_n18014 = ~new_n9495 & new_n18013;
  assign new_n18015 = new_n18014 ^ n105;
  assign new_n18016 = new_n18015 ^ new_n18011;
  assign new_n18017 = new_n18016 ^ new_n18008;
  assign new_n18018 = new_n18017 ^ new_n18000;
  assign new_n18019 = new_n17880 ^ new_n17867;
  assign new_n18020 = ~new_n18019 & new_n17874;
  assign new_n18021 = new_n18020 ^ new_n17880;
  assign new_n18022 = new_n18021 ^ new_n18018;
  assign new_n18023 = new_n18022 ^ new_n17992;
  assign new_n18024 = new_n18023 ^ new_n17980;
  assign new_n18025 = new_n18024 ^ new_n17968;
  assign new_n18026 = new_n17883 ^ new_n17831;
  assign new_n18027 = ~new_n18026 & new_n17835;
  assign new_n18028 = new_n18027 ^ new_n17834;
  assign new_n18029 = new_n18028 ^ new_n18025;
  assign new_n18030 = new_n18029 ^ new_n17960;
  assign new_n18031 = new_n17884 ^ new_n17819;
  assign new_n18032 = ~new_n18031 & new_n17823;
  assign new_n18033 = new_n18032 ^ new_n17822;
  assign new_n18034 = new_n18033 ^ new_n18030;
  assign new_n18035 = new_n18034 ^ new_n17952;
  assign new_n18036 = new_n17897 ^ new_n17893;
  assign new_n18037 = new_n17894 & new_n18036;
  assign new_n18038 = new_n18037 ^ new_n17885;
  assign new_n18039 = new_n18038 ^ new_n18035;
  assign new_n18040 = new_n17910 ^ new_n17898;
  assign new_n18041 = ~new_n17902 & new_n18040;
  assign new_n18042 = new_n18041 ^ new_n17901;
  assign new_n18043 = new_n18042 ^ new_n18039;
  assign new_n18044 = n127 & new_n4206;
  assign new_n18045 = new_n4201 & new_n10010;
  assign new_n18046 = new_n18045 ^ new_n18044;
  assign new_n18047 = ~new_n4212 & n128;
  assign new_n18048 = new_n18047 ^ new_n18046;
  assign new_n18049 = new_n18048 ^ n42;
  assign new_n18050 = new_n18049 ^ new_n18043;
  assign new_n18051 = new_n18050 ^ new_n17944;
  assign new_n18052 = ~new_n17943 & new_n18050;
  assign new_n18053 = new_n17923 ^ new_n17811;
  assign new_n18054 = ~new_n18053 & new_n17927;
  assign new_n18055 = new_n18054 ^ new_n17926;
  assign new_n18056 = ~new_n18052 & new_n18055;
  assign new_n18057 = ~new_n17930 & new_n18050;
  assign new_n18058 = ~new_n17936 & ~new_n18057;
  assign new_n18059 = new_n17811 & new_n18058;
  assign new_n18060 = ~new_n18050 & new_n17935;
  assign new_n18061 = ~new_n18059 & ~new_n18060;
  assign new_n18062 = ~new_n18056 & new_n18061;
  assign new_n18063 = n128 & new_n4206;
  assign new_n18064 = new_n4201 & new_n11133;
  assign new_n18065 = new_n18064 ^ new_n18063;
  assign new_n18066 = new_n18065 ^ n42;
  assign new_n18067 = new_n18038 ^ new_n18034;
  assign new_n18068 = ~new_n18035 & new_n18067;
  assign new_n18069 = new_n18068 ^ new_n17952;
  assign new_n18070 = new_n18069 ^ new_n18066;
  assign new_n18071 = ~new_n4804 & n126;
  assign new_n18072 = new_n4799 & new_n10304;
  assign new_n18073 = new_n18072 ^ new_n18071;
  assign new_n18074 = n127 & new_n4798;
  assign new_n18075 = n125 & new_n4810;
  assign new_n18076 = new_n18075 ^ new_n18074;
  assign new_n18077 = new_n18076 ^ new_n18073;
  assign new_n18078 = new_n18077 ^ n45;
  assign new_n18079 = ~new_n6110 & n120;
  assign new_n18080 = new_n6105 & new_n8560;
  assign new_n18081 = new_n18080 ^ new_n18079;
  assign new_n18082 = n121 & new_n6104;
  assign new_n18083 = n119 & new_n6347;
  assign new_n18084 = new_n18083 ^ new_n18082;
  assign new_n18085 = new_n18084 ^ new_n18081;
  assign new_n18086 = new_n18085 ^ n51;
  assign new_n18087 = new_n18023 ^ new_n17976;
  assign new_n18088 = new_n17980 & new_n18087;
  assign new_n18089 = new_n18088 ^ new_n17979;
  assign new_n18090 = new_n18089 ^ new_n18086;
  assign new_n18091 = ~new_n6805 & n117;
  assign new_n18092 = ~new_n7761 & new_n6800;
  assign new_n18093 = new_n18092 ^ new_n18091;
  assign new_n18094 = n118 & new_n6799;
  assign new_n18095 = n116 & new_n6811;
  assign new_n18096 = new_n18095 ^ new_n18094;
  assign new_n18097 = new_n18096 ^ new_n18093;
  assign new_n18098 = new_n18097 ^ n54;
  assign new_n18099 = new_n18022 ^ new_n17991;
  assign new_n18100 = new_n17992 & new_n18099;
  assign new_n18101 = new_n18100 ^ new_n17988;
  assign new_n18102 = new_n18101 ^ new_n18098;
  assign new_n18103 = n114 & new_n7553;
  assign new_n18104 = ~new_n7013 & new_n7543;
  assign new_n18105 = new_n18104 ^ new_n18103;
  assign new_n18106 = n115 & new_n7542;
  assign new_n18107 = n113 & new_n7547;
  assign new_n18108 = new_n18107 ^ new_n18106;
  assign new_n18109 = new_n18108 ^ new_n18105;
  assign new_n18110 = new_n18109 ^ n57;
  assign new_n18111 = new_n18021 ^ new_n18000;
  assign new_n18112 = ~new_n18018 & ~new_n18111;
  assign new_n18113 = new_n18112 ^ new_n18021;
  assign new_n18114 = new_n18113 ^ new_n18110;
  assign new_n18115 = n111 & new_n8355;
  assign new_n18116 = ~new_n6284 & new_n8345;
  assign new_n18117 = new_n18116 ^ new_n18115;
  assign new_n18118 = n112 & new_n8344;
  assign new_n18119 = n110 & new_n8349;
  assign new_n18120 = new_n18119 ^ new_n18118;
  assign new_n18121 = new_n18120 ^ new_n18117;
  assign new_n18122 = new_n18121 ^ n60;
  assign new_n18123 = n64 & n105;
  assign new_n18124 = new_n18123 ^ n106;
  assign new_n18125 = ~new_n9495 & new_n18124;
  assign new_n18126 = new_n18125 ^ n106;
  assign new_n18127 = new_n18011 ^ new_n18008;
  assign new_n18128 = new_n18016 & new_n18127;
  assign new_n18129 = new_n18128 ^ new_n18126;
  assign new_n18130 = n108 & new_n9195;
  assign new_n18131 = new_n5604 & new_n9185;
  assign new_n18132 = new_n18131 ^ new_n18130;
  assign new_n18133 = n109 & new_n9184;
  assign new_n18134 = n107 & new_n9189;
  assign new_n18135 = new_n18134 ^ new_n18133;
  assign new_n18136 = new_n18135 ^ new_n18132;
  assign new_n18137 = new_n18136 ^ n63;
  assign new_n18138 = new_n18137 ^ new_n18129;
  assign new_n18139 = new_n18138 ^ new_n18122;
  assign new_n18140 = new_n18139 ^ new_n18114;
  assign new_n18141 = new_n18140 ^ new_n18102;
  assign new_n18142 = new_n18141 ^ new_n18090;
  assign new_n18143 = new_n18028 ^ new_n18024;
  assign new_n18144 = ~new_n18025 & new_n18143;
  assign new_n18145 = new_n18144 ^ new_n17968;
  assign new_n18146 = new_n18145 ^ new_n18142;
  assign new_n18147 = ~new_n5424 & n123;
  assign new_n18148 = ~new_n9405 & new_n5419;
  assign new_n18149 = new_n18148 ^ new_n18147;
  assign new_n18150 = n124 & new_n5418;
  assign new_n18151 = n122 & new_n5648;
  assign new_n18152 = new_n18151 ^ new_n18150;
  assign new_n18153 = new_n18152 ^ new_n18149;
  assign new_n18154 = new_n18153 ^ n48;
  assign new_n18155 = new_n18154 ^ new_n18146;
  assign new_n18156 = new_n18033 ^ new_n18029;
  assign new_n18157 = ~new_n18030 & new_n18156;
  assign new_n18158 = new_n18157 ^ new_n17960;
  assign new_n18159 = new_n18158 ^ new_n18155;
  assign new_n18160 = new_n18159 ^ new_n18078;
  assign new_n18161 = new_n18160 ^ new_n18070;
  assign new_n18162 = new_n18049 ^ new_n18039;
  assign new_n18163 = ~new_n18043 & new_n18162;
  assign new_n18164 = new_n18163 ^ new_n18042;
  assign new_n18165 = new_n18164 ^ new_n18161;
  assign new_n18166 = new_n18165 ^ new_n18062;
  assign new_n18167 = ~new_n4804 & n127;
  assign new_n18168 = new_n4799 & new_n10581;
  assign new_n18169 = new_n18168 ^ new_n18167;
  assign new_n18170 = n128 & new_n4798;
  assign new_n18171 = n126 & new_n4810;
  assign new_n18172 = new_n18171 ^ new_n18170;
  assign new_n18173 = new_n18172 ^ new_n18169;
  assign new_n18174 = new_n18173 ^ n45;
  assign new_n18175 = ~new_n5424 & n124;
  assign new_n18176 = new_n5419 & new_n9700;
  assign new_n18177 = new_n18176 ^ new_n18175;
  assign new_n18178 = n125 & new_n5418;
  assign new_n18179 = n123 & new_n5648;
  assign new_n18180 = new_n18179 ^ new_n18178;
  assign new_n18181 = new_n18180 ^ new_n18177;
  assign new_n18182 = new_n18181 ^ n48;
  assign new_n18183 = ~new_n6110 & n121;
  assign new_n18184 = new_n6105 & new_n8850;
  assign new_n18185 = new_n18184 ^ new_n18183;
  assign new_n18186 = n122 & new_n6104;
  assign new_n18187 = n120 & new_n6347;
  assign new_n18188 = new_n18187 ^ new_n18186;
  assign new_n18189 = new_n18188 ^ new_n18185;
  assign new_n18190 = new_n18189 ^ n51;
  assign new_n18191 = new_n18141 ^ new_n18086;
  assign new_n18192 = new_n18090 & new_n18191;
  assign new_n18193 = new_n18192 ^ new_n18089;
  assign new_n18194 = new_n18193 ^ new_n18190;
  assign new_n18195 = ~new_n6805 & n118;
  assign new_n18196 = ~new_n8019 & new_n6800;
  assign new_n18197 = new_n18196 ^ new_n18195;
  assign new_n18198 = n119 & new_n6799;
  assign new_n18199 = n117 & new_n6811;
  assign new_n18200 = new_n18199 ^ new_n18198;
  assign new_n18201 = new_n18200 ^ new_n18197;
  assign new_n18202 = new_n18201 ^ n54;
  assign new_n18203 = new_n18140 ^ new_n18101;
  assign new_n18204 = new_n18102 & new_n18203;
  assign new_n18205 = new_n18204 ^ new_n18098;
  assign new_n18206 = new_n18205 ^ new_n18202;
  assign new_n18207 = n115 & new_n7553;
  assign new_n18208 = ~new_n7256 & new_n7543;
  assign new_n18209 = new_n18208 ^ new_n18207;
  assign new_n18210 = n116 & new_n7542;
  assign new_n18211 = n114 & new_n7547;
  assign new_n18212 = new_n18211 ^ new_n18210;
  assign new_n18213 = new_n18212 ^ new_n18209;
  assign new_n18214 = new_n18213 ^ n57;
  assign new_n18215 = n112 & new_n8355;
  assign new_n18216 = ~new_n6518 & new_n8345;
  assign new_n18217 = new_n18216 ^ new_n18215;
  assign new_n18218 = n113 & new_n8344;
  assign new_n18219 = n111 & new_n8349;
  assign new_n18220 = new_n18219 ^ new_n18218;
  assign new_n18221 = new_n18220 ^ new_n18217;
  assign new_n18222 = new_n18221 ^ n60;
  assign new_n18223 = n109 & new_n9195;
  assign new_n18224 = new_n5825 & new_n9185;
  assign new_n18225 = new_n18224 ^ new_n18223;
  assign new_n18226 = n110 & new_n9184;
  assign new_n18227 = n108 & new_n9189;
  assign new_n18228 = new_n18227 ^ new_n18226;
  assign new_n18229 = new_n18228 ^ new_n18225;
  assign new_n18230 = new_n18229 ^ n63;
  assign new_n18231 = new_n18126 ^ new_n18015;
  assign new_n18232 = ~new_n18231 & new_n18128;
  assign new_n18233 = new_n18232 ^ new_n18015;
  assign new_n18234 = new_n18233 ^ new_n18230;
  assign new_n18235 = n64 & n106;
  assign new_n18236 = new_n18235 ^ n107;
  assign new_n18237 = ~new_n9495 & new_n18236;
  assign new_n18238 = new_n18237 ^ n107;
  assign new_n18239 = new_n18238 ^ new_n18015;
  assign new_n18240 = new_n18239 ^ n42;
  assign new_n18241 = new_n18240 ^ new_n18234;
  assign new_n18242 = new_n18241 ^ new_n18222;
  assign new_n18243 = new_n18129 ^ new_n18122;
  assign new_n18244 = ~new_n18138 & new_n18243;
  assign new_n18245 = new_n18244 ^ new_n18122;
  assign new_n18246 = new_n18245 ^ new_n18242;
  assign new_n18247 = new_n18246 ^ new_n18214;
  assign new_n18248 = new_n18139 ^ new_n18113;
  assign new_n18249 = ~new_n18114 & new_n18248;
  assign new_n18250 = new_n18249 ^ new_n18110;
  assign new_n18251 = new_n18250 ^ new_n18247;
  assign new_n18252 = new_n18251 ^ new_n18206;
  assign new_n18253 = new_n18252 ^ new_n18194;
  assign new_n18254 = new_n18253 ^ new_n18182;
  assign new_n18255 = new_n18154 ^ new_n18142;
  assign new_n18256 = ~new_n18146 & new_n18255;
  assign new_n18257 = new_n18256 ^ new_n18145;
  assign new_n18258 = new_n18257 ^ new_n18254;
  assign new_n18259 = new_n18258 ^ new_n18174;
  assign new_n18260 = new_n18158 ^ new_n18078;
  assign new_n18261 = new_n18159 & new_n18260;
  assign new_n18262 = new_n18261 ^ new_n18078;
  assign new_n18263 = new_n18262 ^ new_n18259;
  assign new_n18264 = new_n18160 ^ new_n18066;
  assign new_n18265 = ~new_n18160 & new_n18066;
  assign new_n18266 = new_n18069 & new_n18265;
  assign new_n18267 = new_n18266 ^ new_n18264;
  assign new_n18268 = new_n18070 & new_n18264;
  assign new_n18269 = new_n18268 ^ new_n18267;
  assign new_n18270 = ~new_n18164 & new_n18269;
  assign new_n18271 = new_n18164 & new_n18266;
  assign new_n18272 = new_n18271 ^ new_n18270;
  assign new_n18273 = new_n18268 ^ new_n18069;
  assign new_n18274 = new_n18266 ^ new_n18164;
  assign new_n18275 = new_n18274 ^ new_n18271;
  assign new_n18276 = new_n18273 & new_n18275;
  assign new_n18277 = new_n18276 ^ new_n18165;
  assign new_n18278 = new_n18277 ^ new_n18272;
  assign new_n18279 = new_n18278 ^ new_n18276;
  assign new_n18280 = ~new_n18062 & ~new_n18279;
  assign new_n18281 = new_n18280 ^ new_n18278;
  assign new_n18282 = ~new_n18272 & new_n18281;
  assign new_n18283 = new_n18282 ^ new_n18263;
  assign new_n18284 = ~new_n18263 & ~new_n18276;
  assign new_n18285 = ~new_n18270 & ~new_n18284;
  assign new_n18286 = ~new_n18062 & new_n18285;
  assign new_n18287 = new_n18263 & new_n18278;
  assign new_n18288 = ~new_n18271 & ~new_n18287;
  assign new_n18289 = ~new_n18286 & new_n18288;
  assign new_n18290 = ~new_n5424 & n125;
  assign new_n18291 = new_n5419 & new_n9987;
  assign new_n18292 = new_n18291 ^ new_n18290;
  assign new_n18293 = n126 & new_n5418;
  assign new_n18294 = n124 & new_n5648;
  assign new_n18295 = new_n18294 ^ new_n18293;
  assign new_n18296 = new_n18295 ^ new_n18292;
  assign new_n18297 = new_n18296 ^ n48;
  assign new_n18298 = new_n18252 ^ new_n18190;
  assign new_n18299 = ~new_n18298 & new_n18194;
  assign new_n18300 = new_n18299 ^ new_n18193;
  assign new_n18301 = new_n18300 ^ new_n18297;
  assign new_n18302 = ~new_n6805 & n119;
  assign new_n18303 = new_n6800 & new_n8286;
  assign new_n18304 = new_n18303 ^ new_n18302;
  assign new_n18305 = n120 & new_n6799;
  assign new_n18306 = n118 & new_n6811;
  assign new_n18307 = new_n18306 ^ new_n18305;
  assign new_n18308 = new_n18307 ^ new_n18304;
  assign new_n18309 = new_n18308 ^ n54;
  assign new_n18310 = n116 & new_n7553;
  assign new_n18311 = ~new_n7503 & new_n7543;
  assign new_n18312 = new_n18311 ^ new_n18310;
  assign new_n18313 = n117 & new_n7542;
  assign new_n18314 = n115 & new_n7547;
  assign new_n18315 = new_n18314 ^ new_n18313;
  assign new_n18316 = new_n18315 ^ new_n18312;
  assign new_n18317 = new_n18316 ^ n57;
  assign new_n18318 = new_n18245 ^ new_n18222;
  assign new_n18319 = ~new_n18242 & new_n18318;
  assign new_n18320 = new_n18319 ^ new_n18245;
  assign new_n18321 = new_n18320 ^ new_n18317;
  assign new_n18322 = n113 & new_n8355;
  assign new_n18323 = ~new_n6764 & new_n8345;
  assign new_n18324 = new_n18323 ^ new_n18322;
  assign new_n18325 = n114 & new_n8344;
  assign new_n18326 = n112 & new_n8349;
  assign new_n18327 = new_n18326 ^ new_n18325;
  assign new_n18328 = new_n18327 ^ new_n18324;
  assign new_n18329 = new_n18328 ^ n60;
  assign new_n18330 = new_n18240 ^ new_n18230;
  assign new_n18331 = ~new_n18234 & new_n18330;
  assign new_n18332 = new_n18331 ^ new_n18233;
  assign new_n18333 = new_n18332 ^ new_n18329;
  assign new_n18334 = n110 & new_n9195;
  assign new_n18335 = new_n6049 & new_n9185;
  assign new_n18336 = new_n18335 ^ new_n18334;
  assign new_n18337 = n111 & new_n9184;
  assign new_n18338 = n109 & new_n9189;
  assign new_n18339 = new_n18338 ^ new_n18337;
  assign new_n18340 = new_n18339 ^ new_n18336;
  assign new_n18341 = new_n18340 ^ n63;
  assign new_n18342 = n64 & n107;
  assign new_n18343 = new_n18342 ^ n108;
  assign new_n18344 = ~new_n9495 & new_n18343;
  assign new_n18345 = new_n18344 ^ n108;
  assign new_n18346 = new_n18015 ^ n42;
  assign new_n18347 = ~new_n18239 & ~new_n18346;
  assign new_n18348 = new_n18347 ^ n42;
  assign new_n18349 = new_n18348 ^ new_n18345;
  assign new_n18350 = new_n18349 ^ new_n18341;
  assign new_n18351 = new_n18350 ^ new_n18333;
  assign new_n18352 = new_n18351 ^ new_n18321;
  assign new_n18353 = new_n18352 ^ new_n18309;
  assign new_n18354 = new_n18250 ^ new_n18214;
  assign new_n18355 = ~new_n18247 & new_n18354;
  assign new_n18356 = new_n18355 ^ new_n18250;
  assign new_n18357 = new_n18356 ^ new_n18353;
  assign new_n18358 = new_n18251 ^ new_n18202;
  assign new_n18359 = ~new_n18358 & new_n18206;
  assign new_n18360 = new_n18359 ^ new_n18205;
  assign new_n18361 = new_n18360 ^ new_n18357;
  assign new_n18362 = ~new_n6110 & n122;
  assign new_n18363 = ~new_n9116 & new_n6105;
  assign new_n18364 = new_n18363 ^ new_n18362;
  assign new_n18365 = n123 & new_n6104;
  assign new_n18366 = n121 & new_n6347;
  assign new_n18367 = new_n18366 ^ new_n18365;
  assign new_n18368 = new_n18367 ^ new_n18364;
  assign new_n18369 = new_n18368 ^ n51;
  assign new_n18370 = new_n18369 ^ new_n18361;
  assign new_n18371 = new_n18370 ^ new_n18301;
  assign new_n18372 = new_n18257 ^ new_n18182;
  assign new_n18373 = ~new_n18254 & new_n18372;
  assign new_n18374 = new_n18373 ^ new_n18257;
  assign new_n18375 = new_n18374 ^ new_n18371;
  assign new_n18376 = n127 & new_n4810;
  assign new_n18377 = new_n4799 & new_n10010;
  assign new_n18378 = new_n18377 ^ new_n18376;
  assign new_n18379 = ~new_n4804 & n128;
  assign new_n18380 = new_n18379 ^ new_n18378;
  assign new_n18381 = new_n18380 ^ n45;
  assign new_n18382 = new_n18381 ^ new_n18375;
  assign new_n18383 = new_n18262 ^ new_n18174;
  assign new_n18384 = ~new_n18259 & new_n18383;
  assign new_n18385 = new_n18384 ^ new_n18262;
  assign new_n18386 = new_n18385 ^ new_n18382;
  assign new_n18387 = new_n18386 ^ new_n18289;
  assign new_n18388 = ~new_n4809 & n128;
  assign new_n18389 = ~n45 & ~new_n18388;
  assign new_n18390 = new_n18389 ^ n44;
  assign new_n18391 = new_n4409 & new_n11133;
  assign new_n18392 = new_n18391 ^ new_n18388;
  assign new_n18393 = ~new_n18390 & ~new_n18392;
  assign new_n18394 = new_n18393 ^ n44;
  assign new_n18395 = new_n18370 ^ new_n18300;
  assign new_n18396 = new_n18301 & new_n18395;
  assign new_n18397 = new_n18396 ^ new_n18297;
  assign new_n18398 = new_n18397 ^ new_n18394;
  assign new_n18399 = ~new_n5424 & n126;
  assign new_n18400 = new_n5419 & new_n10304;
  assign new_n18401 = new_n18400 ^ new_n18399;
  assign new_n18402 = n127 & new_n5418;
  assign new_n18403 = n125 & new_n5648;
  assign new_n18404 = new_n18403 ^ new_n18402;
  assign new_n18405 = new_n18404 ^ new_n18401;
  assign new_n18406 = new_n18405 ^ n48;
  assign new_n18407 = ~new_n6110 & n123;
  assign new_n18408 = ~new_n9405 & new_n6105;
  assign new_n18409 = new_n18408 ^ new_n18407;
  assign new_n18410 = n124 & new_n6104;
  assign new_n18411 = n122 & new_n6347;
  assign new_n18412 = new_n18411 ^ new_n18410;
  assign new_n18413 = new_n18412 ^ new_n18409;
  assign new_n18414 = new_n18413 ^ n51;
  assign new_n18415 = ~new_n6805 & n120;
  assign new_n18416 = new_n6800 & new_n8560;
  assign new_n18417 = new_n18416 ^ new_n18415;
  assign new_n18418 = n121 & new_n6799;
  assign new_n18419 = n119 & new_n6811;
  assign new_n18420 = new_n18419 ^ new_n18418;
  assign new_n18421 = new_n18420 ^ new_n18417;
  assign new_n18422 = new_n18421 ^ n54;
  assign new_n18423 = n117 & new_n7553;
  assign new_n18424 = ~new_n7761 & new_n7543;
  assign new_n18425 = new_n18424 ^ new_n18423;
  assign new_n18426 = n118 & new_n7542;
  assign new_n18427 = n116 & new_n7547;
  assign new_n18428 = new_n18427 ^ new_n18426;
  assign new_n18429 = new_n18428 ^ new_n18425;
  assign new_n18430 = new_n18429 ^ n57;
  assign new_n18431 = n114 & new_n8355;
  assign new_n18432 = ~new_n7013 & new_n8345;
  assign new_n18433 = new_n18432 ^ new_n18431;
  assign new_n18434 = n115 & new_n8344;
  assign new_n18435 = n113 & new_n8349;
  assign new_n18436 = new_n18435 ^ new_n18434;
  assign new_n18437 = new_n18436 ^ new_n18433;
  assign new_n18438 = new_n18437 ^ n60;
  assign new_n18439 = n111 & new_n9195;
  assign new_n18440 = ~new_n6284 & new_n9185;
  assign new_n18441 = new_n18440 ^ new_n18439;
  assign new_n18442 = n112 & new_n9184;
  assign new_n18443 = n110 & new_n9189;
  assign new_n18444 = new_n18443 ^ new_n18442;
  assign new_n18445 = new_n18444 ^ new_n18441;
  assign new_n18446 = new_n5177 ^ n63;
  assign new_n18447 = n64 & new_n4974;
  assign new_n18448 = new_n18447 ^ new_n5177;
  assign new_n18449 = ~new_n9495 & new_n18448;
  assign new_n18450 = new_n18449 ^ new_n18446;
  assign new_n18451 = new_n18450 ^ new_n18445;
  assign new_n18452 = new_n18348 ^ new_n18341;
  assign new_n18453 = ~new_n18349 & ~new_n18452;
  assign new_n18454 = new_n18453 ^ new_n18341;
  assign new_n18455 = new_n18454 ^ new_n18451;
  assign new_n18456 = new_n18455 ^ new_n18438;
  assign new_n18457 = new_n18456 ^ new_n18430;
  assign new_n18458 = new_n18350 ^ new_n18332;
  assign new_n18459 = ~new_n18333 & new_n18458;
  assign new_n18460 = new_n18459 ^ new_n18329;
  assign new_n18461 = new_n18460 ^ new_n18457;
  assign new_n18462 = new_n18461 ^ new_n18422;
  assign new_n18463 = new_n18351 ^ new_n18320;
  assign new_n18464 = new_n18321 & new_n18463;
  assign new_n18465 = new_n18464 ^ new_n18317;
  assign new_n18466 = new_n18465 ^ new_n18462;
  assign new_n18467 = new_n18466 ^ new_n18414;
  assign new_n18468 = new_n18356 ^ new_n18352;
  assign new_n18469 = ~new_n18353 & new_n18468;
  assign new_n18470 = new_n18469 ^ new_n18309;
  assign new_n18471 = new_n18470 ^ new_n18467;
  assign new_n18472 = new_n18471 ^ new_n18406;
  assign new_n18473 = new_n18369 ^ new_n18357;
  assign new_n18474 = ~new_n18361 & new_n18473;
  assign new_n18475 = new_n18474 ^ new_n18360;
  assign new_n18476 = new_n18475 ^ new_n18472;
  assign new_n18477 = new_n18476 ^ new_n18398;
  assign new_n18478 = new_n18381 ^ new_n18371;
  assign new_n18479 = ~new_n18375 & new_n18478;
  assign new_n18480 = new_n18479 ^ new_n18374;
  assign new_n18481 = new_n18480 ^ new_n18477;
  assign new_n18482 = new_n18382 ^ new_n18289;
  assign new_n18483 = ~new_n18386 & ~new_n18482;
  assign new_n18484 = new_n18483 ^ new_n18385;
  assign new_n18485 = new_n18484 ^ new_n18481;
  assign new_n18486 = new_n18397 & new_n18480;
  assign new_n18487 = new_n18480 ^ new_n18397;
  assign new_n18488 = new_n18487 ^ new_n18486;
  assign new_n18489 = new_n18476 ^ new_n18394;
  assign new_n18490 = ~new_n18476 & new_n18394;
  assign new_n18491 = new_n18490 ^ new_n18489;
  assign new_n18492 = ~new_n18488 & new_n18491;
  assign new_n18493 = new_n18486 ^ new_n18484;
  assign new_n18494 = new_n18491 ^ new_n18486;
  assign new_n18495 = ~new_n18493 & new_n18494;
  assign new_n18496 = new_n18495 ^ new_n18492;
  assign new_n18497 = new_n18486 & new_n18490;
  assign new_n18498 = new_n18488 ^ new_n18484;
  assign new_n18499 = new_n18490 ^ new_n18488;
  assign new_n18500 = ~new_n18498 & ~new_n18499;
  assign new_n18501 = new_n18500 ^ new_n18497;
  assign new_n18502 = new_n18501 ^ new_n18496;
  assign new_n18503 = ~new_n5424 & n127;
  assign new_n18504 = new_n5419 & new_n10581;
  assign new_n18505 = new_n18504 ^ new_n18503;
  assign new_n18506 = n128 & new_n5418;
  assign new_n18507 = n126 & new_n5648;
  assign new_n18508 = new_n18507 ^ new_n18506;
  assign new_n18509 = new_n18508 ^ new_n18505;
  assign new_n18510 = new_n18509 ^ n48;
  assign new_n18511 = ~new_n6110 & n124;
  assign new_n18512 = new_n6105 & new_n9700;
  assign new_n18513 = new_n18512 ^ new_n18511;
  assign new_n18514 = n125 & new_n6104;
  assign new_n18515 = n123 & new_n6347;
  assign new_n18516 = new_n18515 ^ new_n18514;
  assign new_n18517 = new_n18516 ^ new_n18513;
  assign new_n18518 = new_n18517 ^ n51;
  assign new_n18519 = ~new_n6805 & n121;
  assign new_n18520 = new_n6800 & new_n8850;
  assign new_n18521 = new_n18520 ^ new_n18519;
  assign new_n18522 = n122 & new_n6799;
  assign new_n18523 = n120 & new_n6811;
  assign new_n18524 = new_n18523 ^ new_n18522;
  assign new_n18525 = new_n18524 ^ new_n18521;
  assign new_n18526 = new_n18525 ^ n54;
  assign new_n18527 = new_n18465 ^ new_n18461;
  assign new_n18528 = ~new_n18462 & new_n18527;
  assign new_n18529 = new_n18528 ^ new_n18422;
  assign new_n18530 = new_n18529 ^ new_n18526;
  assign new_n18531 = n115 & new_n8355;
  assign new_n18532 = ~new_n7256 & new_n8345;
  assign new_n18533 = new_n18532 ^ new_n18531;
  assign new_n18534 = n116 & new_n8344;
  assign new_n18535 = n114 & new_n8349;
  assign new_n18536 = new_n18535 ^ new_n18534;
  assign new_n18537 = new_n18536 ^ new_n18533;
  assign new_n18538 = new_n18537 ^ n60;
  assign new_n18539 = new_n18454 ^ new_n18438;
  assign new_n18540 = new_n18455 & new_n18539;
  assign new_n18541 = new_n18540 ^ new_n18438;
  assign new_n18542 = new_n18541 ^ new_n18538;
  assign new_n18543 = ~n109 & n108;
  assign new_n18544 = new_n18543 ^ new_n5177;
  assign new_n18545 = ~new_n18544 & new_n11491;
  assign new_n18546 = ~n63 & ~n64;
  assign new_n18547 = new_n18546 ^ n63;
  assign new_n18548 = ~new_n18547 & new_n18544;
  assign new_n18549 = new_n18548 ^ n63;
  assign new_n18550 = new_n18549 ^ new_n18545;
  assign new_n18551 = new_n18549 ^ new_n18543;
  assign new_n18552 = new_n18549 ^ new_n18445;
  assign new_n18553 = ~new_n18552 & new_n18549;
  assign new_n18554 = new_n18553 ^ new_n18549;
  assign new_n18555 = new_n18551 & new_n18554;
  assign new_n18556 = new_n18555 ^ new_n18553;
  assign new_n18557 = new_n18556 ^ new_n18549;
  assign new_n18558 = new_n18557 ^ new_n18445;
  assign new_n18559 = ~new_n18550 & ~new_n18558;
  assign new_n18560 = new_n18559 ^ new_n18545;
  assign new_n18561 = new_n18445 ^ n108;
  assign new_n18562 = ~new_n4974 & ~new_n18561;
  assign new_n18563 = new_n18562 ^ n108;
  assign new_n18564 = new_n18563 ^ new_n18543;
  assign new_n18565 = ~new_n18564 & n63;
  assign new_n18566 = new_n18565 ^ new_n18543;
  assign new_n18567 = n64 & new_n18566;
  assign new_n18568 = ~new_n18560 & ~new_n18567;
  assign new_n18569 = n112 & new_n9195;
  assign new_n18570 = ~new_n6518 & new_n9185;
  assign new_n18571 = new_n18570 ^ new_n18569;
  assign new_n18572 = n113 & new_n9184;
  assign new_n18573 = n111 & new_n9189;
  assign new_n18574 = new_n18573 ^ new_n18572;
  assign new_n18575 = new_n18574 ^ new_n18571;
  assign new_n18576 = new_n18575 ^ n63;
  assign new_n18577 = n64 & n109;
  assign new_n18578 = new_n18577 ^ n110;
  assign new_n18579 = ~new_n9495 & new_n18578;
  assign new_n18580 = new_n18579 ^ n110;
  assign new_n18581 = new_n18580 ^ new_n18345;
  assign new_n18582 = new_n18581 ^ n45;
  assign new_n18583 = new_n18582 ^ new_n18576;
  assign new_n18584 = new_n18583 ^ new_n18568;
  assign new_n18585 = new_n18584 ^ new_n18542;
  assign new_n18586 = n118 & new_n7553;
  assign new_n18587 = ~new_n8019 & new_n7543;
  assign new_n18588 = new_n18587 ^ new_n18586;
  assign new_n18589 = n119 & new_n7542;
  assign new_n18590 = n117 & new_n7547;
  assign new_n18591 = new_n18590 ^ new_n18589;
  assign new_n18592 = new_n18591 ^ new_n18588;
  assign new_n18593 = new_n18592 ^ n57;
  assign new_n18594 = new_n18593 ^ new_n18585;
  assign new_n18595 = new_n18460 ^ new_n18456;
  assign new_n18596 = ~new_n18457 & new_n18595;
  assign new_n18597 = new_n18596 ^ new_n18430;
  assign new_n18598 = new_n18597 ^ new_n18594;
  assign new_n18599 = new_n18598 ^ new_n18530;
  assign new_n18600 = new_n18599 ^ new_n18518;
  assign new_n18601 = new_n18470 ^ new_n18466;
  assign new_n18602 = ~new_n18467 & new_n18601;
  assign new_n18603 = new_n18602 ^ new_n18414;
  assign new_n18604 = new_n18603 ^ new_n18600;
  assign new_n18605 = new_n18604 ^ new_n18510;
  assign new_n18606 = new_n18475 ^ new_n18471;
  assign new_n18607 = ~new_n18472 & new_n18606;
  assign new_n18608 = new_n18607 ^ new_n18406;
  assign new_n18609 = new_n18608 ^ new_n18605;
  assign new_n18610 = new_n18609 ^ new_n18502;
  assign new_n18611 = ~new_n18609 & new_n18488;
  assign new_n18612 = ~new_n18490 & ~new_n18611;
  assign new_n18613 = ~new_n18484 & new_n18612;
  assign new_n18614 = new_n18486 ^ new_n18476;
  assign new_n18615 = ~new_n18489 & new_n18614;
  assign new_n18616 = new_n18615 ^ new_n18394;
  assign new_n18617 = ~new_n18616 & new_n18609;
  assign new_n18618 = ~new_n18613 & ~new_n18617;
  assign new_n18619 = ~new_n18491 & ~new_n18609;
  assign new_n18620 = new_n18484 ^ new_n18480;
  assign new_n18621 = new_n18487 & new_n18620;
  assign new_n18622 = new_n18621 ^ new_n18480;
  assign new_n18623 = ~new_n18619 & ~new_n18622;
  assign new_n18624 = ~new_n18623 & new_n18618;
  assign new_n18625 = n127 & new_n5648;
  assign new_n18626 = new_n5419 & new_n10010;
  assign new_n18627 = new_n18626 ^ new_n18625;
  assign new_n18628 = ~new_n5424 & n128;
  assign new_n18629 = new_n18628 ^ new_n18627;
  assign new_n18630 = new_n18629 ^ n48;
  assign new_n18631 = ~new_n6110 & n125;
  assign new_n18632 = new_n6105 & new_n9987;
  assign new_n18633 = new_n18632 ^ new_n18631;
  assign new_n18634 = n126 & new_n6104;
  assign new_n18635 = n124 & new_n6347;
  assign new_n18636 = new_n18635 ^ new_n18634;
  assign new_n18637 = new_n18636 ^ new_n18633;
  assign new_n18638 = new_n18637 ^ n51;
  assign new_n18639 = ~new_n6805 & n122;
  assign new_n18640 = ~new_n9116 & new_n6800;
  assign new_n18641 = new_n18640 ^ new_n18639;
  assign new_n18642 = n123 & new_n6799;
  assign new_n18643 = n121 & new_n6811;
  assign new_n18644 = new_n18643 ^ new_n18642;
  assign new_n18645 = new_n18644 ^ new_n18641;
  assign new_n18646 = new_n18645 ^ n54;
  assign new_n18647 = n119 & new_n7553;
  assign new_n18648 = new_n7543 & new_n8286;
  assign new_n18649 = new_n18648 ^ new_n18647;
  assign new_n18650 = n120 & new_n7542;
  assign new_n18651 = n118 & new_n7547;
  assign new_n18652 = new_n18651 ^ new_n18650;
  assign new_n18653 = new_n18652 ^ new_n18649;
  assign new_n18654 = new_n18653 ^ n57;
  assign new_n18655 = n116 & new_n8355;
  assign new_n18656 = ~new_n7503 & new_n8345;
  assign new_n18657 = new_n18656 ^ new_n18655;
  assign new_n18658 = n117 & new_n8344;
  assign new_n18659 = n115 & new_n8349;
  assign new_n18660 = new_n18659 ^ new_n18658;
  assign new_n18661 = new_n18660 ^ new_n18657;
  assign new_n18662 = new_n18661 ^ n60;
  assign new_n18663 = n110 & new_n11492;
  assign new_n18664 = n111 & new_n9495;
  assign new_n18665 = new_n18664 ^ new_n18663;
  assign new_n18666 = n113 & new_n9195;
  assign new_n18667 = ~new_n6764 & new_n9185;
  assign new_n18668 = new_n18667 ^ new_n18666;
  assign new_n18669 = n114 & new_n9184;
  assign new_n18670 = n112 & new_n9189;
  assign new_n18671 = new_n18670 ^ new_n18669;
  assign new_n18672 = new_n18671 ^ new_n18668;
  assign new_n18673 = new_n18672 ^ n63;
  assign new_n18674 = new_n18345 ^ n45;
  assign new_n18675 = ~new_n18581 & ~new_n18674;
  assign new_n18676 = new_n18675 ^ n45;
  assign new_n18677 = new_n18676 ^ new_n18673;
  assign new_n18678 = new_n18677 ^ new_n18665;
  assign new_n18679 = new_n18678 ^ new_n18662;
  assign new_n18680 = new_n18576 ^ new_n18568;
  assign new_n18681 = new_n18583 & new_n18680;
  assign new_n18682 = new_n18681 ^ new_n18568;
  assign new_n18683 = new_n18682 ^ new_n18679;
  assign new_n18684 = new_n18683 ^ new_n18654;
  assign new_n18685 = new_n18584 ^ new_n18538;
  assign new_n18686 = new_n18542 & new_n18685;
  assign new_n18687 = new_n18686 ^ new_n18541;
  assign new_n18688 = new_n18687 ^ new_n18684;
  assign new_n18689 = new_n18688 ^ new_n18646;
  assign new_n18690 = new_n18597 ^ new_n18585;
  assign new_n18691 = ~new_n18690 & new_n18594;
  assign new_n18692 = new_n18691 ^ new_n18597;
  assign new_n18693 = new_n18692 ^ new_n18689;
  assign new_n18694 = new_n18693 ^ new_n18638;
  assign new_n18695 = new_n18598 ^ new_n18526;
  assign new_n18696 = new_n18530 & new_n18695;
  assign new_n18697 = new_n18696 ^ new_n18529;
  assign new_n18698 = new_n18697 ^ new_n18694;
  assign new_n18699 = new_n18698 ^ new_n18630;
  assign new_n18700 = new_n18603 ^ new_n18518;
  assign new_n18701 = new_n18600 & new_n18700;
  assign new_n18702 = new_n18701 ^ new_n18603;
  assign new_n18703 = new_n18702 ^ new_n18699;
  assign new_n18704 = new_n18608 ^ new_n18510;
  assign new_n18705 = new_n18605 & new_n18704;
  assign new_n18706 = new_n18705 ^ new_n18608;
  assign new_n18707 = new_n18706 ^ new_n18703;
  assign new_n18708 = new_n18707 ^ new_n18624;
  assign new_n18709 = ~new_n18630 & ~new_n18698;
  assign new_n18710 = new_n18709 ^ new_n18699;
  assign new_n18711 = new_n18706 ^ new_n18702;
  assign new_n18712 = ~new_n18702 & ~new_n18706;
  assign new_n18713 = new_n18712 ^ new_n18711;
  assign new_n18714 = ~new_n18710 & new_n18713;
  assign new_n18715 = new_n18713 ^ new_n18709;
  assign new_n18716 = new_n18709 ^ new_n18624;
  assign new_n18717 = new_n18715 & new_n18716;
  assign new_n18718 = new_n18717 ^ new_n18714;
  assign new_n18719 = ~new_n18712 & new_n18709;
  assign new_n18720 = new_n18712 ^ new_n18710;
  assign new_n18721 = new_n18710 ^ new_n18624;
  assign new_n18722 = new_n18720 & new_n18721;
  assign new_n18723 = new_n18722 ^ new_n18719;
  assign new_n18724 = new_n18723 ^ new_n18718;
  assign new_n18725 = ~new_n6110 & n126;
  assign new_n18726 = new_n6105 & new_n10304;
  assign new_n18727 = new_n18726 ^ new_n18725;
  assign new_n18728 = n127 & new_n6104;
  assign new_n18729 = n125 & new_n6347;
  assign new_n18730 = new_n18729 ^ new_n18728;
  assign new_n18731 = new_n18730 ^ new_n18727;
  assign new_n18732 = new_n18731 ^ n51;
  assign new_n18733 = ~new_n6805 & n123;
  assign new_n18734 = ~new_n9405 & new_n6800;
  assign new_n18735 = new_n18734 ^ new_n18733;
  assign new_n18736 = n124 & new_n6799;
  assign new_n18737 = n122 & new_n6811;
  assign new_n18738 = new_n18737 ^ new_n18736;
  assign new_n18739 = new_n18738 ^ new_n18735;
  assign new_n18740 = new_n18739 ^ n54;
  assign new_n18741 = n120 & new_n7553;
  assign new_n18742 = new_n7543 & new_n8560;
  assign new_n18743 = new_n18742 ^ new_n18741;
  assign new_n18744 = n121 & new_n7542;
  assign new_n18745 = n119 & new_n7547;
  assign new_n18746 = new_n18745 ^ new_n18744;
  assign new_n18747 = new_n18746 ^ new_n18743;
  assign new_n18748 = new_n18747 ^ n57;
  assign new_n18749 = new_n18682 ^ new_n18678;
  assign new_n18750 = ~new_n18749 & new_n18679;
  assign new_n18751 = new_n18750 ^ new_n18662;
  assign new_n18752 = new_n18751 ^ new_n18748;
  assign new_n18753 = n117 & new_n8355;
  assign new_n18754 = ~new_n7761 & new_n8345;
  assign new_n18755 = new_n18754 ^ new_n18753;
  assign new_n18756 = n118 & new_n8344;
  assign new_n18757 = n116 & new_n8349;
  assign new_n18758 = new_n18757 ^ new_n18756;
  assign new_n18759 = new_n18758 ^ new_n18755;
  assign new_n18760 = new_n18759 ^ n60;
  assign new_n18761 = n114 & new_n9195;
  assign new_n18762 = ~new_n7013 & new_n9185;
  assign new_n18763 = new_n18762 ^ new_n18761;
  assign new_n18764 = n115 & new_n9184;
  assign new_n18765 = n113 & new_n9189;
  assign new_n18766 = new_n18765 ^ new_n18764;
  assign new_n18767 = new_n18766 ^ new_n18763;
  assign new_n18768 = new_n18767 ^ n63;
  assign new_n18769 = new_n18768 ^ new_n18760;
  assign new_n18770 = new_n18676 ^ new_n18665;
  assign new_n18771 = ~new_n18677 & ~new_n18770;
  assign new_n18772 = new_n18771 ^ new_n18673;
  assign new_n18773 = ~n112 & new_n9495;
  assign new_n18774 = new_n18773 ^ new_n18663;
  assign new_n18775 = n111 & new_n18774;
  assign new_n18776 = new_n18775 ^ new_n18663;
  assign new_n18777 = n112 ^ n111;
  assign new_n18778 = new_n9495 ^ n111;
  assign new_n18779 = new_n11789 ^ n110;
  assign new_n18780 = new_n18779 ^ new_n18774;
  assign new_n18781 = new_n18780 ^ n110;
  assign new_n18782 = new_n18778 & new_n18781;
  assign new_n18783 = new_n18782 ^ new_n18777;
  assign new_n18784 = new_n18783 ^ new_n18776;
  assign new_n18785 = new_n18784 ^ new_n18777;
  assign new_n18786 = new_n18785 ^ new_n18772;
  assign new_n18787 = new_n18786 ^ new_n18769;
  assign new_n18788 = new_n18787 ^ new_n18752;
  assign new_n18789 = new_n18788 ^ new_n18740;
  assign new_n18790 = new_n18687 ^ new_n18683;
  assign new_n18791 = ~new_n18790 & new_n18684;
  assign new_n18792 = new_n18791 ^ new_n18654;
  assign new_n18793 = new_n18792 ^ new_n18789;
  assign new_n18794 = new_n18793 ^ new_n18732;
  assign new_n18795 = new_n18692 ^ new_n18688;
  assign new_n18796 = ~new_n18795 & new_n18689;
  assign new_n18797 = new_n18796 ^ new_n18646;
  assign new_n18798 = new_n18797 ^ new_n18794;
  assign new_n18799 = ~new_n5647 & n128;
  assign new_n18800 = ~n48 & ~new_n18799;
  assign new_n18801 = new_n18800 ^ n47;
  assign new_n18802 = new_n5015 & new_n11133;
  assign new_n18803 = new_n18802 ^ new_n18799;
  assign new_n18804 = ~new_n18801 & ~new_n18803;
  assign new_n18805 = new_n18804 ^ n47;
  assign new_n18806 = new_n18805 ^ new_n18798;
  assign new_n18807 = new_n18697 ^ new_n18693;
  assign new_n18808 = ~new_n18807 & new_n18694;
  assign new_n18809 = new_n18808 ^ new_n18638;
  assign new_n18810 = new_n18809 ^ new_n18806;
  assign new_n18811 = new_n18810 ^ new_n18724;
  assign new_n18812 = ~new_n18709 & ~new_n18713;
  assign new_n18813 = ~new_n18812 & new_n18810;
  assign new_n18814 = ~new_n18813 & new_n18624;
  assign new_n18815 = ~new_n18712 & ~new_n18810;
  assign new_n18816 = ~new_n18815 & new_n18710;
  assign new_n18817 = ~new_n18814 & new_n18816;
  assign new_n18818 = ~new_n18709 & ~new_n18810;
  assign new_n18819 = new_n18706 ^ new_n18624;
  assign new_n18820 = new_n18711 & new_n18819;
  assign new_n18821 = new_n18820 ^ new_n18706;
  assign new_n18822 = ~new_n18818 & ~new_n18821;
  assign new_n18823 = ~new_n18817 & ~new_n18822;
  assign new_n18824 = new_n18809 ^ new_n18798;
  assign new_n18825 = ~new_n18806 & new_n18824;
  assign new_n18826 = new_n18825 ^ new_n18805;
  assign new_n18827 = new_n18797 ^ new_n18793;
  assign new_n18828 = ~new_n18794 & new_n18827;
  assign new_n18829 = new_n18828 ^ new_n18732;
  assign new_n18830 = new_n18829 ^ new_n18826;
  assign new_n18831 = ~new_n6110 & n127;
  assign new_n18832 = new_n6105 & new_n10581;
  assign new_n18833 = new_n18832 ^ new_n18831;
  assign new_n18834 = n128 & new_n6104;
  assign new_n18835 = n126 & new_n6347;
  assign new_n18836 = new_n18835 ^ new_n18834;
  assign new_n18837 = new_n18836 ^ new_n18833;
  assign new_n18838 = new_n18837 ^ n51;
  assign new_n18839 = ~new_n6805 & n124;
  assign new_n18840 = new_n6800 & new_n9700;
  assign new_n18841 = new_n18840 ^ new_n18839;
  assign new_n18842 = n125 & new_n6799;
  assign new_n18843 = n123 & new_n6811;
  assign new_n18844 = new_n18843 ^ new_n18842;
  assign new_n18845 = new_n18844 ^ new_n18841;
  assign new_n18846 = new_n18845 ^ n54;
  assign new_n18847 = n118 & new_n8355;
  assign new_n18848 = ~new_n8019 & new_n8345;
  assign new_n18849 = new_n18848 ^ new_n18847;
  assign new_n18850 = n119 & new_n8344;
  assign new_n18851 = n117 & new_n8349;
  assign new_n18852 = new_n18851 ^ new_n18850;
  assign new_n18853 = new_n18852 ^ new_n18849;
  assign new_n18854 = new_n18853 ^ n60;
  assign new_n18855 = new_n18786 ^ new_n18768;
  assign new_n18856 = new_n18769 & new_n18855;
  assign new_n18857 = new_n18856 ^ new_n18760;
  assign new_n18858 = new_n18857 ^ new_n18854;
  assign new_n18859 = ~new_n18772 & ~new_n18776;
  assign new_n18860 = ~new_n18782 & ~new_n18859;
  assign new_n18861 = n115 & new_n9195;
  assign new_n18862 = ~new_n7256 & new_n9185;
  assign new_n18863 = new_n18862 ^ new_n18861;
  assign new_n18864 = n116 & new_n9184;
  assign new_n18865 = n114 & new_n9189;
  assign new_n18866 = new_n18865 ^ new_n18864;
  assign new_n18867 = new_n18866 ^ new_n18863;
  assign new_n18868 = new_n18867 ^ n63;
  assign new_n18869 = n113 ^ n111;
  assign new_n18870 = ~new_n11492 & new_n18869;
  assign new_n18871 = new_n18870 ^ n111;
  assign new_n18872 = new_n18871 ^ n112;
  assign new_n18873 = new_n11789 & new_n18872;
  assign new_n18874 = new_n18873 ^ n48;
  assign new_n18875 = new_n18874 ^ new_n18868;
  assign new_n18876 = new_n18875 ^ new_n18860;
  assign new_n18877 = new_n18876 ^ new_n18858;
  assign new_n18878 = n121 & new_n7553;
  assign new_n18879 = new_n7543 & new_n8850;
  assign new_n18880 = new_n18879 ^ new_n18878;
  assign new_n18881 = n122 & new_n7542;
  assign new_n18882 = n120 & new_n7547;
  assign new_n18883 = new_n18882 ^ new_n18881;
  assign new_n18884 = new_n18883 ^ new_n18880;
  assign new_n18885 = new_n18884 ^ n57;
  assign new_n18886 = new_n18885 ^ new_n18877;
  assign new_n18887 = new_n18787 ^ new_n18748;
  assign new_n18888 = new_n18752 & new_n18887;
  assign new_n18889 = new_n18888 ^ new_n18751;
  assign new_n18890 = new_n18889 ^ new_n18886;
  assign new_n18891 = new_n18890 ^ new_n18846;
  assign new_n18892 = new_n18792 ^ new_n18788;
  assign new_n18893 = ~new_n18789 & new_n18892;
  assign new_n18894 = new_n18893 ^ new_n18740;
  assign new_n18895 = new_n18894 ^ new_n18891;
  assign new_n18896 = new_n18895 ^ new_n18838;
  assign new_n18897 = new_n18896 ^ new_n18830;
  assign new_n18898 = new_n18897 ^ new_n18823;
  assign new_n18899 = ~new_n18895 & new_n18838;
  assign new_n18900 = new_n18899 ^ new_n18896;
  assign new_n18901 = new_n18900 ^ new_n18823;
  assign new_n18902 = ~new_n18826 & ~new_n18829;
  assign new_n18903 = new_n18902 ^ new_n18830;
  assign new_n18904 = new_n18902 ^ new_n18900;
  assign new_n18905 = new_n18904 ^ new_n18903;
  assign new_n18906 = ~new_n18901 & new_n18905;
  assign new_n18907 = new_n18906 ^ new_n18903;
  assign new_n18908 = ~new_n18823 & ~new_n18899;
  assign new_n18909 = new_n18908 ^ new_n18907;
  assign new_n18910 = new_n18830 & new_n18899;
  assign new_n18911 = new_n18910 ^ new_n18909;
  assign new_n18912 = ~new_n6805 & n125;
  assign new_n18913 = new_n6800 & new_n9987;
  assign new_n18914 = new_n18913 ^ new_n18912;
  assign new_n18915 = n126 & new_n6799;
  assign new_n18916 = n124 & new_n6811;
  assign new_n18917 = new_n18916 ^ new_n18915;
  assign new_n18918 = new_n18917 ^ new_n18914;
  assign new_n18919 = new_n18918 ^ n54;
  assign new_n18920 = new_n18889 ^ new_n18885;
  assign new_n18921 = ~new_n18886 & ~new_n18920;
  assign new_n18922 = new_n18921 ^ new_n18877;
  assign new_n18923 = new_n18922 ^ new_n18919;
  assign new_n18924 = n122 & new_n7553;
  assign new_n18925 = ~new_n9116 & new_n7543;
  assign new_n18926 = new_n18925 ^ new_n18924;
  assign new_n18927 = n123 & new_n7542;
  assign new_n18928 = n121 & new_n7547;
  assign new_n18929 = new_n18928 ^ new_n18927;
  assign new_n18930 = new_n18929 ^ new_n18926;
  assign new_n18931 = new_n18930 ^ n57;
  assign new_n18932 = new_n18876 ^ new_n18854;
  assign new_n18933 = new_n18858 & new_n18932;
  assign new_n18934 = new_n18933 ^ new_n18857;
  assign new_n18935 = new_n18934 ^ new_n18931;
  assign new_n18936 = n119 & new_n8355;
  assign new_n18937 = new_n8286 & new_n8345;
  assign new_n18938 = new_n18937 ^ new_n18936;
  assign new_n18939 = n120 & new_n8344;
  assign new_n18940 = n118 & new_n8349;
  assign new_n18941 = new_n18940 ^ new_n18939;
  assign new_n18942 = new_n18941 ^ new_n18938;
  assign new_n18943 = new_n18942 ^ n60;
  assign new_n18944 = n116 & new_n9195;
  assign new_n18945 = ~new_n7503 & new_n9185;
  assign new_n18946 = new_n18945 ^ new_n18944;
  assign new_n18947 = n117 & new_n9184;
  assign new_n18948 = n115 & new_n9189;
  assign new_n18949 = new_n18948 ^ new_n18947;
  assign new_n18950 = new_n18949 ^ new_n18946;
  assign new_n18951 = new_n18950 ^ n63;
  assign new_n18952 = n112 ^ n48;
  assign new_n18953 = ~new_n18952 & new_n18872;
  assign new_n18954 = new_n18953 ^ n112;
  assign new_n18955 = new_n11789 & new_n18954;
  assign new_n18956 = n64 & n113;
  assign new_n18957 = new_n18956 ^ n114;
  assign new_n18958 = ~new_n9495 & new_n18957;
  assign new_n18959 = new_n18958 ^ n114;
  assign new_n18960 = new_n18959 ^ new_n18955;
  assign new_n18961 = new_n18960 ^ new_n18951;
  assign new_n18962 = new_n18961 ^ new_n18943;
  assign new_n18963 = new_n18868 ^ new_n18860;
  assign new_n18964 = new_n18875 & new_n18963;
  assign new_n18965 = new_n18964 ^ new_n18860;
  assign new_n18966 = new_n18965 ^ new_n18962;
  assign new_n18967 = new_n18966 ^ new_n18935;
  assign new_n18968 = new_n18967 ^ new_n18923;
  assign new_n18969 = new_n18894 ^ new_n18846;
  assign new_n18970 = new_n18891 & new_n18969;
  assign new_n18971 = new_n18970 ^ new_n18894;
  assign new_n18972 = new_n18971 ^ new_n18968;
  assign new_n18973 = n127 & new_n6347;
  assign new_n18974 = new_n6105 & new_n10010;
  assign new_n18975 = new_n18974 ^ new_n18973;
  assign new_n18976 = ~new_n6110 & n128;
  assign new_n18977 = new_n18976 ^ new_n18975;
  assign new_n18978 = new_n18977 ^ n51;
  assign new_n18979 = new_n18978 ^ new_n18972;
  assign new_n18980 = new_n18979 ^ new_n18911;
  assign new_n18981 = ~new_n18979 & new_n18903;
  assign new_n18982 = ~new_n18900 & ~new_n18981;
  assign new_n18983 = ~new_n18908 & new_n18982;
  assign new_n18984 = ~new_n18899 & ~new_n18979;
  assign new_n18985 = ~new_n18902 & ~new_n18984;
  assign new_n18986 = new_n18823 & new_n18985;
  assign new_n18987 = new_n18900 ^ new_n18829;
  assign new_n18988 = new_n18830 & new_n18987;
  assign new_n18989 = new_n18988 ^ new_n18826;
  assign new_n18990 = new_n18979 & new_n18989;
  assign new_n18991 = ~new_n18986 & ~new_n18990;
  assign new_n18992 = ~new_n18983 & new_n18991;
  assign new_n18993 = ~new_n6805 & n126;
  assign new_n18994 = new_n6800 & new_n10304;
  assign new_n18995 = new_n18994 ^ new_n18993;
  assign new_n18996 = n127 & new_n6799;
  assign new_n18997 = n125 & new_n6811;
  assign new_n18998 = new_n18997 ^ new_n18996;
  assign new_n18999 = new_n18998 ^ new_n18995;
  assign new_n19000 = new_n18999 ^ n54;
  assign new_n19001 = new_n18966 ^ new_n18931;
  assign new_n19002 = new_n18935 & new_n19001;
  assign new_n19003 = new_n19002 ^ new_n18934;
  assign new_n19004 = new_n19003 ^ new_n19000;
  assign new_n19005 = n123 & new_n7553;
  assign new_n19006 = ~new_n9405 & new_n7543;
  assign new_n19007 = new_n19006 ^ new_n19005;
  assign new_n19008 = n124 & new_n7542;
  assign new_n19009 = n122 & new_n7547;
  assign new_n19010 = new_n19009 ^ new_n19008;
  assign new_n19011 = new_n19010 ^ new_n19007;
  assign new_n19012 = new_n19011 ^ n57;
  assign new_n19013 = n120 & new_n8355;
  assign new_n19014 = new_n8345 & new_n8560;
  assign new_n19015 = new_n19014 ^ new_n19013;
  assign new_n19016 = n121 & new_n8344;
  assign new_n19017 = n119 & new_n8349;
  assign new_n19018 = new_n19017 ^ new_n19016;
  assign new_n19019 = new_n19018 ^ new_n19015;
  assign new_n19020 = new_n19019 ^ n60;
  assign new_n19021 = n117 & new_n9195;
  assign new_n19022 = ~new_n7761 & new_n9185;
  assign new_n19023 = new_n19022 ^ new_n19021;
  assign new_n19024 = n118 & new_n9184;
  assign new_n19025 = n116 & new_n9189;
  assign new_n19026 = new_n19025 ^ new_n19024;
  assign new_n19027 = new_n19026 ^ new_n19023;
  assign new_n19028 = n115 ^ n114;
  assign new_n19029 = new_n19028 ^ n63;
  assign new_n19030 = n114 ^ n113;
  assign new_n19031 = n64 & new_n19030;
  assign new_n19032 = new_n19031 ^ new_n19028;
  assign new_n19033 = ~new_n9495 & new_n19032;
  assign new_n19034 = new_n19033 ^ new_n19029;
  assign new_n19035 = new_n19034 ^ new_n19027;
  assign new_n19036 = new_n18955 ^ new_n18951;
  assign new_n19037 = new_n18960 & new_n19036;
  assign new_n19038 = new_n19037 ^ new_n18951;
  assign new_n19039 = new_n19038 ^ new_n19035;
  assign new_n19040 = new_n19039 ^ new_n19020;
  assign new_n19041 = new_n19040 ^ new_n19012;
  assign new_n19042 = new_n18965 ^ new_n18943;
  assign new_n19043 = new_n18962 & new_n19042;
  assign new_n19044 = new_n19043 ^ new_n18965;
  assign new_n19045 = new_n19044 ^ new_n19041;
  assign new_n19046 = new_n19045 ^ new_n19004;
  assign new_n19047 = new_n18978 ^ new_n18968;
  assign new_n19048 = ~new_n19047 & new_n18972;
  assign new_n19049 = new_n19048 ^ new_n18971;
  assign new_n19050 = new_n19049 ^ new_n19046;
  assign new_n19051 = ~new_n6346 & n128;
  assign new_n19052 = ~n51 & ~new_n19051;
  assign new_n19053 = new_n19052 ^ n50;
  assign new_n19054 = new_n5640 & new_n11133;
  assign new_n19055 = new_n19054 ^ new_n19051;
  assign new_n19056 = ~new_n19053 & ~new_n19055;
  assign new_n19057 = new_n19056 ^ n50;
  assign new_n19058 = new_n18967 ^ new_n18922;
  assign new_n19059 = ~new_n18923 & ~new_n19058;
  assign new_n19060 = new_n19059 ^ new_n18919;
  assign new_n19061 = new_n19060 ^ new_n19057;
  assign new_n19062 = new_n19061 ^ new_n19050;
  assign new_n19063 = new_n19062 ^ new_n18992;
  assign new_n19064 = ~new_n19057 & ~new_n19060;
  assign new_n19065 = new_n19064 ^ new_n19061;
  assign new_n19066 = new_n19065 ^ new_n18992;
  assign new_n19067 = ~new_n19046 & new_n19049;
  assign new_n19068 = new_n19067 ^ new_n19050;
  assign new_n19069 = new_n19067 ^ new_n19065;
  assign new_n19070 = new_n19069 ^ new_n19068;
  assign new_n19071 = new_n19066 & new_n19070;
  assign new_n19072 = new_n19071 ^ new_n19068;
  assign new_n19073 = ~new_n18992 & ~new_n19064;
  assign new_n19074 = new_n19073 ^ new_n19072;
  assign new_n19075 = ~new_n19050 & new_n19064;
  assign new_n19076 = new_n19075 ^ new_n19074;
  assign new_n19077 = ~new_n6805 & n127;
  assign new_n19078 = new_n6800 & new_n10581;
  assign new_n19079 = new_n19078 ^ new_n19077;
  assign new_n19080 = n128 & new_n6799;
  assign new_n19081 = n126 & new_n6811;
  assign new_n19082 = new_n19081 ^ new_n19080;
  assign new_n19083 = new_n19082 ^ new_n19079;
  assign new_n19084 = new_n19083 ^ n54;
  assign new_n19085 = n124 & new_n7553;
  assign new_n19086 = new_n7543 & new_n9700;
  assign new_n19087 = new_n19086 ^ new_n19085;
  assign new_n19088 = n125 & new_n7542;
  assign new_n19089 = n123 & new_n7547;
  assign new_n19090 = new_n19089 ^ new_n19088;
  assign new_n19091 = new_n19090 ^ new_n19087;
  assign new_n19092 = new_n19091 ^ n57;
  assign new_n19093 = n121 & new_n8355;
  assign new_n19094 = new_n8345 & new_n8850;
  assign new_n19095 = new_n19094 ^ new_n19093;
  assign new_n19096 = n122 & new_n8344;
  assign new_n19097 = n120 & new_n8349;
  assign new_n19098 = new_n19097 ^ new_n19096;
  assign new_n19099 = new_n19098 ^ new_n19095;
  assign new_n19100 = new_n19099 ^ n60;
  assign new_n19101 = new_n19038 ^ new_n19020;
  assign new_n19102 = new_n19039 & new_n19101;
  assign new_n19103 = new_n19102 ^ new_n19020;
  assign new_n19104 = new_n19103 ^ new_n19100;
  assign new_n19105 = n118 & new_n9195;
  assign new_n19106 = ~new_n8019 & new_n9185;
  assign new_n19107 = new_n19106 ^ new_n19105;
  assign new_n19108 = n119 & new_n9184;
  assign new_n19109 = n117 & new_n9189;
  assign new_n19110 = new_n19109 ^ new_n19108;
  assign new_n19111 = new_n19110 ^ new_n19107;
  assign new_n19112 = new_n19111 ^ n63;
  assign new_n19113 = n64 & n115;
  assign new_n19114 = new_n19113 ^ n116;
  assign new_n19115 = ~new_n9495 & new_n19114;
  assign new_n19116 = new_n19115 ^ n116;
  assign new_n19117 = new_n19116 ^ n51;
  assign new_n19118 = new_n19117 ^ new_n18959;
  assign new_n19119 = new_n19118 ^ new_n19112;
  assign new_n19120 = new_n19027 ^ n63;
  assign new_n19121 = ~n114 & new_n19030;
  assign new_n19122 = n114 & new_n19030;
  assign new_n19123 = new_n19122 ^ new_n19121;
  assign new_n19124 = ~new_n19120 & ~new_n19123;
  assign new_n19125 = new_n19124 ^ new_n19121;
  assign new_n19126 = ~n115 & n114;
  assign new_n19127 = ~n114 & n115;
  assign new_n19128 = new_n19127 ^ new_n19126;
  assign new_n19129 = ~new_n19120 & ~new_n19128;
  assign new_n19130 = new_n19129 ^ new_n19126;
  assign new_n19131 = new_n19130 ^ new_n19125;
  assign new_n19132 = ~new_n9495 & new_n19131;
  assign new_n19133 = new_n19132 ^ new_n19130;
  assign new_n19134 = new_n19130 ^ new_n19120;
  assign new_n19135 = ~new_n9495 & ~new_n19134;
  assign new_n19136 = new_n19135 ^ new_n19130;
  assign new_n19137 = new_n19136 ^ new_n19133;
  assign new_n19138 = ~n63 & new_n19137;
  assign new_n19139 = new_n19138 ^ new_n19133;
  assign new_n19140 = new_n19139 ^ new_n19119;
  assign new_n19141 = new_n19140 ^ new_n19104;
  assign new_n19142 = new_n19141 ^ new_n19092;
  assign new_n19143 = new_n19044 ^ new_n19040;
  assign new_n19144 = ~new_n19041 & new_n19143;
  assign new_n19145 = new_n19144 ^ new_n19012;
  assign new_n19146 = new_n19145 ^ new_n19142;
  assign new_n19147 = new_n19146 ^ new_n19084;
  assign new_n19148 = new_n19045 ^ new_n19003;
  assign new_n19149 = new_n19004 & new_n19148;
  assign new_n19150 = new_n19149 ^ new_n19000;
  assign new_n19151 = new_n19150 ^ new_n19147;
  assign new_n19152 = new_n19151 ^ new_n19076;
  assign new_n19153 = ~new_n19068 & new_n19151;
  assign new_n19154 = ~new_n19153 & new_n19065;
  assign new_n19155 = ~new_n19073 & new_n19154;
  assign new_n19156 = ~new_n19064 & new_n19151;
  assign new_n19157 = ~new_n19067 & ~new_n19156;
  assign new_n19158 = new_n18992 & new_n19157;
  assign new_n19159 = new_n19065 ^ new_n19046;
  assign new_n19160 = ~new_n19050 & ~new_n19159;
  assign new_n19161 = new_n19160 ^ new_n19049;
  assign new_n19162 = ~new_n19151 & ~new_n19161;
  assign new_n19163 = ~new_n19158 & ~new_n19162;
  assign new_n19164 = ~new_n19155 & new_n19163;
  assign new_n19165 = n125 & new_n7553;
  assign new_n19166 = new_n7543 & new_n9987;
  assign new_n19167 = new_n19166 ^ new_n19165;
  assign new_n19168 = n126 & new_n7542;
  assign new_n19169 = n124 & new_n7547;
  assign new_n19170 = new_n19169 ^ new_n19168;
  assign new_n19171 = new_n19170 ^ new_n19167;
  assign new_n19172 = new_n19171 ^ n57;
  assign new_n19173 = new_n19140 ^ new_n19100;
  assign new_n19174 = ~new_n19173 & new_n19104;
  assign new_n19175 = new_n19174 ^ new_n19103;
  assign new_n19176 = new_n19175 ^ new_n19172;
  assign new_n19177 = n122 & new_n8355;
  assign new_n19178 = ~new_n9116 & new_n8345;
  assign new_n19179 = new_n19178 ^ new_n19177;
  assign new_n19180 = n123 & new_n8344;
  assign new_n19181 = n121 & new_n8349;
  assign new_n19182 = new_n19181 ^ new_n19180;
  assign new_n19183 = new_n19182 ^ new_n19179;
  assign new_n19184 = new_n19183 ^ n60;
  assign new_n19185 = n117 & new_n9495;
  assign new_n19186 = n116 & new_n11492;
  assign new_n19187 = new_n19186 ^ new_n19185;
  assign new_n19188 = n119 & new_n9195;
  assign new_n19189 = new_n8286 & new_n9185;
  assign new_n19190 = new_n19189 ^ new_n19188;
  assign new_n19191 = n120 & new_n9184;
  assign new_n19192 = n118 & new_n9189;
  assign new_n19193 = new_n19192 ^ new_n19191;
  assign new_n19194 = new_n19193 ^ new_n19190;
  assign new_n19195 = new_n19194 ^ n63;
  assign new_n19196 = new_n18959 ^ n51;
  assign new_n19197 = new_n19116 ^ new_n18959;
  assign new_n19198 = ~new_n19196 & ~new_n19197;
  assign new_n19199 = new_n19198 ^ n51;
  assign new_n19200 = new_n19199 ^ new_n19195;
  assign new_n19201 = new_n19200 ^ new_n19187;
  assign new_n19202 = new_n19201 ^ new_n19184;
  assign new_n19203 = new_n19139 ^ new_n19112;
  assign new_n19204 = ~new_n19203 & new_n19119;
  assign new_n19205 = new_n19204 ^ new_n19139;
  assign new_n19206 = new_n19205 ^ new_n19202;
  assign new_n19207 = new_n19206 ^ new_n19176;
  assign new_n19208 = new_n19145 ^ new_n19092;
  assign new_n19209 = ~new_n19142 & new_n19208;
  assign new_n19210 = new_n19209 ^ new_n19145;
  assign new_n19211 = new_n19210 ^ new_n19207;
  assign new_n19212 = n127 & new_n6811;
  assign new_n19213 = new_n6800 & new_n10010;
  assign new_n19214 = new_n19213 ^ new_n19212;
  assign new_n19215 = ~new_n6805 & n128;
  assign new_n19216 = new_n19215 ^ new_n19214;
  assign new_n19217 = new_n19216 ^ n54;
  assign new_n19218 = new_n19217 ^ new_n19211;
  assign new_n19219 = new_n19150 ^ new_n19084;
  assign new_n19220 = ~new_n19147 & new_n19219;
  assign new_n19221 = new_n19220 ^ new_n19150;
  assign new_n19222 = new_n19221 ^ new_n19218;
  assign new_n19223 = new_n19222 ^ new_n19164;
  assign new_n19224 = new_n19218 ^ new_n19164;
  assign new_n19225 = ~new_n19222 & new_n19224;
  assign new_n19226 = new_n19225 ^ new_n19221;
  assign new_n19227 = n126 & new_n7553;
  assign new_n19228 = new_n7543 & new_n10304;
  assign new_n19229 = new_n19228 ^ new_n19227;
  assign new_n19230 = n127 & new_n7542;
  assign new_n19231 = n125 & new_n7547;
  assign new_n19232 = new_n19231 ^ new_n19230;
  assign new_n19233 = new_n19232 ^ new_n19229;
  assign new_n19234 = new_n19233 ^ n57;
  assign new_n19235 = n123 & new_n8355;
  assign new_n19236 = ~new_n9405 & new_n8345;
  assign new_n19237 = new_n19236 ^ new_n19235;
  assign new_n19238 = n124 & new_n8344;
  assign new_n19239 = n122 & new_n8349;
  assign new_n19240 = new_n19239 ^ new_n19238;
  assign new_n19241 = new_n19240 ^ new_n19237;
  assign new_n19242 = new_n19241 ^ n60;
  assign new_n19243 = n120 & new_n9195;
  assign new_n19244 = new_n8560 & new_n9185;
  assign new_n19245 = new_n19244 ^ new_n19243;
  assign new_n19246 = n121 & new_n9184;
  assign new_n19247 = n119 & new_n9189;
  assign new_n19248 = new_n19247 ^ new_n19246;
  assign new_n19249 = new_n19248 ^ new_n19245;
  assign new_n19250 = new_n19249 ^ n63;
  assign new_n19251 = new_n19250 ^ new_n19242;
  assign new_n19252 = new_n19199 ^ new_n19187;
  assign new_n19253 = ~new_n19200 & ~new_n19252;
  assign new_n19254 = new_n19253 ^ new_n19195;
  assign new_n19255 = ~n118 & new_n9495;
  assign new_n19256 = new_n19255 ^ new_n19186;
  assign new_n19257 = n117 & new_n19256;
  assign new_n19258 = new_n9495 ^ n117;
  assign new_n19259 = new_n11789 ^ n116;
  assign new_n19260 = new_n19259 ^ new_n19256;
  assign new_n19261 = new_n19260 ^ n116;
  assign new_n19262 = new_n19258 & new_n19261;
  assign new_n19263 = new_n19262 ^ new_n19186;
  assign new_n19264 = new_n19263 ^ new_n19257;
  assign new_n19265 = new_n19264 ^ new_n19254;
  assign new_n19266 = new_n19265 ^ new_n19251;
  assign new_n19267 = new_n19205 ^ new_n19201;
  assign new_n19268 = new_n19202 & new_n19267;
  assign new_n19269 = new_n19268 ^ new_n19184;
  assign new_n19270 = new_n19269 ^ new_n19266;
  assign new_n19271 = new_n19270 ^ new_n19234;
  assign new_n19272 = ~new_n6810 & n128;
  assign new_n19273 = ~n54 & ~new_n19272;
  assign new_n19274 = new_n19273 ^ n53;
  assign new_n19275 = new_n6352 & new_n11133;
  assign new_n19276 = new_n19275 ^ new_n19272;
  assign new_n19277 = ~new_n19274 & ~new_n19276;
  assign new_n19278 = new_n19277 ^ n53;
  assign new_n19279 = new_n19278 ^ new_n19271;
  assign new_n19280 = new_n19206 ^ new_n19175;
  assign new_n19281 = new_n19176 & new_n19280;
  assign new_n19282 = new_n19281 ^ new_n19172;
  assign new_n19283 = new_n19282 ^ new_n19279;
  assign new_n19284 = new_n19217 ^ new_n19207;
  assign new_n19285 = ~new_n19211 & new_n19284;
  assign new_n19286 = new_n19285 ^ new_n19210;
  assign new_n19287 = new_n19286 ^ new_n19283;
  assign new_n19288 = new_n19287 ^ new_n19226;
  assign new_n19289 = new_n19282 ^ new_n19271;
  assign new_n19290 = ~new_n19279 & new_n19289;
  assign new_n19291 = new_n19290 ^ new_n19278;
  assign new_n19292 = new_n19269 ^ new_n19234;
  assign new_n19293 = new_n19270 & new_n19292;
  assign new_n19294 = new_n19293 ^ new_n19234;
  assign new_n19295 = new_n19294 ^ new_n19291;
  assign new_n19296 = n124 & new_n8355;
  assign new_n19297 = new_n8345 & new_n9700;
  assign new_n19298 = new_n19297 ^ new_n19296;
  assign new_n19299 = n125 & new_n8344;
  assign new_n19300 = n123 & new_n8349;
  assign new_n19301 = new_n19300 ^ new_n19299;
  assign new_n19302 = new_n19301 ^ new_n19298;
  assign new_n19303 = new_n19302 ^ n60;
  assign new_n19304 = new_n19265 ^ new_n19250;
  assign new_n19305 = new_n19251 & new_n19304;
  assign new_n19306 = new_n19305 ^ new_n19242;
  assign new_n19307 = new_n19306 ^ new_n19303;
  assign new_n19308 = n121 & new_n9195;
  assign new_n19309 = new_n8850 & new_n9185;
  assign new_n19310 = new_n19309 ^ new_n19308;
  assign new_n19311 = n122 & new_n9184;
  assign new_n19312 = n120 & new_n9189;
  assign new_n19313 = new_n19312 ^ new_n19311;
  assign new_n19314 = new_n19313 ^ new_n19310;
  assign new_n19315 = new_n19314 ^ n63;
  assign new_n19316 = n119 ^ n117;
  assign new_n19317 = ~new_n11492 & new_n19316;
  assign new_n19318 = new_n19317 ^ n117;
  assign new_n19319 = new_n19318 ^ n118;
  assign new_n19320 = new_n11789 & new_n19319;
  assign new_n19321 = new_n19320 ^ n54;
  assign new_n19322 = new_n19321 ^ new_n19315;
  assign new_n19323 = ~new_n19254 & ~new_n19264;
  assign new_n19324 = new_n19323 ^ new_n19262;
  assign new_n19325 = new_n19324 ^ new_n19322;
  assign new_n19326 = new_n19325 ^ new_n19307;
  assign new_n19327 = n127 & new_n7553;
  assign new_n19328 = new_n7543 & new_n10581;
  assign new_n19329 = new_n19328 ^ new_n19327;
  assign new_n19330 = n128 & new_n7542;
  assign new_n19331 = n126 & new_n7547;
  assign new_n19332 = new_n19331 ^ new_n19330;
  assign new_n19333 = new_n19332 ^ new_n19329;
  assign new_n19334 = new_n19333 ^ n57;
  assign new_n19335 = new_n19334 ^ new_n19326;
  assign new_n19336 = new_n19335 ^ new_n19295;
  assign new_n19337 = new_n19283 ^ new_n19226;
  assign new_n19338 = ~new_n19287 & new_n19337;
  assign new_n19339 = new_n19338 ^ new_n19286;
  assign new_n19340 = new_n19339 ^ new_n19336;
  assign new_n19341 = ~new_n19326 & ~new_n19334;
  assign new_n19342 = new_n19341 ^ new_n19335;
  assign new_n19343 = ~new_n19339 & new_n19342;
  assign new_n19344 = ~new_n19291 & ~new_n19294;
  assign new_n19345 = ~new_n19342 & ~new_n19344;
  assign new_n19346 = new_n19344 ^ new_n19295;
  assign new_n19347 = ~new_n19345 & new_n19346;
  assign new_n19348 = ~new_n19341 & ~new_n19347;
  assign new_n19349 = new_n19347 ^ new_n19341;
  assign new_n19350 = new_n19349 ^ new_n19348;
  assign new_n19351 = ~new_n19344 & new_n19350;
  assign new_n19352 = ~new_n19351 & new_n19343;
  assign new_n19353 = new_n19339 & new_n19348;
  assign new_n19354 = new_n19350 ^ new_n19345;
  assign new_n19355 = ~new_n19295 & ~new_n19354;
  assign new_n19356 = ~new_n19353 & ~new_n19355;
  assign new_n19357 = ~new_n19352 & new_n19356;
  assign new_n19358 = n125 & new_n8355;
  assign new_n19359 = new_n8345 & new_n9987;
  assign new_n19360 = new_n19359 ^ new_n19358;
  assign new_n19361 = n126 & new_n8344;
  assign new_n19362 = n124 & new_n8349;
  assign new_n19363 = new_n19362 ^ new_n19361;
  assign new_n19364 = new_n19363 ^ new_n19360;
  assign new_n19365 = new_n19364 ^ n60;
  assign new_n19366 = new_n19324 ^ new_n19315;
  assign new_n19367 = ~new_n19366 & new_n19322;
  assign new_n19368 = new_n19367 ^ new_n19324;
  assign new_n19369 = new_n19368 ^ new_n19365;
  assign new_n19370 = n122 & new_n9195;
  assign new_n19371 = ~new_n9116 & new_n9185;
  assign new_n19372 = new_n19371 ^ new_n19370;
  assign new_n19373 = n123 & new_n9184;
  assign new_n19374 = n121 & new_n9189;
  assign new_n19375 = new_n19374 ^ new_n19373;
  assign new_n19376 = new_n19375 ^ new_n19372;
  assign new_n19377 = new_n19376 ^ n63;
  assign new_n19378 = n119 ^ n64;
  assign new_n19379 = n119 & new_n19378;
  assign new_n19380 = new_n19379 ^ n119;
  assign new_n19381 = new_n19380 ^ n120;
  assign new_n19382 = ~new_n9495 & new_n19381;
  assign new_n19383 = new_n19382 ^ n120;
  assign new_n19384 = n118 ^ n54;
  assign new_n19385 = ~new_n19384 & new_n19319;
  assign new_n19386 = new_n19385 ^ n118;
  assign new_n19387 = new_n11789 & new_n19386;
  assign new_n19388 = new_n19387 ^ new_n19383;
  assign new_n19389 = new_n19388 ^ new_n19377;
  assign new_n19390 = new_n19389 ^ new_n19369;
  assign new_n19391 = new_n19325 ^ new_n19303;
  assign new_n19392 = ~new_n19391 & new_n19307;
  assign new_n19393 = new_n19392 ^ new_n19306;
  assign new_n19394 = new_n19393 ^ new_n19390;
  assign new_n19395 = n127 & new_n7547;
  assign new_n19396 = new_n7543 & new_n10010;
  assign new_n19397 = new_n19396 ^ new_n19395;
  assign new_n19398 = n128 & new_n7553;
  assign new_n19399 = new_n19398 ^ new_n19397;
  assign new_n19400 = new_n19399 ^ n57;
  assign new_n19401 = new_n19400 ^ new_n19394;
  assign new_n19402 = new_n19401 ^ new_n19357;
  assign new_n19403 = ~new_n19401 & new_n19346;
  assign new_n19404 = ~new_n19341 & ~new_n19403;
  assign new_n19405 = ~new_n19343 & new_n19404;
  assign new_n19406 = ~new_n19401 & new_n19342;
  assign new_n19407 = ~new_n19344 & ~new_n19406;
  assign new_n19408 = new_n19339 & new_n19407;
  assign new_n19409 = new_n19351 & new_n19401;
  assign new_n19410 = ~new_n19408 & ~new_n19409;
  assign new_n19411 = ~new_n19405 & new_n19410;
  assign new_n19412 = n126 & new_n8355;
  assign new_n19413 = new_n8345 & new_n10304;
  assign new_n19414 = new_n19413 ^ new_n19412;
  assign new_n19415 = n127 & new_n8344;
  assign new_n19416 = n125 & new_n8349;
  assign new_n19417 = new_n19416 ^ new_n19415;
  assign new_n19418 = new_n19417 ^ new_n19414;
  assign new_n19419 = new_n19418 ^ n60;
  assign new_n19420 = n123 & new_n9195;
  assign new_n19421 = ~new_n9405 & new_n9185;
  assign new_n19422 = new_n19421 ^ new_n19420;
  assign new_n19423 = n124 & new_n9184;
  assign new_n19424 = n122 & new_n9189;
  assign new_n19425 = new_n19424 ^ new_n19423;
  assign new_n19426 = new_n19425 ^ new_n19422;
  assign new_n19427 = new_n19426 ^ n63;
  assign new_n19428 = n121 ^ n120;
  assign new_n19429 = new_n19428 ^ new_n7778;
  assign new_n19430 = new_n19429 ^ n64;
  assign new_n19431 = new_n19430 ^ new_n19429;
  assign new_n19432 = new_n19429 ^ new_n19428;
  assign new_n19433 = ~new_n19431 & new_n19432;
  assign new_n19434 = new_n19433 ^ new_n19429;
  assign new_n19435 = ~new_n9495 & new_n19434;
  assign new_n19436 = new_n19435 ^ new_n19428;
  assign new_n19437 = new_n19436 ^ new_n19427;
  assign new_n19438 = new_n19387 ^ new_n19377;
  assign new_n19439 = new_n19388 & new_n19438;
  assign new_n19440 = new_n19439 ^ new_n19377;
  assign new_n19441 = new_n19440 ^ new_n19437;
  assign new_n19442 = new_n19441 ^ new_n19419;
  assign new_n19443 = new_n19400 ^ new_n19390;
  assign new_n19444 = ~new_n19443 & new_n19394;
  assign new_n19445 = new_n19444 ^ new_n19393;
  assign new_n19446 = new_n19445 ^ new_n19442;
  assign new_n19447 = n128 & new_n7547;
  assign new_n19448 = new_n7543 & new_n11133;
  assign new_n19449 = new_n19448 ^ new_n19447;
  assign new_n19450 = new_n19449 ^ n57;
  assign new_n19451 = new_n19389 ^ new_n19365;
  assign new_n19452 = ~new_n19369 & new_n19451;
  assign new_n19453 = new_n19452 ^ new_n19368;
  assign new_n19454 = new_n19453 ^ new_n19450;
  assign new_n19455 = new_n19454 ^ new_n19446;
  assign new_n19456 = new_n19455 ^ new_n19411;
  assign new_n19457 = ~new_n19450 & new_n19453;
  assign new_n19458 = new_n19457 ^ new_n19454;
  assign new_n19459 = ~new_n19411 & new_n19458;
  assign new_n19460 = new_n19458 ^ new_n19411;
  assign new_n19461 = new_n19460 ^ new_n19459;
  assign new_n19462 = ~new_n19461 & new_n19457;
  assign new_n19463 = n127 & new_n8355;
  assign new_n19464 = new_n8345 & new_n10581;
  assign new_n19465 = new_n19464 ^ new_n19463;
  assign new_n19466 = n128 & new_n8344;
  assign new_n19467 = n126 & new_n8349;
  assign new_n19468 = new_n19467 ^ new_n19466;
  assign new_n19469 = new_n19468 ^ new_n19465;
  assign new_n19470 = new_n19469 ^ n60;
  assign new_n19471 = new_n19440 ^ new_n19419;
  assign new_n19472 = new_n19441 & new_n19471;
  assign new_n19473 = new_n19472 ^ new_n19419;
  assign new_n19474 = new_n19473 ^ new_n19470;
  assign new_n19475 = n124 & new_n9195;
  assign new_n19476 = new_n9185 & new_n9700;
  assign new_n19477 = new_n19476 ^ new_n19475;
  assign new_n19478 = n125 & new_n9184;
  assign new_n19479 = n123 & new_n9189;
  assign new_n19480 = new_n19479 ^ new_n19478;
  assign new_n19481 = new_n19480 ^ new_n19477;
  assign new_n19482 = new_n19481 ^ n63;
  assign new_n19483 = n64 & n121;
  assign new_n19484 = new_n19483 ^ n122;
  assign new_n19485 = ~new_n9495 & new_n19484;
  assign new_n19486 = new_n19485 ^ n122;
  assign new_n19487 = new_n19486 ^ n57;
  assign new_n19488 = new_n19487 ^ new_n19383;
  assign new_n19489 = new_n19488 ^ new_n19482;
  assign new_n19490 = ~n119 & n120;
  assign new_n19491 = new_n19490 ^ new_n8041;
  assign new_n19492 = new_n19491 ^ new_n8041;
  assign new_n19493 = n64 & new_n19492;
  assign new_n19494 = new_n19493 ^ new_n8041;
  assign new_n19495 = ~new_n9495 & new_n19494;
  assign new_n19496 = new_n19495 ^ new_n8041;
  assign new_n19497 = ~new_n19436 & new_n19427;
  assign new_n19498 = new_n19497 ^ new_n19496;
  assign new_n19499 = new_n19498 ^ new_n19489;
  assign new_n19500 = new_n19499 ^ new_n19474;
  assign new_n19501 = new_n19500 ^ new_n19462;
  assign new_n19502 = new_n19446 ^ new_n19411;
  assign new_n19503 = ~new_n19502 & new_n19460;
  assign new_n19504 = new_n19503 ^ new_n19446;
  assign new_n19505 = new_n19457 ^ new_n19442;
  assign new_n19506 = ~new_n19446 & ~new_n19505;
  assign new_n19507 = new_n19506 ^ new_n19445;
  assign new_n19508 = new_n19507 ^ new_n19504;
  assign new_n19509 = new_n19508 ^ new_n19501;
  assign new_n19510 = ~new_n19445 & new_n19442;
  assign new_n19511 = new_n19510 ^ new_n19446;
  assign new_n19512 = ~new_n19511 & new_n19500;
  assign new_n19513 = ~new_n19457 & ~new_n19512;
  assign new_n19514 = ~new_n19461 & new_n19513;
  assign new_n19515 = ~new_n19458 & new_n19500;
  assign new_n19516 = ~new_n19510 & ~new_n19515;
  assign new_n19517 = ~new_n19411 & new_n19516;
  assign new_n19518 = ~new_n19500 & new_n19507;
  assign new_n19519 = ~new_n19517 & ~new_n19518;
  assign new_n19520 = ~new_n19514 & new_n19519;
  assign new_n19521 = n127 & new_n8349;
  assign new_n19522 = new_n8345 & new_n10010;
  assign new_n19523 = new_n19522 ^ new_n19521;
  assign new_n19524 = n128 & new_n8355;
  assign new_n19525 = new_n19524 ^ new_n19523;
  assign new_n19526 = new_n19525 ^ n60;
  assign new_n19527 = n122 & new_n11492;
  assign new_n19528 = n123 & new_n9495;
  assign new_n19529 = new_n19528 ^ new_n19527;
  assign new_n19530 = n125 & new_n9195;
  assign new_n19531 = new_n9185 & new_n9987;
  assign new_n19532 = new_n19531 ^ new_n19530;
  assign new_n19533 = n126 & new_n9184;
  assign new_n19534 = n124 & new_n9189;
  assign new_n19535 = new_n19534 ^ new_n19533;
  assign new_n19536 = new_n19535 ^ new_n19532;
  assign new_n19537 = new_n19536 ^ n63;
  assign new_n19538 = new_n19383 ^ n57;
  assign new_n19539 = new_n19486 ^ new_n19383;
  assign new_n19540 = ~new_n19538 & ~new_n19539;
  assign new_n19541 = new_n19540 ^ n57;
  assign new_n19542 = new_n19541 ^ new_n19537;
  assign new_n19543 = new_n19542 ^ new_n19529;
  assign new_n19544 = new_n19498 ^ new_n19482;
  assign new_n19545 = new_n19489 & new_n19544;
  assign new_n19546 = new_n19545 ^ new_n19498;
  assign new_n19547 = new_n19546 ^ new_n19543;
  assign new_n19548 = new_n19547 ^ new_n19526;
  assign new_n19549 = new_n19499 ^ new_n19470;
  assign new_n19550 = new_n19474 & new_n19549;
  assign new_n19551 = new_n19550 ^ new_n19473;
  assign new_n19552 = new_n19551 ^ new_n19548;
  assign new_n19553 = new_n19552 ^ new_n19520;
  assign new_n19554 = n128 & new_n8349;
  assign new_n19555 = new_n8345 & new_n11133;
  assign new_n19556 = new_n19555 ^ new_n19554;
  assign new_n19557 = new_n19556 ^ n60;
  assign new_n19558 = new_n19546 ^ new_n19526;
  assign new_n19559 = ~new_n19547 & new_n19558;
  assign new_n19560 = new_n19559 ^ new_n19526;
  assign new_n19561 = new_n19560 ^ new_n19557;
  assign new_n19562 = new_n19541 ^ new_n19529;
  assign new_n19563 = ~new_n19542 & ~new_n19562;
  assign new_n19564 = new_n19563 ^ new_n19537;
  assign new_n19565 = ~n124 & new_n9495;
  assign new_n19566 = new_n19565 ^ new_n19527;
  assign new_n19567 = n123 & new_n19566;
  assign new_n19568 = new_n9495 ^ n123;
  assign new_n19569 = new_n11789 ^ n122;
  assign new_n19570 = new_n19569 ^ new_n19566;
  assign new_n19571 = new_n19570 ^ n122;
  assign new_n19572 = new_n19568 & new_n19571;
  assign new_n19573 = new_n19572 ^ new_n19527;
  assign new_n19574 = new_n19573 ^ new_n19567;
  assign new_n19575 = new_n19574 ^ new_n19564;
  assign new_n19576 = n126 & new_n9195;
  assign new_n19577 = new_n9185 & new_n10304;
  assign new_n19578 = new_n19577 ^ new_n19576;
  assign new_n19579 = n127 & new_n9184;
  assign new_n19580 = n125 & new_n9189;
  assign new_n19581 = new_n19580 ^ new_n19579;
  assign new_n19582 = new_n19581 ^ new_n19578;
  assign new_n19583 = new_n19582 ^ n63;
  assign new_n19584 = new_n19583 ^ new_n19575;
  assign new_n19585 = new_n19584 ^ new_n19561;
  assign new_n19586 = new_n19551 ^ new_n19520;
  assign new_n19587 = ~new_n19552 & ~new_n19586;
  assign new_n19588 = new_n19587 ^ new_n19520;
  assign new_n19589 = new_n19588 ^ new_n19585;
  assign new_n19590 = ~new_n19583 & new_n19575;
  assign new_n19591 = new_n19590 ^ new_n19584;
  assign new_n19592 = ~new_n19557 & ~new_n19560;
  assign new_n19593 = new_n19592 ^ new_n19561;
  assign new_n19594 = ~new_n19593 & new_n19591;
  assign new_n19595 = new_n19590 ^ new_n19588;
  assign new_n19596 = new_n19593 ^ new_n19590;
  assign new_n19597 = ~new_n19595 & ~new_n19596;
  assign new_n19598 = new_n19597 ^ new_n19594;
  assign new_n19599 = new_n19590 & new_n19592;
  assign new_n19600 = new_n19591 ^ new_n19588;
  assign new_n19601 = new_n19592 ^ new_n19591;
  assign new_n19602 = new_n19600 & new_n19601;
  assign new_n19603 = new_n19602 ^ new_n19599;
  assign new_n19604 = new_n19603 ^ new_n19598;
  assign new_n19605 = n127 & new_n9195;
  assign new_n19606 = new_n9185 & new_n10581;
  assign new_n19607 = new_n19606 ^ new_n19605;
  assign new_n19608 = n128 & new_n9184;
  assign new_n19609 = n126 & new_n9189;
  assign new_n19610 = new_n19609 ^ new_n19608;
  assign new_n19611 = new_n19610 ^ new_n19607;
  assign new_n19612 = new_n19611 ^ n63;
  assign new_n19613 = n125 ^ n123;
  assign new_n19614 = ~new_n11492 & new_n19613;
  assign new_n19615 = new_n19614 ^ n123;
  assign new_n19616 = new_n19615 ^ n124;
  assign new_n19617 = new_n11789 & new_n19616;
  assign new_n19618 = new_n19617 ^ n60;
  assign new_n19619 = new_n19618 ^ new_n19612;
  assign new_n19620 = ~new_n19564 & ~new_n19574;
  assign new_n19621 = new_n19620 ^ new_n19572;
  assign new_n19622 = new_n19621 ^ new_n19619;
  assign new_n19623 = new_n19622 ^ new_n19604;
  assign new_n19624 = ~new_n19622 & new_n19593;
  assign new_n19625 = ~new_n19590 & ~new_n19624;
  assign new_n19626 = ~new_n19592 & new_n19591;
  assign new_n19627 = ~new_n19592 & new_n19622;
  assign new_n19628 = ~new_n19626 & ~new_n19627;
  assign new_n19629 = ~new_n19625 & new_n19628;
  assign new_n19630 = ~new_n19588 & ~new_n19629;
  assign new_n19631 = ~new_n19624 & new_n19591;
  assign new_n19632 = new_n19590 & new_n19593;
  assign new_n19633 = ~new_n19632 & new_n19627;
  assign new_n19634 = ~new_n19631 & ~new_n19633;
  assign new_n19635 = ~new_n19630 & new_n19634;
  assign new_n19636 = n127 & new_n9189;
  assign new_n19637 = new_n9185 & new_n10010;
  assign new_n19638 = new_n19637 ^ new_n19636;
  assign new_n19639 = n128 & new_n9195;
  assign new_n19640 = new_n19639 ^ new_n19638;
  assign new_n19641 = new_n19640 ^ n63;
  assign new_n19642 = n124 ^ n60;
  assign new_n19643 = ~new_n19642 & new_n19616;
  assign new_n19644 = new_n19643 ^ n124;
  assign new_n19645 = new_n11789 & new_n19644;
  assign new_n19646 = new_n19645 ^ new_n19641;
  assign new_n19647 = new_n9423 & new_n11492;
  assign new_n19648 = n64 & n126;
  assign new_n19649 = n126 & new_n11491;
  assign new_n19650 = new_n19649 ^ new_n19648;
  assign new_n19651 = new_n19650 ^ new_n19647;
  assign new_n19652 = new_n19651 ^ new_n19646;
  assign new_n19653 = new_n19621 ^ new_n19612;
  assign new_n19654 = ~new_n19653 & new_n19619;
  assign new_n19655 = new_n19654 ^ new_n19621;
  assign new_n19656 = new_n19655 ^ new_n19652;
  assign new_n19657 = new_n19656 ^ new_n19635;
  assign new_n19658 = n128 & new_n9189;
  assign new_n19659 = new_n9185 & new_n11133;
  assign new_n19660 = new_n19659 ^ new_n19658;
  assign new_n19661 = new_n19647 ^ n64;
  assign new_n19662 = ~new_n9718 & new_n9495;
  assign new_n19663 = new_n19662 ^ new_n19661;
  assign new_n19664 = new_n19663 ^ new_n19660;
  assign new_n19665 = new_n19651 ^ new_n19645;
  assign new_n19666 = new_n19646 & new_n19665;
  assign new_n19667 = new_n19666 ^ new_n19641;
  assign new_n19668 = new_n19667 ^ new_n19664;
  assign new_n19669 = new_n19652 ^ new_n19635;
  assign new_n19670 = ~new_n19669 & new_n19656;
  assign new_n19671 = new_n19670 ^ new_n19655;
  assign new_n19672 = new_n19671 ^ new_n19668;
  assign new_n19673 = new_n19660 ^ n126;
  assign new_n19674 = ~new_n9423 & ~new_n19673;
  assign new_n19675 = new_n19674 ^ n126;
  assign new_n19676 = new_n19660 ^ n127;
  assign new_n19677 = new_n9718 & new_n19676;
  assign new_n19678 = new_n19677 ^ new_n19673;
  assign new_n19679 = new_n19678 ^ n127;
  assign new_n19680 = new_n19679 ^ new_n19675;
  assign new_n19681 = ~n64 & ~new_n19680;
  assign new_n19682 = new_n19681 ^ new_n19675;
  assign new_n19683 = n64 & new_n19677;
  assign new_n19684 = new_n19683 ^ new_n19660;
  assign new_n19685 = new_n19684 ^ new_n19682;
  assign new_n19686 = n63 & new_n19685;
  assign new_n19687 = new_n19686 ^ new_n19684;
  assign new_n19688 = n128 ^ n126;
  assign new_n19689 = new_n19688 ^ n63;
  assign new_n19690 = n127 ^ n125;
  assign new_n19691 = new_n19690 ^ new_n19688;
  assign new_n19692 = new_n19691 ^ new_n19688;
  assign new_n19693 = n64 & new_n19692;
  assign new_n19694 = new_n19693 ^ new_n19688;
  assign new_n19695 = ~new_n9495 & new_n19694;
  assign new_n19696 = new_n19695 ^ new_n19689;
  assign new_n19697 = new_n19696 ^ new_n19687;
  assign new_n19698 = new_n19671 ^ new_n19667;
  assign new_n19699 = ~new_n19698 & new_n19668;
  assign new_n19700 = new_n19699 ^ new_n19671;
  assign new_n19701 = new_n19700 ^ new_n19697;
  assign new_n19702 = ~n126 & ~n128;
  assign new_n19703 = ~new_n19702 & n64;
  assign new_n19704 = new_n19703 ^ new_n19649;
  assign new_n19705 = n125 & n127;
  assign new_n19706 = new_n11492 & new_n19705;
  assign new_n19707 = ~n128 & n126;
  assign new_n19708 = n63 & new_n19707;
  assign new_n19709 = new_n19708 ^ new_n19706;
  assign new_n19710 = new_n19709 ^ new_n19704;
  assign new_n19711 = new_n19700 ^ new_n19687;
  assign new_n19712 = ~new_n19711 & new_n19697;
  assign new_n19713 = new_n19712 ^ new_n19700;
  assign new_n19714 = new_n19713 ^ new_n19710;
  assign po0 = new_n129;
  assign po1 = new_n132;
  assign po2 = new_n148;
  assign po3 = new_n179;
  assign po4 = new_n205;
  assign po5 = new_n257;
  assign po6 = new_n289;
  assign po7 = ~new_n334;
  assign po8 = ~new_n383;
  assign po9 = new_n436;
  assign po10 = new_n493;
  assign po11 = new_n565;
  assign po12 = new_n626;
  assign po13 = ~new_n690;
  assign po14 = new_n767;
  assign po15 = new_n842;
  assign po16 = new_n922;
  assign po17 = new_n1015;
  assign po18 = new_n1099;
  assign po19 = new_n1190;
  assign po20 = new_n1296;
  assign po21 = new_n1393;
  assign po22 = new_n1498;
  assign po23 = new_n1614;
  assign po24 = new_n1724;
  assign po25 = new_n1841;
  assign po26 = new_n1970;
  assign po27 = ~new_n2093;
  assign po28 = new_n2225;
  assign po29 = new_n2373;
  assign po30 = new_n2514;
  assign po31 = new_n2660;
  assign po32 = new_n2815;
  assign po33 = new_n2968;
  assign po34 = new_n3135;
  assign po35 = new_n3303;
  assign po36 = new_n3464;
  assign po37 = new_n3638;
  assign po38 = new_n3827;
  assign po39 = new_n4005;
  assign po40 = new_n4190;
  assign po41 = new_n4398;
  assign po42 = ~new_n4587;
  assign po43 = new_n4784;
  assign po44 = new_n4993;
  assign po45 = new_n5198;
  assign po46 = new_n5411;
  assign po47 = ~new_n5637;
  assign po48 = ~new_n5856;
  assign po49 = new_n6079;
  assign po50 = new_n6315;
  assign po51 = new_n6549;
  assign po52 = ~new_n6797;
  assign po53 = new_n7046;
  assign po54 = new_n7286;
  assign po55 = new_n7532;
  assign po56 = new_n7792;
  assign po57 = ~new_n8057;
  assign po58 = new_n8318;
  assign po59 = new_n8601;
  assign po60 = new_n8872;
  assign po61 = ~new_n9154;
  assign po62 = ~new_n9455;
  assign po63 = ~new_n9747;
  assign po64 = new_n10039;
  assign po65 = ~new_n10325;
  assign po66 = new_n10597;
  assign po67 = new_n10872;
  assign po68 = ~new_n11150;
  assign po69 = new_n11430;
  assign po70 = new_n11697;
  assign po71 = ~new_n11975;
  assign po72 = ~new_n12230;
  assign po73 = ~new_n12483;
  assign po74 = ~new_n12745;
  assign po75 = ~new_n12981;
  assign po76 = ~new_n13212;
  assign po77 = new_n13443;
  assign po78 = new_n13683;
  assign po79 = ~new_n13915;
  assign po80 = ~new_n14147;
  assign po81 = ~new_n14383;
  assign po82 = ~new_n14593;
  assign po83 = ~new_n14807;
  assign po84 = new_n15013;
  assign po85 = new_n15214;
  assign po86 = ~new_n15403;
  assign po87 = new_n15588;
  assign po88 = new_n15768;
  assign po89 = new_n15956;
  assign po90 = ~new_n16134;
  assign po91 = new_n16310;
  assign po92 = ~new_n16477;
  assign po93 = ~new_n16639;
  assign po94 = ~new_n16793;
  assign po95 = new_n16979;
  assign po96 = ~new_n17122;
  assign po97 = new_n17268;
  assign po98 = new_n17410;
  assign po99 = ~new_n17550;
  assign po100 = new_n17677;
  assign po101 = ~new_n17808;
  assign po102 = ~new_n17929;
  assign po103 = ~new_n18051;
  assign po104 = new_n18166;
  assign po105 = new_n18283;
  assign po106 = new_n18387;
  assign po107 = ~new_n18485;
  assign po108 = new_n18610;
  assign po109 = new_n18708;
  assign po110 = ~new_n18811;
  assign po111 = ~new_n18898;
  assign po112 = new_n18980;
  assign po113 = new_n19063;
  assign po114 = ~new_n19152;
  assign po115 = ~new_n19223;
  assign po116 = ~new_n19288;
  assign po117 = new_n19340;
  assign po118 = new_n19402;
  assign po119 = ~new_n19456;
  assign po120 = ~new_n19509;
  assign po121 = ~new_n19553;
  assign po122 = new_n19589;
  assign po123 = ~new_n19623;
  assign po124 = ~new_n19657;
  assign po125 = new_n19672;
  assign po126 = new_n19701;
  assign po127 = new_n19714;
endmodule


