module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 ;
  assign n82 = x4 & x7 ;
  assign n83 = n82 ^ x7 ;
  assign n101 = x1 & x2 ;
  assign n102 = n101 ^ x1 ;
  assign n103 = n83 & n102 ;
  assign n104 = n103 ^ n102 ;
  assign n73 = x3 & x4 ;
  assign n105 = x4 & x8 ;
  assign n106 = n73 & n105 ;
  assign n107 = n106 ^ n73 ;
  assign n108 = n107 ^ n105 ;
  assign n109 = n104 & ~n108 ;
  assign n110 = x7 & x8 ;
  assign n111 = n110 ^ x7 ;
  assign n112 = n111 ^ x8 ;
  assign n113 = n101 ^ x2 ;
  assign n114 = ~n112 & n113 ;
  assign n115 = x9 & n114 ;
  assign n116 = n115 ^ x9 ;
  assign n117 = n116 ^ n114 ;
  assign n118 = n109 & ~n117 ;
  assign n119 = n118 ^ n117 ;
  assign n91 = x5 & x6 ;
  assign n92 = n91 ^ x6 ;
  assign n93 = x9 & ~n92 ;
  assign n120 = n91 ^ x5 ;
  assign n125 = n93 & n120 ;
  assign n126 = n119 & n125 ;
  assign n12 = ~x6 & ~x7 ;
  assign n60 = x1 & x4 ;
  assign n56 = x8 ^ x1 ;
  assign n57 = x4 & n56 ;
  assign n58 = n57 ^ x8 ;
  assign n61 = n60 ^ n58 ;
  assign n62 = n61 ^ n58 ;
  assign n59 = n58 ^ x0 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n59 ^ n58 ;
  assign n65 = n63 & ~n64 ;
  assign n66 = n65 ^ n59 ;
  assign n67 = n12 & n66 ;
  assign n51 = x4 & ~x5 ;
  assign n52 = x8 & n51 ;
  assign n53 = n52 ^ x5 ;
  assign n77 = x2 & x7 ;
  assign n78 = n77 ^ x2 ;
  assign n79 = n78 ^ x7 ;
  assign n80 = x1 & x5 ;
  assign n81 = ~n79 & n80 ;
  assign n84 = n83 ^ n81 ;
  assign n85 = x3 & x8 ;
  assign n86 = n85 ^ x3 ;
  assign n87 = n84 & n86 ;
  assign n74 = n73 ^ x4 ;
  assign n75 = x7 & ~x8 ;
  assign n76 = n74 & n75 ;
  assign n88 = n87 ^ n76 ;
  assign n96 = ~n53 & n88 ;
  assign n97 = n96 ^ n53 ;
  assign n98 = n67 & ~n97 ;
  assign n99 = n98 ^ n97 ;
  assign n47 = x4 & x5 ;
  assign n48 = n47 ^ x5 ;
  assign n49 = x8 & n48 ;
  assign n50 = x5 & ~n49 ;
  assign n95 = n50 & ~n88 ;
  assign n100 = n99 ^ n95 ;
  assign n121 = ~x9 & n120 ;
  assign n122 = ~n119 & n121 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = ~n100 & n123 ;
  assign n127 = n126 ^ n124 ;
  assign n54 = n53 ^ n50 ;
  assign n68 = n67 ^ n54 ;
  assign n55 = n54 ^ n53 ;
  assign n69 = n68 ^ n55 ;
  assign n70 = n55 ^ n54 ;
  assign n71 = ~n69 & ~n70 ;
  assign n72 = n71 ^ n55 ;
  assign n89 = ~x9 & ~n88 ;
  assign n90 = n72 & n89 ;
  assign n94 = n93 ^ n90 ;
  assign n128 = n127 ^ n94 ;
  assign n133 = x10 & n128 ;
  assign n134 = n133 ^ n128 ;
  assign n14 = x10 ^ x8 ;
  assign n15 = n14 ^ x10 ;
  assign n20 = n15 ^ x10 ;
  assign n16 = x10 ^ x9 ;
  assign n17 = n16 ^ x10 ;
  assign n18 = n17 ^ n15 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = x3 ^ x2 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = x10 ^ x7 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n23 & ~n25 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n21 & ~n28 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n22 ;
  assign n19 = n18 ^ n15 ;
  assign n32 = n31 ^ n19 ;
  assign n33 = n20 ^ n15 ;
  assign n35 = n22 ^ n18 ;
  assign n34 = n24 ^ n20 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n33 & n36 ;
  assign n38 = n37 ^ n29 ;
  assign n39 = n38 ^ n26 ;
  assign n40 = ~n32 & n39 ;
  assign n41 = n40 ^ n24 ;
  assign n42 = n41 ^ x10 ;
  assign n43 = n42 ^ n24 ;
  assign n129 = x6 & ~x10 ;
  assign n130 = ~n43 & n129 ;
  assign n131 = n130 ^ n129 ;
  assign n132 = n128 & n131 ;
  assign n135 = n134 ^ n132 ;
  assign n44 = x6 & x10 ;
  assign n45 = ~n43 & n44 ;
  assign n13 = x10 & n12 ;
  assign n46 = n45 ^ n13 ;
  assign n136 = n135 ^ n46 ;
  assign n185 = x4 & x9 ;
  assign n186 = n185 ^ x4 ;
  assign n187 = n186 ^ x9 ;
  assign n188 = ~n79 & ~n187 ;
  assign n189 = n188 ^ n79 ;
  assign n190 = n189 ^ n187 ;
  assign n140 = x8 & x9 ;
  assign n141 = n140 ^ x8 ;
  assign n191 = x1 & n141 ;
  assign n192 = n191 ^ x1 ;
  assign n193 = n192 ^ n141 ;
  assign n194 = ~n190 & ~n193 ;
  assign n195 = n194 ^ n193 ;
  assign n196 = n195 ^ n141 ;
  assign n197 = x0 & x2 ;
  assign n198 = n197 ^ x2 ;
  assign n199 = n82 ^ x4 ;
  assign n200 = n198 & n199 ;
  assign n201 = n200 ^ n199 ;
  assign n208 = x0 & x6 ;
  assign n209 = n208 ^ x0 ;
  assign n210 = n101 & n209 ;
  assign n211 = n210 ^ n209 ;
  assign n212 = n201 & n211 ;
  assign n213 = ~n196 & n212 ;
  assign n214 = n213 ^ n212 ;
  assign n202 = x6 & n201 ;
  assign n203 = n202 ^ x6 ;
  assign n204 = n203 ^ n201 ;
  assign n205 = ~n196 & ~n204 ;
  assign n206 = n205 ^ n204 ;
  assign n207 = n206 ^ x6 ;
  assign n215 = n214 ^ n207 ;
  assign n168 = n105 ^ x8 ;
  assign n169 = n168 ^ x7 ;
  assign n170 = x9 & n169 ;
  assign n171 = n170 ^ x9 ;
  assign n172 = n171 ^ n168 ;
  assign n216 = n172 ^ x6 ;
  assign n217 = ~x5 & ~x10 ;
  assign n218 = n217 ^ x6 ;
  assign n219 = ~n217 & n218 ;
  assign n220 = n219 ^ n217 ;
  assign n221 = n220 ^ n172 ;
  assign n222 = ~n216 & ~n221 ;
  assign n223 = n222 ^ n219 ;
  assign n224 = n223 ^ n172 ;
  assign n142 = n141 ^ x9 ;
  assign n225 = x7 & ~n142 ;
  assign n226 = x7 & x9 ;
  assign n227 = n226 ^ x9 ;
  assign n228 = ~n73 & ~n227 ;
  assign n229 = n225 & n228 ;
  assign n230 = n229 ^ n227 ;
  assign n231 = n230 ^ n224 ;
  assign n232 = n224 & n231 ;
  assign n233 = n232 ^ n230 ;
  assign n234 = n233 ^ n215 ;
  assign n235 = n215 & n234 ;
  assign n236 = n235 ^ n232 ;
  assign n237 = n236 ^ n230 ;
  assign n173 = x6 & ~n172 ;
  assign n174 = n173 ^ x6 ;
  assign n175 = n174 ^ n172 ;
  assign n150 = x7 ^ x4 ;
  assign n151 = x9 & n150 ;
  assign n152 = n151 ^ n150 ;
  assign n153 = n152 ^ x7 ;
  assign n163 = ~x3 & x6 ;
  assign n164 = n142 & n163 ;
  assign n165 = n153 & n164 ;
  assign n166 = n165 ^ x3 ;
  assign n146 = ~x4 & ~x6 ;
  assign n137 = x7 & n101 ;
  assign n147 = n137 ^ n101 ;
  assign n148 = n146 & n147 ;
  assign n138 = n137 ^ x7 ;
  assign n139 = n138 ^ n101 ;
  assign n143 = x4 & ~n142 ;
  assign n144 = ~n139 & n143 ;
  assign n145 = n144 ^ n143 ;
  assign n149 = n148 ^ n145 ;
  assign n160 = x3 & n149 ;
  assign n161 = n160 ^ x3 ;
  assign n154 = x3 & x6 ;
  assign n155 = ~n142 & n154 ;
  assign n156 = n155 ^ n154 ;
  assign n157 = n153 & n156 ;
  assign n158 = n149 & n157 ;
  assign n159 = n158 ^ n157 ;
  assign n162 = n161 ^ n159 ;
  assign n167 = n166 ^ n162 ;
  assign n176 = n175 ^ n167 ;
  assign n177 = x5 & ~x10 ;
  assign n178 = n177 ^ n175 ;
  assign n179 = ~n177 & ~n178 ;
  assign n180 = n179 ^ n175 ;
  assign n181 = n176 & n180 ;
  assign n182 = n181 ^ n179 ;
  assign n183 = n182 ^ n167 ;
  assign n184 = n183 ^ x10 ;
  assign n238 = n237 ^ n184 ;
  assign n252 = ~x4 & x6 ;
  assign n253 = ~x9 & n252 ;
  assign n250 = ~x3 & x5 ;
  assign n251 = ~x6 & n250 ;
  assign n254 = n253 ^ n251 ;
  assign n255 = ~x2 & n254 ;
  assign n247 = x6 & ~x9 ;
  assign n248 = x2 & n73 ;
  assign n249 = n247 & n248 ;
  assign n256 = n255 ^ n249 ;
  assign n257 = ~x4 & n247 ;
  assign n261 = ~x1 & ~x3 ;
  assign n262 = n120 & n261 ;
  assign n263 = ~n257 & n262 ;
  assign n264 = ~n256 & n263 ;
  assign n258 = ~x3 & n257 ;
  assign n259 = ~n256 & n258 ;
  assign n260 = n259 ^ n256 ;
  assign n265 = n264 ^ n260 ;
  assign n239 = x8 & x10 ;
  assign n240 = x6 & x7 ;
  assign n241 = ~x9 & n240 ;
  assign n242 = n239 & n241 ;
  assign n243 = ~x8 & ~n240 ;
  assign n266 = ~x7 & ~x10 ;
  assign n267 = n243 & n266 ;
  assign n268 = ~n242 & n267 ;
  assign n269 = n265 & n268 ;
  assign n244 = x10 & n243 ;
  assign n245 = ~n242 & n244 ;
  assign n246 = n245 ^ n242 ;
  assign n270 = n269 ^ n246 ;
  assign n271 = n238 & n270 ;
  assign n272 = n271 ^ n238 ;
  assign n318 = x7 ^ x6 ;
  assign n320 = x7 ^ x3 ;
  assign n319 = n22 ^ x3 ;
  assign n321 = n320 ^ n319 ;
  assign n322 = n320 ^ x3 ;
  assign n323 = n321 & n322 ;
  assign n324 = n323 ^ n321 ;
  assign n325 = n324 ^ n320 ;
  assign n326 = n318 & n325 ;
  assign n327 = n326 ^ n318 ;
  assign n328 = n327 ^ n240 ;
  assign n329 = n47 & n328 ;
  assign n330 = n329 ^ n47 ;
  assign n331 = n330 ^ n328 ;
  assign n332 = n331 ^ n47 ;
  assign n333 = n332 ^ n327 ;
  assign n273 = n240 ^ x6 ;
  assign n274 = n47 & n273 ;
  assign n275 = n274 ^ n273 ;
  assign n276 = n275 ^ x6 ;
  assign n277 = n276 ^ x7 ;
  assign n334 = n277 ^ x8 ;
  assign n335 = x9 & x10 ;
  assign n336 = n335 ^ x9 ;
  assign n337 = n336 ^ x10 ;
  assign n338 = n337 ^ x8 ;
  assign n339 = ~n337 & ~n338 ;
  assign n340 = n339 ^ n337 ;
  assign n341 = n340 ^ n338 ;
  assign n342 = n341 ^ n337 ;
  assign n343 = n342 ^ n277 ;
  assign n344 = n334 & n343 ;
  assign n345 = n344 ^ n334 ;
  assign n346 = n345 ^ n341 ;
  assign n347 = n346 ^ n277 ;
  assign n348 = n333 & ~n347 ;
  assign n349 = n348 ^ n333 ;
  assign n350 = n349 ^ n347 ;
  assign n372 = x8 & n350 ;
  assign n283 = x0 & x1 ;
  assign n284 = n73 & n283 ;
  assign n285 = n284 ^ n73 ;
  assign n286 = n285 ^ n146 ;
  assign n295 = x2 & ~x5 ;
  assign n296 = n286 & n295 ;
  assign n314 = x7 & n296 ;
  assign n287 = x5 & n286 ;
  assign n288 = n287 ^ n286 ;
  assign n290 = n74 & n209 ;
  assign n289 = x3 & n48 ;
  assign n291 = n290 ^ n289 ;
  assign n312 = n137 & n291 ;
  assign n313 = ~n288 & n312 ;
  assign n315 = n314 ^ n313 ;
  assign n292 = n101 & n291 ;
  assign n293 = n288 & n292 ;
  assign n294 = n293 ^ n292 ;
  assign n297 = n296 ^ n294 ;
  assign n316 = n315 ^ n297 ;
  assign n298 = x6 ^ x5 ;
  assign n300 = n298 ^ x2 ;
  assign n299 = n298 ^ x6 ;
  assign n301 = n300 ^ n299 ;
  assign n302 = n299 ^ n298 ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = n303 ^ n299 ;
  assign n305 = x3 & n304 ;
  assign n306 = n305 ^ n298 ;
  assign n307 = n306 ^ x6 ;
  assign n308 = n199 & ~n307 ;
  assign n309 = n308 ^ n199 ;
  assign n310 = n297 & n309 ;
  assign n311 = n310 ^ n309 ;
  assign n317 = n316 ^ n311 ;
  assign n363 = n73 & n91 ;
  assign n364 = n363 ^ n91 ;
  assign n365 = x8 & n364 ;
  assign n366 = n365 ^ x8 ;
  assign n367 = n366 ^ n364 ;
  assign n353 = x6 ^ x2 ;
  assign n351 = x2 ^ x1 ;
  assign n352 = n351 ^ x2 ;
  assign n354 = n353 ^ n352 ;
  assign n355 = n353 ^ x2 ;
  assign n356 = n354 & n355 ;
  assign n357 = n356 ^ n354 ;
  assign n358 = n357 ^ n353 ;
  assign n359 = n298 & n358 ;
  assign n360 = n359 ^ n298 ;
  assign n361 = ~x8 & n73 ;
  assign n362 = n360 & n361 ;
  assign n368 = n367 ^ n362 ;
  assign n369 = n350 & ~n368 ;
  assign n370 = n317 & n369 ;
  assign n371 = n370 ^ n369 ;
  assign n373 = n372 ^ n371 ;
  assign n278 = x8 & ~n277 ;
  assign n279 = n278 ^ x8 ;
  assign n280 = x9 & ~x10 ;
  assign n281 = ~n279 & n280 ;
  assign n282 = n281 ^ x10 ;
  assign n374 = n373 ^ n282 ;
  assign n375 = x5 & ~x8 ;
  assign n376 = x9 & n375 ;
  assign n377 = ~n239 & ~n376 ;
  assign n378 = n240 & ~n377 ;
  assign n379 = x5 & x7 ;
  assign n380 = x8 & ~n379 ;
  assign n381 = ~x10 & ~n380 ;
  assign n382 = x9 & ~n381 ;
  assign n383 = ~n378 & ~n382 ;
  assign n384 = n374 & n383 ;
  assign n385 = x7 & n91 ;
  assign n386 = ~x2 & n105 ;
  assign n387 = n385 & n386 ;
  assign n388 = ~x5 & ~x6 ;
  assign n389 = ~x4 & ~x7 ;
  assign n390 = ~x8 & n389 ;
  assign n391 = n388 & n390 ;
  assign n392 = ~n387 & ~n391 ;
  assign n393 = ~x3 & ~n337 ;
  assign n394 = ~n392 & n393 ;
  assign n399 = x3 & ~x7 ;
  assign n400 = n101 & n399 ;
  assign n395 = ~x5 & ~x7 ;
  assign n401 = ~n91 & ~n395 ;
  assign n402 = n400 & n401 ;
  assign n396 = x3 & n91 ;
  assign n397 = ~n395 & n396 ;
  assign n398 = n397 ^ n395 ;
  assign n403 = n402 ^ n398 ;
  assign n405 = ~x4 & ~n273 ;
  assign n406 = n403 & n405 ;
  assign n404 = ~n273 & ~n403 ;
  assign n407 = n406 ^ n404 ;
  assign n409 = n283 & n388 ;
  assign n410 = ~n274 & ~n409 ;
  assign n411 = x2 & x3 ;
  assign n412 = ~x8 & n411 ;
  assign n413 = ~n410 & n412 ;
  assign n414 = ~n407 & n413 ;
  assign n408 = ~x8 & n407 ;
  assign n415 = n414 ^ n408 ;
  assign n416 = n91 & n110 ;
  assign n417 = x9 & ~n416 ;
  assign n425 = ~x10 & ~n417 ;
  assign n426 = ~n415 & n425 ;
  assign n418 = n47 & n241 ;
  assign n419 = x2 & ~x3 ;
  assign n420 = ~n85 & ~n419 ;
  assign n421 = ~x10 & ~n420 ;
  assign n422 = n418 & n421 ;
  assign n423 = ~n417 & n422 ;
  assign n424 = ~n415 & n423 ;
  assign n427 = n426 ^ n424 ;
  assign n428 = n427 ^ x10 ;
  assign n430 = n86 & n283 ;
  assign n431 = n395 & n430 ;
  assign n432 = x2 & ~n416 ;
  assign n433 = ~n431 & n432 ;
  assign n434 = n433 ^ x2 ;
  assign n429 = n85 & n385 ;
  assign n435 = n434 ^ n429 ;
  assign n436 = n429 ^ x4 ;
  assign n437 = ~x4 & n436 ;
  assign n438 = n437 ^ x4 ;
  assign n439 = n438 ^ n434 ;
  assign n440 = n435 & n439 ;
  assign n441 = n440 ^ n437 ;
  assign n442 = n441 ^ n434 ;
  assign n443 = n91 & n248 ;
  assign n444 = ~n112 & ~n388 ;
  assign n445 = ~n443 & n444 ;
  assign n446 = ~n337 & ~n445 ;
  assign n447 = n442 & n446 ;
  assign n448 = n447 ^ n446 ;
  assign n449 = ~n112 & ~n337 ;
  assign n450 = ~n443 & n449 ;
  assign y0 = ~n136 ;
  assign y1 = n272 ;
  assign y2 = ~n384 ;
  assign y3 = ~n394 ;
  assign y4 = n428 ;
  assign y5 = ~n448 ;
  assign y6 = ~n450 ;
endmodule
