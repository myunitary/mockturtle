module point_and_ary_16( a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, b11, b12, b13, b14, b15, d0 );
  input a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15;
  input b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, b11, b12, b13, b14, b15;
  output d0;
  wire e0, e1, e2, e3, e4, e5, e6, e7, e8, e9, e10, e11, e12, e13, e14, e15,c0, c1, c2, c3, c4, c5, c6, c7, c8, c9, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c20, c21, c22, c23, c24, c25, c26, c27;
  assign e0 = a0 ^ b0;
  assign e1 = a1 ^ b1;
  assign e2 = a2 ^ b2;
  assign e3 = a3 ^ b3;
  assign e4 = a4 ^ b4;
  assign e5 = a5 ^ b5;
  assign e6 = a6 ^ b6;
  assign e7 = a7 ^ b7;
  assign e8 = a8 ^ b8;
  assign e9 = a9 ^ b9;
  assign e10 = a10 ^ b10;
  assign e11 = a11 ^ b11;
  assign e12 = a12 ^ b12;
  assign e13 = a13 ^ b13;
  assign e14 = a14 ^ b14;
  assign e15 = a15 ^ b15;
  assign c0 = e0 & e1;
  assign c1 = e2 & e3;
  assign c2 = e4 & e5;
  assign c3 = e6 & e7;
  assign c4 = e8 & e9;
  assign c5 = e10 & e11;
  assign c6 = e12 & e13;
  assign c7 = e14 & e15;
  assign c8 = c0 & c1;
  assign c9 = c2 & c3;
  assign c10 = c4 & c5;
  assign c11 = c6 & c7;
  assign c12 = c8 & c9;
  assign c13 = c10 & c11;
  assign d0 = c12 & c13;
endmodule
