module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 ;
  assign n50 = x8 ^ x0 ;
  assign n54 = x9 ^ x1 ;
  assign n55 = n50 & n54 ;
  assign n56 = n55 ^ n50 ;
  assign n57 = n56 ^ n54 ;
  assign n59 = x10 ^ x2 ;
  assign n67 = x11 ^ x3 ;
  assign n68 = n59 & n67 ;
  assign n69 = n68 ^ n59 ;
  assign n70 = n69 ^ n67 ;
  assign n71 = ~n57 & ~n70 ;
  assign n73 = x12 ^ x4 ;
  assign n77 = x13 ^ x5 ;
  assign n78 = n73 & n77 ;
  assign n79 = n78 ^ n73 ;
  assign n80 = n79 ^ n77 ;
  assign n82 = x14 ^ x6 ;
  assign n92 = x15 ^ x7 ;
  assign n93 = n82 & n92 ;
  assign n94 = n93 ^ n82 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = ~n80 & ~n95 ;
  assign n97 = n71 & n96 ;
  assign n83 = x7 & x15 ;
  assign n84 = n83 ^ x7 ;
  assign n85 = n82 & n84 ;
  assign n86 = n85 ^ n84 ;
  assign n81 = x6 & ~x14 ;
  assign n87 = n86 ^ n81 ;
  assign n88 = ~n80 & n87 ;
  assign n74 = x5 & ~x13 ;
  assign n75 = ~n73 & n74 ;
  assign n72 = x4 & ~x12 ;
  assign n76 = n75 ^ n72 ;
  assign n89 = n88 ^ n76 ;
  assign n90 = n71 & n89 ;
  assign n60 = x3 & x11 ;
  assign n61 = n60 ^ x3 ;
  assign n62 = n59 & n61 ;
  assign n63 = n62 ^ n61 ;
  assign n58 = x2 & ~x10 ;
  assign n64 = n63 ^ n58 ;
  assign n65 = ~n57 & n64 ;
  assign n51 = x1 & ~x9 ;
  assign n52 = ~n50 & n51 ;
  assign n49 = x0 & ~x8 ;
  assign n53 = n52 ^ n49 ;
  assign n66 = n65 ^ n53 ;
  assign n91 = n90 ^ n66 ;
  assign n98 = n97 ^ n91 ;
  assign n103 = x0 & n98 ;
  assign n100 = x8 & n98 ;
  assign n102 = n100 ^ x8 ;
  assign n104 = n103 ^ n102 ;
  assign n106 = n104 ^ x16 ;
  assign n109 = x1 & n98 ;
  assign n107 = x9 & n98 ;
  assign n108 = n107 ^ x9 ;
  assign n110 = n109 ^ n108 ;
  assign n114 = n110 ^ x17 ;
  assign n115 = n106 & n114 ;
  assign n116 = n115 ^ n106 ;
  assign n117 = n116 ^ n114 ;
  assign n120 = x2 & n98 ;
  assign n118 = x10 & n98 ;
  assign n119 = n118 ^ x10 ;
  assign n121 = n120 ^ n119 ;
  assign n123 = n121 ^ x18 ;
  assign n126 = x3 & n98 ;
  assign n124 = x11 & n98 ;
  assign n125 = n124 ^ x11 ;
  assign n127 = n126 ^ n125 ;
  assign n135 = n127 ^ x19 ;
  assign n136 = n123 & n135 ;
  assign n137 = n136 ^ n123 ;
  assign n138 = n137 ^ n135 ;
  assign n139 = ~n117 & ~n138 ;
  assign n142 = x4 & n98 ;
  assign n140 = x12 & n98 ;
  assign n141 = n140 ^ x12 ;
  assign n143 = n142 ^ n141 ;
  assign n145 = n143 ^ x20 ;
  assign n148 = x5 & n98 ;
  assign n146 = x13 & n98 ;
  assign n147 = n146 ^ x13 ;
  assign n149 = n148 ^ n147 ;
  assign n155 = n149 ^ x21 ;
  assign n156 = n145 & n155 ;
  assign n157 = n156 ^ n145 ;
  assign n158 = n157 ^ n155 ;
  assign n161 = x6 & n98 ;
  assign n159 = x14 & n98 ;
  assign n160 = n159 ^ x14 ;
  assign n162 = n161 ^ n160 ;
  assign n165 = n162 ^ x22 ;
  assign n179 = x7 & n66 ;
  assign n180 = n179 ^ x7 ;
  assign n177 = x7 & n97 ;
  assign n178 = n177 ^ x7 ;
  assign n181 = n180 ^ n178 ;
  assign n175 = x7 & n71 ;
  assign n176 = n89 & n175 ;
  assign n182 = n181 ^ n176 ;
  assign n170 = x15 & n66 ;
  assign n171 = n170 ^ x15 ;
  assign n168 = x15 & n97 ;
  assign n169 = n168 ^ x15 ;
  assign n172 = n171 ^ n169 ;
  assign n166 = x15 & n71 ;
  assign n167 = n89 & n166 ;
  assign n173 = n172 ^ n167 ;
  assign n174 = n173 ^ x15 ;
  assign n183 = n182 ^ n174 ;
  assign n193 = n183 ^ x23 ;
  assign n194 = n165 & n193 ;
  assign n195 = n194 ^ n165 ;
  assign n196 = n195 ^ n193 ;
  assign n197 = ~n158 & ~n196 ;
  assign n198 = n139 & n197 ;
  assign n184 = x23 & n183 ;
  assign n185 = n184 ^ n183 ;
  assign n186 = n165 & n185 ;
  assign n187 = n186 ^ n185 ;
  assign n163 = x22 & n162 ;
  assign n164 = n163 ^ n162 ;
  assign n188 = n187 ^ n164 ;
  assign n189 = ~n158 & n188 ;
  assign n150 = x21 & n149 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = n145 & n151 ;
  assign n153 = n152 ^ n151 ;
  assign n144 = ~x20 & n143 ;
  assign n154 = n153 ^ n144 ;
  assign n190 = n189 ^ n154 ;
  assign n191 = n139 & n190 ;
  assign n128 = x19 & n127 ;
  assign n129 = n128 ^ n127 ;
  assign n130 = n123 & n129 ;
  assign n131 = n130 ^ n129 ;
  assign n122 = ~x18 & n121 ;
  assign n132 = n131 ^ n122 ;
  assign n133 = ~n117 & n132 ;
  assign n111 = ~x17 & n110 ;
  assign n112 = ~n106 & n111 ;
  assign n105 = ~x16 & n104 ;
  assign n113 = n112 ^ n105 ;
  assign n134 = n133 ^ n113 ;
  assign n192 = n191 ^ n134 ;
  assign n199 = n198 ^ n192 ;
  assign n202 = x16 & n199 ;
  assign n310 = n202 ^ x16 ;
  assign n200 = n104 & n199 ;
  assign n311 = n310 ^ n200 ;
  assign n313 = n311 ^ x24 ;
  assign n208 = x17 & n199 ;
  assign n314 = n208 ^ x17 ;
  assign n206 = n110 & n199 ;
  assign n315 = n314 ^ n206 ;
  assign n319 = n315 ^ x25 ;
  assign n320 = n313 & n319 ;
  assign n321 = n320 ^ n313 ;
  assign n322 = n321 ^ n319 ;
  assign n223 = x18 & n199 ;
  assign n323 = n223 ^ x18 ;
  assign n221 = n121 & n199 ;
  assign n324 = n323 ^ n221 ;
  assign n326 = n324 ^ x26 ;
  assign n231 = x19 & n199 ;
  assign n327 = n231 ^ x19 ;
  assign n229 = n127 & n199 ;
  assign n328 = n327 ^ n229 ;
  assign n336 = n328 ^ x27 ;
  assign n337 = n326 & n336 ;
  assign n338 = n337 ^ n326 ;
  assign n339 = n338 ^ n336 ;
  assign n340 = ~n322 & ~n339 ;
  assign n249 = x20 & n199 ;
  assign n341 = n249 ^ x20 ;
  assign n247 = n143 & n199 ;
  assign n342 = n341 ^ n247 ;
  assign n344 = n342 ^ x28 ;
  assign n257 = x21 & n199 ;
  assign n345 = n257 ^ x21 ;
  assign n255 = n149 & n199 ;
  assign n346 = n345 ^ n255 ;
  assign n352 = n346 ^ x29 ;
  assign n353 = n344 & n352 ;
  assign n354 = n353 ^ n344 ;
  assign n355 = n354 ^ n352 ;
  assign n272 = x22 & n199 ;
  assign n369 = n272 ^ x22 ;
  assign n270 = n162 & n199 ;
  assign n382 = n369 ^ n270 ;
  assign n383 = n382 ^ x30 ;
  assign n295 = x23 & n199 ;
  assign n364 = n295 ^ x23 ;
  assign n293 = n183 & n199 ;
  assign n365 = n364 ^ n293 ;
  assign n384 = n365 ^ x31 ;
  assign n385 = n383 & n384 ;
  assign n386 = n385 ^ n383 ;
  assign n387 = n386 ^ n384 ;
  assign n388 = ~n355 & ~n387 ;
  assign n389 = n340 & n388 ;
  assign n374 = x22 & ~x30 ;
  assign n375 = ~n199 & n374 ;
  assign n360 = x23 & x31 ;
  assign n361 = n199 & n360 ;
  assign n362 = n361 ^ n360 ;
  assign n358 = x31 & n183 ;
  assign n359 = n199 & n358 ;
  assign n363 = n362 ^ n359 ;
  assign n366 = n365 ^ n363 ;
  assign n370 = n366 & n369 ;
  assign n368 = n270 & n366 ;
  assign n371 = n370 ^ n368 ;
  assign n367 = x30 & n366 ;
  assign n372 = n371 ^ n367 ;
  assign n373 = n372 ^ n366 ;
  assign n376 = n375 ^ n373 ;
  assign n356 = ~x30 & n162 ;
  assign n357 = n199 & n356 ;
  assign n377 = n376 ^ n357 ;
  assign n378 = ~n355 & n377 ;
  assign n347 = x29 & n346 ;
  assign n348 = n347 ^ n346 ;
  assign n349 = n344 & n348 ;
  assign n350 = n349 ^ n348 ;
  assign n343 = ~x28 & n342 ;
  assign n351 = n350 ^ n343 ;
  assign n379 = n378 ^ n351 ;
  assign n380 = n340 & n379 ;
  assign n329 = x27 & n328 ;
  assign n330 = n329 ^ n328 ;
  assign n331 = n326 & n330 ;
  assign n332 = n331 ^ n330 ;
  assign n325 = ~x26 & n324 ;
  assign n333 = n332 ^ n325 ;
  assign n334 = ~n322 & n333 ;
  assign n316 = ~x25 & n315 ;
  assign n317 = ~n313 & n316 ;
  assign n312 = ~x24 & n311 ;
  assign n318 = n317 ^ n312 ;
  assign n335 = n334 ^ n318 ;
  assign n381 = n380 ^ n335 ;
  assign n390 = n389 ^ n381 ;
  assign n577 = n311 & n390 ;
  assign n576 = x24 & ~n390 ;
  assign n578 = n577 ^ n576 ;
  assign n580 = n578 ^ x32 ;
  assign n582 = n315 & n390 ;
  assign n581 = x25 & ~n390 ;
  assign n583 = n582 ^ n581 ;
  assign n587 = n583 ^ x33 ;
  assign n588 = ~n580 & ~n587 ;
  assign n590 = n324 & n390 ;
  assign n589 = x26 & ~n390 ;
  assign n591 = n590 ^ n589 ;
  assign n593 = n591 ^ x34 ;
  assign n595 = n328 & n390 ;
  assign n594 = x27 & ~n390 ;
  assign n596 = n595 ^ n594 ;
  assign n602 = n596 ^ x35 ;
  assign n603 = ~n593 & ~n602 ;
  assign n604 = n588 & n603 ;
  assign n606 = n342 & n390 ;
  assign n605 = x28 & ~n390 ;
  assign n607 = n606 ^ n605 ;
  assign n609 = n607 ^ x36 ;
  assign n611 = n346 & n390 ;
  assign n610 = x29 & ~n390 ;
  assign n612 = n611 ^ n610 ;
  assign n616 = n612 ^ x37 ;
  assign n617 = ~n609 & ~n616 ;
  assign n631 = x30 & ~n390 ;
  assign n629 = n382 & n390 ;
  assign n644 = n631 ^ n629 ;
  assign n645 = n644 ^ x38 ;
  assign n458 = x31 & n390 ;
  assign n625 = n458 ^ x31 ;
  assign n456 = n365 & n390 ;
  assign n626 = n625 ^ n456 ;
  assign n646 = n626 ^ x39 ;
  assign n647 = ~n645 & ~n646 ;
  assign n648 = n617 & n647 ;
  assign n649 = n604 & n648 ;
  assign n636 = x30 & ~x38 ;
  assign n637 = ~n390 & n636 ;
  assign n622 = x31 & x39 ;
  assign n623 = ~n390 & n622 ;
  assign n620 = x39 & n365 ;
  assign n621 = n390 & n620 ;
  assign n624 = n623 ^ n621 ;
  assign n627 = n626 ^ n624 ;
  assign n632 = n627 & n631 ;
  assign n630 = n627 & n629 ;
  assign n633 = n632 ^ n630 ;
  assign n628 = x38 & n627 ;
  assign n634 = n633 ^ n628 ;
  assign n635 = n634 ^ n627 ;
  assign n638 = n637 ^ n635 ;
  assign n618 = ~x38 & n382 ;
  assign n619 = n390 & n618 ;
  assign n639 = n638 ^ n619 ;
  assign n640 = n617 & n639 ;
  assign n613 = ~x37 & n612 ;
  assign n614 = ~n609 & n613 ;
  assign n608 = ~x36 & n607 ;
  assign n615 = n614 ^ n608 ;
  assign n641 = n640 ^ n615 ;
  assign n642 = n604 & n641 ;
  assign n597 = ~x35 & n596 ;
  assign n598 = ~n593 & n597 ;
  assign n592 = ~x34 & n591 ;
  assign n599 = n598 ^ n592 ;
  assign n600 = n588 & n599 ;
  assign n584 = ~x33 & n583 ;
  assign n585 = ~n580 & n584 ;
  assign n579 = ~x32 & n578 ;
  assign n586 = n585 ^ n579 ;
  assign n601 = n600 ^ n586 ;
  assign n643 = n642 ^ n601 ;
  assign n650 = n649 ^ n643 ;
  assign n925 = n578 & n650 ;
  assign n924 = x32 & ~n650 ;
  assign n926 = n925 ^ n924 ;
  assign n928 = n926 ^ x40 ;
  assign n930 = n583 & n650 ;
  assign n929 = x33 & ~n650 ;
  assign n931 = n930 ^ n929 ;
  assign n935 = n931 ^ x41 ;
  assign n936 = ~n928 & ~n935 ;
  assign n938 = n591 & n650 ;
  assign n937 = x34 & ~n650 ;
  assign n939 = n938 ^ n937 ;
  assign n941 = n939 ^ x42 ;
  assign n943 = n596 & n650 ;
  assign n942 = x35 & ~n650 ;
  assign n944 = n943 ^ n942 ;
  assign n950 = n944 ^ x43 ;
  assign n951 = ~n941 & ~n950 ;
  assign n952 = n936 & n951 ;
  assign n954 = n607 & n650 ;
  assign n953 = x36 & ~n650 ;
  assign n955 = n954 ^ n953 ;
  assign n957 = n955 ^ x44 ;
  assign n959 = n612 & n650 ;
  assign n958 = x37 & ~n650 ;
  assign n960 = n959 ^ n958 ;
  assign n964 = n960 ^ x45 ;
  assign n965 = ~n957 & ~n964 ;
  assign n979 = x38 & ~n650 ;
  assign n977 = n644 & n650 ;
  assign n992 = n979 ^ n977 ;
  assign n993 = n992 ^ x46 ;
  assign n718 = x39 & n650 ;
  assign n973 = n718 ^ x39 ;
  assign n716 = n626 & n650 ;
  assign n974 = n973 ^ n716 ;
  assign n994 = n974 ^ x47 ;
  assign n995 = ~n993 & ~n994 ;
  assign n996 = n965 & n995 ;
  assign n997 = n952 & n996 ;
  assign n984 = x38 & ~x46 ;
  assign n985 = ~n650 & n984 ;
  assign n970 = x39 & x47 ;
  assign n971 = ~n650 & n970 ;
  assign n968 = x47 & n626 ;
  assign n969 = n650 & n968 ;
  assign n972 = n971 ^ n969 ;
  assign n975 = n974 ^ n972 ;
  assign n980 = n975 & n979 ;
  assign n978 = n975 & n977 ;
  assign n981 = n980 ^ n978 ;
  assign n976 = x46 & n975 ;
  assign n982 = n981 ^ n976 ;
  assign n983 = n982 ^ n975 ;
  assign n986 = n985 ^ n983 ;
  assign n966 = ~x46 & n644 ;
  assign n967 = n650 & n966 ;
  assign n987 = n986 ^ n967 ;
  assign n988 = n965 & n987 ;
  assign n961 = ~x45 & n960 ;
  assign n962 = ~n957 & n961 ;
  assign n956 = ~x44 & n955 ;
  assign n963 = n962 ^ n956 ;
  assign n989 = n988 ^ n963 ;
  assign n990 = n952 & n989 ;
  assign n945 = ~x43 & n944 ;
  assign n946 = ~n941 & n945 ;
  assign n940 = ~x42 & n939 ;
  assign n947 = n946 ^ n940 ;
  assign n948 = n936 & n947 ;
  assign n932 = ~x41 & n931 ;
  assign n933 = ~n928 & n932 ;
  assign n927 = ~x40 & n926 ;
  assign n934 = n933 ^ n927 ;
  assign n949 = n948 ^ n934 ;
  assign n991 = n990 ^ n949 ;
  assign n998 = n997 ^ n991 ;
  assign n1000 = x40 & n998 ;
  assign n999 = n926 & ~n998 ;
  assign n1001 = n1000 ^ n999 ;
  assign n99 = x0 & ~n98 ;
  assign n101 = n100 ^ n99 ;
  assign n201 = n200 ^ n104 ;
  assign n203 = n202 ^ n201 ;
  assign n205 = n203 ^ n101 ;
  assign n210 = x1 & ~n98 ;
  assign n211 = n210 ^ n107 ;
  assign n207 = n206 ^ n110 ;
  assign n209 = n208 ^ n207 ;
  assign n215 = n211 ^ n209 ;
  assign n216 = n205 & n215 ;
  assign n217 = n216 ^ n205 ;
  assign n218 = n217 ^ n215 ;
  assign n222 = n221 ^ n121 ;
  assign n224 = n223 ^ n222 ;
  assign n219 = x2 & ~n98 ;
  assign n220 = n219 ^ n118 ;
  assign n226 = n224 ^ n220 ;
  assign n230 = n229 ^ n127 ;
  assign n232 = n231 ^ n230 ;
  assign n227 = x3 & ~n98 ;
  assign n228 = n227 ^ n124 ;
  assign n240 = n232 ^ n228 ;
  assign n241 = n226 & n240 ;
  assign n242 = n241 ^ n226 ;
  assign n243 = n242 ^ n240 ;
  assign n244 = ~n218 & ~n243 ;
  assign n248 = n247 ^ n143 ;
  assign n250 = n249 ^ n248 ;
  assign n245 = x4 & ~n98 ;
  assign n246 = n245 ^ n140 ;
  assign n252 = n250 ^ n246 ;
  assign n256 = n255 ^ n149 ;
  assign n258 = n257 ^ n256 ;
  assign n253 = x5 & ~n98 ;
  assign n254 = n253 ^ n146 ;
  assign n264 = n258 ^ n254 ;
  assign n265 = n252 & n264 ;
  assign n266 = n265 ^ n252 ;
  assign n267 = n266 ^ n264 ;
  assign n271 = n270 ^ n162 ;
  assign n273 = n272 ^ n271 ;
  assign n268 = x6 & ~n98 ;
  assign n269 = n268 ^ n159 ;
  assign n276 = n273 ^ n269 ;
  assign n294 = n293 ^ n183 ;
  assign n296 = n295 ^ n294 ;
  assign n277 = x7 & ~n98 ;
  assign n278 = n277 ^ n173 ;
  assign n297 = n296 ^ n278 ;
  assign n298 = n276 & n297 ;
  assign n299 = n298 ^ n276 ;
  assign n300 = n299 ^ n297 ;
  assign n301 = ~n267 & ~n300 ;
  assign n302 = n244 & n301 ;
  assign n282 = x23 & n278 ;
  assign n283 = n199 & n282 ;
  assign n279 = n183 & n278 ;
  assign n280 = n199 & n279 ;
  assign n281 = n280 ^ n279 ;
  assign n284 = n283 ^ n281 ;
  assign n285 = n284 ^ n278 ;
  assign n286 = n276 & n285 ;
  assign n287 = n286 ^ n285 ;
  assign n274 = n269 & n273 ;
  assign n275 = n274 ^ n269 ;
  assign n288 = n287 ^ n275 ;
  assign n289 = ~n267 & n288 ;
  assign n259 = n254 & n258 ;
  assign n260 = n259 ^ n254 ;
  assign n261 = n252 & n260 ;
  assign n262 = n261 ^ n260 ;
  assign n251 = n246 & ~n250 ;
  assign n263 = n262 ^ n251 ;
  assign n290 = n289 ^ n263 ;
  assign n291 = n244 & n290 ;
  assign n233 = n228 & n232 ;
  assign n234 = n233 ^ n228 ;
  assign n235 = n226 & n234 ;
  assign n236 = n235 ^ n234 ;
  assign n225 = n220 & ~n224 ;
  assign n237 = n236 ^ n225 ;
  assign n238 = ~n218 & n237 ;
  assign n212 = ~n209 & n211 ;
  assign n213 = ~n205 & n212 ;
  assign n204 = n101 & ~n203 ;
  assign n214 = n213 ^ n204 ;
  assign n239 = n238 ^ n214 ;
  assign n292 = n291 ^ n239 ;
  assign n303 = n302 ^ n292 ;
  assign n308 = n101 & n303 ;
  assign n307 = n203 & ~n303 ;
  assign n309 = n308 ^ n307 ;
  assign n392 = x24 & n390 ;
  assign n391 = n311 & ~n390 ;
  assign n393 = n392 ^ n391 ;
  assign n395 = n393 ^ n309 ;
  assign n400 = n211 & n303 ;
  assign n399 = n209 & ~n303 ;
  assign n401 = n400 ^ n399 ;
  assign n397 = x25 & n390 ;
  assign n396 = n315 & ~n390 ;
  assign n398 = n397 ^ n396 ;
  assign n405 = n401 ^ n398 ;
  assign n406 = ~n395 & ~n405 ;
  assign n411 = x26 & n390 ;
  assign n410 = n324 & ~n390 ;
  assign n412 = n411 ^ n410 ;
  assign n408 = n220 & n303 ;
  assign n407 = n224 & ~n303 ;
  assign n409 = n408 ^ n407 ;
  assign n414 = n412 ^ n409 ;
  assign n419 = x27 & n390 ;
  assign n418 = n328 & ~n390 ;
  assign n420 = n419 ^ n418 ;
  assign n416 = n228 & n303 ;
  assign n415 = n232 & ~n303 ;
  assign n417 = n416 ^ n415 ;
  assign n426 = n420 ^ n417 ;
  assign n427 = ~n414 & ~n426 ;
  assign n428 = n406 & n427 ;
  assign n433 = x28 & n390 ;
  assign n432 = n342 & ~n390 ;
  assign n434 = n433 ^ n432 ;
  assign n430 = n246 & n303 ;
  assign n429 = n250 & ~n303 ;
  assign n431 = n430 ^ n429 ;
  assign n436 = n434 ^ n431 ;
  assign n441 = x29 & n390 ;
  assign n440 = n346 & ~n390 ;
  assign n442 = n441 ^ n440 ;
  assign n438 = n254 & n303 ;
  assign n437 = n258 & ~n303 ;
  assign n439 = n438 ^ n437 ;
  assign n446 = n442 ^ n439 ;
  assign n447 = ~n436 & ~n446 ;
  assign n452 = x30 & n390 ;
  assign n451 = n382 & ~n390 ;
  assign n453 = n452 ^ n451 ;
  assign n449 = n269 & n303 ;
  assign n448 = n273 & ~n303 ;
  assign n450 = n449 ^ n448 ;
  assign n455 = n453 ^ n450 ;
  assign n462 = n278 & n303 ;
  assign n460 = n296 & n303 ;
  assign n461 = n460 ^ n296 ;
  assign n463 = n462 ^ n461 ;
  assign n457 = n456 ^ n365 ;
  assign n459 = n458 ^ n457 ;
  assign n473 = n463 ^ n459 ;
  assign n474 = ~n455 & ~n473 ;
  assign n475 = n447 & n474 ;
  assign n476 = n428 & n475 ;
  assign n464 = n459 & n463 ;
  assign n465 = n464 ^ n463 ;
  assign n466 = n455 & n465 ;
  assign n467 = n466 ^ n465 ;
  assign n454 = n450 & ~n453 ;
  assign n468 = n467 ^ n454 ;
  assign n469 = n447 & n468 ;
  assign n443 = n439 & ~n442 ;
  assign n444 = ~n436 & n443 ;
  assign n435 = n431 & ~n434 ;
  assign n445 = n444 ^ n435 ;
  assign n470 = n469 ^ n445 ;
  assign n471 = n428 & n470 ;
  assign n421 = n417 & ~n420 ;
  assign n422 = ~n414 & n421 ;
  assign n413 = n409 & ~n412 ;
  assign n423 = n422 ^ n413 ;
  assign n424 = n406 & n423 ;
  assign n402 = ~n398 & n401 ;
  assign n403 = ~n395 & n402 ;
  assign n394 = n309 & ~n393 ;
  assign n404 = n403 ^ n394 ;
  assign n425 = n424 ^ n404 ;
  assign n472 = n471 ^ n425 ;
  assign n477 = n476 ^ n472 ;
  assign n574 = n309 & n477 ;
  assign n573 = n393 & ~n477 ;
  assign n575 = n574 ^ n573 ;
  assign n652 = x32 & n650 ;
  assign n651 = n578 & ~n650 ;
  assign n653 = n652 ^ n651 ;
  assign n655 = n653 ^ n575 ;
  assign n660 = n401 & n477 ;
  assign n659 = n398 & ~n477 ;
  assign n661 = n660 ^ n659 ;
  assign n657 = x33 & n650 ;
  assign n656 = n583 & ~n650 ;
  assign n658 = n657 ^ n656 ;
  assign n665 = n661 ^ n658 ;
  assign n666 = ~n655 & ~n665 ;
  assign n671 = x34 & n650 ;
  assign n670 = n591 & ~n650 ;
  assign n672 = n671 ^ n670 ;
  assign n668 = n409 & n477 ;
  assign n667 = n412 & ~n477 ;
  assign n669 = n668 ^ n667 ;
  assign n674 = n672 ^ n669 ;
  assign n679 = x35 & n650 ;
  assign n678 = n596 & ~n650 ;
  assign n680 = n679 ^ n678 ;
  assign n676 = n417 & n477 ;
  assign n675 = n420 & ~n477 ;
  assign n677 = n676 ^ n675 ;
  assign n686 = n680 ^ n677 ;
  assign n687 = ~n674 & ~n686 ;
  assign n688 = n666 & n687 ;
  assign n693 = x36 & n650 ;
  assign n692 = n607 & ~n650 ;
  assign n694 = n693 ^ n692 ;
  assign n690 = n431 & n477 ;
  assign n689 = n434 & ~n477 ;
  assign n691 = n690 ^ n689 ;
  assign n696 = n694 ^ n691 ;
  assign n701 = x37 & n650 ;
  assign n700 = n612 & ~n650 ;
  assign n702 = n701 ^ n700 ;
  assign n698 = n439 & n477 ;
  assign n697 = n442 & ~n477 ;
  assign n699 = n698 ^ n697 ;
  assign n706 = n702 ^ n699 ;
  assign n707 = ~n696 & ~n706 ;
  assign n712 = x38 & n650 ;
  assign n711 = n644 & ~n650 ;
  assign n713 = n712 ^ n711 ;
  assign n709 = n450 & n477 ;
  assign n708 = n453 & ~n477 ;
  assign n710 = n709 ^ n708 ;
  assign n715 = n713 ^ n710 ;
  assign n560 = n459 & n477 ;
  assign n720 = n560 ^ n459 ;
  assign n558 = n463 & n477 ;
  assign n721 = n720 ^ n558 ;
  assign n717 = n716 ^ n626 ;
  assign n719 = n718 ^ n717 ;
  assign n731 = n721 ^ n719 ;
  assign n732 = ~n715 & ~n731 ;
  assign n733 = n707 & n732 ;
  assign n734 = n688 & n733 ;
  assign n722 = n719 & n721 ;
  assign n723 = n722 ^ n721 ;
  assign n724 = n715 & n723 ;
  assign n725 = n724 ^ n723 ;
  assign n714 = n710 & ~n713 ;
  assign n726 = n725 ^ n714 ;
  assign n727 = n707 & n726 ;
  assign n703 = n699 & ~n702 ;
  assign n704 = ~n696 & n703 ;
  assign n695 = n691 & ~n694 ;
  assign n705 = n704 ^ n695 ;
  assign n728 = n727 ^ n705 ;
  assign n729 = n688 & n728 ;
  assign n681 = n677 & ~n680 ;
  assign n682 = ~n674 & n681 ;
  assign n673 = n669 & ~n672 ;
  assign n683 = n682 ^ n673 ;
  assign n684 = n666 & n683 ;
  assign n662 = ~n658 & n661 ;
  assign n663 = ~n655 & n662 ;
  assign n654 = n575 & ~n653 ;
  assign n664 = n663 ^ n654 ;
  assign n685 = n684 ^ n664 ;
  assign n730 = n729 ^ n685 ;
  assign n735 = n734 ^ n730 ;
  assign n922 = n575 & n735 ;
  assign n921 = n653 & ~n735 ;
  assign n923 = n922 ^ n921 ;
  assign n1003 = n1001 ^ n923 ;
  assign n1008 = x41 & n998 ;
  assign n1007 = n931 & ~n998 ;
  assign n1009 = n1008 ^ n1007 ;
  assign n1005 = n661 & n735 ;
  assign n1004 = n658 & ~n735 ;
  assign n1006 = n1005 ^ n1004 ;
  assign n1013 = n1009 ^ n1006 ;
  assign n1014 = ~n1003 & ~n1013 ;
  assign n1019 = x42 & n998 ;
  assign n1018 = n939 & ~n998 ;
  assign n1020 = n1019 ^ n1018 ;
  assign n1016 = n669 & n735 ;
  assign n1015 = n672 & ~n735 ;
  assign n1017 = n1016 ^ n1015 ;
  assign n1022 = n1020 ^ n1017 ;
  assign n1027 = x43 & n998 ;
  assign n1026 = n944 & ~n998 ;
  assign n1028 = n1027 ^ n1026 ;
  assign n1024 = n677 & n735 ;
  assign n1023 = n680 & ~n735 ;
  assign n1025 = n1024 ^ n1023 ;
  assign n1034 = n1028 ^ n1025 ;
  assign n1035 = ~n1022 & ~n1034 ;
  assign n1036 = n1014 & n1035 ;
  assign n1041 = x44 & n998 ;
  assign n1040 = n955 & ~n998 ;
  assign n1042 = n1041 ^ n1040 ;
  assign n1038 = n691 & n735 ;
  assign n1037 = n694 & ~n735 ;
  assign n1039 = n1038 ^ n1037 ;
  assign n1044 = n1042 ^ n1039 ;
  assign n1049 = x45 & n998 ;
  assign n1048 = n960 & ~n998 ;
  assign n1050 = n1049 ^ n1048 ;
  assign n1046 = n699 & n735 ;
  assign n1045 = n702 & ~n735 ;
  assign n1047 = n1046 ^ n1045 ;
  assign n1054 = n1050 ^ n1047 ;
  assign n1055 = ~n1044 & ~n1054 ;
  assign n1060 = x46 & n998 ;
  assign n1059 = n992 & ~n998 ;
  assign n1061 = n1060 ^ n1059 ;
  assign n1057 = n710 & n735 ;
  assign n1056 = n713 & ~n735 ;
  assign n1058 = n1057 ^ n1056 ;
  assign n1063 = n1061 ^ n1058 ;
  assign n1068 = x47 & n998 ;
  assign n1066 = n974 & n998 ;
  assign n1067 = n1066 ^ n974 ;
  assign n1069 = n1068 ^ n1067 ;
  assign n803 = n719 & n735 ;
  assign n1064 = n803 ^ n719 ;
  assign n801 = n721 & n735 ;
  assign n1065 = n1064 ^ n801 ;
  assign n1079 = n1069 ^ n1065 ;
  assign n1080 = ~n1063 & ~n1079 ;
  assign n1081 = n1055 & n1080 ;
  assign n1082 = n1036 & n1081 ;
  assign n1070 = n1065 & n1069 ;
  assign n1071 = n1070 ^ n1065 ;
  assign n1072 = n1063 & n1071 ;
  assign n1073 = n1072 ^ n1071 ;
  assign n1062 = n1058 & ~n1061 ;
  assign n1074 = n1073 ^ n1062 ;
  assign n1075 = n1055 & n1074 ;
  assign n1051 = n1047 & ~n1050 ;
  assign n1052 = ~n1044 & n1051 ;
  assign n1043 = n1039 & ~n1042 ;
  assign n1053 = n1052 ^ n1043 ;
  assign n1076 = n1075 ^ n1053 ;
  assign n1077 = n1036 & n1076 ;
  assign n1029 = n1025 & ~n1028 ;
  assign n1030 = ~n1022 & n1029 ;
  assign n1021 = n1017 & ~n1020 ;
  assign n1031 = n1030 ^ n1021 ;
  assign n1032 = n1014 & n1031 ;
  assign n1010 = n1006 & ~n1009 ;
  assign n1011 = ~n1003 & n1010 ;
  assign n1002 = n923 & ~n1001 ;
  assign n1012 = n1011 ^ n1002 ;
  assign n1033 = n1032 ^ n1012 ;
  assign n1078 = n1077 ^ n1033 ;
  assign n1083 = n1082 ^ n1078 ;
  assign n1085 = n1001 & n1083 ;
  assign n1084 = n923 & ~n1083 ;
  assign n1086 = n1085 ^ n1084 ;
  assign n305 = n203 & n303 ;
  assign n304 = n101 & ~n303 ;
  assign n306 = n305 ^ n304 ;
  assign n479 = n393 & n477 ;
  assign n478 = n309 & ~n477 ;
  assign n480 = n479 ^ n478 ;
  assign n482 = n480 ^ n306 ;
  assign n487 = n209 & n303 ;
  assign n486 = n211 & ~n303 ;
  assign n488 = n487 ^ n486 ;
  assign n484 = n398 & n477 ;
  assign n483 = n401 & ~n477 ;
  assign n485 = n484 ^ n483 ;
  assign n492 = n488 ^ n485 ;
  assign n493 = ~n482 & ~n492 ;
  assign n498 = n412 & n477 ;
  assign n497 = n409 & ~n477 ;
  assign n499 = n498 ^ n497 ;
  assign n495 = n224 & n303 ;
  assign n494 = n220 & ~n303 ;
  assign n496 = n495 ^ n494 ;
  assign n501 = n499 ^ n496 ;
  assign n506 = n420 & n477 ;
  assign n505 = n417 & ~n477 ;
  assign n507 = n506 ^ n505 ;
  assign n503 = n232 & n303 ;
  assign n502 = n228 & ~n303 ;
  assign n504 = n503 ^ n502 ;
  assign n513 = n507 ^ n504 ;
  assign n514 = ~n501 & ~n513 ;
  assign n515 = n493 & n514 ;
  assign n520 = n434 & n477 ;
  assign n519 = n431 & ~n477 ;
  assign n521 = n520 ^ n519 ;
  assign n517 = n250 & n303 ;
  assign n516 = n246 & ~n303 ;
  assign n518 = n517 ^ n516 ;
  assign n523 = n521 ^ n518 ;
  assign n528 = n442 & n477 ;
  assign n527 = n439 & ~n477 ;
  assign n529 = n528 ^ n527 ;
  assign n525 = n258 & n303 ;
  assign n524 = n254 & ~n303 ;
  assign n526 = n525 ^ n524 ;
  assign n533 = n529 ^ n526 ;
  assign n534 = ~n523 & ~n533 ;
  assign n539 = n453 & n477 ;
  assign n538 = n450 & ~n477 ;
  assign n540 = n539 ^ n538 ;
  assign n536 = n273 & n303 ;
  assign n535 = n269 & ~n303 ;
  assign n537 = n536 ^ n535 ;
  assign n542 = n540 ^ n537 ;
  assign n559 = n558 ^ n463 ;
  assign n561 = n560 ^ n559 ;
  assign n543 = n278 & ~n303 ;
  assign n544 = n543 ^ n460 ;
  assign n562 = n561 ^ n544 ;
  assign n563 = ~n542 & ~n562 ;
  assign n564 = n534 & n563 ;
  assign n565 = n515 & n564 ;
  assign n547 = n459 & n544 ;
  assign n548 = n477 & n547 ;
  assign n545 = n463 & n544 ;
  assign n546 = ~n477 & n545 ;
  assign n549 = n548 ^ n546 ;
  assign n550 = n549 ^ n544 ;
  assign n551 = n542 & n550 ;
  assign n552 = n551 ^ n550 ;
  assign n541 = n537 & ~n540 ;
  assign n553 = n552 ^ n541 ;
  assign n554 = n534 & n553 ;
  assign n530 = n526 & ~n529 ;
  assign n531 = ~n523 & n530 ;
  assign n522 = n518 & ~n521 ;
  assign n532 = n531 ^ n522 ;
  assign n555 = n554 ^ n532 ;
  assign n556 = n515 & n555 ;
  assign n508 = n504 & ~n507 ;
  assign n509 = ~n501 & n508 ;
  assign n500 = n496 & ~n499 ;
  assign n510 = n509 ^ n500 ;
  assign n511 = n493 & n510 ;
  assign n489 = ~n485 & n488 ;
  assign n490 = ~n482 & n489 ;
  assign n481 = n306 & ~n480 ;
  assign n491 = n490 ^ n481 ;
  assign n512 = n511 ^ n491 ;
  assign n557 = n556 ^ n512 ;
  assign n566 = n565 ^ n557 ;
  assign n571 = n306 & n566 ;
  assign n570 = n480 & ~n566 ;
  assign n572 = n571 ^ n570 ;
  assign n737 = n653 & n735 ;
  assign n736 = n575 & ~n735 ;
  assign n738 = n737 ^ n736 ;
  assign n740 = n738 ^ n572 ;
  assign n745 = n488 & n566 ;
  assign n744 = n485 & ~n566 ;
  assign n746 = n745 ^ n744 ;
  assign n742 = n658 & n735 ;
  assign n741 = n661 & ~n735 ;
  assign n743 = n742 ^ n741 ;
  assign n750 = n746 ^ n743 ;
  assign n751 = ~n740 & ~n750 ;
  assign n756 = n672 & n735 ;
  assign n755 = n669 & ~n735 ;
  assign n757 = n756 ^ n755 ;
  assign n753 = n496 & n566 ;
  assign n752 = n499 & ~n566 ;
  assign n754 = n753 ^ n752 ;
  assign n759 = n757 ^ n754 ;
  assign n764 = n680 & n735 ;
  assign n763 = n677 & ~n735 ;
  assign n765 = n764 ^ n763 ;
  assign n761 = n504 & n566 ;
  assign n760 = n507 & ~n566 ;
  assign n762 = n761 ^ n760 ;
  assign n771 = n765 ^ n762 ;
  assign n772 = ~n759 & ~n771 ;
  assign n773 = n751 & n772 ;
  assign n778 = n694 & n735 ;
  assign n777 = n691 & ~n735 ;
  assign n779 = n778 ^ n777 ;
  assign n775 = n518 & n566 ;
  assign n774 = n521 & ~n566 ;
  assign n776 = n775 ^ n774 ;
  assign n781 = n779 ^ n776 ;
  assign n786 = n702 & n735 ;
  assign n785 = n699 & ~n735 ;
  assign n787 = n786 ^ n785 ;
  assign n783 = n526 & n566 ;
  assign n782 = n529 & ~n566 ;
  assign n784 = n783 ^ n782 ;
  assign n791 = n787 ^ n784 ;
  assign n792 = ~n781 & ~n791 ;
  assign n797 = n713 & n735 ;
  assign n796 = n710 & ~n735 ;
  assign n798 = n797 ^ n796 ;
  assign n794 = n537 & n566 ;
  assign n793 = n540 & ~n566 ;
  assign n795 = n794 ^ n793 ;
  assign n800 = n798 ^ n795 ;
  assign n807 = n544 & n566 ;
  assign n805 = n561 & n566 ;
  assign n806 = n805 ^ n561 ;
  assign n808 = n807 ^ n806 ;
  assign n802 = n801 ^ n721 ;
  assign n804 = n803 ^ n802 ;
  assign n818 = n808 ^ n804 ;
  assign n819 = ~n800 & ~n818 ;
  assign n820 = n792 & n819 ;
  assign n821 = n773 & n820 ;
  assign n809 = n804 & n808 ;
  assign n810 = n809 ^ n808 ;
  assign n811 = n800 & n810 ;
  assign n812 = n811 ^ n810 ;
  assign n799 = n795 & ~n798 ;
  assign n813 = n812 ^ n799 ;
  assign n814 = n792 & n813 ;
  assign n788 = n784 & ~n787 ;
  assign n789 = ~n781 & n788 ;
  assign n780 = n776 & ~n779 ;
  assign n790 = n789 ^ n780 ;
  assign n815 = n814 ^ n790 ;
  assign n816 = n773 & n815 ;
  assign n766 = n762 & ~n765 ;
  assign n767 = ~n759 & n766 ;
  assign n758 = n754 & ~n757 ;
  assign n768 = n767 ^ n758 ;
  assign n769 = n751 & n768 ;
  assign n747 = ~n743 & n746 ;
  assign n748 = ~n740 & n747 ;
  assign n739 = n572 & ~n738 ;
  assign n749 = n748 ^ n739 ;
  assign n770 = n769 ^ n749 ;
  assign n817 = n816 ^ n770 ;
  assign n822 = n821 ^ n817 ;
  assign n919 = n572 & n822 ;
  assign n918 = n738 & ~n822 ;
  assign n920 = n919 ^ n918 ;
  assign n1088 = n1086 ^ n920 ;
  assign n1093 = n1009 & n1083 ;
  assign n1092 = n1006 & ~n1083 ;
  assign n1094 = n1093 ^ n1092 ;
  assign n1090 = n746 & n822 ;
  assign n1089 = n743 & ~n822 ;
  assign n1091 = n1090 ^ n1089 ;
  assign n1098 = n1094 ^ n1091 ;
  assign n1099 = ~n1088 & ~n1098 ;
  assign n1104 = n1020 & n1083 ;
  assign n1103 = n1017 & ~n1083 ;
  assign n1105 = n1104 ^ n1103 ;
  assign n1101 = n754 & n822 ;
  assign n1100 = n757 & ~n822 ;
  assign n1102 = n1101 ^ n1100 ;
  assign n1107 = n1105 ^ n1102 ;
  assign n1112 = n1028 & n1083 ;
  assign n1111 = n1025 & ~n1083 ;
  assign n1113 = n1112 ^ n1111 ;
  assign n1109 = n762 & n822 ;
  assign n1108 = n765 & ~n822 ;
  assign n1110 = n1109 ^ n1108 ;
  assign n1119 = n1113 ^ n1110 ;
  assign n1120 = ~n1107 & ~n1119 ;
  assign n1121 = n1099 & n1120 ;
  assign n1126 = n1042 & n1083 ;
  assign n1125 = n1039 & ~n1083 ;
  assign n1127 = n1126 ^ n1125 ;
  assign n1123 = n776 & n822 ;
  assign n1122 = n779 & ~n822 ;
  assign n1124 = n1123 ^ n1122 ;
  assign n1129 = n1127 ^ n1124 ;
  assign n1134 = n1050 & n1083 ;
  assign n1133 = n1047 & ~n1083 ;
  assign n1135 = n1134 ^ n1133 ;
  assign n1131 = n784 & n822 ;
  assign n1130 = n787 & ~n822 ;
  assign n1132 = n1131 ^ n1130 ;
  assign n1139 = n1135 ^ n1132 ;
  assign n1140 = ~n1129 & ~n1139 ;
  assign n1145 = n1061 & n1083 ;
  assign n1144 = n1058 & ~n1083 ;
  assign n1146 = n1145 ^ n1144 ;
  assign n1142 = n795 & n822 ;
  assign n1141 = n798 & ~n822 ;
  assign n1143 = n1142 ^ n1141 ;
  assign n1148 = n1146 ^ n1143 ;
  assign n1153 = n1069 & n1083 ;
  assign n1151 = n1065 & n1083 ;
  assign n1152 = n1151 ^ n1065 ;
  assign n1154 = n1153 ^ n1152 ;
  assign n905 = n804 & n822 ;
  assign n1149 = n905 ^ n804 ;
  assign n903 = n808 & n822 ;
  assign n1150 = n1149 ^ n903 ;
  assign n1164 = n1154 ^ n1150 ;
  assign n1165 = ~n1148 & ~n1164 ;
  assign n1166 = n1140 & n1165 ;
  assign n1167 = n1121 & n1166 ;
  assign n1155 = n1150 & n1154 ;
  assign n1156 = n1155 ^ n1150 ;
  assign n1157 = n1148 & n1156 ;
  assign n1158 = n1157 ^ n1156 ;
  assign n1147 = n1143 & ~n1146 ;
  assign n1159 = n1158 ^ n1147 ;
  assign n1160 = n1140 & n1159 ;
  assign n1136 = n1132 & ~n1135 ;
  assign n1137 = ~n1129 & n1136 ;
  assign n1128 = n1124 & ~n1127 ;
  assign n1138 = n1137 ^ n1128 ;
  assign n1161 = n1160 ^ n1138 ;
  assign n1162 = n1121 & n1161 ;
  assign n1114 = n1110 & ~n1113 ;
  assign n1115 = ~n1107 & n1114 ;
  assign n1106 = n1102 & ~n1105 ;
  assign n1116 = n1115 ^ n1106 ;
  assign n1117 = n1099 & n1116 ;
  assign n1095 = n1091 & ~n1094 ;
  assign n1096 = ~n1088 & n1095 ;
  assign n1087 = n920 & ~n1086 ;
  assign n1097 = n1096 ^ n1087 ;
  assign n1118 = n1117 ^ n1097 ;
  assign n1163 = n1162 ^ n1118 ;
  assign n1168 = n1167 ^ n1163 ;
  assign n1170 = n1086 & n1168 ;
  assign n1169 = n920 & ~n1168 ;
  assign n1171 = n1170 ^ n1169 ;
  assign n568 = n480 & n566 ;
  assign n567 = n306 & ~n566 ;
  assign n569 = n568 ^ n567 ;
  assign n824 = n738 & n822 ;
  assign n823 = n572 & ~n822 ;
  assign n825 = n824 ^ n823 ;
  assign n827 = n825 ^ n569 ;
  assign n832 = n485 & n566 ;
  assign n831 = n488 & ~n566 ;
  assign n833 = n832 ^ n831 ;
  assign n829 = n743 & n822 ;
  assign n828 = n746 & ~n822 ;
  assign n830 = n829 ^ n828 ;
  assign n837 = n833 ^ n830 ;
  assign n838 = ~n827 & ~n837 ;
  assign n843 = n757 & n822 ;
  assign n842 = n754 & ~n822 ;
  assign n844 = n843 ^ n842 ;
  assign n840 = n499 & n566 ;
  assign n839 = n496 & ~n566 ;
  assign n841 = n840 ^ n839 ;
  assign n846 = n844 ^ n841 ;
  assign n851 = n765 & n822 ;
  assign n850 = n762 & ~n822 ;
  assign n852 = n851 ^ n850 ;
  assign n848 = n507 & n566 ;
  assign n847 = n504 & ~n566 ;
  assign n849 = n848 ^ n847 ;
  assign n858 = n852 ^ n849 ;
  assign n859 = ~n846 & ~n858 ;
  assign n860 = n838 & n859 ;
  assign n865 = n779 & n822 ;
  assign n864 = n776 & ~n822 ;
  assign n866 = n865 ^ n864 ;
  assign n862 = n521 & n566 ;
  assign n861 = n518 & ~n566 ;
  assign n863 = n862 ^ n861 ;
  assign n868 = n866 ^ n863 ;
  assign n873 = n787 & n822 ;
  assign n872 = n784 & ~n822 ;
  assign n874 = n873 ^ n872 ;
  assign n870 = n529 & n566 ;
  assign n869 = n526 & ~n566 ;
  assign n871 = n870 ^ n869 ;
  assign n878 = n874 ^ n871 ;
  assign n879 = ~n868 & ~n878 ;
  assign n884 = n798 & n822 ;
  assign n883 = n795 & ~n822 ;
  assign n885 = n884 ^ n883 ;
  assign n881 = n540 & n566 ;
  assign n880 = n537 & ~n566 ;
  assign n882 = n881 ^ n880 ;
  assign n887 = n885 ^ n882 ;
  assign n904 = n903 ^ n808 ;
  assign n906 = n905 ^ n904 ;
  assign n888 = n544 & ~n566 ;
  assign n889 = n888 ^ n805 ;
  assign n907 = n906 ^ n889 ;
  assign n908 = ~n887 & ~n907 ;
  assign n909 = n879 & n908 ;
  assign n910 = n860 & n909 ;
  assign n892 = n804 & n889 ;
  assign n893 = n822 & n892 ;
  assign n890 = n808 & n889 ;
  assign n891 = ~n822 & n890 ;
  assign n894 = n893 ^ n891 ;
  assign n895 = n894 ^ n889 ;
  assign n896 = n887 & n895 ;
  assign n897 = n896 ^ n895 ;
  assign n886 = n882 & ~n885 ;
  assign n898 = n897 ^ n886 ;
  assign n899 = n879 & n898 ;
  assign n875 = n871 & ~n874 ;
  assign n876 = ~n868 & n875 ;
  assign n867 = n863 & ~n866 ;
  assign n877 = n876 ^ n867 ;
  assign n900 = n899 ^ n877 ;
  assign n901 = n860 & n900 ;
  assign n853 = n849 & ~n852 ;
  assign n854 = ~n846 & n853 ;
  assign n845 = n841 & ~n844 ;
  assign n855 = n854 ^ n845 ;
  assign n856 = n838 & n855 ;
  assign n834 = ~n830 & n833 ;
  assign n835 = ~n827 & n834 ;
  assign n826 = n569 & ~n825 ;
  assign n836 = n835 ^ n826 ;
  assign n857 = n856 ^ n836 ;
  assign n902 = n901 ^ n857 ;
  assign n911 = n910 ^ n902 ;
  assign n916 = n569 & n911 ;
  assign n915 = n825 & ~n911 ;
  assign n917 = n916 ^ n915 ;
  assign n1173 = n1171 ^ n917 ;
  assign n1178 = n1094 & n1168 ;
  assign n1177 = n1091 & ~n1168 ;
  assign n1179 = n1178 ^ n1177 ;
  assign n1175 = n833 & n911 ;
  assign n1174 = n830 & ~n911 ;
  assign n1176 = n1175 ^ n1174 ;
  assign n1183 = n1179 ^ n1176 ;
  assign n1184 = ~n1173 & ~n1183 ;
  assign n1189 = n1105 & n1168 ;
  assign n1188 = n1102 & ~n1168 ;
  assign n1190 = n1189 ^ n1188 ;
  assign n1186 = n841 & n911 ;
  assign n1185 = n844 & ~n911 ;
  assign n1187 = n1186 ^ n1185 ;
  assign n1192 = n1190 ^ n1187 ;
  assign n1197 = n1113 & n1168 ;
  assign n1196 = n1110 & ~n1168 ;
  assign n1198 = n1197 ^ n1196 ;
  assign n1194 = n849 & n911 ;
  assign n1193 = n852 & ~n911 ;
  assign n1195 = n1194 ^ n1193 ;
  assign n1204 = n1198 ^ n1195 ;
  assign n1205 = ~n1192 & ~n1204 ;
  assign n1206 = n1184 & n1205 ;
  assign n1211 = n1127 & n1168 ;
  assign n1210 = n1124 & ~n1168 ;
  assign n1212 = n1211 ^ n1210 ;
  assign n1208 = n863 & n911 ;
  assign n1207 = n866 & ~n911 ;
  assign n1209 = n1208 ^ n1207 ;
  assign n1214 = n1212 ^ n1209 ;
  assign n1219 = n1135 & n1168 ;
  assign n1218 = n1132 & ~n1168 ;
  assign n1220 = n1219 ^ n1218 ;
  assign n1216 = n871 & n911 ;
  assign n1215 = n874 & ~n911 ;
  assign n1217 = n1216 ^ n1215 ;
  assign n1224 = n1220 ^ n1217 ;
  assign n1225 = ~n1214 & ~n1224 ;
  assign n1230 = n1146 & n1168 ;
  assign n1229 = n1143 & ~n1168 ;
  assign n1231 = n1230 ^ n1229 ;
  assign n1227 = n882 & n911 ;
  assign n1226 = n885 & ~n911 ;
  assign n1228 = n1227 ^ n1226 ;
  assign n1233 = n1231 ^ n1228 ;
  assign n1240 = n1154 & n1168 ;
  assign n1238 = n1150 & n1168 ;
  assign n1239 = n1238 ^ n1150 ;
  assign n1241 = n1240 ^ n1239 ;
  assign n1236 = n889 & n911 ;
  assign n1234 = n906 & n911 ;
  assign n1235 = n1234 ^ n906 ;
  assign n1237 = n1236 ^ n1235 ;
  assign n1251 = n1241 ^ n1237 ;
  assign n1252 = ~n1233 & ~n1251 ;
  assign n1253 = n1225 & n1252 ;
  assign n1254 = n1206 & n1253 ;
  assign n1242 = n1237 & n1241 ;
  assign n1243 = n1242 ^ n1237 ;
  assign n1244 = n1233 & n1243 ;
  assign n1245 = n1244 ^ n1243 ;
  assign n1232 = n1228 & ~n1231 ;
  assign n1246 = n1245 ^ n1232 ;
  assign n1247 = n1225 & n1246 ;
  assign n1221 = n1217 & ~n1220 ;
  assign n1222 = ~n1214 & n1221 ;
  assign n1213 = n1209 & ~n1212 ;
  assign n1223 = n1222 ^ n1213 ;
  assign n1248 = n1247 ^ n1223 ;
  assign n1249 = n1206 & n1248 ;
  assign n1199 = n1195 & ~n1198 ;
  assign n1200 = ~n1192 & n1199 ;
  assign n1191 = n1187 & ~n1190 ;
  assign n1201 = n1200 ^ n1191 ;
  assign n1202 = n1184 & n1201 ;
  assign n1180 = n1176 & ~n1179 ;
  assign n1181 = ~n1173 & n1180 ;
  assign n1172 = n917 & ~n1171 ;
  assign n1182 = n1181 ^ n1172 ;
  assign n1203 = n1202 ^ n1182 ;
  assign n1250 = n1249 ^ n1203 ;
  assign n1255 = n1254 ^ n1250 ;
  assign n1258 = n1171 & n1255 ;
  assign n1256 = n917 & n1255 ;
  assign n1257 = n1256 ^ n917 ;
  assign n1259 = n1258 ^ n1257 ;
  assign n913 = n825 & n911 ;
  assign n912 = n569 & ~n911 ;
  assign n914 = n913 ^ n912 ;
  assign n1261 = n1259 ^ n914 ;
  assign n1267 = n1179 & n1255 ;
  assign n1265 = n1176 & n1255 ;
  assign n1266 = n1265 ^ n1176 ;
  assign n1268 = n1267 ^ n1266 ;
  assign n1263 = n830 & n911 ;
  assign n1262 = n833 & ~n911 ;
  assign n1264 = n1263 ^ n1262 ;
  assign n1272 = n1268 ^ n1264 ;
  assign n1273 = n1261 & n1272 ;
  assign n1274 = n1273 ^ n1261 ;
  assign n1275 = n1274 ^ n1272 ;
  assign n1281 = n1190 & n1255 ;
  assign n1279 = n1187 & n1255 ;
  assign n1280 = n1279 ^ n1187 ;
  assign n1282 = n1281 ^ n1280 ;
  assign n1277 = n844 & n911 ;
  assign n1276 = n841 & ~n911 ;
  assign n1278 = n1277 ^ n1276 ;
  assign n1284 = n1282 ^ n1278 ;
  assign n1290 = n1198 & n1255 ;
  assign n1288 = n1195 & n1255 ;
  assign n1289 = n1288 ^ n1195 ;
  assign n1291 = n1290 ^ n1289 ;
  assign n1286 = n852 & n911 ;
  assign n1285 = n849 & ~n911 ;
  assign n1287 = n1286 ^ n1285 ;
  assign n1299 = n1291 ^ n1287 ;
  assign n1300 = n1284 & n1299 ;
  assign n1301 = n1300 ^ n1284 ;
  assign n1302 = n1301 ^ n1299 ;
  assign n1303 = ~n1275 & ~n1302 ;
  assign n1309 = n1212 & n1255 ;
  assign n1307 = n1209 & n1255 ;
  assign n1308 = n1307 ^ n1209 ;
  assign n1310 = n1309 ^ n1308 ;
  assign n1305 = n866 & n911 ;
  assign n1304 = n863 & ~n911 ;
  assign n1306 = n1305 ^ n1304 ;
  assign n1312 = n1310 ^ n1306 ;
  assign n1318 = n1220 & n1255 ;
  assign n1316 = n1217 & n1255 ;
  assign n1317 = n1316 ^ n1217 ;
  assign n1319 = n1318 ^ n1317 ;
  assign n1314 = n874 & n911 ;
  assign n1313 = n871 & ~n911 ;
  assign n1315 = n1314 ^ n1313 ;
  assign n1325 = n1319 ^ n1315 ;
  assign n1326 = n1312 & n1325 ;
  assign n1327 = n1326 ^ n1312 ;
  assign n1328 = n1327 ^ n1325 ;
  assign n1334 = n1231 & n1255 ;
  assign n1332 = n1228 & n1255 ;
  assign n1333 = n1332 ^ n1228 ;
  assign n1335 = n1334 ^ n1333 ;
  assign n1330 = n885 & n911 ;
  assign n1329 = n882 & ~n911 ;
  assign n1331 = n1330 ^ n1329 ;
  assign n1338 = n1335 ^ n1331 ;
  assign n1356 = n1237 & n1255 ;
  assign n1357 = n1356 ^ n1237 ;
  assign n1355 = n1241 & n1255 ;
  assign n1358 = n1357 ^ n1355 ;
  assign n1339 = n889 & ~n911 ;
  assign n1340 = n1339 ^ n1234 ;
  assign n1359 = n1358 ^ n1340 ;
  assign n1360 = n1338 & n1359 ;
  assign n1361 = n1360 ^ n1338 ;
  assign n1362 = n1361 ^ n1359 ;
  assign n1363 = ~n1328 & ~n1362 ;
  assign n1364 = n1303 & n1363 ;
  assign n1343 = n1237 & n1340 ;
  assign n1344 = n1255 & n1343 ;
  assign n1345 = n1344 ^ n1343 ;
  assign n1341 = n1241 & n1340 ;
  assign n1342 = n1255 & n1341 ;
  assign n1346 = n1345 ^ n1342 ;
  assign n1347 = n1346 ^ n1340 ;
  assign n1348 = n1338 & n1347 ;
  assign n1349 = n1348 ^ n1347 ;
  assign n1336 = n1331 & n1335 ;
  assign n1337 = n1336 ^ n1331 ;
  assign n1350 = n1349 ^ n1337 ;
  assign n1351 = ~n1328 & n1350 ;
  assign n1320 = n1315 & n1319 ;
  assign n1321 = n1320 ^ n1315 ;
  assign n1322 = n1312 & n1321 ;
  assign n1323 = n1322 ^ n1321 ;
  assign n1311 = n1306 & ~n1310 ;
  assign n1324 = n1323 ^ n1311 ;
  assign n1352 = n1351 ^ n1324 ;
  assign n1353 = n1303 & n1352 ;
  assign n1292 = n1287 & n1291 ;
  assign n1293 = n1292 ^ n1287 ;
  assign n1294 = n1284 & n1293 ;
  assign n1295 = n1294 ^ n1293 ;
  assign n1283 = n1278 & ~n1282 ;
  assign n1296 = n1295 ^ n1283 ;
  assign n1297 = ~n1275 & n1296 ;
  assign n1269 = n1264 & ~n1268 ;
  assign n1270 = ~n1261 & n1269 ;
  assign n1260 = n914 & ~n1259 ;
  assign n1271 = n1270 ^ n1260 ;
  assign n1298 = n1297 ^ n1271 ;
  assign n1354 = n1353 ^ n1298 ;
  assign n1365 = n1364 ^ n1354 ;
  assign n1368 = n1259 & n1365 ;
  assign n1366 = n914 & n1365 ;
  assign n1367 = n1366 ^ n914 ;
  assign n1369 = n1368 ^ n1367 ;
  assign n1372 = n1268 & n1365 ;
  assign n1370 = n1264 & n1365 ;
  assign n1371 = n1370 ^ n1264 ;
  assign n1373 = n1372 ^ n1371 ;
  assign n1376 = n1282 & n1365 ;
  assign n1374 = n1278 & n1365 ;
  assign n1375 = n1374 ^ n1278 ;
  assign n1377 = n1376 ^ n1375 ;
  assign n1380 = n1291 & n1365 ;
  assign n1378 = n1287 & n1365 ;
  assign n1379 = n1378 ^ n1287 ;
  assign n1381 = n1380 ^ n1379 ;
  assign n1384 = n1310 & n1365 ;
  assign n1382 = n1306 & n1365 ;
  assign n1383 = n1382 ^ n1306 ;
  assign n1385 = n1384 ^ n1383 ;
  assign n1388 = n1319 & n1365 ;
  assign n1386 = n1315 & n1365 ;
  assign n1387 = n1386 ^ n1315 ;
  assign n1389 = n1388 ^ n1387 ;
  assign n1392 = n1335 & n1365 ;
  assign n1390 = n1331 & n1365 ;
  assign n1391 = n1390 ^ n1331 ;
  assign n1393 = n1392 ^ n1391 ;
  assign n1396 = n1358 & n1365 ;
  assign n1394 = n1340 & n1365 ;
  assign n1395 = n1394 ^ n1340 ;
  assign n1397 = n1396 ^ n1395 ;
  assign n1398 = n1368 ^ n1259 ;
  assign n1399 = n1398 ^ n1366 ;
  assign n1400 = n1372 ^ n1268 ;
  assign n1401 = n1400 ^ n1370 ;
  assign n1402 = n1376 ^ n1282 ;
  assign n1403 = n1402 ^ n1374 ;
  assign n1404 = n1380 ^ n1291 ;
  assign n1405 = n1404 ^ n1378 ;
  assign n1406 = n1384 ^ n1310 ;
  assign n1407 = n1406 ^ n1382 ;
  assign n1408 = n1388 ^ n1319 ;
  assign n1409 = n1408 ^ n1386 ;
  assign n1410 = n1392 ^ n1335 ;
  assign n1411 = n1410 ^ n1390 ;
  assign n1412 = n1396 ^ n1358 ;
  assign n1413 = n1412 ^ n1394 ;
  assign n1414 = n1171 & ~n1255 ;
  assign n1415 = n1414 ^ n1256 ;
  assign n1416 = n1179 & ~n1255 ;
  assign n1417 = n1416 ^ n1265 ;
  assign n1418 = n1190 & ~n1255 ;
  assign n1419 = n1418 ^ n1279 ;
  assign n1420 = n1198 & ~n1255 ;
  assign n1421 = n1420 ^ n1288 ;
  assign n1422 = n1212 & ~n1255 ;
  assign n1423 = n1422 ^ n1307 ;
  assign n1424 = n1220 & ~n1255 ;
  assign n1425 = n1424 ^ n1316 ;
  assign n1426 = n1231 & ~n1255 ;
  assign n1427 = n1426 ^ n1332 ;
  assign n1428 = n1241 & ~n1255 ;
  assign n1429 = n1428 ^ n1356 ;
  assign n1431 = n920 & n1168 ;
  assign n1430 = n1086 & ~n1168 ;
  assign n1432 = n1431 ^ n1430 ;
  assign n1434 = n1091 & n1168 ;
  assign n1433 = n1094 & ~n1168 ;
  assign n1435 = n1434 ^ n1433 ;
  assign n1437 = n1102 & n1168 ;
  assign n1436 = n1105 & ~n1168 ;
  assign n1438 = n1437 ^ n1436 ;
  assign n1440 = n1110 & n1168 ;
  assign n1439 = n1113 & ~n1168 ;
  assign n1441 = n1440 ^ n1439 ;
  assign n1443 = n1124 & n1168 ;
  assign n1442 = n1127 & ~n1168 ;
  assign n1444 = n1443 ^ n1442 ;
  assign n1446 = n1132 & n1168 ;
  assign n1445 = n1135 & ~n1168 ;
  assign n1447 = n1446 ^ n1445 ;
  assign n1449 = n1143 & n1168 ;
  assign n1448 = n1146 & ~n1168 ;
  assign n1450 = n1449 ^ n1448 ;
  assign n1451 = n1154 & ~n1168 ;
  assign n1452 = n1451 ^ n1238 ;
  assign n1454 = n923 & n1083 ;
  assign n1453 = n1001 & ~n1083 ;
  assign n1455 = n1454 ^ n1453 ;
  assign n1457 = n1006 & n1083 ;
  assign n1456 = n1009 & ~n1083 ;
  assign n1458 = n1457 ^ n1456 ;
  assign n1460 = n1017 & n1083 ;
  assign n1459 = n1020 & ~n1083 ;
  assign n1461 = n1460 ^ n1459 ;
  assign n1463 = n1025 & n1083 ;
  assign n1462 = n1028 & ~n1083 ;
  assign n1464 = n1463 ^ n1462 ;
  assign n1466 = n1039 & n1083 ;
  assign n1465 = n1042 & ~n1083 ;
  assign n1467 = n1466 ^ n1465 ;
  assign n1469 = n1047 & n1083 ;
  assign n1468 = n1050 & ~n1083 ;
  assign n1470 = n1469 ^ n1468 ;
  assign n1472 = n1058 & n1083 ;
  assign n1471 = n1061 & ~n1083 ;
  assign n1473 = n1472 ^ n1471 ;
  assign n1474 = n1069 & ~n1083 ;
  assign n1475 = n1474 ^ n1151 ;
  assign n1477 = n926 & n998 ;
  assign n1476 = x40 & ~n998 ;
  assign n1478 = n1477 ^ n1476 ;
  assign n1480 = n931 & n998 ;
  assign n1479 = x41 & ~n998 ;
  assign n1481 = n1480 ^ n1479 ;
  assign n1483 = n939 & n998 ;
  assign n1482 = x42 & ~n998 ;
  assign n1484 = n1483 ^ n1482 ;
  assign n1486 = n944 & n998 ;
  assign n1485 = x43 & ~n998 ;
  assign n1487 = n1486 ^ n1485 ;
  assign n1489 = n955 & n998 ;
  assign n1488 = x44 & ~n998 ;
  assign n1490 = n1489 ^ n1488 ;
  assign n1492 = n960 & n998 ;
  assign n1491 = x45 & ~n998 ;
  assign n1493 = n1492 ^ n1491 ;
  assign n1495 = n992 & n998 ;
  assign n1494 = x46 & ~n998 ;
  assign n1496 = n1495 ^ n1494 ;
  assign n1497 = x47 & ~n998 ;
  assign n1498 = n1497 ^ n1066 ;
  assign y0 = n1369 ;
  assign y1 = n1373 ;
  assign y2 = n1377 ;
  assign y3 = n1381 ;
  assign y4 = n1385 ;
  assign y5 = n1389 ;
  assign y6 = n1393 ;
  assign y7 = n1397 ;
  assign y8 = n1399 ;
  assign y9 = n1401 ;
  assign y10 = n1403 ;
  assign y11 = n1405 ;
  assign y12 = n1407 ;
  assign y13 = n1409 ;
  assign y14 = n1411 ;
  assign y15 = n1413 ;
  assign y16 = n1415 ;
  assign y17 = n1417 ;
  assign y18 = n1419 ;
  assign y19 = n1421 ;
  assign y20 = n1423 ;
  assign y21 = n1425 ;
  assign y22 = n1427 ;
  assign y23 = n1429 ;
  assign y24 = n1432 ;
  assign y25 = n1435 ;
  assign y26 = n1438 ;
  assign y27 = n1441 ;
  assign y28 = n1444 ;
  assign y29 = n1447 ;
  assign y30 = n1450 ;
  assign y31 = n1452 ;
  assign y32 = n1455 ;
  assign y33 = n1458 ;
  assign y34 = n1461 ;
  assign y35 = n1464 ;
  assign y36 = n1467 ;
  assign y37 = n1470 ;
  assign y38 = n1473 ;
  assign y39 = n1475 ;
  assign y40 = n1478 ;
  assign y41 = n1481 ;
  assign y42 = n1484 ;
  assign y43 = n1487 ;
  assign y44 = n1490 ;
  assign y45 = n1493 ;
  assign y46 = n1496 ;
  assign y47 = n1498 ;
endmodule
