module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 ;
  assign n65 = ~x47 & x63 ;
  assign n66 = x47 & ~x63 ;
  assign n67 = ~x46 & x62 ;
  assign n68 = x46 & ~x62 ;
  assign n69 = ~x45 & x61 ;
  assign n70 = x45 & ~x61 ;
  assign n71 = ~x44 & x60 ;
  assign n72 = x44 & ~x60 ;
  assign n73 = ~x43 & x59 ;
  assign n74 = x43 & ~x59 ;
  assign n75 = ~x42 & x58 ;
  assign n76 = x42 & ~x58 ;
  assign n77 = ~x41 & x57 ;
  assign n78 = x41 & ~x57 ;
  assign n79 = ~x40 & x56 ;
  assign n80 = x40 & ~x56 ;
  assign n81 = ~x39 & x55 ;
  assign n82 = x39 & ~x55 ;
  assign n83 = ~x38 & x54 ;
  assign n84 = x38 & ~x54 ;
  assign n85 = ~x37 & x53 ;
  assign n86 = x37 & ~x53 ;
  assign n87 = ~x36 & x52 ;
  assign n88 = x36 & ~x52 ;
  assign n89 = ~x35 & x51 ;
  assign n90 = x35 & ~x51 ;
  assign n91 = ~x34 & x50 ;
  assign n92 = x34 & ~x50 ;
  assign n93 = ~x33 & x49 ;
  assign n94 = x33 & ~x49 ;
  assign n95 = x32 & ~x48 ;
  assign n96 = ~n94 & ~n95 ;
  assign n97 = ~n93 & ~n96 ;
  assign n98 = ~n92 & ~n97 ;
  assign n99 = ~n91 & ~n98 ;
  assign n100 = ~n90 & ~n99 ;
  assign n101 = ~n89 & ~n100 ;
  assign n102 = ~n88 & ~n101 ;
  assign n103 = ~n87 & ~n102 ;
  assign n104 = ~n86 & ~n103 ;
  assign n105 = ~n85 & ~n104 ;
  assign n106 = ~n84 & ~n105 ;
  assign n107 = ~n83 & ~n106 ;
  assign n108 = ~n82 & ~n107 ;
  assign n109 = ~n81 & ~n108 ;
  assign n110 = ~n80 & ~n109 ;
  assign n111 = ~n79 & ~n110 ;
  assign n112 = ~n78 & ~n111 ;
  assign n113 = ~n77 & ~n112 ;
  assign n114 = ~n76 & ~n113 ;
  assign n115 = ~n75 & ~n114 ;
  assign n116 = ~n74 & ~n115 ;
  assign n117 = ~n73 & ~n116 ;
  assign n118 = ~n72 & ~n117 ;
  assign n119 = ~n71 & ~n118 ;
  assign n120 = ~n70 & ~n119 ;
  assign n121 = ~n69 & ~n120 ;
  assign n122 = ~n68 & ~n121 ;
  assign n123 = ~n67 & ~n122 ;
  assign n124 = ~n66 & ~n123 ;
  assign n125 = ~n65 & ~n124 ;
  assign n126 = ~x47 & ~x63 ;
  assign n127 = ~x15 & ~x31 ;
  assign n128 = ~n126 & n127 ;
  assign n129 = n126 & ~n127 ;
  assign n130 = x62 & ~n125 ;
  assign n131 = x46 & n125 ;
  assign n132 = ~n130 & ~n131 ;
  assign n133 = ~x15 & x31 ;
  assign n134 = x15 & ~x31 ;
  assign n135 = ~x14 & x30 ;
  assign n136 = x14 & ~x30 ;
  assign n137 = ~x13 & x29 ;
  assign n138 = x13 & ~x29 ;
  assign n139 = ~x12 & x28 ;
  assign n140 = x12 & ~x28 ;
  assign n141 = ~x11 & x27 ;
  assign n142 = x11 & ~x27 ;
  assign n143 = ~x10 & x26 ;
  assign n144 = x10 & ~x26 ;
  assign n145 = ~x9 & x25 ;
  assign n146 = x9 & ~x25 ;
  assign n147 = ~x8 & x24 ;
  assign n148 = x8 & ~x24 ;
  assign n149 = ~x7 & x23 ;
  assign n150 = x7 & ~x23 ;
  assign n151 = ~x6 & x22 ;
  assign n152 = x6 & ~x22 ;
  assign n153 = ~x5 & x21 ;
  assign n154 = x5 & ~x21 ;
  assign n155 = ~x4 & x20 ;
  assign n156 = x4 & ~x20 ;
  assign n157 = ~x3 & x19 ;
  assign n158 = x3 & ~x19 ;
  assign n159 = ~x2 & x18 ;
  assign n160 = x2 & ~x18 ;
  assign n161 = ~x1 & x17 ;
  assign n162 = x1 & ~x17 ;
  assign n163 = x0 & ~x16 ;
  assign n164 = ~n162 & ~n163 ;
  assign n165 = ~n161 & ~n164 ;
  assign n166 = ~n160 & ~n165 ;
  assign n167 = ~n159 & ~n166 ;
  assign n168 = ~n158 & ~n167 ;
  assign n169 = ~n157 & ~n168 ;
  assign n170 = ~n156 & ~n169 ;
  assign n171 = ~n155 & ~n170 ;
  assign n172 = ~n154 & ~n171 ;
  assign n173 = ~n153 & ~n172 ;
  assign n174 = ~n152 & ~n173 ;
  assign n175 = ~n151 & ~n174 ;
  assign n176 = ~n150 & ~n175 ;
  assign n177 = ~n149 & ~n176 ;
  assign n178 = ~n148 & ~n177 ;
  assign n179 = ~n147 & ~n178 ;
  assign n180 = ~n146 & ~n179 ;
  assign n181 = ~n145 & ~n180 ;
  assign n182 = ~n144 & ~n181 ;
  assign n183 = ~n143 & ~n182 ;
  assign n184 = ~n142 & ~n183 ;
  assign n185 = ~n141 & ~n184 ;
  assign n186 = ~n140 & ~n185 ;
  assign n187 = ~n139 & ~n186 ;
  assign n188 = ~n138 & ~n187 ;
  assign n189 = ~n137 & ~n188 ;
  assign n190 = ~n136 & ~n189 ;
  assign n191 = ~n135 & ~n190 ;
  assign n192 = ~n134 & ~n191 ;
  assign n193 = ~n133 & ~n192 ;
  assign n194 = x30 & ~n193 ;
  assign n195 = x14 & n193 ;
  assign n196 = ~n194 & ~n195 ;
  assign n197 = ~n132 & n196 ;
  assign n198 = x49 & ~n125 ;
  assign n199 = x33 & n125 ;
  assign n200 = ~n198 & ~n199 ;
  assign n201 = x17 & ~n193 ;
  assign n202 = x1 & n193 ;
  assign n203 = ~n201 & ~n202 ;
  assign n204 = ~n200 & n203 ;
  assign n205 = x48 & ~n125 ;
  assign n206 = x32 & n125 ;
  assign n207 = ~n205 & ~n206 ;
  assign n208 = x16 & ~n193 ;
  assign n209 = x0 & n193 ;
  assign n210 = ~n208 & ~n209 ;
  assign n211 = n207 & ~n210 ;
  assign n212 = ~n204 & n211 ;
  assign n213 = x50 & ~n125 ;
  assign n214 = x34 & n125 ;
  assign n215 = ~n213 & ~n214 ;
  assign n216 = x18 & ~n193 ;
  assign n217 = x2 & n193 ;
  assign n218 = ~n216 & ~n217 ;
  assign n219 = n215 & ~n218 ;
  assign n220 = n200 & ~n203 ;
  assign n221 = ~n219 & ~n220 ;
  assign n222 = ~n212 & n221 ;
  assign n223 = x51 & ~n125 ;
  assign n224 = x35 & n125 ;
  assign n225 = ~n223 & ~n224 ;
  assign n226 = x19 & ~n193 ;
  assign n227 = x3 & n193 ;
  assign n228 = ~n226 & ~n227 ;
  assign n229 = ~n225 & n228 ;
  assign n230 = ~n215 & n218 ;
  assign n231 = ~n229 & ~n230 ;
  assign n232 = ~n222 & n231 ;
  assign n233 = x52 & ~n125 ;
  assign n234 = x36 & n125 ;
  assign n235 = ~n233 & ~n234 ;
  assign n236 = x20 & ~n193 ;
  assign n237 = x4 & n193 ;
  assign n238 = ~n236 & ~n237 ;
  assign n239 = n235 & ~n238 ;
  assign n240 = n225 & ~n228 ;
  assign n241 = ~n239 & ~n240 ;
  assign n242 = ~n232 & n241 ;
  assign n243 = ~n235 & n238 ;
  assign n244 = x53 & ~n125 ;
  assign n245 = x37 & n125 ;
  assign n246 = ~n244 & ~n245 ;
  assign n247 = x21 & ~n193 ;
  assign n248 = x5 & n193 ;
  assign n249 = ~n247 & ~n248 ;
  assign n250 = ~n246 & n249 ;
  assign n251 = ~n243 & ~n250 ;
  assign n252 = ~n242 & n251 ;
  assign n253 = x54 & ~n125 ;
  assign n254 = x38 & n125 ;
  assign n255 = ~n253 & ~n254 ;
  assign n256 = x22 & ~n193 ;
  assign n257 = x6 & n193 ;
  assign n258 = ~n256 & ~n257 ;
  assign n259 = n255 & ~n258 ;
  assign n260 = n246 & ~n249 ;
  assign n261 = ~n259 & ~n260 ;
  assign n262 = ~n252 & n261 ;
  assign n263 = x23 & ~n193 ;
  assign n264 = x7 & n193 ;
  assign n265 = ~n263 & ~n264 ;
  assign n266 = x55 & ~n125 ;
  assign n267 = x39 & n125 ;
  assign n268 = ~n266 & ~n267 ;
  assign n269 = n265 & ~n268 ;
  assign n270 = ~n255 & n258 ;
  assign n271 = ~n269 & ~n270 ;
  assign n272 = ~n262 & n271 ;
  assign n273 = ~n265 & n268 ;
  assign n274 = x56 & ~n125 ;
  assign n275 = x40 & n125 ;
  assign n276 = ~n274 & ~n275 ;
  assign n277 = x24 & ~n193 ;
  assign n278 = x8 & n193 ;
  assign n279 = ~n277 & ~n278 ;
  assign n280 = n276 & ~n279 ;
  assign n281 = ~n273 & ~n280 ;
  assign n282 = ~n272 & n281 ;
  assign n283 = ~n276 & n279 ;
  assign n284 = x57 & ~n125 ;
  assign n285 = x41 & n125 ;
  assign n286 = ~n284 & ~n285 ;
  assign n287 = x25 & ~n193 ;
  assign n288 = x9 & n193 ;
  assign n289 = ~n287 & ~n288 ;
  assign n290 = ~n286 & n289 ;
  assign n291 = ~n283 & ~n290 ;
  assign n292 = ~n282 & n291 ;
  assign n293 = n286 & ~n289 ;
  assign n294 = x26 & ~n193 ;
  assign n295 = x10 & n193 ;
  assign n296 = ~n294 & ~n295 ;
  assign n297 = x58 & ~n125 ;
  assign n298 = x42 & n125 ;
  assign n299 = ~n297 & ~n298 ;
  assign n300 = ~n296 & n299 ;
  assign n301 = ~n293 & ~n300 ;
  assign n302 = ~n292 & n301 ;
  assign n303 = x27 & ~n193 ;
  assign n304 = x11 & n193 ;
  assign n305 = ~n303 & ~n304 ;
  assign n306 = x59 & ~n125 ;
  assign n307 = x43 & n125 ;
  assign n308 = ~n306 & ~n307 ;
  assign n309 = n305 & ~n308 ;
  assign n310 = n296 & ~n299 ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = ~n302 & n311 ;
  assign n313 = x60 & ~n125 ;
  assign n314 = x44 & n125 ;
  assign n315 = ~n313 & ~n314 ;
  assign n316 = x28 & ~n193 ;
  assign n317 = x12 & n193 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = n315 & ~n318 ;
  assign n320 = ~n305 & n308 ;
  assign n321 = ~n319 & ~n320 ;
  assign n322 = ~n312 & n321 ;
  assign n323 = ~n315 & n318 ;
  assign n324 = x61 & ~n125 ;
  assign n325 = x45 & n125 ;
  assign n326 = ~n324 & ~n325 ;
  assign n327 = x29 & ~n193 ;
  assign n328 = x13 & n193 ;
  assign n329 = ~n327 & ~n328 ;
  assign n330 = ~n326 & n329 ;
  assign n331 = ~n323 & ~n330 ;
  assign n332 = ~n322 & n331 ;
  assign n333 = n132 & ~n196 ;
  assign n334 = n326 & ~n329 ;
  assign n335 = ~n333 & ~n334 ;
  assign n336 = ~n332 & n335 ;
  assign n337 = ~n197 & ~n336 ;
  assign n338 = ~n129 & ~n337 ;
  assign n339 = ~n128 & ~n338 ;
  assign n340 = ~n125 & ~n339 ;
  assign n341 = ~n193 & n339 ;
  assign n342 = ~n340 & ~n341 ;
  assign n343 = ~n210 & n339 ;
  assign n344 = ~n207 & ~n339 ;
  assign n345 = ~n343 & ~n344 ;
  assign n346 = ~n203 & n339 ;
  assign n347 = ~n200 & ~n339 ;
  assign n348 = ~n346 & ~n347 ;
  assign n349 = ~n218 & n339 ;
  assign n350 = ~n215 & ~n339 ;
  assign n351 = ~n349 & ~n350 ;
  assign n352 = ~n228 & n339 ;
  assign n353 = ~n225 & ~n339 ;
  assign n354 = ~n352 & ~n353 ;
  assign n355 = ~n238 & n339 ;
  assign n356 = ~n235 & ~n339 ;
  assign n357 = ~n355 & ~n356 ;
  assign n358 = ~n249 & n339 ;
  assign n359 = ~n246 & ~n339 ;
  assign n360 = ~n358 & ~n359 ;
  assign n361 = ~n258 & n339 ;
  assign n362 = ~n255 & ~n339 ;
  assign n363 = ~n361 & ~n362 ;
  assign n364 = ~n265 & n339 ;
  assign n365 = ~n268 & ~n339 ;
  assign n366 = ~n364 & ~n365 ;
  assign n367 = ~n279 & n339 ;
  assign n368 = ~n276 & ~n339 ;
  assign n369 = ~n367 & ~n368 ;
  assign n370 = ~n289 & n339 ;
  assign n371 = ~n286 & ~n339 ;
  assign n372 = ~n370 & ~n371 ;
  assign n373 = ~n296 & n339 ;
  assign n374 = ~n299 & ~n339 ;
  assign n375 = ~n373 & ~n374 ;
  assign n376 = ~n305 & n339 ;
  assign n377 = ~n308 & ~n339 ;
  assign n378 = ~n376 & ~n377 ;
  assign n379 = ~n318 & n339 ;
  assign n380 = ~n315 & ~n339 ;
  assign n381 = ~n379 & ~n380 ;
  assign n382 = ~n329 & n339 ;
  assign n383 = ~n326 & ~n339 ;
  assign n384 = ~n382 & ~n383 ;
  assign n385 = ~n196 & n339 ;
  assign n386 = ~n132 & ~n339 ;
  assign n387 = ~n385 & ~n386 ;
  assign n388 = n126 & n127 ;
  assign y0 = ~n342 ;
  assign y1 = ~n339 ;
  assign y2 = ~n345 ;
  assign y3 = ~n348 ;
  assign y4 = ~n351 ;
  assign y5 = ~n354 ;
  assign y6 = ~n357 ;
  assign y7 = ~n360 ;
  assign y8 = ~n363 ;
  assign y9 = ~n366 ;
  assign y10 = ~n369 ;
  assign y11 = ~n372 ;
  assign y12 = ~n375 ;
  assign y13 = ~n378 ;
  assign y14 = ~n381 ;
  assign y15 = ~n384 ;
  assign y16 = ~n387 ;
  assign y17 = ~n388 ;
endmodule
