module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 ;
  assign n289 = ~x30 & ~x286 ;
  assign n290 = x30 & x286 ;
  assign n291 = ~n289 & ~n290 ;
  assign n292 = ~x29 & ~x285 ;
  assign n293 = x29 & x285 ;
  assign n294 = ~n292 & ~n293 ;
  assign n295 = n291 & n294 ;
  assign n296 = ~n291 & ~n294 ;
  assign n297 = ~n295 & ~n296 ;
  assign n298 = ~x31 & ~x287 ;
  assign n299 = x31 & x287 ;
  assign n300 = ~n298 & ~n299 ;
  assign n301 = ~n297 & ~n300 ;
  assign n302 = n297 & n300 ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = ~x25 & ~x281 ;
  assign n305 = x25 & x281 ;
  assign n306 = ~n304 & ~n305 ;
  assign n307 = ~n303 & ~n306 ;
  assign n308 = n303 & n306 ;
  assign n309 = ~n307 & ~n308 ;
  assign n310 = ~x27 & ~x283 ;
  assign n311 = x27 & x283 ;
  assign n312 = ~n310 & ~n311 ;
  assign n313 = ~x26 & ~x282 ;
  assign n314 = x26 & x282 ;
  assign n315 = ~n313 & ~n314 ;
  assign n316 = ~n312 & ~n315 ;
  assign n317 = n312 & n315 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = ~x28 & ~x284 ;
  assign n320 = x28 & x284 ;
  assign n321 = ~n319 & ~n320 ;
  assign n322 = ~n318 & ~n321 ;
  assign n323 = n318 & n321 ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = n309 & ~n324 ;
  assign n326 = ~n307 & ~n325 ;
  assign n327 = ~n295 & ~n302 ;
  assign n328 = ~n326 & n327 ;
  assign n329 = n326 & ~n327 ;
  assign n330 = ~n328 & ~n329 ;
  assign n331 = ~n317 & ~n323 ;
  assign n332 = n330 & n331 ;
  assign n333 = ~n328 & ~n332 ;
  assign n334 = ~n330 & ~n331 ;
  assign n335 = ~n332 & ~n334 ;
  assign n336 = ~n309 & n324 ;
  assign n337 = ~n325 & ~n336 ;
  assign n338 = ~x17 & ~x273 ;
  assign n339 = x17 & x273 ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = n337 & ~n340 ;
  assign n342 = ~x23 & ~x279 ;
  assign n343 = x23 & x279 ;
  assign n344 = ~n342 & ~n343 ;
  assign n345 = ~x22 & ~x278 ;
  assign n346 = x22 & x278 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = ~n344 & ~n347 ;
  assign n349 = n344 & n347 ;
  assign n350 = ~n348 & ~n349 ;
  assign n351 = ~x24 & ~x280 ;
  assign n352 = x24 & x280 ;
  assign n353 = ~n351 & ~n352 ;
  assign n354 = ~n350 & ~n353 ;
  assign n355 = n350 & n353 ;
  assign n356 = ~n354 & ~n355 ;
  assign n357 = ~x18 & ~x274 ;
  assign n358 = x18 & x274 ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = ~n356 & ~n359 ;
  assign n361 = n356 & n359 ;
  assign n362 = ~n360 & ~n361 ;
  assign n363 = ~x20 & ~x276 ;
  assign n364 = x20 & x276 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = ~x19 & ~x275 ;
  assign n367 = x19 & x275 ;
  assign n368 = ~n366 & ~n367 ;
  assign n369 = ~n365 & ~n368 ;
  assign n370 = n365 & n368 ;
  assign n371 = ~n369 & ~n370 ;
  assign n372 = ~x21 & ~x277 ;
  assign n373 = x21 & x277 ;
  assign n374 = ~n372 & ~n373 ;
  assign n375 = ~n371 & ~n374 ;
  assign n376 = n371 & n374 ;
  assign n377 = ~n375 & ~n376 ;
  assign n378 = n362 & ~n377 ;
  assign n379 = ~n362 & n377 ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = ~n337 & n340 ;
  assign n382 = ~n341 & ~n381 ;
  assign n383 = n380 & n382 ;
  assign n384 = ~n341 & ~n383 ;
  assign n385 = n335 & ~n384 ;
  assign n386 = ~n360 & ~n378 ;
  assign n387 = ~n349 & ~n355 ;
  assign n388 = ~n386 & n387 ;
  assign n389 = n386 & ~n387 ;
  assign n390 = ~n388 & ~n389 ;
  assign n391 = ~n370 & ~n376 ;
  assign n392 = n390 & n391 ;
  assign n393 = ~n390 & ~n391 ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = ~n335 & n384 ;
  assign n396 = ~n385 & ~n395 ;
  assign n397 = n394 & n396 ;
  assign n398 = ~n385 & ~n397 ;
  assign n399 = ~n333 & ~n398 ;
  assign n400 = n333 & n398 ;
  assign n401 = ~n399 & ~n400 ;
  assign n402 = ~n388 & ~n392 ;
  assign n403 = n401 & ~n402 ;
  assign n404 = ~n399 & ~n403 ;
  assign n405 = ~n401 & n402 ;
  assign n406 = ~n403 & ~n405 ;
  assign n407 = ~n394 & ~n396 ;
  assign n408 = ~n397 & ~n407 ;
  assign n409 = ~n380 & ~n382 ;
  assign n410 = ~n383 & ~n409 ;
  assign n411 = ~x1 & ~x257 ;
  assign n412 = x1 & x257 ;
  assign n413 = ~n411 & ~n412 ;
  assign n414 = n410 & ~n413 ;
  assign n415 = ~x8 & ~x264 ;
  assign n416 = x8 & x264 ;
  assign n417 = ~n415 & ~n416 ;
  assign n418 = ~x7 & ~x263 ;
  assign n419 = x7 & x263 ;
  assign n420 = ~n418 & ~n419 ;
  assign n421 = ~n417 & ~n420 ;
  assign n422 = n417 & n420 ;
  assign n423 = ~n421 & ~n422 ;
  assign n424 = ~x9 & ~x265 ;
  assign n425 = x9 & x265 ;
  assign n426 = ~n424 & ~n425 ;
  assign n427 = ~n423 & ~n426 ;
  assign n428 = n423 & n426 ;
  assign n429 = ~n427 & ~n428 ;
  assign n430 = ~x3 & ~x259 ;
  assign n431 = x3 & x259 ;
  assign n432 = ~n430 & ~n431 ;
  assign n433 = ~n429 & ~n432 ;
  assign n434 = n429 & n432 ;
  assign n435 = ~n433 & ~n434 ;
  assign n436 = ~x5 & ~x261 ;
  assign n437 = x5 & x261 ;
  assign n438 = ~n436 & ~n437 ;
  assign n439 = ~x4 & ~x260 ;
  assign n440 = x4 & x260 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = ~n438 & ~n441 ;
  assign n443 = n438 & n441 ;
  assign n444 = ~n442 & ~n443 ;
  assign n445 = ~x6 & ~x262 ;
  assign n446 = x6 & x262 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = ~n444 & ~n447 ;
  assign n449 = n444 & n447 ;
  assign n450 = ~n448 & ~n449 ;
  assign n451 = n435 & ~n450 ;
  assign n452 = ~n435 & n450 ;
  assign n453 = ~n451 & ~n452 ;
  assign n454 = ~x15 & ~x271 ;
  assign n455 = x15 & x271 ;
  assign n456 = ~n454 & ~n455 ;
  assign n457 = ~x14 & ~x270 ;
  assign n458 = x14 & x270 ;
  assign n459 = ~n457 & ~n458 ;
  assign n460 = ~n456 & ~n459 ;
  assign n461 = n456 & n459 ;
  assign n462 = ~n460 & ~n461 ;
  assign n463 = ~x16 & ~x272 ;
  assign n464 = x16 & x272 ;
  assign n465 = ~n463 & ~n464 ;
  assign n466 = ~n462 & ~n465 ;
  assign n467 = n462 & n465 ;
  assign n468 = ~n466 & ~n467 ;
  assign n469 = ~x10 & ~x266 ;
  assign n470 = x10 & x266 ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = ~n468 & ~n471 ;
  assign n473 = n468 & n471 ;
  assign n474 = ~n472 & ~n473 ;
  assign n475 = ~x12 & ~x268 ;
  assign n476 = x12 & x268 ;
  assign n477 = ~n475 & ~n476 ;
  assign n478 = ~x11 & ~x267 ;
  assign n479 = x11 & x267 ;
  assign n480 = ~n478 & ~n479 ;
  assign n481 = ~n477 & ~n480 ;
  assign n482 = n477 & n480 ;
  assign n483 = ~n481 & ~n482 ;
  assign n484 = ~x13 & ~x269 ;
  assign n485 = x13 & x269 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = ~n483 & ~n486 ;
  assign n488 = n483 & n486 ;
  assign n489 = ~n487 & ~n488 ;
  assign n490 = n474 & ~n489 ;
  assign n491 = ~n474 & n489 ;
  assign n492 = ~n490 & ~n491 ;
  assign n493 = ~x2 & ~x258 ;
  assign n494 = x2 & x258 ;
  assign n495 = ~n493 & ~n494 ;
  assign n496 = n492 & ~n495 ;
  assign n497 = ~n492 & n495 ;
  assign n498 = ~n496 & ~n497 ;
  assign n499 = n453 & n498 ;
  assign n500 = ~n453 & ~n498 ;
  assign n501 = ~n499 & ~n500 ;
  assign n502 = ~n410 & n413 ;
  assign n503 = ~n414 & ~n502 ;
  assign n504 = n501 & n503 ;
  assign n505 = ~n414 & ~n504 ;
  assign n506 = n408 & ~n505 ;
  assign n507 = ~n433 & ~n451 ;
  assign n508 = ~n422 & ~n428 ;
  assign n509 = ~n507 & n508 ;
  assign n510 = n507 & ~n508 ;
  assign n511 = ~n509 & ~n510 ;
  assign n512 = ~n443 & ~n449 ;
  assign n513 = n511 & n512 ;
  assign n514 = ~n511 & ~n512 ;
  assign n515 = ~n513 & ~n514 ;
  assign n516 = ~n472 & ~n490 ;
  assign n517 = ~n461 & ~n467 ;
  assign n518 = ~n516 & n517 ;
  assign n519 = n516 & ~n517 ;
  assign n520 = ~n518 & ~n519 ;
  assign n521 = ~n482 & ~n488 ;
  assign n522 = n520 & n521 ;
  assign n523 = ~n520 & ~n521 ;
  assign n524 = ~n522 & ~n523 ;
  assign n525 = ~n496 & ~n499 ;
  assign n526 = n524 & ~n525 ;
  assign n527 = ~n524 & n525 ;
  assign n528 = ~n526 & ~n527 ;
  assign n529 = n515 & n528 ;
  assign n530 = ~n515 & ~n528 ;
  assign n531 = ~n529 & ~n530 ;
  assign n532 = ~n408 & n505 ;
  assign n533 = ~n506 & ~n532 ;
  assign n534 = n531 & n533 ;
  assign n535 = ~n506 & ~n534 ;
  assign n536 = n406 & ~n535 ;
  assign n537 = ~n518 & ~n522 ;
  assign n538 = ~n526 & ~n529 ;
  assign n539 = ~n537 & ~n538 ;
  assign n540 = n537 & n538 ;
  assign n541 = ~n539 & ~n540 ;
  assign n542 = ~n509 & ~n513 ;
  assign n543 = n541 & ~n542 ;
  assign n544 = ~n541 & n542 ;
  assign n545 = ~n543 & ~n544 ;
  assign n546 = ~n406 & n535 ;
  assign n547 = ~n536 & ~n546 ;
  assign n548 = n545 & n547 ;
  assign n549 = ~n536 & ~n548 ;
  assign n550 = ~n404 & ~n549 ;
  assign n551 = n404 & n549 ;
  assign n552 = ~n550 & ~n551 ;
  assign n553 = ~n539 & ~n543 ;
  assign n554 = n552 & ~n553 ;
  assign n555 = ~n552 & n553 ;
  assign n556 = ~n554 & ~n555 ;
  assign n557 = ~n545 & ~n547 ;
  assign n558 = ~n548 & ~n557 ;
  assign n559 = ~n531 & ~n533 ;
  assign n560 = ~n534 & ~n559 ;
  assign n561 = ~n501 & ~n503 ;
  assign n562 = ~n504 & ~n561 ;
  assign n563 = ~x0 & ~x256 ;
  assign n564 = x0 & x256 ;
  assign n565 = ~n563 & ~n564 ;
  assign n566 = ~n562 & n565 ;
  assign n567 = ~n560 & n566 ;
  assign n568 = ~n558 & n567 ;
  assign n569 = ~n556 & n568 ;
  assign n570 = ~n550 & ~n554 ;
  assign n571 = n569 & n570 ;
  assign n572 = ~x47 & ~x271 ;
  assign n573 = x47 & x271 ;
  assign n574 = ~n572 & ~n573 ;
  assign n575 = ~x46 & ~x270 ;
  assign n576 = x46 & x270 ;
  assign n577 = ~n575 & ~n576 ;
  assign n578 = ~n574 & ~n577 ;
  assign n579 = n574 & n577 ;
  assign n580 = ~n578 & ~n579 ;
  assign n581 = ~x48 & ~x272 ;
  assign n582 = x48 & x272 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = ~n580 & ~n583 ;
  assign n585 = n580 & n583 ;
  assign n586 = ~n584 & ~n585 ;
  assign n587 = ~x42 & ~x266 ;
  assign n588 = x42 & x266 ;
  assign n589 = ~n587 & ~n588 ;
  assign n590 = ~n586 & ~n589 ;
  assign n591 = n586 & n589 ;
  assign n592 = ~n590 & ~n591 ;
  assign n593 = ~x44 & ~x268 ;
  assign n594 = x44 & x268 ;
  assign n595 = ~n593 & ~n594 ;
  assign n596 = ~x43 & ~x267 ;
  assign n597 = x43 & x267 ;
  assign n598 = ~n596 & ~n597 ;
  assign n599 = ~n595 & ~n598 ;
  assign n600 = n595 & n598 ;
  assign n601 = ~n599 & ~n600 ;
  assign n602 = ~x45 & ~x269 ;
  assign n603 = x45 & x269 ;
  assign n604 = ~n602 & ~n603 ;
  assign n605 = ~n601 & ~n604 ;
  assign n606 = n601 & n604 ;
  assign n607 = ~n605 & ~n606 ;
  assign n608 = n592 & ~n607 ;
  assign n609 = ~n590 & ~n608 ;
  assign n610 = ~n579 & ~n585 ;
  assign n611 = ~n609 & n610 ;
  assign n612 = n609 & ~n610 ;
  assign n613 = ~n611 & ~n612 ;
  assign n614 = ~n600 & ~n606 ;
  assign n615 = n613 & n614 ;
  assign n616 = ~n611 & ~n615 ;
  assign n617 = ~n613 & ~n614 ;
  assign n618 = ~n615 & ~n617 ;
  assign n619 = ~n592 & n607 ;
  assign n620 = ~n608 & ~n619 ;
  assign n621 = ~x34 & ~x258 ;
  assign n622 = x34 & x258 ;
  assign n623 = ~n621 & ~n622 ;
  assign n624 = n620 & ~n623 ;
  assign n625 = ~x40 & ~x264 ;
  assign n626 = x40 & x264 ;
  assign n627 = ~n625 & ~n626 ;
  assign n628 = ~x39 & ~x263 ;
  assign n629 = x39 & x263 ;
  assign n630 = ~n628 & ~n629 ;
  assign n631 = ~n627 & ~n630 ;
  assign n632 = n627 & n630 ;
  assign n633 = ~n631 & ~n632 ;
  assign n634 = ~x41 & ~x265 ;
  assign n635 = x41 & x265 ;
  assign n636 = ~n634 & ~n635 ;
  assign n637 = ~n633 & ~n636 ;
  assign n638 = n633 & n636 ;
  assign n639 = ~n637 & ~n638 ;
  assign n640 = ~x35 & ~x259 ;
  assign n641 = x35 & x259 ;
  assign n642 = ~n640 & ~n641 ;
  assign n643 = ~n639 & ~n642 ;
  assign n644 = n639 & n642 ;
  assign n645 = ~n643 & ~n644 ;
  assign n646 = ~x37 & ~x261 ;
  assign n647 = x37 & x261 ;
  assign n648 = ~n646 & ~n647 ;
  assign n649 = ~x36 & ~x260 ;
  assign n650 = x36 & x260 ;
  assign n651 = ~n649 & ~n650 ;
  assign n652 = ~n648 & ~n651 ;
  assign n653 = n648 & n651 ;
  assign n654 = ~n652 & ~n653 ;
  assign n655 = ~x38 & ~x262 ;
  assign n656 = x38 & x262 ;
  assign n657 = ~n655 & ~n656 ;
  assign n658 = ~n654 & ~n657 ;
  assign n659 = n654 & n657 ;
  assign n660 = ~n658 & ~n659 ;
  assign n661 = n645 & ~n660 ;
  assign n662 = ~n645 & n660 ;
  assign n663 = ~n661 & ~n662 ;
  assign n664 = ~n620 & n623 ;
  assign n665 = ~n624 & ~n664 ;
  assign n666 = n663 & n665 ;
  assign n667 = ~n624 & ~n666 ;
  assign n668 = n618 & ~n667 ;
  assign n669 = ~n643 & ~n661 ;
  assign n670 = ~n632 & ~n638 ;
  assign n671 = ~n669 & n670 ;
  assign n672 = n669 & ~n670 ;
  assign n673 = ~n671 & ~n672 ;
  assign n674 = ~n653 & ~n659 ;
  assign n675 = n673 & n674 ;
  assign n676 = ~n673 & ~n674 ;
  assign n677 = ~n675 & ~n676 ;
  assign n678 = ~n618 & n667 ;
  assign n679 = ~n668 & ~n678 ;
  assign n680 = n677 & n679 ;
  assign n681 = ~n668 & ~n680 ;
  assign n682 = ~n616 & ~n681 ;
  assign n683 = n616 & n681 ;
  assign n684 = ~n682 & ~n683 ;
  assign n685 = ~n671 & ~n675 ;
  assign n686 = n684 & ~n685 ;
  assign n687 = ~n684 & n685 ;
  assign n688 = ~n686 & ~n687 ;
  assign n689 = ~x62 & ~x286 ;
  assign n690 = x62 & x286 ;
  assign n691 = ~n689 & ~n690 ;
  assign n692 = ~x61 & ~x285 ;
  assign n693 = x61 & x285 ;
  assign n694 = ~n692 & ~n693 ;
  assign n695 = n691 & n694 ;
  assign n696 = ~n691 & ~n694 ;
  assign n697 = ~n695 & ~n696 ;
  assign n698 = ~x63 & ~x287 ;
  assign n699 = x63 & x287 ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = ~n697 & ~n700 ;
  assign n702 = n697 & n700 ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = ~x57 & ~x281 ;
  assign n705 = x57 & x281 ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = ~n703 & ~n706 ;
  assign n708 = n703 & n706 ;
  assign n709 = ~n707 & ~n708 ;
  assign n710 = ~x59 & ~x283 ;
  assign n711 = x59 & x283 ;
  assign n712 = ~n710 & ~n711 ;
  assign n713 = ~x58 & ~x282 ;
  assign n714 = x58 & x282 ;
  assign n715 = ~n713 & ~n714 ;
  assign n716 = ~n712 & ~n715 ;
  assign n717 = n712 & n715 ;
  assign n718 = ~n716 & ~n717 ;
  assign n719 = ~x60 & ~x284 ;
  assign n720 = x60 & x284 ;
  assign n721 = ~n719 & ~n720 ;
  assign n722 = ~n718 & ~n721 ;
  assign n723 = n718 & n721 ;
  assign n724 = ~n722 & ~n723 ;
  assign n725 = n709 & ~n724 ;
  assign n726 = ~n707 & ~n725 ;
  assign n727 = ~n695 & ~n702 ;
  assign n728 = ~n726 & n727 ;
  assign n729 = n726 & ~n727 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = ~n717 & ~n723 ;
  assign n732 = n730 & n731 ;
  assign n733 = ~n728 & ~n732 ;
  assign n734 = ~n730 & ~n731 ;
  assign n735 = ~n732 & ~n734 ;
  assign n736 = ~n709 & n724 ;
  assign n737 = ~n725 & ~n736 ;
  assign n738 = ~x49 & ~x273 ;
  assign n739 = x49 & x273 ;
  assign n740 = ~n738 & ~n739 ;
  assign n741 = n737 & ~n740 ;
  assign n742 = ~x55 & ~x279 ;
  assign n743 = x55 & x279 ;
  assign n744 = ~n742 & ~n743 ;
  assign n745 = ~x54 & ~x278 ;
  assign n746 = x54 & x278 ;
  assign n747 = ~n745 & ~n746 ;
  assign n748 = ~n744 & ~n747 ;
  assign n749 = n744 & n747 ;
  assign n750 = ~n748 & ~n749 ;
  assign n751 = ~x56 & ~x280 ;
  assign n752 = x56 & x280 ;
  assign n753 = ~n751 & ~n752 ;
  assign n754 = ~n750 & ~n753 ;
  assign n755 = n750 & n753 ;
  assign n756 = ~n754 & ~n755 ;
  assign n757 = ~x50 & ~x274 ;
  assign n758 = x50 & x274 ;
  assign n759 = ~n757 & ~n758 ;
  assign n760 = ~n756 & ~n759 ;
  assign n761 = n756 & n759 ;
  assign n762 = ~n760 & ~n761 ;
  assign n763 = ~x52 & ~x276 ;
  assign n764 = x52 & x276 ;
  assign n765 = ~n763 & ~n764 ;
  assign n766 = ~x51 & ~x275 ;
  assign n767 = x51 & x275 ;
  assign n768 = ~n766 & ~n767 ;
  assign n769 = ~n765 & ~n768 ;
  assign n770 = n765 & n768 ;
  assign n771 = ~n769 & ~n770 ;
  assign n772 = ~x53 & ~x277 ;
  assign n773 = x53 & x277 ;
  assign n774 = ~n772 & ~n773 ;
  assign n775 = ~n771 & ~n774 ;
  assign n776 = n771 & n774 ;
  assign n777 = ~n775 & ~n776 ;
  assign n778 = n762 & ~n777 ;
  assign n779 = ~n762 & n777 ;
  assign n780 = ~n778 & ~n779 ;
  assign n781 = ~n737 & n740 ;
  assign n782 = ~n741 & ~n781 ;
  assign n783 = n780 & n782 ;
  assign n784 = ~n741 & ~n783 ;
  assign n785 = n735 & ~n784 ;
  assign n786 = ~n760 & ~n778 ;
  assign n787 = ~n749 & ~n755 ;
  assign n788 = ~n786 & n787 ;
  assign n789 = n786 & ~n787 ;
  assign n790 = ~n788 & ~n789 ;
  assign n791 = ~n770 & ~n776 ;
  assign n792 = n790 & n791 ;
  assign n793 = ~n790 & ~n791 ;
  assign n794 = ~n792 & ~n793 ;
  assign n795 = ~n735 & n784 ;
  assign n796 = ~n785 & ~n795 ;
  assign n797 = n794 & n796 ;
  assign n798 = ~n785 & ~n797 ;
  assign n799 = ~n733 & ~n798 ;
  assign n800 = n733 & n798 ;
  assign n801 = ~n799 & ~n800 ;
  assign n802 = ~n788 & ~n792 ;
  assign n803 = n801 & ~n802 ;
  assign n804 = ~n801 & n802 ;
  assign n805 = ~n803 & ~n804 ;
  assign n806 = ~n794 & ~n796 ;
  assign n807 = ~n797 & ~n806 ;
  assign n808 = ~n780 & ~n782 ;
  assign n809 = ~n783 & ~n808 ;
  assign n810 = ~x33 & ~x257 ;
  assign n811 = x33 & x257 ;
  assign n812 = ~n810 & ~n811 ;
  assign n813 = n809 & ~n812 ;
  assign n814 = ~n663 & ~n665 ;
  assign n815 = ~n666 & ~n814 ;
  assign n816 = ~n809 & n812 ;
  assign n817 = ~n813 & ~n816 ;
  assign n818 = n815 & n817 ;
  assign n819 = ~n813 & ~n818 ;
  assign n820 = n807 & ~n819 ;
  assign n821 = ~n677 & ~n679 ;
  assign n822 = ~n680 & ~n821 ;
  assign n823 = ~n807 & n819 ;
  assign n824 = ~n820 & ~n823 ;
  assign n825 = n822 & n824 ;
  assign n826 = ~n820 & ~n825 ;
  assign n827 = n805 & ~n826 ;
  assign n828 = ~n805 & n826 ;
  assign n829 = ~n827 & ~n828 ;
  assign n830 = n688 & n829 ;
  assign n831 = ~n688 & ~n829 ;
  assign n832 = ~n830 & ~n831 ;
  assign n833 = ~n822 & ~n824 ;
  assign n834 = ~n825 & ~n833 ;
  assign n835 = ~n815 & ~n817 ;
  assign n836 = ~n818 & ~n835 ;
  assign n837 = ~x32 & ~x256 ;
  assign n838 = x32 & x256 ;
  assign n839 = ~n837 & ~n838 ;
  assign n840 = ~n836 & n839 ;
  assign n841 = ~n834 & n840 ;
  assign n842 = ~n832 & n841 ;
  assign n843 = ~n799 & ~n803 ;
  assign n844 = ~n827 & ~n830 ;
  assign n845 = ~n843 & ~n844 ;
  assign n846 = n843 & n844 ;
  assign n847 = ~n845 & ~n846 ;
  assign n848 = ~n682 & ~n686 ;
  assign n849 = n847 & ~n848 ;
  assign n850 = ~n847 & n848 ;
  assign n851 = ~n849 & ~n850 ;
  assign n852 = n842 & ~n851 ;
  assign n853 = ~n845 & ~n849 ;
  assign n854 = n852 & n853 ;
  assign n855 = ~x79 & ~x271 ;
  assign n856 = x79 & x271 ;
  assign n857 = ~n855 & ~n856 ;
  assign n858 = ~x78 & ~x270 ;
  assign n859 = x78 & x270 ;
  assign n860 = ~n858 & ~n859 ;
  assign n861 = ~n857 & ~n860 ;
  assign n862 = n857 & n860 ;
  assign n863 = ~n861 & ~n862 ;
  assign n864 = ~x80 & ~x272 ;
  assign n865 = x80 & x272 ;
  assign n866 = ~n864 & ~n865 ;
  assign n867 = ~n863 & ~n866 ;
  assign n868 = n863 & n866 ;
  assign n869 = ~n867 & ~n868 ;
  assign n870 = ~x74 & ~x266 ;
  assign n871 = x74 & x266 ;
  assign n872 = ~n870 & ~n871 ;
  assign n873 = ~n869 & ~n872 ;
  assign n874 = n869 & n872 ;
  assign n875 = ~n873 & ~n874 ;
  assign n876 = ~x76 & ~x268 ;
  assign n877 = x76 & x268 ;
  assign n878 = ~n876 & ~n877 ;
  assign n879 = ~x75 & ~x267 ;
  assign n880 = x75 & x267 ;
  assign n881 = ~n879 & ~n880 ;
  assign n882 = ~n878 & ~n881 ;
  assign n883 = n878 & n881 ;
  assign n884 = ~n882 & ~n883 ;
  assign n885 = ~x77 & ~x269 ;
  assign n886 = x77 & x269 ;
  assign n887 = ~n885 & ~n886 ;
  assign n888 = ~n884 & ~n887 ;
  assign n889 = n884 & n887 ;
  assign n890 = ~n888 & ~n889 ;
  assign n891 = n875 & ~n890 ;
  assign n892 = ~n873 & ~n891 ;
  assign n893 = ~n862 & ~n868 ;
  assign n894 = ~n892 & n893 ;
  assign n895 = n892 & ~n893 ;
  assign n896 = ~n894 & ~n895 ;
  assign n897 = ~n883 & ~n889 ;
  assign n898 = n896 & n897 ;
  assign n899 = ~n894 & ~n898 ;
  assign n900 = ~n896 & ~n897 ;
  assign n901 = ~n898 & ~n900 ;
  assign n902 = ~n875 & n890 ;
  assign n903 = ~n891 & ~n902 ;
  assign n904 = ~x66 & ~x258 ;
  assign n905 = x66 & x258 ;
  assign n906 = ~n904 & ~n905 ;
  assign n907 = n903 & ~n906 ;
  assign n908 = ~x72 & ~x264 ;
  assign n909 = x72 & x264 ;
  assign n910 = ~n908 & ~n909 ;
  assign n911 = ~x71 & ~x263 ;
  assign n912 = x71 & x263 ;
  assign n913 = ~n911 & ~n912 ;
  assign n914 = ~n910 & ~n913 ;
  assign n915 = n910 & n913 ;
  assign n916 = ~n914 & ~n915 ;
  assign n917 = ~x73 & ~x265 ;
  assign n918 = x73 & x265 ;
  assign n919 = ~n917 & ~n918 ;
  assign n920 = ~n916 & ~n919 ;
  assign n921 = n916 & n919 ;
  assign n922 = ~n920 & ~n921 ;
  assign n923 = ~x67 & ~x259 ;
  assign n924 = x67 & x259 ;
  assign n925 = ~n923 & ~n924 ;
  assign n926 = ~n922 & ~n925 ;
  assign n927 = n922 & n925 ;
  assign n928 = ~n926 & ~n927 ;
  assign n929 = ~x69 & ~x261 ;
  assign n930 = x69 & x261 ;
  assign n931 = ~n929 & ~n930 ;
  assign n932 = ~x68 & ~x260 ;
  assign n933 = x68 & x260 ;
  assign n934 = ~n932 & ~n933 ;
  assign n935 = ~n931 & ~n934 ;
  assign n936 = n931 & n934 ;
  assign n937 = ~n935 & ~n936 ;
  assign n938 = ~x70 & ~x262 ;
  assign n939 = x70 & x262 ;
  assign n940 = ~n938 & ~n939 ;
  assign n941 = ~n937 & ~n940 ;
  assign n942 = n937 & n940 ;
  assign n943 = ~n941 & ~n942 ;
  assign n944 = n928 & ~n943 ;
  assign n945 = ~n928 & n943 ;
  assign n946 = ~n944 & ~n945 ;
  assign n947 = ~n903 & n906 ;
  assign n948 = ~n907 & ~n947 ;
  assign n949 = n946 & n948 ;
  assign n950 = ~n907 & ~n949 ;
  assign n951 = n901 & ~n950 ;
  assign n952 = ~n926 & ~n944 ;
  assign n953 = ~n915 & ~n921 ;
  assign n954 = ~n952 & n953 ;
  assign n955 = n952 & ~n953 ;
  assign n956 = ~n954 & ~n955 ;
  assign n957 = ~n936 & ~n942 ;
  assign n958 = n956 & n957 ;
  assign n959 = ~n956 & ~n957 ;
  assign n960 = ~n958 & ~n959 ;
  assign n961 = ~n901 & n950 ;
  assign n962 = ~n951 & ~n961 ;
  assign n963 = n960 & n962 ;
  assign n964 = ~n951 & ~n963 ;
  assign n965 = ~n899 & ~n964 ;
  assign n966 = n899 & n964 ;
  assign n967 = ~n965 & ~n966 ;
  assign n968 = ~n954 & ~n958 ;
  assign n969 = n967 & ~n968 ;
  assign n970 = ~n967 & n968 ;
  assign n971 = ~n969 & ~n970 ;
  assign n972 = ~x94 & ~x286 ;
  assign n973 = x94 & x286 ;
  assign n974 = ~n972 & ~n973 ;
  assign n975 = ~x93 & ~x285 ;
  assign n976 = x93 & x285 ;
  assign n977 = ~n975 & ~n976 ;
  assign n978 = n974 & n977 ;
  assign n979 = ~n974 & ~n977 ;
  assign n980 = ~n978 & ~n979 ;
  assign n981 = ~x95 & ~x287 ;
  assign n982 = x95 & x287 ;
  assign n983 = ~n981 & ~n982 ;
  assign n984 = ~n980 & ~n983 ;
  assign n985 = n980 & n983 ;
  assign n986 = ~n984 & ~n985 ;
  assign n987 = ~x89 & ~x281 ;
  assign n988 = x89 & x281 ;
  assign n989 = ~n987 & ~n988 ;
  assign n990 = ~n986 & ~n989 ;
  assign n991 = n986 & n989 ;
  assign n992 = ~n990 & ~n991 ;
  assign n993 = ~x91 & ~x283 ;
  assign n994 = x91 & x283 ;
  assign n995 = ~n993 & ~n994 ;
  assign n996 = ~x90 & ~x282 ;
  assign n997 = x90 & x282 ;
  assign n998 = ~n996 & ~n997 ;
  assign n999 = ~n995 & ~n998 ;
  assign n1000 = n995 & n998 ;
  assign n1001 = ~n999 & ~n1000 ;
  assign n1002 = ~x92 & ~x284 ;
  assign n1003 = x92 & x284 ;
  assign n1004 = ~n1002 & ~n1003 ;
  assign n1005 = ~n1001 & ~n1004 ;
  assign n1006 = n1001 & n1004 ;
  assign n1007 = ~n1005 & ~n1006 ;
  assign n1008 = n992 & ~n1007 ;
  assign n1009 = ~n990 & ~n1008 ;
  assign n1010 = ~n978 & ~n985 ;
  assign n1011 = ~n1009 & n1010 ;
  assign n1012 = n1009 & ~n1010 ;
  assign n1013 = ~n1011 & ~n1012 ;
  assign n1014 = ~n1000 & ~n1006 ;
  assign n1015 = n1013 & n1014 ;
  assign n1016 = ~n1011 & ~n1015 ;
  assign n1017 = ~n1013 & ~n1014 ;
  assign n1018 = ~n1015 & ~n1017 ;
  assign n1019 = ~n992 & n1007 ;
  assign n1020 = ~n1008 & ~n1019 ;
  assign n1021 = ~x81 & ~x273 ;
  assign n1022 = x81 & x273 ;
  assign n1023 = ~n1021 & ~n1022 ;
  assign n1024 = n1020 & ~n1023 ;
  assign n1025 = ~x87 & ~x279 ;
  assign n1026 = x87 & x279 ;
  assign n1027 = ~n1025 & ~n1026 ;
  assign n1028 = ~x86 & ~x278 ;
  assign n1029 = x86 & x278 ;
  assign n1030 = ~n1028 & ~n1029 ;
  assign n1031 = ~n1027 & ~n1030 ;
  assign n1032 = n1027 & n1030 ;
  assign n1033 = ~n1031 & ~n1032 ;
  assign n1034 = ~x88 & ~x280 ;
  assign n1035 = x88 & x280 ;
  assign n1036 = ~n1034 & ~n1035 ;
  assign n1037 = ~n1033 & ~n1036 ;
  assign n1038 = n1033 & n1036 ;
  assign n1039 = ~n1037 & ~n1038 ;
  assign n1040 = ~x82 & ~x274 ;
  assign n1041 = x82 & x274 ;
  assign n1042 = ~n1040 & ~n1041 ;
  assign n1043 = ~n1039 & ~n1042 ;
  assign n1044 = n1039 & n1042 ;
  assign n1045 = ~n1043 & ~n1044 ;
  assign n1046 = ~x84 & ~x276 ;
  assign n1047 = x84 & x276 ;
  assign n1048 = ~n1046 & ~n1047 ;
  assign n1049 = ~x83 & ~x275 ;
  assign n1050 = x83 & x275 ;
  assign n1051 = ~n1049 & ~n1050 ;
  assign n1052 = ~n1048 & ~n1051 ;
  assign n1053 = n1048 & n1051 ;
  assign n1054 = ~n1052 & ~n1053 ;
  assign n1055 = ~x85 & ~x277 ;
  assign n1056 = x85 & x277 ;
  assign n1057 = ~n1055 & ~n1056 ;
  assign n1058 = ~n1054 & ~n1057 ;
  assign n1059 = n1054 & n1057 ;
  assign n1060 = ~n1058 & ~n1059 ;
  assign n1061 = n1045 & ~n1060 ;
  assign n1062 = ~n1045 & n1060 ;
  assign n1063 = ~n1061 & ~n1062 ;
  assign n1064 = ~n1020 & n1023 ;
  assign n1065 = ~n1024 & ~n1064 ;
  assign n1066 = n1063 & n1065 ;
  assign n1067 = ~n1024 & ~n1066 ;
  assign n1068 = n1018 & ~n1067 ;
  assign n1069 = ~n1043 & ~n1061 ;
  assign n1070 = ~n1032 & ~n1038 ;
  assign n1071 = ~n1069 & n1070 ;
  assign n1072 = n1069 & ~n1070 ;
  assign n1073 = ~n1071 & ~n1072 ;
  assign n1074 = ~n1053 & ~n1059 ;
  assign n1075 = n1073 & n1074 ;
  assign n1076 = ~n1073 & ~n1074 ;
  assign n1077 = ~n1075 & ~n1076 ;
  assign n1078 = ~n1018 & n1067 ;
  assign n1079 = ~n1068 & ~n1078 ;
  assign n1080 = n1077 & n1079 ;
  assign n1081 = ~n1068 & ~n1080 ;
  assign n1082 = ~n1016 & ~n1081 ;
  assign n1083 = n1016 & n1081 ;
  assign n1084 = ~n1082 & ~n1083 ;
  assign n1085 = ~n1071 & ~n1075 ;
  assign n1086 = n1084 & ~n1085 ;
  assign n1087 = ~n1084 & n1085 ;
  assign n1088 = ~n1086 & ~n1087 ;
  assign n1089 = ~n1077 & ~n1079 ;
  assign n1090 = ~n1080 & ~n1089 ;
  assign n1091 = ~n1063 & ~n1065 ;
  assign n1092 = ~n1066 & ~n1091 ;
  assign n1093 = ~x65 & ~x257 ;
  assign n1094 = x65 & x257 ;
  assign n1095 = ~n1093 & ~n1094 ;
  assign n1096 = n1092 & ~n1095 ;
  assign n1097 = ~n946 & ~n948 ;
  assign n1098 = ~n949 & ~n1097 ;
  assign n1099 = ~n1092 & n1095 ;
  assign n1100 = ~n1096 & ~n1099 ;
  assign n1101 = n1098 & n1100 ;
  assign n1102 = ~n1096 & ~n1101 ;
  assign n1103 = n1090 & ~n1102 ;
  assign n1104 = ~n960 & ~n962 ;
  assign n1105 = ~n963 & ~n1104 ;
  assign n1106 = ~n1090 & n1102 ;
  assign n1107 = ~n1103 & ~n1106 ;
  assign n1108 = n1105 & n1107 ;
  assign n1109 = ~n1103 & ~n1108 ;
  assign n1110 = n1088 & ~n1109 ;
  assign n1111 = ~n1088 & n1109 ;
  assign n1112 = ~n1110 & ~n1111 ;
  assign n1113 = n971 & n1112 ;
  assign n1114 = ~n971 & ~n1112 ;
  assign n1115 = ~n1113 & ~n1114 ;
  assign n1116 = ~n1105 & ~n1107 ;
  assign n1117 = ~n1108 & ~n1116 ;
  assign n1118 = ~n1098 & ~n1100 ;
  assign n1119 = ~n1101 & ~n1118 ;
  assign n1120 = ~x64 & ~x256 ;
  assign n1121 = x64 & x256 ;
  assign n1122 = ~n1120 & ~n1121 ;
  assign n1123 = ~n1119 & n1122 ;
  assign n1124 = ~n1117 & n1123 ;
  assign n1125 = ~n1115 & n1124 ;
  assign n1126 = ~n1082 & ~n1086 ;
  assign n1127 = ~n1110 & ~n1113 ;
  assign n1128 = ~n1126 & ~n1127 ;
  assign n1129 = n1126 & n1127 ;
  assign n1130 = ~n1128 & ~n1129 ;
  assign n1131 = ~n965 & ~n969 ;
  assign n1132 = n1130 & ~n1131 ;
  assign n1133 = ~n1130 & n1131 ;
  assign n1134 = ~n1132 & ~n1133 ;
  assign n1135 = n1125 & ~n1134 ;
  assign n1136 = ~n1128 & ~n1132 ;
  assign n1137 = n1135 & n1136 ;
  assign n1138 = ~x111 & ~x271 ;
  assign n1139 = x111 & x271 ;
  assign n1140 = ~n1138 & ~n1139 ;
  assign n1141 = ~x110 & ~x270 ;
  assign n1142 = x110 & x270 ;
  assign n1143 = ~n1141 & ~n1142 ;
  assign n1144 = ~n1140 & ~n1143 ;
  assign n1145 = n1140 & n1143 ;
  assign n1146 = ~n1144 & ~n1145 ;
  assign n1147 = ~x112 & ~x272 ;
  assign n1148 = x112 & x272 ;
  assign n1149 = ~n1147 & ~n1148 ;
  assign n1150 = ~n1146 & ~n1149 ;
  assign n1151 = n1146 & n1149 ;
  assign n1152 = ~n1150 & ~n1151 ;
  assign n1153 = ~x106 & ~x266 ;
  assign n1154 = x106 & x266 ;
  assign n1155 = ~n1153 & ~n1154 ;
  assign n1156 = ~n1152 & ~n1155 ;
  assign n1157 = n1152 & n1155 ;
  assign n1158 = ~n1156 & ~n1157 ;
  assign n1159 = ~x108 & ~x268 ;
  assign n1160 = x108 & x268 ;
  assign n1161 = ~n1159 & ~n1160 ;
  assign n1162 = ~x107 & ~x267 ;
  assign n1163 = x107 & x267 ;
  assign n1164 = ~n1162 & ~n1163 ;
  assign n1165 = ~n1161 & ~n1164 ;
  assign n1166 = n1161 & n1164 ;
  assign n1167 = ~n1165 & ~n1166 ;
  assign n1168 = ~x109 & ~x269 ;
  assign n1169 = x109 & x269 ;
  assign n1170 = ~n1168 & ~n1169 ;
  assign n1171 = ~n1167 & ~n1170 ;
  assign n1172 = n1167 & n1170 ;
  assign n1173 = ~n1171 & ~n1172 ;
  assign n1174 = n1158 & ~n1173 ;
  assign n1175 = ~n1156 & ~n1174 ;
  assign n1176 = ~n1145 & ~n1151 ;
  assign n1177 = ~n1175 & n1176 ;
  assign n1178 = n1175 & ~n1176 ;
  assign n1179 = ~n1177 & ~n1178 ;
  assign n1180 = ~n1166 & ~n1172 ;
  assign n1181 = n1179 & n1180 ;
  assign n1182 = ~n1177 & ~n1181 ;
  assign n1183 = ~n1179 & ~n1180 ;
  assign n1184 = ~n1181 & ~n1183 ;
  assign n1185 = ~n1158 & n1173 ;
  assign n1186 = ~n1174 & ~n1185 ;
  assign n1187 = ~x98 & ~x258 ;
  assign n1188 = x98 & x258 ;
  assign n1189 = ~n1187 & ~n1188 ;
  assign n1190 = n1186 & ~n1189 ;
  assign n1191 = ~x104 & ~x264 ;
  assign n1192 = x104 & x264 ;
  assign n1193 = ~n1191 & ~n1192 ;
  assign n1194 = ~x103 & ~x263 ;
  assign n1195 = x103 & x263 ;
  assign n1196 = ~n1194 & ~n1195 ;
  assign n1197 = ~n1193 & ~n1196 ;
  assign n1198 = n1193 & n1196 ;
  assign n1199 = ~n1197 & ~n1198 ;
  assign n1200 = ~x105 & ~x265 ;
  assign n1201 = x105 & x265 ;
  assign n1202 = ~n1200 & ~n1201 ;
  assign n1203 = ~n1199 & ~n1202 ;
  assign n1204 = n1199 & n1202 ;
  assign n1205 = ~n1203 & ~n1204 ;
  assign n1206 = ~x99 & ~x259 ;
  assign n1207 = x99 & x259 ;
  assign n1208 = ~n1206 & ~n1207 ;
  assign n1209 = ~n1205 & ~n1208 ;
  assign n1210 = n1205 & n1208 ;
  assign n1211 = ~n1209 & ~n1210 ;
  assign n1212 = ~x101 & ~x261 ;
  assign n1213 = x101 & x261 ;
  assign n1214 = ~n1212 & ~n1213 ;
  assign n1215 = ~x100 & ~x260 ;
  assign n1216 = x100 & x260 ;
  assign n1217 = ~n1215 & ~n1216 ;
  assign n1218 = ~n1214 & ~n1217 ;
  assign n1219 = n1214 & n1217 ;
  assign n1220 = ~n1218 & ~n1219 ;
  assign n1221 = ~x102 & ~x262 ;
  assign n1222 = x102 & x262 ;
  assign n1223 = ~n1221 & ~n1222 ;
  assign n1224 = ~n1220 & ~n1223 ;
  assign n1225 = n1220 & n1223 ;
  assign n1226 = ~n1224 & ~n1225 ;
  assign n1227 = n1211 & ~n1226 ;
  assign n1228 = ~n1211 & n1226 ;
  assign n1229 = ~n1227 & ~n1228 ;
  assign n1230 = ~n1186 & n1189 ;
  assign n1231 = ~n1190 & ~n1230 ;
  assign n1232 = n1229 & n1231 ;
  assign n1233 = ~n1190 & ~n1232 ;
  assign n1234 = n1184 & ~n1233 ;
  assign n1235 = ~n1209 & ~n1227 ;
  assign n1236 = ~n1198 & ~n1204 ;
  assign n1237 = ~n1235 & n1236 ;
  assign n1238 = n1235 & ~n1236 ;
  assign n1239 = ~n1237 & ~n1238 ;
  assign n1240 = ~n1219 & ~n1225 ;
  assign n1241 = n1239 & n1240 ;
  assign n1242 = ~n1239 & ~n1240 ;
  assign n1243 = ~n1241 & ~n1242 ;
  assign n1244 = ~n1184 & n1233 ;
  assign n1245 = ~n1234 & ~n1244 ;
  assign n1246 = n1243 & n1245 ;
  assign n1247 = ~n1234 & ~n1246 ;
  assign n1248 = ~n1182 & ~n1247 ;
  assign n1249 = n1182 & n1247 ;
  assign n1250 = ~n1248 & ~n1249 ;
  assign n1251 = ~n1237 & ~n1241 ;
  assign n1252 = n1250 & ~n1251 ;
  assign n1253 = ~n1250 & n1251 ;
  assign n1254 = ~n1252 & ~n1253 ;
  assign n1255 = ~x126 & ~x286 ;
  assign n1256 = x126 & x286 ;
  assign n1257 = ~n1255 & ~n1256 ;
  assign n1258 = ~x125 & ~x285 ;
  assign n1259 = x125 & x285 ;
  assign n1260 = ~n1258 & ~n1259 ;
  assign n1261 = n1257 & n1260 ;
  assign n1262 = ~n1257 & ~n1260 ;
  assign n1263 = ~n1261 & ~n1262 ;
  assign n1264 = ~x127 & ~x287 ;
  assign n1265 = x127 & x287 ;
  assign n1266 = ~n1264 & ~n1265 ;
  assign n1267 = ~n1263 & ~n1266 ;
  assign n1268 = n1263 & n1266 ;
  assign n1269 = ~n1267 & ~n1268 ;
  assign n1270 = ~x121 & ~x281 ;
  assign n1271 = x121 & x281 ;
  assign n1272 = ~n1270 & ~n1271 ;
  assign n1273 = ~n1269 & ~n1272 ;
  assign n1274 = n1269 & n1272 ;
  assign n1275 = ~n1273 & ~n1274 ;
  assign n1276 = ~x123 & ~x283 ;
  assign n1277 = x123 & x283 ;
  assign n1278 = ~n1276 & ~n1277 ;
  assign n1279 = ~x122 & ~x282 ;
  assign n1280 = x122 & x282 ;
  assign n1281 = ~n1279 & ~n1280 ;
  assign n1282 = ~n1278 & ~n1281 ;
  assign n1283 = n1278 & n1281 ;
  assign n1284 = ~n1282 & ~n1283 ;
  assign n1285 = ~x124 & ~x284 ;
  assign n1286 = x124 & x284 ;
  assign n1287 = ~n1285 & ~n1286 ;
  assign n1288 = ~n1284 & ~n1287 ;
  assign n1289 = n1284 & n1287 ;
  assign n1290 = ~n1288 & ~n1289 ;
  assign n1291 = n1275 & ~n1290 ;
  assign n1292 = ~n1273 & ~n1291 ;
  assign n1293 = ~n1261 & ~n1268 ;
  assign n1294 = ~n1292 & n1293 ;
  assign n1295 = n1292 & ~n1293 ;
  assign n1296 = ~n1294 & ~n1295 ;
  assign n1297 = ~n1283 & ~n1289 ;
  assign n1298 = n1296 & n1297 ;
  assign n1299 = ~n1294 & ~n1298 ;
  assign n1300 = ~n1296 & ~n1297 ;
  assign n1301 = ~n1298 & ~n1300 ;
  assign n1302 = ~n1275 & n1290 ;
  assign n1303 = ~n1291 & ~n1302 ;
  assign n1304 = ~x113 & ~x273 ;
  assign n1305 = x113 & x273 ;
  assign n1306 = ~n1304 & ~n1305 ;
  assign n1307 = n1303 & ~n1306 ;
  assign n1308 = ~x119 & ~x279 ;
  assign n1309 = x119 & x279 ;
  assign n1310 = ~n1308 & ~n1309 ;
  assign n1311 = ~x118 & ~x278 ;
  assign n1312 = x118 & x278 ;
  assign n1313 = ~n1311 & ~n1312 ;
  assign n1314 = ~n1310 & ~n1313 ;
  assign n1315 = n1310 & n1313 ;
  assign n1316 = ~n1314 & ~n1315 ;
  assign n1317 = ~x120 & ~x280 ;
  assign n1318 = x120 & x280 ;
  assign n1319 = ~n1317 & ~n1318 ;
  assign n1320 = ~n1316 & ~n1319 ;
  assign n1321 = n1316 & n1319 ;
  assign n1322 = ~n1320 & ~n1321 ;
  assign n1323 = ~x114 & ~x274 ;
  assign n1324 = x114 & x274 ;
  assign n1325 = ~n1323 & ~n1324 ;
  assign n1326 = ~n1322 & ~n1325 ;
  assign n1327 = n1322 & n1325 ;
  assign n1328 = ~n1326 & ~n1327 ;
  assign n1329 = ~x116 & ~x276 ;
  assign n1330 = x116 & x276 ;
  assign n1331 = ~n1329 & ~n1330 ;
  assign n1332 = ~x115 & ~x275 ;
  assign n1333 = x115 & x275 ;
  assign n1334 = ~n1332 & ~n1333 ;
  assign n1335 = ~n1331 & ~n1334 ;
  assign n1336 = n1331 & n1334 ;
  assign n1337 = ~n1335 & ~n1336 ;
  assign n1338 = ~x117 & ~x277 ;
  assign n1339 = x117 & x277 ;
  assign n1340 = ~n1338 & ~n1339 ;
  assign n1341 = ~n1337 & ~n1340 ;
  assign n1342 = n1337 & n1340 ;
  assign n1343 = ~n1341 & ~n1342 ;
  assign n1344 = n1328 & ~n1343 ;
  assign n1345 = ~n1328 & n1343 ;
  assign n1346 = ~n1344 & ~n1345 ;
  assign n1347 = ~n1303 & n1306 ;
  assign n1348 = ~n1307 & ~n1347 ;
  assign n1349 = n1346 & n1348 ;
  assign n1350 = ~n1307 & ~n1349 ;
  assign n1351 = n1301 & ~n1350 ;
  assign n1352 = ~n1326 & ~n1344 ;
  assign n1353 = ~n1315 & ~n1321 ;
  assign n1354 = ~n1352 & n1353 ;
  assign n1355 = n1352 & ~n1353 ;
  assign n1356 = ~n1354 & ~n1355 ;
  assign n1357 = ~n1336 & ~n1342 ;
  assign n1358 = n1356 & n1357 ;
  assign n1359 = ~n1356 & ~n1357 ;
  assign n1360 = ~n1358 & ~n1359 ;
  assign n1361 = ~n1301 & n1350 ;
  assign n1362 = ~n1351 & ~n1361 ;
  assign n1363 = n1360 & n1362 ;
  assign n1364 = ~n1351 & ~n1363 ;
  assign n1365 = ~n1299 & ~n1364 ;
  assign n1366 = n1299 & n1364 ;
  assign n1367 = ~n1365 & ~n1366 ;
  assign n1368 = ~n1354 & ~n1358 ;
  assign n1369 = n1367 & ~n1368 ;
  assign n1370 = ~n1367 & n1368 ;
  assign n1371 = ~n1369 & ~n1370 ;
  assign n1372 = ~n1360 & ~n1362 ;
  assign n1373 = ~n1363 & ~n1372 ;
  assign n1374 = ~n1346 & ~n1348 ;
  assign n1375 = ~n1349 & ~n1374 ;
  assign n1376 = ~x97 & ~x257 ;
  assign n1377 = x97 & x257 ;
  assign n1378 = ~n1376 & ~n1377 ;
  assign n1379 = n1375 & ~n1378 ;
  assign n1380 = ~n1229 & ~n1231 ;
  assign n1381 = ~n1232 & ~n1380 ;
  assign n1382 = ~n1375 & n1378 ;
  assign n1383 = ~n1379 & ~n1382 ;
  assign n1384 = n1381 & n1383 ;
  assign n1385 = ~n1379 & ~n1384 ;
  assign n1386 = n1373 & ~n1385 ;
  assign n1387 = ~n1243 & ~n1245 ;
  assign n1388 = ~n1246 & ~n1387 ;
  assign n1389 = ~n1373 & n1385 ;
  assign n1390 = ~n1386 & ~n1389 ;
  assign n1391 = n1388 & n1390 ;
  assign n1392 = ~n1386 & ~n1391 ;
  assign n1393 = n1371 & ~n1392 ;
  assign n1394 = ~n1371 & n1392 ;
  assign n1395 = ~n1393 & ~n1394 ;
  assign n1396 = n1254 & n1395 ;
  assign n1397 = ~n1254 & ~n1395 ;
  assign n1398 = ~n1396 & ~n1397 ;
  assign n1399 = ~n1388 & ~n1390 ;
  assign n1400 = ~n1391 & ~n1399 ;
  assign n1401 = ~n1381 & ~n1383 ;
  assign n1402 = ~n1384 & ~n1401 ;
  assign n1403 = ~x96 & ~x256 ;
  assign n1404 = x96 & x256 ;
  assign n1405 = ~n1403 & ~n1404 ;
  assign n1406 = ~n1402 & n1405 ;
  assign n1407 = ~n1400 & n1406 ;
  assign n1408 = ~n1398 & n1407 ;
  assign n1409 = ~n1365 & ~n1369 ;
  assign n1410 = ~n1393 & ~n1396 ;
  assign n1411 = ~n1409 & ~n1410 ;
  assign n1412 = n1409 & n1410 ;
  assign n1413 = ~n1411 & ~n1412 ;
  assign n1414 = ~n1248 & ~n1252 ;
  assign n1415 = n1413 & ~n1414 ;
  assign n1416 = ~n1413 & n1414 ;
  assign n1417 = ~n1415 & ~n1416 ;
  assign n1418 = n1408 & ~n1417 ;
  assign n1419 = ~n1411 & ~n1415 ;
  assign n1420 = n1418 & n1419 ;
  assign n1421 = ~x175 & ~x271 ;
  assign n1422 = x175 & x271 ;
  assign n1423 = ~n1421 & ~n1422 ;
  assign n1424 = ~x174 & ~x270 ;
  assign n1425 = x174 & x270 ;
  assign n1426 = ~n1424 & ~n1425 ;
  assign n1427 = ~n1423 & ~n1426 ;
  assign n1428 = n1423 & n1426 ;
  assign n1429 = ~n1427 & ~n1428 ;
  assign n1430 = ~x176 & ~x272 ;
  assign n1431 = x176 & x272 ;
  assign n1432 = ~n1430 & ~n1431 ;
  assign n1433 = ~n1429 & ~n1432 ;
  assign n1434 = n1429 & n1432 ;
  assign n1435 = ~n1433 & ~n1434 ;
  assign n1436 = ~x170 & ~x266 ;
  assign n1437 = x170 & x266 ;
  assign n1438 = ~n1436 & ~n1437 ;
  assign n1439 = ~n1435 & ~n1438 ;
  assign n1440 = n1435 & n1438 ;
  assign n1441 = ~n1439 & ~n1440 ;
  assign n1442 = ~x172 & ~x268 ;
  assign n1443 = x172 & x268 ;
  assign n1444 = ~n1442 & ~n1443 ;
  assign n1445 = ~x171 & ~x267 ;
  assign n1446 = x171 & x267 ;
  assign n1447 = ~n1445 & ~n1446 ;
  assign n1448 = ~n1444 & ~n1447 ;
  assign n1449 = n1444 & n1447 ;
  assign n1450 = ~n1448 & ~n1449 ;
  assign n1451 = ~x173 & ~x269 ;
  assign n1452 = x173 & x269 ;
  assign n1453 = ~n1451 & ~n1452 ;
  assign n1454 = ~n1450 & ~n1453 ;
  assign n1455 = n1450 & n1453 ;
  assign n1456 = ~n1454 & ~n1455 ;
  assign n1457 = n1441 & ~n1456 ;
  assign n1458 = ~n1439 & ~n1457 ;
  assign n1459 = ~n1428 & ~n1434 ;
  assign n1460 = ~n1458 & n1459 ;
  assign n1461 = n1458 & ~n1459 ;
  assign n1462 = ~n1460 & ~n1461 ;
  assign n1463 = ~n1449 & ~n1455 ;
  assign n1464 = n1462 & n1463 ;
  assign n1465 = ~n1460 & ~n1464 ;
  assign n1466 = ~n1462 & ~n1463 ;
  assign n1467 = ~n1464 & ~n1466 ;
  assign n1468 = ~n1441 & n1456 ;
  assign n1469 = ~n1457 & ~n1468 ;
  assign n1470 = ~x162 & ~x258 ;
  assign n1471 = x162 & x258 ;
  assign n1472 = ~n1470 & ~n1471 ;
  assign n1473 = n1469 & ~n1472 ;
  assign n1474 = ~x168 & ~x264 ;
  assign n1475 = x168 & x264 ;
  assign n1476 = ~n1474 & ~n1475 ;
  assign n1477 = ~x167 & ~x263 ;
  assign n1478 = x167 & x263 ;
  assign n1479 = ~n1477 & ~n1478 ;
  assign n1480 = ~n1476 & ~n1479 ;
  assign n1481 = n1476 & n1479 ;
  assign n1482 = ~n1480 & ~n1481 ;
  assign n1483 = ~x169 & ~x265 ;
  assign n1484 = x169 & x265 ;
  assign n1485 = ~n1483 & ~n1484 ;
  assign n1486 = ~n1482 & ~n1485 ;
  assign n1487 = n1482 & n1485 ;
  assign n1488 = ~n1486 & ~n1487 ;
  assign n1489 = ~x163 & ~x259 ;
  assign n1490 = x163 & x259 ;
  assign n1491 = ~n1489 & ~n1490 ;
  assign n1492 = ~n1488 & ~n1491 ;
  assign n1493 = n1488 & n1491 ;
  assign n1494 = ~n1492 & ~n1493 ;
  assign n1495 = ~x165 & ~x261 ;
  assign n1496 = x165 & x261 ;
  assign n1497 = ~n1495 & ~n1496 ;
  assign n1498 = ~x164 & ~x260 ;
  assign n1499 = x164 & x260 ;
  assign n1500 = ~n1498 & ~n1499 ;
  assign n1501 = ~n1497 & ~n1500 ;
  assign n1502 = n1497 & n1500 ;
  assign n1503 = ~n1501 & ~n1502 ;
  assign n1504 = ~x166 & ~x262 ;
  assign n1505 = x166 & x262 ;
  assign n1506 = ~n1504 & ~n1505 ;
  assign n1507 = ~n1503 & ~n1506 ;
  assign n1508 = n1503 & n1506 ;
  assign n1509 = ~n1507 & ~n1508 ;
  assign n1510 = n1494 & ~n1509 ;
  assign n1511 = ~n1494 & n1509 ;
  assign n1512 = ~n1510 & ~n1511 ;
  assign n1513 = ~n1469 & n1472 ;
  assign n1514 = ~n1473 & ~n1513 ;
  assign n1515 = n1512 & n1514 ;
  assign n1516 = ~n1473 & ~n1515 ;
  assign n1517 = n1467 & ~n1516 ;
  assign n1518 = ~n1492 & ~n1510 ;
  assign n1519 = ~n1481 & ~n1487 ;
  assign n1520 = ~n1518 & n1519 ;
  assign n1521 = n1518 & ~n1519 ;
  assign n1522 = ~n1520 & ~n1521 ;
  assign n1523 = ~n1502 & ~n1508 ;
  assign n1524 = n1522 & n1523 ;
  assign n1525 = ~n1522 & ~n1523 ;
  assign n1526 = ~n1524 & ~n1525 ;
  assign n1527 = ~n1467 & n1516 ;
  assign n1528 = ~n1517 & ~n1527 ;
  assign n1529 = n1526 & n1528 ;
  assign n1530 = ~n1517 & ~n1529 ;
  assign n1531 = ~n1465 & ~n1530 ;
  assign n1532 = n1465 & n1530 ;
  assign n1533 = ~n1531 & ~n1532 ;
  assign n1534 = ~n1520 & ~n1524 ;
  assign n1535 = n1533 & ~n1534 ;
  assign n1536 = ~n1533 & n1534 ;
  assign n1537 = ~n1535 & ~n1536 ;
  assign n1538 = ~x190 & ~x286 ;
  assign n1539 = x190 & x286 ;
  assign n1540 = ~n1538 & ~n1539 ;
  assign n1541 = ~x189 & ~x285 ;
  assign n1542 = x189 & x285 ;
  assign n1543 = ~n1541 & ~n1542 ;
  assign n1544 = n1540 & n1543 ;
  assign n1545 = ~n1540 & ~n1543 ;
  assign n1546 = ~n1544 & ~n1545 ;
  assign n1547 = ~x191 & ~x287 ;
  assign n1548 = x191 & x287 ;
  assign n1549 = ~n1547 & ~n1548 ;
  assign n1550 = ~n1546 & ~n1549 ;
  assign n1551 = n1546 & n1549 ;
  assign n1552 = ~n1550 & ~n1551 ;
  assign n1553 = ~x185 & ~x281 ;
  assign n1554 = x185 & x281 ;
  assign n1555 = ~n1553 & ~n1554 ;
  assign n1556 = ~n1552 & ~n1555 ;
  assign n1557 = n1552 & n1555 ;
  assign n1558 = ~n1556 & ~n1557 ;
  assign n1559 = ~x187 & ~x283 ;
  assign n1560 = x187 & x283 ;
  assign n1561 = ~n1559 & ~n1560 ;
  assign n1562 = ~x186 & ~x282 ;
  assign n1563 = x186 & x282 ;
  assign n1564 = ~n1562 & ~n1563 ;
  assign n1565 = ~n1561 & ~n1564 ;
  assign n1566 = n1561 & n1564 ;
  assign n1567 = ~n1565 & ~n1566 ;
  assign n1568 = ~x188 & ~x284 ;
  assign n1569 = x188 & x284 ;
  assign n1570 = ~n1568 & ~n1569 ;
  assign n1571 = ~n1567 & ~n1570 ;
  assign n1572 = n1567 & n1570 ;
  assign n1573 = ~n1571 & ~n1572 ;
  assign n1574 = n1558 & ~n1573 ;
  assign n1575 = ~n1556 & ~n1574 ;
  assign n1576 = ~n1544 & ~n1551 ;
  assign n1577 = ~n1575 & n1576 ;
  assign n1578 = n1575 & ~n1576 ;
  assign n1579 = ~n1577 & ~n1578 ;
  assign n1580 = ~n1566 & ~n1572 ;
  assign n1581 = n1579 & n1580 ;
  assign n1582 = ~n1577 & ~n1581 ;
  assign n1583 = ~n1579 & ~n1580 ;
  assign n1584 = ~n1581 & ~n1583 ;
  assign n1585 = ~n1558 & n1573 ;
  assign n1586 = ~n1574 & ~n1585 ;
  assign n1587 = ~x177 & ~x273 ;
  assign n1588 = x177 & x273 ;
  assign n1589 = ~n1587 & ~n1588 ;
  assign n1590 = n1586 & ~n1589 ;
  assign n1591 = ~x183 & ~x279 ;
  assign n1592 = x183 & x279 ;
  assign n1593 = ~n1591 & ~n1592 ;
  assign n1594 = ~x182 & ~x278 ;
  assign n1595 = x182 & x278 ;
  assign n1596 = ~n1594 & ~n1595 ;
  assign n1597 = ~n1593 & ~n1596 ;
  assign n1598 = n1593 & n1596 ;
  assign n1599 = ~n1597 & ~n1598 ;
  assign n1600 = ~x184 & ~x280 ;
  assign n1601 = x184 & x280 ;
  assign n1602 = ~n1600 & ~n1601 ;
  assign n1603 = ~n1599 & ~n1602 ;
  assign n1604 = n1599 & n1602 ;
  assign n1605 = ~n1603 & ~n1604 ;
  assign n1606 = ~x178 & ~x274 ;
  assign n1607 = x178 & x274 ;
  assign n1608 = ~n1606 & ~n1607 ;
  assign n1609 = ~n1605 & ~n1608 ;
  assign n1610 = n1605 & n1608 ;
  assign n1611 = ~n1609 & ~n1610 ;
  assign n1612 = ~x180 & ~x276 ;
  assign n1613 = x180 & x276 ;
  assign n1614 = ~n1612 & ~n1613 ;
  assign n1615 = ~x179 & ~x275 ;
  assign n1616 = x179 & x275 ;
  assign n1617 = ~n1615 & ~n1616 ;
  assign n1618 = ~n1614 & ~n1617 ;
  assign n1619 = n1614 & n1617 ;
  assign n1620 = ~n1618 & ~n1619 ;
  assign n1621 = ~x181 & ~x277 ;
  assign n1622 = x181 & x277 ;
  assign n1623 = ~n1621 & ~n1622 ;
  assign n1624 = ~n1620 & ~n1623 ;
  assign n1625 = n1620 & n1623 ;
  assign n1626 = ~n1624 & ~n1625 ;
  assign n1627 = n1611 & ~n1626 ;
  assign n1628 = ~n1611 & n1626 ;
  assign n1629 = ~n1627 & ~n1628 ;
  assign n1630 = ~n1586 & n1589 ;
  assign n1631 = ~n1590 & ~n1630 ;
  assign n1632 = n1629 & n1631 ;
  assign n1633 = ~n1590 & ~n1632 ;
  assign n1634 = n1584 & ~n1633 ;
  assign n1635 = ~n1609 & ~n1627 ;
  assign n1636 = ~n1598 & ~n1604 ;
  assign n1637 = ~n1635 & n1636 ;
  assign n1638 = n1635 & ~n1636 ;
  assign n1639 = ~n1637 & ~n1638 ;
  assign n1640 = ~n1619 & ~n1625 ;
  assign n1641 = n1639 & n1640 ;
  assign n1642 = ~n1639 & ~n1640 ;
  assign n1643 = ~n1641 & ~n1642 ;
  assign n1644 = ~n1584 & n1633 ;
  assign n1645 = ~n1634 & ~n1644 ;
  assign n1646 = n1643 & n1645 ;
  assign n1647 = ~n1634 & ~n1646 ;
  assign n1648 = ~n1582 & ~n1647 ;
  assign n1649 = n1582 & n1647 ;
  assign n1650 = ~n1648 & ~n1649 ;
  assign n1651 = ~n1637 & ~n1641 ;
  assign n1652 = n1650 & ~n1651 ;
  assign n1653 = ~n1650 & n1651 ;
  assign n1654 = ~n1652 & ~n1653 ;
  assign n1655 = ~n1643 & ~n1645 ;
  assign n1656 = ~n1646 & ~n1655 ;
  assign n1657 = ~n1629 & ~n1631 ;
  assign n1658 = ~n1632 & ~n1657 ;
  assign n1659 = ~x161 & ~x257 ;
  assign n1660 = x161 & x257 ;
  assign n1661 = ~n1659 & ~n1660 ;
  assign n1662 = n1658 & ~n1661 ;
  assign n1663 = ~n1512 & ~n1514 ;
  assign n1664 = ~n1515 & ~n1663 ;
  assign n1665 = ~n1658 & n1661 ;
  assign n1666 = ~n1662 & ~n1665 ;
  assign n1667 = n1664 & n1666 ;
  assign n1668 = ~n1662 & ~n1667 ;
  assign n1669 = n1656 & ~n1668 ;
  assign n1670 = ~n1526 & ~n1528 ;
  assign n1671 = ~n1529 & ~n1670 ;
  assign n1672 = ~n1656 & n1668 ;
  assign n1673 = ~n1669 & ~n1672 ;
  assign n1674 = n1671 & n1673 ;
  assign n1675 = ~n1669 & ~n1674 ;
  assign n1676 = n1654 & ~n1675 ;
  assign n1677 = ~n1654 & n1675 ;
  assign n1678 = ~n1676 & ~n1677 ;
  assign n1679 = n1537 & n1678 ;
  assign n1680 = ~n1537 & ~n1678 ;
  assign n1681 = ~n1679 & ~n1680 ;
  assign n1682 = ~n1671 & ~n1673 ;
  assign n1683 = ~n1674 & ~n1682 ;
  assign n1684 = ~n1664 & ~n1666 ;
  assign n1685 = ~n1667 & ~n1684 ;
  assign n1686 = ~x160 & ~x256 ;
  assign n1687 = x160 & x256 ;
  assign n1688 = ~n1686 & ~n1687 ;
  assign n1689 = ~n1685 & n1688 ;
  assign n1690 = ~n1683 & n1689 ;
  assign n1691 = ~n1681 & n1690 ;
  assign n1692 = ~n1648 & ~n1652 ;
  assign n1693 = ~n1676 & ~n1679 ;
  assign n1694 = ~n1692 & ~n1693 ;
  assign n1695 = n1692 & n1693 ;
  assign n1696 = ~n1694 & ~n1695 ;
  assign n1697 = ~n1531 & ~n1535 ;
  assign n1698 = n1696 & ~n1697 ;
  assign n1699 = ~n1696 & n1697 ;
  assign n1700 = ~n1698 & ~n1699 ;
  assign n1701 = n1691 & ~n1700 ;
  assign n1702 = ~n1694 & ~n1698 ;
  assign n1703 = n1701 & n1702 ;
  assign n1704 = ~x254 & ~x286 ;
  assign n1705 = x254 & x286 ;
  assign n1706 = ~n1704 & ~n1705 ;
  assign n1707 = ~x253 & ~x285 ;
  assign n1708 = x253 & x285 ;
  assign n1709 = ~n1707 & ~n1708 ;
  assign n1710 = n1706 & n1709 ;
  assign n1711 = ~n1706 & ~n1709 ;
  assign n1712 = ~n1710 & ~n1711 ;
  assign n1713 = ~x255 & ~x287 ;
  assign n1714 = x255 & x287 ;
  assign n1715 = ~n1713 & ~n1714 ;
  assign n1716 = n1712 & n1715 ;
  assign n1717 = ~n1710 & ~n1716 ;
  assign n1718 = ~n1712 & ~n1715 ;
  assign n1719 = ~n1716 & ~n1718 ;
  assign n1720 = ~x249 & ~x281 ;
  assign n1721 = x249 & x281 ;
  assign n1722 = ~n1720 & ~n1721 ;
  assign n1723 = n1719 & n1722 ;
  assign n1724 = ~n1719 & ~n1722 ;
  assign n1725 = ~x251 & ~x283 ;
  assign n1726 = x251 & x283 ;
  assign n1727 = ~n1725 & ~n1726 ;
  assign n1728 = ~x250 & ~x282 ;
  assign n1729 = x250 & x282 ;
  assign n1730 = ~n1728 & ~n1729 ;
  assign n1731 = ~n1727 & ~n1730 ;
  assign n1732 = n1727 & n1730 ;
  assign n1733 = ~n1731 & ~n1732 ;
  assign n1734 = ~x252 & ~x284 ;
  assign n1735 = x252 & x284 ;
  assign n1736 = ~n1734 & ~n1735 ;
  assign n1737 = ~n1733 & ~n1736 ;
  assign n1738 = n1733 & n1736 ;
  assign n1739 = ~n1737 & ~n1738 ;
  assign n1740 = ~n1724 & n1739 ;
  assign n1741 = ~n1723 & ~n1740 ;
  assign n1742 = n1717 & n1741 ;
  assign n1743 = ~n1717 & ~n1741 ;
  assign n1744 = ~n1742 & ~n1743 ;
  assign n1745 = ~n1732 & ~n1738 ;
  assign n1746 = n1744 & n1745 ;
  assign n1747 = ~n1742 & ~n1746 ;
  assign n1748 = ~n1744 & ~n1745 ;
  assign n1749 = ~n1746 & ~n1748 ;
  assign n1750 = ~n1723 & ~n1724 ;
  assign n1751 = ~n1739 & n1750 ;
  assign n1752 = n1739 & ~n1750 ;
  assign n1753 = ~n1751 & ~n1752 ;
  assign n1754 = ~x241 & ~x273 ;
  assign n1755 = x241 & x273 ;
  assign n1756 = ~n1754 & ~n1755 ;
  assign n1757 = ~n1753 & n1756 ;
  assign n1758 = n1753 & ~n1756 ;
  assign n1759 = ~x247 & ~x279 ;
  assign n1760 = x247 & x279 ;
  assign n1761 = ~n1759 & ~n1760 ;
  assign n1762 = ~x246 & ~x278 ;
  assign n1763 = x246 & x278 ;
  assign n1764 = ~n1762 & ~n1763 ;
  assign n1765 = ~n1761 & ~n1764 ;
  assign n1766 = n1761 & n1764 ;
  assign n1767 = ~n1765 & ~n1766 ;
  assign n1768 = ~x248 & ~x280 ;
  assign n1769 = x248 & x280 ;
  assign n1770 = ~n1768 & ~n1769 ;
  assign n1771 = ~n1767 & ~n1770 ;
  assign n1772 = n1767 & n1770 ;
  assign n1773 = ~n1771 & ~n1772 ;
  assign n1774 = ~x242 & ~x274 ;
  assign n1775 = x242 & x274 ;
  assign n1776 = ~n1774 & ~n1775 ;
  assign n1777 = ~n1773 & ~n1776 ;
  assign n1778 = n1773 & n1776 ;
  assign n1779 = ~n1777 & ~n1778 ;
  assign n1780 = ~x244 & ~x276 ;
  assign n1781 = x244 & x276 ;
  assign n1782 = ~n1780 & ~n1781 ;
  assign n1783 = ~x243 & ~x275 ;
  assign n1784 = x243 & x275 ;
  assign n1785 = ~n1783 & ~n1784 ;
  assign n1786 = ~n1782 & ~n1785 ;
  assign n1787 = n1782 & n1785 ;
  assign n1788 = ~n1786 & ~n1787 ;
  assign n1789 = ~x245 & ~x277 ;
  assign n1790 = x245 & x277 ;
  assign n1791 = ~n1789 & ~n1790 ;
  assign n1792 = ~n1788 & ~n1791 ;
  assign n1793 = n1788 & n1791 ;
  assign n1794 = ~n1792 & ~n1793 ;
  assign n1795 = n1779 & ~n1794 ;
  assign n1796 = ~n1779 & n1794 ;
  assign n1797 = ~n1795 & ~n1796 ;
  assign n1798 = ~n1758 & ~n1797 ;
  assign n1799 = ~n1757 & ~n1798 ;
  assign n1800 = n1749 & n1799 ;
  assign n1801 = ~n1749 & ~n1799 ;
  assign n1802 = ~n1777 & ~n1795 ;
  assign n1803 = ~n1766 & ~n1772 ;
  assign n1804 = ~n1802 & n1803 ;
  assign n1805 = n1802 & ~n1803 ;
  assign n1806 = ~n1804 & ~n1805 ;
  assign n1807 = ~n1787 & ~n1793 ;
  assign n1808 = n1806 & n1807 ;
  assign n1809 = ~n1806 & ~n1807 ;
  assign n1810 = ~n1808 & ~n1809 ;
  assign n1811 = ~n1801 & n1810 ;
  assign n1812 = ~n1800 & ~n1811 ;
  assign n1813 = ~n1747 & ~n1812 ;
  assign n1814 = n1747 & n1812 ;
  assign n1815 = ~n1813 & ~n1814 ;
  assign n1816 = ~n1804 & ~n1808 ;
  assign n1817 = n1815 & ~n1816 ;
  assign n1818 = ~n1813 & ~n1817 ;
  assign n1819 = ~n1815 & n1816 ;
  assign n1820 = ~n1817 & ~n1819 ;
  assign n1821 = ~x225 & ~x257 ;
  assign n1822 = x225 & x257 ;
  assign n1823 = ~n1821 & ~n1822 ;
  assign n1824 = ~n1757 & ~n1758 ;
  assign n1825 = ~n1797 & n1824 ;
  assign n1826 = n1797 & ~n1824 ;
  assign n1827 = ~n1825 & ~n1826 ;
  assign n1828 = ~n1823 & ~n1827 ;
  assign n1829 = n1823 & n1827 ;
  assign n1830 = ~x232 & ~x264 ;
  assign n1831 = x232 & x264 ;
  assign n1832 = ~n1830 & ~n1831 ;
  assign n1833 = ~x231 & ~x263 ;
  assign n1834 = x231 & x263 ;
  assign n1835 = ~n1833 & ~n1834 ;
  assign n1836 = ~n1832 & ~n1835 ;
  assign n1837 = n1832 & n1835 ;
  assign n1838 = ~n1836 & ~n1837 ;
  assign n1839 = ~x233 & ~x265 ;
  assign n1840 = x233 & x265 ;
  assign n1841 = ~n1839 & ~n1840 ;
  assign n1842 = ~n1838 & ~n1841 ;
  assign n1843 = n1838 & n1841 ;
  assign n1844 = ~n1842 & ~n1843 ;
  assign n1845 = ~x227 & ~x259 ;
  assign n1846 = x227 & x259 ;
  assign n1847 = ~n1845 & ~n1846 ;
  assign n1848 = ~n1844 & ~n1847 ;
  assign n1849 = n1844 & n1847 ;
  assign n1850 = ~n1848 & ~n1849 ;
  assign n1851 = ~x229 & ~x261 ;
  assign n1852 = x229 & x261 ;
  assign n1853 = ~n1851 & ~n1852 ;
  assign n1854 = ~x228 & ~x260 ;
  assign n1855 = x228 & x260 ;
  assign n1856 = ~n1854 & ~n1855 ;
  assign n1857 = ~n1853 & ~n1856 ;
  assign n1858 = n1853 & n1856 ;
  assign n1859 = ~n1857 & ~n1858 ;
  assign n1860 = ~x230 & ~x262 ;
  assign n1861 = x230 & x262 ;
  assign n1862 = ~n1860 & ~n1861 ;
  assign n1863 = ~n1859 & ~n1862 ;
  assign n1864 = n1859 & n1862 ;
  assign n1865 = ~n1863 & ~n1864 ;
  assign n1866 = n1850 & ~n1865 ;
  assign n1867 = ~n1850 & n1865 ;
  assign n1868 = ~n1866 & ~n1867 ;
  assign n1869 = ~x239 & ~x271 ;
  assign n1870 = x239 & x271 ;
  assign n1871 = ~n1869 & ~n1870 ;
  assign n1872 = ~x238 & ~x270 ;
  assign n1873 = x238 & x270 ;
  assign n1874 = ~n1872 & ~n1873 ;
  assign n1875 = ~n1871 & ~n1874 ;
  assign n1876 = n1871 & n1874 ;
  assign n1877 = ~n1875 & ~n1876 ;
  assign n1878 = ~x240 & ~x272 ;
  assign n1879 = x240 & x272 ;
  assign n1880 = ~n1878 & ~n1879 ;
  assign n1881 = ~n1877 & ~n1880 ;
  assign n1882 = n1877 & n1880 ;
  assign n1883 = ~n1881 & ~n1882 ;
  assign n1884 = ~x234 & ~x266 ;
  assign n1885 = x234 & x266 ;
  assign n1886 = ~n1884 & ~n1885 ;
  assign n1887 = ~n1883 & ~n1886 ;
  assign n1888 = n1883 & n1886 ;
  assign n1889 = ~n1887 & ~n1888 ;
  assign n1890 = ~x236 & ~x268 ;
  assign n1891 = x236 & x268 ;
  assign n1892 = ~n1890 & ~n1891 ;
  assign n1893 = ~x235 & ~x267 ;
  assign n1894 = x235 & x267 ;
  assign n1895 = ~n1893 & ~n1894 ;
  assign n1896 = ~n1892 & ~n1895 ;
  assign n1897 = n1892 & n1895 ;
  assign n1898 = ~n1896 & ~n1897 ;
  assign n1899 = ~x237 & ~x269 ;
  assign n1900 = x237 & x269 ;
  assign n1901 = ~n1899 & ~n1900 ;
  assign n1902 = ~n1898 & ~n1901 ;
  assign n1903 = n1898 & n1901 ;
  assign n1904 = ~n1902 & ~n1903 ;
  assign n1905 = n1889 & ~n1904 ;
  assign n1906 = ~n1889 & n1904 ;
  assign n1907 = ~n1905 & ~n1906 ;
  assign n1908 = ~x226 & ~x258 ;
  assign n1909 = x226 & x258 ;
  assign n1910 = ~n1908 & ~n1909 ;
  assign n1911 = n1907 & ~n1910 ;
  assign n1912 = ~n1907 & n1910 ;
  assign n1913 = ~n1911 & ~n1912 ;
  assign n1914 = n1868 & n1913 ;
  assign n1915 = ~n1868 & ~n1913 ;
  assign n1916 = ~n1914 & ~n1915 ;
  assign n1917 = ~n1829 & n1916 ;
  assign n1918 = ~n1828 & ~n1917 ;
  assign n1919 = ~n1800 & ~n1801 ;
  assign n1920 = ~n1810 & n1919 ;
  assign n1921 = n1810 & ~n1919 ;
  assign n1922 = ~n1920 & ~n1921 ;
  assign n1923 = n1918 & n1922 ;
  assign n1924 = ~n1918 & ~n1922 ;
  assign n1925 = ~n1848 & ~n1866 ;
  assign n1926 = ~n1837 & ~n1843 ;
  assign n1927 = ~n1925 & n1926 ;
  assign n1928 = n1925 & ~n1926 ;
  assign n1929 = ~n1927 & ~n1928 ;
  assign n1930 = ~n1858 & ~n1864 ;
  assign n1931 = n1929 & n1930 ;
  assign n1932 = ~n1929 & ~n1930 ;
  assign n1933 = ~n1931 & ~n1932 ;
  assign n1934 = ~n1887 & ~n1905 ;
  assign n1935 = ~n1876 & ~n1882 ;
  assign n1936 = ~n1934 & n1935 ;
  assign n1937 = n1934 & ~n1935 ;
  assign n1938 = ~n1936 & ~n1937 ;
  assign n1939 = ~n1897 & ~n1903 ;
  assign n1940 = n1938 & n1939 ;
  assign n1941 = ~n1938 & ~n1939 ;
  assign n1942 = ~n1940 & ~n1941 ;
  assign n1943 = ~n1911 & ~n1914 ;
  assign n1944 = n1942 & ~n1943 ;
  assign n1945 = ~n1942 & n1943 ;
  assign n1946 = ~n1944 & ~n1945 ;
  assign n1947 = n1933 & n1946 ;
  assign n1948 = ~n1933 & ~n1946 ;
  assign n1949 = ~n1947 & ~n1948 ;
  assign n1950 = ~n1924 & ~n1949 ;
  assign n1951 = ~n1923 & ~n1950 ;
  assign n1952 = ~n1820 & ~n1951 ;
  assign n1953 = n1820 & n1951 ;
  assign n1954 = ~n1933 & ~n1944 ;
  assign n1955 = ~n1945 & ~n1954 ;
  assign n1956 = ~n1936 & ~n1940 ;
  assign n1957 = n1955 & ~n1956 ;
  assign n1958 = ~n1955 & n1956 ;
  assign n1959 = ~n1957 & ~n1958 ;
  assign n1960 = ~n1927 & ~n1931 ;
  assign n1961 = n1959 & ~n1960 ;
  assign n1962 = ~n1959 & n1960 ;
  assign n1963 = ~n1961 & ~n1962 ;
  assign n1964 = ~n1953 & ~n1963 ;
  assign n1965 = ~n1952 & ~n1964 ;
  assign n1966 = ~n1818 & n1965 ;
  assign n1967 = n1818 & ~n1965 ;
  assign n1968 = ~n1966 & ~n1967 ;
  assign n1969 = ~n1957 & ~n1961 ;
  assign n1970 = n1968 & ~n1969 ;
  assign n1971 = ~n1968 & n1969 ;
  assign n1972 = ~n1970 & ~n1971 ;
  assign n1973 = ~x224 & ~x256 ;
  assign n1974 = x224 & x256 ;
  assign n1975 = ~n1973 & ~n1974 ;
  assign n1976 = ~n1828 & ~n1829 ;
  assign n1977 = n1916 & n1976 ;
  assign n1978 = ~n1916 & ~n1976 ;
  assign n1979 = ~n1977 & ~n1978 ;
  assign n1980 = n1975 & ~n1979 ;
  assign n1981 = ~n1923 & ~n1924 ;
  assign n1982 = ~n1949 & n1981 ;
  assign n1983 = n1949 & ~n1981 ;
  assign n1984 = ~n1982 & ~n1983 ;
  assign n1985 = n1980 & n1984 ;
  assign n1986 = ~n1952 & ~n1953 ;
  assign n1987 = ~n1963 & n1986 ;
  assign n1988 = n1963 & ~n1986 ;
  assign n1989 = ~n1987 & ~n1988 ;
  assign n1990 = n1985 & n1989 ;
  assign n1991 = ~n1972 & n1990 ;
  assign n1992 = ~n1966 & ~n1970 ;
  assign n1993 = n1991 & n1992 ;
  assign n1994 = ~x222 & ~x286 ;
  assign n1995 = x222 & x286 ;
  assign n1996 = ~n1994 & ~n1995 ;
  assign n1997 = ~x221 & ~x285 ;
  assign n1998 = x221 & x285 ;
  assign n1999 = ~n1997 & ~n1998 ;
  assign n2000 = n1996 & n1999 ;
  assign n2001 = ~n1996 & ~n1999 ;
  assign n2002 = ~n2000 & ~n2001 ;
  assign n2003 = ~x223 & ~x287 ;
  assign n2004 = x223 & x287 ;
  assign n2005 = ~n2003 & ~n2004 ;
  assign n2006 = n2002 & n2005 ;
  assign n2007 = ~n2000 & ~n2006 ;
  assign n2008 = ~n2002 & ~n2005 ;
  assign n2009 = ~n2006 & ~n2008 ;
  assign n2010 = ~x217 & ~x281 ;
  assign n2011 = x217 & x281 ;
  assign n2012 = ~n2010 & ~n2011 ;
  assign n2013 = n2009 & n2012 ;
  assign n2014 = ~n2009 & ~n2012 ;
  assign n2015 = ~x219 & ~x283 ;
  assign n2016 = x219 & x283 ;
  assign n2017 = ~n2015 & ~n2016 ;
  assign n2018 = ~x218 & ~x282 ;
  assign n2019 = x218 & x282 ;
  assign n2020 = ~n2018 & ~n2019 ;
  assign n2021 = ~n2017 & ~n2020 ;
  assign n2022 = n2017 & n2020 ;
  assign n2023 = ~n2021 & ~n2022 ;
  assign n2024 = ~x220 & ~x284 ;
  assign n2025 = x220 & x284 ;
  assign n2026 = ~n2024 & ~n2025 ;
  assign n2027 = ~n2023 & ~n2026 ;
  assign n2028 = n2023 & n2026 ;
  assign n2029 = ~n2027 & ~n2028 ;
  assign n2030 = ~n2014 & n2029 ;
  assign n2031 = ~n2013 & ~n2030 ;
  assign n2032 = n2007 & n2031 ;
  assign n2033 = ~n2007 & ~n2031 ;
  assign n2034 = ~n2032 & ~n2033 ;
  assign n2035 = ~n2022 & ~n2028 ;
  assign n2036 = n2034 & n2035 ;
  assign n2037 = ~n2032 & ~n2036 ;
  assign n2038 = ~n2034 & ~n2035 ;
  assign n2039 = ~n2036 & ~n2038 ;
  assign n2040 = ~n2013 & ~n2014 ;
  assign n2041 = ~n2029 & n2040 ;
  assign n2042 = n2029 & ~n2040 ;
  assign n2043 = ~n2041 & ~n2042 ;
  assign n2044 = ~x209 & ~x273 ;
  assign n2045 = x209 & x273 ;
  assign n2046 = ~n2044 & ~n2045 ;
  assign n2047 = ~n2043 & n2046 ;
  assign n2048 = n2043 & ~n2046 ;
  assign n2049 = ~x215 & ~x279 ;
  assign n2050 = x215 & x279 ;
  assign n2051 = ~n2049 & ~n2050 ;
  assign n2052 = ~x214 & ~x278 ;
  assign n2053 = x214 & x278 ;
  assign n2054 = ~n2052 & ~n2053 ;
  assign n2055 = ~n2051 & ~n2054 ;
  assign n2056 = n2051 & n2054 ;
  assign n2057 = ~n2055 & ~n2056 ;
  assign n2058 = ~x216 & ~x280 ;
  assign n2059 = x216 & x280 ;
  assign n2060 = ~n2058 & ~n2059 ;
  assign n2061 = ~n2057 & ~n2060 ;
  assign n2062 = n2057 & n2060 ;
  assign n2063 = ~n2061 & ~n2062 ;
  assign n2064 = ~x210 & ~x274 ;
  assign n2065 = x210 & x274 ;
  assign n2066 = ~n2064 & ~n2065 ;
  assign n2067 = ~n2063 & ~n2066 ;
  assign n2068 = n2063 & n2066 ;
  assign n2069 = ~n2067 & ~n2068 ;
  assign n2070 = ~x212 & ~x276 ;
  assign n2071 = x212 & x276 ;
  assign n2072 = ~n2070 & ~n2071 ;
  assign n2073 = ~x211 & ~x275 ;
  assign n2074 = x211 & x275 ;
  assign n2075 = ~n2073 & ~n2074 ;
  assign n2076 = ~n2072 & ~n2075 ;
  assign n2077 = n2072 & n2075 ;
  assign n2078 = ~n2076 & ~n2077 ;
  assign n2079 = ~x213 & ~x277 ;
  assign n2080 = x213 & x277 ;
  assign n2081 = ~n2079 & ~n2080 ;
  assign n2082 = ~n2078 & ~n2081 ;
  assign n2083 = n2078 & n2081 ;
  assign n2084 = ~n2082 & ~n2083 ;
  assign n2085 = n2069 & ~n2084 ;
  assign n2086 = ~n2069 & n2084 ;
  assign n2087 = ~n2085 & ~n2086 ;
  assign n2088 = ~n2048 & ~n2087 ;
  assign n2089 = ~n2047 & ~n2088 ;
  assign n2090 = n2039 & n2089 ;
  assign n2091 = ~n2039 & ~n2089 ;
  assign n2092 = ~n2067 & ~n2085 ;
  assign n2093 = ~n2056 & ~n2062 ;
  assign n2094 = ~n2092 & n2093 ;
  assign n2095 = n2092 & ~n2093 ;
  assign n2096 = ~n2094 & ~n2095 ;
  assign n2097 = ~n2077 & ~n2083 ;
  assign n2098 = n2096 & n2097 ;
  assign n2099 = ~n2096 & ~n2097 ;
  assign n2100 = ~n2098 & ~n2099 ;
  assign n2101 = ~n2091 & n2100 ;
  assign n2102 = ~n2090 & ~n2101 ;
  assign n2103 = ~n2037 & ~n2102 ;
  assign n2104 = n2037 & n2102 ;
  assign n2105 = ~n2103 & ~n2104 ;
  assign n2106 = ~n2094 & ~n2098 ;
  assign n2107 = n2105 & ~n2106 ;
  assign n2108 = ~n2103 & ~n2107 ;
  assign n2109 = ~n2105 & n2106 ;
  assign n2110 = ~n2107 & ~n2109 ;
  assign n2111 = ~x193 & ~x257 ;
  assign n2112 = x193 & x257 ;
  assign n2113 = ~n2111 & ~n2112 ;
  assign n2114 = ~n2047 & ~n2048 ;
  assign n2115 = ~n2087 & n2114 ;
  assign n2116 = n2087 & ~n2114 ;
  assign n2117 = ~n2115 & ~n2116 ;
  assign n2118 = ~n2113 & ~n2117 ;
  assign n2119 = n2113 & n2117 ;
  assign n2120 = ~x200 & ~x264 ;
  assign n2121 = x200 & x264 ;
  assign n2122 = ~n2120 & ~n2121 ;
  assign n2123 = ~x199 & ~x263 ;
  assign n2124 = x199 & x263 ;
  assign n2125 = ~n2123 & ~n2124 ;
  assign n2126 = ~n2122 & ~n2125 ;
  assign n2127 = n2122 & n2125 ;
  assign n2128 = ~n2126 & ~n2127 ;
  assign n2129 = ~x201 & ~x265 ;
  assign n2130 = x201 & x265 ;
  assign n2131 = ~n2129 & ~n2130 ;
  assign n2132 = ~n2128 & ~n2131 ;
  assign n2133 = n2128 & n2131 ;
  assign n2134 = ~n2132 & ~n2133 ;
  assign n2135 = ~x195 & ~x259 ;
  assign n2136 = x195 & x259 ;
  assign n2137 = ~n2135 & ~n2136 ;
  assign n2138 = ~n2134 & ~n2137 ;
  assign n2139 = n2134 & n2137 ;
  assign n2140 = ~n2138 & ~n2139 ;
  assign n2141 = ~x197 & ~x261 ;
  assign n2142 = x197 & x261 ;
  assign n2143 = ~n2141 & ~n2142 ;
  assign n2144 = ~x196 & ~x260 ;
  assign n2145 = x196 & x260 ;
  assign n2146 = ~n2144 & ~n2145 ;
  assign n2147 = ~n2143 & ~n2146 ;
  assign n2148 = n2143 & n2146 ;
  assign n2149 = ~n2147 & ~n2148 ;
  assign n2150 = ~x198 & ~x262 ;
  assign n2151 = x198 & x262 ;
  assign n2152 = ~n2150 & ~n2151 ;
  assign n2153 = ~n2149 & ~n2152 ;
  assign n2154 = n2149 & n2152 ;
  assign n2155 = ~n2153 & ~n2154 ;
  assign n2156 = n2140 & ~n2155 ;
  assign n2157 = ~n2140 & n2155 ;
  assign n2158 = ~n2156 & ~n2157 ;
  assign n2159 = ~x207 & ~x271 ;
  assign n2160 = x207 & x271 ;
  assign n2161 = ~n2159 & ~n2160 ;
  assign n2162 = ~x206 & ~x270 ;
  assign n2163 = x206 & x270 ;
  assign n2164 = ~n2162 & ~n2163 ;
  assign n2165 = ~n2161 & ~n2164 ;
  assign n2166 = n2161 & n2164 ;
  assign n2167 = ~n2165 & ~n2166 ;
  assign n2168 = ~x208 & ~x272 ;
  assign n2169 = x208 & x272 ;
  assign n2170 = ~n2168 & ~n2169 ;
  assign n2171 = ~n2167 & ~n2170 ;
  assign n2172 = n2167 & n2170 ;
  assign n2173 = ~n2171 & ~n2172 ;
  assign n2174 = ~x202 & ~x266 ;
  assign n2175 = x202 & x266 ;
  assign n2176 = ~n2174 & ~n2175 ;
  assign n2177 = ~n2173 & ~n2176 ;
  assign n2178 = n2173 & n2176 ;
  assign n2179 = ~n2177 & ~n2178 ;
  assign n2180 = ~x204 & ~x268 ;
  assign n2181 = x204 & x268 ;
  assign n2182 = ~n2180 & ~n2181 ;
  assign n2183 = ~x203 & ~x267 ;
  assign n2184 = x203 & x267 ;
  assign n2185 = ~n2183 & ~n2184 ;
  assign n2186 = ~n2182 & ~n2185 ;
  assign n2187 = n2182 & n2185 ;
  assign n2188 = ~n2186 & ~n2187 ;
  assign n2189 = ~x205 & ~x269 ;
  assign n2190 = x205 & x269 ;
  assign n2191 = ~n2189 & ~n2190 ;
  assign n2192 = ~n2188 & ~n2191 ;
  assign n2193 = n2188 & n2191 ;
  assign n2194 = ~n2192 & ~n2193 ;
  assign n2195 = n2179 & ~n2194 ;
  assign n2196 = ~n2179 & n2194 ;
  assign n2197 = ~n2195 & ~n2196 ;
  assign n2198 = ~x194 & ~x258 ;
  assign n2199 = x194 & x258 ;
  assign n2200 = ~n2198 & ~n2199 ;
  assign n2201 = n2197 & ~n2200 ;
  assign n2202 = ~n2197 & n2200 ;
  assign n2203 = ~n2201 & ~n2202 ;
  assign n2204 = n2158 & n2203 ;
  assign n2205 = ~n2158 & ~n2203 ;
  assign n2206 = ~n2204 & ~n2205 ;
  assign n2207 = ~n2119 & n2206 ;
  assign n2208 = ~n2118 & ~n2207 ;
  assign n2209 = ~n2090 & ~n2091 ;
  assign n2210 = ~n2100 & n2209 ;
  assign n2211 = n2100 & ~n2209 ;
  assign n2212 = ~n2210 & ~n2211 ;
  assign n2213 = n2208 & n2212 ;
  assign n2214 = ~n2208 & ~n2212 ;
  assign n2215 = ~n2138 & ~n2156 ;
  assign n2216 = ~n2127 & ~n2133 ;
  assign n2217 = ~n2215 & n2216 ;
  assign n2218 = n2215 & ~n2216 ;
  assign n2219 = ~n2217 & ~n2218 ;
  assign n2220 = ~n2148 & ~n2154 ;
  assign n2221 = n2219 & n2220 ;
  assign n2222 = ~n2219 & ~n2220 ;
  assign n2223 = ~n2221 & ~n2222 ;
  assign n2224 = ~n2177 & ~n2195 ;
  assign n2225 = ~n2166 & ~n2172 ;
  assign n2226 = ~n2224 & n2225 ;
  assign n2227 = n2224 & ~n2225 ;
  assign n2228 = ~n2226 & ~n2227 ;
  assign n2229 = ~n2187 & ~n2193 ;
  assign n2230 = n2228 & n2229 ;
  assign n2231 = ~n2228 & ~n2229 ;
  assign n2232 = ~n2230 & ~n2231 ;
  assign n2233 = ~n2201 & ~n2204 ;
  assign n2234 = n2232 & ~n2233 ;
  assign n2235 = ~n2232 & n2233 ;
  assign n2236 = ~n2234 & ~n2235 ;
  assign n2237 = n2223 & n2236 ;
  assign n2238 = ~n2223 & ~n2236 ;
  assign n2239 = ~n2237 & ~n2238 ;
  assign n2240 = ~n2214 & ~n2239 ;
  assign n2241 = ~n2213 & ~n2240 ;
  assign n2242 = ~n2110 & ~n2241 ;
  assign n2243 = n2110 & n2241 ;
  assign n2244 = ~n2223 & ~n2234 ;
  assign n2245 = ~n2235 & ~n2244 ;
  assign n2246 = ~n2226 & ~n2230 ;
  assign n2247 = n2245 & ~n2246 ;
  assign n2248 = ~n2245 & n2246 ;
  assign n2249 = ~n2247 & ~n2248 ;
  assign n2250 = ~n2217 & ~n2221 ;
  assign n2251 = n2249 & ~n2250 ;
  assign n2252 = ~n2249 & n2250 ;
  assign n2253 = ~n2251 & ~n2252 ;
  assign n2254 = ~n2243 & ~n2253 ;
  assign n2255 = ~n2242 & ~n2254 ;
  assign n2256 = ~n2108 & n2255 ;
  assign n2257 = n2108 & ~n2255 ;
  assign n2258 = ~n2256 & ~n2257 ;
  assign n2259 = ~n2247 & ~n2251 ;
  assign n2260 = n2258 & ~n2259 ;
  assign n2261 = ~n2258 & n2259 ;
  assign n2262 = ~n2260 & ~n2261 ;
  assign n2263 = ~x192 & ~x256 ;
  assign n2264 = x192 & x256 ;
  assign n2265 = ~n2263 & ~n2264 ;
  assign n2266 = ~n2118 & ~n2119 ;
  assign n2267 = n2206 & n2266 ;
  assign n2268 = ~n2206 & ~n2266 ;
  assign n2269 = ~n2267 & ~n2268 ;
  assign n2270 = n2265 & ~n2269 ;
  assign n2271 = ~n2213 & ~n2214 ;
  assign n2272 = ~n2239 & n2271 ;
  assign n2273 = n2239 & ~n2271 ;
  assign n2274 = ~n2272 & ~n2273 ;
  assign n2275 = n2270 & n2274 ;
  assign n2276 = ~n2242 & ~n2243 ;
  assign n2277 = ~n2253 & n2276 ;
  assign n2278 = n2253 & ~n2276 ;
  assign n2279 = ~n2277 & ~n2278 ;
  assign n2280 = n2275 & n2279 ;
  assign n2281 = ~n2262 & n2280 ;
  assign n2282 = ~n2256 & ~n2260 ;
  assign n2283 = n2281 & n2282 ;
  assign n2284 = ~n1993 & ~n2283 ;
  assign n2285 = n1703 & ~n2284 ;
  assign n2286 = n1993 & n2283 ;
  assign n2287 = ~n1703 & n2286 ;
  assign n2288 = ~n2285 & ~n2287 ;
  assign n2289 = ~x136 & ~x264 ;
  assign n2290 = x136 & x264 ;
  assign n2291 = ~n2289 & ~n2290 ;
  assign n2292 = ~x135 & ~x263 ;
  assign n2293 = x135 & x263 ;
  assign n2294 = ~n2292 & ~n2293 ;
  assign n2295 = ~n2291 & ~n2294 ;
  assign n2296 = n2291 & n2294 ;
  assign n2297 = ~n2295 & ~n2296 ;
  assign n2298 = ~x137 & ~x265 ;
  assign n2299 = x137 & x265 ;
  assign n2300 = ~n2298 & ~n2299 ;
  assign n2301 = ~n2297 & ~n2300 ;
  assign n2302 = n2297 & n2300 ;
  assign n2303 = ~n2301 & ~n2302 ;
  assign n2304 = ~x131 & ~x259 ;
  assign n2305 = x131 & x259 ;
  assign n2306 = ~n2304 & ~n2305 ;
  assign n2307 = ~n2303 & ~n2306 ;
  assign n2308 = n2303 & n2306 ;
  assign n2309 = ~n2307 & ~n2308 ;
  assign n2310 = ~x133 & ~x261 ;
  assign n2311 = x133 & x261 ;
  assign n2312 = ~n2310 & ~n2311 ;
  assign n2313 = ~x132 & ~x260 ;
  assign n2314 = x132 & x260 ;
  assign n2315 = ~n2313 & ~n2314 ;
  assign n2316 = ~n2312 & ~n2315 ;
  assign n2317 = n2312 & n2315 ;
  assign n2318 = ~n2316 & ~n2317 ;
  assign n2319 = ~x134 & ~x262 ;
  assign n2320 = x134 & x262 ;
  assign n2321 = ~n2319 & ~n2320 ;
  assign n2322 = ~n2318 & ~n2321 ;
  assign n2323 = n2318 & n2321 ;
  assign n2324 = ~n2322 & ~n2323 ;
  assign n2325 = n2309 & ~n2324 ;
  assign n2326 = ~n2307 & ~n2325 ;
  assign n2327 = ~n2296 & ~n2302 ;
  assign n2328 = ~n2326 & n2327 ;
  assign n2329 = n2326 & ~n2327 ;
  assign n2330 = ~n2328 & ~n2329 ;
  assign n2331 = ~n2317 & ~n2323 ;
  assign n2332 = n2330 & n2331 ;
  assign n2333 = ~n2330 & ~n2331 ;
  assign n2334 = ~n2332 & ~n2333 ;
  assign n2335 = ~x143 & ~x271 ;
  assign n2336 = x143 & x271 ;
  assign n2337 = ~n2335 & ~n2336 ;
  assign n2338 = ~x142 & ~x270 ;
  assign n2339 = x142 & x270 ;
  assign n2340 = ~n2338 & ~n2339 ;
  assign n2341 = ~n2337 & ~n2340 ;
  assign n2342 = n2337 & n2340 ;
  assign n2343 = ~n2341 & ~n2342 ;
  assign n2344 = ~x144 & ~x272 ;
  assign n2345 = x144 & x272 ;
  assign n2346 = ~n2344 & ~n2345 ;
  assign n2347 = ~n2343 & ~n2346 ;
  assign n2348 = n2343 & n2346 ;
  assign n2349 = ~n2347 & ~n2348 ;
  assign n2350 = ~x138 & ~x266 ;
  assign n2351 = x138 & x266 ;
  assign n2352 = ~n2350 & ~n2351 ;
  assign n2353 = ~n2349 & ~n2352 ;
  assign n2354 = n2349 & n2352 ;
  assign n2355 = ~n2353 & ~n2354 ;
  assign n2356 = ~x140 & ~x268 ;
  assign n2357 = x140 & x268 ;
  assign n2358 = ~n2356 & ~n2357 ;
  assign n2359 = ~x139 & ~x267 ;
  assign n2360 = x139 & x267 ;
  assign n2361 = ~n2359 & ~n2360 ;
  assign n2362 = ~n2358 & ~n2361 ;
  assign n2363 = n2358 & n2361 ;
  assign n2364 = ~n2362 & ~n2363 ;
  assign n2365 = ~x141 & ~x269 ;
  assign n2366 = x141 & x269 ;
  assign n2367 = ~n2365 & ~n2366 ;
  assign n2368 = ~n2364 & ~n2367 ;
  assign n2369 = n2364 & n2367 ;
  assign n2370 = ~n2368 & ~n2369 ;
  assign n2371 = n2355 & ~n2370 ;
  assign n2372 = ~n2353 & ~n2371 ;
  assign n2373 = ~n2342 & ~n2348 ;
  assign n2374 = ~n2372 & n2373 ;
  assign n2375 = n2372 & ~n2373 ;
  assign n2376 = ~n2374 & ~n2375 ;
  assign n2377 = ~n2363 & ~n2369 ;
  assign n2378 = n2376 & n2377 ;
  assign n2379 = ~n2376 & ~n2377 ;
  assign n2380 = ~n2378 & ~n2379 ;
  assign n2381 = ~n2355 & n2370 ;
  assign n2382 = ~n2371 & ~n2381 ;
  assign n2383 = ~x130 & ~x258 ;
  assign n2384 = x130 & x258 ;
  assign n2385 = ~n2383 & ~n2384 ;
  assign n2386 = n2382 & ~n2385 ;
  assign n2387 = ~n2309 & n2324 ;
  assign n2388 = ~n2325 & ~n2387 ;
  assign n2389 = ~n2382 & n2385 ;
  assign n2390 = ~n2386 & ~n2389 ;
  assign n2391 = n2388 & n2390 ;
  assign n2392 = ~n2386 & ~n2391 ;
  assign n2393 = n2380 & ~n2392 ;
  assign n2394 = ~n2380 & n2392 ;
  assign n2395 = ~n2393 & ~n2394 ;
  assign n2396 = n2334 & n2395 ;
  assign n2397 = ~n2334 & ~n2395 ;
  assign n2398 = ~n2396 & ~n2397 ;
  assign n2399 = ~x151 & ~x279 ;
  assign n2400 = x151 & x279 ;
  assign n2401 = ~n2399 & ~n2400 ;
  assign n2402 = ~x150 & ~x278 ;
  assign n2403 = x150 & x278 ;
  assign n2404 = ~n2402 & ~n2403 ;
  assign n2405 = ~n2401 & ~n2404 ;
  assign n2406 = n2401 & n2404 ;
  assign n2407 = ~n2405 & ~n2406 ;
  assign n2408 = ~x152 & ~x280 ;
  assign n2409 = x152 & x280 ;
  assign n2410 = ~n2408 & ~n2409 ;
  assign n2411 = ~n2407 & ~n2410 ;
  assign n2412 = n2407 & n2410 ;
  assign n2413 = ~n2411 & ~n2412 ;
  assign n2414 = ~x146 & ~x274 ;
  assign n2415 = x146 & x274 ;
  assign n2416 = ~n2414 & ~n2415 ;
  assign n2417 = ~n2413 & ~n2416 ;
  assign n2418 = n2413 & n2416 ;
  assign n2419 = ~n2417 & ~n2418 ;
  assign n2420 = ~x148 & ~x276 ;
  assign n2421 = x148 & x276 ;
  assign n2422 = ~n2420 & ~n2421 ;
  assign n2423 = ~x147 & ~x275 ;
  assign n2424 = x147 & x275 ;
  assign n2425 = ~n2423 & ~n2424 ;
  assign n2426 = ~n2422 & ~n2425 ;
  assign n2427 = n2422 & n2425 ;
  assign n2428 = ~n2426 & ~n2427 ;
  assign n2429 = ~x149 & ~x277 ;
  assign n2430 = x149 & x277 ;
  assign n2431 = ~n2429 & ~n2430 ;
  assign n2432 = ~n2428 & ~n2431 ;
  assign n2433 = n2428 & n2431 ;
  assign n2434 = ~n2432 & ~n2433 ;
  assign n2435 = n2419 & ~n2434 ;
  assign n2436 = ~n2417 & ~n2435 ;
  assign n2437 = ~n2406 & ~n2412 ;
  assign n2438 = ~n2436 & n2437 ;
  assign n2439 = n2436 & ~n2437 ;
  assign n2440 = ~n2438 & ~n2439 ;
  assign n2441 = ~n2427 & ~n2433 ;
  assign n2442 = n2440 & n2441 ;
  assign n2443 = ~n2440 & ~n2441 ;
  assign n2444 = ~n2442 & ~n2443 ;
  assign n2445 = ~x158 & ~x286 ;
  assign n2446 = x158 & x286 ;
  assign n2447 = ~n2445 & ~n2446 ;
  assign n2448 = ~x157 & ~x285 ;
  assign n2449 = x157 & x285 ;
  assign n2450 = ~n2448 & ~n2449 ;
  assign n2451 = n2447 & n2450 ;
  assign n2452 = ~n2447 & ~n2450 ;
  assign n2453 = ~n2451 & ~n2452 ;
  assign n2454 = ~x159 & ~x287 ;
  assign n2455 = x159 & x287 ;
  assign n2456 = ~n2454 & ~n2455 ;
  assign n2457 = ~n2453 & ~n2456 ;
  assign n2458 = n2453 & n2456 ;
  assign n2459 = ~n2457 & ~n2458 ;
  assign n2460 = ~x153 & ~x281 ;
  assign n2461 = x153 & x281 ;
  assign n2462 = ~n2460 & ~n2461 ;
  assign n2463 = ~n2459 & ~n2462 ;
  assign n2464 = n2459 & n2462 ;
  assign n2465 = ~n2463 & ~n2464 ;
  assign n2466 = ~x155 & ~x283 ;
  assign n2467 = x155 & x283 ;
  assign n2468 = ~n2466 & ~n2467 ;
  assign n2469 = ~x154 & ~x282 ;
  assign n2470 = x154 & x282 ;
  assign n2471 = ~n2469 & ~n2470 ;
  assign n2472 = ~n2468 & ~n2471 ;
  assign n2473 = n2468 & n2471 ;
  assign n2474 = ~n2472 & ~n2473 ;
  assign n2475 = ~x156 & ~x284 ;
  assign n2476 = x156 & x284 ;
  assign n2477 = ~n2475 & ~n2476 ;
  assign n2478 = ~n2474 & ~n2477 ;
  assign n2479 = n2474 & n2477 ;
  assign n2480 = ~n2478 & ~n2479 ;
  assign n2481 = n2465 & ~n2480 ;
  assign n2482 = ~n2463 & ~n2481 ;
  assign n2483 = ~n2451 & ~n2458 ;
  assign n2484 = ~n2482 & n2483 ;
  assign n2485 = n2482 & ~n2483 ;
  assign n2486 = ~n2484 & ~n2485 ;
  assign n2487 = ~n2473 & ~n2479 ;
  assign n2488 = n2486 & n2487 ;
  assign n2489 = ~n2486 & ~n2487 ;
  assign n2490 = ~n2488 & ~n2489 ;
  assign n2491 = ~n2465 & n2480 ;
  assign n2492 = ~n2481 & ~n2491 ;
  assign n2493 = ~x145 & ~x273 ;
  assign n2494 = x145 & x273 ;
  assign n2495 = ~n2493 & ~n2494 ;
  assign n2496 = n2492 & ~n2495 ;
  assign n2497 = ~n2419 & n2434 ;
  assign n2498 = ~n2435 & ~n2497 ;
  assign n2499 = ~n2492 & n2495 ;
  assign n2500 = ~n2496 & ~n2499 ;
  assign n2501 = n2498 & n2500 ;
  assign n2502 = ~n2496 & ~n2501 ;
  assign n2503 = n2490 & ~n2502 ;
  assign n2504 = ~n2490 & n2502 ;
  assign n2505 = ~n2503 & ~n2504 ;
  assign n2506 = n2444 & n2505 ;
  assign n2507 = ~n2444 & ~n2505 ;
  assign n2508 = ~n2506 & ~n2507 ;
  assign n2509 = ~n2498 & ~n2500 ;
  assign n2510 = ~n2501 & ~n2509 ;
  assign n2511 = ~x129 & ~x257 ;
  assign n2512 = x129 & x257 ;
  assign n2513 = ~n2511 & ~n2512 ;
  assign n2514 = n2510 & ~n2513 ;
  assign n2515 = ~n2388 & ~n2390 ;
  assign n2516 = ~n2391 & ~n2515 ;
  assign n2517 = ~n2510 & n2513 ;
  assign n2518 = ~n2514 & ~n2517 ;
  assign n2519 = n2516 & n2518 ;
  assign n2520 = ~n2514 & ~n2519 ;
  assign n2521 = n2508 & ~n2520 ;
  assign n2522 = ~n2508 & n2520 ;
  assign n2523 = ~n2521 & ~n2522 ;
  assign n2524 = n2398 & n2523 ;
  assign n2525 = ~n2398 & ~n2523 ;
  assign n2526 = ~n2524 & ~n2525 ;
  assign n2527 = ~n2516 & ~n2518 ;
  assign n2528 = ~n2519 & ~n2527 ;
  assign n2529 = ~x128 & ~x256 ;
  assign n2530 = x128 & x256 ;
  assign n2531 = ~n2529 & ~n2530 ;
  assign n2532 = ~n2528 & n2531 ;
  assign n2533 = ~n2526 & n2532 ;
  assign n2534 = ~n2374 & ~n2378 ;
  assign n2535 = ~n2393 & ~n2396 ;
  assign n2536 = ~n2534 & ~n2535 ;
  assign n2537 = n2534 & n2535 ;
  assign n2538 = ~n2536 & ~n2537 ;
  assign n2539 = ~n2328 & ~n2332 ;
  assign n2540 = n2538 & ~n2539 ;
  assign n2541 = ~n2538 & n2539 ;
  assign n2542 = ~n2540 & ~n2541 ;
  assign n2543 = ~n2484 & ~n2488 ;
  assign n2544 = ~n2503 & ~n2506 ;
  assign n2545 = ~n2543 & ~n2544 ;
  assign n2546 = n2543 & n2544 ;
  assign n2547 = ~n2545 & ~n2546 ;
  assign n2548 = ~n2438 & ~n2442 ;
  assign n2549 = n2547 & ~n2548 ;
  assign n2550 = ~n2547 & n2548 ;
  assign n2551 = ~n2549 & ~n2550 ;
  assign n2552 = ~n2521 & ~n2524 ;
  assign n2553 = n2551 & ~n2552 ;
  assign n2554 = ~n2551 & n2552 ;
  assign n2555 = ~n2553 & ~n2554 ;
  assign n2556 = n2542 & n2555 ;
  assign n2557 = ~n2542 & ~n2555 ;
  assign n2558 = ~n2556 & ~n2557 ;
  assign n2559 = n2533 & ~n2558 ;
  assign n2560 = ~n2545 & ~n2549 ;
  assign n2561 = ~n2553 & ~n2556 ;
  assign n2562 = ~n2560 & ~n2561 ;
  assign n2563 = n2560 & n2561 ;
  assign n2564 = ~n2562 & ~n2563 ;
  assign n2565 = ~n2536 & ~n2540 ;
  assign n2566 = n2564 & ~n2565 ;
  assign n2567 = ~n2564 & n2565 ;
  assign n2568 = ~n2566 & ~n2567 ;
  assign n2569 = n2559 & ~n2568 ;
  assign n2570 = ~n2562 & ~n2566 ;
  assign n2571 = n2569 & n2570 ;
  assign n2572 = ~n2288 & n2571 ;
  assign n2573 = n1703 & n2286 ;
  assign n2574 = ~n2571 & n2573 ;
  assign n2575 = ~n2572 & ~n2574 ;
  assign n2576 = n1420 & ~n2575 ;
  assign n2577 = n2571 & n2573 ;
  assign n2578 = ~n2576 & ~n2577 ;
  assign n2579 = n1137 & ~n2578 ;
  assign n2580 = n2576 & n2577 ;
  assign n2581 = ~n1137 & n2580 ;
  assign n2582 = ~n2579 & ~n2581 ;
  assign n2583 = n854 & ~n2582 ;
  assign n2584 = n1137 & n2580 ;
  assign n2585 = ~n854 & n2584 ;
  assign n2586 = ~n2583 & ~n2585 ;
  assign n2587 = n571 & ~n2586 ;
  assign n2588 = n854 & n2584 ;
  assign n2589 = ~n2587 & n2588 ;
  assign n2590 = ~n1980 & ~n1984 ;
  assign n2591 = ~n1985 & ~n2590 ;
  assign n2592 = n1993 & ~n2283 ;
  assign n2593 = n2262 & ~n2280 ;
  assign n2594 = ~n2281 & ~n2593 ;
  assign n2595 = n1972 & ~n1990 ;
  assign n2596 = ~n1991 & ~n2595 ;
  assign n2597 = n2594 & ~n2596 ;
  assign n2598 = ~n1985 & ~n1989 ;
  assign n2599 = ~n1990 & ~n2598 ;
  assign n2600 = ~n2275 & ~n2279 ;
  assign n2601 = ~n2280 & ~n2600 ;
  assign n2602 = ~n2599 & n2601 ;
  assign n2603 = n2599 & ~n2601 ;
  assign n2604 = ~n2270 & ~n2274 ;
  assign n2605 = ~n2275 & ~n2604 ;
  assign n2606 = ~n2591 & n2605 ;
  assign n2607 = ~n2274 & n2591 ;
  assign n2608 = ~n2265 & n2269 ;
  assign n2609 = ~n2270 & ~n2608 ;
  assign n2610 = ~n1975 & n1979 ;
  assign n2611 = ~n1980 & ~n2610 ;
  assign n2612 = n2609 & ~n2611 ;
  assign n2613 = ~n2607 & n2612 ;
  assign n2614 = ~n2606 & ~n2613 ;
  assign n2615 = ~n2603 & ~n2614 ;
  assign n2616 = ~n2602 & ~n2615 ;
  assign n2617 = ~n2597 & n2616 ;
  assign n2618 = ~n1991 & ~n1992 ;
  assign n2619 = ~n1993 & ~n2618 ;
  assign n2620 = ~n2281 & ~n2282 ;
  assign n2621 = ~n2283 & ~n2620 ;
  assign n2622 = n2619 & ~n2621 ;
  assign n2623 = ~n2594 & n2596 ;
  assign n2624 = ~n2622 & ~n2623 ;
  assign n2625 = ~n2617 & n2624 ;
  assign n2626 = ~n2619 & n2621 ;
  assign n2627 = ~n1993 & n2283 ;
  assign n2628 = ~n2626 & ~n2627 ;
  assign n2629 = ~n2625 & n2628 ;
  assign n2630 = ~n2592 & ~n2629 ;
  assign n2631 = ~n2591 & ~n2630 ;
  assign n2632 = ~n2605 & n2630 ;
  assign n2633 = ~n2631 & ~n2632 ;
  assign n2634 = n1683 & ~n1689 ;
  assign n2635 = ~n1690 & ~n2634 ;
  assign n2636 = ~n2633 & n2635 ;
  assign n2637 = n1685 & ~n1688 ;
  assign n2638 = ~n1689 & ~n2637 ;
  assign n2639 = ~n2611 & ~n2630 ;
  assign n2640 = ~n2609 & n2630 ;
  assign n2641 = ~n2639 & ~n2640 ;
  assign n2642 = n2638 & ~n2641 ;
  assign n2643 = ~n2636 & ~n2642 ;
  assign n2644 = n1683 & n2633 ;
  assign n2645 = n1681 & ~n1690 ;
  assign n2646 = ~n1691 & ~n2645 ;
  assign n2647 = ~n2599 & ~n2630 ;
  assign n2648 = ~n2601 & n2630 ;
  assign n2649 = ~n2647 & ~n2648 ;
  assign n2650 = ~n2646 & n2649 ;
  assign n2651 = ~n2644 & ~n2650 ;
  assign n2652 = ~n2643 & n2651 ;
  assign n2653 = ~n1691 & n1700 ;
  assign n2654 = ~n1701 & ~n2653 ;
  assign n2655 = n2597 & ~n2630 ;
  assign n2656 = ~n2597 & ~n2623 ;
  assign n2657 = ~n2630 & ~n2656 ;
  assign n2658 = ~n2594 & ~n2657 ;
  assign n2659 = ~n2655 & ~n2658 ;
  assign n2660 = n2654 & ~n2659 ;
  assign n2661 = n2646 & ~n2649 ;
  assign n2662 = ~n2660 & ~n2661 ;
  assign n2663 = ~n2652 & n2662 ;
  assign n2664 = ~n2654 & n2659 ;
  assign n2665 = ~n1701 & ~n1702 ;
  assign n2666 = ~n1703 & ~n2665 ;
  assign n2667 = ~n2622 & ~n2626 ;
  assign n2668 = ~n2630 & ~n2667 ;
  assign n2669 = ~n2621 & ~n2668 ;
  assign n2670 = n2592 & ~n2620 ;
  assign n2671 = ~n2669 & ~n2670 ;
  assign n2672 = ~n2666 & n2671 ;
  assign n2673 = ~n1703 & ~n2284 ;
  assign n2674 = ~n2672 & ~n2673 ;
  assign n2675 = ~n2664 & n2674 ;
  assign n2676 = ~n2663 & n2675 ;
  assign n2677 = ~n1703 & n2671 ;
  assign n2678 = n2284 & ~n2665 ;
  assign n2679 = ~n2677 & n2678 ;
  assign n2680 = ~n2676 & ~n2679 ;
  assign n2681 = n2633 & ~n2680 ;
  assign n2682 = n2635 & n2680 ;
  assign n2683 = ~n2681 & ~n2682 ;
  assign n2684 = n2285 & ~n2286 ;
  assign n2685 = n2605 & ~n2630 ;
  assign n2686 = n2591 & n2630 ;
  assign n2687 = ~n2685 & ~n2686 ;
  assign n2688 = n2683 & ~n2687 ;
  assign n2689 = ~n2638 & n2680 ;
  assign n2690 = ~n2641 & ~n2680 ;
  assign n2691 = ~n2689 & ~n2690 ;
  assign n2692 = n2609 & ~n2630 ;
  assign n2693 = n2611 & n2630 ;
  assign n2694 = ~n2692 & ~n2693 ;
  assign n2695 = n2691 & n2694 ;
  assign n2696 = ~n2688 & n2695 ;
  assign n2697 = ~n2683 & n2687 ;
  assign n2698 = n2601 & ~n2630 ;
  assign n2699 = n2599 & n2630 ;
  assign n2700 = ~n2698 & ~n2699 ;
  assign n2701 = n2646 & n2680 ;
  assign n2702 = n2649 & ~n2680 ;
  assign n2703 = ~n2701 & ~n2702 ;
  assign n2704 = n2700 & ~n2703 ;
  assign n2705 = ~n2697 & ~n2704 ;
  assign n2706 = ~n2696 & n2705 ;
  assign n2707 = n2596 & ~n2657 ;
  assign n2708 = ~n2655 & ~n2707 ;
  assign n2709 = n2654 & n2680 ;
  assign n2710 = n2659 & ~n2680 ;
  assign n2711 = ~n2709 & ~n2710 ;
  assign n2712 = ~n2708 & n2711 ;
  assign n2713 = ~n2700 & n2703 ;
  assign n2714 = ~n2712 & ~n2713 ;
  assign n2715 = ~n2706 & n2714 ;
  assign n2716 = n2708 & ~n2711 ;
  assign n2717 = n2619 & ~n2668 ;
  assign n2718 = ~n2670 & ~n2717 ;
  assign n2719 = n2666 & n2680 ;
  assign n2720 = n2671 & ~n2680 ;
  assign n2721 = ~n2719 & ~n2720 ;
  assign n2722 = n2718 & ~n2721 ;
  assign n2723 = ~n2716 & ~n2722 ;
  assign n2724 = ~n2715 & n2723 ;
  assign n2725 = ~n2718 & n2721 ;
  assign n2726 = ~n2287 & ~n2725 ;
  assign n2727 = ~n2724 & n2726 ;
  assign n2728 = ~n2684 & ~n2727 ;
  assign n2729 = ~n2683 & n2728 ;
  assign n2730 = ~n2687 & ~n2728 ;
  assign n2731 = ~n2729 & ~n2730 ;
  assign n2732 = n2572 & ~n2573 ;
  assign n2733 = ~n2687 & n2728 ;
  assign n2734 = ~n2683 & ~n2728 ;
  assign n2735 = ~n2733 & ~n2734 ;
  assign n2736 = n2528 & ~n2531 ;
  assign n2737 = ~n2532 & ~n2736 ;
  assign n2738 = ~n2694 & n2728 ;
  assign n2739 = n2691 & ~n2728 ;
  assign n2740 = ~n2738 & ~n2739 ;
  assign n2741 = n2737 & n2740 ;
  assign n2742 = ~n2526 & n2741 ;
  assign n2743 = ~n2735 & ~n2742 ;
  assign n2744 = n2526 & ~n2532 ;
  assign n2745 = ~n2533 & ~n2744 ;
  assign n2746 = ~n2741 & ~n2745 ;
  assign n2747 = ~n2533 & n2558 ;
  assign n2748 = ~n2559 & ~n2747 ;
  assign n2749 = ~n2700 & n2728 ;
  assign n2750 = ~n2703 & ~n2728 ;
  assign n2751 = ~n2749 & ~n2750 ;
  assign n2752 = ~n2748 & ~n2751 ;
  assign n2753 = ~n2746 & ~n2752 ;
  assign n2754 = ~n2743 & n2753 ;
  assign n2755 = n2748 & n2751 ;
  assign n2756 = ~n2559 & n2568 ;
  assign n2757 = ~n2569 & ~n2756 ;
  assign n2758 = n2716 & n2728 ;
  assign n2759 = ~n2712 & ~n2716 ;
  assign n2760 = n2728 & ~n2759 ;
  assign n2761 = n2711 & ~n2760 ;
  assign n2762 = ~n2758 & ~n2761 ;
  assign n2763 = n2757 & ~n2762 ;
  assign n2764 = ~n2755 & ~n2763 ;
  assign n2765 = ~n2754 & n2764 ;
  assign n2766 = ~n2569 & ~n2570 ;
  assign n2767 = ~n2571 & ~n2766 ;
  assign n2768 = n2722 & n2728 ;
  assign n2769 = ~n2722 & ~n2725 ;
  assign n2770 = n2728 & ~n2769 ;
  assign n2771 = n2721 & ~n2770 ;
  assign n2772 = ~n2768 & ~n2771 ;
  assign n2773 = ~n2767 & n2772 ;
  assign n2774 = ~n2757 & n2762 ;
  assign n2775 = ~n2288 & ~n2571 ;
  assign n2776 = ~n2774 & ~n2775 ;
  assign n2777 = ~n2773 & n2776 ;
  assign n2778 = ~n2765 & n2777 ;
  assign n2779 = ~n2571 & n2772 ;
  assign n2780 = n2288 & ~n2766 ;
  assign n2781 = ~n2779 & n2780 ;
  assign n2782 = ~n2778 & ~n2781 ;
  assign n2783 = ~n2735 & ~n2782 ;
  assign n2784 = n2745 & n2782 ;
  assign n2785 = ~n2783 & ~n2784 ;
  assign n2786 = ~n2731 & n2785 ;
  assign n2787 = ~n2691 & n2728 ;
  assign n2788 = n2694 & ~n2728 ;
  assign n2789 = ~n2787 & ~n2788 ;
  assign n2790 = ~n2737 & n2782 ;
  assign n2791 = n2740 & ~n2782 ;
  assign n2792 = ~n2790 & ~n2791 ;
  assign n2793 = ~n2789 & n2792 ;
  assign n2794 = ~n2786 & n2793 ;
  assign n2795 = n2731 & ~n2785 ;
  assign n2796 = n2700 & ~n2728 ;
  assign n2797 = n2703 & n2728 ;
  assign n2798 = ~n2796 & ~n2797 ;
  assign n2799 = ~n2751 & ~n2782 ;
  assign n2800 = n2748 & n2782 ;
  assign n2801 = ~n2799 & ~n2800 ;
  assign n2802 = ~n2798 & ~n2801 ;
  assign n2803 = ~n2795 & ~n2802 ;
  assign n2804 = ~n2794 & n2803 ;
  assign n2805 = ~n2708 & ~n2760 ;
  assign n2806 = ~n2758 & ~n2805 ;
  assign n2807 = n2757 & n2782 ;
  assign n2808 = n2762 & ~n2782 ;
  assign n2809 = ~n2807 & ~n2808 ;
  assign n2810 = ~n2806 & n2809 ;
  assign n2811 = n2798 & n2801 ;
  assign n2812 = ~n2810 & ~n2811 ;
  assign n2813 = ~n2804 & n2812 ;
  assign n2814 = n2806 & ~n2809 ;
  assign n2815 = ~n2718 & ~n2770 ;
  assign n2816 = ~n2768 & ~n2815 ;
  assign n2817 = n2767 & n2782 ;
  assign n2818 = n2772 & ~n2782 ;
  assign n2819 = ~n2817 & ~n2818 ;
  assign n2820 = n2816 & ~n2819 ;
  assign n2821 = ~n2814 & ~n2820 ;
  assign n2822 = ~n2813 & n2821 ;
  assign n2823 = ~n2816 & n2819 ;
  assign n2824 = ~n2574 & ~n2823 ;
  assign n2825 = ~n2822 & n2824 ;
  assign n2826 = ~n2732 & ~n2825 ;
  assign n2827 = n2731 & ~n2826 ;
  assign n2828 = n2785 & n2826 ;
  assign n2829 = ~n2827 & ~n2828 ;
  assign n2830 = n2576 & ~n2577 ;
  assign n2831 = ~n2785 & ~n2826 ;
  assign n2832 = ~n2731 & n2826 ;
  assign n2833 = ~n2831 & ~n2832 ;
  assign n2834 = n1400 & ~n1406 ;
  assign n2835 = ~n1407 & ~n2834 ;
  assign n2836 = n2833 & n2835 ;
  assign n2837 = n1402 & ~n1405 ;
  assign n2838 = ~n1406 & ~n2837 ;
  assign n2839 = ~n2789 & n2826 ;
  assign n2840 = ~n2792 & ~n2826 ;
  assign n2841 = ~n2839 & ~n2840 ;
  assign n2842 = n2838 & ~n2841 ;
  assign n2843 = ~n2836 & ~n2842 ;
  assign n2844 = n1400 & ~n2833 ;
  assign n2845 = n1398 & ~n1407 ;
  assign n2846 = ~n1408 & ~n2845 ;
  assign n2847 = ~n2798 & n2826 ;
  assign n2848 = n2801 & ~n2826 ;
  assign n2849 = ~n2847 & ~n2848 ;
  assign n2850 = ~n2846 & n2849 ;
  assign n2851 = ~n2844 & ~n2850 ;
  assign n2852 = ~n2843 & n2851 ;
  assign n2853 = ~n1408 & n1417 ;
  assign n2854 = ~n1418 & ~n2853 ;
  assign n2855 = n2814 & n2826 ;
  assign n2856 = ~n2810 & ~n2814 ;
  assign n2857 = n2826 & ~n2856 ;
  assign n2858 = n2809 & ~n2857 ;
  assign n2859 = ~n2855 & ~n2858 ;
  assign n2860 = n2854 & ~n2859 ;
  assign n2861 = n2846 & ~n2849 ;
  assign n2862 = ~n2860 & ~n2861 ;
  assign n2863 = ~n2852 & n2862 ;
  assign n2864 = ~n2854 & n2859 ;
  assign n2865 = ~n1418 & ~n1419 ;
  assign n2866 = ~n1420 & ~n2865 ;
  assign n2867 = n2820 & n2826 ;
  assign n2868 = ~n2820 & ~n2823 ;
  assign n2869 = n2826 & ~n2868 ;
  assign n2870 = n2819 & ~n2869 ;
  assign n2871 = ~n2867 & ~n2870 ;
  assign n2872 = ~n2866 & n2871 ;
  assign n2873 = ~n1420 & ~n2575 ;
  assign n2874 = ~n2872 & ~n2873 ;
  assign n2875 = ~n2864 & n2874 ;
  assign n2876 = ~n2863 & n2875 ;
  assign n2877 = ~n1420 & n2871 ;
  assign n2878 = n2575 & ~n2865 ;
  assign n2879 = ~n2877 & n2878 ;
  assign n2880 = ~n2876 & ~n2879 ;
  assign n2881 = ~n2833 & ~n2880 ;
  assign n2882 = n2835 & n2880 ;
  assign n2883 = ~n2881 & ~n2882 ;
  assign n2884 = n2829 & n2883 ;
  assign n2885 = n2789 & ~n2826 ;
  assign n2886 = n2792 & n2826 ;
  assign n2887 = ~n2885 & ~n2886 ;
  assign n2888 = ~n2838 & n2880 ;
  assign n2889 = ~n2841 & ~n2880 ;
  assign n2890 = ~n2888 & ~n2889 ;
  assign n2891 = n2887 & n2890 ;
  assign n2892 = ~n2884 & n2891 ;
  assign n2893 = ~n2829 & ~n2883 ;
  assign n2894 = ~n2801 & n2826 ;
  assign n2895 = n2798 & ~n2826 ;
  assign n2896 = ~n2894 & ~n2895 ;
  assign n2897 = n2846 & n2880 ;
  assign n2898 = n2849 & ~n2880 ;
  assign n2899 = ~n2897 & ~n2898 ;
  assign n2900 = n2896 & ~n2899 ;
  assign n2901 = ~n2893 & ~n2900 ;
  assign n2902 = ~n2892 & n2901 ;
  assign n2903 = ~n2806 & ~n2857 ;
  assign n2904 = ~n2855 & ~n2903 ;
  assign n2905 = n2854 & n2880 ;
  assign n2906 = n2859 & ~n2880 ;
  assign n2907 = ~n2905 & ~n2906 ;
  assign n2908 = ~n2904 & n2907 ;
  assign n2909 = ~n2896 & n2899 ;
  assign n2910 = ~n2908 & ~n2909 ;
  assign n2911 = ~n2902 & n2910 ;
  assign n2912 = n2904 & ~n2907 ;
  assign n2913 = ~n2816 & ~n2869 ;
  assign n2914 = ~n2867 & ~n2913 ;
  assign n2915 = n2866 & n2880 ;
  assign n2916 = n2871 & ~n2880 ;
  assign n2917 = ~n2915 & ~n2916 ;
  assign n2918 = n2914 & ~n2917 ;
  assign n2919 = ~n2912 & ~n2918 ;
  assign n2920 = ~n2911 & n2919 ;
  assign n2921 = ~n2914 & n2917 ;
  assign n2922 = ~n2576 & n2577 ;
  assign n2923 = ~n2921 & ~n2922 ;
  assign n2924 = ~n2920 & n2923 ;
  assign n2925 = ~n2830 & ~n2924 ;
  assign n2926 = ~n2829 & ~n2925 ;
  assign n2927 = n2883 & n2925 ;
  assign n2928 = ~n2926 & ~n2927 ;
  assign n2929 = n2579 & ~n2580 ;
  assign n2930 = ~n2829 & n2925 ;
  assign n2931 = n2883 & ~n2925 ;
  assign n2932 = ~n2930 & ~n2931 ;
  assign n2933 = n1117 & ~n1123 ;
  assign n2934 = ~n1124 & ~n2933 ;
  assign n2935 = ~n2932 & n2934 ;
  assign n2936 = n1119 & ~n1122 ;
  assign n2937 = ~n1123 & ~n2936 ;
  assign n2938 = ~n2887 & n2925 ;
  assign n2939 = n2890 & ~n2925 ;
  assign n2940 = ~n2938 & ~n2939 ;
  assign n2941 = n2937 & n2940 ;
  assign n2942 = ~n2935 & ~n2941 ;
  assign n2943 = n1117 & n2932 ;
  assign n2944 = n1115 & ~n1124 ;
  assign n2945 = ~n1125 & ~n2944 ;
  assign n2946 = ~n2896 & n2925 ;
  assign n2947 = ~n2899 & ~n2925 ;
  assign n2948 = ~n2946 & ~n2947 ;
  assign n2949 = ~n2945 & ~n2948 ;
  assign n2950 = ~n2943 & ~n2949 ;
  assign n2951 = ~n2942 & n2950 ;
  assign n2952 = ~n1125 & n1134 ;
  assign n2953 = ~n1135 & ~n2952 ;
  assign n2954 = n2912 & n2925 ;
  assign n2955 = ~n2908 & ~n2912 ;
  assign n2956 = n2925 & ~n2955 ;
  assign n2957 = n2907 & ~n2956 ;
  assign n2958 = ~n2954 & ~n2957 ;
  assign n2959 = n2953 & ~n2958 ;
  assign n2960 = n2945 & n2948 ;
  assign n2961 = ~n2959 & ~n2960 ;
  assign n2962 = ~n2951 & n2961 ;
  assign n2963 = ~n2953 & n2958 ;
  assign n2964 = ~n1135 & ~n1136 ;
  assign n2965 = ~n1137 & ~n2964 ;
  assign n2966 = n2918 & n2925 ;
  assign n2967 = ~n2918 & ~n2921 ;
  assign n2968 = n2925 & ~n2967 ;
  assign n2969 = n2917 & ~n2968 ;
  assign n2970 = ~n2966 & ~n2969 ;
  assign n2971 = ~n2965 & n2970 ;
  assign n2972 = ~n1137 & ~n2578 ;
  assign n2973 = ~n2971 & ~n2972 ;
  assign n2974 = ~n2963 & n2973 ;
  assign n2975 = ~n2962 & n2974 ;
  assign n2976 = ~n1137 & n2970 ;
  assign n2977 = n2578 & ~n2964 ;
  assign n2978 = ~n2976 & n2977 ;
  assign n2979 = ~n2975 & ~n2978 ;
  assign n2980 = n2932 & ~n2979 ;
  assign n2981 = n2934 & n2979 ;
  assign n2982 = ~n2980 & ~n2981 ;
  assign n2983 = n2928 & n2982 ;
  assign n2984 = n2887 & ~n2925 ;
  assign n2985 = ~n2890 & n2925 ;
  assign n2986 = ~n2984 & ~n2985 ;
  assign n2987 = ~n2937 & n2979 ;
  assign n2988 = n2940 & ~n2979 ;
  assign n2989 = ~n2987 & ~n2988 ;
  assign n2990 = ~n2986 & n2989 ;
  assign n2991 = ~n2983 & n2990 ;
  assign n2992 = ~n2928 & ~n2982 ;
  assign n2993 = n2896 & ~n2925 ;
  assign n2994 = n2899 & n2925 ;
  assign n2995 = ~n2993 & ~n2994 ;
  assign n2996 = ~n2948 & ~n2979 ;
  assign n2997 = n2945 & n2979 ;
  assign n2998 = ~n2996 & ~n2997 ;
  assign n2999 = ~n2995 & ~n2998 ;
  assign n3000 = ~n2992 & ~n2999 ;
  assign n3001 = ~n2991 & n3000 ;
  assign n3002 = ~n2904 & ~n2956 ;
  assign n3003 = ~n2954 & ~n3002 ;
  assign n3004 = n2953 & n2979 ;
  assign n3005 = n2958 & ~n2979 ;
  assign n3006 = ~n3004 & ~n3005 ;
  assign n3007 = ~n3003 & n3006 ;
  assign n3008 = n2995 & n2998 ;
  assign n3009 = ~n3007 & ~n3008 ;
  assign n3010 = ~n3001 & n3009 ;
  assign n3011 = n3003 & ~n3006 ;
  assign n3012 = ~n2914 & ~n2968 ;
  assign n3013 = ~n2966 & ~n3012 ;
  assign n3014 = n2965 & n2979 ;
  assign n3015 = n2970 & ~n2979 ;
  assign n3016 = ~n3014 & ~n3015 ;
  assign n3017 = n3013 & ~n3016 ;
  assign n3018 = ~n3011 & ~n3017 ;
  assign n3019 = ~n3010 & n3018 ;
  assign n3020 = ~n3013 & n3016 ;
  assign n3021 = ~n2581 & ~n3020 ;
  assign n3022 = ~n3019 & n3021 ;
  assign n3023 = ~n2929 & ~n3022 ;
  assign n3024 = ~n2928 & n3023 ;
  assign n3025 = n2982 & ~n3023 ;
  assign n3026 = ~n3024 & ~n3025 ;
  assign n3027 = n834 & ~n840 ;
  assign n3028 = ~n841 & ~n3027 ;
  assign n3029 = ~n3026 & n3028 ;
  assign n3030 = n836 & ~n839 ;
  assign n3031 = ~n840 & ~n3030 ;
  assign n3032 = n2989 & ~n3023 ;
  assign n3033 = n2986 & n3023 ;
  assign n3034 = ~n3032 & ~n3033 ;
  assign n3035 = n3031 & n3034 ;
  assign n3036 = ~n3029 & ~n3035 ;
  assign n3037 = n834 & n3026 ;
  assign n3038 = n832 & ~n841 ;
  assign n3039 = ~n842 & ~n3038 ;
  assign n3040 = ~n2995 & n3023 ;
  assign n3041 = n2998 & ~n3023 ;
  assign n3042 = ~n3040 & ~n3041 ;
  assign n3043 = ~n3039 & n3042 ;
  assign n3044 = ~n3037 & ~n3043 ;
  assign n3045 = ~n3036 & n3044 ;
  assign n3046 = ~n842 & n851 ;
  assign n3047 = ~n852 & ~n3046 ;
  assign n3048 = n3011 & n3023 ;
  assign n3049 = ~n3007 & ~n3011 ;
  assign n3050 = n3023 & ~n3049 ;
  assign n3051 = n3006 & ~n3050 ;
  assign n3052 = ~n3048 & ~n3051 ;
  assign n3053 = n3047 & ~n3052 ;
  assign n3054 = n3039 & ~n3042 ;
  assign n3055 = ~n3053 & ~n3054 ;
  assign n3056 = ~n3045 & n3055 ;
  assign n3057 = ~n3047 & n3052 ;
  assign n3058 = ~n852 & ~n853 ;
  assign n3059 = ~n854 & ~n3058 ;
  assign n3060 = n3017 & n3023 ;
  assign n3061 = ~n3017 & ~n3020 ;
  assign n3062 = n3023 & ~n3061 ;
  assign n3063 = n3016 & ~n3062 ;
  assign n3064 = ~n3060 & ~n3063 ;
  assign n3065 = ~n3059 & n3064 ;
  assign n3066 = ~n854 & ~n2582 ;
  assign n3067 = ~n3065 & ~n3066 ;
  assign n3068 = ~n3057 & n3067 ;
  assign n3069 = ~n3056 & n3068 ;
  assign n3070 = ~n854 & n3064 ;
  assign n3071 = n2582 & ~n3058 ;
  assign n3072 = ~n3070 & n3071 ;
  assign n3073 = ~n3069 & ~n3072 ;
  assign n3074 = n3026 & ~n3073 ;
  assign n3075 = n3028 & n3073 ;
  assign n3076 = ~n3074 & ~n3075 ;
  assign n3077 = n2583 & ~n2584 ;
  assign n3078 = ~n2928 & ~n3023 ;
  assign n3079 = n2982 & n3023 ;
  assign n3080 = ~n3078 & ~n3079 ;
  assign n3081 = n3076 & n3080 ;
  assign n3082 = ~n3031 & n3073 ;
  assign n3083 = n3034 & ~n3073 ;
  assign n3084 = ~n3082 & ~n3083 ;
  assign n3085 = ~n2986 & ~n3023 ;
  assign n3086 = ~n2989 & n3023 ;
  assign n3087 = ~n3085 & ~n3086 ;
  assign n3088 = n3084 & ~n3087 ;
  assign n3089 = ~n3081 & n3088 ;
  assign n3090 = ~n3076 & ~n3080 ;
  assign n3091 = ~n2998 & n3023 ;
  assign n3092 = n2995 & ~n3023 ;
  assign n3093 = ~n3091 & ~n3092 ;
  assign n3094 = n3039 & n3073 ;
  assign n3095 = n3042 & ~n3073 ;
  assign n3096 = ~n3094 & ~n3095 ;
  assign n3097 = n3093 & ~n3096 ;
  assign n3098 = ~n3090 & ~n3097 ;
  assign n3099 = ~n3089 & n3098 ;
  assign n3100 = ~n3003 & ~n3050 ;
  assign n3101 = ~n3048 & ~n3100 ;
  assign n3102 = n3047 & n3073 ;
  assign n3103 = n3052 & ~n3073 ;
  assign n3104 = ~n3102 & ~n3103 ;
  assign n3105 = ~n3101 & n3104 ;
  assign n3106 = ~n3093 & n3096 ;
  assign n3107 = ~n3105 & ~n3106 ;
  assign n3108 = ~n3099 & n3107 ;
  assign n3109 = n3101 & ~n3104 ;
  assign n3110 = ~n3013 & ~n3062 ;
  assign n3111 = ~n3060 & ~n3110 ;
  assign n3112 = n3059 & n3073 ;
  assign n3113 = n3064 & ~n3073 ;
  assign n3114 = ~n3112 & ~n3113 ;
  assign n3115 = n3111 & ~n3114 ;
  assign n3116 = ~n3109 & ~n3115 ;
  assign n3117 = ~n3108 & n3116 ;
  assign n3118 = ~n3111 & n3114 ;
  assign n3119 = ~n2585 & ~n3118 ;
  assign n3120 = ~n3117 & n3119 ;
  assign n3121 = ~n3077 & ~n3120 ;
  assign n3122 = ~n3076 & n3121 ;
  assign n3123 = n3080 & ~n3121 ;
  assign n3124 = ~n3122 & ~n3123 ;
  assign n3125 = ~n3087 & n3121 ;
  assign n3126 = ~n3084 & ~n3121 ;
  assign n3127 = ~n3125 & ~n3126 ;
  assign n3128 = n560 & ~n566 ;
  assign n3129 = ~n567 & ~n3128 ;
  assign n3130 = ~n3080 & n3121 ;
  assign n3131 = n3076 & ~n3121 ;
  assign n3132 = ~n3130 & ~n3131 ;
  assign n3133 = n3129 & ~n3132 ;
  assign n3134 = n562 & ~n565 ;
  assign n3135 = ~n566 & ~n3134 ;
  assign n3136 = ~n3127 & n3135 ;
  assign n3137 = ~n3133 & ~n3136 ;
  assign n3138 = n560 & n3132 ;
  assign n3139 = n558 & ~n567 ;
  assign n3140 = ~n568 & ~n3139 ;
  assign n3141 = ~n3093 & n3121 ;
  assign n3142 = ~n3096 & ~n3121 ;
  assign n3143 = ~n3141 & ~n3142 ;
  assign n3144 = ~n3140 & ~n3143 ;
  assign n3145 = ~n3138 & ~n3144 ;
  assign n3146 = ~n3137 & n3145 ;
  assign n3147 = n3109 & n3121 ;
  assign n3148 = ~n3105 & ~n3109 ;
  assign n3149 = n3121 & ~n3148 ;
  assign n3150 = n3104 & ~n3149 ;
  assign n3151 = ~n3147 & ~n3150 ;
  assign n3152 = n556 & ~n568 ;
  assign n3153 = ~n569 & ~n3152 ;
  assign n3154 = ~n3151 & n3153 ;
  assign n3155 = n3140 & n3143 ;
  assign n3156 = ~n3154 & ~n3155 ;
  assign n3157 = ~n3146 & n3156 ;
  assign n3158 = n3151 & ~n3153 ;
  assign n3159 = n3115 & n3121 ;
  assign n3160 = ~n3115 & ~n3118 ;
  assign n3161 = n3121 & ~n3160 ;
  assign n3162 = n3114 & ~n3161 ;
  assign n3163 = ~n3159 & ~n3162 ;
  assign n3164 = ~n569 & ~n570 ;
  assign n3165 = ~n571 & ~n3164 ;
  assign n3166 = n3163 & ~n3165 ;
  assign n3167 = ~n571 & ~n2586 ;
  assign n3168 = ~n3166 & ~n3167 ;
  assign n3169 = ~n3158 & n3168 ;
  assign n3170 = ~n3157 & n3169 ;
  assign n3171 = ~n571 & n3163 ;
  assign n3172 = n2586 & ~n3164 ;
  assign n3173 = ~n3171 & n3172 ;
  assign n3174 = ~n3170 & ~n3173 ;
  assign n3175 = ~n3127 & ~n3174 ;
  assign n3176 = ~n3135 & n3174 ;
  assign n3177 = n3084 & n3121 ;
  assign n3178 = n3087 & ~n3121 ;
  assign n3179 = ~n3177 & ~n3178 ;
  assign n3180 = ~n3176 & n3179 ;
  assign n3181 = ~n3175 & n3180 ;
  assign n3182 = ~n3129 & n3174 ;
  assign n3183 = ~n3132 & ~n3174 ;
  assign n3184 = ~n3182 & ~n3183 ;
  assign n3185 = n3181 & n3184 ;
  assign n3186 = ~n3124 & ~n3185 ;
  assign n3187 = ~n3096 & n3121 ;
  assign n3188 = ~n3093 & ~n3121 ;
  assign n3189 = ~n3187 & ~n3188 ;
  assign n3190 = ~n3143 & ~n3174 ;
  assign n3191 = n3140 & n3174 ;
  assign n3192 = ~n3190 & ~n3191 ;
  assign n3193 = ~n3189 & n3192 ;
  assign n3194 = ~n3181 & ~n3184 ;
  assign n3195 = ~n3193 & ~n3194 ;
  assign n3196 = ~n3186 & n3195 ;
  assign n3197 = ~n3101 & ~n3149 ;
  assign n3198 = ~n3147 & ~n3197 ;
  assign n3199 = ~n3151 & ~n3174 ;
  assign n3200 = ~n3153 & n3174 ;
  assign n3201 = ~n3199 & ~n3200 ;
  assign n3202 = n3198 & n3201 ;
  assign n3203 = n3189 & ~n3192 ;
  assign n3204 = ~n3202 & ~n3203 ;
  assign n3205 = ~n3196 & n3204 ;
  assign n3206 = ~n3111 & ~n3161 ;
  assign n3207 = ~n3159 & ~n3206 ;
  assign n3208 = n3163 & ~n3174 ;
  assign n3209 = n3165 & n3174 ;
  assign n3210 = ~n3208 & ~n3209 ;
  assign n3211 = ~n3207 & n3210 ;
  assign n3212 = ~n3198 & ~n3201 ;
  assign n3213 = ~n3211 & ~n3212 ;
  assign n3214 = ~n3205 & n3213 ;
  assign n3215 = n2587 & ~n2588 ;
  assign n3216 = n3207 & ~n3210 ;
  assign n3217 = ~n3215 & ~n3216 ;
  assign n3218 = ~n3214 & n3217 ;
  assign n3219 = ~n2589 & ~n3218 ;
  assign n3220 = x192 & ~n2630 ;
  assign n3221 = x224 & n2630 ;
  assign n3222 = ~n3220 & ~n3221 ;
  assign n3223 = ~n2728 & ~n3222 ;
  assign n3224 = ~x224 & ~n2630 ;
  assign n3225 = ~x192 & n2630 ;
  assign n3226 = ~n3224 & ~n3225 ;
  assign n3227 = ~n2680 & ~n3226 ;
  assign n3228 = ~x160 & n2680 ;
  assign n3229 = ~n3227 & ~n3228 ;
  assign n3230 = n2728 & n3229 ;
  assign n3231 = ~n3223 & ~n3230 ;
  assign n3232 = ~n2826 & ~n3231 ;
  assign n3233 = n2728 & ~n3222 ;
  assign n3234 = ~n2728 & n3229 ;
  assign n3235 = ~n3233 & ~n3234 ;
  assign n3236 = ~n2782 & ~n3235 ;
  assign n3237 = x128 & n2782 ;
  assign n3238 = ~n3236 & ~n3237 ;
  assign n3239 = n2826 & ~n3238 ;
  assign n3240 = ~n3232 & ~n3239 ;
  assign n3241 = ~n2925 & ~n3240 ;
  assign n3242 = n2826 & ~n3231 ;
  assign n3243 = ~n2826 & ~n3238 ;
  assign n3244 = ~n3242 & ~n3243 ;
  assign n3245 = ~n2880 & ~n3244 ;
  assign n3246 = x96 & n2880 ;
  assign n3247 = ~n3245 & ~n3246 ;
  assign n3248 = n2925 & ~n3247 ;
  assign n3249 = ~n3241 & ~n3248 ;
  assign n3250 = ~n3023 & ~n3249 ;
  assign n3251 = n2925 & ~n3240 ;
  assign n3252 = ~n2925 & ~n3247 ;
  assign n3253 = ~n3251 & ~n3252 ;
  assign n3254 = ~n2979 & ~n3253 ;
  assign n3255 = x64 & n2979 ;
  assign n3256 = ~n3254 & ~n3255 ;
  assign n3257 = n3023 & ~n3256 ;
  assign n3258 = ~n3250 & ~n3257 ;
  assign n3259 = ~n3121 & ~n3258 ;
  assign n3260 = n3023 & ~n3249 ;
  assign n3261 = ~n3023 & ~n3256 ;
  assign n3262 = ~n3260 & ~n3261 ;
  assign n3263 = ~n3073 & ~n3262 ;
  assign n3264 = x32 & n3073 ;
  assign n3265 = ~n3263 & ~n3264 ;
  assign n3266 = n3121 & ~n3265 ;
  assign n3267 = ~n3259 & ~n3266 ;
  assign n3268 = n3219 & ~n3267 ;
  assign n3269 = n3121 & ~n3258 ;
  assign n3270 = ~n3121 & ~n3265 ;
  assign n3271 = ~n3269 & ~n3270 ;
  assign n3272 = ~n3174 & ~n3271 ;
  assign n3273 = x0 & n3174 ;
  assign n3274 = ~n3272 & ~n3273 ;
  assign n3275 = ~n3219 & ~n3274 ;
  assign n3276 = ~n3268 & ~n3275 ;
  assign n3277 = x193 & ~n2630 ;
  assign n3278 = x225 & n2630 ;
  assign n3279 = ~n3277 & ~n3278 ;
  assign n3280 = ~n2728 & ~n3279 ;
  assign n3281 = ~x225 & ~n2630 ;
  assign n3282 = ~x193 & n2630 ;
  assign n3283 = ~n3281 & ~n3282 ;
  assign n3284 = ~n2680 & ~n3283 ;
  assign n3285 = ~x161 & n2680 ;
  assign n3286 = ~n3284 & ~n3285 ;
  assign n3287 = n2728 & n3286 ;
  assign n3288 = ~n3280 & ~n3287 ;
  assign n3289 = ~n2826 & ~n3288 ;
  assign n3290 = n2728 & ~n3279 ;
  assign n3291 = ~n2728 & n3286 ;
  assign n3292 = ~n3290 & ~n3291 ;
  assign n3293 = ~n2782 & ~n3292 ;
  assign n3294 = x129 & n2782 ;
  assign n3295 = ~n3293 & ~n3294 ;
  assign n3296 = n2826 & ~n3295 ;
  assign n3297 = ~n3289 & ~n3296 ;
  assign n3298 = ~n2925 & ~n3297 ;
  assign n3299 = n2826 & ~n3288 ;
  assign n3300 = ~n2826 & ~n3295 ;
  assign n3301 = ~n3299 & ~n3300 ;
  assign n3302 = ~n2880 & ~n3301 ;
  assign n3303 = x97 & n2880 ;
  assign n3304 = ~n3302 & ~n3303 ;
  assign n3305 = n2925 & ~n3304 ;
  assign n3306 = ~n3298 & ~n3305 ;
  assign n3307 = ~n3023 & ~n3306 ;
  assign n3308 = n2925 & ~n3297 ;
  assign n3309 = ~n2925 & ~n3304 ;
  assign n3310 = ~n3308 & ~n3309 ;
  assign n3311 = ~n2979 & ~n3310 ;
  assign n3312 = x65 & n2979 ;
  assign n3313 = ~n3311 & ~n3312 ;
  assign n3314 = n3023 & ~n3313 ;
  assign n3315 = ~n3307 & ~n3314 ;
  assign n3316 = ~n3121 & ~n3315 ;
  assign n3317 = n3023 & ~n3306 ;
  assign n3318 = ~n3023 & ~n3313 ;
  assign n3319 = ~n3317 & ~n3318 ;
  assign n3320 = ~n3073 & ~n3319 ;
  assign n3321 = x33 & n3073 ;
  assign n3322 = ~n3320 & ~n3321 ;
  assign n3323 = n3121 & ~n3322 ;
  assign n3324 = ~n3316 & ~n3323 ;
  assign n3325 = n3219 & ~n3324 ;
  assign n3326 = n3121 & ~n3315 ;
  assign n3327 = ~n3121 & ~n3322 ;
  assign n3328 = ~n3326 & ~n3327 ;
  assign n3329 = ~n3174 & ~n3328 ;
  assign n3330 = x1 & n3174 ;
  assign n3331 = ~n3329 & ~n3330 ;
  assign n3332 = ~n3219 & ~n3331 ;
  assign n3333 = ~n3325 & ~n3332 ;
  assign n3334 = x194 & ~n2630 ;
  assign n3335 = x226 & n2630 ;
  assign n3336 = ~n3334 & ~n3335 ;
  assign n3337 = ~n2728 & ~n3336 ;
  assign n3338 = ~x226 & ~n2630 ;
  assign n3339 = ~x194 & n2630 ;
  assign n3340 = ~n3338 & ~n3339 ;
  assign n3341 = ~n2680 & ~n3340 ;
  assign n3342 = ~x162 & n2680 ;
  assign n3343 = ~n3341 & ~n3342 ;
  assign n3344 = n2728 & n3343 ;
  assign n3345 = ~n3337 & ~n3344 ;
  assign n3346 = ~n2826 & ~n3345 ;
  assign n3347 = n2728 & ~n3336 ;
  assign n3348 = ~n2728 & n3343 ;
  assign n3349 = ~n3347 & ~n3348 ;
  assign n3350 = ~n2782 & ~n3349 ;
  assign n3351 = x130 & n2782 ;
  assign n3352 = ~n3350 & ~n3351 ;
  assign n3353 = n2826 & ~n3352 ;
  assign n3354 = ~n3346 & ~n3353 ;
  assign n3355 = ~n2925 & ~n3354 ;
  assign n3356 = n2826 & ~n3345 ;
  assign n3357 = ~n2826 & ~n3352 ;
  assign n3358 = ~n3356 & ~n3357 ;
  assign n3359 = ~n2880 & ~n3358 ;
  assign n3360 = x98 & n2880 ;
  assign n3361 = ~n3359 & ~n3360 ;
  assign n3362 = n2925 & ~n3361 ;
  assign n3363 = ~n3355 & ~n3362 ;
  assign n3364 = ~n3023 & ~n3363 ;
  assign n3365 = n2925 & ~n3354 ;
  assign n3366 = ~n2925 & ~n3361 ;
  assign n3367 = ~n3365 & ~n3366 ;
  assign n3368 = ~n2979 & ~n3367 ;
  assign n3369 = x66 & n2979 ;
  assign n3370 = ~n3368 & ~n3369 ;
  assign n3371 = n3023 & ~n3370 ;
  assign n3372 = ~n3364 & ~n3371 ;
  assign n3373 = ~n3121 & ~n3372 ;
  assign n3374 = n3023 & ~n3363 ;
  assign n3375 = ~n3023 & ~n3370 ;
  assign n3376 = ~n3374 & ~n3375 ;
  assign n3377 = ~n3073 & ~n3376 ;
  assign n3378 = x34 & n3073 ;
  assign n3379 = ~n3377 & ~n3378 ;
  assign n3380 = n3121 & ~n3379 ;
  assign n3381 = ~n3373 & ~n3380 ;
  assign n3382 = n3219 & ~n3381 ;
  assign n3383 = n3121 & ~n3372 ;
  assign n3384 = ~n3121 & ~n3379 ;
  assign n3385 = ~n3383 & ~n3384 ;
  assign n3386 = ~n3174 & ~n3385 ;
  assign n3387 = x2 & n3174 ;
  assign n3388 = ~n3386 & ~n3387 ;
  assign n3389 = ~n3219 & ~n3388 ;
  assign n3390 = ~n3382 & ~n3389 ;
  assign n3391 = x195 & ~n2630 ;
  assign n3392 = x227 & n2630 ;
  assign n3393 = ~n3391 & ~n3392 ;
  assign n3394 = ~n2728 & ~n3393 ;
  assign n3395 = ~x227 & ~n2630 ;
  assign n3396 = ~x195 & n2630 ;
  assign n3397 = ~n3395 & ~n3396 ;
  assign n3398 = ~n2680 & ~n3397 ;
  assign n3399 = ~x163 & n2680 ;
  assign n3400 = ~n3398 & ~n3399 ;
  assign n3401 = n2728 & n3400 ;
  assign n3402 = ~n3394 & ~n3401 ;
  assign n3403 = ~n2826 & ~n3402 ;
  assign n3404 = n2728 & ~n3393 ;
  assign n3405 = ~n2728 & n3400 ;
  assign n3406 = ~n3404 & ~n3405 ;
  assign n3407 = ~n2782 & ~n3406 ;
  assign n3408 = x131 & n2782 ;
  assign n3409 = ~n3407 & ~n3408 ;
  assign n3410 = n2826 & ~n3409 ;
  assign n3411 = ~n3403 & ~n3410 ;
  assign n3412 = ~n2925 & ~n3411 ;
  assign n3413 = n2826 & ~n3402 ;
  assign n3414 = ~n2826 & ~n3409 ;
  assign n3415 = ~n3413 & ~n3414 ;
  assign n3416 = ~n2880 & ~n3415 ;
  assign n3417 = x99 & n2880 ;
  assign n3418 = ~n3416 & ~n3417 ;
  assign n3419 = n2925 & ~n3418 ;
  assign n3420 = ~n3412 & ~n3419 ;
  assign n3421 = ~n3023 & ~n3420 ;
  assign n3422 = n2925 & ~n3411 ;
  assign n3423 = ~n2925 & ~n3418 ;
  assign n3424 = ~n3422 & ~n3423 ;
  assign n3425 = ~n2979 & ~n3424 ;
  assign n3426 = x67 & n2979 ;
  assign n3427 = ~n3425 & ~n3426 ;
  assign n3428 = n3023 & ~n3427 ;
  assign n3429 = ~n3421 & ~n3428 ;
  assign n3430 = ~n3121 & ~n3429 ;
  assign n3431 = n3023 & ~n3420 ;
  assign n3432 = ~n3023 & ~n3427 ;
  assign n3433 = ~n3431 & ~n3432 ;
  assign n3434 = ~n3073 & ~n3433 ;
  assign n3435 = x35 & n3073 ;
  assign n3436 = ~n3434 & ~n3435 ;
  assign n3437 = n3121 & ~n3436 ;
  assign n3438 = ~n3430 & ~n3437 ;
  assign n3439 = n3219 & ~n3438 ;
  assign n3440 = n3121 & ~n3429 ;
  assign n3441 = ~n3121 & ~n3436 ;
  assign n3442 = ~n3440 & ~n3441 ;
  assign n3443 = ~n3174 & ~n3442 ;
  assign n3444 = x3 & n3174 ;
  assign n3445 = ~n3443 & ~n3444 ;
  assign n3446 = ~n3219 & ~n3445 ;
  assign n3447 = ~n3439 & ~n3446 ;
  assign n3448 = x196 & ~n2630 ;
  assign n3449 = x228 & n2630 ;
  assign n3450 = ~n3448 & ~n3449 ;
  assign n3451 = ~n2728 & ~n3450 ;
  assign n3452 = ~x228 & ~n2630 ;
  assign n3453 = ~x196 & n2630 ;
  assign n3454 = ~n3452 & ~n3453 ;
  assign n3455 = ~n2680 & ~n3454 ;
  assign n3456 = ~x164 & n2680 ;
  assign n3457 = ~n3455 & ~n3456 ;
  assign n3458 = n2728 & n3457 ;
  assign n3459 = ~n3451 & ~n3458 ;
  assign n3460 = ~n2826 & ~n3459 ;
  assign n3461 = n2728 & ~n3450 ;
  assign n3462 = ~n2728 & n3457 ;
  assign n3463 = ~n3461 & ~n3462 ;
  assign n3464 = ~n2782 & ~n3463 ;
  assign n3465 = x132 & n2782 ;
  assign n3466 = ~n3464 & ~n3465 ;
  assign n3467 = n2826 & ~n3466 ;
  assign n3468 = ~n3460 & ~n3467 ;
  assign n3469 = ~n2925 & ~n3468 ;
  assign n3470 = n2826 & ~n3459 ;
  assign n3471 = ~n2826 & ~n3466 ;
  assign n3472 = ~n3470 & ~n3471 ;
  assign n3473 = ~n2880 & ~n3472 ;
  assign n3474 = x100 & n2880 ;
  assign n3475 = ~n3473 & ~n3474 ;
  assign n3476 = n2925 & ~n3475 ;
  assign n3477 = ~n3469 & ~n3476 ;
  assign n3478 = ~n3023 & ~n3477 ;
  assign n3479 = n2925 & ~n3468 ;
  assign n3480 = ~n2925 & ~n3475 ;
  assign n3481 = ~n3479 & ~n3480 ;
  assign n3482 = ~n2979 & ~n3481 ;
  assign n3483 = x68 & n2979 ;
  assign n3484 = ~n3482 & ~n3483 ;
  assign n3485 = n3023 & ~n3484 ;
  assign n3486 = ~n3478 & ~n3485 ;
  assign n3487 = ~n3121 & ~n3486 ;
  assign n3488 = n3023 & ~n3477 ;
  assign n3489 = ~n3023 & ~n3484 ;
  assign n3490 = ~n3488 & ~n3489 ;
  assign n3491 = ~n3073 & ~n3490 ;
  assign n3492 = x36 & n3073 ;
  assign n3493 = ~n3491 & ~n3492 ;
  assign n3494 = n3121 & ~n3493 ;
  assign n3495 = ~n3487 & ~n3494 ;
  assign n3496 = n3219 & ~n3495 ;
  assign n3497 = n3121 & ~n3486 ;
  assign n3498 = ~n3121 & ~n3493 ;
  assign n3499 = ~n3497 & ~n3498 ;
  assign n3500 = ~n3174 & ~n3499 ;
  assign n3501 = x4 & n3174 ;
  assign n3502 = ~n3500 & ~n3501 ;
  assign n3503 = ~n3219 & ~n3502 ;
  assign n3504 = ~n3496 & ~n3503 ;
  assign n3505 = x197 & ~n2630 ;
  assign n3506 = x229 & n2630 ;
  assign n3507 = ~n3505 & ~n3506 ;
  assign n3508 = ~n2728 & ~n3507 ;
  assign n3509 = ~x229 & ~n2630 ;
  assign n3510 = ~x197 & n2630 ;
  assign n3511 = ~n3509 & ~n3510 ;
  assign n3512 = ~n2680 & ~n3511 ;
  assign n3513 = ~x165 & n2680 ;
  assign n3514 = ~n3512 & ~n3513 ;
  assign n3515 = n2728 & n3514 ;
  assign n3516 = ~n3508 & ~n3515 ;
  assign n3517 = ~n2826 & ~n3516 ;
  assign n3518 = n2728 & ~n3507 ;
  assign n3519 = ~n2728 & n3514 ;
  assign n3520 = ~n3518 & ~n3519 ;
  assign n3521 = ~n2782 & ~n3520 ;
  assign n3522 = x133 & n2782 ;
  assign n3523 = ~n3521 & ~n3522 ;
  assign n3524 = n2826 & ~n3523 ;
  assign n3525 = ~n3517 & ~n3524 ;
  assign n3526 = ~n2925 & ~n3525 ;
  assign n3527 = n2826 & ~n3516 ;
  assign n3528 = ~n2826 & ~n3523 ;
  assign n3529 = ~n3527 & ~n3528 ;
  assign n3530 = ~n2880 & ~n3529 ;
  assign n3531 = x101 & n2880 ;
  assign n3532 = ~n3530 & ~n3531 ;
  assign n3533 = n2925 & ~n3532 ;
  assign n3534 = ~n3526 & ~n3533 ;
  assign n3535 = ~n3023 & ~n3534 ;
  assign n3536 = n2925 & ~n3525 ;
  assign n3537 = ~n2925 & ~n3532 ;
  assign n3538 = ~n3536 & ~n3537 ;
  assign n3539 = ~n2979 & ~n3538 ;
  assign n3540 = x69 & n2979 ;
  assign n3541 = ~n3539 & ~n3540 ;
  assign n3542 = n3023 & ~n3541 ;
  assign n3543 = ~n3535 & ~n3542 ;
  assign n3544 = ~n3121 & ~n3543 ;
  assign n3545 = n3023 & ~n3534 ;
  assign n3546 = ~n3023 & ~n3541 ;
  assign n3547 = ~n3545 & ~n3546 ;
  assign n3548 = ~n3073 & ~n3547 ;
  assign n3549 = x37 & n3073 ;
  assign n3550 = ~n3548 & ~n3549 ;
  assign n3551 = n3121 & ~n3550 ;
  assign n3552 = ~n3544 & ~n3551 ;
  assign n3553 = n3219 & ~n3552 ;
  assign n3554 = n3121 & ~n3543 ;
  assign n3555 = ~n3121 & ~n3550 ;
  assign n3556 = ~n3554 & ~n3555 ;
  assign n3557 = ~n3174 & ~n3556 ;
  assign n3558 = x5 & n3174 ;
  assign n3559 = ~n3557 & ~n3558 ;
  assign n3560 = ~n3219 & ~n3559 ;
  assign n3561 = ~n3553 & ~n3560 ;
  assign n3562 = x198 & ~n2630 ;
  assign n3563 = x230 & n2630 ;
  assign n3564 = ~n3562 & ~n3563 ;
  assign n3565 = ~n2728 & ~n3564 ;
  assign n3566 = ~x230 & ~n2630 ;
  assign n3567 = ~x198 & n2630 ;
  assign n3568 = ~n3566 & ~n3567 ;
  assign n3569 = ~n2680 & ~n3568 ;
  assign n3570 = ~x166 & n2680 ;
  assign n3571 = ~n3569 & ~n3570 ;
  assign n3572 = n2728 & n3571 ;
  assign n3573 = ~n3565 & ~n3572 ;
  assign n3574 = ~n2826 & ~n3573 ;
  assign n3575 = n2728 & ~n3564 ;
  assign n3576 = ~n2728 & n3571 ;
  assign n3577 = ~n3575 & ~n3576 ;
  assign n3578 = ~n2782 & ~n3577 ;
  assign n3579 = x134 & n2782 ;
  assign n3580 = ~n3578 & ~n3579 ;
  assign n3581 = n2826 & ~n3580 ;
  assign n3582 = ~n3574 & ~n3581 ;
  assign n3583 = ~n2925 & ~n3582 ;
  assign n3584 = n2826 & ~n3573 ;
  assign n3585 = ~n2826 & ~n3580 ;
  assign n3586 = ~n3584 & ~n3585 ;
  assign n3587 = ~n2880 & ~n3586 ;
  assign n3588 = x102 & n2880 ;
  assign n3589 = ~n3587 & ~n3588 ;
  assign n3590 = n2925 & ~n3589 ;
  assign n3591 = ~n3583 & ~n3590 ;
  assign n3592 = ~n3023 & ~n3591 ;
  assign n3593 = n2925 & ~n3582 ;
  assign n3594 = ~n2925 & ~n3589 ;
  assign n3595 = ~n3593 & ~n3594 ;
  assign n3596 = ~n2979 & ~n3595 ;
  assign n3597 = x70 & n2979 ;
  assign n3598 = ~n3596 & ~n3597 ;
  assign n3599 = n3023 & ~n3598 ;
  assign n3600 = ~n3592 & ~n3599 ;
  assign n3601 = ~n3121 & ~n3600 ;
  assign n3602 = n3023 & ~n3591 ;
  assign n3603 = ~n3023 & ~n3598 ;
  assign n3604 = ~n3602 & ~n3603 ;
  assign n3605 = ~n3073 & ~n3604 ;
  assign n3606 = x38 & n3073 ;
  assign n3607 = ~n3605 & ~n3606 ;
  assign n3608 = n3121 & ~n3607 ;
  assign n3609 = ~n3601 & ~n3608 ;
  assign n3610 = n3219 & ~n3609 ;
  assign n3611 = n3121 & ~n3600 ;
  assign n3612 = ~n3121 & ~n3607 ;
  assign n3613 = ~n3611 & ~n3612 ;
  assign n3614 = ~n3174 & ~n3613 ;
  assign n3615 = x6 & n3174 ;
  assign n3616 = ~n3614 & ~n3615 ;
  assign n3617 = ~n3219 & ~n3616 ;
  assign n3618 = ~n3610 & ~n3617 ;
  assign n3619 = x199 & ~n2630 ;
  assign n3620 = x231 & n2630 ;
  assign n3621 = ~n3619 & ~n3620 ;
  assign n3622 = ~n2728 & ~n3621 ;
  assign n3623 = ~x231 & ~n2630 ;
  assign n3624 = ~x199 & n2630 ;
  assign n3625 = ~n3623 & ~n3624 ;
  assign n3626 = ~n2680 & ~n3625 ;
  assign n3627 = ~x167 & n2680 ;
  assign n3628 = ~n3626 & ~n3627 ;
  assign n3629 = n2728 & n3628 ;
  assign n3630 = ~n3622 & ~n3629 ;
  assign n3631 = ~n2826 & ~n3630 ;
  assign n3632 = n2728 & ~n3621 ;
  assign n3633 = ~n2728 & n3628 ;
  assign n3634 = ~n3632 & ~n3633 ;
  assign n3635 = ~n2782 & ~n3634 ;
  assign n3636 = x135 & n2782 ;
  assign n3637 = ~n3635 & ~n3636 ;
  assign n3638 = n2826 & ~n3637 ;
  assign n3639 = ~n3631 & ~n3638 ;
  assign n3640 = ~n2925 & ~n3639 ;
  assign n3641 = n2826 & ~n3630 ;
  assign n3642 = ~n2826 & ~n3637 ;
  assign n3643 = ~n3641 & ~n3642 ;
  assign n3644 = ~n2880 & ~n3643 ;
  assign n3645 = x103 & n2880 ;
  assign n3646 = ~n3644 & ~n3645 ;
  assign n3647 = n2925 & ~n3646 ;
  assign n3648 = ~n3640 & ~n3647 ;
  assign n3649 = ~n3023 & ~n3648 ;
  assign n3650 = n2925 & ~n3639 ;
  assign n3651 = ~n2925 & ~n3646 ;
  assign n3652 = ~n3650 & ~n3651 ;
  assign n3653 = ~n2979 & ~n3652 ;
  assign n3654 = x71 & n2979 ;
  assign n3655 = ~n3653 & ~n3654 ;
  assign n3656 = n3023 & ~n3655 ;
  assign n3657 = ~n3649 & ~n3656 ;
  assign n3658 = ~n3121 & ~n3657 ;
  assign n3659 = n3023 & ~n3648 ;
  assign n3660 = ~n3023 & ~n3655 ;
  assign n3661 = ~n3659 & ~n3660 ;
  assign n3662 = ~n3073 & ~n3661 ;
  assign n3663 = x39 & n3073 ;
  assign n3664 = ~n3662 & ~n3663 ;
  assign n3665 = n3121 & ~n3664 ;
  assign n3666 = ~n3658 & ~n3665 ;
  assign n3667 = n3219 & ~n3666 ;
  assign n3668 = n3121 & ~n3657 ;
  assign n3669 = ~n3121 & ~n3664 ;
  assign n3670 = ~n3668 & ~n3669 ;
  assign n3671 = ~n3174 & ~n3670 ;
  assign n3672 = x7 & n3174 ;
  assign n3673 = ~n3671 & ~n3672 ;
  assign n3674 = ~n3219 & ~n3673 ;
  assign n3675 = ~n3667 & ~n3674 ;
  assign n3676 = x200 & ~n2630 ;
  assign n3677 = x232 & n2630 ;
  assign n3678 = ~n3676 & ~n3677 ;
  assign n3679 = ~n2728 & ~n3678 ;
  assign n3680 = ~x232 & ~n2630 ;
  assign n3681 = ~x200 & n2630 ;
  assign n3682 = ~n3680 & ~n3681 ;
  assign n3683 = ~n2680 & ~n3682 ;
  assign n3684 = ~x168 & n2680 ;
  assign n3685 = ~n3683 & ~n3684 ;
  assign n3686 = n2728 & n3685 ;
  assign n3687 = ~n3679 & ~n3686 ;
  assign n3688 = ~n2826 & ~n3687 ;
  assign n3689 = n2728 & ~n3678 ;
  assign n3690 = ~n2728 & n3685 ;
  assign n3691 = ~n3689 & ~n3690 ;
  assign n3692 = ~n2782 & ~n3691 ;
  assign n3693 = x136 & n2782 ;
  assign n3694 = ~n3692 & ~n3693 ;
  assign n3695 = n2826 & ~n3694 ;
  assign n3696 = ~n3688 & ~n3695 ;
  assign n3697 = ~n2925 & ~n3696 ;
  assign n3698 = n2826 & ~n3687 ;
  assign n3699 = ~n2826 & ~n3694 ;
  assign n3700 = ~n3698 & ~n3699 ;
  assign n3701 = ~n2880 & ~n3700 ;
  assign n3702 = x104 & n2880 ;
  assign n3703 = ~n3701 & ~n3702 ;
  assign n3704 = n2925 & ~n3703 ;
  assign n3705 = ~n3697 & ~n3704 ;
  assign n3706 = ~n3023 & ~n3705 ;
  assign n3707 = n2925 & ~n3696 ;
  assign n3708 = ~n2925 & ~n3703 ;
  assign n3709 = ~n3707 & ~n3708 ;
  assign n3710 = ~n2979 & ~n3709 ;
  assign n3711 = x72 & n2979 ;
  assign n3712 = ~n3710 & ~n3711 ;
  assign n3713 = n3023 & ~n3712 ;
  assign n3714 = ~n3706 & ~n3713 ;
  assign n3715 = ~n3121 & ~n3714 ;
  assign n3716 = n3023 & ~n3705 ;
  assign n3717 = ~n3023 & ~n3712 ;
  assign n3718 = ~n3716 & ~n3717 ;
  assign n3719 = ~n3073 & ~n3718 ;
  assign n3720 = x40 & n3073 ;
  assign n3721 = ~n3719 & ~n3720 ;
  assign n3722 = n3121 & ~n3721 ;
  assign n3723 = ~n3715 & ~n3722 ;
  assign n3724 = n3219 & ~n3723 ;
  assign n3725 = n3121 & ~n3714 ;
  assign n3726 = ~n3121 & ~n3721 ;
  assign n3727 = ~n3725 & ~n3726 ;
  assign n3728 = ~n3174 & ~n3727 ;
  assign n3729 = x8 & n3174 ;
  assign n3730 = ~n3728 & ~n3729 ;
  assign n3731 = ~n3219 & ~n3730 ;
  assign n3732 = ~n3724 & ~n3731 ;
  assign n3733 = x201 & ~n2630 ;
  assign n3734 = x233 & n2630 ;
  assign n3735 = ~n3733 & ~n3734 ;
  assign n3736 = ~n2728 & ~n3735 ;
  assign n3737 = ~x233 & ~n2630 ;
  assign n3738 = ~x201 & n2630 ;
  assign n3739 = ~n3737 & ~n3738 ;
  assign n3740 = ~n2680 & ~n3739 ;
  assign n3741 = ~x169 & n2680 ;
  assign n3742 = ~n3740 & ~n3741 ;
  assign n3743 = n2728 & n3742 ;
  assign n3744 = ~n3736 & ~n3743 ;
  assign n3745 = ~n2826 & ~n3744 ;
  assign n3746 = n2728 & ~n3735 ;
  assign n3747 = ~n2728 & n3742 ;
  assign n3748 = ~n3746 & ~n3747 ;
  assign n3749 = ~n2782 & ~n3748 ;
  assign n3750 = x137 & n2782 ;
  assign n3751 = ~n3749 & ~n3750 ;
  assign n3752 = n2826 & ~n3751 ;
  assign n3753 = ~n3745 & ~n3752 ;
  assign n3754 = ~n2925 & ~n3753 ;
  assign n3755 = n2826 & ~n3744 ;
  assign n3756 = ~n2826 & ~n3751 ;
  assign n3757 = ~n3755 & ~n3756 ;
  assign n3758 = ~n2880 & ~n3757 ;
  assign n3759 = x105 & n2880 ;
  assign n3760 = ~n3758 & ~n3759 ;
  assign n3761 = n2925 & ~n3760 ;
  assign n3762 = ~n3754 & ~n3761 ;
  assign n3763 = ~n3023 & ~n3762 ;
  assign n3764 = n2925 & ~n3753 ;
  assign n3765 = ~n2925 & ~n3760 ;
  assign n3766 = ~n3764 & ~n3765 ;
  assign n3767 = ~n2979 & ~n3766 ;
  assign n3768 = x73 & n2979 ;
  assign n3769 = ~n3767 & ~n3768 ;
  assign n3770 = n3023 & ~n3769 ;
  assign n3771 = ~n3763 & ~n3770 ;
  assign n3772 = ~n3121 & ~n3771 ;
  assign n3773 = n3023 & ~n3762 ;
  assign n3774 = ~n3023 & ~n3769 ;
  assign n3775 = ~n3773 & ~n3774 ;
  assign n3776 = ~n3073 & ~n3775 ;
  assign n3777 = x41 & n3073 ;
  assign n3778 = ~n3776 & ~n3777 ;
  assign n3779 = n3121 & ~n3778 ;
  assign n3780 = ~n3772 & ~n3779 ;
  assign n3781 = n3219 & ~n3780 ;
  assign n3782 = n3121 & ~n3771 ;
  assign n3783 = ~n3121 & ~n3778 ;
  assign n3784 = ~n3782 & ~n3783 ;
  assign n3785 = ~n3174 & ~n3784 ;
  assign n3786 = x9 & n3174 ;
  assign n3787 = ~n3785 & ~n3786 ;
  assign n3788 = ~n3219 & ~n3787 ;
  assign n3789 = ~n3781 & ~n3788 ;
  assign n3790 = x202 & ~n2630 ;
  assign n3791 = x234 & n2630 ;
  assign n3792 = ~n3790 & ~n3791 ;
  assign n3793 = ~n2728 & ~n3792 ;
  assign n3794 = ~x234 & ~n2630 ;
  assign n3795 = ~x202 & n2630 ;
  assign n3796 = ~n3794 & ~n3795 ;
  assign n3797 = ~n2680 & ~n3796 ;
  assign n3798 = ~x170 & n2680 ;
  assign n3799 = ~n3797 & ~n3798 ;
  assign n3800 = n2728 & n3799 ;
  assign n3801 = ~n3793 & ~n3800 ;
  assign n3802 = ~n2826 & ~n3801 ;
  assign n3803 = n2728 & ~n3792 ;
  assign n3804 = ~n2728 & n3799 ;
  assign n3805 = ~n3803 & ~n3804 ;
  assign n3806 = ~n2782 & ~n3805 ;
  assign n3807 = x138 & n2782 ;
  assign n3808 = ~n3806 & ~n3807 ;
  assign n3809 = n2826 & ~n3808 ;
  assign n3810 = ~n3802 & ~n3809 ;
  assign n3811 = ~n2925 & ~n3810 ;
  assign n3812 = n2826 & ~n3801 ;
  assign n3813 = ~n2826 & ~n3808 ;
  assign n3814 = ~n3812 & ~n3813 ;
  assign n3815 = ~n2880 & ~n3814 ;
  assign n3816 = x106 & n2880 ;
  assign n3817 = ~n3815 & ~n3816 ;
  assign n3818 = n2925 & ~n3817 ;
  assign n3819 = ~n3811 & ~n3818 ;
  assign n3820 = ~n3023 & ~n3819 ;
  assign n3821 = n2925 & ~n3810 ;
  assign n3822 = ~n2925 & ~n3817 ;
  assign n3823 = ~n3821 & ~n3822 ;
  assign n3824 = ~n2979 & ~n3823 ;
  assign n3825 = x74 & n2979 ;
  assign n3826 = ~n3824 & ~n3825 ;
  assign n3827 = n3023 & ~n3826 ;
  assign n3828 = ~n3820 & ~n3827 ;
  assign n3829 = ~n3121 & ~n3828 ;
  assign n3830 = n3023 & ~n3819 ;
  assign n3831 = ~n3023 & ~n3826 ;
  assign n3832 = ~n3830 & ~n3831 ;
  assign n3833 = ~n3073 & ~n3832 ;
  assign n3834 = x42 & n3073 ;
  assign n3835 = ~n3833 & ~n3834 ;
  assign n3836 = n3121 & ~n3835 ;
  assign n3837 = ~n3829 & ~n3836 ;
  assign n3838 = n3219 & ~n3837 ;
  assign n3839 = n3121 & ~n3828 ;
  assign n3840 = ~n3121 & ~n3835 ;
  assign n3841 = ~n3839 & ~n3840 ;
  assign n3842 = ~n3174 & ~n3841 ;
  assign n3843 = x10 & n3174 ;
  assign n3844 = ~n3842 & ~n3843 ;
  assign n3845 = ~n3219 & ~n3844 ;
  assign n3846 = ~n3838 & ~n3845 ;
  assign n3847 = x203 & ~n2630 ;
  assign n3848 = x235 & n2630 ;
  assign n3849 = ~n3847 & ~n3848 ;
  assign n3850 = ~n2728 & ~n3849 ;
  assign n3851 = ~x235 & ~n2630 ;
  assign n3852 = ~x203 & n2630 ;
  assign n3853 = ~n3851 & ~n3852 ;
  assign n3854 = ~n2680 & ~n3853 ;
  assign n3855 = ~x171 & n2680 ;
  assign n3856 = ~n3854 & ~n3855 ;
  assign n3857 = n2728 & n3856 ;
  assign n3858 = ~n3850 & ~n3857 ;
  assign n3859 = ~n2826 & ~n3858 ;
  assign n3860 = n2728 & ~n3849 ;
  assign n3861 = ~n2728 & n3856 ;
  assign n3862 = ~n3860 & ~n3861 ;
  assign n3863 = ~n2782 & ~n3862 ;
  assign n3864 = x139 & n2782 ;
  assign n3865 = ~n3863 & ~n3864 ;
  assign n3866 = n2826 & ~n3865 ;
  assign n3867 = ~n3859 & ~n3866 ;
  assign n3868 = ~n2925 & ~n3867 ;
  assign n3869 = n2826 & ~n3858 ;
  assign n3870 = ~n2826 & ~n3865 ;
  assign n3871 = ~n3869 & ~n3870 ;
  assign n3872 = ~n2880 & ~n3871 ;
  assign n3873 = x107 & n2880 ;
  assign n3874 = ~n3872 & ~n3873 ;
  assign n3875 = n2925 & ~n3874 ;
  assign n3876 = ~n3868 & ~n3875 ;
  assign n3877 = ~n3023 & ~n3876 ;
  assign n3878 = n2925 & ~n3867 ;
  assign n3879 = ~n2925 & ~n3874 ;
  assign n3880 = ~n3878 & ~n3879 ;
  assign n3881 = ~n2979 & ~n3880 ;
  assign n3882 = x75 & n2979 ;
  assign n3883 = ~n3881 & ~n3882 ;
  assign n3884 = n3023 & ~n3883 ;
  assign n3885 = ~n3877 & ~n3884 ;
  assign n3886 = ~n3121 & ~n3885 ;
  assign n3887 = n3023 & ~n3876 ;
  assign n3888 = ~n3023 & ~n3883 ;
  assign n3889 = ~n3887 & ~n3888 ;
  assign n3890 = ~n3073 & ~n3889 ;
  assign n3891 = x43 & n3073 ;
  assign n3892 = ~n3890 & ~n3891 ;
  assign n3893 = n3121 & ~n3892 ;
  assign n3894 = ~n3886 & ~n3893 ;
  assign n3895 = n3219 & ~n3894 ;
  assign n3896 = n3121 & ~n3885 ;
  assign n3897 = ~n3121 & ~n3892 ;
  assign n3898 = ~n3896 & ~n3897 ;
  assign n3899 = ~n3174 & ~n3898 ;
  assign n3900 = x11 & n3174 ;
  assign n3901 = ~n3899 & ~n3900 ;
  assign n3902 = ~n3219 & ~n3901 ;
  assign n3903 = ~n3895 & ~n3902 ;
  assign n3904 = x204 & ~n2630 ;
  assign n3905 = x236 & n2630 ;
  assign n3906 = ~n3904 & ~n3905 ;
  assign n3907 = ~n2728 & ~n3906 ;
  assign n3908 = ~x236 & ~n2630 ;
  assign n3909 = ~x204 & n2630 ;
  assign n3910 = ~n3908 & ~n3909 ;
  assign n3911 = ~n2680 & ~n3910 ;
  assign n3912 = ~x172 & n2680 ;
  assign n3913 = ~n3911 & ~n3912 ;
  assign n3914 = n2728 & n3913 ;
  assign n3915 = ~n3907 & ~n3914 ;
  assign n3916 = ~n2826 & ~n3915 ;
  assign n3917 = n2728 & ~n3906 ;
  assign n3918 = ~n2728 & n3913 ;
  assign n3919 = ~n3917 & ~n3918 ;
  assign n3920 = ~n2782 & ~n3919 ;
  assign n3921 = x140 & n2782 ;
  assign n3922 = ~n3920 & ~n3921 ;
  assign n3923 = n2826 & ~n3922 ;
  assign n3924 = ~n3916 & ~n3923 ;
  assign n3925 = ~n2925 & ~n3924 ;
  assign n3926 = n2826 & ~n3915 ;
  assign n3927 = ~n2826 & ~n3922 ;
  assign n3928 = ~n3926 & ~n3927 ;
  assign n3929 = ~n2880 & ~n3928 ;
  assign n3930 = x108 & n2880 ;
  assign n3931 = ~n3929 & ~n3930 ;
  assign n3932 = n2925 & ~n3931 ;
  assign n3933 = ~n3925 & ~n3932 ;
  assign n3934 = ~n3023 & ~n3933 ;
  assign n3935 = n2925 & ~n3924 ;
  assign n3936 = ~n2925 & ~n3931 ;
  assign n3937 = ~n3935 & ~n3936 ;
  assign n3938 = ~n2979 & ~n3937 ;
  assign n3939 = x76 & n2979 ;
  assign n3940 = ~n3938 & ~n3939 ;
  assign n3941 = n3023 & ~n3940 ;
  assign n3942 = ~n3934 & ~n3941 ;
  assign n3943 = ~n3121 & ~n3942 ;
  assign n3944 = n3023 & ~n3933 ;
  assign n3945 = ~n3023 & ~n3940 ;
  assign n3946 = ~n3944 & ~n3945 ;
  assign n3947 = ~n3073 & ~n3946 ;
  assign n3948 = x44 & n3073 ;
  assign n3949 = ~n3947 & ~n3948 ;
  assign n3950 = n3121 & ~n3949 ;
  assign n3951 = ~n3943 & ~n3950 ;
  assign n3952 = n3219 & ~n3951 ;
  assign n3953 = n3121 & ~n3942 ;
  assign n3954 = ~n3121 & ~n3949 ;
  assign n3955 = ~n3953 & ~n3954 ;
  assign n3956 = ~n3174 & ~n3955 ;
  assign n3957 = x12 & n3174 ;
  assign n3958 = ~n3956 & ~n3957 ;
  assign n3959 = ~n3219 & ~n3958 ;
  assign n3960 = ~n3952 & ~n3959 ;
  assign n3961 = x205 & ~n2630 ;
  assign n3962 = x237 & n2630 ;
  assign n3963 = ~n3961 & ~n3962 ;
  assign n3964 = ~n2728 & ~n3963 ;
  assign n3965 = ~x237 & ~n2630 ;
  assign n3966 = ~x205 & n2630 ;
  assign n3967 = ~n3965 & ~n3966 ;
  assign n3968 = ~n2680 & ~n3967 ;
  assign n3969 = ~x173 & n2680 ;
  assign n3970 = ~n3968 & ~n3969 ;
  assign n3971 = n2728 & n3970 ;
  assign n3972 = ~n3964 & ~n3971 ;
  assign n3973 = ~n2826 & ~n3972 ;
  assign n3974 = n2728 & ~n3963 ;
  assign n3975 = ~n2728 & n3970 ;
  assign n3976 = ~n3974 & ~n3975 ;
  assign n3977 = ~n2782 & ~n3976 ;
  assign n3978 = x141 & n2782 ;
  assign n3979 = ~n3977 & ~n3978 ;
  assign n3980 = n2826 & ~n3979 ;
  assign n3981 = ~n3973 & ~n3980 ;
  assign n3982 = ~n2925 & ~n3981 ;
  assign n3983 = n2826 & ~n3972 ;
  assign n3984 = ~n2826 & ~n3979 ;
  assign n3985 = ~n3983 & ~n3984 ;
  assign n3986 = ~n2880 & ~n3985 ;
  assign n3987 = x109 & n2880 ;
  assign n3988 = ~n3986 & ~n3987 ;
  assign n3989 = n2925 & ~n3988 ;
  assign n3990 = ~n3982 & ~n3989 ;
  assign n3991 = ~n3023 & ~n3990 ;
  assign n3992 = n2925 & ~n3981 ;
  assign n3993 = ~n2925 & ~n3988 ;
  assign n3994 = ~n3992 & ~n3993 ;
  assign n3995 = ~n2979 & ~n3994 ;
  assign n3996 = x77 & n2979 ;
  assign n3997 = ~n3995 & ~n3996 ;
  assign n3998 = n3023 & ~n3997 ;
  assign n3999 = ~n3991 & ~n3998 ;
  assign n4000 = ~n3121 & ~n3999 ;
  assign n4001 = n3023 & ~n3990 ;
  assign n4002 = ~n3023 & ~n3997 ;
  assign n4003 = ~n4001 & ~n4002 ;
  assign n4004 = ~n3073 & ~n4003 ;
  assign n4005 = x45 & n3073 ;
  assign n4006 = ~n4004 & ~n4005 ;
  assign n4007 = n3121 & ~n4006 ;
  assign n4008 = ~n4000 & ~n4007 ;
  assign n4009 = n3219 & ~n4008 ;
  assign n4010 = n3121 & ~n3999 ;
  assign n4011 = ~n3121 & ~n4006 ;
  assign n4012 = ~n4010 & ~n4011 ;
  assign n4013 = ~n3174 & ~n4012 ;
  assign n4014 = x13 & n3174 ;
  assign n4015 = ~n4013 & ~n4014 ;
  assign n4016 = ~n3219 & ~n4015 ;
  assign n4017 = ~n4009 & ~n4016 ;
  assign n4018 = x206 & ~n2630 ;
  assign n4019 = x238 & n2630 ;
  assign n4020 = ~n4018 & ~n4019 ;
  assign n4021 = ~n2728 & ~n4020 ;
  assign n4022 = ~x238 & ~n2630 ;
  assign n4023 = ~x206 & n2630 ;
  assign n4024 = ~n4022 & ~n4023 ;
  assign n4025 = ~n2680 & ~n4024 ;
  assign n4026 = ~x174 & n2680 ;
  assign n4027 = ~n4025 & ~n4026 ;
  assign n4028 = n2728 & n4027 ;
  assign n4029 = ~n4021 & ~n4028 ;
  assign n4030 = ~n2826 & ~n4029 ;
  assign n4031 = n2728 & ~n4020 ;
  assign n4032 = ~n2728 & n4027 ;
  assign n4033 = ~n4031 & ~n4032 ;
  assign n4034 = ~n2782 & ~n4033 ;
  assign n4035 = x142 & n2782 ;
  assign n4036 = ~n4034 & ~n4035 ;
  assign n4037 = n2826 & ~n4036 ;
  assign n4038 = ~n4030 & ~n4037 ;
  assign n4039 = ~n2925 & ~n4038 ;
  assign n4040 = n2826 & ~n4029 ;
  assign n4041 = ~n2826 & ~n4036 ;
  assign n4042 = ~n4040 & ~n4041 ;
  assign n4043 = ~n2880 & ~n4042 ;
  assign n4044 = x110 & n2880 ;
  assign n4045 = ~n4043 & ~n4044 ;
  assign n4046 = n2925 & ~n4045 ;
  assign n4047 = ~n4039 & ~n4046 ;
  assign n4048 = ~n3023 & ~n4047 ;
  assign n4049 = n2925 & ~n4038 ;
  assign n4050 = ~n2925 & ~n4045 ;
  assign n4051 = ~n4049 & ~n4050 ;
  assign n4052 = ~n2979 & ~n4051 ;
  assign n4053 = x78 & n2979 ;
  assign n4054 = ~n4052 & ~n4053 ;
  assign n4055 = n3023 & ~n4054 ;
  assign n4056 = ~n4048 & ~n4055 ;
  assign n4057 = ~n3121 & ~n4056 ;
  assign n4058 = n3023 & ~n4047 ;
  assign n4059 = ~n3023 & ~n4054 ;
  assign n4060 = ~n4058 & ~n4059 ;
  assign n4061 = ~n3073 & ~n4060 ;
  assign n4062 = x46 & n3073 ;
  assign n4063 = ~n4061 & ~n4062 ;
  assign n4064 = n3121 & ~n4063 ;
  assign n4065 = ~n4057 & ~n4064 ;
  assign n4066 = n3219 & ~n4065 ;
  assign n4067 = n3121 & ~n4056 ;
  assign n4068 = ~n3121 & ~n4063 ;
  assign n4069 = ~n4067 & ~n4068 ;
  assign n4070 = ~n3174 & ~n4069 ;
  assign n4071 = x14 & n3174 ;
  assign n4072 = ~n4070 & ~n4071 ;
  assign n4073 = ~n3219 & ~n4072 ;
  assign n4074 = ~n4066 & ~n4073 ;
  assign n4075 = x207 & ~n2630 ;
  assign n4076 = x239 & n2630 ;
  assign n4077 = ~n4075 & ~n4076 ;
  assign n4078 = ~n2728 & ~n4077 ;
  assign n4079 = ~x239 & ~n2630 ;
  assign n4080 = ~x207 & n2630 ;
  assign n4081 = ~n4079 & ~n4080 ;
  assign n4082 = ~n2680 & ~n4081 ;
  assign n4083 = ~x175 & n2680 ;
  assign n4084 = ~n4082 & ~n4083 ;
  assign n4085 = n2728 & n4084 ;
  assign n4086 = ~n4078 & ~n4085 ;
  assign n4087 = ~n2826 & ~n4086 ;
  assign n4088 = n2728 & ~n4077 ;
  assign n4089 = ~n2728 & n4084 ;
  assign n4090 = ~n4088 & ~n4089 ;
  assign n4091 = ~n2782 & ~n4090 ;
  assign n4092 = x143 & n2782 ;
  assign n4093 = ~n4091 & ~n4092 ;
  assign n4094 = n2826 & ~n4093 ;
  assign n4095 = ~n4087 & ~n4094 ;
  assign n4096 = ~n2925 & ~n4095 ;
  assign n4097 = n2826 & ~n4086 ;
  assign n4098 = ~n2826 & ~n4093 ;
  assign n4099 = ~n4097 & ~n4098 ;
  assign n4100 = ~n2880 & ~n4099 ;
  assign n4101 = x111 & n2880 ;
  assign n4102 = ~n4100 & ~n4101 ;
  assign n4103 = n2925 & ~n4102 ;
  assign n4104 = ~n4096 & ~n4103 ;
  assign n4105 = ~n3023 & ~n4104 ;
  assign n4106 = n2925 & ~n4095 ;
  assign n4107 = ~n2925 & ~n4102 ;
  assign n4108 = ~n4106 & ~n4107 ;
  assign n4109 = ~n2979 & ~n4108 ;
  assign n4110 = x79 & n2979 ;
  assign n4111 = ~n4109 & ~n4110 ;
  assign n4112 = n3023 & ~n4111 ;
  assign n4113 = ~n4105 & ~n4112 ;
  assign n4114 = ~n3121 & ~n4113 ;
  assign n4115 = n3023 & ~n4104 ;
  assign n4116 = ~n3023 & ~n4111 ;
  assign n4117 = ~n4115 & ~n4116 ;
  assign n4118 = ~n3073 & ~n4117 ;
  assign n4119 = x47 & n3073 ;
  assign n4120 = ~n4118 & ~n4119 ;
  assign n4121 = n3121 & ~n4120 ;
  assign n4122 = ~n4114 & ~n4121 ;
  assign n4123 = n3219 & ~n4122 ;
  assign n4124 = n3121 & ~n4113 ;
  assign n4125 = ~n3121 & ~n4120 ;
  assign n4126 = ~n4124 & ~n4125 ;
  assign n4127 = ~n3174 & ~n4126 ;
  assign n4128 = x15 & n3174 ;
  assign n4129 = ~n4127 & ~n4128 ;
  assign n4130 = ~n3219 & ~n4129 ;
  assign n4131 = ~n4123 & ~n4130 ;
  assign n4132 = x208 & ~n2630 ;
  assign n4133 = x240 & n2630 ;
  assign n4134 = ~n4132 & ~n4133 ;
  assign n4135 = ~n2728 & ~n4134 ;
  assign n4136 = ~x240 & ~n2630 ;
  assign n4137 = ~x208 & n2630 ;
  assign n4138 = ~n4136 & ~n4137 ;
  assign n4139 = ~n2680 & ~n4138 ;
  assign n4140 = ~x176 & n2680 ;
  assign n4141 = ~n4139 & ~n4140 ;
  assign n4142 = n2728 & n4141 ;
  assign n4143 = ~n4135 & ~n4142 ;
  assign n4144 = ~n2826 & ~n4143 ;
  assign n4145 = n2728 & ~n4134 ;
  assign n4146 = ~n2728 & n4141 ;
  assign n4147 = ~n4145 & ~n4146 ;
  assign n4148 = ~n2782 & ~n4147 ;
  assign n4149 = x144 & n2782 ;
  assign n4150 = ~n4148 & ~n4149 ;
  assign n4151 = n2826 & ~n4150 ;
  assign n4152 = ~n4144 & ~n4151 ;
  assign n4153 = ~n2925 & ~n4152 ;
  assign n4154 = n2826 & ~n4143 ;
  assign n4155 = ~n2826 & ~n4150 ;
  assign n4156 = ~n4154 & ~n4155 ;
  assign n4157 = ~n2880 & ~n4156 ;
  assign n4158 = x112 & n2880 ;
  assign n4159 = ~n4157 & ~n4158 ;
  assign n4160 = n2925 & ~n4159 ;
  assign n4161 = ~n4153 & ~n4160 ;
  assign n4162 = ~n3023 & ~n4161 ;
  assign n4163 = n2925 & ~n4152 ;
  assign n4164 = ~n2925 & ~n4159 ;
  assign n4165 = ~n4163 & ~n4164 ;
  assign n4166 = ~n2979 & ~n4165 ;
  assign n4167 = x80 & n2979 ;
  assign n4168 = ~n4166 & ~n4167 ;
  assign n4169 = n3023 & ~n4168 ;
  assign n4170 = ~n4162 & ~n4169 ;
  assign n4171 = ~n3121 & ~n4170 ;
  assign n4172 = n3023 & ~n4161 ;
  assign n4173 = ~n3023 & ~n4168 ;
  assign n4174 = ~n4172 & ~n4173 ;
  assign n4175 = ~n3073 & ~n4174 ;
  assign n4176 = x48 & n3073 ;
  assign n4177 = ~n4175 & ~n4176 ;
  assign n4178 = n3121 & ~n4177 ;
  assign n4179 = ~n4171 & ~n4178 ;
  assign n4180 = n3219 & ~n4179 ;
  assign n4181 = n3121 & ~n4170 ;
  assign n4182 = ~n3121 & ~n4177 ;
  assign n4183 = ~n4181 & ~n4182 ;
  assign n4184 = ~n3174 & ~n4183 ;
  assign n4185 = x16 & n3174 ;
  assign n4186 = ~n4184 & ~n4185 ;
  assign n4187 = ~n3219 & ~n4186 ;
  assign n4188 = ~n4180 & ~n4187 ;
  assign n4189 = x209 & ~n2630 ;
  assign n4190 = x241 & n2630 ;
  assign n4191 = ~n4189 & ~n4190 ;
  assign n4192 = ~n2728 & ~n4191 ;
  assign n4193 = ~x241 & ~n2630 ;
  assign n4194 = ~x209 & n2630 ;
  assign n4195 = ~n4193 & ~n4194 ;
  assign n4196 = ~n2680 & ~n4195 ;
  assign n4197 = ~x177 & n2680 ;
  assign n4198 = ~n4196 & ~n4197 ;
  assign n4199 = n2728 & n4198 ;
  assign n4200 = ~n4192 & ~n4199 ;
  assign n4201 = ~n2826 & ~n4200 ;
  assign n4202 = n2728 & ~n4191 ;
  assign n4203 = ~n2728 & n4198 ;
  assign n4204 = ~n4202 & ~n4203 ;
  assign n4205 = ~n2782 & ~n4204 ;
  assign n4206 = x145 & n2782 ;
  assign n4207 = ~n4205 & ~n4206 ;
  assign n4208 = n2826 & ~n4207 ;
  assign n4209 = ~n4201 & ~n4208 ;
  assign n4210 = ~n2925 & ~n4209 ;
  assign n4211 = n2826 & ~n4200 ;
  assign n4212 = ~n2826 & ~n4207 ;
  assign n4213 = ~n4211 & ~n4212 ;
  assign n4214 = ~n2880 & ~n4213 ;
  assign n4215 = x113 & n2880 ;
  assign n4216 = ~n4214 & ~n4215 ;
  assign n4217 = n2925 & ~n4216 ;
  assign n4218 = ~n4210 & ~n4217 ;
  assign n4219 = ~n3023 & ~n4218 ;
  assign n4220 = n2925 & ~n4209 ;
  assign n4221 = ~n2925 & ~n4216 ;
  assign n4222 = ~n4220 & ~n4221 ;
  assign n4223 = ~n2979 & ~n4222 ;
  assign n4224 = x81 & n2979 ;
  assign n4225 = ~n4223 & ~n4224 ;
  assign n4226 = n3023 & ~n4225 ;
  assign n4227 = ~n4219 & ~n4226 ;
  assign n4228 = ~n3121 & ~n4227 ;
  assign n4229 = n3023 & ~n4218 ;
  assign n4230 = ~n3023 & ~n4225 ;
  assign n4231 = ~n4229 & ~n4230 ;
  assign n4232 = ~n3073 & ~n4231 ;
  assign n4233 = x49 & n3073 ;
  assign n4234 = ~n4232 & ~n4233 ;
  assign n4235 = n3121 & ~n4234 ;
  assign n4236 = ~n4228 & ~n4235 ;
  assign n4237 = n3219 & ~n4236 ;
  assign n4238 = n3121 & ~n4227 ;
  assign n4239 = ~n3121 & ~n4234 ;
  assign n4240 = ~n4238 & ~n4239 ;
  assign n4241 = ~n3174 & ~n4240 ;
  assign n4242 = x17 & n3174 ;
  assign n4243 = ~n4241 & ~n4242 ;
  assign n4244 = ~n3219 & ~n4243 ;
  assign n4245 = ~n4237 & ~n4244 ;
  assign n4246 = x210 & ~n2630 ;
  assign n4247 = x242 & n2630 ;
  assign n4248 = ~n4246 & ~n4247 ;
  assign n4249 = ~n2728 & ~n4248 ;
  assign n4250 = ~x242 & ~n2630 ;
  assign n4251 = ~x210 & n2630 ;
  assign n4252 = ~n4250 & ~n4251 ;
  assign n4253 = ~n2680 & ~n4252 ;
  assign n4254 = ~x178 & n2680 ;
  assign n4255 = ~n4253 & ~n4254 ;
  assign n4256 = n2728 & n4255 ;
  assign n4257 = ~n4249 & ~n4256 ;
  assign n4258 = ~n2826 & ~n4257 ;
  assign n4259 = n2728 & ~n4248 ;
  assign n4260 = ~n2728 & n4255 ;
  assign n4261 = ~n4259 & ~n4260 ;
  assign n4262 = ~n2782 & ~n4261 ;
  assign n4263 = x146 & n2782 ;
  assign n4264 = ~n4262 & ~n4263 ;
  assign n4265 = n2826 & ~n4264 ;
  assign n4266 = ~n4258 & ~n4265 ;
  assign n4267 = ~n2925 & ~n4266 ;
  assign n4268 = n2826 & ~n4257 ;
  assign n4269 = ~n2826 & ~n4264 ;
  assign n4270 = ~n4268 & ~n4269 ;
  assign n4271 = ~n2880 & ~n4270 ;
  assign n4272 = x114 & n2880 ;
  assign n4273 = ~n4271 & ~n4272 ;
  assign n4274 = n2925 & ~n4273 ;
  assign n4275 = ~n4267 & ~n4274 ;
  assign n4276 = ~n3023 & ~n4275 ;
  assign n4277 = n2925 & ~n4266 ;
  assign n4278 = ~n2925 & ~n4273 ;
  assign n4279 = ~n4277 & ~n4278 ;
  assign n4280 = ~n2979 & ~n4279 ;
  assign n4281 = x82 & n2979 ;
  assign n4282 = ~n4280 & ~n4281 ;
  assign n4283 = n3023 & ~n4282 ;
  assign n4284 = ~n4276 & ~n4283 ;
  assign n4285 = ~n3121 & ~n4284 ;
  assign n4286 = n3023 & ~n4275 ;
  assign n4287 = ~n3023 & ~n4282 ;
  assign n4288 = ~n4286 & ~n4287 ;
  assign n4289 = ~n3073 & ~n4288 ;
  assign n4290 = x50 & n3073 ;
  assign n4291 = ~n4289 & ~n4290 ;
  assign n4292 = n3121 & ~n4291 ;
  assign n4293 = ~n4285 & ~n4292 ;
  assign n4294 = n3219 & ~n4293 ;
  assign n4295 = n3121 & ~n4284 ;
  assign n4296 = ~n3121 & ~n4291 ;
  assign n4297 = ~n4295 & ~n4296 ;
  assign n4298 = ~n3174 & ~n4297 ;
  assign n4299 = x18 & n3174 ;
  assign n4300 = ~n4298 & ~n4299 ;
  assign n4301 = ~n3219 & ~n4300 ;
  assign n4302 = ~n4294 & ~n4301 ;
  assign n4303 = x211 & ~n2630 ;
  assign n4304 = x243 & n2630 ;
  assign n4305 = ~n4303 & ~n4304 ;
  assign n4306 = ~n2728 & ~n4305 ;
  assign n4307 = ~x243 & ~n2630 ;
  assign n4308 = ~x211 & n2630 ;
  assign n4309 = ~n4307 & ~n4308 ;
  assign n4310 = ~n2680 & ~n4309 ;
  assign n4311 = ~x179 & n2680 ;
  assign n4312 = ~n4310 & ~n4311 ;
  assign n4313 = n2728 & n4312 ;
  assign n4314 = ~n4306 & ~n4313 ;
  assign n4315 = ~n2826 & ~n4314 ;
  assign n4316 = n2728 & ~n4305 ;
  assign n4317 = ~n2728 & n4312 ;
  assign n4318 = ~n4316 & ~n4317 ;
  assign n4319 = ~n2782 & ~n4318 ;
  assign n4320 = x147 & n2782 ;
  assign n4321 = ~n4319 & ~n4320 ;
  assign n4322 = n2826 & ~n4321 ;
  assign n4323 = ~n4315 & ~n4322 ;
  assign n4324 = ~n2925 & ~n4323 ;
  assign n4325 = n2826 & ~n4314 ;
  assign n4326 = ~n2826 & ~n4321 ;
  assign n4327 = ~n4325 & ~n4326 ;
  assign n4328 = ~n2880 & ~n4327 ;
  assign n4329 = x115 & n2880 ;
  assign n4330 = ~n4328 & ~n4329 ;
  assign n4331 = n2925 & ~n4330 ;
  assign n4332 = ~n4324 & ~n4331 ;
  assign n4333 = ~n3023 & ~n4332 ;
  assign n4334 = n2925 & ~n4323 ;
  assign n4335 = ~n2925 & ~n4330 ;
  assign n4336 = ~n4334 & ~n4335 ;
  assign n4337 = ~n2979 & ~n4336 ;
  assign n4338 = x83 & n2979 ;
  assign n4339 = ~n4337 & ~n4338 ;
  assign n4340 = n3023 & ~n4339 ;
  assign n4341 = ~n4333 & ~n4340 ;
  assign n4342 = ~n3121 & ~n4341 ;
  assign n4343 = n3023 & ~n4332 ;
  assign n4344 = ~n3023 & ~n4339 ;
  assign n4345 = ~n4343 & ~n4344 ;
  assign n4346 = ~n3073 & ~n4345 ;
  assign n4347 = x51 & n3073 ;
  assign n4348 = ~n4346 & ~n4347 ;
  assign n4349 = n3121 & ~n4348 ;
  assign n4350 = ~n4342 & ~n4349 ;
  assign n4351 = n3219 & ~n4350 ;
  assign n4352 = n3121 & ~n4341 ;
  assign n4353 = ~n3121 & ~n4348 ;
  assign n4354 = ~n4352 & ~n4353 ;
  assign n4355 = ~n3174 & ~n4354 ;
  assign n4356 = x19 & n3174 ;
  assign n4357 = ~n4355 & ~n4356 ;
  assign n4358 = ~n3219 & ~n4357 ;
  assign n4359 = ~n4351 & ~n4358 ;
  assign n4360 = x212 & ~n2630 ;
  assign n4361 = x244 & n2630 ;
  assign n4362 = ~n4360 & ~n4361 ;
  assign n4363 = ~n2728 & ~n4362 ;
  assign n4364 = ~x244 & ~n2630 ;
  assign n4365 = ~x212 & n2630 ;
  assign n4366 = ~n4364 & ~n4365 ;
  assign n4367 = ~n2680 & ~n4366 ;
  assign n4368 = ~x180 & n2680 ;
  assign n4369 = ~n4367 & ~n4368 ;
  assign n4370 = n2728 & n4369 ;
  assign n4371 = ~n4363 & ~n4370 ;
  assign n4372 = ~n2826 & ~n4371 ;
  assign n4373 = n2728 & ~n4362 ;
  assign n4374 = ~n2728 & n4369 ;
  assign n4375 = ~n4373 & ~n4374 ;
  assign n4376 = ~n2782 & ~n4375 ;
  assign n4377 = x148 & n2782 ;
  assign n4378 = ~n4376 & ~n4377 ;
  assign n4379 = n2826 & ~n4378 ;
  assign n4380 = ~n4372 & ~n4379 ;
  assign n4381 = ~n2925 & ~n4380 ;
  assign n4382 = n2826 & ~n4371 ;
  assign n4383 = ~n2826 & ~n4378 ;
  assign n4384 = ~n4382 & ~n4383 ;
  assign n4385 = ~n2880 & ~n4384 ;
  assign n4386 = x116 & n2880 ;
  assign n4387 = ~n4385 & ~n4386 ;
  assign n4388 = n2925 & ~n4387 ;
  assign n4389 = ~n4381 & ~n4388 ;
  assign n4390 = ~n3023 & ~n4389 ;
  assign n4391 = n2925 & ~n4380 ;
  assign n4392 = ~n2925 & ~n4387 ;
  assign n4393 = ~n4391 & ~n4392 ;
  assign n4394 = ~n2979 & ~n4393 ;
  assign n4395 = x84 & n2979 ;
  assign n4396 = ~n4394 & ~n4395 ;
  assign n4397 = n3023 & ~n4396 ;
  assign n4398 = ~n4390 & ~n4397 ;
  assign n4399 = ~n3121 & ~n4398 ;
  assign n4400 = n3023 & ~n4389 ;
  assign n4401 = ~n3023 & ~n4396 ;
  assign n4402 = ~n4400 & ~n4401 ;
  assign n4403 = ~n3073 & ~n4402 ;
  assign n4404 = x52 & n3073 ;
  assign n4405 = ~n4403 & ~n4404 ;
  assign n4406 = n3121 & ~n4405 ;
  assign n4407 = ~n4399 & ~n4406 ;
  assign n4408 = n3219 & ~n4407 ;
  assign n4409 = n3121 & ~n4398 ;
  assign n4410 = ~n3121 & ~n4405 ;
  assign n4411 = ~n4409 & ~n4410 ;
  assign n4412 = ~n3174 & ~n4411 ;
  assign n4413 = x20 & n3174 ;
  assign n4414 = ~n4412 & ~n4413 ;
  assign n4415 = ~n3219 & ~n4414 ;
  assign n4416 = ~n4408 & ~n4415 ;
  assign n4417 = x213 & ~n2630 ;
  assign n4418 = x245 & n2630 ;
  assign n4419 = ~n4417 & ~n4418 ;
  assign n4420 = ~n2728 & ~n4419 ;
  assign n4421 = ~x245 & ~n2630 ;
  assign n4422 = ~x213 & n2630 ;
  assign n4423 = ~n4421 & ~n4422 ;
  assign n4424 = ~n2680 & ~n4423 ;
  assign n4425 = ~x181 & n2680 ;
  assign n4426 = ~n4424 & ~n4425 ;
  assign n4427 = n2728 & n4426 ;
  assign n4428 = ~n4420 & ~n4427 ;
  assign n4429 = ~n2826 & ~n4428 ;
  assign n4430 = n2728 & ~n4419 ;
  assign n4431 = ~n2728 & n4426 ;
  assign n4432 = ~n4430 & ~n4431 ;
  assign n4433 = ~n2782 & ~n4432 ;
  assign n4434 = x149 & n2782 ;
  assign n4435 = ~n4433 & ~n4434 ;
  assign n4436 = n2826 & ~n4435 ;
  assign n4437 = ~n4429 & ~n4436 ;
  assign n4438 = ~n2925 & ~n4437 ;
  assign n4439 = n2826 & ~n4428 ;
  assign n4440 = ~n2826 & ~n4435 ;
  assign n4441 = ~n4439 & ~n4440 ;
  assign n4442 = ~n2880 & ~n4441 ;
  assign n4443 = x117 & n2880 ;
  assign n4444 = ~n4442 & ~n4443 ;
  assign n4445 = n2925 & ~n4444 ;
  assign n4446 = ~n4438 & ~n4445 ;
  assign n4447 = ~n3023 & ~n4446 ;
  assign n4448 = n2925 & ~n4437 ;
  assign n4449 = ~n2925 & ~n4444 ;
  assign n4450 = ~n4448 & ~n4449 ;
  assign n4451 = ~n2979 & ~n4450 ;
  assign n4452 = x85 & n2979 ;
  assign n4453 = ~n4451 & ~n4452 ;
  assign n4454 = n3023 & ~n4453 ;
  assign n4455 = ~n4447 & ~n4454 ;
  assign n4456 = ~n3121 & ~n4455 ;
  assign n4457 = n3023 & ~n4446 ;
  assign n4458 = ~n3023 & ~n4453 ;
  assign n4459 = ~n4457 & ~n4458 ;
  assign n4460 = ~n3073 & ~n4459 ;
  assign n4461 = x53 & n3073 ;
  assign n4462 = ~n4460 & ~n4461 ;
  assign n4463 = n3121 & ~n4462 ;
  assign n4464 = ~n4456 & ~n4463 ;
  assign n4465 = n3219 & ~n4464 ;
  assign n4466 = n3121 & ~n4455 ;
  assign n4467 = ~n3121 & ~n4462 ;
  assign n4468 = ~n4466 & ~n4467 ;
  assign n4469 = ~n3174 & ~n4468 ;
  assign n4470 = x21 & n3174 ;
  assign n4471 = ~n4469 & ~n4470 ;
  assign n4472 = ~n3219 & ~n4471 ;
  assign n4473 = ~n4465 & ~n4472 ;
  assign n4474 = x214 & ~n2630 ;
  assign n4475 = x246 & n2630 ;
  assign n4476 = ~n4474 & ~n4475 ;
  assign n4477 = ~n2728 & ~n4476 ;
  assign n4478 = ~x246 & ~n2630 ;
  assign n4479 = ~x214 & n2630 ;
  assign n4480 = ~n4478 & ~n4479 ;
  assign n4481 = ~n2680 & ~n4480 ;
  assign n4482 = ~x182 & n2680 ;
  assign n4483 = ~n4481 & ~n4482 ;
  assign n4484 = n2728 & n4483 ;
  assign n4485 = ~n4477 & ~n4484 ;
  assign n4486 = ~n2826 & ~n4485 ;
  assign n4487 = n2728 & ~n4476 ;
  assign n4488 = ~n2728 & n4483 ;
  assign n4489 = ~n4487 & ~n4488 ;
  assign n4490 = ~n2782 & ~n4489 ;
  assign n4491 = x150 & n2782 ;
  assign n4492 = ~n4490 & ~n4491 ;
  assign n4493 = n2826 & ~n4492 ;
  assign n4494 = ~n4486 & ~n4493 ;
  assign n4495 = ~n2925 & ~n4494 ;
  assign n4496 = n2826 & ~n4485 ;
  assign n4497 = ~n2826 & ~n4492 ;
  assign n4498 = ~n4496 & ~n4497 ;
  assign n4499 = ~n2880 & ~n4498 ;
  assign n4500 = x118 & n2880 ;
  assign n4501 = ~n4499 & ~n4500 ;
  assign n4502 = n2925 & ~n4501 ;
  assign n4503 = ~n4495 & ~n4502 ;
  assign n4504 = ~n3023 & ~n4503 ;
  assign n4505 = n2925 & ~n4494 ;
  assign n4506 = ~n2925 & ~n4501 ;
  assign n4507 = ~n4505 & ~n4506 ;
  assign n4508 = ~n2979 & ~n4507 ;
  assign n4509 = x86 & n2979 ;
  assign n4510 = ~n4508 & ~n4509 ;
  assign n4511 = n3023 & ~n4510 ;
  assign n4512 = ~n4504 & ~n4511 ;
  assign n4513 = ~n3121 & ~n4512 ;
  assign n4514 = n3023 & ~n4503 ;
  assign n4515 = ~n3023 & ~n4510 ;
  assign n4516 = ~n4514 & ~n4515 ;
  assign n4517 = ~n3073 & ~n4516 ;
  assign n4518 = x54 & n3073 ;
  assign n4519 = ~n4517 & ~n4518 ;
  assign n4520 = n3121 & ~n4519 ;
  assign n4521 = ~n4513 & ~n4520 ;
  assign n4522 = n3219 & ~n4521 ;
  assign n4523 = n3121 & ~n4512 ;
  assign n4524 = ~n3121 & ~n4519 ;
  assign n4525 = ~n4523 & ~n4524 ;
  assign n4526 = ~n3174 & ~n4525 ;
  assign n4527 = x22 & n3174 ;
  assign n4528 = ~n4526 & ~n4527 ;
  assign n4529 = ~n3219 & ~n4528 ;
  assign n4530 = ~n4522 & ~n4529 ;
  assign n4531 = x215 & ~n2630 ;
  assign n4532 = x247 & n2630 ;
  assign n4533 = ~n4531 & ~n4532 ;
  assign n4534 = ~n2728 & ~n4533 ;
  assign n4535 = ~x247 & ~n2630 ;
  assign n4536 = ~x215 & n2630 ;
  assign n4537 = ~n4535 & ~n4536 ;
  assign n4538 = ~n2680 & ~n4537 ;
  assign n4539 = ~x183 & n2680 ;
  assign n4540 = ~n4538 & ~n4539 ;
  assign n4541 = n2728 & n4540 ;
  assign n4542 = ~n4534 & ~n4541 ;
  assign n4543 = ~n2826 & ~n4542 ;
  assign n4544 = n2728 & ~n4533 ;
  assign n4545 = ~n2728 & n4540 ;
  assign n4546 = ~n4544 & ~n4545 ;
  assign n4547 = ~n2782 & ~n4546 ;
  assign n4548 = x151 & n2782 ;
  assign n4549 = ~n4547 & ~n4548 ;
  assign n4550 = n2826 & ~n4549 ;
  assign n4551 = ~n4543 & ~n4550 ;
  assign n4552 = ~n2925 & ~n4551 ;
  assign n4553 = n2826 & ~n4542 ;
  assign n4554 = ~n2826 & ~n4549 ;
  assign n4555 = ~n4553 & ~n4554 ;
  assign n4556 = ~n2880 & ~n4555 ;
  assign n4557 = x119 & n2880 ;
  assign n4558 = ~n4556 & ~n4557 ;
  assign n4559 = n2925 & ~n4558 ;
  assign n4560 = ~n4552 & ~n4559 ;
  assign n4561 = ~n3023 & ~n4560 ;
  assign n4562 = n2925 & ~n4551 ;
  assign n4563 = ~n2925 & ~n4558 ;
  assign n4564 = ~n4562 & ~n4563 ;
  assign n4565 = ~n2979 & ~n4564 ;
  assign n4566 = x87 & n2979 ;
  assign n4567 = ~n4565 & ~n4566 ;
  assign n4568 = n3023 & ~n4567 ;
  assign n4569 = ~n4561 & ~n4568 ;
  assign n4570 = ~n3121 & ~n4569 ;
  assign n4571 = n3023 & ~n4560 ;
  assign n4572 = ~n3023 & ~n4567 ;
  assign n4573 = ~n4571 & ~n4572 ;
  assign n4574 = ~n3073 & ~n4573 ;
  assign n4575 = x55 & n3073 ;
  assign n4576 = ~n4574 & ~n4575 ;
  assign n4577 = n3121 & ~n4576 ;
  assign n4578 = ~n4570 & ~n4577 ;
  assign n4579 = n3219 & ~n4578 ;
  assign n4580 = n3121 & ~n4569 ;
  assign n4581 = ~n3121 & ~n4576 ;
  assign n4582 = ~n4580 & ~n4581 ;
  assign n4583 = ~n3174 & ~n4582 ;
  assign n4584 = x23 & n3174 ;
  assign n4585 = ~n4583 & ~n4584 ;
  assign n4586 = ~n3219 & ~n4585 ;
  assign n4587 = ~n4579 & ~n4586 ;
  assign n4588 = x216 & ~n2630 ;
  assign n4589 = x248 & n2630 ;
  assign n4590 = ~n4588 & ~n4589 ;
  assign n4591 = ~n2728 & ~n4590 ;
  assign n4592 = ~x248 & ~n2630 ;
  assign n4593 = ~x216 & n2630 ;
  assign n4594 = ~n4592 & ~n4593 ;
  assign n4595 = ~n2680 & ~n4594 ;
  assign n4596 = ~x184 & n2680 ;
  assign n4597 = ~n4595 & ~n4596 ;
  assign n4598 = n2728 & n4597 ;
  assign n4599 = ~n4591 & ~n4598 ;
  assign n4600 = ~n2826 & ~n4599 ;
  assign n4601 = n2728 & ~n4590 ;
  assign n4602 = ~n2728 & n4597 ;
  assign n4603 = ~n4601 & ~n4602 ;
  assign n4604 = ~n2782 & ~n4603 ;
  assign n4605 = x152 & n2782 ;
  assign n4606 = ~n4604 & ~n4605 ;
  assign n4607 = n2826 & ~n4606 ;
  assign n4608 = ~n4600 & ~n4607 ;
  assign n4609 = ~n2925 & ~n4608 ;
  assign n4610 = n2826 & ~n4599 ;
  assign n4611 = ~n2826 & ~n4606 ;
  assign n4612 = ~n4610 & ~n4611 ;
  assign n4613 = ~n2880 & ~n4612 ;
  assign n4614 = x120 & n2880 ;
  assign n4615 = ~n4613 & ~n4614 ;
  assign n4616 = n2925 & ~n4615 ;
  assign n4617 = ~n4609 & ~n4616 ;
  assign n4618 = ~n3023 & ~n4617 ;
  assign n4619 = n2925 & ~n4608 ;
  assign n4620 = ~n2925 & ~n4615 ;
  assign n4621 = ~n4619 & ~n4620 ;
  assign n4622 = ~n2979 & ~n4621 ;
  assign n4623 = x88 & n2979 ;
  assign n4624 = ~n4622 & ~n4623 ;
  assign n4625 = n3023 & ~n4624 ;
  assign n4626 = ~n4618 & ~n4625 ;
  assign n4627 = ~n3121 & ~n4626 ;
  assign n4628 = n3023 & ~n4617 ;
  assign n4629 = ~n3023 & ~n4624 ;
  assign n4630 = ~n4628 & ~n4629 ;
  assign n4631 = ~n3073 & ~n4630 ;
  assign n4632 = x56 & n3073 ;
  assign n4633 = ~n4631 & ~n4632 ;
  assign n4634 = n3121 & ~n4633 ;
  assign n4635 = ~n4627 & ~n4634 ;
  assign n4636 = n3219 & ~n4635 ;
  assign n4637 = n3121 & ~n4626 ;
  assign n4638 = ~n3121 & ~n4633 ;
  assign n4639 = ~n4637 & ~n4638 ;
  assign n4640 = ~n3174 & ~n4639 ;
  assign n4641 = x24 & n3174 ;
  assign n4642 = ~n4640 & ~n4641 ;
  assign n4643 = ~n3219 & ~n4642 ;
  assign n4644 = ~n4636 & ~n4643 ;
  assign n4645 = x217 & ~n2630 ;
  assign n4646 = x249 & n2630 ;
  assign n4647 = ~n4645 & ~n4646 ;
  assign n4648 = ~n2728 & ~n4647 ;
  assign n4649 = ~x249 & ~n2630 ;
  assign n4650 = ~x217 & n2630 ;
  assign n4651 = ~n4649 & ~n4650 ;
  assign n4652 = ~n2680 & ~n4651 ;
  assign n4653 = ~x185 & n2680 ;
  assign n4654 = ~n4652 & ~n4653 ;
  assign n4655 = n2728 & n4654 ;
  assign n4656 = ~n4648 & ~n4655 ;
  assign n4657 = ~n2826 & ~n4656 ;
  assign n4658 = n2728 & ~n4647 ;
  assign n4659 = ~n2728 & n4654 ;
  assign n4660 = ~n4658 & ~n4659 ;
  assign n4661 = ~n2782 & ~n4660 ;
  assign n4662 = x153 & n2782 ;
  assign n4663 = ~n4661 & ~n4662 ;
  assign n4664 = n2826 & ~n4663 ;
  assign n4665 = ~n4657 & ~n4664 ;
  assign n4666 = ~n2925 & ~n4665 ;
  assign n4667 = n2826 & ~n4656 ;
  assign n4668 = ~n2826 & ~n4663 ;
  assign n4669 = ~n4667 & ~n4668 ;
  assign n4670 = ~n2880 & ~n4669 ;
  assign n4671 = x121 & n2880 ;
  assign n4672 = ~n4670 & ~n4671 ;
  assign n4673 = n2925 & ~n4672 ;
  assign n4674 = ~n4666 & ~n4673 ;
  assign n4675 = ~n3023 & ~n4674 ;
  assign n4676 = n2925 & ~n4665 ;
  assign n4677 = ~n2925 & ~n4672 ;
  assign n4678 = ~n4676 & ~n4677 ;
  assign n4679 = ~n2979 & ~n4678 ;
  assign n4680 = x89 & n2979 ;
  assign n4681 = ~n4679 & ~n4680 ;
  assign n4682 = n3023 & ~n4681 ;
  assign n4683 = ~n4675 & ~n4682 ;
  assign n4684 = ~n3121 & ~n4683 ;
  assign n4685 = n3023 & ~n4674 ;
  assign n4686 = ~n3023 & ~n4681 ;
  assign n4687 = ~n4685 & ~n4686 ;
  assign n4688 = ~n3073 & ~n4687 ;
  assign n4689 = x57 & n3073 ;
  assign n4690 = ~n4688 & ~n4689 ;
  assign n4691 = n3121 & ~n4690 ;
  assign n4692 = ~n4684 & ~n4691 ;
  assign n4693 = n3219 & ~n4692 ;
  assign n4694 = n3121 & ~n4683 ;
  assign n4695 = ~n3121 & ~n4690 ;
  assign n4696 = ~n4694 & ~n4695 ;
  assign n4697 = ~n3174 & ~n4696 ;
  assign n4698 = x25 & n3174 ;
  assign n4699 = ~n4697 & ~n4698 ;
  assign n4700 = ~n3219 & ~n4699 ;
  assign n4701 = ~n4693 & ~n4700 ;
  assign n4702 = x218 & ~n2630 ;
  assign n4703 = x250 & n2630 ;
  assign n4704 = ~n4702 & ~n4703 ;
  assign n4705 = ~n2728 & ~n4704 ;
  assign n4706 = ~x250 & ~n2630 ;
  assign n4707 = ~x218 & n2630 ;
  assign n4708 = ~n4706 & ~n4707 ;
  assign n4709 = ~n2680 & ~n4708 ;
  assign n4710 = ~x186 & n2680 ;
  assign n4711 = ~n4709 & ~n4710 ;
  assign n4712 = n2728 & n4711 ;
  assign n4713 = ~n4705 & ~n4712 ;
  assign n4714 = ~n2826 & ~n4713 ;
  assign n4715 = n2728 & ~n4704 ;
  assign n4716 = ~n2728 & n4711 ;
  assign n4717 = ~n4715 & ~n4716 ;
  assign n4718 = ~n2782 & ~n4717 ;
  assign n4719 = x154 & n2782 ;
  assign n4720 = ~n4718 & ~n4719 ;
  assign n4721 = n2826 & ~n4720 ;
  assign n4722 = ~n4714 & ~n4721 ;
  assign n4723 = ~n2925 & ~n4722 ;
  assign n4724 = n2826 & ~n4713 ;
  assign n4725 = ~n2826 & ~n4720 ;
  assign n4726 = ~n4724 & ~n4725 ;
  assign n4727 = ~n2880 & ~n4726 ;
  assign n4728 = x122 & n2880 ;
  assign n4729 = ~n4727 & ~n4728 ;
  assign n4730 = n2925 & ~n4729 ;
  assign n4731 = ~n4723 & ~n4730 ;
  assign n4732 = ~n3023 & ~n4731 ;
  assign n4733 = n2925 & ~n4722 ;
  assign n4734 = ~n2925 & ~n4729 ;
  assign n4735 = ~n4733 & ~n4734 ;
  assign n4736 = ~n2979 & ~n4735 ;
  assign n4737 = x90 & n2979 ;
  assign n4738 = ~n4736 & ~n4737 ;
  assign n4739 = n3023 & ~n4738 ;
  assign n4740 = ~n4732 & ~n4739 ;
  assign n4741 = ~n3121 & ~n4740 ;
  assign n4742 = n3023 & ~n4731 ;
  assign n4743 = ~n3023 & ~n4738 ;
  assign n4744 = ~n4742 & ~n4743 ;
  assign n4745 = ~n3073 & ~n4744 ;
  assign n4746 = x58 & n3073 ;
  assign n4747 = ~n4745 & ~n4746 ;
  assign n4748 = n3121 & ~n4747 ;
  assign n4749 = ~n4741 & ~n4748 ;
  assign n4750 = n3219 & ~n4749 ;
  assign n4751 = n3121 & ~n4740 ;
  assign n4752 = ~n3121 & ~n4747 ;
  assign n4753 = ~n4751 & ~n4752 ;
  assign n4754 = ~n3174 & ~n4753 ;
  assign n4755 = x26 & n3174 ;
  assign n4756 = ~n4754 & ~n4755 ;
  assign n4757 = ~n3219 & ~n4756 ;
  assign n4758 = ~n4750 & ~n4757 ;
  assign n4759 = x219 & ~n2630 ;
  assign n4760 = x251 & n2630 ;
  assign n4761 = ~n4759 & ~n4760 ;
  assign n4762 = ~n2728 & ~n4761 ;
  assign n4763 = ~x251 & ~n2630 ;
  assign n4764 = ~x219 & n2630 ;
  assign n4765 = ~n4763 & ~n4764 ;
  assign n4766 = ~n2680 & ~n4765 ;
  assign n4767 = ~x187 & n2680 ;
  assign n4768 = ~n4766 & ~n4767 ;
  assign n4769 = n2728 & n4768 ;
  assign n4770 = ~n4762 & ~n4769 ;
  assign n4771 = ~n2826 & ~n4770 ;
  assign n4772 = n2728 & ~n4761 ;
  assign n4773 = ~n2728 & n4768 ;
  assign n4774 = ~n4772 & ~n4773 ;
  assign n4775 = ~n2782 & ~n4774 ;
  assign n4776 = x155 & n2782 ;
  assign n4777 = ~n4775 & ~n4776 ;
  assign n4778 = n2826 & ~n4777 ;
  assign n4779 = ~n4771 & ~n4778 ;
  assign n4780 = ~n2925 & ~n4779 ;
  assign n4781 = n2826 & ~n4770 ;
  assign n4782 = ~n2826 & ~n4777 ;
  assign n4783 = ~n4781 & ~n4782 ;
  assign n4784 = ~n2880 & ~n4783 ;
  assign n4785 = x123 & n2880 ;
  assign n4786 = ~n4784 & ~n4785 ;
  assign n4787 = n2925 & ~n4786 ;
  assign n4788 = ~n4780 & ~n4787 ;
  assign n4789 = ~n3023 & ~n4788 ;
  assign n4790 = n2925 & ~n4779 ;
  assign n4791 = ~n2925 & ~n4786 ;
  assign n4792 = ~n4790 & ~n4791 ;
  assign n4793 = ~n2979 & ~n4792 ;
  assign n4794 = x91 & n2979 ;
  assign n4795 = ~n4793 & ~n4794 ;
  assign n4796 = n3023 & ~n4795 ;
  assign n4797 = ~n4789 & ~n4796 ;
  assign n4798 = ~n3121 & ~n4797 ;
  assign n4799 = n3023 & ~n4788 ;
  assign n4800 = ~n3023 & ~n4795 ;
  assign n4801 = ~n4799 & ~n4800 ;
  assign n4802 = ~n3073 & ~n4801 ;
  assign n4803 = x59 & n3073 ;
  assign n4804 = ~n4802 & ~n4803 ;
  assign n4805 = n3121 & ~n4804 ;
  assign n4806 = ~n4798 & ~n4805 ;
  assign n4807 = n3219 & ~n4806 ;
  assign n4808 = n3121 & ~n4797 ;
  assign n4809 = ~n3121 & ~n4804 ;
  assign n4810 = ~n4808 & ~n4809 ;
  assign n4811 = ~n3174 & ~n4810 ;
  assign n4812 = x27 & n3174 ;
  assign n4813 = ~n4811 & ~n4812 ;
  assign n4814 = ~n3219 & ~n4813 ;
  assign n4815 = ~n4807 & ~n4814 ;
  assign n4816 = x220 & ~n2630 ;
  assign n4817 = x252 & n2630 ;
  assign n4818 = ~n4816 & ~n4817 ;
  assign n4819 = ~n2728 & ~n4818 ;
  assign n4820 = ~x252 & ~n2630 ;
  assign n4821 = ~x220 & n2630 ;
  assign n4822 = ~n4820 & ~n4821 ;
  assign n4823 = ~n2680 & ~n4822 ;
  assign n4824 = ~x188 & n2680 ;
  assign n4825 = ~n4823 & ~n4824 ;
  assign n4826 = n2728 & n4825 ;
  assign n4827 = ~n4819 & ~n4826 ;
  assign n4828 = ~n2826 & ~n4827 ;
  assign n4829 = n2728 & ~n4818 ;
  assign n4830 = ~n2728 & n4825 ;
  assign n4831 = ~n4829 & ~n4830 ;
  assign n4832 = ~n2782 & ~n4831 ;
  assign n4833 = x156 & n2782 ;
  assign n4834 = ~n4832 & ~n4833 ;
  assign n4835 = n2826 & ~n4834 ;
  assign n4836 = ~n4828 & ~n4835 ;
  assign n4837 = ~n2925 & ~n4836 ;
  assign n4838 = n2826 & ~n4827 ;
  assign n4839 = ~n2826 & ~n4834 ;
  assign n4840 = ~n4838 & ~n4839 ;
  assign n4841 = ~n2880 & ~n4840 ;
  assign n4842 = x124 & n2880 ;
  assign n4843 = ~n4841 & ~n4842 ;
  assign n4844 = n2925 & ~n4843 ;
  assign n4845 = ~n4837 & ~n4844 ;
  assign n4846 = ~n3023 & ~n4845 ;
  assign n4847 = n2925 & ~n4836 ;
  assign n4848 = ~n2925 & ~n4843 ;
  assign n4849 = ~n4847 & ~n4848 ;
  assign n4850 = ~n2979 & ~n4849 ;
  assign n4851 = x92 & n2979 ;
  assign n4852 = ~n4850 & ~n4851 ;
  assign n4853 = n3023 & ~n4852 ;
  assign n4854 = ~n4846 & ~n4853 ;
  assign n4855 = ~n3121 & ~n4854 ;
  assign n4856 = n3023 & ~n4845 ;
  assign n4857 = ~n3023 & ~n4852 ;
  assign n4858 = ~n4856 & ~n4857 ;
  assign n4859 = ~n3073 & ~n4858 ;
  assign n4860 = x60 & n3073 ;
  assign n4861 = ~n4859 & ~n4860 ;
  assign n4862 = n3121 & ~n4861 ;
  assign n4863 = ~n4855 & ~n4862 ;
  assign n4864 = n3219 & ~n4863 ;
  assign n4865 = n3121 & ~n4854 ;
  assign n4866 = ~n3121 & ~n4861 ;
  assign n4867 = ~n4865 & ~n4866 ;
  assign n4868 = ~n3174 & ~n4867 ;
  assign n4869 = x28 & n3174 ;
  assign n4870 = ~n4868 & ~n4869 ;
  assign n4871 = ~n3219 & ~n4870 ;
  assign n4872 = ~n4864 & ~n4871 ;
  assign n4873 = x221 & ~n2630 ;
  assign n4874 = x253 & n2630 ;
  assign n4875 = ~n4873 & ~n4874 ;
  assign n4876 = ~n2728 & ~n4875 ;
  assign n4877 = ~x253 & ~n2630 ;
  assign n4878 = ~x221 & n2630 ;
  assign n4879 = ~n4877 & ~n4878 ;
  assign n4880 = ~n2680 & ~n4879 ;
  assign n4881 = ~x189 & n2680 ;
  assign n4882 = ~n4880 & ~n4881 ;
  assign n4883 = n2728 & n4882 ;
  assign n4884 = ~n4876 & ~n4883 ;
  assign n4885 = ~n2826 & ~n4884 ;
  assign n4886 = n2728 & ~n4875 ;
  assign n4887 = ~n2728 & n4882 ;
  assign n4888 = ~n4886 & ~n4887 ;
  assign n4889 = ~n2782 & ~n4888 ;
  assign n4890 = x157 & n2782 ;
  assign n4891 = ~n4889 & ~n4890 ;
  assign n4892 = n2826 & ~n4891 ;
  assign n4893 = ~n4885 & ~n4892 ;
  assign n4894 = ~n2925 & ~n4893 ;
  assign n4895 = n2826 & ~n4884 ;
  assign n4896 = ~n2826 & ~n4891 ;
  assign n4897 = ~n4895 & ~n4896 ;
  assign n4898 = ~n2880 & ~n4897 ;
  assign n4899 = x125 & n2880 ;
  assign n4900 = ~n4898 & ~n4899 ;
  assign n4901 = n2925 & ~n4900 ;
  assign n4902 = ~n4894 & ~n4901 ;
  assign n4903 = ~n3023 & ~n4902 ;
  assign n4904 = n2925 & ~n4893 ;
  assign n4905 = ~n2925 & ~n4900 ;
  assign n4906 = ~n4904 & ~n4905 ;
  assign n4907 = ~n2979 & ~n4906 ;
  assign n4908 = x93 & n2979 ;
  assign n4909 = ~n4907 & ~n4908 ;
  assign n4910 = n3023 & ~n4909 ;
  assign n4911 = ~n4903 & ~n4910 ;
  assign n4912 = ~n3121 & ~n4911 ;
  assign n4913 = n3023 & ~n4902 ;
  assign n4914 = ~n3023 & ~n4909 ;
  assign n4915 = ~n4913 & ~n4914 ;
  assign n4916 = ~n3073 & ~n4915 ;
  assign n4917 = x61 & n3073 ;
  assign n4918 = ~n4916 & ~n4917 ;
  assign n4919 = n3121 & ~n4918 ;
  assign n4920 = ~n4912 & ~n4919 ;
  assign n4921 = n3219 & ~n4920 ;
  assign n4922 = n3121 & ~n4911 ;
  assign n4923 = ~n3121 & ~n4918 ;
  assign n4924 = ~n4922 & ~n4923 ;
  assign n4925 = ~n3174 & ~n4924 ;
  assign n4926 = x29 & n3174 ;
  assign n4927 = ~n4925 & ~n4926 ;
  assign n4928 = ~n3219 & ~n4927 ;
  assign n4929 = ~n4921 & ~n4928 ;
  assign n4930 = x222 & ~n2630 ;
  assign n4931 = x254 & n2630 ;
  assign n4932 = ~n4930 & ~n4931 ;
  assign n4933 = ~n2728 & ~n4932 ;
  assign n4934 = ~x254 & ~n2630 ;
  assign n4935 = ~x222 & n2630 ;
  assign n4936 = ~n4934 & ~n4935 ;
  assign n4937 = ~n2680 & ~n4936 ;
  assign n4938 = ~x190 & n2680 ;
  assign n4939 = ~n4937 & ~n4938 ;
  assign n4940 = n2728 & n4939 ;
  assign n4941 = ~n4933 & ~n4940 ;
  assign n4942 = ~n2826 & ~n4941 ;
  assign n4943 = n2728 & ~n4932 ;
  assign n4944 = ~n2728 & n4939 ;
  assign n4945 = ~n4943 & ~n4944 ;
  assign n4946 = ~n2782 & ~n4945 ;
  assign n4947 = x158 & n2782 ;
  assign n4948 = ~n4946 & ~n4947 ;
  assign n4949 = n2826 & ~n4948 ;
  assign n4950 = ~n4942 & ~n4949 ;
  assign n4951 = ~n2925 & ~n4950 ;
  assign n4952 = n2826 & ~n4941 ;
  assign n4953 = ~n2826 & ~n4948 ;
  assign n4954 = ~n4952 & ~n4953 ;
  assign n4955 = ~n2880 & ~n4954 ;
  assign n4956 = x126 & n2880 ;
  assign n4957 = ~n4955 & ~n4956 ;
  assign n4958 = n2925 & ~n4957 ;
  assign n4959 = ~n4951 & ~n4958 ;
  assign n4960 = ~n3023 & ~n4959 ;
  assign n4961 = n2925 & ~n4950 ;
  assign n4962 = ~n2925 & ~n4957 ;
  assign n4963 = ~n4961 & ~n4962 ;
  assign n4964 = ~n2979 & ~n4963 ;
  assign n4965 = x94 & n2979 ;
  assign n4966 = ~n4964 & ~n4965 ;
  assign n4967 = n3023 & ~n4966 ;
  assign n4968 = ~n4960 & ~n4967 ;
  assign n4969 = ~n3121 & ~n4968 ;
  assign n4970 = n3023 & ~n4959 ;
  assign n4971 = ~n3023 & ~n4966 ;
  assign n4972 = ~n4970 & ~n4971 ;
  assign n4973 = ~n3073 & ~n4972 ;
  assign n4974 = x62 & n3073 ;
  assign n4975 = ~n4973 & ~n4974 ;
  assign n4976 = n3121 & ~n4975 ;
  assign n4977 = ~n4969 & ~n4976 ;
  assign n4978 = n3219 & ~n4977 ;
  assign n4979 = n3121 & ~n4968 ;
  assign n4980 = ~n3121 & ~n4975 ;
  assign n4981 = ~n4979 & ~n4980 ;
  assign n4982 = ~n3174 & ~n4981 ;
  assign n4983 = x30 & n3174 ;
  assign n4984 = ~n4982 & ~n4983 ;
  assign n4985 = ~n3219 & ~n4984 ;
  assign n4986 = ~n4978 & ~n4985 ;
  assign n4987 = x223 & ~n2630 ;
  assign n4988 = x255 & n2630 ;
  assign n4989 = ~n4987 & ~n4988 ;
  assign n4990 = ~n2728 & ~n4989 ;
  assign n4991 = ~x255 & ~n2630 ;
  assign n4992 = ~x223 & n2630 ;
  assign n4993 = ~n4991 & ~n4992 ;
  assign n4994 = ~n2680 & ~n4993 ;
  assign n4995 = ~x191 & n2680 ;
  assign n4996 = ~n4994 & ~n4995 ;
  assign n4997 = n2728 & n4996 ;
  assign n4998 = ~n4990 & ~n4997 ;
  assign n4999 = ~n2826 & ~n4998 ;
  assign n5000 = n2728 & ~n4989 ;
  assign n5001 = ~n2728 & n4996 ;
  assign n5002 = ~n5000 & ~n5001 ;
  assign n5003 = ~n2782 & ~n5002 ;
  assign n5004 = x159 & n2782 ;
  assign n5005 = ~n5003 & ~n5004 ;
  assign n5006 = n2826 & ~n5005 ;
  assign n5007 = ~n4999 & ~n5006 ;
  assign n5008 = ~n2925 & ~n5007 ;
  assign n5009 = n2826 & ~n4998 ;
  assign n5010 = ~n2826 & ~n5005 ;
  assign n5011 = ~n5009 & ~n5010 ;
  assign n5012 = ~n2880 & ~n5011 ;
  assign n5013 = x127 & n2880 ;
  assign n5014 = ~n5012 & ~n5013 ;
  assign n5015 = n2925 & ~n5014 ;
  assign n5016 = ~n5008 & ~n5015 ;
  assign n5017 = ~n3023 & ~n5016 ;
  assign n5018 = n2925 & ~n5007 ;
  assign n5019 = ~n2925 & ~n5014 ;
  assign n5020 = ~n5018 & ~n5019 ;
  assign n5021 = ~n2979 & ~n5020 ;
  assign n5022 = x95 & n2979 ;
  assign n5023 = ~n5021 & ~n5022 ;
  assign n5024 = n3023 & ~n5023 ;
  assign n5025 = ~n5017 & ~n5024 ;
  assign n5026 = ~n3121 & ~n5025 ;
  assign n5027 = n3023 & ~n5016 ;
  assign n5028 = ~n3023 & ~n5023 ;
  assign n5029 = ~n5027 & ~n5028 ;
  assign n5030 = ~n3073 & ~n5029 ;
  assign n5031 = x63 & n3073 ;
  assign n5032 = ~n5030 & ~n5031 ;
  assign n5033 = n3121 & ~n5032 ;
  assign n5034 = ~n5026 & ~n5033 ;
  assign n5035 = n3219 & ~n5034 ;
  assign n5036 = n3121 & ~n5025 ;
  assign n5037 = ~n3121 & ~n5032 ;
  assign n5038 = ~n5036 & ~n5037 ;
  assign n5039 = ~n3174 & ~n5038 ;
  assign n5040 = x31 & n3174 ;
  assign n5041 = ~n5039 & ~n5040 ;
  assign n5042 = ~n3219 & ~n5041 ;
  assign n5043 = ~n5035 & ~n5042 ;
  assign n5044 = ~n3219 & ~n3267 ;
  assign n5045 = n3219 & ~n3274 ;
  assign n5046 = ~n5044 & ~n5045 ;
  assign n5047 = ~n3219 & ~n3324 ;
  assign n5048 = n3219 & ~n3331 ;
  assign n5049 = ~n5047 & ~n5048 ;
  assign n5050 = ~n3219 & ~n3381 ;
  assign n5051 = n3219 & ~n3388 ;
  assign n5052 = ~n5050 & ~n5051 ;
  assign n5053 = ~n3219 & ~n3438 ;
  assign n5054 = n3219 & ~n3445 ;
  assign n5055 = ~n5053 & ~n5054 ;
  assign n5056 = ~n3219 & ~n3495 ;
  assign n5057 = n3219 & ~n3502 ;
  assign n5058 = ~n5056 & ~n5057 ;
  assign n5059 = ~n3219 & ~n3552 ;
  assign n5060 = n3219 & ~n3559 ;
  assign n5061 = ~n5059 & ~n5060 ;
  assign n5062 = ~n3219 & ~n3609 ;
  assign n5063 = n3219 & ~n3616 ;
  assign n5064 = ~n5062 & ~n5063 ;
  assign n5065 = ~n3219 & ~n3666 ;
  assign n5066 = n3219 & ~n3673 ;
  assign n5067 = ~n5065 & ~n5066 ;
  assign n5068 = ~n3219 & ~n3723 ;
  assign n5069 = n3219 & ~n3730 ;
  assign n5070 = ~n5068 & ~n5069 ;
  assign n5071 = ~n3219 & ~n3780 ;
  assign n5072 = n3219 & ~n3787 ;
  assign n5073 = ~n5071 & ~n5072 ;
  assign n5074 = ~n3219 & ~n3837 ;
  assign n5075 = n3219 & ~n3844 ;
  assign n5076 = ~n5074 & ~n5075 ;
  assign n5077 = ~n3219 & ~n3894 ;
  assign n5078 = n3219 & ~n3901 ;
  assign n5079 = ~n5077 & ~n5078 ;
  assign n5080 = ~n3219 & ~n3951 ;
  assign n5081 = n3219 & ~n3958 ;
  assign n5082 = ~n5080 & ~n5081 ;
  assign n5083 = ~n3219 & ~n4008 ;
  assign n5084 = n3219 & ~n4015 ;
  assign n5085 = ~n5083 & ~n5084 ;
  assign n5086 = ~n3219 & ~n4065 ;
  assign n5087 = n3219 & ~n4072 ;
  assign n5088 = ~n5086 & ~n5087 ;
  assign n5089 = ~n3219 & ~n4122 ;
  assign n5090 = n3219 & ~n4129 ;
  assign n5091 = ~n5089 & ~n5090 ;
  assign n5092 = ~n3219 & ~n4179 ;
  assign n5093 = n3219 & ~n4186 ;
  assign n5094 = ~n5092 & ~n5093 ;
  assign n5095 = ~n3219 & ~n4236 ;
  assign n5096 = n3219 & ~n4243 ;
  assign n5097 = ~n5095 & ~n5096 ;
  assign n5098 = ~n3219 & ~n4293 ;
  assign n5099 = n3219 & ~n4300 ;
  assign n5100 = ~n5098 & ~n5099 ;
  assign n5101 = ~n3219 & ~n4350 ;
  assign n5102 = n3219 & ~n4357 ;
  assign n5103 = ~n5101 & ~n5102 ;
  assign n5104 = ~n3219 & ~n4407 ;
  assign n5105 = n3219 & ~n4414 ;
  assign n5106 = ~n5104 & ~n5105 ;
  assign n5107 = ~n3219 & ~n4464 ;
  assign n5108 = n3219 & ~n4471 ;
  assign n5109 = ~n5107 & ~n5108 ;
  assign n5110 = ~n3219 & ~n4521 ;
  assign n5111 = n3219 & ~n4528 ;
  assign n5112 = ~n5110 & ~n5111 ;
  assign n5113 = ~n3219 & ~n4578 ;
  assign n5114 = n3219 & ~n4585 ;
  assign n5115 = ~n5113 & ~n5114 ;
  assign n5116 = ~n3219 & ~n4635 ;
  assign n5117 = n3219 & ~n4642 ;
  assign n5118 = ~n5116 & ~n5117 ;
  assign n5119 = ~n3219 & ~n4692 ;
  assign n5120 = n3219 & ~n4699 ;
  assign n5121 = ~n5119 & ~n5120 ;
  assign n5122 = ~n3219 & ~n4749 ;
  assign n5123 = n3219 & ~n4756 ;
  assign n5124 = ~n5122 & ~n5123 ;
  assign n5125 = ~n3219 & ~n4806 ;
  assign n5126 = n3219 & ~n4813 ;
  assign n5127 = ~n5125 & ~n5126 ;
  assign n5128 = ~n3219 & ~n4863 ;
  assign n5129 = n3219 & ~n4870 ;
  assign n5130 = ~n5128 & ~n5129 ;
  assign n5131 = ~n3219 & ~n4920 ;
  assign n5132 = n3219 & ~n4927 ;
  assign n5133 = ~n5131 & ~n5132 ;
  assign n5134 = ~n3219 & ~n4977 ;
  assign n5135 = n3219 & ~n4984 ;
  assign n5136 = ~n5134 & ~n5135 ;
  assign n5137 = ~n3219 & ~n5034 ;
  assign n5138 = n3219 & ~n5041 ;
  assign n5139 = ~n5137 & ~n5138 ;
  assign y0 = ~n3276 ;
  assign y1 = ~n3333 ;
  assign y2 = ~n3390 ;
  assign y3 = ~n3447 ;
  assign y4 = ~n3504 ;
  assign y5 = ~n3561 ;
  assign y6 = ~n3618 ;
  assign y7 = ~n3675 ;
  assign y8 = ~n3732 ;
  assign y9 = ~n3789 ;
  assign y10 = ~n3846 ;
  assign y11 = ~n3903 ;
  assign y12 = ~n3960 ;
  assign y13 = ~n4017 ;
  assign y14 = ~n4074 ;
  assign y15 = ~n4131 ;
  assign y16 = ~n4188 ;
  assign y17 = ~n4245 ;
  assign y18 = ~n4302 ;
  assign y19 = ~n4359 ;
  assign y20 = ~n4416 ;
  assign y21 = ~n4473 ;
  assign y22 = ~n4530 ;
  assign y23 = ~n4587 ;
  assign y24 = ~n4644 ;
  assign y25 = ~n4701 ;
  assign y26 = ~n4758 ;
  assign y27 = ~n4815 ;
  assign y28 = ~n4872 ;
  assign y29 = ~n4929 ;
  assign y30 = ~n4986 ;
  assign y31 = ~n5043 ;
  assign y32 = ~n5046 ;
  assign y33 = ~n5049 ;
  assign y34 = ~n5052 ;
  assign y35 = ~n5055 ;
  assign y36 = ~n5058 ;
  assign y37 = ~n5061 ;
  assign y38 = ~n5064 ;
  assign y39 = ~n5067 ;
  assign y40 = ~n5070 ;
  assign y41 = ~n5073 ;
  assign y42 = ~n5076 ;
  assign y43 = ~n5079 ;
  assign y44 = ~n5082 ;
  assign y45 = ~n5085 ;
  assign y46 = ~n5088 ;
  assign y47 = ~n5091 ;
  assign y48 = ~n5094 ;
  assign y49 = ~n5097 ;
  assign y50 = ~n5100 ;
  assign y51 = ~n5103 ;
  assign y52 = ~n5106 ;
  assign y53 = ~n5109 ;
  assign y54 = ~n5112 ;
  assign y55 = ~n5115 ;
  assign y56 = ~n5118 ;
  assign y57 = ~n5121 ;
  assign y58 = ~n5124 ;
  assign y59 = ~n5127 ;
  assign y60 = ~n5130 ;
  assign y61 = ~n5133 ;
  assign y62 = ~n5136 ;
  assign y63 = ~n5139 ;
endmodule
