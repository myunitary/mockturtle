module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 ;
  assign n14 = ~x6 & ~x7 ;
  assign n9 = ~x0 & ~x1 ;
  assign n10 = ~x2 & ~x3 ;
  assign n11 = n9 & n10 ;
  assign n12 = ~x4 & ~x5 ;
  assign n13 = n11 & n12 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = x6 & x7 ;
  assign n17 = x4 & x5 ;
  assign n18 = n16 & n17 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = x0 & x1 ;
  assign n22 = x2 & x3 ;
  assign n23 = n21 & n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = ~n20 & ~n25 ;
  assign n29 = n12 ^ n10 ;
  assign n30 = n29 ^ n12 ;
  assign n27 = n12 ^ n9 ;
  assign n28 = n27 ^ n12 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n28 ^ n12 ;
  assign n33 = n31 & n32 ;
  assign n34 = n33 ^ n28 ;
  assign n35 = n26 & n34 ;
  assign n36 = n15 & n35 ;
  assign y0 = n36 ;
endmodule
