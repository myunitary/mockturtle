// Benchmark "cardio" written by ABC on Wed Dec 27 23:19:07 2023

module top ( 
    i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10, i_11, i_12, i_13, i_14,
    i_15, i_16, i_17, i_18, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26,
    i_27, i_28, i_29, i_30, i_31, i_32, i_33, i_34, i_35, i_36, i_37, i_38,
    i_39, i_40, i_41, i_42, i_43, i_44, i_45, i_46, i_47, i_48, i_49, i_50,
    i_51, i_52, i_53, i_54, i_55, i_56, i_57, i_58, i_59, i_60, i_61, i_62,
    i_63, i_64, i_65, i_66, i_67, i_68, i_69, i_70, i_71, i_72, i_73, i_74,
    i_75, i_76, i_77, i_78, i_79, i_80, i_81, i_82, i_83, i_84, i_85, i_86,
    i_87, i_88, i_89, i_90, i_91, i_92, i_93, i_94, i_95, i_96, i_97, i_98,
    i_99, i_100, i_101, i_102, i_103, i_104, i_105, i_106, i_107, i_108,
    i_109, i_110, i_111, i_112, i_113,
    m_0, m_1, m_2, m_3  );
  input  i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10, i_11, i_12, i_13,
    i_14, i_15, i_16, i_17, i_18, i_19, i_20, i_21, i_22, i_23, i_24, i_25,
    i_26, i_27, i_28, i_29, i_30, i_31, i_32, i_33, i_34, i_35, i_36, i_37,
    i_38, i_39, i_40, i_41, i_42, i_43, i_44, i_45, i_46, i_47, i_48, i_49,
    i_50, i_51, i_52, i_53, i_54, i_55, i_56, i_57, i_58, i_59, i_60, i_61,
    i_62, i_63, i_64, i_65, i_66, i_67, i_68, i_69, i_70, i_71, i_72, i_73,
    i_74, i_75, i_76, i_77, i_78, i_79, i_80, i_81, i_82, i_83, i_84, i_85,
    i_86, i_87, i_88, i_89, i_90, i_91, i_92, i_93, i_94, i_95, i_96, i_97,
    i_98, i_99, i_100, i_101, i_102, i_103, i_104, i_105, i_106, i_107,
    i_108, i_109, i_110, i_111, i_112, i_113;
  output m_0, m_1, m_2, m_3;
  wire new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n431_;
  assign new_n117_ = ~i_113 ^ ~i_57;
  assign new_n118_ = ~i_112 ^ ~i_56;
  assign new_n119_ = new_n118_ & new_n117_;
  assign new_n120_ = ~i_111 ^ ~i_55;
  assign new_n121_ = ~new_n120_;
  assign new_n122_ = ~i_110 ^ ~i_54;
  assign new_n123_ = ~new_n122_;
  assign new_n124_ = new_n123_ & new_n121_;
  assign new_n125_ = new_n124_ & new_n119_;
  assign new_n126_ = ~new_n125_;
  assign new_n127_ = new_n123_ & new_n120_;
  assign new_n128_ = ~new_n127_ ^ ~new_n123_;
  assign new_n129_ = ~new_n128_ ^ ~new_n126_;
  assign new_n130_ = ~i_107 ^ ~i_51;
  assign new_n131_ = ~new_n130_;
  assign new_n132_ = ~i_50;
  assign new_n133_ = ~i_106 ^ ~new_n132_;
  assign new_n134_ = new_n133_ & new_n131_;
  assign new_n135_ = ~i_109 ^ ~i_53;
  assign new_n136_ = ~new_n135_;
  assign new_n137_ = ~i_108 ^ ~i_52;
  assign new_n138_ = ~new_n137_;
  assign new_n139_ = new_n138_ & new_n136_;
  assign new_n140_ = new_n139_ & new_n134_;
  assign new_n141_ = new_n140_ & new_n129_;
  assign new_n142_ = ~new_n141_;
  assign new_n143_ = new_n138_ & new_n135_;
  assign new_n144_ = ~new_n143_ ^ ~new_n137_;
  assign new_n145_ = new_n144_ & new_n134_;
  assign new_n146_ = new_n133_ & new_n130_;
  assign new_n147_ = ~new_n146_ ^ ~new_n133_;
  assign new_n148_ = ~new_n147_ ^ ~new_n145_;
  assign new_n149_ = ~new_n148_ ^ ~new_n142_;
  assign new_n150_ = ~i_65 ^ ~i_9;
  assign new_n151_ = ~new_n150_;
  assign new_n152_ = new_n151_ & new_n149_;
  assign new_n153_ = ~new_n148_;
  assign new_n154_ = ~new_n128_;
  assign new_n155_ = new_n140_ & new_n154_;
  assign new_n156_ = ~new_n155_ ^ ~new_n153_;
  assign new_n157_ = new_n156_ & new_n150_;
  assign new_n158_ = ~i_99 ^ ~i_43;
  assign new_n159_ = ~new_n158_;
  assign new_n160_ = ~i_98 ^ ~i_42;
  assign new_n161_ = ~new_n160_;
  assign new_n162_ = new_n161_ & new_n159_;
  assign new_n163_ = ~i_101 ^ ~i_45;
  assign new_n164_ = ~i_100 ^ ~i_44;
  assign new_n165_ = ~new_n164_;
  assign new_n166_ = new_n165_ & new_n163_;
  assign new_n167_ = new_n166_ & new_n162_;
  assign new_n168_ = ~i_103 ^ ~i_47;
  assign new_n169_ = ~i_102 ^ ~i_46;
  assign new_n170_ = new_n169_ & new_n168_;
  assign new_n171_ = ~i_105 ^ ~i_49;
  assign new_n172_ = ~new_n171_;
  assign new_n173_ = ~i_104 ^ ~i_48;
  assign new_n174_ = new_n173_ & new_n172_;
  assign new_n175_ = new_n174_ & new_n170_;
  assign new_n176_ = new_n175_ & new_n167_;
  assign new_n177_ = ~new_n176_;
  assign new_n178_ = new_n173_ & new_n171_;
  assign new_n179_ = new_n178_ & new_n170_;
  assign new_n180_ = new_n179_ & new_n167_;
  assign new_n181_ = new_n164_ & new_n162_;
  assign new_n182_ = new_n161_ & new_n158_;
  assign new_n183_ = ~new_n182_ ^ ~new_n160_;
  assign new_n184_ = ~new_n183_ ^ ~new_n181_;
  assign new_n185_ = ~new_n184_ ^ ~new_n180_;
  assign new_n186_ = ~new_n185_ ^ ~new_n177_;
  assign new_n187_ = ~i_83 ^ ~i_27;
  assign new_n188_ = ~i_91 ^ ~i_35;
  assign new_n189_ = ~i_96 ^ ~i_40;
  assign new_n190_ = ~new_n189_;
  assign new_n191_ = ~i_95 ^ ~i_39;
  assign new_n192_ = new_n191_ & new_n190_;
  assign new_n193_ = ~new_n192_ ^ ~new_n189_;
  assign new_n194_ = ~i_94 ^ ~i_38;
  assign new_n195_ = ~new_n194_;
  assign new_n196_ = new_n195_ & new_n193_;
  assign new_n197_ = ~new_n196_ ^ ~new_n193_;
  assign new_n198_ = ~new_n197_;
  assign new_n199_ = ~i_93 ^ ~i_37;
  assign new_n200_ = new_n199_ & new_n198_;
  assign new_n201_ = ~new_n200_ ^ ~new_n197_;
  assign new_n202_ = ~new_n201_;
  assign new_n203_ = ~i_92 ^ ~i_36;
  assign new_n204_ = new_n203_ & new_n202_;
  assign new_n205_ = ~new_n204_ ^ ~new_n201_;
  assign new_n206_ = ~new_n205_ ^ ~new_n188_;
  assign new_n207_ = ~new_n206_ ^ ~new_n187_;
  assign new_n208_ = ~i_82 ^ ~i_26;
  assign new_n209_ = ~new_n205_;
  assign new_n210_ = new_n209_ & new_n188_;
  assign new_n211_ = ~new_n210_ ^ ~new_n205_;
  assign new_n212_ = ~i_90 ^ ~i_34;
  assign new_n213_ = ~new_n212_ ^ ~new_n211_;
  assign new_n214_ = ~new_n213_ ^ ~new_n208_;
  assign new_n215_ = new_n214_ & new_n207_;
  assign new_n216_ = ~i_84 ^ ~i_28;
  assign new_n217_ = ~new_n203_ ^ ~new_n201_;
  assign new_n218_ = ~new_n217_ ^ ~new_n216_;
  assign new_n219_ = ~i_86 ^ ~i_30;
  assign new_n220_ = ~new_n193_;
  assign new_n221_ = ~new_n194_ ^ ~new_n220_;
  assign new_n222_ = ~new_n221_ ^ ~new_n219_;
  assign new_n223_ = ~i_88 ^ ~i_32;
  assign new_n224_ = ~new_n223_ ^ ~new_n189_;
  assign new_n225_ = ~i_33;
  assign new_n226_ = ~i_89 ^ ~new_n225_;
  assign new_n227_ = ~i_97 ^ ~i_41;
  assign new_n228_ = new_n227_ & new_n226_;
  assign new_n229_ = new_n228_ & new_n224_;
  assign new_n230_ = ~new_n223_;
  assign new_n231_ = new_n230_ & new_n190_;
  assign new_n232_ = ~new_n231_ ^ ~new_n229_;
  assign new_n233_ = ~i_87 ^ ~i_31;
  assign new_n234_ = ~new_n191_ ^ ~new_n189_;
  assign new_n235_ = ~new_n234_ ^ ~new_n233_;
  assign new_n236_ = new_n235_ & new_n232_;
  assign new_n237_ = new_n236_ & new_n222_;
  assign new_n238_ = ~new_n237_;
  assign new_n239_ = ~new_n233_;
  assign new_n240_ = ~new_n234_;
  assign new_n241_ = new_n240_ & new_n239_;
  assign new_n242_ = new_n241_ & new_n222_;
  assign new_n243_ = ~new_n242_;
  assign new_n244_ = ~new_n219_;
  assign new_n245_ = ~new_n221_;
  assign new_n246_ = new_n245_ & new_n244_;
  assign new_n247_ = ~new_n246_ ^ ~new_n243_;
  assign new_n248_ = ~new_n247_ ^ ~new_n238_;
  assign new_n249_ = ~i_85 ^ ~i_29;
  assign new_n250_ = ~new_n199_ ^ ~new_n197_;
  assign new_n251_ = ~new_n250_ ^ ~new_n249_;
  assign new_n252_ = new_n251_ & new_n248_;
  assign new_n253_ = new_n252_ & new_n218_;
  assign new_n254_ = new_n253_ & new_n215_;
  assign new_n255_ = ~new_n249_;
  assign new_n256_ = ~new_n250_;
  assign new_n257_ = new_n256_ & new_n255_;
  assign new_n258_ = new_n257_ & new_n218_;
  assign new_n259_ = ~new_n216_;
  assign new_n260_ = ~new_n217_;
  assign new_n261_ = new_n260_ & new_n259_;
  assign new_n262_ = ~new_n261_ ^ ~new_n258_;
  assign new_n263_ = new_n262_ & new_n215_;
  assign new_n264_ = ~new_n187_;
  assign new_n265_ = ~new_n206_;
  assign new_n266_ = new_n265_ & new_n264_;
  assign new_n267_ = new_n266_ & new_n214_;
  assign new_n268_ = ~new_n208_;
  assign new_n269_ = ~new_n213_;
  assign new_n270_ = new_n269_ & new_n268_;
  assign new_n271_ = ~new_n270_ ^ ~new_n267_;
  assign new_n272_ = ~new_n271_ ^ ~new_n263_;
  assign new_n273_ = ~new_n272_ ^ ~new_n254_;
  assign new_n274_ = ~i_75 ^ ~i_19;
  assign new_n275_ = ~new_n274_;
  assign new_n276_ = ~i_74 ^ ~i_18;
  assign new_n277_ = ~new_n276_;
  assign new_n278_ = new_n277_ & new_n275_;
  assign new_n279_ = ~i_77 ^ ~i_21;
  assign new_n280_ = ~new_n279_;
  assign new_n281_ = ~i_76 ^ ~i_20;
  assign new_n282_ = new_n281_ & new_n280_;
  assign new_n283_ = new_n282_ & new_n278_;
  assign new_n284_ = ~i_79 ^ ~i_23;
  assign new_n285_ = ~new_n284_;
  assign new_n286_ = ~i_78 ^ ~i_22;
  assign new_n287_ = new_n286_ & new_n285_;
  assign new_n288_ = ~i_81 ^ ~i_25;
  assign new_n289_ = ~new_n288_;
  assign new_n290_ = ~i_80 ^ ~i_24;
  assign new_n291_ = ~new_n290_;
  assign new_n292_ = new_n291_ & new_n289_;
  assign new_n293_ = new_n292_ & new_n287_;
  assign new_n294_ = new_n293_ & new_n283_;
  assign new_n295_ = ~new_n294_;
  assign new_n296_ = new_n291_ & new_n288_;
  assign new_n297_ = ~new_n296_ ^ ~new_n290_;
  assign new_n298_ = new_n297_ & new_n287_;
  assign new_n299_ = new_n286_ & new_n284_;
  assign new_n300_ = ~new_n299_ ^ ~new_n298_;
  assign new_n301_ = new_n300_ & new_n283_;
  assign new_n302_ = new_n281_ & new_n279_;
  assign new_n303_ = new_n302_ & new_n278_;
  assign new_n304_ = new_n277_ & new_n274_;
  assign new_n305_ = ~new_n304_ ^ ~new_n276_;
  assign new_n306_ = ~new_n305_ ^ ~new_n303_;
  assign new_n307_ = ~new_n306_ ^ ~new_n301_;
  assign new_n308_ = ~new_n307_ ^ ~new_n295_;
  assign new_n309_ = ~i_61 ^ ~i_5;
  assign new_n310_ = ~i_62 ^ ~i_6;
  assign new_n311_ = ~i_63 ^ ~i_7;
  assign new_n312_ = ~i_64 ^ ~i_8;
  assign new_n313_ = ~i_72 ^ ~i_16;
  assign new_n314_ = ~new_n313_;
  assign new_n315_ = ~i_73 ^ ~i_17;
  assign new_n316_ = new_n315_ & new_n314_;
  assign new_n317_ = ~new_n316_ ^ ~new_n313_;
  assign new_n318_ = ~i_69 ^ ~i_13;
  assign new_n319_ = ~i_68 ^ ~i_12;
  assign new_n320_ = new_n319_ & new_n318_;
  assign new_n321_ = ~i_67 ^ ~i_11;
  assign new_n322_ = ~new_n321_;
  assign new_n323_ = ~i_66 ^ ~i_10;
  assign new_n324_ = ~new_n323_;
  assign new_n325_ = new_n324_ & new_n322_;
  assign new_n326_ = new_n325_ & new_n320_;
  assign new_n327_ = ~i_71 ^ ~i_15;
  assign new_n328_ = ~i_70 ^ ~i_14;
  assign new_n329_ = new_n328_ & new_n327_;
  assign new_n330_ = new_n329_ & new_n326_;
  assign new_n331_ = new_n330_ & new_n317_;
  assign new_n332_ = new_n324_ & new_n321_;
  assign new_n333_ = ~new_n332_ ^ ~new_n323_;
  assign new_n334_ = ~new_n333_ ^ ~new_n331_;
  assign new_n335_ = new_n334_ & new_n151_;
  assign new_n336_ = ~new_n333_;
  assign new_n337_ = ~new_n327_;
  assign new_n338_ = ~new_n328_;
  assign new_n339_ = new_n338_ & new_n337_;
  assign new_n340_ = new_n315_ & new_n313_;
  assign new_n341_ = new_n340_ & new_n339_;
  assign new_n342_ = ~new_n341_;
  assign new_n343_ = new_n338_ & new_n327_;
  assign new_n344_ = ~new_n343_ ^ ~new_n338_;
  assign new_n345_ = ~new_n344_ ^ ~new_n342_;
  assign new_n346_ = new_n345_ & new_n326_;
  assign new_n347_ = ~new_n346_;
  assign new_n348_ = new_n347_ & new_n336_;
  assign new_n349_ = ~new_n348_;
  assign new_n350_ = new_n346_ & new_n333_;
  assign new_n351_ = ~new_n350_;
  assign new_n352_ = new_n351_ & new_n150_;
  assign new_n353_ = new_n352_ & new_n349_;
  assign new_n354_ = ~new_n353_ ^ ~new_n335_;
  assign new_n355_ = ~new_n354_ ^ ~new_n312_;
  assign new_n356_ = ~new_n355_ ^ ~new_n311_;
  assign new_n357_ = ~new_n356_ ^ ~new_n310_;
  assign new_n358_ = ~new_n357_ ^ ~new_n309_;
  assign new_n359_ = ~new_n358_ ^ ~new_n308_;
  assign new_n360_ = ~new_n359_ ^ ~new_n273_;
  assign new_n361_ = ~new_n360_ ^ ~new_n186_;
  assign new_n362_ = ~new_n361_ ^ ~new_n157_;
  assign new_n363_ = new_n362_ & new_n152_;
  assign new_n364_ = new_n361_ & new_n157_;
  assign new_n365_ = ~new_n364_;
  assign new_n366_ = new_n360_ & new_n186_;
  assign new_n367_ = new_n359_ & new_n273_;
  assign new_n368_ = new_n358_ & new_n308_;
  assign new_n369_ = new_n357_ & new_n309_;
  assign new_n370_ = new_n356_ & new_n310_;
  assign new_n371_ = new_n355_ & new_n311_;
  assign new_n372_ = new_n353_ & new_n335_;
  assign new_n373_ = ~new_n372_;
  assign new_n374_ = new_n354_ & new_n312_;
  assign new_n375_ = ~new_n374_ ^ ~new_n373_;
  assign new_n376_ = ~new_n375_ ^ ~new_n371_;
  assign new_n377_ = ~new_n376_ ^ ~new_n370_;
  assign new_n378_ = ~new_n377_ ^ ~new_n369_;
  assign new_n379_ = ~new_n378_ ^ ~new_n368_;
  assign new_n380_ = ~new_n379_ ^ ~new_n367_;
  assign new_n381_ = ~new_n380_ ^ ~new_n366_;
  assign new_n382_ = ~new_n381_ ^ ~new_n365_;
  assign new_n383_ = new_n382_ & new_n363_;
  assign new_n384_ = ~new_n381_;
  assign new_n385_ = new_n384_ & new_n364_;
  assign new_n386_ = ~new_n380_;
  assign new_n387_ = new_n386_ & new_n366_;
  assign new_n388_ = ~new_n379_;
  assign new_n389_ = new_n388_ & new_n367_;
  assign new_n390_ = ~new_n378_;
  assign new_n391_ = new_n390_ & new_n368_;
  assign new_n392_ = ~new_n377_;
  assign new_n393_ = new_n392_ & new_n369_;
  assign new_n394_ = ~new_n376_;
  assign new_n395_ = new_n394_ & new_n370_;
  assign new_n396_ = ~new_n375_;
  assign new_n397_ = new_n396_ & new_n371_;
  assign new_n398_ = ~new_n397_;
  assign new_n399_ = new_n374_ & new_n372_;
  assign new_n400_ = ~new_n399_ ^ ~new_n398_;
  assign new_n401_ = ~new_n400_ ^ ~new_n395_;
  assign new_n402_ = ~new_n401_ ^ ~new_n393_;
  assign new_n403_ = ~new_n402_ ^ ~new_n391_;
  assign new_n404_ = ~new_n403_ ^ ~new_n389_;
  assign new_n405_ = ~new_n404_ ^ ~new_n387_;
  assign new_n406_ = ~new_n405_ ^ ~new_n385_;
  assign new_n407_ = ~new_n406_;
  assign new_n408_ = new_n407_ & new_n383_;
  assign new_n409_ = ~new_n408_;
  assign new_n410_ = ~new_n405_;
  assign new_n411_ = new_n410_ & new_n385_;
  assign new_n412_ = ~new_n404_;
  assign new_n413_ = new_n412_ & new_n387_;
  assign new_n414_ = ~new_n403_;
  assign new_n415_ = new_n414_ & new_n389_;
  assign new_n416_ = ~new_n402_;
  assign new_n417_ = new_n416_ & new_n391_;
  assign new_n418_ = ~new_n401_;
  assign new_n419_ = new_n418_ & new_n393_;
  assign new_n420_ = ~new_n400_;
  assign new_n421_ = new_n420_ & new_n395_;
  assign new_n422_ = ~new_n421_;
  assign new_n423_ = new_n399_ & new_n397_;
  assign new_n424_ = ~new_n423_ ^ ~new_n422_;
  assign new_n425_ = ~new_n424_ ^ ~new_n419_;
  assign new_n426_ = ~new_n425_ ^ ~new_n417_;
  assign new_n427_ = ~new_n426_ ^ ~new_n415_;
  assign new_n428_ = ~new_n427_ ^ ~new_n413_;
  assign new_n429_ = ~new_n428_ ^ ~new_n411_;
  assign m_0 = ~new_n429_ ^ ~new_n409_;
  assign new_n431_ = ~new_n383_;
  assign m_1 = ~new_n406_ ^ ~new_n431_;
  assign m_2 = ~new_n382_ ^ ~new_n363_;
  assign m_3 = ~new_n362_ ^ ~new_n152_;
endmodule


