module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n9 = x0 & ~x1 ;
  assign n10 = x2 & n9 ;
  assign n14 = x1 & x2 ;
  assign n11 = x0 & x1 ;
  assign n12 = n11 ^ x0 ;
  assign n13 = n12 ^ x1 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = x3 & n15 ;
  assign n19 = x3 & x4 ;
  assign n20 = n19 ^ x3 ;
  assign n17 = x2 & x3 ;
  assign n18 = n17 ^ x2 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = ~n15 & n21 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = x4 & ~n23 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = x5 & ~n23 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = x4 & x5 ;
  assign n29 = n28 ^ x4 ;
  assign n30 = x6 & n29 ;
  assign n31 = n30 ^ x6 ;
  assign n32 = ~n23 & n31 ;
  assign n33 = n32 ^ x6 ;
  assign n37 = n29 ^ x5 ;
  assign n38 = x7 & ~n37 ;
  assign n39 = ~n23 & n38 ;
  assign n34 = x5 & x6 ;
  assign n35 = x7 & n34 ;
  assign n36 = ~n23 & n35 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = n40 ^ x7 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = n10 ;
  assign y3 = n16 ;
  assign y4 = n25 ;
  assign y5 = n27 ;
  assign y6 = n33 ;
  assign y7 = n41 ;
endmodule
