module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 ;
  assign n61 = ~x9 & ~x10 ;
  assign n62 = x11 & ~n61 ;
  assign n63 = ~x12 & ~x13 ;
  assign n64 = x14 & x15 ;
  assign n65 = n63 & n64 ;
  assign n66 = ~n62 & n65 ;
  assign n67 = n66 ^ n64 ;
  assign n68 = x16 & n67 ;
  assign n69 = ~x7 & ~x8 ;
  assign n70 = x9 & ~x10 ;
  assign n71 = n69 & n70 ;
  assign n72 = ~x3 & ~x4 ;
  assign n73 = ~x5 & ~x6 ;
  assign n74 = n72 & n73 ;
  assign n75 = n71 & n74 ;
  assign n76 = x24 & x25 ;
  assign n77 = ~x26 & n76 ;
  assign n78 = ~x13 & x14 ;
  assign n79 = ~x18 & x19 ;
  assign n80 = n78 & n79 ;
  assign n81 = n77 & n80 ;
  assign n82 = n75 & n81 ;
  assign n83 = x20 & ~x21 ;
  assign n84 = ~x22 & x23 ;
  assign n85 = ~x1 & ~x2 ;
  assign n86 = n84 & n85 ;
  assign n87 = n83 & n86 ;
  assign n92 = ~x11 & x12 ;
  assign n93 = n61 & n92 ;
  assign n94 = n87 & n93 ;
  assign n95 = n82 & n94 ;
  assign n88 = x11 & ~x12 ;
  assign n89 = ~n61 & n88 ;
  assign n90 = n87 & n89 ;
  assign n91 = n82 & n90 ;
  assign n96 = n95 ^ n91 ;
  assign n97 = ~n68 & n96 ;
  assign n111 = x27 & x28 ;
  assign n112 = x29 & n111 ;
  assign n113 = ~x26 & n112 ;
  assign n107 = x23 & x24 ;
  assign n116 = x25 & n107 ;
  assign n117 = n113 & ~n116 ;
  assign n102 = ~x16 & x17 ;
  assign n98 = x19 & x20 ;
  assign n103 = ~x18 & n98 ;
  assign n104 = n102 & n103 ;
  assign n105 = ~n67 & n104 ;
  assign n99 = ~x17 & ~x18 ;
  assign n100 = n98 & n99 ;
  assign n101 = n100 ^ n98 ;
  assign n106 = n105 ^ n101 ;
  assign n108 = ~x21 & ~x22 ;
  assign n109 = x25 & n108 ;
  assign n110 = n107 & n109 ;
  assign n114 = n110 & n113 ;
  assign n115 = ~n106 & n114 ;
  assign n118 = n117 ^ n115 ;
  assign n119 = n118 ^ n112 ;
  assign n120 = ~n67 & n102 ;
  assign n121 = n120 ^ x17 ;
  assign n122 = x14 & n63 ;
  assign n123 = ~n62 & n122 ;
  assign n124 = n123 ^ x14 ;
  assign n125 = n124 ^ x15 ;
  assign n126 = n121 & ~n125 ;
  assign n127 = n119 & n126 ;
  assign n128 = n97 & n127 ;
  assign n129 = n128 ^ n119 ;
  assign n130 = x19 & x25 ;
  assign n131 = ~x26 & n130 ;
  assign n132 = x15 & ~x16 ;
  assign n133 = n63 & n132 ;
  assign n134 = n131 & n133 ;
  assign n135 = n112 & n134 ;
  assign n136 = n83 & n84 ;
  assign n137 = x0 & x1 ;
  assign n138 = n61 & n137 ;
  assign n139 = n136 & n138 ;
  assign n140 = x6 & x7 ;
  assign n141 = x8 & x11 ;
  assign n142 = n140 & n141 ;
  assign n143 = x2 & x3 ;
  assign n144 = x4 & x5 ;
  assign n145 = n143 & n144 ;
  assign n146 = n142 & n145 ;
  assign n147 = n139 & n146 ;
  assign n148 = n135 & n147 ;
  assign n150 = ~n62 & n63 ;
  assign n151 = n150 ^ x14 ;
  assign n155 = n148 & ~n151 ;
  assign n149 = ~x16 & ~n67 ;
  assign n152 = ~x17 & ~n151 ;
  assign n153 = n149 & n152 ;
  assign n154 = n148 & n153 ;
  assign n156 = n155 ^ n154 ;
  assign n157 = ~x18 & n102 ;
  assign n158 = ~n67 & n157 ;
  assign n159 = n158 ^ n99 ;
  assign n166 = ~x24 & n159 ;
  assign n167 = ~n119 & n166 ;
  assign n168 = n156 & n167 ;
  assign n160 = x23 & n108 ;
  assign n161 = ~n106 & n160 ;
  assign n162 = n161 ^ x23 ;
  assign n163 = n159 & ~n162 ;
  assign n164 = ~n119 & n163 ;
  assign n165 = n156 & n164 ;
  assign n169 = n168 ^ n165 ;
  assign n170 = n169 ^ n119 ;
  assign n171 = ~n129 & n170 ;
  assign n172 = x36 & x37 ;
  assign n173 = x38 & x41 ;
  assign n174 = n172 & n173 ;
  assign n175 = x32 & x33 ;
  assign n176 = x34 & x35 ;
  assign n177 = n175 & n176 ;
  assign n178 = n174 & n177 ;
  assign n179 = x57 & x58 ;
  assign n180 = x59 & n179 ;
  assign n181 = ~x46 & x47 ;
  assign n182 = x50 & ~x56 ;
  assign n183 = n181 & n182 ;
  assign n184 = n180 & n183 ;
  assign n185 = n178 & n184 ;
  assign n186 = ~x39 & ~x40 ;
  assign n188 = ~x41 & ~x42 ;
  assign n189 = ~n186 & n188 ;
  assign n187 = ~x42 & n186 ;
  assign n190 = n189 ^ n187 ;
  assign n191 = ~x43 & x44 ;
  assign n192 = n190 & n191 ;
  assign n193 = n192 ^ x44 ;
  assign n194 = x54 & x55 ;
  assign n195 = x30 & x31 ;
  assign n196 = n194 & n195 ;
  assign n197 = ~x48 & ~x49 ;
  assign n198 = n186 & ~n197 ;
  assign n199 = n196 & n198 ;
  assign n200 = ~n193 & n199 ;
  assign n201 = n185 & n200 ;
  assign n205 = x44 & x45 ;
  assign n206 = ~x46 & n205 ;
  assign n202 = x45 & ~x46 ;
  assign n203 = n191 & n202 ;
  assign n204 = n190 & n203 ;
  assign n207 = n206 ^ n204 ;
  assign n208 = n207 ^ x46 ;
  assign n212 = x47 & x49 ;
  assign n213 = n208 & n212 ;
  assign n209 = x47 & x48 ;
  assign n210 = n208 & n209 ;
  assign n211 = n210 ^ x48 ;
  assign n214 = n213 ^ n211 ;
  assign n223 = n193 ^ x45 ;
  assign n224 = ~n214 & ~n223 ;
  assign n225 = n201 & n224 ;
  assign n215 = x41 & x42 ;
  assign n216 = ~n186 & n215 ;
  assign n217 = ~x44 & x45 ;
  assign n218 = x43 & n217 ;
  assign n219 = n216 & n218 ;
  assign n220 = n219 ^ n217 ;
  assign n221 = ~n214 & ~n220 ;
  assign n222 = n201 & n221 ;
  assign n226 = n225 ^ n222 ;
  assign n236 = x47 & ~x48 ;
  assign n231 = ~x51 & ~x52 ;
  assign n232 = x49 & x50 ;
  assign n237 = n231 & n232 ;
  assign n238 = n236 & n237 ;
  assign n239 = n208 & n238 ;
  assign n233 = x48 & n232 ;
  assign n234 = n231 & n233 ;
  assign n235 = n234 ^ n231 ;
  assign n240 = n239 ^ n235 ;
  assign n241 = x53 & n194 ;
  assign n242 = n180 & n241 ;
  assign n227 = ~x0 & ~x51 ;
  assign n243 = ~x56 & ~n227 ;
  assign n244 = n242 & n243 ;
  assign n245 = ~n240 & n244 ;
  assign n228 = x56 & ~n227 ;
  assign n229 = n180 & n228 ;
  assign n230 = n229 ^ n227 ;
  assign n246 = n245 ^ n230 ;
  assign n247 = n232 & n236 ;
  assign n248 = n208 & n247 ;
  assign n249 = n248 ^ n233 ;
  assign n254 = ~x52 & x53 ;
  assign n255 = ~n249 & n254 ;
  assign n256 = n246 & n255 ;
  assign n257 = n226 & n256 ;
  assign n250 = x52 & ~x53 ;
  assign n251 = n249 & n250 ;
  assign n252 = n246 & n251 ;
  assign n253 = n226 & n252 ;
  assign n258 = n257 ^ n253 ;
  assign n259 = n232 & n254 ;
  assign n260 = ~n209 & n259 ;
  assign n261 = ~x33 & ~x34 ;
  assign n262 = ~x35 & ~x36 ;
  assign n263 = n261 & n262 ;
  assign n264 = ~x31 & ~x32 ;
  assign n265 = n194 & n264 ;
  assign n266 = n263 & n265 ;
  assign n267 = n260 & n266 ;
  assign n268 = x41 & ~x43 ;
  assign n269 = n205 & n268 ;
  assign n270 = ~x37 & ~x38 ;
  assign n271 = x39 & ~x40 ;
  assign n272 = n270 & n271 ;
  assign n273 = n269 & n272 ;
  assign n274 = ~x56 & x57 ;
  assign n275 = ~x46 & ~x51 ;
  assign n276 = n274 & n275 ;
  assign n277 = x41 & ~n186 ;
  assign n278 = n277 ^ x42 ;
  assign n279 = n276 & n278 ;
  assign n280 = n273 & n279 ;
  assign n281 = n267 & n280 ;
  assign n282 = x47 & n208 ;
  assign n298 = x48 & ~n208 ;
  assign n299 = ~n282 & ~n298 ;
  assign n300 = n281 & ~n299 ;
  assign n283 = ~x0 & ~x30 ;
  assign n293 = ~x56 & n180 ;
  assign n294 = n241 & n293 ;
  assign n295 = ~n240 & n294 ;
  assign n292 = x56 & n180 ;
  assign n296 = n295 ^ n292 ;
  assign n301 = n283 & ~n296 ;
  assign n302 = n300 & n301 ;
  assign n303 = ~n258 & n302 ;
  assign n297 = ~n258 & ~n296 ;
  assign n304 = n303 ^ n297 ;
  assign n286 = x48 & n283 ;
  assign n287 = ~n208 & n286 ;
  assign n288 = ~n282 & n287 ;
  assign n289 = n281 & n288 ;
  assign n284 = n282 & n283 ;
  assign n285 = n281 & n284 ;
  assign n290 = n289 ^ n285 ;
  assign n291 = ~n258 & n290 ;
  assign n305 = n304 ^ n291 ;
  assign n321 = ~n119 & ~n305 ;
  assign n313 = n156 & n159 ;
  assign n317 = x24 & ~n119 ;
  assign n315 = x23 & ~n119 ;
  assign n314 = ~n119 & n161 ;
  assign n316 = n315 ^ n314 ;
  assign n318 = n317 ^ n316 ;
  assign n319 = n313 & n318 ;
  assign n320 = ~n305 & n319 ;
  assign n322 = n321 ^ n320 ;
  assign n323 = n322 ^ n305 ;
  assign n307 = ~n68 & ~n125 ;
  assign n308 = n96 & n307 ;
  assign n309 = n119 & n121 ;
  assign n310 = n308 & n309 ;
  assign n311 = n305 & n310 ;
  assign n306 = n119 & n305 ;
  assign n312 = n311 ^ n306 ;
  assign n324 = n323 ^ n312 ;
  assign n325 = x0 & x30 ;
  assign n328 = x48 & ~n325 ;
  assign n329 = ~n208 & n328 ;
  assign n330 = ~n282 & n329 ;
  assign n331 = n281 & n330 ;
  assign n326 = n282 & ~n325 ;
  assign n327 = n281 & n326 ;
  assign n332 = n331 ^ n327 ;
  assign n333 = n296 & ~n332 ;
  assign n334 = ~n129 & n333 ;
  assign n335 = n170 & n334 ;
  assign y0 = ~n171 ;
  assign y1 = n324 ;
  assign y2 = n335 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
