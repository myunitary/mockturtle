module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 ;
  assign n165 = x0 & ~x40 ;
  assign n130 = x40 ^ x0 ;
  assign n163 = x1 & ~x41 ;
  assign n164 = ~n130 & n163 ;
  assign n166 = n165 ^ n164 ;
  assign n131 = x41 ^ x1 ;
  assign n132 = ~n130 & ~n131 ;
  assign n160 = x2 & ~x42 ;
  assign n133 = x42 ^ x2 ;
  assign n158 = x3 & ~x43 ;
  assign n159 = ~n133 & n158 ;
  assign n161 = n160 ^ n159 ;
  assign n162 = n132 & n161 ;
  assign n167 = n166 ^ n162 ;
  assign n134 = x43 ^ x3 ;
  assign n135 = ~n133 & ~n134 ;
  assign n136 = n132 & n135 ;
  assign n154 = x4 & ~x44 ;
  assign n137 = x44 ^ x4 ;
  assign n152 = x5 & ~x45 ;
  assign n153 = ~n137 & n152 ;
  assign n155 = n154 ^ n153 ;
  assign n138 = x45 ^ x5 ;
  assign n139 = ~n137 & ~n138 ;
  assign n149 = x6 & ~x46 ;
  assign n140 = x46 ^ x6 ;
  assign n145 = x7 & x47 ;
  assign n146 = n145 ^ x7 ;
  assign n147 = n140 & n146 ;
  assign n148 = n147 ^ n146 ;
  assign n150 = n149 ^ n148 ;
  assign n151 = n139 & n150 ;
  assign n156 = n155 ^ n151 ;
  assign n157 = n136 & n156 ;
  assign n168 = n167 ^ n157 ;
  assign n141 = x47 ^ x7 ;
  assign n142 = ~n140 & ~n141 ;
  assign n143 = n139 & n142 ;
  assign n144 = n136 & n143 ;
  assign n169 = n168 ^ n144 ;
  assign n587 = x0 & ~x24 ;
  assign n552 = x24 ^ x0 ;
  assign n585 = x1 & ~x25 ;
  assign n586 = ~n552 & n585 ;
  assign n588 = n587 ^ n586 ;
  assign n553 = x25 ^ x1 ;
  assign n554 = ~n552 & ~n553 ;
  assign n582 = x2 & ~x26 ;
  assign n555 = x26 ^ x2 ;
  assign n580 = x3 & ~x27 ;
  assign n581 = ~n555 & n580 ;
  assign n583 = n582 ^ n581 ;
  assign n584 = n554 & n583 ;
  assign n589 = n588 ^ n584 ;
  assign n556 = x27 ^ x3 ;
  assign n557 = ~n555 & ~n556 ;
  assign n558 = n554 & n557 ;
  assign n576 = x4 & ~x28 ;
  assign n559 = x28 ^ x4 ;
  assign n574 = x5 & ~x29 ;
  assign n575 = ~n559 & n574 ;
  assign n577 = n576 ^ n575 ;
  assign n560 = x29 ^ x5 ;
  assign n561 = ~n559 & ~n560 ;
  assign n571 = x6 & ~x30 ;
  assign n562 = x30 ^ x6 ;
  assign n567 = x7 & x31 ;
  assign n568 = n567 ^ x7 ;
  assign n569 = n562 & n568 ;
  assign n570 = n569 ^ n568 ;
  assign n572 = n571 ^ n570 ;
  assign n573 = n561 & n572 ;
  assign n578 = n577 ^ n573 ;
  assign n579 = n558 & n578 ;
  assign n590 = n589 ^ n579 ;
  assign n563 = x31 ^ x7 ;
  assign n564 = ~n562 & ~n563 ;
  assign n565 = n561 & n564 ;
  assign n566 = n558 & n565 ;
  assign n591 = n590 ^ n566 ;
  assign n804 = ~n169 & n591 ;
  assign n395 = x0 & ~x32 ;
  assign n360 = x32 ^ x0 ;
  assign n393 = x1 & ~x33 ;
  assign n394 = ~n360 & n393 ;
  assign n396 = n395 ^ n394 ;
  assign n361 = x33 ^ x1 ;
  assign n362 = ~n360 & ~n361 ;
  assign n390 = x2 & ~x34 ;
  assign n363 = x34 ^ x2 ;
  assign n388 = x3 & ~x35 ;
  assign n389 = ~n363 & n388 ;
  assign n391 = n390 ^ n389 ;
  assign n392 = n362 & n391 ;
  assign n397 = n396 ^ n392 ;
  assign n364 = x35 ^ x3 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = n362 & n365 ;
  assign n384 = x4 & ~x36 ;
  assign n367 = x36 ^ x4 ;
  assign n382 = x5 & ~x37 ;
  assign n383 = ~n367 & n382 ;
  assign n385 = n384 ^ n383 ;
  assign n368 = x37 ^ x5 ;
  assign n369 = ~n367 & ~n368 ;
  assign n379 = x6 & ~x38 ;
  assign n370 = x38 ^ x6 ;
  assign n375 = x7 & x39 ;
  assign n376 = n375 ^ x7 ;
  assign n377 = n370 & n376 ;
  assign n378 = n377 ^ n376 ;
  assign n380 = n379 ^ n378 ;
  assign n381 = n369 & n380 ;
  assign n386 = n385 ^ n381 ;
  assign n387 = n366 & n386 ;
  assign n398 = n397 ^ n387 ;
  assign n371 = x39 ^ x7 ;
  assign n372 = ~n370 & ~n371 ;
  assign n373 = n369 & n372 ;
  assign n374 = n366 & n373 ;
  assign n399 = n398 ^ n374 ;
  assign n803 = ~n399 & n591 ;
  assign n805 = n804 ^ n803 ;
  assign n793 = n399 ^ n169 ;
  assign n798 = n591 & n793 ;
  assign n806 = n805 ^ n798 ;
  assign n760 = x0 & ~x8 ;
  assign n725 = x8 ^ x0 ;
  assign n758 = x1 & ~x9 ;
  assign n759 = ~n725 & n758 ;
  assign n761 = n760 ^ n759 ;
  assign n726 = x9 ^ x1 ;
  assign n727 = ~n725 & ~n726 ;
  assign n755 = x2 & ~x10 ;
  assign n728 = x10 ^ x2 ;
  assign n753 = x3 & ~x11 ;
  assign n754 = ~n728 & n753 ;
  assign n756 = n755 ^ n754 ;
  assign n757 = n727 & n756 ;
  assign n762 = n761 ^ n757 ;
  assign n729 = x11 ^ x3 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = n727 & n730 ;
  assign n749 = x4 & ~x12 ;
  assign n732 = x12 ^ x4 ;
  assign n747 = x5 & ~x13 ;
  assign n748 = ~n732 & n747 ;
  assign n750 = n749 ^ n748 ;
  assign n733 = x13 ^ x5 ;
  assign n734 = ~n732 & ~n733 ;
  assign n744 = x6 & ~x14 ;
  assign n735 = x14 ^ x6 ;
  assign n740 = x7 & x15 ;
  assign n741 = n740 ^ x7 ;
  assign n742 = n735 & n741 ;
  assign n743 = n742 ^ n741 ;
  assign n745 = n744 ^ n743 ;
  assign n746 = n734 & n745 ;
  assign n751 = n750 ^ n746 ;
  assign n752 = n731 & n751 ;
  assign n763 = n762 ^ n752 ;
  assign n736 = x15 ^ x7 ;
  assign n737 = ~n735 & ~n736 ;
  assign n738 = n734 & n737 ;
  assign n739 = n731 & n738 ;
  assign n764 = n763 ^ n739 ;
  assign n653 = x0 & ~x16 ;
  assign n618 = x16 ^ x0 ;
  assign n651 = x1 & ~x17 ;
  assign n652 = ~n618 & n651 ;
  assign n654 = n653 ^ n652 ;
  assign n619 = x17 ^ x1 ;
  assign n620 = ~n618 & ~n619 ;
  assign n648 = x2 & ~x18 ;
  assign n621 = x18 ^ x2 ;
  assign n646 = x3 & ~x19 ;
  assign n647 = ~n621 & n646 ;
  assign n649 = n648 ^ n647 ;
  assign n650 = n620 & n649 ;
  assign n655 = n654 ^ n650 ;
  assign n622 = x19 ^ x3 ;
  assign n623 = ~n621 & ~n622 ;
  assign n624 = n620 & n623 ;
  assign n642 = x4 & ~x20 ;
  assign n625 = x20 ^ x4 ;
  assign n640 = x5 & ~x21 ;
  assign n641 = ~n625 & n640 ;
  assign n643 = n642 ^ n641 ;
  assign n626 = x21 ^ x5 ;
  assign n627 = ~n625 & ~n626 ;
  assign n637 = x6 & ~x22 ;
  assign n628 = x22 ^ x6 ;
  assign n633 = x7 & x23 ;
  assign n634 = n633 ^ x7 ;
  assign n635 = n628 & n634 ;
  assign n636 = n635 ^ n634 ;
  assign n638 = n637 ^ n636 ;
  assign n639 = n627 & n638 ;
  assign n644 = n643 ^ n639 ;
  assign n645 = n624 & n644 ;
  assign n656 = n655 ^ n645 ;
  assign n629 = x23 ^ x7 ;
  assign n630 = ~n628 & ~n629 ;
  assign n631 = n627 & n630 ;
  assign n632 = n624 & n631 ;
  assign n657 = n656 ^ n632 ;
  assign n792 = n764 ^ n657 ;
  assign n794 = n793 ^ n591 ;
  assign n795 = n792 & n794 ;
  assign n791 = n657 & n764 ;
  assign n796 = n795 ^ n791 ;
  assign n797 = n169 & n399 ;
  assign n799 = n798 ^ n797 ;
  assign n800 = n799 ^ n795 ;
  assign n801 = n796 & n800 ;
  assign n802 = n801 ^ n795 ;
  assign n807 = n806 ^ n802 ;
  assign n808 = n799 ^ n796 ;
  assign n809 = n794 ^ n792 ;
  assign n810 = x0 & n809 ;
  assign n811 = n810 ^ x0 ;
  assign n812 = n808 & n811 ;
  assign n813 = n812 ^ n811 ;
  assign n814 = n807 & n813 ;
  assign n815 = n814 ^ n813 ;
  assign n124 = x8 & ~x40 ;
  assign n89 = x40 ^ x8 ;
  assign n122 = x9 & ~x41 ;
  assign n123 = ~n89 & n122 ;
  assign n125 = n124 ^ n123 ;
  assign n90 = x41 ^ x9 ;
  assign n91 = ~n89 & ~n90 ;
  assign n119 = x10 & ~x42 ;
  assign n92 = x42 ^ x10 ;
  assign n117 = x11 & ~x43 ;
  assign n118 = ~n92 & n117 ;
  assign n120 = n119 ^ n118 ;
  assign n121 = n91 & n120 ;
  assign n126 = n125 ^ n121 ;
  assign n93 = x43 ^ x11 ;
  assign n94 = ~n92 & ~n93 ;
  assign n95 = n91 & n94 ;
  assign n113 = x12 & ~x44 ;
  assign n96 = x44 ^ x12 ;
  assign n111 = x13 & ~x45 ;
  assign n112 = ~n96 & n111 ;
  assign n114 = n113 ^ n112 ;
  assign n97 = x45 ^ x13 ;
  assign n98 = ~n96 & ~n97 ;
  assign n108 = x14 & ~x46 ;
  assign n99 = x46 ^ x14 ;
  assign n104 = x15 & x47 ;
  assign n105 = n104 ^ x15 ;
  assign n106 = n99 & n105 ;
  assign n107 = n106 ^ n105 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = n98 & n109 ;
  assign n115 = n114 ^ n110 ;
  assign n116 = n95 & n115 ;
  assign n127 = n126 ^ n116 ;
  assign n100 = x47 ^ x15 ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = n98 & n101 ;
  assign n103 = n95 & n102 ;
  assign n128 = n127 ^ n103 ;
  assign n546 = x8 & ~x24 ;
  assign n511 = x24 ^ x8 ;
  assign n544 = x9 & ~x25 ;
  assign n545 = ~n511 & n544 ;
  assign n547 = n546 ^ n545 ;
  assign n512 = x25 ^ x9 ;
  assign n513 = ~n511 & ~n512 ;
  assign n541 = x10 & ~x26 ;
  assign n514 = x26 ^ x10 ;
  assign n539 = x11 & ~x27 ;
  assign n540 = ~n514 & n539 ;
  assign n542 = n541 ^ n540 ;
  assign n543 = n513 & n542 ;
  assign n548 = n547 ^ n543 ;
  assign n515 = x27 ^ x11 ;
  assign n516 = ~n514 & ~n515 ;
  assign n517 = n513 & n516 ;
  assign n535 = x12 & ~x28 ;
  assign n518 = x28 ^ x12 ;
  assign n533 = x13 & ~x29 ;
  assign n534 = ~n518 & n533 ;
  assign n536 = n535 ^ n534 ;
  assign n519 = x29 ^ x13 ;
  assign n520 = ~n518 & ~n519 ;
  assign n530 = x14 & ~x30 ;
  assign n521 = x30 ^ x14 ;
  assign n526 = x15 & x31 ;
  assign n527 = n526 ^ x15 ;
  assign n528 = n521 & n527 ;
  assign n529 = n528 ^ n527 ;
  assign n531 = n530 ^ n529 ;
  assign n532 = n520 & n531 ;
  assign n537 = n536 ^ n532 ;
  assign n538 = n517 & n537 ;
  assign n549 = n548 ^ n538 ;
  assign n522 = x31 ^ x15 ;
  assign n523 = ~n521 & ~n522 ;
  assign n524 = n520 & n523 ;
  assign n525 = n517 & n524 ;
  assign n550 = n549 ^ n525 ;
  assign n780 = ~n128 & n550 ;
  assign n354 = x8 & ~x32 ;
  assign n319 = x32 ^ x8 ;
  assign n352 = x9 & ~x33 ;
  assign n353 = ~n319 & n352 ;
  assign n355 = n354 ^ n353 ;
  assign n320 = x33 ^ x9 ;
  assign n321 = ~n319 & ~n320 ;
  assign n349 = x10 & ~x34 ;
  assign n322 = x34 ^ x10 ;
  assign n347 = x11 & ~x35 ;
  assign n348 = ~n322 & n347 ;
  assign n350 = n349 ^ n348 ;
  assign n351 = n321 & n350 ;
  assign n356 = n355 ^ n351 ;
  assign n323 = x35 ^ x11 ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = n321 & n324 ;
  assign n343 = x12 & ~x36 ;
  assign n326 = x36 ^ x12 ;
  assign n341 = x13 & ~x37 ;
  assign n342 = ~n326 & n341 ;
  assign n344 = n343 ^ n342 ;
  assign n327 = x37 ^ x13 ;
  assign n328 = ~n326 & ~n327 ;
  assign n338 = x14 & ~x38 ;
  assign n329 = x38 ^ x14 ;
  assign n334 = x15 & x39 ;
  assign n335 = n334 ^ x15 ;
  assign n336 = n329 & n335 ;
  assign n337 = n336 ^ n335 ;
  assign n339 = n338 ^ n337 ;
  assign n340 = n328 & n339 ;
  assign n345 = n344 ^ n340 ;
  assign n346 = n325 & n345 ;
  assign n357 = n356 ^ n346 ;
  assign n330 = x39 ^ x15 ;
  assign n331 = ~n329 & ~n330 ;
  assign n332 = n328 & n331 ;
  assign n333 = n325 & n332 ;
  assign n358 = n357 ^ n333 ;
  assign n779 = ~n358 & n550 ;
  assign n781 = n780 ^ n779 ;
  assign n768 = n358 ^ n128 ;
  assign n774 = n550 & n768 ;
  assign n782 = n781 ^ n774 ;
  assign n693 = x8 & ~x16 ;
  assign n658 = x16 ^ x8 ;
  assign n691 = x9 & ~x17 ;
  assign n692 = ~n658 & n691 ;
  assign n694 = n693 ^ n692 ;
  assign n659 = x17 ^ x9 ;
  assign n660 = ~n658 & ~n659 ;
  assign n688 = x10 & ~x18 ;
  assign n661 = x18 ^ x10 ;
  assign n686 = x11 & ~x19 ;
  assign n687 = ~n661 & n686 ;
  assign n689 = n688 ^ n687 ;
  assign n690 = n660 & n689 ;
  assign n695 = n694 ^ n690 ;
  assign n662 = x19 ^ x11 ;
  assign n663 = ~n661 & ~n662 ;
  assign n664 = n660 & n663 ;
  assign n682 = x12 & ~x20 ;
  assign n665 = x20 ^ x12 ;
  assign n680 = x13 & ~x21 ;
  assign n681 = ~n665 & n680 ;
  assign n683 = n682 ^ n681 ;
  assign n666 = x21 ^ x13 ;
  assign n667 = ~n665 & ~n666 ;
  assign n677 = x14 & ~x22 ;
  assign n668 = x22 ^ x14 ;
  assign n673 = x15 & x23 ;
  assign n674 = n673 ^ x15 ;
  assign n675 = n668 & n674 ;
  assign n676 = n675 ^ n674 ;
  assign n678 = n677 ^ n676 ;
  assign n679 = n667 & n678 ;
  assign n684 = n683 ^ n679 ;
  assign n685 = n664 & n684 ;
  assign n696 = n695 ^ n685 ;
  assign n669 = x23 ^ x15 ;
  assign n670 = ~n668 & ~n669 ;
  assign n671 = n667 & n670 ;
  assign n672 = n664 & n671 ;
  assign n697 = n696 ^ n672 ;
  assign n767 = n764 ^ n697 ;
  assign n769 = n768 ^ n550 ;
  assign n770 = n767 & n769 ;
  assign n771 = n770 ^ n769 ;
  assign n765 = n697 & n764 ;
  assign n766 = n765 ^ n697 ;
  assign n772 = n771 ^ n766 ;
  assign n773 = n128 & n358 ;
  assign n775 = n774 ^ n773 ;
  assign n776 = n775 ^ n771 ;
  assign n777 = n772 & n776 ;
  assign n778 = n777 ^ n771 ;
  assign n783 = n782 ^ n778 ;
  assign n784 = n775 ^ n772 ;
  assign n785 = n769 ^ n767 ;
  assign n786 = x8 & n785 ;
  assign n787 = n784 & n786 ;
  assign n788 = n787 ^ n786 ;
  assign n789 = n783 & n788 ;
  assign n790 = n789 ^ n788 ;
  assign n816 = n815 ^ n790 ;
  assign n84 = x16 & ~x40 ;
  assign n49 = x40 ^ x16 ;
  assign n82 = x17 & ~x41 ;
  assign n83 = ~n49 & n82 ;
  assign n85 = n84 ^ n83 ;
  assign n50 = x41 ^ x17 ;
  assign n51 = ~n49 & ~n50 ;
  assign n79 = x18 & ~x42 ;
  assign n52 = x42 ^ x18 ;
  assign n77 = x19 & ~x43 ;
  assign n78 = ~n52 & n77 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n51 & n80 ;
  assign n86 = n85 ^ n81 ;
  assign n53 = x43 ^ x19 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n51 & n54 ;
  assign n73 = x20 & ~x44 ;
  assign n56 = x44 ^ x20 ;
  assign n71 = x21 & ~x45 ;
  assign n72 = ~n56 & n71 ;
  assign n74 = n73 ^ n72 ;
  assign n57 = x45 ^ x21 ;
  assign n58 = ~n56 & ~n57 ;
  assign n68 = x22 & ~x46 ;
  assign n59 = x46 ^ x22 ;
  assign n64 = x23 & x47 ;
  assign n65 = n64 ^ x23 ;
  assign n66 = n59 & n65 ;
  assign n67 = n66 ^ n65 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n58 & n69 ;
  assign n75 = n74 ^ n70 ;
  assign n76 = n55 & n75 ;
  assign n87 = n86 ^ n76 ;
  assign n60 = x47 ^ x23 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = n58 & n61 ;
  assign n63 = n55 & n62 ;
  assign n88 = n87 ^ n63 ;
  assign n506 = x16 & ~x24 ;
  assign n471 = x24 ^ x16 ;
  assign n504 = x17 & ~x25 ;
  assign n505 = ~n471 & n504 ;
  assign n507 = n506 ^ n505 ;
  assign n472 = x25 ^ x17 ;
  assign n473 = ~n471 & ~n472 ;
  assign n501 = x18 & ~x26 ;
  assign n474 = x26 ^ x18 ;
  assign n499 = x19 & ~x27 ;
  assign n500 = ~n474 & n499 ;
  assign n502 = n501 ^ n500 ;
  assign n503 = n473 & n502 ;
  assign n508 = n507 ^ n503 ;
  assign n475 = x27 ^ x19 ;
  assign n476 = ~n474 & ~n475 ;
  assign n477 = n473 & n476 ;
  assign n495 = x20 & ~x28 ;
  assign n478 = x28 ^ x20 ;
  assign n493 = x21 & ~x29 ;
  assign n494 = ~n478 & n493 ;
  assign n496 = n495 ^ n494 ;
  assign n479 = x29 ^ x21 ;
  assign n480 = ~n478 & ~n479 ;
  assign n490 = x22 & ~x30 ;
  assign n481 = x30 ^ x22 ;
  assign n486 = x23 & x31 ;
  assign n487 = n486 ^ x23 ;
  assign n488 = n481 & n487 ;
  assign n489 = n488 ^ n487 ;
  assign n491 = n490 ^ n489 ;
  assign n492 = n480 & n491 ;
  assign n497 = n496 ^ n492 ;
  assign n498 = n477 & n497 ;
  assign n509 = n508 ^ n498 ;
  assign n482 = x31 ^ x23 ;
  assign n483 = ~n481 & ~n482 ;
  assign n484 = n480 & n483 ;
  assign n485 = n477 & n484 ;
  assign n510 = n509 ^ n485 ;
  assign n713 = ~n88 & n510 ;
  assign n314 = x16 & ~x32 ;
  assign n279 = x32 ^ x16 ;
  assign n312 = x17 & ~x33 ;
  assign n313 = ~n279 & n312 ;
  assign n315 = n314 ^ n313 ;
  assign n280 = x33 ^ x17 ;
  assign n281 = ~n279 & ~n280 ;
  assign n309 = x18 & ~x34 ;
  assign n282 = x34 ^ x18 ;
  assign n307 = x19 & ~x35 ;
  assign n308 = ~n282 & n307 ;
  assign n310 = n309 ^ n308 ;
  assign n311 = n281 & n310 ;
  assign n316 = n315 ^ n311 ;
  assign n283 = x35 ^ x19 ;
  assign n284 = ~n282 & ~n283 ;
  assign n285 = n281 & n284 ;
  assign n303 = x20 & ~x36 ;
  assign n286 = x36 ^ x20 ;
  assign n301 = x21 & ~x37 ;
  assign n302 = ~n286 & n301 ;
  assign n304 = n303 ^ n302 ;
  assign n287 = x37 ^ x21 ;
  assign n288 = ~n286 & ~n287 ;
  assign n298 = x22 & ~x38 ;
  assign n289 = x38 ^ x22 ;
  assign n294 = x23 & x39 ;
  assign n295 = n294 ^ x23 ;
  assign n296 = n289 & n295 ;
  assign n297 = n296 ^ n295 ;
  assign n299 = n298 ^ n297 ;
  assign n300 = n288 & n299 ;
  assign n305 = n304 ^ n300 ;
  assign n306 = n285 & n305 ;
  assign n317 = n316 ^ n306 ;
  assign n290 = x39 ^ x23 ;
  assign n291 = ~n289 & ~n290 ;
  assign n292 = n288 & n291 ;
  assign n293 = n285 & n292 ;
  assign n318 = n317 ^ n293 ;
  assign n712 = ~n318 & n510 ;
  assign n714 = n713 ^ n712 ;
  assign n702 = n318 ^ n88 ;
  assign n707 = n510 & n702 ;
  assign n715 = n714 ^ n707 ;
  assign n701 = n697 ^ n657 ;
  assign n703 = n702 ^ n510 ;
  assign n704 = n701 & n703 ;
  assign n698 = n657 & n697 ;
  assign n699 = n698 ^ n657 ;
  assign n700 = n699 ^ n697 ;
  assign n705 = n704 ^ n700 ;
  assign n706 = n88 & n318 ;
  assign n708 = n707 ^ n706 ;
  assign n709 = n708 ^ n704 ;
  assign n710 = ~n705 & n709 ;
  assign n711 = n710 ^ n704 ;
  assign n716 = n715 ^ n711 ;
  assign n717 = n708 ^ n705 ;
  assign n718 = n703 ^ n701 ;
  assign n719 = x16 & n718 ;
  assign n720 = n719 ^ x16 ;
  assign n721 = ~n717 & n720 ;
  assign n722 = n721 ^ n720 ;
  assign n723 = n716 & n722 ;
  assign n724 = n723 ^ n722 ;
  assign n817 = n816 ^ n724 ;
  assign n607 = ~n510 & ~n591 ;
  assign n606 = ~n550 & ~n591 ;
  assign n608 = n607 ^ n606 ;
  assign n551 = n550 ^ n510 ;
  assign n598 = n551 & n591 ;
  assign n599 = n598 ^ n551 ;
  assign n609 = n608 ^ n599 ;
  assign n595 = n510 & n550 ;
  assign n596 = n595 ^ n510 ;
  assign n597 = n596 ^ n550 ;
  assign n600 = n599 ^ n597 ;
  assign n436 = x24 & ~x32 ;
  assign n401 = x32 ^ x24 ;
  assign n434 = x25 & ~x33 ;
  assign n435 = ~n401 & n434 ;
  assign n437 = n436 ^ n435 ;
  assign n402 = x33 ^ x25 ;
  assign n403 = ~n401 & ~n402 ;
  assign n431 = x26 & ~x34 ;
  assign n404 = x34 ^ x26 ;
  assign n429 = x27 & ~x35 ;
  assign n430 = ~n404 & n429 ;
  assign n432 = n431 ^ n430 ;
  assign n433 = n403 & n432 ;
  assign n438 = n437 ^ n433 ;
  assign n405 = x35 ^ x27 ;
  assign n406 = ~n404 & ~n405 ;
  assign n407 = n403 & n406 ;
  assign n425 = x28 & ~x36 ;
  assign n408 = x36 ^ x28 ;
  assign n423 = x29 & ~x37 ;
  assign n424 = ~n408 & n423 ;
  assign n426 = n425 ^ n424 ;
  assign n409 = x37 ^ x29 ;
  assign n410 = ~n408 & ~n409 ;
  assign n420 = x30 & ~x38 ;
  assign n411 = x38 ^ x30 ;
  assign n416 = x31 & x39 ;
  assign n417 = n416 ^ x31 ;
  assign n418 = n411 & n417 ;
  assign n419 = n418 ^ n417 ;
  assign n421 = n420 ^ n419 ;
  assign n422 = n410 & n421 ;
  assign n427 = n426 ^ n422 ;
  assign n428 = n407 & n427 ;
  assign n439 = n438 ^ n428 ;
  assign n412 = x39 ^ x31 ;
  assign n413 = ~n411 & ~n412 ;
  assign n414 = n410 & n413 ;
  assign n415 = n407 & n414 ;
  assign n440 = n439 ^ n415 ;
  assign n246 = x24 & ~x40 ;
  assign n211 = x40 ^ x24 ;
  assign n244 = x25 & ~x41 ;
  assign n245 = ~n211 & n244 ;
  assign n247 = n246 ^ n245 ;
  assign n212 = x41 ^ x25 ;
  assign n213 = ~n211 & ~n212 ;
  assign n241 = x26 & ~x42 ;
  assign n214 = x42 ^ x26 ;
  assign n239 = x27 & ~x43 ;
  assign n240 = ~n214 & n239 ;
  assign n242 = n241 ^ n240 ;
  assign n243 = n213 & n242 ;
  assign n248 = n247 ^ n243 ;
  assign n215 = x43 ^ x27 ;
  assign n216 = ~n214 & ~n215 ;
  assign n217 = n213 & n216 ;
  assign n235 = x28 & ~x44 ;
  assign n218 = x44 ^ x28 ;
  assign n233 = x29 & ~x45 ;
  assign n234 = ~n218 & n233 ;
  assign n236 = n235 ^ n234 ;
  assign n219 = x45 ^ x29 ;
  assign n220 = ~n218 & ~n219 ;
  assign n230 = x30 & ~x46 ;
  assign n221 = x46 ^ x30 ;
  assign n226 = x31 & x47 ;
  assign n227 = n226 ^ x31 ;
  assign n228 = n221 & n227 ;
  assign n229 = n228 ^ n227 ;
  assign n231 = n230 ^ n229 ;
  assign n232 = n220 & n231 ;
  assign n237 = n236 ^ n232 ;
  assign n238 = n217 & n237 ;
  assign n249 = n248 ^ n238 ;
  assign n222 = x47 ^ x31 ;
  assign n223 = ~n221 & ~n222 ;
  assign n224 = n220 & n223 ;
  assign n225 = n217 & n224 ;
  assign n250 = n249 ^ n225 ;
  assign n470 = n440 ^ n250 ;
  assign n592 = n591 ^ n551 ;
  assign n593 = n470 & n592 ;
  assign n594 = n593 ^ n470 ;
  assign n601 = n600 ^ n594 ;
  assign n602 = n250 & n440 ;
  assign n603 = n602 ^ n594 ;
  assign n604 = ~n601 & n603 ;
  assign n605 = n604 ^ n594 ;
  assign n610 = n609 ^ n605 ;
  assign n611 = n602 ^ n601 ;
  assign n612 = n592 ^ n470 ;
  assign n613 = x24 & n612 ;
  assign n614 = ~n611 & n613 ;
  assign n615 = n614 ^ n613 ;
  assign n616 = n610 & n615 ;
  assign n617 = n616 ^ n615 ;
  assign n818 = n817 ^ n617 ;
  assign n458 = ~n318 & ~n399 ;
  assign n457 = ~n358 & ~n399 ;
  assign n459 = n458 ^ n457 ;
  assign n359 = n358 ^ n318 ;
  assign n448 = n359 & n399 ;
  assign n449 = n448 ^ n359 ;
  assign n460 = n459 ^ n449 ;
  assign n445 = n318 & n358 ;
  assign n446 = n445 ^ n318 ;
  assign n447 = n446 ^ n358 ;
  assign n450 = n449 ^ n447 ;
  assign n400 = n399 ^ n359 ;
  assign n206 = x32 & ~x40 ;
  assign n171 = x40 ^ x32 ;
  assign n204 = x33 & ~x41 ;
  assign n205 = ~n171 & n204 ;
  assign n207 = n206 ^ n205 ;
  assign n172 = x41 ^ x33 ;
  assign n173 = ~n171 & ~n172 ;
  assign n201 = x34 & ~x42 ;
  assign n174 = x42 ^ x34 ;
  assign n199 = x35 & ~x43 ;
  assign n200 = ~n174 & n199 ;
  assign n202 = n201 ^ n200 ;
  assign n203 = n173 & n202 ;
  assign n208 = n207 ^ n203 ;
  assign n175 = x43 ^ x35 ;
  assign n176 = ~n174 & ~n175 ;
  assign n177 = n173 & n176 ;
  assign n195 = x36 & ~x44 ;
  assign n178 = x44 ^ x36 ;
  assign n193 = x37 & ~x45 ;
  assign n194 = ~n178 & n193 ;
  assign n196 = n195 ^ n194 ;
  assign n179 = x45 ^ x37 ;
  assign n180 = ~n178 & ~n179 ;
  assign n190 = x38 & ~x46 ;
  assign n181 = x46 ^ x38 ;
  assign n186 = x39 & x47 ;
  assign n187 = n186 ^ x39 ;
  assign n188 = n181 & n187 ;
  assign n189 = n188 ^ n187 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = n180 & n191 ;
  assign n197 = n196 ^ n192 ;
  assign n198 = n177 & n197 ;
  assign n209 = n208 ^ n198 ;
  assign n182 = x47 ^ x39 ;
  assign n183 = ~n181 & ~n182 ;
  assign n184 = n180 & n183 ;
  assign n185 = n177 & n184 ;
  assign n210 = n209 ^ n185 ;
  assign n441 = n440 ^ n210 ;
  assign n442 = n400 & n441 ;
  assign n443 = n442 ^ n400 ;
  assign n444 = n443 ^ n441 ;
  assign n451 = n450 ^ n444 ;
  assign n452 = n210 & n440 ;
  assign n453 = n452 ^ n210 ;
  assign n454 = n453 ^ n444 ;
  assign n455 = n451 & ~n454 ;
  assign n456 = n455 ^ n444 ;
  assign n461 = n460 ^ n456 ;
  assign n462 = n453 ^ n451 ;
  assign n463 = n441 ^ n400 ;
  assign n464 = x32 & n463 ;
  assign n465 = n464 ^ x32 ;
  assign n466 = n462 & n465 ;
  assign n467 = n466 ^ n465 ;
  assign n468 = ~n461 & n467 ;
  assign n469 = n468 ^ n467 ;
  assign n819 = n818 ^ n469 ;
  assign n268 = ~n88 & ~n169 ;
  assign n267 = ~n128 & ~n169 ;
  assign n269 = n268 ^ n267 ;
  assign n129 = n128 ^ n88 ;
  assign n257 = n129 & n169 ;
  assign n258 = n257 ^ n129 ;
  assign n270 = n269 ^ n258 ;
  assign n254 = n88 & n128 ;
  assign n255 = n254 ^ n88 ;
  assign n256 = n255 ^ n128 ;
  assign n259 = n258 ^ n256 ;
  assign n170 = n169 ^ n129 ;
  assign n251 = n250 ^ n210 ;
  assign n252 = n170 & n251 ;
  assign n253 = n252 ^ n251 ;
  assign n260 = n259 ^ n253 ;
  assign n261 = n210 & n250 ;
  assign n262 = n261 ^ n210 ;
  assign n263 = n262 ^ n250 ;
  assign n264 = n263 ^ n253 ;
  assign n265 = ~n260 & ~n264 ;
  assign n266 = n265 ^ n253 ;
  assign n271 = n270 ^ n266 ;
  assign n272 = n263 ^ n260 ;
  assign n273 = n251 ^ n170 ;
  assign n274 = x40 & n273 ;
  assign n275 = n272 & n274 ;
  assign n276 = n275 ^ n274 ;
  assign n277 = n271 & n276 ;
  assign n278 = n277 ^ n276 ;
  assign n820 = n819 ^ n278 ;
  assign n848 = x1 & n809 ;
  assign n849 = n848 ^ x1 ;
  assign n850 = n808 & n849 ;
  assign n851 = n850 ^ n849 ;
  assign n852 = n807 & n851 ;
  assign n853 = n852 ^ n851 ;
  assign n843 = x9 & n785 ;
  assign n844 = n784 & n843 ;
  assign n845 = n844 ^ n843 ;
  assign n846 = n783 & n845 ;
  assign n847 = n846 ^ n845 ;
  assign n854 = n853 ^ n847 ;
  assign n837 = x17 & n718 ;
  assign n838 = n837 ^ x17 ;
  assign n839 = ~n717 & n838 ;
  assign n840 = n839 ^ n838 ;
  assign n841 = n716 & n840 ;
  assign n842 = n841 ^ n840 ;
  assign n855 = n854 ^ n842 ;
  assign n832 = x25 & n612 ;
  assign n833 = ~n611 & n832 ;
  assign n834 = n833 ^ n832 ;
  assign n835 = n610 & n834 ;
  assign n836 = n835 ^ n834 ;
  assign n856 = n855 ^ n836 ;
  assign n826 = x33 & n463 ;
  assign n827 = n826 ^ x33 ;
  assign n828 = n462 & n827 ;
  assign n829 = n828 ^ n827 ;
  assign n830 = ~n461 & n829 ;
  assign n831 = n830 ^ n829 ;
  assign n857 = n856 ^ n831 ;
  assign n821 = x41 & n273 ;
  assign n822 = n272 & n821 ;
  assign n823 = n822 ^ n821 ;
  assign n824 = n271 & n823 ;
  assign n825 = n824 ^ n823 ;
  assign n858 = n857 ^ n825 ;
  assign n886 = x2 & n809 ;
  assign n887 = n886 ^ x2 ;
  assign n888 = n808 & n887 ;
  assign n889 = n888 ^ n887 ;
  assign n890 = n807 & n889 ;
  assign n891 = n890 ^ n889 ;
  assign n881 = x10 & n785 ;
  assign n882 = n784 & n881 ;
  assign n883 = n882 ^ n881 ;
  assign n884 = n783 & n883 ;
  assign n885 = n884 ^ n883 ;
  assign n892 = n891 ^ n885 ;
  assign n875 = x18 & n718 ;
  assign n876 = n875 ^ x18 ;
  assign n877 = ~n717 & n876 ;
  assign n878 = n877 ^ n876 ;
  assign n879 = n716 & n878 ;
  assign n880 = n879 ^ n878 ;
  assign n893 = n892 ^ n880 ;
  assign n870 = x26 & n612 ;
  assign n871 = ~n611 & n870 ;
  assign n872 = n871 ^ n870 ;
  assign n873 = n610 & n872 ;
  assign n874 = n873 ^ n872 ;
  assign n894 = n893 ^ n874 ;
  assign n864 = x34 & n463 ;
  assign n865 = n864 ^ x34 ;
  assign n866 = n462 & n865 ;
  assign n867 = n866 ^ n865 ;
  assign n868 = ~n461 & n867 ;
  assign n869 = n868 ^ n867 ;
  assign n895 = n894 ^ n869 ;
  assign n859 = x42 & n273 ;
  assign n860 = n272 & n859 ;
  assign n861 = n860 ^ n859 ;
  assign n862 = n271 & n861 ;
  assign n863 = n862 ^ n861 ;
  assign n896 = n895 ^ n863 ;
  assign n924 = x3 & n809 ;
  assign n925 = n924 ^ x3 ;
  assign n926 = n808 & n925 ;
  assign n927 = n926 ^ n925 ;
  assign n928 = n807 & n927 ;
  assign n929 = n928 ^ n927 ;
  assign n919 = x11 & n785 ;
  assign n920 = n784 & n919 ;
  assign n921 = n920 ^ n919 ;
  assign n922 = n783 & n921 ;
  assign n923 = n922 ^ n921 ;
  assign n930 = n929 ^ n923 ;
  assign n913 = x19 & n718 ;
  assign n914 = n913 ^ x19 ;
  assign n915 = ~n717 & n914 ;
  assign n916 = n915 ^ n914 ;
  assign n917 = n716 & n916 ;
  assign n918 = n917 ^ n916 ;
  assign n931 = n930 ^ n918 ;
  assign n908 = x27 & n612 ;
  assign n909 = ~n611 & n908 ;
  assign n910 = n909 ^ n908 ;
  assign n911 = n610 & n910 ;
  assign n912 = n911 ^ n910 ;
  assign n932 = n931 ^ n912 ;
  assign n902 = x35 & n463 ;
  assign n903 = n902 ^ x35 ;
  assign n904 = n462 & n903 ;
  assign n905 = n904 ^ n903 ;
  assign n906 = ~n461 & n905 ;
  assign n907 = n906 ^ n905 ;
  assign n933 = n932 ^ n907 ;
  assign n897 = x43 & n273 ;
  assign n898 = n272 & n897 ;
  assign n899 = n898 ^ n897 ;
  assign n900 = n271 & n899 ;
  assign n901 = n900 ^ n899 ;
  assign n934 = n933 ^ n901 ;
  assign n962 = x4 & n809 ;
  assign n963 = n962 ^ x4 ;
  assign n964 = n808 & n963 ;
  assign n965 = n964 ^ n963 ;
  assign n966 = n807 & n965 ;
  assign n967 = n966 ^ n965 ;
  assign n957 = x12 & n785 ;
  assign n958 = n784 & n957 ;
  assign n959 = n958 ^ n957 ;
  assign n960 = n783 & n959 ;
  assign n961 = n960 ^ n959 ;
  assign n968 = n967 ^ n961 ;
  assign n951 = x20 & n718 ;
  assign n952 = n951 ^ x20 ;
  assign n953 = ~n717 & n952 ;
  assign n954 = n953 ^ n952 ;
  assign n955 = n716 & n954 ;
  assign n956 = n955 ^ n954 ;
  assign n969 = n968 ^ n956 ;
  assign n946 = x28 & n612 ;
  assign n947 = ~n611 & n946 ;
  assign n948 = n947 ^ n946 ;
  assign n949 = n610 & n948 ;
  assign n950 = n949 ^ n948 ;
  assign n970 = n969 ^ n950 ;
  assign n940 = x36 & n463 ;
  assign n941 = n940 ^ x36 ;
  assign n942 = n462 & n941 ;
  assign n943 = n942 ^ n941 ;
  assign n944 = ~n461 & n943 ;
  assign n945 = n944 ^ n943 ;
  assign n971 = n970 ^ n945 ;
  assign n935 = x44 & n273 ;
  assign n936 = n272 & n935 ;
  assign n937 = n936 ^ n935 ;
  assign n938 = n271 & n937 ;
  assign n939 = n938 ^ n937 ;
  assign n972 = n971 ^ n939 ;
  assign n1000 = x5 & n809 ;
  assign n1001 = n1000 ^ x5 ;
  assign n1002 = n808 & n1001 ;
  assign n1003 = n1002 ^ n1001 ;
  assign n1004 = n807 & n1003 ;
  assign n1005 = n1004 ^ n1003 ;
  assign n995 = x13 & n785 ;
  assign n996 = n784 & n995 ;
  assign n997 = n996 ^ n995 ;
  assign n998 = n783 & n997 ;
  assign n999 = n998 ^ n997 ;
  assign n1006 = n1005 ^ n999 ;
  assign n989 = x21 & n718 ;
  assign n990 = n989 ^ x21 ;
  assign n991 = ~n717 & n990 ;
  assign n992 = n991 ^ n990 ;
  assign n993 = n716 & n992 ;
  assign n994 = n993 ^ n992 ;
  assign n1007 = n1006 ^ n994 ;
  assign n984 = x29 & n612 ;
  assign n985 = ~n611 & n984 ;
  assign n986 = n985 ^ n984 ;
  assign n987 = n610 & n986 ;
  assign n988 = n987 ^ n986 ;
  assign n1008 = n1007 ^ n988 ;
  assign n978 = x37 & n463 ;
  assign n979 = n978 ^ x37 ;
  assign n980 = n462 & n979 ;
  assign n981 = n980 ^ n979 ;
  assign n982 = ~n461 & n981 ;
  assign n983 = n982 ^ n981 ;
  assign n1009 = n1008 ^ n983 ;
  assign n973 = x45 & n273 ;
  assign n974 = n272 & n973 ;
  assign n975 = n974 ^ n973 ;
  assign n976 = n271 & n975 ;
  assign n977 = n976 ^ n975 ;
  assign n1010 = n1009 ^ n977 ;
  assign n1038 = x6 & n809 ;
  assign n1039 = n1038 ^ x6 ;
  assign n1040 = n808 & n1039 ;
  assign n1041 = n1040 ^ n1039 ;
  assign n1042 = n807 & n1041 ;
  assign n1043 = n1042 ^ n1041 ;
  assign n1033 = x14 & n785 ;
  assign n1034 = n784 & n1033 ;
  assign n1035 = n1034 ^ n1033 ;
  assign n1036 = n783 & n1035 ;
  assign n1037 = n1036 ^ n1035 ;
  assign n1044 = n1043 ^ n1037 ;
  assign n1027 = x22 & n718 ;
  assign n1028 = n1027 ^ x22 ;
  assign n1029 = ~n717 & n1028 ;
  assign n1030 = n1029 ^ n1028 ;
  assign n1031 = n716 & n1030 ;
  assign n1032 = n1031 ^ n1030 ;
  assign n1045 = n1044 ^ n1032 ;
  assign n1022 = x30 & n612 ;
  assign n1023 = ~n611 & n1022 ;
  assign n1024 = n1023 ^ n1022 ;
  assign n1025 = n610 & n1024 ;
  assign n1026 = n1025 ^ n1024 ;
  assign n1046 = n1045 ^ n1026 ;
  assign n1016 = x38 & n463 ;
  assign n1017 = n1016 ^ x38 ;
  assign n1018 = n462 & n1017 ;
  assign n1019 = n1018 ^ n1017 ;
  assign n1020 = ~n461 & n1019 ;
  assign n1021 = n1020 ^ n1019 ;
  assign n1047 = n1046 ^ n1021 ;
  assign n1011 = x46 & n273 ;
  assign n1012 = n272 & n1011 ;
  assign n1013 = n1012 ^ n1011 ;
  assign n1014 = n271 & n1013 ;
  assign n1015 = n1014 ^ n1013 ;
  assign n1048 = n1047 ^ n1015 ;
  assign n1076 = x7 & n809 ;
  assign n1077 = n1076 ^ x7 ;
  assign n1078 = n808 & n1077 ;
  assign n1079 = n1078 ^ n1077 ;
  assign n1080 = n807 & n1079 ;
  assign n1081 = n1080 ^ n1079 ;
  assign n1071 = x15 & n785 ;
  assign n1072 = n784 & n1071 ;
  assign n1073 = n1072 ^ n1071 ;
  assign n1074 = n783 & n1073 ;
  assign n1075 = n1074 ^ n1073 ;
  assign n1082 = n1081 ^ n1075 ;
  assign n1065 = x23 & n718 ;
  assign n1066 = n1065 ^ x23 ;
  assign n1067 = ~n717 & n1066 ;
  assign n1068 = n1067 ^ n1066 ;
  assign n1069 = n716 & n1068 ;
  assign n1070 = n1069 ^ n1068 ;
  assign n1083 = n1082 ^ n1070 ;
  assign n1060 = x31 & n612 ;
  assign n1061 = ~n611 & n1060 ;
  assign n1062 = n1061 ^ n1060 ;
  assign n1063 = n610 & n1062 ;
  assign n1064 = n1063 ^ n1062 ;
  assign n1084 = n1083 ^ n1064 ;
  assign n1054 = x39 & n463 ;
  assign n1055 = n1054 ^ x39 ;
  assign n1056 = n462 & n1055 ;
  assign n1057 = n1056 ^ n1055 ;
  assign n1058 = ~n461 & n1057 ;
  assign n1059 = n1058 ^ n1057 ;
  assign n1085 = n1084 ^ n1059 ;
  assign n1049 = x47 & n273 ;
  assign n1050 = n272 & n1049 ;
  assign n1051 = n1050 ^ n1049 ;
  assign n1052 = n271 & n1051 ;
  assign n1053 = n1052 ^ n1051 ;
  assign n1086 = n1085 ^ n1053 ;
  assign n1110 = n808 & n810 ;
  assign n1111 = n1110 ^ n810 ;
  assign n1112 = n807 & n1111 ;
  assign n1113 = n1112 ^ n1111 ;
  assign n1105 = n786 ^ x8 ;
  assign n1106 = n784 & n1105 ;
  assign n1107 = n1106 ^ n1105 ;
  assign n1108 = n783 & n1107 ;
  assign n1109 = n1108 ^ n1107 ;
  assign n1114 = n1113 ^ n1109 ;
  assign n1101 = ~n717 & n719 ;
  assign n1102 = n1101 ^ n719 ;
  assign n1103 = n716 & n1102 ;
  assign n1104 = n1103 ^ n1102 ;
  assign n1115 = n1114 ^ n1104 ;
  assign n1096 = n613 ^ x24 ;
  assign n1097 = ~n611 & n1096 ;
  assign n1098 = n1097 ^ n1096 ;
  assign n1099 = n610 & n1098 ;
  assign n1100 = n1099 ^ n1098 ;
  assign n1116 = n1115 ^ n1100 ;
  assign n1092 = n462 & n464 ;
  assign n1093 = n1092 ^ n464 ;
  assign n1094 = ~n461 & n1093 ;
  assign n1095 = n1094 ^ n1093 ;
  assign n1117 = n1116 ^ n1095 ;
  assign n1087 = n274 ^ x40 ;
  assign n1088 = n272 & n1087 ;
  assign n1089 = n1088 ^ n1087 ;
  assign n1090 = n271 & n1089 ;
  assign n1091 = n1090 ^ n1089 ;
  assign n1118 = n1117 ^ n1091 ;
  assign n1142 = n808 & n848 ;
  assign n1143 = n1142 ^ n848 ;
  assign n1144 = n807 & n1143 ;
  assign n1145 = n1144 ^ n1143 ;
  assign n1137 = n843 ^ x9 ;
  assign n1138 = n784 & n1137 ;
  assign n1139 = n1138 ^ n1137 ;
  assign n1140 = n783 & n1139 ;
  assign n1141 = n1140 ^ n1139 ;
  assign n1146 = n1145 ^ n1141 ;
  assign n1133 = ~n717 & n837 ;
  assign n1134 = n1133 ^ n837 ;
  assign n1135 = n716 & n1134 ;
  assign n1136 = n1135 ^ n1134 ;
  assign n1147 = n1146 ^ n1136 ;
  assign n1128 = n832 ^ x25 ;
  assign n1129 = ~n611 & n1128 ;
  assign n1130 = n1129 ^ n1128 ;
  assign n1131 = n610 & n1130 ;
  assign n1132 = n1131 ^ n1130 ;
  assign n1148 = n1147 ^ n1132 ;
  assign n1124 = n462 & n826 ;
  assign n1125 = n1124 ^ n826 ;
  assign n1126 = ~n461 & n1125 ;
  assign n1127 = n1126 ^ n1125 ;
  assign n1149 = n1148 ^ n1127 ;
  assign n1119 = n821 ^ x41 ;
  assign n1120 = n272 & n1119 ;
  assign n1121 = n1120 ^ n1119 ;
  assign n1122 = n271 & n1121 ;
  assign n1123 = n1122 ^ n1121 ;
  assign n1150 = n1149 ^ n1123 ;
  assign n1174 = n808 & n886 ;
  assign n1175 = n1174 ^ n886 ;
  assign n1176 = n807 & n1175 ;
  assign n1177 = n1176 ^ n1175 ;
  assign n1169 = n881 ^ x10 ;
  assign n1170 = n784 & n1169 ;
  assign n1171 = n1170 ^ n1169 ;
  assign n1172 = n783 & n1171 ;
  assign n1173 = n1172 ^ n1171 ;
  assign n1178 = n1177 ^ n1173 ;
  assign n1165 = ~n717 & n875 ;
  assign n1166 = n1165 ^ n875 ;
  assign n1167 = n716 & n1166 ;
  assign n1168 = n1167 ^ n1166 ;
  assign n1179 = n1178 ^ n1168 ;
  assign n1160 = n870 ^ x26 ;
  assign n1161 = ~n611 & n1160 ;
  assign n1162 = n1161 ^ n1160 ;
  assign n1163 = n610 & n1162 ;
  assign n1164 = n1163 ^ n1162 ;
  assign n1180 = n1179 ^ n1164 ;
  assign n1156 = n462 & n864 ;
  assign n1157 = n1156 ^ n864 ;
  assign n1158 = ~n461 & n1157 ;
  assign n1159 = n1158 ^ n1157 ;
  assign n1181 = n1180 ^ n1159 ;
  assign n1151 = n859 ^ x42 ;
  assign n1152 = n272 & n1151 ;
  assign n1153 = n1152 ^ n1151 ;
  assign n1154 = n271 & n1153 ;
  assign n1155 = n1154 ^ n1153 ;
  assign n1182 = n1181 ^ n1155 ;
  assign n1206 = n808 & n924 ;
  assign n1207 = n1206 ^ n924 ;
  assign n1208 = n807 & n1207 ;
  assign n1209 = n1208 ^ n1207 ;
  assign n1201 = n919 ^ x11 ;
  assign n1202 = n784 & n1201 ;
  assign n1203 = n1202 ^ n1201 ;
  assign n1204 = n783 & n1203 ;
  assign n1205 = n1204 ^ n1203 ;
  assign n1210 = n1209 ^ n1205 ;
  assign n1197 = ~n717 & n913 ;
  assign n1198 = n1197 ^ n913 ;
  assign n1199 = n716 & n1198 ;
  assign n1200 = n1199 ^ n1198 ;
  assign n1211 = n1210 ^ n1200 ;
  assign n1192 = n908 ^ x27 ;
  assign n1193 = ~n611 & n1192 ;
  assign n1194 = n1193 ^ n1192 ;
  assign n1195 = n610 & n1194 ;
  assign n1196 = n1195 ^ n1194 ;
  assign n1212 = n1211 ^ n1196 ;
  assign n1188 = n462 & n902 ;
  assign n1189 = n1188 ^ n902 ;
  assign n1190 = ~n461 & n1189 ;
  assign n1191 = n1190 ^ n1189 ;
  assign n1213 = n1212 ^ n1191 ;
  assign n1183 = n897 ^ x43 ;
  assign n1184 = n272 & n1183 ;
  assign n1185 = n1184 ^ n1183 ;
  assign n1186 = n271 & n1185 ;
  assign n1187 = n1186 ^ n1185 ;
  assign n1214 = n1213 ^ n1187 ;
  assign n1238 = n808 & n962 ;
  assign n1239 = n1238 ^ n962 ;
  assign n1240 = n807 & n1239 ;
  assign n1241 = n1240 ^ n1239 ;
  assign n1233 = n957 ^ x12 ;
  assign n1234 = n784 & n1233 ;
  assign n1235 = n1234 ^ n1233 ;
  assign n1236 = n783 & n1235 ;
  assign n1237 = n1236 ^ n1235 ;
  assign n1242 = n1241 ^ n1237 ;
  assign n1229 = ~n717 & n951 ;
  assign n1230 = n1229 ^ n951 ;
  assign n1231 = n716 & n1230 ;
  assign n1232 = n1231 ^ n1230 ;
  assign n1243 = n1242 ^ n1232 ;
  assign n1224 = n946 ^ x28 ;
  assign n1225 = ~n611 & n1224 ;
  assign n1226 = n1225 ^ n1224 ;
  assign n1227 = n610 & n1226 ;
  assign n1228 = n1227 ^ n1226 ;
  assign n1244 = n1243 ^ n1228 ;
  assign n1220 = n462 & n940 ;
  assign n1221 = n1220 ^ n940 ;
  assign n1222 = ~n461 & n1221 ;
  assign n1223 = n1222 ^ n1221 ;
  assign n1245 = n1244 ^ n1223 ;
  assign n1215 = n935 ^ x44 ;
  assign n1216 = n272 & n1215 ;
  assign n1217 = n1216 ^ n1215 ;
  assign n1218 = n271 & n1217 ;
  assign n1219 = n1218 ^ n1217 ;
  assign n1246 = n1245 ^ n1219 ;
  assign n1270 = n808 & n1000 ;
  assign n1271 = n1270 ^ n1000 ;
  assign n1272 = n807 & n1271 ;
  assign n1273 = n1272 ^ n1271 ;
  assign n1265 = n995 ^ x13 ;
  assign n1266 = n784 & n1265 ;
  assign n1267 = n1266 ^ n1265 ;
  assign n1268 = n783 & n1267 ;
  assign n1269 = n1268 ^ n1267 ;
  assign n1274 = n1273 ^ n1269 ;
  assign n1261 = ~n717 & n989 ;
  assign n1262 = n1261 ^ n989 ;
  assign n1263 = n716 & n1262 ;
  assign n1264 = n1263 ^ n1262 ;
  assign n1275 = n1274 ^ n1264 ;
  assign n1256 = n984 ^ x29 ;
  assign n1257 = ~n611 & n1256 ;
  assign n1258 = n1257 ^ n1256 ;
  assign n1259 = n610 & n1258 ;
  assign n1260 = n1259 ^ n1258 ;
  assign n1276 = n1275 ^ n1260 ;
  assign n1252 = n462 & n978 ;
  assign n1253 = n1252 ^ n978 ;
  assign n1254 = ~n461 & n1253 ;
  assign n1255 = n1254 ^ n1253 ;
  assign n1277 = n1276 ^ n1255 ;
  assign n1247 = n973 ^ x45 ;
  assign n1248 = n272 & n1247 ;
  assign n1249 = n1248 ^ n1247 ;
  assign n1250 = n271 & n1249 ;
  assign n1251 = n1250 ^ n1249 ;
  assign n1278 = n1277 ^ n1251 ;
  assign n1302 = n808 & n1038 ;
  assign n1303 = n1302 ^ n1038 ;
  assign n1304 = n807 & n1303 ;
  assign n1305 = n1304 ^ n1303 ;
  assign n1297 = n1033 ^ x14 ;
  assign n1298 = n784 & n1297 ;
  assign n1299 = n1298 ^ n1297 ;
  assign n1300 = n783 & n1299 ;
  assign n1301 = n1300 ^ n1299 ;
  assign n1306 = n1305 ^ n1301 ;
  assign n1293 = ~n717 & n1027 ;
  assign n1294 = n1293 ^ n1027 ;
  assign n1295 = n716 & n1294 ;
  assign n1296 = n1295 ^ n1294 ;
  assign n1307 = n1306 ^ n1296 ;
  assign n1288 = n1022 ^ x30 ;
  assign n1289 = ~n611 & n1288 ;
  assign n1290 = n1289 ^ n1288 ;
  assign n1291 = n610 & n1290 ;
  assign n1292 = n1291 ^ n1290 ;
  assign n1308 = n1307 ^ n1292 ;
  assign n1284 = n462 & n1016 ;
  assign n1285 = n1284 ^ n1016 ;
  assign n1286 = ~n461 & n1285 ;
  assign n1287 = n1286 ^ n1285 ;
  assign n1309 = n1308 ^ n1287 ;
  assign n1279 = n1011 ^ x46 ;
  assign n1280 = n272 & n1279 ;
  assign n1281 = n1280 ^ n1279 ;
  assign n1282 = n271 & n1281 ;
  assign n1283 = n1282 ^ n1281 ;
  assign n1310 = n1309 ^ n1283 ;
  assign n1334 = n808 & n1076 ;
  assign n1335 = n1334 ^ n1076 ;
  assign n1336 = n807 & n1335 ;
  assign n1337 = n1336 ^ n1335 ;
  assign n1329 = n1071 ^ x15 ;
  assign n1330 = n784 & n1329 ;
  assign n1331 = n1330 ^ n1329 ;
  assign n1332 = n783 & n1331 ;
  assign n1333 = n1332 ^ n1331 ;
  assign n1338 = n1337 ^ n1333 ;
  assign n1325 = ~n717 & n1065 ;
  assign n1326 = n1325 ^ n1065 ;
  assign n1327 = n716 & n1326 ;
  assign n1328 = n1327 ^ n1326 ;
  assign n1339 = n1338 ^ n1328 ;
  assign n1320 = n1060 ^ x31 ;
  assign n1321 = ~n611 & n1320 ;
  assign n1322 = n1321 ^ n1320 ;
  assign n1323 = n610 & n1322 ;
  assign n1324 = n1323 ^ n1322 ;
  assign n1340 = n1339 ^ n1324 ;
  assign n1316 = n462 & n1054 ;
  assign n1317 = n1316 ^ n1054 ;
  assign n1318 = ~n461 & n1317 ;
  assign n1319 = n1318 ^ n1317 ;
  assign n1341 = n1340 ^ n1319 ;
  assign n1311 = n1049 ^ x47 ;
  assign n1312 = n272 & n1311 ;
  assign n1313 = n1312 ^ n1311 ;
  assign n1314 = n271 & n1313 ;
  assign n1315 = n1314 ^ n1313 ;
  assign n1342 = n1341 ^ n1315 ;
  assign n1353 = n807 & n812 ;
  assign n1354 = n1353 ^ n812 ;
  assign n1351 = n783 & n787 ;
  assign n1352 = n1351 ^ n787 ;
  assign n1355 = n1354 ^ n1352 ;
  assign n1349 = n716 & n721 ;
  assign n1350 = n1349 ^ n721 ;
  assign n1356 = n1355 ^ n1350 ;
  assign n1347 = n610 & n614 ;
  assign n1348 = n1347 ^ n614 ;
  assign n1357 = n1356 ^ n1348 ;
  assign n1345 = ~n461 & n466 ;
  assign n1346 = n1345 ^ n466 ;
  assign n1358 = n1357 ^ n1346 ;
  assign n1343 = n271 & n275 ;
  assign n1344 = n1343 ^ n275 ;
  assign n1359 = n1358 ^ n1344 ;
  assign n1370 = n807 & n850 ;
  assign n1371 = n1370 ^ n850 ;
  assign n1368 = n783 & n844 ;
  assign n1369 = n1368 ^ n844 ;
  assign n1372 = n1371 ^ n1369 ;
  assign n1366 = n716 & n839 ;
  assign n1367 = n1366 ^ n839 ;
  assign n1373 = n1372 ^ n1367 ;
  assign n1364 = n610 & n833 ;
  assign n1365 = n1364 ^ n833 ;
  assign n1374 = n1373 ^ n1365 ;
  assign n1362 = ~n461 & n828 ;
  assign n1363 = n1362 ^ n828 ;
  assign n1375 = n1374 ^ n1363 ;
  assign n1360 = n271 & n822 ;
  assign n1361 = n1360 ^ n822 ;
  assign n1376 = n1375 ^ n1361 ;
  assign n1387 = n807 & n888 ;
  assign n1388 = n1387 ^ n888 ;
  assign n1385 = n783 & n882 ;
  assign n1386 = n1385 ^ n882 ;
  assign n1389 = n1388 ^ n1386 ;
  assign n1383 = n716 & n877 ;
  assign n1384 = n1383 ^ n877 ;
  assign n1390 = n1389 ^ n1384 ;
  assign n1381 = n610 & n871 ;
  assign n1382 = n1381 ^ n871 ;
  assign n1391 = n1390 ^ n1382 ;
  assign n1379 = ~n461 & n866 ;
  assign n1380 = n1379 ^ n866 ;
  assign n1392 = n1391 ^ n1380 ;
  assign n1377 = n271 & n860 ;
  assign n1378 = n1377 ^ n860 ;
  assign n1393 = n1392 ^ n1378 ;
  assign n1404 = n807 & n926 ;
  assign n1405 = n1404 ^ n926 ;
  assign n1402 = n783 & n920 ;
  assign n1403 = n1402 ^ n920 ;
  assign n1406 = n1405 ^ n1403 ;
  assign n1400 = n716 & n915 ;
  assign n1401 = n1400 ^ n915 ;
  assign n1407 = n1406 ^ n1401 ;
  assign n1398 = n610 & n909 ;
  assign n1399 = n1398 ^ n909 ;
  assign n1408 = n1407 ^ n1399 ;
  assign n1396 = ~n461 & n904 ;
  assign n1397 = n1396 ^ n904 ;
  assign n1409 = n1408 ^ n1397 ;
  assign n1394 = n271 & n898 ;
  assign n1395 = n1394 ^ n898 ;
  assign n1410 = n1409 ^ n1395 ;
  assign n1421 = n807 & n964 ;
  assign n1422 = n1421 ^ n964 ;
  assign n1419 = n783 & n958 ;
  assign n1420 = n1419 ^ n958 ;
  assign n1423 = n1422 ^ n1420 ;
  assign n1417 = n716 & n953 ;
  assign n1418 = n1417 ^ n953 ;
  assign n1424 = n1423 ^ n1418 ;
  assign n1415 = n610 & n947 ;
  assign n1416 = n1415 ^ n947 ;
  assign n1425 = n1424 ^ n1416 ;
  assign n1413 = ~n461 & n942 ;
  assign n1414 = n1413 ^ n942 ;
  assign n1426 = n1425 ^ n1414 ;
  assign n1411 = n271 & n936 ;
  assign n1412 = n1411 ^ n936 ;
  assign n1427 = n1426 ^ n1412 ;
  assign n1438 = n807 & n1002 ;
  assign n1439 = n1438 ^ n1002 ;
  assign n1436 = n783 & n996 ;
  assign n1437 = n1436 ^ n996 ;
  assign n1440 = n1439 ^ n1437 ;
  assign n1434 = n716 & n991 ;
  assign n1435 = n1434 ^ n991 ;
  assign n1441 = n1440 ^ n1435 ;
  assign n1432 = n610 & n985 ;
  assign n1433 = n1432 ^ n985 ;
  assign n1442 = n1441 ^ n1433 ;
  assign n1430 = ~n461 & n980 ;
  assign n1431 = n1430 ^ n980 ;
  assign n1443 = n1442 ^ n1431 ;
  assign n1428 = n271 & n974 ;
  assign n1429 = n1428 ^ n974 ;
  assign n1444 = n1443 ^ n1429 ;
  assign n1455 = n807 & n1040 ;
  assign n1456 = n1455 ^ n1040 ;
  assign n1453 = n783 & n1034 ;
  assign n1454 = n1453 ^ n1034 ;
  assign n1457 = n1456 ^ n1454 ;
  assign n1451 = n716 & n1029 ;
  assign n1452 = n1451 ^ n1029 ;
  assign n1458 = n1457 ^ n1452 ;
  assign n1449 = n610 & n1023 ;
  assign n1450 = n1449 ^ n1023 ;
  assign n1459 = n1458 ^ n1450 ;
  assign n1447 = ~n461 & n1018 ;
  assign n1448 = n1447 ^ n1018 ;
  assign n1460 = n1459 ^ n1448 ;
  assign n1445 = n271 & n1012 ;
  assign n1446 = n1445 ^ n1012 ;
  assign n1461 = n1460 ^ n1446 ;
  assign n1472 = n807 & n1078 ;
  assign n1473 = n1472 ^ n1078 ;
  assign n1470 = n783 & n1072 ;
  assign n1471 = n1470 ^ n1072 ;
  assign n1474 = n1473 ^ n1471 ;
  assign n1468 = n716 & n1067 ;
  assign n1469 = n1468 ^ n1067 ;
  assign n1475 = n1474 ^ n1469 ;
  assign n1466 = n610 & n1061 ;
  assign n1467 = n1466 ^ n1061 ;
  assign n1476 = n1475 ^ n1467 ;
  assign n1464 = ~n461 & n1056 ;
  assign n1465 = n1464 ^ n1056 ;
  assign n1477 = n1476 ^ n1465 ;
  assign n1462 = n271 & n1050 ;
  assign n1463 = n1462 ^ n1050 ;
  assign n1478 = n1477 ^ n1463 ;
  assign n1489 = n807 & n1110 ;
  assign n1490 = n1489 ^ n1110 ;
  assign n1487 = n783 & n1106 ;
  assign n1488 = n1487 ^ n1106 ;
  assign n1491 = n1490 ^ n1488 ;
  assign n1485 = n716 & n1101 ;
  assign n1486 = n1485 ^ n1101 ;
  assign n1492 = n1491 ^ n1486 ;
  assign n1483 = n610 & n1097 ;
  assign n1484 = n1483 ^ n1097 ;
  assign n1493 = n1492 ^ n1484 ;
  assign n1481 = ~n461 & n1092 ;
  assign n1482 = n1481 ^ n1092 ;
  assign n1494 = n1493 ^ n1482 ;
  assign n1479 = n271 & n1088 ;
  assign n1480 = n1479 ^ n1088 ;
  assign n1495 = n1494 ^ n1480 ;
  assign n1506 = n807 & n1142 ;
  assign n1507 = n1506 ^ n1142 ;
  assign n1504 = n783 & n1138 ;
  assign n1505 = n1504 ^ n1138 ;
  assign n1508 = n1507 ^ n1505 ;
  assign n1502 = n716 & n1133 ;
  assign n1503 = n1502 ^ n1133 ;
  assign n1509 = n1508 ^ n1503 ;
  assign n1500 = n610 & n1129 ;
  assign n1501 = n1500 ^ n1129 ;
  assign n1510 = n1509 ^ n1501 ;
  assign n1498 = ~n461 & n1124 ;
  assign n1499 = n1498 ^ n1124 ;
  assign n1511 = n1510 ^ n1499 ;
  assign n1496 = n271 & n1120 ;
  assign n1497 = n1496 ^ n1120 ;
  assign n1512 = n1511 ^ n1497 ;
  assign n1523 = n807 & n1174 ;
  assign n1524 = n1523 ^ n1174 ;
  assign n1521 = n783 & n1170 ;
  assign n1522 = n1521 ^ n1170 ;
  assign n1525 = n1524 ^ n1522 ;
  assign n1519 = n716 & n1165 ;
  assign n1520 = n1519 ^ n1165 ;
  assign n1526 = n1525 ^ n1520 ;
  assign n1517 = n610 & n1161 ;
  assign n1518 = n1517 ^ n1161 ;
  assign n1527 = n1526 ^ n1518 ;
  assign n1515 = ~n461 & n1156 ;
  assign n1516 = n1515 ^ n1156 ;
  assign n1528 = n1527 ^ n1516 ;
  assign n1513 = n271 & n1152 ;
  assign n1514 = n1513 ^ n1152 ;
  assign n1529 = n1528 ^ n1514 ;
  assign n1540 = n807 & n1206 ;
  assign n1541 = n1540 ^ n1206 ;
  assign n1538 = n783 & n1202 ;
  assign n1539 = n1538 ^ n1202 ;
  assign n1542 = n1541 ^ n1539 ;
  assign n1536 = n716 & n1197 ;
  assign n1537 = n1536 ^ n1197 ;
  assign n1543 = n1542 ^ n1537 ;
  assign n1534 = n610 & n1193 ;
  assign n1535 = n1534 ^ n1193 ;
  assign n1544 = n1543 ^ n1535 ;
  assign n1532 = ~n461 & n1188 ;
  assign n1533 = n1532 ^ n1188 ;
  assign n1545 = n1544 ^ n1533 ;
  assign n1530 = n271 & n1184 ;
  assign n1531 = n1530 ^ n1184 ;
  assign n1546 = n1545 ^ n1531 ;
  assign n1557 = n807 & n1238 ;
  assign n1558 = n1557 ^ n1238 ;
  assign n1555 = n783 & n1234 ;
  assign n1556 = n1555 ^ n1234 ;
  assign n1559 = n1558 ^ n1556 ;
  assign n1553 = n716 & n1229 ;
  assign n1554 = n1553 ^ n1229 ;
  assign n1560 = n1559 ^ n1554 ;
  assign n1551 = n610 & n1225 ;
  assign n1552 = n1551 ^ n1225 ;
  assign n1561 = n1560 ^ n1552 ;
  assign n1549 = ~n461 & n1220 ;
  assign n1550 = n1549 ^ n1220 ;
  assign n1562 = n1561 ^ n1550 ;
  assign n1547 = n271 & n1216 ;
  assign n1548 = n1547 ^ n1216 ;
  assign n1563 = n1562 ^ n1548 ;
  assign n1574 = n807 & n1270 ;
  assign n1575 = n1574 ^ n1270 ;
  assign n1572 = n783 & n1266 ;
  assign n1573 = n1572 ^ n1266 ;
  assign n1576 = n1575 ^ n1573 ;
  assign n1570 = n716 & n1261 ;
  assign n1571 = n1570 ^ n1261 ;
  assign n1577 = n1576 ^ n1571 ;
  assign n1568 = n610 & n1257 ;
  assign n1569 = n1568 ^ n1257 ;
  assign n1578 = n1577 ^ n1569 ;
  assign n1566 = ~n461 & n1252 ;
  assign n1567 = n1566 ^ n1252 ;
  assign n1579 = n1578 ^ n1567 ;
  assign n1564 = n271 & n1248 ;
  assign n1565 = n1564 ^ n1248 ;
  assign n1580 = n1579 ^ n1565 ;
  assign n1591 = n807 & n1302 ;
  assign n1592 = n1591 ^ n1302 ;
  assign n1589 = n783 & n1298 ;
  assign n1590 = n1589 ^ n1298 ;
  assign n1593 = n1592 ^ n1590 ;
  assign n1587 = n716 & n1293 ;
  assign n1588 = n1587 ^ n1293 ;
  assign n1594 = n1593 ^ n1588 ;
  assign n1585 = n610 & n1289 ;
  assign n1586 = n1585 ^ n1289 ;
  assign n1595 = n1594 ^ n1586 ;
  assign n1583 = ~n461 & n1284 ;
  assign n1584 = n1583 ^ n1284 ;
  assign n1596 = n1595 ^ n1584 ;
  assign n1581 = n271 & n1280 ;
  assign n1582 = n1581 ^ n1280 ;
  assign n1597 = n1596 ^ n1582 ;
  assign n1608 = n807 & n1334 ;
  assign n1609 = n1608 ^ n1334 ;
  assign n1606 = n783 & n1330 ;
  assign n1607 = n1606 ^ n1330 ;
  assign n1610 = n1609 ^ n1607 ;
  assign n1604 = n716 & n1325 ;
  assign n1605 = n1604 ^ n1325 ;
  assign n1611 = n1610 ^ n1605 ;
  assign n1602 = n610 & n1321 ;
  assign n1603 = n1602 ^ n1321 ;
  assign n1612 = n1611 ^ n1603 ;
  assign n1600 = ~n461 & n1316 ;
  assign n1601 = n1600 ^ n1316 ;
  assign n1613 = n1612 ^ n1601 ;
  assign n1598 = n271 & n1312 ;
  assign n1599 = n1598 ^ n1312 ;
  assign n1614 = n1613 ^ n1599 ;
  assign n1615 = n814 ^ n789 ;
  assign n1616 = n1615 ^ n723 ;
  assign n1617 = n1616 ^ n616 ;
  assign n1618 = n1617 ^ n468 ;
  assign n1619 = n1618 ^ n277 ;
  assign n1620 = n852 ^ n846 ;
  assign n1621 = n1620 ^ n841 ;
  assign n1622 = n1621 ^ n835 ;
  assign n1623 = n1622 ^ n830 ;
  assign n1624 = n1623 ^ n824 ;
  assign n1625 = n890 ^ n884 ;
  assign n1626 = n1625 ^ n879 ;
  assign n1627 = n1626 ^ n873 ;
  assign n1628 = n1627 ^ n868 ;
  assign n1629 = n1628 ^ n862 ;
  assign n1630 = n928 ^ n922 ;
  assign n1631 = n1630 ^ n917 ;
  assign n1632 = n1631 ^ n911 ;
  assign n1633 = n1632 ^ n906 ;
  assign n1634 = n1633 ^ n900 ;
  assign n1635 = n966 ^ n960 ;
  assign n1636 = n1635 ^ n955 ;
  assign n1637 = n1636 ^ n949 ;
  assign n1638 = n1637 ^ n944 ;
  assign n1639 = n1638 ^ n938 ;
  assign n1640 = n1004 ^ n998 ;
  assign n1641 = n1640 ^ n993 ;
  assign n1642 = n1641 ^ n987 ;
  assign n1643 = n1642 ^ n982 ;
  assign n1644 = n1643 ^ n976 ;
  assign n1645 = n1042 ^ n1036 ;
  assign n1646 = n1645 ^ n1031 ;
  assign n1647 = n1646 ^ n1025 ;
  assign n1648 = n1647 ^ n1020 ;
  assign n1649 = n1648 ^ n1014 ;
  assign n1650 = n1080 ^ n1074 ;
  assign n1651 = n1650 ^ n1069 ;
  assign n1652 = n1651 ^ n1063 ;
  assign n1653 = n1652 ^ n1058 ;
  assign n1654 = n1653 ^ n1052 ;
  assign n1655 = n1112 ^ n1108 ;
  assign n1656 = n1655 ^ n1103 ;
  assign n1657 = n1656 ^ n1099 ;
  assign n1658 = n1657 ^ n1094 ;
  assign n1659 = n1658 ^ n1090 ;
  assign n1660 = n1144 ^ n1140 ;
  assign n1661 = n1660 ^ n1135 ;
  assign n1662 = n1661 ^ n1131 ;
  assign n1663 = n1662 ^ n1126 ;
  assign n1664 = n1663 ^ n1122 ;
  assign n1665 = n1176 ^ n1172 ;
  assign n1666 = n1665 ^ n1167 ;
  assign n1667 = n1666 ^ n1163 ;
  assign n1668 = n1667 ^ n1158 ;
  assign n1669 = n1668 ^ n1154 ;
  assign n1670 = n1208 ^ n1204 ;
  assign n1671 = n1670 ^ n1199 ;
  assign n1672 = n1671 ^ n1195 ;
  assign n1673 = n1672 ^ n1190 ;
  assign n1674 = n1673 ^ n1186 ;
  assign n1675 = n1240 ^ n1236 ;
  assign n1676 = n1675 ^ n1231 ;
  assign n1677 = n1676 ^ n1227 ;
  assign n1678 = n1677 ^ n1222 ;
  assign n1679 = n1678 ^ n1218 ;
  assign n1680 = n1272 ^ n1268 ;
  assign n1681 = n1680 ^ n1263 ;
  assign n1682 = n1681 ^ n1259 ;
  assign n1683 = n1682 ^ n1254 ;
  assign n1684 = n1683 ^ n1250 ;
  assign n1685 = n1304 ^ n1300 ;
  assign n1686 = n1685 ^ n1295 ;
  assign n1687 = n1686 ^ n1291 ;
  assign n1688 = n1687 ^ n1286 ;
  assign n1689 = n1688 ^ n1282 ;
  assign n1690 = n1336 ^ n1332 ;
  assign n1691 = n1690 ^ n1327 ;
  assign n1692 = n1691 ^ n1323 ;
  assign n1693 = n1692 ^ n1318 ;
  assign n1694 = n1693 ^ n1314 ;
  assign y0 = n820 ;
  assign y1 = n858 ;
  assign y2 = n896 ;
  assign y3 = n934 ;
  assign y4 = n972 ;
  assign y5 = n1010 ;
  assign y6 = n1048 ;
  assign y7 = n1086 ;
  assign y8 = n1118 ;
  assign y9 = n1150 ;
  assign y10 = n1182 ;
  assign y11 = n1214 ;
  assign y12 = n1246 ;
  assign y13 = n1278 ;
  assign y14 = n1310 ;
  assign y15 = n1342 ;
  assign y16 = n1359 ;
  assign y17 = n1376 ;
  assign y18 = n1393 ;
  assign y19 = n1410 ;
  assign y20 = n1427 ;
  assign y21 = n1444 ;
  assign y22 = n1461 ;
  assign y23 = n1478 ;
  assign y24 = n1495 ;
  assign y25 = n1512 ;
  assign y26 = n1529 ;
  assign y27 = n1546 ;
  assign y28 = n1563 ;
  assign y29 = n1580 ;
  assign y30 = n1597 ;
  assign y31 = n1614 ;
  assign y32 = n1619 ;
  assign y33 = n1624 ;
  assign y34 = n1629 ;
  assign y35 = n1634 ;
  assign y36 = n1639 ;
  assign y37 = n1644 ;
  assign y38 = n1649 ;
  assign y39 = n1654 ;
  assign y40 = n1659 ;
  assign y41 = n1664 ;
  assign y42 = n1669 ;
  assign y43 = n1674 ;
  assign y44 = n1679 ;
  assign y45 = n1684 ;
  assign y46 = n1689 ;
  assign y47 = n1694 ;
endmodule
