module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n9 = x2 & x3 ;
  assign n10 = ~x2 & ~x3 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = x4 & n11 ;
  assign n13 = ~n9 & ~n12 ;
  assign n14 = x5 & x6 ;
  assign n15 = ~x5 & ~x6 ;
  assign n16 = ~n14 & ~n15 ;
  assign n17 = x7 & n16 ;
  assign n18 = ~n14 & ~n17 ;
  assign n19 = ~x7 & ~n16 ;
  assign n20 = ~n17 & ~n19 ;
  assign n21 = ~x1 & ~n20 ;
  assign n22 = x1 & n20 ;
  assign n23 = ~x4 & ~n11 ;
  assign n24 = ~n12 & ~n23 ;
  assign n25 = ~n22 & ~n24 ;
  assign n26 = ~n21 & ~n25 ;
  assign n27 = n18 & ~n26 ;
  assign n28 = n13 & n27 ;
  assign n29 = ~n21 & ~n22 ;
  assign n30 = ~n24 & n29 ;
  assign n31 = n24 & ~n29 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = x0 & ~n32 ;
  assign n34 = ~n28 & n33 ;
  assign n35 = ~n18 & n26 ;
  assign n36 = n13 & ~n35 ;
  assign n37 = ~n27 & ~n36 ;
  assign n38 = ~n34 & ~n37 ;
  assign y0 = ~n38 ;
endmodule
