module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 ;
  assign n16 = x2 & ~x8 ;
  assign n17 = x9 & n16 ;
  assign n11 = ~x1 & ~x8 ;
  assign n12 = ~x9 & n11 ;
  assign n13 = ~x2 & x6 ;
  assign n14 = x3 & ~n13 ;
  assign n15 = n12 & ~n14 ;
  assign n18 = n17 ^ n15 ;
  assign n22 = ~x1 & x9 ;
  assign n23 = x2 & ~x3 ;
  assign n24 = n22 & n23 ;
  assign n25 = x1 & ~x8 ;
  assign n26 = ~x0 & ~x5 ;
  assign n27 = ~n25 & n26 ;
  assign n28 = ~n24 & n27 ;
  assign n29 = ~n18 & n28 ;
  assign n19 = x0 & ~x5 ;
  assign n20 = ~n18 & n19 ;
  assign n21 = n20 ^ x5 ;
  assign n30 = n29 ^ n21 ;
  assign n31 = x8 & n30 ;
  assign n38 = ~x0 & x9 ;
  assign n39 = x1 & ~x3 ;
  assign n40 = ~n38 & n39 ;
  assign n32 = ~x2 & x5 ;
  assign n33 = x0 & ~x9 ;
  assign n41 = n32 & ~n33 ;
  assign n42 = n40 & n41 ;
  assign n36 = x5 & x6 ;
  assign n34 = x6 & ~n33 ;
  assign n35 = n32 & n34 ;
  assign n37 = n36 ^ n35 ;
  assign n43 = n42 ^ n37 ;
  assign n46 = ~x0 & ~x3 ;
  assign n47 = x6 & n46 ;
  assign n51 = x2 & x9 ;
  assign n52 = n47 & n51 ;
  assign n53 = ~n43 & n52 ;
  assign n44 = x1 & ~x9 ;
  assign n45 = ~x2 & n44 ;
  assign n48 = n45 & n47 ;
  assign n49 = ~n43 & n48 ;
  assign n50 = n49 ^ n43 ;
  assign n54 = n53 ^ n50 ;
  assign n67 = n31 & n54 ;
  assign n58 = ~x1 & ~x9 ;
  assign n59 = ~x8 & n58 ;
  assign n60 = ~x2 & ~x3 ;
  assign n61 = ~x0 & n60 ;
  assign n62 = n59 & n61 ;
  assign n63 = n30 & ~n62 ;
  assign n68 = n67 ^ n63 ;
  assign n69 = ~x0 & ~x2 ;
  assign n70 = n22 & n69 ;
  assign n71 = ~x5 & x6 ;
  assign n72 = ~n70 & n71 ;
  assign n73 = n72 ^ x6 ;
  assign n75 = x1 & x5 ;
  assign n76 = x2 & n75 ;
  assign n77 = x9 ^ x0 ;
  assign n78 = x8 & ~n77 ;
  assign n79 = n76 & n78 ;
  assign n80 = ~n73 & n79 ;
  assign n74 = x8 & n73 ;
  assign n81 = n80 ^ n74 ;
  assign n86 = x0 & ~x1 ;
  assign n87 = x2 & ~x9 ;
  assign n88 = n86 & n87 ;
  assign n82 = ~x0 & ~x1 ;
  assign n83 = ~x8 & x9 ;
  assign n84 = n82 & n83 ;
  assign n85 = n84 ^ n25 ;
  assign n89 = n88 ^ n85 ;
  assign n90 = x3 & ~x7 ;
  assign n91 = ~x5 & n90 ;
  assign n92 = n89 & n91 ;
  assign n93 = n92 ^ n90 ;
  assign n94 = ~n81 & n93 ;
  assign n95 = n68 & n94 ;
  assign n55 = ~x3 & ~x7 ;
  assign n64 = n55 & n63 ;
  assign n56 = n54 & n55 ;
  assign n57 = n31 & n56 ;
  assign n65 = n64 ^ n57 ;
  assign n66 = n65 ^ x7 ;
  assign n96 = n95 ^ n66 ;
  assign n128 = x1 & ~x7 ;
  assign n129 = x9 & n128 ;
  assign n116 = ~x3 & ~x5 ;
  assign n117 = ~n22 & n116 ;
  assign n126 = ~x1 & n117 ;
  assign n121 = ~x0 & x1 ;
  assign n122 = x7 & x9 ;
  assign n123 = n121 & n122 ;
  assign n124 = n117 & n123 ;
  assign n118 = ~x7 & ~x9 ;
  assign n119 = n86 & n118 ;
  assign n120 = ~n117 & n119 ;
  assign n125 = n124 ^ n120 ;
  assign n127 = n126 ^ n125 ;
  assign n130 = n129 ^ n127 ;
  assign n131 = ~x2 & n130 ;
  assign n136 = x3 & ~x9 ;
  assign n137 = n82 & n136 ;
  assign n138 = n137 ^ x3 ;
  assign n132 = ~x3 & x9 ;
  assign n133 = ~x1 & x2 ;
  assign n134 = n132 & n133 ;
  assign n135 = n134 ^ x1 ;
  assign n139 = n138 ^ n135 ;
  assign n147 = ~x7 & n139 ;
  assign n148 = ~x8 & ~n147 ;
  assign n140 = n118 & ~n139 ;
  assign n143 = x5 & n69 ;
  assign n141 = x2 & n86 ;
  assign n142 = n141 ^ x2 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = ~x8 & n144 ;
  assign n146 = n140 & n145 ;
  assign n149 = n148 ^ n146 ;
  assign n150 = ~n131 & n149 ;
  assign n151 = n150 ^ x8 ;
  assign n159 = x1 & ~x5 ;
  assign n160 = x7 & x8 ;
  assign n161 = n159 & n160 ;
  assign n162 = n161 ^ n129 ;
  assign n163 = ~x5 & ~x9 ;
  assign n164 = ~n128 & n163 ;
  assign n165 = ~n162 & ~n164 ;
  assign n152 = ~x5 & x7 ;
  assign n153 = x8 & n152 ;
  assign n154 = n82 & n87 ;
  assign n155 = n153 & n154 ;
  assign n166 = x0 & ~x2 ;
  assign n167 = ~x3 & n166 ;
  assign n168 = ~n155 & n167 ;
  assign n169 = ~n165 & n168 ;
  assign n170 = n151 & n169 ;
  assign n156 = ~x3 & n155 ;
  assign n157 = n151 & n156 ;
  assign n158 = n157 ^ n151 ;
  assign n171 = n170 ^ n158 ;
  assign n97 = ~x6 & x8 ;
  assign n98 = x5 & ~n97 ;
  assign n99 = ~x6 & ~x9 ;
  assign n100 = x4 & x8 ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = n98 & ~n101 ;
  assign n103 = x6 & ~x9 ;
  assign n104 = x4 & x9 ;
  assign n105 = ~n103 & ~n104 ;
  assign n106 = ~x8 & ~n36 ;
  assign n107 = ~n105 & n106 ;
  assign n108 = ~n102 & ~n107 ;
  assign n109 = ~x1 & ~x3 ;
  assign n110 = ~x7 & n69 ;
  assign n111 = n109 & n110 ;
  assign n112 = ~n108 & n111 ;
  assign n172 = ~x4 & ~x6 ;
  assign n173 = ~n112 & n172 ;
  assign n174 = ~n171 & n173 ;
  assign n175 = n96 & n174 ;
  assign n113 = ~x4 & ~n112 ;
  assign n114 = ~n96 & n113 ;
  assign n115 = n114 ^ n112 ;
  assign n176 = n175 ^ n115 ;
  assign n182 = x3 & x8 ;
  assign n183 = ~x2 & ~n182 ;
  assign n187 = n82 & ~n183 ;
  assign n188 = n187 ^ x1 ;
  assign n178 = x5 ^ x0 ;
  assign n184 = n121 & ~n178 ;
  assign n185 = n183 & n184 ;
  assign n177 = x0 & x1 ;
  assign n179 = ~x2 & x8 ;
  assign n180 = ~n178 & ~n179 ;
  assign n181 = n177 & n180 ;
  assign n186 = n185 ^ n181 ;
  assign n189 = n188 ^ n186 ;
  assign n190 = ~x2 & ~x8 ;
  assign n191 = x5 & n190 ;
  assign n196 = x5 & x8 ;
  assign n195 = x3 & ~x8 ;
  assign n197 = n196 ^ n195 ;
  assign n198 = n86 & n197 ;
  assign n199 = ~n191 & n198 ;
  assign n200 = ~n189 & n199 ;
  assign n192 = ~x1 & n191 ;
  assign n193 = ~n189 & n192 ;
  assign n194 = n193 ^ n189 ;
  assign n201 = n200 ^ n194 ;
  assign n202 = ~x6 & n201 ;
  assign n203 = ~x0 & x8 ;
  assign n204 = ~x2 & ~n203 ;
  assign n205 = ~x1 & ~x6 ;
  assign n206 = ~n177 & ~n205 ;
  assign n207 = n204 & n206 ;
  assign n212 = ~x1 & ~x2 ;
  assign n213 = ~x8 & n212 ;
  assign n210 = x6 & x8 ;
  assign n211 = n133 & n210 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = n214 ^ x2 ;
  assign n216 = x3 & ~x5 ;
  assign n217 = ~x9 & n216 ;
  assign n218 = ~n215 & n217 ;
  assign n219 = ~n207 & n218 ;
  assign n208 = n163 & n207 ;
  assign n209 = n208 ^ x9 ;
  assign n220 = n219 ^ n209 ;
  assign n221 = ~n202 & ~n220 ;
  assign n222 = ~x1 & x3 ;
  assign n223 = n190 & n222 ;
  assign n224 = n223 ^ n75 ;
  assign n225 = x0 & n224 ;
  assign n227 = x1 & x2 ;
  assign n228 = n216 & n227 ;
  assign n226 = x5 & n60 ;
  assign n229 = n228 ^ n226 ;
  assign n230 = n229 ^ x5 ;
  assign n231 = x6 & ~n230 ;
  assign n232 = ~n225 & n231 ;
  assign n233 = n232 ^ x6 ;
  assign n234 = x5 & ~x8 ;
  assign n235 = x3 & n227 ;
  assign n236 = n234 & n235 ;
  assign n237 = ~x4 & x9 ;
  assign n238 = ~n236 & n237 ;
  assign n239 = ~n233 & n238 ;
  assign n240 = n239 ^ x4 ;
  assign n241 = ~n221 & ~n240 ;
  assign n279 = n19 & n97 ;
  assign n276 = ~x0 & x5 ;
  assign n277 = n83 & n276 ;
  assign n246 = x0 & x6 ;
  assign n247 = n83 & n246 ;
  assign n278 = n277 ^ n247 ;
  assign n280 = n279 ^ n278 ;
  assign n281 = ~x2 & n280 ;
  assign n287 = ~x6 & ~x8 ;
  assign n288 = ~x9 & n287 ;
  assign n282 = ~x0 & x6 ;
  assign n283 = ~x2 & ~n282 ;
  assign n284 = ~x5 & x8 ;
  assign n285 = ~x9 & n284 ;
  assign n286 = ~n283 & n285 ;
  assign n289 = n288 ^ n286 ;
  assign n290 = ~n281 & ~n289 ;
  assign n243 = ~x6 & n26 ;
  assign n242 = x8 & x9 ;
  assign n269 = n133 & n242 ;
  assign n270 = n243 & n269 ;
  assign n252 = x5 & ~x9 ;
  assign n250 = x8 & ~x9 ;
  assign n251 = n19 & n250 ;
  assign n253 = n252 ^ n251 ;
  assign n267 = n133 & n253 ;
  assign n245 = ~x6 & x9 ;
  assign n248 = n247 ^ n245 ;
  assign n266 = n133 & ~n248 ;
  assign n268 = n267 ^ n266 ;
  assign n271 = n270 ^ n268 ;
  assign n257 = ~x0 & ~x9 ;
  assign n258 = n190 & n257 ;
  assign n255 = x0 & x8 ;
  assign n256 = n51 & n255 ;
  assign n259 = n258 ^ n256 ;
  assign n263 = ~x1 & x5 ;
  assign n264 = n259 & n263 ;
  assign n244 = n242 & n243 ;
  assign n249 = n248 ^ n244 ;
  assign n254 = n253 ^ n249 ;
  assign n260 = x5 & n133 ;
  assign n261 = n259 & n260 ;
  assign n262 = ~n254 & n261 ;
  assign n265 = n264 ^ n262 ;
  assign n272 = n271 ^ n265 ;
  assign n273 = n87 & n97 ;
  assign n291 = x1 & ~x4 ;
  assign n292 = ~n273 & n291 ;
  assign n293 = ~n272 & n292 ;
  assign n294 = ~n290 & n293 ;
  assign n274 = ~n272 & ~n273 ;
  assign n275 = ~x4 & ~n274 ;
  assign n295 = n294 ^ n275 ;
  assign n296 = ~x2 & n82 ;
  assign n297 = ~n100 & ~n234 ;
  assign n298 = n99 & ~n297 ;
  assign n299 = x6 & x9 ;
  assign n300 = x4 & n299 ;
  assign n301 = ~n298 & ~n300 ;
  assign n302 = n296 & ~n301 ;
  assign n329 = n55 & ~n302 ;
  assign n330 = ~n295 & n329 ;
  assign n331 = n330 ^ n90 ;
  assign n332 = ~n241 & n331 ;
  assign n333 = n332 ^ x7 ;
  assign n313 = ~x2 & x9 ;
  assign n314 = n86 & n313 ;
  assign n315 = n314 ^ n69 ;
  assign n320 = ~x8 & ~n315 ;
  assign n318 = n44 & n179 ;
  assign n316 = n16 & ~n82 ;
  assign n317 = ~n315 & n316 ;
  assign n319 = n318 ^ n317 ;
  assign n321 = n320 ^ n319 ;
  assign n323 = ~x7 & ~n154 ;
  assign n324 = n321 & n323 ;
  assign n322 = ~n154 & ~n321 ;
  assign n325 = n324 ^ n322 ;
  assign n303 = ~x6 & n116 ;
  assign n304 = ~x4 & n303 ;
  assign n326 = x7 & n304 ;
  assign n327 = ~n325 & n326 ;
  assign n305 = ~x7 & n154 ;
  assign n306 = n304 & n305 ;
  assign n310 = x3 & n306 ;
  assign n307 = ~x3 & n306 ;
  assign n308 = ~n302 & n307 ;
  assign n309 = ~n295 & n308 ;
  assign n311 = n310 ^ n309 ;
  assign n312 = ~n241 & n311 ;
  assign n328 = n327 ^ n312 ;
  assign n334 = n333 ^ n328 ;
  assign n406 = x2 & ~n97 ;
  assign n407 = x1 & ~n406 ;
  assign n408 = x5 & ~n183 ;
  assign n409 = ~n407 & n408 ;
  assign n410 = ~n44 & ~n195 ;
  assign n411 = ~x6 & ~n136 ;
  assign n412 = ~n410 & n411 ;
  assign n413 = x1 & n132 ;
  assign n414 = x6 & ~x8 ;
  assign n415 = ~x4 & n414 ;
  assign n416 = n413 & n415 ;
  assign n417 = n416 ^ x4 ;
  assign n418 = ~n412 & ~n417 ;
  assign n419 = ~n409 & n418 ;
  assign n426 = x3 & x5 ;
  assign n424 = ~x5 & ~x8 ;
  assign n422 = ~x2 & x3 ;
  assign n423 = x8 & n422 ;
  assign n425 = n424 ^ n423 ;
  assign n427 = n426 ^ n425 ;
  assign n428 = n44 & ~n427 ;
  assign n420 = ~x3 & n71 ;
  assign n421 = n12 & n420 ;
  assign n429 = n428 ^ n421 ;
  assign n438 = ~x8 & n22 ;
  assign n430 = x1 & x8 ;
  assign n432 = n99 & ~n430 ;
  assign n431 = ~x9 & n430 ;
  assign n433 = n432 ^ n431 ;
  assign n436 = ~x2 & ~n433 ;
  assign n434 = n22 & n190 ;
  assign n435 = ~n433 & n434 ;
  assign n437 = n436 ^ n435 ;
  assign n439 = n438 ^ n437 ;
  assign n440 = x3 & n439 ;
  assign n441 = ~n429 & ~n440 ;
  assign n442 = n419 & n441 ;
  assign n347 = ~x1 & x6 ;
  assign n348 = x8 & n347 ;
  assign n346 = n227 & n299 ;
  assign n349 = n348 ^ n346 ;
  assign n352 = x2 & x3 ;
  assign n353 = ~x9 & n352 ;
  assign n354 = ~n349 & n353 ;
  assign n350 = n195 & ~n349 ;
  assign n351 = n350 ^ x3 ;
  assign n355 = n354 ^ n351 ;
  assign n359 = x1 & ~x6 ;
  assign n360 = n359 ^ n22 ;
  assign n361 = n360 ^ n99 ;
  assign n362 = n179 & ~n361 ;
  assign n356 = x9 ^ x1 ;
  assign n357 = ~x8 & ~n356 ;
  assign n358 = n60 & n357 ;
  assign n363 = n362 ^ n358 ;
  assign n364 = n19 & ~n363 ;
  assign n365 = ~n355 & n364 ;
  assign n366 = n365 ^ n19 ;
  assign n367 = ~x4 & n366 ;
  assign n445 = ~x7 & ~n367 ;
  assign n369 = x5 & x9 ;
  assign n370 = ~n255 & n369 ;
  assign n368 = ~x9 & n196 ;
  assign n371 = n370 ^ n368 ;
  assign n372 = ~n51 & n159 ;
  assign n373 = n372 ^ x1 ;
  assign n374 = ~n371 & n373 ;
  assign n376 = x9 ^ x8 ;
  assign n377 = ~n58 & ~n376 ;
  assign n378 = n23 & ~n377 ;
  assign n379 = ~n374 & n378 ;
  assign n375 = ~x3 & n374 ;
  assign n380 = n379 ^ n375 ;
  assign n381 = x5 & ~n222 ;
  assign n382 = ~x8 & ~x9 ;
  assign n387 = ~x2 & n382 ;
  assign n388 = ~n381 & n387 ;
  assign n389 = x9 & ~n60 ;
  assign n390 = ~x1 & x8 ;
  assign n391 = x0 & n390 ;
  assign n392 = n389 & n391 ;
  assign n393 = ~n388 & n392 ;
  assign n394 = ~n380 & n393 ;
  assign n383 = n166 & n382 ;
  assign n384 = ~n381 & n383 ;
  assign n385 = ~n380 & n384 ;
  assign n386 = n385 ^ n380 ;
  assign n395 = n394 ^ n386 ;
  assign n399 = ~n19 & n172 ;
  assign n396 = n19 & n172 ;
  assign n397 = ~n363 & n396 ;
  assign n398 = ~n355 & n397 ;
  assign n400 = n399 ^ n398 ;
  assign n443 = ~x7 & n400 ;
  assign n444 = n395 & n443 ;
  assign n446 = n445 ^ n444 ;
  assign n336 = x1 & ~n38 ;
  assign n337 = x0 & x7 ;
  assign n338 = n242 & n337 ;
  assign n339 = n338 ^ x0 ;
  assign n340 = n336 & ~n339 ;
  assign n335 = n11 & n33 ;
  assign n341 = n340 ^ n335 ;
  assign n342 = ~x5 & ~x6 ;
  assign n343 = ~x4 & n60 ;
  assign n344 = n342 & n343 ;
  assign n345 = n341 & n344 ;
  assign n447 = n287 ^ n250 ;
  assign n448 = ~x5 & ~n447 ;
  assign n449 = ~x2 & x4 ;
  assign n450 = n109 & n449 ;
  assign n451 = ~n448 & n450 ;
  assign n452 = n451 ^ x4 ;
  assign n453 = ~x0 & ~n452 ;
  assign n454 = ~n345 & n453 ;
  assign n455 = n446 & n454 ;
  assign n456 = ~n442 & n455 ;
  assign n401 = n395 & n400 ;
  assign n402 = n401 ^ n367 ;
  assign n403 = ~x7 & n402 ;
  assign n404 = ~n345 & n403 ;
  assign n405 = n404 ^ n345 ;
  assign n457 = n456 ^ n405 ;
  assign n557 = n116 & n414 ;
  assign n555 = n97 & n426 ;
  assign n556 = n555 ^ n216 ;
  assign n558 = n557 ^ n556 ;
  assign n562 = ~x2 & n291 ;
  assign n563 = ~n558 & n562 ;
  assign n552 = ~x8 & n163 ;
  assign n551 = n97 & n369 ;
  assign n553 = n552 ^ n551 ;
  assign n554 = ~n71 & ~n553 ;
  assign n559 = x2 & n291 ;
  assign n560 = ~n558 & n559 ;
  assign n561 = n554 & n560 ;
  assign n564 = n563 ^ n561 ;
  assign n545 = x6 & ~n60 ;
  assign n546 = ~n136 & ~n545 ;
  assign n547 = x2 & n71 ;
  assign n548 = ~x1 & ~x4 ;
  assign n549 = ~n547 & n548 ;
  assign n550 = n546 & n549 ;
  assign n565 = n564 ^ n550 ;
  assign n579 = n565 ^ x4 ;
  assign n567 = ~x3 & x4 ;
  assign n568 = n212 & n567 ;
  assign n569 = x6 ^ x5 ;
  assign n571 = ~x5 & ~n569 ;
  assign n572 = ~n242 & n571 ;
  assign n573 = n568 & n572 ;
  assign n570 = n568 & ~n569 ;
  assign n574 = n573 ^ n570 ;
  assign n580 = ~x0 & ~n574 ;
  assign n581 = n579 & n580 ;
  assign n582 = n581 ^ x0 ;
  assign n528 = ~n163 & ~n287 ;
  assign n529 = ~x2 & ~n528 ;
  assign n531 = x5 & ~x6 ;
  assign n532 = n250 & n531 ;
  assign n530 = n159 & n245 ;
  assign n533 = n532 ^ n530 ;
  assign n534 = x3 & ~n533 ;
  assign n535 = ~n529 & n534 ;
  assign n536 = n535 ^ x3 ;
  assign n539 = ~x9 & n71 ;
  assign n540 = n430 & n539 ;
  assign n541 = ~n536 & n540 ;
  assign n519 = n60 & n71 ;
  assign n518 = ~x6 & n352 ;
  assign n520 = n519 ^ n518 ;
  assign n521 = n520 ^ n71 ;
  assign n514 = x3 & ~x6 ;
  assign n523 = n83 & n514 ;
  assign n524 = ~n521 & n523 ;
  assign n522 = x9 & ~n521 ;
  assign n525 = n524 ^ n522 ;
  assign n515 = ~n71 & ~n514 ;
  assign n516 = n382 & n515 ;
  assign n517 = n516 ^ n250 ;
  assign n526 = n525 ^ n517 ;
  assign n527 = ~x1 & ~n526 ;
  assign n537 = n527 & ~n536 ;
  assign n538 = n537 ^ n536 ;
  assign n542 = n541 ^ n538 ;
  assign n566 = ~x0 & ~x4 ;
  assign n575 = n566 & ~n574 ;
  assign n576 = n565 & n575 ;
  assign n458 = x0 & ~x4 ;
  assign n577 = n576 ^ n458 ;
  assign n578 = n542 & n577 ;
  assign n583 = n582 ^ n578 ;
  assign n584 = ~x7 & ~n583 ;
  assign n461 = ~x3 & x5 ;
  assign n468 = n83 & n461 ;
  assign n495 = n216 & n468 ;
  assign n493 = n97 & n216 ;
  assign n494 = n468 & n493 ;
  assign n496 = n495 ^ n494 ;
  assign n469 = n468 ^ x3 ;
  assign n467 = ~x6 & ~n195 ;
  assign n474 = n32 & n250 ;
  assign n466 = n87 & ~n197 ;
  assign n475 = n474 ^ n466 ;
  assign n491 = n467 & n475 ;
  assign n492 = ~n469 & n491 ;
  assign n497 = n496 ^ n492 ;
  assign n487 = n467 & ~n475 ;
  assign n473 = x2 & n216 ;
  assign n488 = ~n469 & n473 ;
  assign n489 = n487 & n488 ;
  assign n485 = x2 & ~n216 ;
  assign n486 = n467 & n485 ;
  assign n490 = n489 ^ n486 ;
  assign n498 = n497 ^ n490 ;
  assign n480 = ~x2 & ~x6 ;
  assign n481 = ~n195 & n480 ;
  assign n482 = ~n469 & n481 ;
  assign n479 = n469 & n473 ;
  assign n483 = n482 ^ n479 ;
  assign n476 = ~n467 & n475 ;
  assign n477 = n473 & n476 ;
  assign n470 = n467 & n469 ;
  assign n471 = n466 & n470 ;
  assign n460 = ~x2 & n216 ;
  assign n463 = ~x9 & n23 ;
  assign n462 = n250 & n461 ;
  assign n464 = n463 ^ n462 ;
  assign n465 = n460 & n464 ;
  assign n472 = n471 ^ n465 ;
  assign n478 = n477 ^ n472 ;
  assign n484 = n483 ^ n478 ;
  assign n499 = n498 ^ n484 ;
  assign n502 = n191 & n205 ;
  assign n508 = n58 & ~n420 ;
  assign n509 = ~n502 & n508 ;
  assign n510 = ~n499 & n509 ;
  assign n503 = ~x3 & ~x9 ;
  assign n504 = n71 & n503 ;
  assign n505 = n504 ^ x9 ;
  assign n506 = ~n502 & ~n505 ;
  assign n507 = n499 & n506 ;
  assign n511 = n510 ^ n507 ;
  assign n459 = x1 & x9 ;
  assign n500 = n459 & ~n499 ;
  assign n501 = n500 ^ x9 ;
  assign n512 = n511 ^ n501 ;
  assign n513 = n458 & ~n512 ;
  assign n543 = ~x7 & ~n542 ;
  assign n544 = n513 & n543 ;
  assign n585 = n584 ^ n544 ;
  assign n586 = x2 & ~n82 ;
  assign n587 = ~x4 & n586 ;
  assign n588 = x4 ^ x3 ;
  assign n589 = n296 & n588 ;
  assign n590 = ~n587 & ~n589 ;
  assign n591 = ~x7 & n36 ;
  assign n592 = ~n590 & n591 ;
  assign n593 = x3 & ~x4 ;
  assign n594 = ~n296 & n593 ;
  assign n595 = n296 & n567 ;
  assign n596 = ~n594 & ~n595 ;
  assign n597 = n591 & ~n596 ;
  assign n665 = x9 & n75 ;
  assign n666 = n255 & n665 ;
  assign n661 = ~x1 & ~x5 ;
  assign n662 = x2 & ~n661 ;
  assign n663 = n99 & n255 ;
  assign n664 = ~n662 & n663 ;
  assign n667 = n666 ^ n664 ;
  assign n650 = ~x0 & x2 ;
  assign n659 = ~n163 & n650 ;
  assign n660 = x8 & n659 ;
  assign n668 = n667 ^ n660 ;
  assign n653 = x8 ^ x2 ;
  assign n654 = x6 & ~n376 ;
  assign n655 = ~n653 & n654 ;
  assign n671 = ~x7 & ~n655 ;
  assign n672 = ~n668 & n671 ;
  assign n673 = n672 ^ x7 ;
  assign n674 = n342 & n673 ;
  assign n651 = x9 & n650 ;
  assign n652 = n651 ^ n12 ;
  assign n656 = x5 & ~x7 ;
  assign n657 = ~n655 & n656 ;
  assign n658 = n652 & n657 ;
  assign n669 = n342 & ~n668 ;
  assign n670 = n658 & n669 ;
  assign n675 = n674 ^ n670 ;
  assign n680 = n44 & n69 ;
  assign n676 = x2 & n82 ;
  assign n677 = x7 & ~x9 ;
  assign n678 = x8 & ~n677 ;
  assign n679 = n676 & ~n678 ;
  assign n681 = n680 ^ n679 ;
  assign n682 = ~x2 & x7 ;
  assign n683 = n255 & n459 ;
  assign n684 = n683 ^ n382 ;
  assign n685 = n682 & n684 ;
  assign n686 = ~n681 & ~n685 ;
  assign n696 = n675 & ~n686 ;
  assign n689 = n658 & ~n668 ;
  assign n690 = n689 ^ n673 ;
  assign n697 = n696 ^ n690 ;
  assign n698 = ~x3 & x7 ;
  assign n699 = ~n697 & n698 ;
  assign n617 = x2 & x8 ;
  assign n618 = n38 & n617 ;
  assign n619 = ~x0 & ~n414 ;
  assign n620 = ~x2 & ~x9 ;
  assign n621 = ~n196 & n620 ;
  assign n622 = ~n619 & n621 ;
  assign n623 = ~n618 & ~n622 ;
  assign n624 = ~x1 & n623 ;
  assign n602 = x2 & ~x5 ;
  assign n603 = ~x6 & ~n602 ;
  assign n598 = ~x0 & ~x8 ;
  assign n604 = x9 & n598 ;
  assign n605 = ~n603 & n604 ;
  assign n600 = n32 & n83 ;
  assign n599 = n32 & n598 ;
  assign n601 = n600 ^ n599 ;
  assign n606 = n605 ^ n601 ;
  assign n607 = x9 & n255 ;
  assign n611 = x2 & x6 ;
  assign n612 = ~n382 & n611 ;
  assign n613 = ~n607 & n612 ;
  assign n614 = ~n606 & n613 ;
  assign n608 = x6 & n607 ;
  assign n609 = ~n606 & n608 ;
  assign n610 = n609 ^ n606 ;
  assign n615 = n614 ^ n610 ;
  assign n616 = x1 & ~n615 ;
  assign n625 = n624 ^ n616 ;
  assign n691 = n55 & n690 ;
  assign n687 = n55 & ~n686 ;
  assign n688 = n675 & n687 ;
  assign n692 = n691 ^ n688 ;
  assign n693 = n625 & n692 ;
  assign n635 = n86 & n382 ;
  assign n634 = x9 & n177 ;
  assign n636 = n635 ^ n634 ;
  assign n626 = ~x0 & ~x6 ;
  assign n629 = n227 & ~n626 ;
  assign n627 = n11 & n626 ;
  assign n628 = n627 ^ n626 ;
  assign n630 = n629 ^ n628 ;
  assign n632 = x9 & n630 ;
  assign n631 = x1 & n630 ;
  assign n633 = n632 ^ n631 ;
  assign n637 = n636 ^ n633 ;
  assign n638 = ~x5 & n637 ;
  assign n642 = n166 & n210 ;
  assign n641 = n16 & n121 ;
  assign n643 = n642 ^ n641 ;
  assign n644 = n643 ^ n25 ;
  assign n645 = x9 & n644 ;
  assign n639 = ~n19 & ~n598 ;
  assign n640 = n44 & n639 ;
  assign n646 = n645 ^ n640 ;
  assign n647 = n90 & ~n646 ;
  assign n648 = ~n638 & n647 ;
  assign n649 = n625 & n648 ;
  assign n694 = n693 ^ n649 ;
  assign n695 = n694 ^ x7 ;
  assign n700 = n699 ^ n695 ;
  assign n701 = x4 & n82 ;
  assign n702 = n60 & n701 ;
  assign n703 = ~n36 & ~n702 ;
  assign n704 = ~x7 & ~n703 ;
  assign n705 = ~x4 & ~n704 ;
  assign n706 = ~n700 & n705 ;
  assign n707 = n706 ^ n704 ;
  assign n750 = ~x3 & ~x6 ;
  assign n751 = x8 & n750 ;
  assign n752 = n751 ^ x6 ;
  assign n748 = ~x9 & n414 ;
  assign n746 = x9 & n203 ;
  assign n744 = ~x6 & n46 ;
  assign n745 = n250 & n744 ;
  assign n747 = n746 ^ n745 ;
  assign n749 = n748 ^ n747 ;
  assign n753 = n752 ^ n749 ;
  assign n725 = ~x3 & ~x8 ;
  assign n740 = n99 & n725 ;
  assign n754 = ~x2 & ~n740 ;
  assign n755 = ~n753 & n754 ;
  assign n736 = x3 & ~n242 ;
  assign n737 = ~n255 & ~n736 ;
  assign n738 = ~x6 & ~n737 ;
  assign n739 = ~x3 & n242 ;
  assign n741 = x2 & ~n740 ;
  assign n742 = ~n739 & n741 ;
  assign n743 = ~n738 & n742 ;
  assign n756 = n755 ^ n743 ;
  assign n729 = x3 & n190 ;
  assign n730 = n103 & n729 ;
  assign n757 = n159 & ~n730 ;
  assign n758 = n756 & n757 ;
  assign n720 = n99 & n650 ;
  assign n721 = n720 ^ n257 ;
  assign n718 = n83 & n480 ;
  assign n717 = x8 & n282 ;
  assign n719 = n718 ^ n717 ;
  assign n722 = n721 ^ n719 ;
  assign n723 = x3 & n722 ;
  assign n724 = x2 & ~n382 ;
  assign n726 = ~x6 & ~n725 ;
  assign n727 = n724 & ~n726 ;
  assign n728 = ~n723 & ~n727 ;
  assign n731 = n33 & n210 ;
  assign n732 = n731 ^ n258 ;
  assign n733 = n661 & ~n732 ;
  assign n734 = ~n730 & n733 ;
  assign n735 = n728 & n734 ;
  assign n759 = n758 ^ n735 ;
  assign n760 = n759 ^ x5 ;
  assign n785 = n26 & n250 ;
  assign n786 = n785 ^ n250 ;
  assign n782 = x2 & x5 ;
  assign n783 = n83 & n782 ;
  assign n781 = x8 & n166 ;
  assign n784 = n783 ^ n781 ;
  assign n787 = n786 ^ n784 ;
  assign n794 = ~x3 & n787 ;
  assign n795 = n426 & n620 ;
  assign n796 = ~n794 & ~n795 ;
  assign n773 = ~n87 & ~n426 ;
  assign n779 = ~x0 & ~n773 ;
  assign n777 = x3 & n32 ;
  assign n774 = ~x0 & x3 ;
  assign n775 = n32 & n774 ;
  assign n776 = ~n773 & n775 ;
  assign n778 = n777 ^ n776 ;
  assign n780 = n779 ^ n778 ;
  assign n790 = ~x8 & n620 ;
  assign n791 = n426 & n790 ;
  assign n788 = n725 & n787 ;
  assign n789 = n788 ^ x8 ;
  assign n792 = n791 ^ n789 ;
  assign n793 = n780 & ~n792 ;
  assign n797 = n796 ^ n793 ;
  assign n769 = x8 & n369 ;
  assign n770 = n352 & n769 ;
  assign n798 = n359 & ~n770 ;
  assign n799 = n797 & n798 ;
  assign n761 = x0 & x3 ;
  assign n762 = x2 & n382 ;
  assign n763 = n761 & n762 ;
  assign n764 = ~n352 & n376 ;
  assign n765 = n32 & ~n761 ;
  assign n766 = n765 ^ x5 ;
  assign n767 = ~n764 & n766 ;
  assign n768 = ~n763 & ~n767 ;
  assign n771 = n205 & ~n770 ;
  assign n772 = n768 & n771 ;
  assign n800 = n799 ^ n772 ;
  assign n801 = n800 ^ x6 ;
  assign n710 = n376 & n650 ;
  assign n708 = x8 & n677 ;
  assign n709 = n166 & n708 ;
  assign n711 = n710 ^ n709 ;
  assign n712 = n109 & n342 ;
  assign n802 = ~x4 & ~x7 ;
  assign n803 = n712 & n802 ;
  assign n804 = n711 & n803 ;
  assign n805 = n804 ^ n802 ;
  assign n806 = n801 & n805 ;
  assign n807 = n760 & n806 ;
  assign n713 = n711 & n712 ;
  assign n714 = ~x4 & x7 ;
  assign n715 = ~n713 & n714 ;
  assign n716 = n715 ^ x4 ;
  assign n808 = n807 ^ n716 ;
  assign n809 = ~x5 & ~x7 ;
  assign n810 = n595 & n809 ;
  assign n811 = ~x6 & n810 ;
  assign n812 = n808 & ~n811 ;
  assign n884 = ~x8 & n650 ;
  assign n882 = ~x9 & n179 ;
  assign n883 = n882 ^ n257 ;
  assign n885 = n884 ^ n883 ;
  assign n886 = ~x1 & n885 ;
  assign n880 = ~x0 & n190 ;
  assign n881 = n459 & n880 ;
  assign n887 = n886 ^ n881 ;
  assign n888 = n304 & n887 ;
  assign n889 = ~n810 & n888 ;
  assign n892 = x7 & n889 ;
  assign n834 = n227 & ~n426 ;
  assign n849 = n234 & n834 ;
  assign n850 = n849 ^ x8 ;
  assign n851 = ~x9 & ~n850 ;
  assign n841 = n116 & n166 ;
  assign n839 = n212 & n426 ;
  assign n837 = n86 & n461 ;
  assign n836 = n23 & n86 ;
  assign n838 = n837 ^ n836 ;
  assign n840 = n839 ^ n838 ;
  assign n842 = n841 ^ n840 ;
  assign n843 = ~x9 & ~n842 ;
  assign n845 = x8 & n19 ;
  assign n846 = n834 & n845 ;
  assign n847 = n843 & ~n846 ;
  assign n835 = x8 & ~n834 ;
  assign n844 = ~n835 & n843 ;
  assign n848 = n847 ^ n844 ;
  assign n852 = n851 ^ n848 ;
  assign n824 = ~n426 & ~n602 ;
  assign n825 = x1 & x3 ;
  assign n826 = ~n179 & n825 ;
  assign n827 = n826 ^ x1 ;
  assign n828 = ~n824 & n827 ;
  assign n829 = n179 & ~n276 ;
  assign n830 = x9 & n222 ;
  assign n831 = n829 & n830 ;
  assign n832 = n831 ^ x9 ;
  assign n833 = ~n828 & n832 ;
  assign n853 = n852 ^ n833 ;
  assign n856 = ~x6 & ~n853 ;
  assign n813 = n263 ^ n116 ;
  assign n814 = ~x2 & ~n58 ;
  assign n815 = ~n132 & n814 ;
  assign n816 = n813 & n815 ;
  assign n817 = n32 & n58 ;
  assign n818 = n817 ^ n413 ;
  assign n819 = ~x0 & n818 ;
  assign n820 = n356 & ~n661 ;
  assign n821 = n23 & ~n820 ;
  assign n822 = ~n819 & ~n821 ;
  assign n823 = ~n816 & n822 ;
  assign n854 = n287 & n853 ;
  assign n855 = ~n823 & n854 ;
  assign n857 = n856 ^ n855 ;
  assign n862 = n103 & n203 ;
  assign n860 = ~x9 & n347 ;
  assign n858 = x1 & x6 ;
  assign n859 = ~n203 & n858 ;
  assign n861 = n860 ^ n859 ;
  assign n863 = n862 ^ n861 ;
  assign n864 = n460 & ~n863 ;
  assign n865 = n864 ^ n216 ;
  assign n872 = ~x7 & ~n865 ;
  assign n866 = n86 & ~n382 ;
  assign n867 = n866 ^ x0 ;
  assign n868 = ~x6 & ~x7 ;
  assign n869 = ~n25 & n868 ;
  assign n870 = ~n867 & n869 ;
  assign n871 = n865 & n870 ;
  assign n873 = n872 ^ n871 ;
  assign n890 = n873 & n889 ;
  assign n891 = ~n857 & n890 ;
  assign n893 = n892 ^ n891 ;
  assign n874 = ~x4 & ~n810 ;
  assign n877 = ~x7 & n874 ;
  assign n875 = n873 & n874 ;
  assign n876 = ~n857 & n875 ;
  assign n878 = n877 ^ n876 ;
  assign n879 = n878 ^ n810 ;
  assign n894 = n893 ^ n879 ;
  assign n895 = ~x1 & ~n382 ;
  assign n896 = x2 & n514 ;
  assign n897 = n19 & n896 ;
  assign n898 = ~x7 & ~n897 ;
  assign n899 = ~n895 & ~n898 ;
  assign n900 = ~x2 & n109 ;
  assign n901 = ~x7 & ~n900 ;
  assign n902 = x0 & ~n901 ;
  assign n903 = ~x5 & ~n23 ;
  assign n904 = x6 & ~n903 ;
  assign n905 = n450 ^ x4 ;
  assign n906 = x7 & ~n23 ;
  assign n907 = ~n905 & ~n906 ;
  assign n908 = ~n904 & n907 ;
  assign n909 = ~n902 & n908 ;
  assign n910 = ~n899 & n909 ;
  assign n926 = n163 & ~n203 ;
  assign n927 = n60 & n926 ;
  assign n924 = n203 & n299 ;
  assign n925 = n422 & n924 ;
  assign n928 = n927 ^ n925 ;
  assign n929 = n928 ^ n60 ;
  assign n931 = n551 ^ x6 ;
  assign n932 = ~x3 & n931 ;
  assign n918 = ~x5 & ~n242 ;
  assign n930 = n518 & n918 ;
  assign n933 = n932 ^ n930 ;
  assign n934 = ~n929 & ~n933 ;
  assign n935 = x1 & n934 ;
  assign n936 = n910 & n935 ;
  assign n911 = x3 & ~n299 ;
  assign n912 = ~x6 & ~n369 ;
  assign n913 = n203 & ~n912 ;
  assign n914 = n911 & ~n913 ;
  assign n915 = ~n342 & n567 ;
  assign n916 = ~x2 & ~n915 ;
  assign n917 = ~n914 & n916 ;
  assign n919 = n23 & ~n382 ;
  assign n920 = ~n918 & n919 ;
  assign n921 = ~x1 & ~n920 ;
  assign n922 = ~n917 & n921 ;
  assign n923 = n910 & n922 ;
  assign n937 = n936 ^ n923 ;
  assign n938 = ~x7 & n342 ;
  assign n939 = x8 & ~n336 ;
  assign n940 = ~x1 & ~n33 ;
  assign n941 = x2 & n593 ;
  assign n942 = ~n940 & n941 ;
  assign n943 = ~n939 & n942 ;
  assign n944 = ~n595 & ~n943 ;
  assign n945 = n938 & ~n944 ;
  assign y0 = n176 ;
  assign y1 = ~n334 ;
  assign y2 = n457 ;
  assign y3 = n585 ;
  assign y4 = n592 ;
  assign y5 = n597 ;
  assign y6 = ~n707 ;
  assign y7 = n812 ;
  assign y8 = ~n894 ;
  assign y9 = n937 ;
  assign y10 = n945 ;
endmodule
