module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 ;
  assign n33 = ~x24 & ~x25 ;
  assign n34 = ~x26 & ~x27 ;
  assign n35 = n33 & n34 ;
  assign n36 = ~x22 & ~x23 ;
  assign n37 = ~x20 & ~x21 ;
  assign n38 = n36 & n37 ;
  assign n39 = n35 & n38 ;
  assign n40 = ~x8 & ~x9 ;
  assign n41 = ~x10 & ~x11 ;
  assign n42 = n40 & n41 ;
  assign n43 = ~x28 & ~x29 ;
  assign n44 = ~x30 & ~x31 ;
  assign n45 = n43 & n44 ;
  assign n46 = n42 & n45 ;
  assign n47 = n39 & n46 ;
  assign n48 = ~x0 & ~x1 ;
  assign n49 = ~x2 & ~x3 ;
  assign n50 = n48 & n49 ;
  assign n51 = ~x4 & ~x5 ;
  assign n52 = ~x6 & ~x7 ;
  assign n53 = n51 & n52 ;
  assign n54 = n50 & n53 ;
  assign n55 = ~x14 & ~x15 ;
  assign n56 = ~x12 & ~x13 ;
  assign n57 = n55 & n56 ;
  assign n58 = ~x16 & ~x17 ;
  assign n59 = ~x18 & ~x19 ;
  assign n60 = n58 & n59 ;
  assign n61 = n57 & n60 ;
  assign n62 = n54 & n61 ;
  assign n63 = n47 & n62 ;
  assign n89 = ~x0 & x1 ;
  assign n90 = n89 ^ x0 ;
  assign n86 = ~x2 & x3 ;
  assign n87 = n86 ^ x2 ;
  assign n88 = n48 & n87 ;
  assign n91 = n90 ^ n88 ;
  assign n82 = ~x4 & x5 ;
  assign n83 = n82 ^ x4 ;
  assign n79 = ~x6 & x7 ;
  assign n80 = n79 ^ x6 ;
  assign n81 = n51 & n80 ;
  assign n84 = n83 ^ n81 ;
  assign n85 = n50 & n84 ;
  assign n92 = n91 ^ n85 ;
  assign n74 = ~x8 & x9 ;
  assign n75 = n74 ^ x8 ;
  assign n71 = ~x10 & x11 ;
  assign n72 = n71 ^ x10 ;
  assign n73 = n40 & n72 ;
  assign n76 = n75 ^ n73 ;
  assign n67 = ~x12 & x13 ;
  assign n68 = n67 ^ x12 ;
  assign n64 = ~x14 & x15 ;
  assign n65 = n64 ^ x14 ;
  assign n66 = n56 & n65 ;
  assign n69 = n68 ^ n66 ;
  assign n70 = n42 & n69 ;
  assign n77 = n76 ^ n70 ;
  assign n78 = n54 & n77 ;
  assign n93 = n92 ^ n78 ;
  assign n136 = x16 & ~n93 ;
  assign n135 = x0 & n93 ;
  assign n137 = n136 ^ n135 ;
  assign n139 = x17 & ~n93 ;
  assign n138 = x1 & n93 ;
  assign n140 = n139 ^ n138 ;
  assign n141 = ~n137 & n140 ;
  assign n142 = n141 ^ n137 ;
  assign n117 = n48 & n92 ;
  assign n118 = n117 ^ n78 ;
  assign n116 = n58 & ~n93 ;
  assign n119 = n118 ^ n116 ;
  assign n131 = x18 & ~n93 ;
  assign n130 = x2 & n93 ;
  assign n132 = n131 ^ n130 ;
  assign n127 = ~x18 & x19 ;
  assign n128 = ~n93 & n127 ;
  assign n126 = n86 & n93 ;
  assign n129 = n128 ^ n126 ;
  assign n133 = n132 ^ n129 ;
  assign n134 = n119 & n133 ;
  assign n143 = n142 ^ n134 ;
  assign n112 = x20 & ~n93 ;
  assign n111 = x4 & n93 ;
  assign n113 = n112 ^ n111 ;
  assign n108 = ~x20 & x21 ;
  assign n109 = ~n93 & n108 ;
  assign n107 = n82 & n93 ;
  assign n110 = n109 ^ n107 ;
  assign n114 = n113 ^ n110 ;
  assign n99 = x22 & ~n93 ;
  assign n98 = x6 & n93 ;
  assign n100 = n99 ^ n98 ;
  assign n95 = ~x22 & x23 ;
  assign n96 = ~n93 & n95 ;
  assign n94 = n79 & n93 ;
  assign n97 = n96 ^ n94 ;
  assign n101 = n100 ^ n97 ;
  assign n104 = n37 & ~n93 ;
  assign n102 = n51 & n92 ;
  assign n103 = n102 ^ n78 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n101 & n105 ;
  assign n115 = n114 ^ n106 ;
  assign n122 = n59 & ~n93 ;
  assign n120 = n49 & n92 ;
  assign n121 = n120 ^ n78 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = n119 & n123 ;
  assign n125 = n115 & n124 ;
  assign n144 = n143 ^ n125 ;
  assign n166 = x24 & ~n93 ;
  assign n165 = x8 & n93 ;
  assign n167 = n166 ^ n165 ;
  assign n168 = ~n144 & n167 ;
  assign n164 = n137 & n144 ;
  assign n169 = n168 ^ n164 ;
  assign n172 = x25 & ~n93 ;
  assign n171 = x9 & n93 ;
  assign n173 = n172 ^ n171 ;
  assign n174 = ~n144 & n173 ;
  assign n170 = n140 & n144 ;
  assign n175 = n174 ^ n170 ;
  assign n178 = ~n169 & n175 ;
  assign n179 = n178 ^ n169 ;
  assign n156 = x27 & ~n93 ;
  assign n155 = x11 & n93 ;
  assign n157 = n156 ^ n155 ;
  assign n160 = ~n132 & n157 ;
  assign n161 = ~n144 & n160 ;
  assign n149 = x26 & ~n93 ;
  assign n148 = x10 & n93 ;
  assign n150 = n149 ^ n148 ;
  assign n158 = n150 & n157 ;
  assign n159 = ~n144 & n158 ;
  assign n162 = n161 ^ n159 ;
  assign n146 = x19 & ~n93 ;
  assign n145 = x3 & n93 ;
  assign n147 = n146 ^ n145 ;
  assign n153 = ~n132 & ~n147 ;
  assign n151 = ~n147 & n150 ;
  assign n152 = ~n144 & n151 ;
  assign n154 = n153 ^ n152 ;
  assign n163 = n162 ^ n154 ;
  assign n176 = ~n169 & ~n175 ;
  assign n177 = ~n163 & n176 ;
  assign n180 = n179 ^ n177 ;
  assign n183 = x28 & ~n93 ;
  assign n182 = x12 & n93 ;
  assign n184 = n183 ^ n182 ;
  assign n185 = ~n144 & n184 ;
  assign n181 = n113 & n144 ;
  assign n186 = n185 ^ n181 ;
  assign n187 = n163 & n186 ;
  assign n188 = n176 & n187 ;
  assign n189 = n188 ^ n169 ;
  assign n195 = x29 & ~n93 ;
  assign n194 = x13 & n93 ;
  assign n196 = n195 ^ n194 ;
  assign n197 = ~n144 & n196 ;
  assign n191 = x21 & ~n93 ;
  assign n190 = x5 & n93 ;
  assign n192 = n191 ^ n190 ;
  assign n193 = n144 & n192 ;
  assign n198 = n197 ^ n193 ;
  assign n199 = n163 & n198 ;
  assign n200 = n176 & n199 ;
  assign n201 = n200 ^ n175 ;
  assign n202 = ~n189 & n201 ;
  assign n203 = n202 ^ n189 ;
  assign n212 = ~n175 & ~n187 ;
  assign n213 = ~n144 & n150 ;
  assign n214 = n213 ^ n132 ;
  assign n215 = ~n169 & n214 ;
  assign n216 = ~n199 & n215 ;
  assign n217 = n212 & n216 ;
  assign n206 = x30 & ~n93 ;
  assign n205 = x14 & n93 ;
  assign n207 = n206 ^ n205 ;
  assign n208 = ~n144 & n207 ;
  assign n204 = n100 & n144 ;
  assign n209 = n208 ^ n204 ;
  assign n210 = ~n180 & n209 ;
  assign n211 = ~n203 & n210 ;
  assign n218 = n217 ^ n211 ;
  assign n219 = n218 ^ n189 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = 1'b0 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = n63 ;
  assign y27 = ~n93 ;
  assign y28 = ~n144 ;
  assign y29 = ~n180 ;
  assign y30 = ~n203 ;
  assign y31 = ~n219 ;
endmodule
