module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409, y63, n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419, y62, n_420, n_421, n_422, n_423, n_424, n_425, y61, n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, y60, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487, y59, n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521, y58, n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567, y57, n_568, n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616, y56, n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670, y55, n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742, n_743, y54, n_744, n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814, n_815, y53, n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892, y52, n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967, y51, n_968, n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, y50, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, y49, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, y48, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, y47, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, y46, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, y45, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, y44, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, y43, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, y42, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, y41, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, y40, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, y39, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, y38, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, y37, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, y36, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, y35, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, y34, n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, y33, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, y32, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, y31, n_3928, n_3929, n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985, n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, n_4012, n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, n_4021, n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4029, n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4048, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, n_4057, n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077, n_4078, n_4079, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085, n_4086, n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, n_4093, n_4094, n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, n_4102, n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, n_4141, y30, n_4142, n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157, n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165, n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220, n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, n_4227, n_4228, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, n_4236, n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, n_4255, n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, n_4264, n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281, n_4282, n_4283, n_4284, n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, n_4291, n_4292, n_4293, n_4294, n_4295, n_4296, n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, n_4303, n_4304, n_4305, n_4306, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312, n_4313, n_4314, n_4315, n_4316, n_4317, n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330, n_4331, n_4332, n_4333, n_4334, n_4335, n_4336, n_4337, n_4338, n_4339, n_4340, n_4341, n_4342, n_4343, n_4344, n_4345, y29, n_4346, n_4347, n_4348, n_4349, n_4350, n_4351, n_4352, n_4353, n_4354, n_4355, n_4356, n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, n_4363, n_4364, n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372, n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380, n_4381, n_4382, n_4383, n_4384, n_4385, n_4386, n_4387, n_4388, n_4389, n_4390, n_4391, n_4392, n_4393, n_4394, n_4395, n_4396, n_4397, n_4398, n_4399, n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4407, n_4408, n_4409, n_4410, n_4411, n_4412, n_4413, n_4414, n_4415, n_4416, n_4417, n_4418, n_4419, n_4420, n_4421, n_4422, n_4423, n_4424, n_4425, n_4426, n_4427, n_4428, n_4429, n_4430, n_4431, n_4432, n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439, n_4440, n_4441, n_4442, n_4443, n_4444, n_4445, n_4446, n_4447, n_4448, n_4449, n_4450, n_4451, n_4452, n_4453, n_4454, n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461, n_4462, n_4463, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469, n_4470, n_4471, n_4472, n_4473, n_4474, n_4475, n_4476, n_4477, n_4478, n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485, n_4486, n_4487, n_4488, n_4489, n_4490, n_4491, n_4492, n_4493, n_4494, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500, n_4501, n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509, n_4510, n_4511, n_4512, n_4513, n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525, n_4526, n_4527, n_4528, n_4529, n_4530, n_4531, n_4532, n_4533, n_4534, n_4535, n_4536, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4543, n_4544, n_4545, n_4546, n_4547, n_4548, n_4549, n_4550, n_4551, n_4552, n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559, n_4560, n_4561, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568, n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575, n_4576, n_4577, n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584, y28, n_4585, n_4586, n_4587, n_4588, n_4589, n_4590, n_4591, n_4592, n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600, n_4601, n_4602, n_4603, n_4604, n_4605, n_4606, n_4607, n_4608, n_4609, n_4610, n_4611, n_4612, n_4613, n_4614, n_4615, n_4616, n_4617, n_4618, n_4619, n_4620, n_4621, n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4629, n_4630, n_4631, n_4632, n_4633, n_4634, n_4635, n_4636, n_4637, n_4638, n_4639, n_4640, n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648, n_4649, n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656, n_4657, n_4658, n_4659, n_4660, n_4661, n_4662, n_4663, n_4664, n_4665, n_4666, n_4667, n_4668, n_4669, n_4670, n_4671, n_4672, n_4673, n_4674, n_4675, n_4676, n_4677, n_4678, n_4679, n_4680, n_4681, n_4682, n_4683, n_4684, n_4685, n_4686, n_4687, n_4688, n_4689, n_4690, n_4691, n_4692, n_4693, n_4694, n_4695, n_4696, n_4697, n_4698, n_4699, n_4700, n_4701, n_4702, n_4703, n_4704, n_4705, n_4706, n_4707, n_4708, n_4709, n_4710, n_4711, n_4712, n_4713, n_4714, n_4715, n_4716, n_4717, n_4718, n_4719, n_4720, n_4721, n_4722, n_4723, n_4724, n_4725, n_4726, n_4727, n_4728, n_4729, n_4730, n_4731, n_4732, n_4733, n_4734, n_4735, n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750, n_4751, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4758, n_4759, n_4760, n_4761, n_4762, n_4763, n_4764, n_4765, n_4766, n_4767, n_4768, n_4769, n_4770, n_4771, n_4772, n_4773, n_4774, n_4775, n_4776, n_4777, n_4778, n_4779, n_4780, n_4781, n_4782, n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790, n_4791, n_4792, n_4793, n_4794, n_4795, n_4796, n_4797, n_4798, n_4799, n_4800, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806, n_4807, n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814, n_4815, n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823, n_4824, n_4825, n_4826, n_4827, n_4828, n_4829, n_4830, n_4831, n_4832, n_4833, n_4834, n_4835, n_4836, n_4837, n_4838, n_4839, n_4840, n_4841, y27, n_4842, n_4843, n_4844, n_4845, n_4846, n_4847, n_4848, n_4849, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855, n_4856, n_4857, n_4858, n_4859, n_4860, n_4861, n_4862, n_4863, n_4864, n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872, n_4873, n_4874, n_4875, n_4876, n_4877, n_4878, n_4879, n_4880, n_4881, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887, n_4888, n_4889, n_4890, n_4891, n_4892, n_4893, n_4894, n_4895, n_4896, n_4897, n_4898, n_4899, n_4900, n_4901, n_4902, n_4903, n_4904, n_4905, n_4906, n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913, n_4914, n_4915, n_4916, n_4917, n_4918, n_4919, n_4920, n_4921, n_4922, n_4923, n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930, n_4931, n_4932, n_4933, n_4934, n_4935, n_4936, n_4937, n_4938, n_4939, n_4940, n_4941, n_4942, n_4943, n_4944, n_4945, n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953, n_4954, n_4955, n_4956, n_4957, n_4958, n_4959, n_4960, n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, n_4969, n_4970, n_4971, n_4972, n_4973, n_4974, n_4975, n_4976, n_4977, n_4978, n_4979, n_4980, n_4981, n_4982, n_4983, n_4984, n_4985, n_4986, n_4987, n_4988, n_4989, n_4990, n_4991, n_4992, n_4993, n_4994, n_4995, n_4996, n_4997, n_4998, n_4999, n_5000, n_5001, n_5002, n_5003, n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010, n_5011, n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018, n_5019, n_5020, n_5021, n_5022, n_5023, n_5024, n_5025, n_5026, n_5027, n_5028, n_5029, n_5030, n_5031, n_5032, n_5033, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040, n_5041, n_5042, n_5043, n_5044, n_5045, n_5046, n_5047, n_5048, n_5049, n_5050, n_5051, n_5052, n_5053, n_5054, n_5055, n_5056, n_5057, n_5058, n_5059, n_5060, n_5061, n_5062, n_5063, n_5064, n_5065, n_5066, n_5067, n_5068, n_5069, n_5070, n_5071, n_5072, n_5073, n_5074, n_5075, n_5076, n_5077, n_5078, n_5079, n_5080, n_5081, n_5082, n_5083, n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091, n_5092, n_5093, n_5094, n_5095, n_5096, n_5097, n_5098, n_5099, n_5100, n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107, y26, n_5108, n_5109, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115, n_5116, n_5117, n_5118, n_5119, n_5120, n_5121, n_5122, n_5123, n_5124, n_5125, n_5126, n_5127, n_5128, n_5129, n_5130, n_5131, n_5132, n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139, n_5140, n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147, n_5148, n_5149, n_5150, n_5151, n_5152, n_5153, n_5154, n_5155, n_5156, n_5157, n_5158, n_5159, n_5160, n_5161, n_5162, n_5163, n_5164, n_5165, n_5166, n_5167, n_5168, n_5169, n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5176, n_5177, n_5178, n_5179, n_5180, n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192, n_5193, n_5194, n_5195, n_5196, n_5197, n_5198, n_5199, n_5200, n_5201, n_5202, n_5203, n_5204, n_5205, n_5206, n_5207, n_5208, n_5209, n_5210, n_5211, n_5212, n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, n_5219, n_5220, n_5221, n_5222, n_5223, n_5224, n_5225, n_5226, n_5227, n_5228, n_5229, n_5230, n_5231, n_5232, n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240, n_5241, n_5242, n_5243, n_5244, n_5245, n_5246, n_5247, n_5248, n_5249, n_5250, n_5251, n_5252, n_5253, n_5254, n_5255, n_5256, n_5257, n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264, n_5265, n_5266, n_5267, n_5268, n_5269, n_5270, n_5271, n_5272, n_5273, n_5274, n_5275, n_5276, n_5277, n_5278, n_5279, n_5280, n_5281, n_5282, n_5283, n_5284, n_5285, n_5286, n_5287, n_5288, n_5289, n_5290, n_5291, n_5292, n_5293, n_5294, n_5295, n_5296, n_5297, n_5298, n_5299, n_5300, n_5301, n_5302, n_5303, n_5304, n_5305, n_5306, n_5307, n_5308, n_5309, n_5310, n_5311, n_5312, n_5313, n_5314, n_5315, n_5316, n_5317, n_5318, n_5319, n_5320, n_5321, n_5322, n_5323, n_5324, n_5325, n_5326, n_5327, n_5328, n_5329, n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, n_5336, n_5337, n_5338, n_5339, n_5340, n_5341, n_5342, n_5343, n_5344, n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5351, n_5352, n_5353, n_5354, n_5355, n_5356, n_5357, n_5358, n_5359, n_5360, n_5361, y25, n_5362, n_5363, n_5364, n_5365, n_5366, n_5367, n_5368, n_5369, n_5370, n_5371, n_5372, n_5373, n_5374, n_5375, n_5376, n_5377, n_5378, n_5379, n_5380, n_5381, n_5382, n_5383, n_5384, n_5385, n_5386, n_5387, n_5388, n_5389, n_5390, n_5391, n_5392, n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5399, n_5400, n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407, n_5408, n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415, n_5416, n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423, n_5424, n_5425, n_5426, n_5427, n_5428, n_5429, n_5430, n_5431, n_5432, n_5433, n_5434, n_5435, n_5436, n_5437, n_5438, n_5439, n_5440, n_5441, n_5442, n_5443, n_5444, n_5445, n_5446, n_5447, n_5448, n_5449, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456, n_5457, n_5458, n_5459, n_5460, n_5461, n_5462, n_5463, n_5464, n_5465, n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472, n_5473, n_5474, n_5475, n_5476, n_5477, n_5478, n_5479, n_5480, n_5481, n_5482, n_5483, n_5484, n_5485, n_5486, n_5487, n_5488, n_5489, n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, n_5496, n_5497, n_5498, n_5499, n_5500, n_5501, n_5502, n_5503, n_5504, n_5505, n_5506, n_5507, n_5508, n_5509, n_5510, n_5511, n_5512, n_5513, n_5514, n_5515, n_5516, n_5517, n_5518, n_5519, n_5520, n_5521, n_5522, n_5523, n_5524, n_5525, n_5526, n_5527, n_5528, n_5529, n_5530, n_5531, n_5532, n_5533, n_5534, n_5535, n_5536, n_5537, n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544, n_5545, n_5546, n_5547, n_5548, n_5549, n_5550, n_5551, n_5552, n_5553, n_5554, n_5555, n_5556, n_5557, n_5558, n_5559, n_5560, n_5561, n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568, n_5569, n_5570, n_5571, n_5572, n_5573, n_5574, n_5575, n_5576, n_5577, n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584, n_5585, n_5586, n_5587, n_5588, n_5589, n_5590, n_5591, n_5592, n_5593, n_5594, n_5595, n_5596, n_5597, n_5598, n_5599, n_5600, n_5601, n_5602, n_5603, n_5604, n_5605, n_5606, n_5607, n_5608, n_5609, y24, n_5610, n_5611, n_5612, n_5613, n_5614, n_5615, n_5616, n_5617, n_5618, n_5619, n_5620, n_5621, n_5622, n_5623, n_5624, n_5625, n_5626, n_5627, n_5628, n_5629, n_5630, n_5631, n_5632, n_5633, n_5634, n_5635, n_5636, n_5637, n_5638, n_5639, n_5640, n_5641, n_5642, n_5643, n_5644, n_5645, n_5646, n_5647, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653, n_5654, n_5655, n_5656, n_5657, n_5658, n_5659, n_5660, n_5661, n_5662, n_5663, n_5664, n_5665, n_5666, n_5667, n_5668, n_5669, n_5670, n_5671, n_5672, n_5673, n_5674, n_5675, n_5676, n_5677, n_5678, n_5679, n_5680, n_5681, n_5682, n_5683, n_5684, n_5685, n_5686, n_5687, n_5688, n_5689, n_5690, n_5691, n_5692, n_5693, n_5694, n_5695, n_5696, n_5697, n_5698, n_5699, n_5700, n_5701, n_5702, n_5703, n_5704, n_5705, n_5706, n_5707, n_5708, n_5709, n_5710, n_5711, n_5712, n_5713, n_5714, n_5715, n_5716, n_5717, n_5718, n_5719, n_5720, n_5721, n_5722, n_5723, n_5724, n_5725, n_5726, n_5727, n_5728, n_5729, n_5730, n_5731, n_5732, n_5733, n_5734, n_5735, n_5736, n_5737, n_5738, n_5739, n_5740, n_5741, n_5742, n_5743, n_5744, n_5745, n_5746, n_5747, n_5748, n_5749, n_5750, n_5751, n_5752, n_5753, n_5754, n_5755, n_5756, n_5757, n_5758, n_5759, n_5760, n_5761, n_5762, n_5763, n_5764, n_5765, n_5766, n_5767, n_5768, n_5769, n_5770, n_5771, n_5772, n_5773, n_5774, n_5775, n_5776, n_5777, n_5778, n_5779, n_5780, n_5781, n_5782, n_5783, n_5784, n_5785, n_5786, n_5787, n_5788, n_5789, n_5790, n_5791, n_5792, n_5793, n_5794, n_5795, n_5796, n_5797, n_5798, n_5799, n_5800, n_5801, n_5802, n_5803, n_5804, n_5805, n_5806, n_5807, n_5808, n_5809, n_5810, n_5811, n_5812, n_5813, n_5814, n_5815, n_5816, n_5817, n_5818, n_5819, n_5820, n_5821, n_5822, n_5823, n_5824, n_5825, n_5826, n_5827, n_5828, n_5829, n_5830, n_5831, n_5832, n_5833, n_5834, n_5835, n_5836, n_5837, n_5838, n_5839, n_5840, n_5841, n_5842, n_5843, n_5844, n_5845, n_5846, n_5847, n_5848, n_5849, n_5850, n_5851, n_5852, n_5853, n_5854, n_5855, n_5856, n_5857, n_5858, n_5859, n_5860, n_5861, n_5862, n_5863, n_5864, n_5865, n_5866, n_5867, n_5868, n_5869, n_5870, n_5871, n_5872, n_5873, n_5874, n_5875, n_5876, n_5877, n_5878, n_5879, n_5880, n_5881, y23, n_5882, n_5883, n_5884, n_5885, n_5886, n_5887, n_5888, n_5889, n_5890, n_5891, n_5892, n_5893, n_5894, n_5895, n_5896, n_5897, n_5898, n_5899, n_5900, n_5901, n_5902, n_5903, n_5904, n_5905, n_5906, n_5907, n_5908, n_5909, n_5910, n_5911, n_5912, n_5913, n_5914, n_5915, n_5916, n_5917, n_5918, n_5919, n_5920, n_5921, n_5922, n_5923, n_5924, n_5925, n_5926, n_5927, n_5928, n_5929, n_5930, n_5931, n_5932, n_5933, n_5934, n_5935, n_5936, n_5937, n_5938, n_5939, n_5940, n_5941, n_5942, n_5943, n_5944, n_5945, n_5946, n_5947, n_5948, n_5949, n_5950, n_5951, n_5952, n_5953, n_5954, n_5955, n_5956, n_5957, n_5958, n_5959, n_5960, n_5961, n_5962, n_5963, n_5964, n_5965, n_5966, n_5967, n_5968, n_5969, n_5970, n_5971, n_5972, n_5973, n_5974, n_5975, n_5976, n_5977, n_5978, n_5979, n_5980, n_5981, n_5982, n_5983, n_5984, n_5985, n_5986, n_5987, n_5988, n_5989, n_5990, n_5991, n_5992, n_5993, n_5994, n_5995, n_5996, n_5997, n_5998, n_5999, n_6000, n_6001, n_6002, n_6003, n_6004, n_6005, n_6006, n_6007, n_6008, n_6009, n_6010, n_6011, n_6012, n_6013, n_6014, n_6015, n_6016, n_6017, n_6018, n_6019, n_6020, n_6021, n_6022, n_6023, n_6024, n_6025, n_6026, n_6027, n_6028, n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, n_6035, n_6036, n_6037, n_6038, n_6039, n_6040, n_6041, n_6042, n_6043, n_6044, n_6045, n_6046, n_6047, n_6048, n_6049, n_6050, n_6051, n_6052, n_6053, n_6054, n_6055, n_6056, n_6057, n_6058, n_6059, n_6060, n_6061, n_6062, n_6063, n_6064, n_6065, n_6066, n_6067, n_6068, n_6069, n_6070, n_6071, n_6072, n_6073, n_6074, n_6075, n_6076, n_6077, n_6078, n_6079, n_6080, n_6081, n_6082, n_6083, n_6084, n_6085, n_6086, n_6087, n_6088, n_6089, n_6090, n_6091, n_6092, n_6093, n_6094, n_6095, n_6096, n_6097, n_6098, n_6099, n_6100, n_6101, n_6102, n_6103, n_6104, n_6105, n_6106, n_6107, n_6108, n_6109, n_6110, n_6111, n_6112, n_6113, n_6114, n_6115, n_6116, n_6117, n_6118, n_6119, n_6120, n_6121, n_6122, n_6123, n_6124, n_6125, n_6126, n_6127, n_6128, n_6129, n_6130, n_6131, n_6132, n_6133, n_6134, n_6135, n_6136, n_6137, n_6138, n_6139, n_6140, n_6141, n_6142, n_6143, n_6144, n_6145, n_6146, n_6147, n_6148, n_6149, n_6150, n_6151, n_6152, n_6153, n_6154, n_6155, n_6156, n_6157, n_6158, y22, n_6159, n_6160, n_6161, n_6162, n_6163, n_6164, n_6165, n_6166, n_6167, n_6168, n_6169, n_6170, n_6171, n_6172, n_6173, n_6174, n_6175, n_6176, n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183, n_6184, n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191, n_6192, n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199, n_6200, n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207, n_6208, n_6209, n_6210, n_6211, n_6212, n_6213, n_6214, n_6215, n_6216, n_6217, n_6218, n_6219, n_6220, n_6221, n_6222, n_6223, n_6224, n_6225, n_6226, n_6227, n_6228, n_6229, n_6230, n_6231, n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239, n_6240, n_6241, n_6242, n_6243, n_6244, n_6245, n_6246, n_6247, n_6248, n_6249, n_6250, n_6251, n_6252, n_6253, n_6254, n_6255, n_6256, n_6257, n_6258, n_6259, n_6260, n_6261, n_6262, n_6263, n_6264, n_6265, n_6266, n_6267, n_6268, n_6269, n_6270, n_6271, n_6272, n_6273, n_6274, n_6275, n_6276, n_6277, n_6278, n_6279, n_6280, n_6281, n_6282, n_6283, n_6284, n_6285, n_6286, n_6287, n_6288, n_6289, n_6290, n_6291, n_6292, n_6293, n_6294, n_6295, n_6296, n_6297, n_6298, n_6299, n_6300, n_6301, n_6302, n_6303, n_6304, n_6305, n_6306, n_6307, n_6308, n_6309, n_6310, n_6311, n_6312, n_6313, n_6314, n_6315, n_6316, n_6317, n_6318, n_6319, n_6320, n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, n_6327, n_6328, n_6329, n_6330, n_6331, n_6332, n_6333, n_6334, n_6335, n_6336, n_6337, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343, n_6344, n_6345, n_6346, n_6347, n_6348, n_6349, n_6350, n_6351, n_6352, n_6353, n_6354, n_6355, n_6356, n_6357, n_6358, n_6359, n_6360, n_6361, n_6362, n_6363, n_6364, n_6365, n_6366, n_6367, n_6368, n_6369, n_6370, n_6371, n_6372, n_6373, n_6374, n_6375, n_6376, n_6377, n_6378, n_6379, n_6380, n_6381, n_6382, n_6383, n_6384, n_6385, n_6386, n_6387, n_6388, n_6389, n_6390, n_6391, n_6392, n_6393, n_6394, n_6395, n_6396, n_6397, n_6398, n_6399, n_6400, n_6401, n_6402, n_6403, n_6404, n_6405, n_6406, n_6407, n_6408, n_6409, n_6410, n_6411, n_6412, n_6413, n_6414, n_6415, n_6416, n_6417, n_6418, n_6419, n_6420, n_6421, n_6422, n_6423, n_6424, n_6425, n_6426, n_6427, n_6428, n_6429, n_6430, n_6431, n_6432, n_6433, n_6434, n_6435, n_6436, n_6437, n_6438, n_6439, n_6440, n_6441, n_6442, n_6443, n_6444, n_6445, n_6446, n_6447, n_6448, n_6449, n_6450, n_6451, n_6452, n_6453, n_6454, n_6455, n_6456, n_6457, n_6458, n_6459, n_6460, n_6461, n_6462, n_6463, n_6464, y21, n_6465, n_6466, n_6467, n_6468, n_6469, n_6470, n_6471, n_6472, n_6473, n_6474, n_6475, n_6476, n_6477, n_6478, n_6479, n_6480, n_6481, n_6482, n_6483, n_6484, n_6485, n_6486, n_6487, n_6488, n_6489, n_6490, n_6491, n_6492, n_6493, n_6494, n_6495, n_6496, n_6497, n_6498, n_6499, n_6500, n_6501, n_6502, n_6503, n_6504, n_6505, n_6506, n_6507, n_6508, n_6509, n_6510, n_6511, n_6512, n_6513, n_6514, n_6515, n_6516, n_6517, n_6518, n_6519, n_6520, n_6521, n_6522, n_6523, n_6524, n_6525, n_6526, n_6527, n_6528, n_6529, n_6530, n_6531, n_6532, n_6533, n_6534, n_6535, n_6536, n_6537, n_6538, n_6539, n_6540, n_6541, n_6542, n_6543, n_6544, n_6545, n_6546, n_6547, n_6548, n_6549, n_6550, n_6551, n_6552, n_6553, n_6554, n_6555, n_6556, n_6557, n_6558, n_6559, n_6560, n_6561, n_6562, n_6563, n_6564, n_6565, n_6566, n_6567, n_6568, n_6569, n_6570, n_6571, n_6572, n_6573, n_6574, n_6575, n_6576, n_6577, n_6578, n_6579, n_6580, n_6581, n_6582, n_6583, n_6584, n_6585, n_6586, n_6587, n_6588, n_6589, n_6590, n_6591, n_6592, n_6593, n_6594, n_6595, n_6596, n_6597, n_6598, n_6599, n_6600, n_6601, n_6602, n_6603, n_6604, n_6605, n_6606, n_6607, n_6608, n_6609, n_6610, n_6611, n_6612, n_6613, n_6614, n_6615, n_6616, n_6617, n_6618, n_6619, n_6620, n_6621, n_6622, n_6623, n_6624, n_6625, n_6626, n_6627, n_6628, n_6629, n_6630, n_6631, n_6632, n_6633, n_6634, n_6635, n_6636, n_6637, n_6638, n_6639, n_6640, n_6641, n_6642, n_6643, n_6644, n_6645, n_6646, n_6647, n_6648, n_6649, n_6650, n_6651, n_6652, n_6653, n_6654, n_6655, n_6656, n_6657, n_6658, n_6659, n_6660, n_6661, n_6662, n_6663, n_6664, n_6665, n_6666, n_6667, n_6668, n_6669, n_6670, n_6671, n_6672, n_6673, n_6674, n_6675, n_6676, n_6677, n_6678, n_6679, n_6680, n_6681, n_6682, n_6683, n_6684, n_6685, n_6686, n_6687, n_6688, n_6689, n_6690, n_6691, n_6692, n_6693, n_6694, n_6695, n_6696, n_6697, n_6698, n_6699, n_6700, n_6701, n_6702, n_6703, n_6704, n_6705, n_6706, n_6707, n_6708, n_6709, n_6710, n_6711, n_6712, n_6713, n_6714, n_6715, n_6716, n_6717, n_6718, n_6719, n_6720, n_6721, n_6722, n_6723, n_6724, n_6725, n_6726, n_6727, n_6728, n_6729, n_6730, n_6731, n_6732, n_6733, n_6734, n_6735, n_6736, n_6737, n_6738, n_6739, n_6740, n_6741, n_6742, n_6743, n_6744, n_6745, n_6746, n_6747, n_6748, n_6749, n_6750, n_6751, n_6752, n_6753, n_6754, n_6755, n_6756, n_6757, n_6758, n_6759, y20, n_6760, n_6761, n_6762, n_6763, n_6764, n_6765, n_6766, n_6767, n_6768, n_6769, n_6770, n_6771, n_6772, n_6773, n_6774, n_6775, n_6776, n_6777, n_6778, n_6779, n_6780, n_6781, n_6782, n_6783, n_6784, n_6785, n_6786, n_6787, n_6788, n_6789, n_6790, n_6791, n_6792, n_6793, n_6794, n_6795, n_6796, n_6797, n_6798, n_6799, n_6800, n_6801, n_6802, n_6803, n_6804, n_6805, n_6806, n_6807, n_6808, n_6809, n_6810, n_6811, n_6812, n_6813, n_6814, n_6815, n_6816, n_6817, n_6818, n_6819, n_6820, n_6821, n_6822, n_6823, n_6824, n_6825, n_6826, n_6827, n_6828, n_6829, n_6830, n_6831, n_6832, n_6833, n_6834, n_6835, n_6836, n_6837, n_6838, n_6839, n_6840, n_6841, n_6842, n_6843, n_6844, n_6845, n_6846, n_6847, n_6848, n_6849, n_6850, n_6851, n_6852, n_6853, n_6854, n_6855, n_6856, n_6857, n_6858, n_6859, n_6860, n_6861, n_6862, n_6863, n_6864, n_6865, n_6866, n_6867, n_6868, n_6869, n_6870, n_6871, n_6872, n_6873, n_6874, n_6875, n_6876, n_6877, n_6878, n_6879, n_6880, n_6881, n_6882, n_6883, n_6884, n_6885, n_6886, n_6887, n_6888, n_6889, n_6890, n_6891, n_6892, n_6893, n_6894, n_6895, n_6896, n_6897, n_6898, n_6899, n_6900, n_6901, n_6902, n_6903, n_6904, n_6905, n_6906, n_6907, n_6908, n_6909, n_6910, n_6911, n_6912, n_6913, n_6914, n_6915, n_6916, n_6917, n_6918, n_6919, n_6920, n_6921, n_6922, n_6923, n_6924, n_6925, n_6926, n_6927, n_6928, n_6929, n_6930, n_6931, n_6932, n_6933, n_6934, n_6935, n_6936, n_6937, n_6938, n_6939, n_6940, n_6941, n_6942, n_6943, n_6944, n_6945, n_6946, n_6947, n_6948, n_6949, n_6950, n_6951, n_6952, n_6953, n_6954, n_6955, n_6956, n_6957, n_6958, n_6959, n_6960, n_6961, n_6962, n_6963, n_6964, n_6965, n_6966, n_6967, n_6968, n_6969, n_6970, n_6971, n_6972, n_6973, n_6974, n_6975, n_6976, n_6977, n_6978, n_6979, n_6980, n_6981, n_6982, n_6983, n_6984, n_6985, n_6986, n_6987, n_6988, n_6989, n_6990, n_6991, n_6992, n_6993, n_6994, n_6995, n_6996, n_6997, n_6998, n_6999, n_7000, n_7001, n_7002, n_7003, n_7004, n_7005, n_7006, n_7007, n_7008, n_7009, n_7010, n_7011, n_7012, n_7013, n_7014, n_7015, n_7016, n_7017, n_7018, n_7019, n_7020, n_7021, n_7022, n_7023, n_7024, n_7025, n_7026, n_7027, n_7028, n_7029, n_7030, n_7031, n_7032, n_7033, n_7034, n_7035, n_7036, n_7037, n_7038, n_7039, n_7040, n_7041, n_7042, n_7043, n_7044, n_7045, n_7046, n_7047, n_7048, n_7049, n_7050, n_7051, n_7052, y19, n_7053, n_7054, n_7055, n_7056, n_7057, n_7058, n_7059, n_7060, n_7061, n_7062, n_7063, n_7064, n_7065, n_7066, n_7067, n_7068, n_7069, n_7070, n_7071, n_7072, n_7073, n_7074, n_7075, n_7076, n_7077, n_7078, n_7079, n_7080, n_7081, n_7082, n_7083, n_7084, n_7085, n_7086, n_7087, n_7088, n_7089, n_7090, n_7091, n_7092, n_7093, n_7094, n_7095, n_7096, n_7097, n_7098, n_7099, n_7100, n_7101, n_7102, n_7103, n_7104, n_7105, n_7106, n_7107, n_7108, n_7109, n_7110, n_7111, n_7112, n_7113, n_7114, n_7115, n_7116, n_7117, n_7118, n_7119, n_7120, n_7121, n_7122, n_7123, n_7124, n_7125, n_7126, n_7127, n_7128, n_7129, n_7130, n_7131, n_7132, n_7133, n_7134, n_7135, n_7136, n_7137, n_7138, n_7139, n_7140, n_7141, n_7142, n_7143, n_7144, n_7145, n_7146, n_7147, n_7148, n_7149, n_7150, n_7151, n_7152, n_7153, n_7154, n_7155, n_7156, n_7157, n_7158, n_7159, n_7160, n_7161, n_7162, n_7163, n_7164, n_7165, n_7166, n_7167, n_7168, n_7169, n_7170, n_7171, n_7172, n_7173, n_7174, n_7175, n_7176, n_7177, n_7178, n_7179, n_7180, n_7181, n_7182, n_7183, n_7184, n_7185, n_7186, n_7187, n_7188, n_7189, n_7190, n_7191, n_7192, n_7193, n_7194, n_7195, n_7196, n_7197, n_7198, n_7199, n_7200, n_7201, n_7202, n_7203, n_7204, n_7205, n_7206, n_7207, n_7208, n_7209, n_7210, n_7211, n_7212, n_7213, n_7214, n_7215, n_7216, n_7217, n_7218, n_7219, n_7220, n_7221, n_7222, n_7223, n_7224, n_7225, n_7226, n_7227, n_7228, n_7229, n_7230, n_7231, n_7232, n_7233, n_7234, n_7235, n_7236, n_7237, n_7238, n_7239, n_7240, n_7241, n_7242, n_7243, n_7244, n_7245, n_7246, n_7247, n_7248, n_7249, n_7250, n_7251, n_7252, n_7253, n_7254, n_7255, n_7256, n_7257, n_7258, n_7259, n_7260, n_7261, n_7262, n_7263, n_7264, n_7265, n_7266, n_7267, n_7268, n_7269, n_7270, n_7271, n_7272, n_7273, n_7274, n_7275, n_7276, n_7277, n_7278, n_7279, n_7280, n_7281, n_7282, n_7283, n_7284, n_7285, n_7286, n_7287, n_7288, n_7289, n_7290, n_7291, n_7292, n_7293, n_7294, n_7295, n_7296, n_7297, n_7298, n_7299, n_7300, n_7301, n_7302, n_7303, n_7304, n_7305, n_7306, n_7307, n_7308, n_7309, n_7310, n_7311, n_7312, n_7313, n_7314, n_7315, n_7316, n_7317, n_7318, n_7319, n_7320, n_7321, n_7322, n_7323, n_7324, n_7325, n_7326, n_7327, n_7328, n_7329, n_7330, n_7331, n_7332, n_7333, n_7334, n_7335, n_7336, n_7337, n_7338, n_7339, n_7340, n_7341, n_7342, n_7343, n_7344, n_7345, n_7346, n_7347, n_7348, n_7349, n_7350, n_7351, n_7352, n_7353, n_7354, y18, n_7355, n_7356, n_7357, n_7358, n_7359, n_7360, n_7361, n_7362, n_7363, n_7364, n_7365, n_7366, n_7367, n_7368, n_7369, n_7370, n_7371, n_7372, n_7373, n_7374, n_7375, n_7376, n_7377, n_7378, n_7379, n_7380, n_7381, n_7382, n_7383, n_7384, n_7385, n_7386, n_7387, n_7388, n_7389, n_7390, n_7391, n_7392, n_7393, n_7394, n_7395, n_7396, n_7397, n_7398, n_7399, n_7400, n_7401, n_7402, n_7403, n_7404, n_7405, n_7406, n_7407, n_7408, n_7409, n_7410, n_7411, n_7412, n_7413, n_7414, n_7415, n_7416, n_7417, n_7418, n_7419, n_7420, n_7421, n_7422, n_7423, n_7424, n_7425, n_7426, n_7427, n_7428, n_7429, n_7430, n_7431, n_7432, n_7433, n_7434, n_7435, n_7436, n_7437, n_7438, n_7439, n_7440, n_7441, n_7442, n_7443, n_7444, n_7445, n_7446, n_7447, n_7448, n_7449, n_7450, n_7451, n_7452, n_7453, n_7454, n_7455, n_7456, n_7457, n_7458, n_7459, n_7460, n_7461, n_7462, n_7463, n_7464, n_7465, n_7466, n_7467, n_7468, n_7469, n_7470, n_7471, n_7472, n_7473, n_7474, n_7475, n_7476, n_7477, n_7478, n_7479, n_7480, n_7481, n_7482, n_7483, n_7484, n_7485, n_7486, n_7487, n_7488, n_7489, n_7490, n_7491, n_7492, n_7493, n_7494, n_7495, n_7496, n_7497, n_7498, n_7499, n_7500, n_7501, n_7502, n_7503, n_7504, n_7505, n_7506, n_7507, n_7508, n_7509, n_7510, n_7511, n_7512, n_7513, n_7514, n_7515, n_7516, n_7517, n_7518, n_7519, n_7520, n_7521, n_7522, n_7523, n_7524, n_7525, n_7526, n_7527, n_7528, n_7529, n_7530, n_7531, n_7532, n_7533, n_7534, n_7535, n_7536, n_7537, n_7538, n_7539, n_7540, n_7541, n_7542, n_7543, n_7544, n_7545, n_7546, n_7547, n_7548, n_7549, n_7550, n_7551, n_7552, n_7553, n_7554, n_7555, n_7556, n_7557, n_7558, n_7559, n_7560, n_7561, n_7562, n_7563, n_7564, n_7565, n_7566, n_7567, n_7568, n_7569, n_7570, n_7571, n_7572, n_7573, n_7574, n_7575, n_7576, n_7577, n_7578, n_7579, n_7580, n_7581, n_7582, n_7583, n_7584, n_7585, n_7586, n_7587, n_7588, n_7589, n_7590, n_7591, n_7592, n_7593, n_7594, n_7595, n_7596, n_7597, n_7598, n_7599, n_7600, n_7601, n_7602, n_7603, n_7604, n_7605, n_7606, n_7607, n_7608, n_7609, n_7610, n_7611, n_7612, n_7613, n_7614, n_7615, n_7616, n_7617, n_7618, n_7619, n_7620, n_7621, n_7622, n_7623, n_7624, n_7625, n_7626, n_7627, n_7628, n_7629, n_7630, n_7631, n_7632, n_7633, n_7634, n_7635, n_7636, n_7637, n_7638, n_7639, n_7640, n_7641, n_7642, n_7643, n_7644, n_7645, n_7646, n_7647, n_7648, n_7649, n_7650, n_7651, n_7652, n_7653, n_7654, n_7655, n_7656, n_7657, n_7658, n_7659, n_7660, n_7661, n_7662, n_7663, n_7664, n_7665, y17, n_7666, n_7667, n_7668, n_7669, n_7670, n_7671, n_7672, n_7673, n_7674, n_7675, n_7676, n_7677, n_7678, n_7679, n_7680, n_7681, n_7682, n_7683, n_7684, n_7685, n_7686, n_7687, n_7688, n_7689, n_7690, n_7691, n_7692, n_7693, n_7694, n_7695, n_7696, n_7697, n_7698, n_7699, n_7700, n_7701, n_7702, n_7703, n_7704, n_7705, n_7706, n_7707, n_7708, n_7709, n_7710, n_7711, n_7712, n_7713, n_7714, n_7715, n_7716, n_7717, n_7718, n_7719, n_7720, n_7721, n_7722, n_7723, n_7724, n_7725, n_7726, n_7727, n_7728, n_7729, n_7730, n_7731, n_7732, n_7733, n_7734, n_7735, n_7736, n_7737, n_7738, n_7739, n_7740, n_7741, n_7742, n_7743, n_7744, n_7745, n_7746, n_7747, n_7748, n_7749, n_7750, n_7751, n_7752, n_7753, n_7754, n_7755, n_7756, n_7757, n_7758, n_7759, n_7760, n_7761, n_7762, n_7763, n_7764, n_7765, n_7766, n_7767, n_7768, n_7769, n_7770, n_7771, n_7772, n_7773, n_7774, n_7775, n_7776, n_7777, n_7778, n_7779, n_7780, n_7781, n_7782, n_7783, n_7784, n_7785, n_7786, n_7787, n_7788, n_7789, n_7790, n_7791, n_7792, n_7793, n_7794, n_7795, n_7796, n_7797, n_7798, n_7799, n_7800, n_7801, n_7802, n_7803, n_7804, n_7805, n_7806, n_7807, n_7808, n_7809, n_7810, n_7811, n_7812, n_7813, n_7814, n_7815, n_7816, n_7817, n_7818, n_7819, n_7820, n_7821, n_7822, n_7823, n_7824, n_7825, n_7826, n_7827, n_7828, n_7829, n_7830, n_7831, n_7832, n_7833, n_7834, n_7835, n_7836, n_7837, n_7838, n_7839, n_7840, n_7841, n_7842, n_7843, n_7844, n_7845, n_7846, n_7847, n_7848, n_7849, n_7850, n_7851, n_7852, n_7853, n_7854, n_7855, n_7856, n_7857, n_7858, n_7859, n_7860, n_7861, n_7862, n_7863, n_7864, n_7865, n_7866, n_7867, n_7868, n_7869, n_7870, n_7871, n_7872, n_7873, n_7874, n_7875, n_7876, n_7877, n_7878, n_7879, n_7880, n_7881, n_7882, n_7883, n_7884, n_7885, n_7886, n_7887, n_7888, n_7889, n_7890, n_7891, n_7892, n_7893, n_7894, n_7895, n_7896, n_7897, n_7898, n_7899, n_7900, n_7901, n_7902, n_7903, n_7904, n_7905, n_7906, n_7907, n_7908, n_7909, n_7910, n_7911, n_7912, n_7913, n_7914, n_7915, n_7916, n_7917, n_7918, n_7919, n_7920, n_7921, n_7922, n_7923, n_7924, n_7925, n_7926, n_7927, n_7928, n_7929, n_7930, n_7931, n_7932, n_7933, n_7934, n_7935, n_7936, n_7937, n_7938, n_7939, n_7940, n_7941, n_7942, n_7943, n_7944, n_7945, n_7946, n_7947, n_7948, n_7949, n_7950, n_7951, n_7952, n_7953, n_7954, n_7955, n_7956, n_7957, n_7958, n_7959, n_7960, n_7961, n_7962, n_7963, n_7964, n_7965, n_7966, n_7967, n_7968, y16, n_7969, n_7970, n_7971, n_7972, n_7973, n_7974, n_7975, n_7976, n_7977, n_7978, n_7979, n_7980, n_7981, n_7982, n_7983, n_7984, n_7985, n_7986, n_7987, n_7988, n_7989, n_7990, n_7991, n_7992, n_7993, n_7994, n_7995, n_7996, n_7997, n_7998, n_7999, n_8000, n_8001, n_8002, n_8003, n_8004, n_8005, n_8006, n_8007, n_8008, n_8009, n_8010, n_8011, n_8012, n_8013, n_8014, n_8015, n_8016, n_8017, n_8018, n_8019, n_8020, n_8021, n_8022, n_8023, n_8024, n_8025, n_8026, n_8027, n_8028, n_8029, n_8030, n_8031, n_8032, n_8033, n_8034, n_8035, n_8036, n_8037, n_8038, n_8039, n_8040, n_8041, n_8042, n_8043, n_8044, n_8045, n_8046, n_8047, n_8048, n_8049, n_8050, n_8051, n_8052, n_8053, n_8054, n_8055, n_8056, n_8057, n_8058, n_8059, n_8060, n_8061, n_8062, n_8063, n_8064, n_8065, n_8066, n_8067, n_8068, n_8069, n_8070, n_8071, n_8072, n_8073, n_8074, n_8075, n_8076, n_8077, n_8078, n_8079, n_8080, n_8081, n_8082, n_8083, n_8084, n_8085, n_8086, n_8087, n_8088, n_8089, n_8090, n_8091, n_8092, n_8093, n_8094, n_8095, n_8096, n_8097, n_8098, n_8099, n_8100, n_8101, n_8102, n_8103, n_8104, n_8105, n_8106, n_8107, n_8108, n_8109, n_8110, n_8111, n_8112, n_8113, n_8114, n_8115, n_8116, n_8117, n_8118, n_8119, n_8120, n_8121, n_8122, n_8123, n_8124, n_8125, n_8126, n_8127, n_8128, n_8129, n_8130, n_8131, n_8132, n_8133, n_8134, n_8135, n_8136, n_8137, n_8138, n_8139, n_8140, n_8141, n_8142, n_8143, n_8144, n_8145, n_8146, n_8147, n_8148, n_8149, n_8150, n_8151, n_8152, n_8153, n_8154, n_8155, n_8156, n_8157, n_8158, n_8159, n_8160, n_8161, n_8162, n_8163, n_8164, n_8165, n_8166, n_8167, n_8168, n_8169, n_8170, n_8171, n_8172, n_8173, n_8174, n_8175, n_8176, n_8177, n_8178, n_8179, n_8180, n_8181, n_8182, n_8183, n_8184, n_8185, n_8186, n_8187, n_8188, n_8189, n_8190, n_8191, n_8192, n_8193, n_8194, n_8195, n_8196, n_8197, n_8198, n_8199, n_8200, n_8201, n_8202, n_8203, n_8204, n_8205, n_8206, n_8207, n_8208, n_8209, n_8210, n_8211, n_8212, n_8213, n_8214, n_8215, n_8216, n_8217, n_8218, n_8219, n_8220, n_8221, n_8222, n_8223, n_8224, n_8225, n_8226, n_8227, n_8228, n_8229, n_8230, n_8231, n_8232, n_8233, n_8234, n_8235, n_8236, n_8237, n_8238, n_8239, n_8240, n_8241, n_8242, n_8243, n_8244, n_8245, n_8246, n_8247, n_8248, n_8249, n_8250, n_8251, n_8252, n_8253, n_8254, n_8255, n_8256, n_8257, n_8258, n_8259, n_8260, n_8261, n_8262, n_8263, n_8264, n_8265, n_8266, n_8267, n_8268, n_8269, n_8270, n_8271, n_8272, n_8273, n_8274, n_8275, n_8276, n_8277, n_8278, n_8279, n_8280, n_8281, n_8282, n_8283, n_8284, n_8285, n_8286, n_8287, n_8288, n_8289, n_8290, n_8291, y15, n_8292, n_8293, n_8294, n_8295, n_8296, n_8297, n_8298, n_8299, n_8300, n_8301, n_8302, n_8303, n_8304, n_8305, n_8306, n_8307, n_8308, n_8309, n_8310, n_8311, n_8312, n_8313, n_8314, n_8315, n_8316, n_8317, n_8318, n_8319, n_8320, n_8321, n_8322, n_8323, n_8324, n_8325, n_8326, n_8327, n_8328, n_8329, n_8330, n_8331, n_8332, n_8333, n_8334, n_8335, n_8336, n_8337, n_8338, n_8339, n_8340, n_8341, n_8342, n_8343, n_8344, n_8345, n_8346, n_8347, n_8348, n_8349, n_8350, n_8351, n_8352, n_8353, n_8354, n_8355, n_8356, n_8357, n_8358, n_8359, n_8360, n_8361, n_8362, n_8363, n_8364, n_8365, n_8366, n_8367, n_8368, n_8369, n_8370, n_8371, n_8372, n_8373, n_8374, n_8375, n_8376, n_8377, n_8378, n_8379, n_8380, n_8381, n_8382, n_8383, n_8384, n_8385, n_8386, n_8387, n_8388, n_8389, n_8390, n_8391, n_8392, n_8393, n_8394, n_8395, n_8396, n_8397, n_8398, n_8399, n_8400, n_8401, n_8402, n_8403, n_8404, n_8405, n_8406, n_8407, n_8408, n_8409, n_8410, n_8411, n_8412, n_8413, n_8414, n_8415, n_8416, n_8417, n_8418, n_8419, n_8420, n_8421, n_8422, n_8423, n_8424, n_8425, n_8426, n_8427, n_8428, n_8429, n_8430, n_8431, n_8432, n_8433, n_8434, n_8435, n_8436, n_8437, n_8438, n_8439, n_8440, n_8441, n_8442, n_8443, n_8444, n_8445, n_8446, n_8447, n_8448, n_8449, n_8450, n_8451, n_8452, n_8453, n_8454, n_8455, n_8456, n_8457, n_8458, n_8459, n_8460, n_8461, n_8462, n_8463, n_8464, n_8465, n_8466, n_8467, n_8468, n_8469, n_8470, n_8471, n_8472, n_8473, n_8474, n_8475, n_8476, n_8477, n_8478, n_8479, n_8480, n_8481, n_8482, n_8483, n_8484, n_8485, n_8486, n_8487, n_8488, n_8489, n_8490, n_8491, n_8492, n_8493, n_8494, n_8495, n_8496, n_8497, n_8498, n_8499, n_8500, n_8501, n_8502, n_8503, n_8504, n_8505, n_8506, n_8507, n_8508, n_8509, n_8510, n_8511, n_8512, n_8513, n_8514, n_8515, n_8516, n_8517, n_8518, n_8519, n_8520, n_8521, n_8522, n_8523, n_8524, n_8525, n_8526, n_8527, n_8528, n_8529, n_8530, n_8531, n_8532, n_8533, n_8534, n_8535, n_8536, n_8537, n_8538, n_8539, n_8540, n_8541, n_8542, n_8543, n_8544, n_8545, n_8546, n_8547, n_8548, n_8549, n_8550, n_8551, n_8552, n_8553, n_8554, n_8555, n_8556, n_8557, n_8558, n_8559, n_8560, n_8561, n_8562, n_8563, n_8564, n_8565, n_8566, n_8567, n_8568, n_8569, n_8570, n_8571, n_8572, n_8573, n_8574, n_8575, n_8576, n_8577, n_8578, n_8579, n_8580, n_8581, n_8582, n_8583, n_8584, n_8585, n_8586, n_8587, n_8588, n_8589, n_8590, n_8591, n_8592, n_8593, n_8594, n_8595, n_8596, n_8597, n_8598, n_8599, n_8600, n_8601, n_8602, n_8603, n_8604, n_8605, n_8606, n_8607, n_8608, n_8609, n_8610, n_8611, n_8612, n_8613, n_8614, n_8615, n_8616, n_8617, n_8618, n_8619, n_8620, n_8621, n_8622, n_8623, n_8624, n_8625, n_8626, y14, n_8627, n_8628, n_8629, n_8630, n_8631, n_8632, n_8633, n_8634, n_8635, n_8636, n_8637, n_8638, n_8639, n_8640, n_8641, n_8642, n_8643, n_8644, n_8645, n_8646, n_8647, n_8648, n_8649, n_8650, n_8651, n_8652, n_8653, n_8654, n_8655, n_8656, n_8657, n_8658, n_8659, n_8660, n_8661, n_8662, n_8663, n_8664, n_8665, n_8666, n_8667, n_8668, n_8669, n_8670, n_8671, n_8672, n_8673, n_8674, n_8675, n_8676, n_8677, n_8678, n_8679, n_8680, n_8681, n_8682, n_8683, n_8684, n_8685, n_8686, n_8687, n_8688, n_8689, n_8690, n_8691, n_8692, n_8693, n_8694, n_8695, n_8696, n_8697, n_8698, n_8699, n_8700, n_8701, n_8702, n_8703, n_8704, n_8705, n_8706, n_8707, n_8708, n_8709, n_8710, n_8711, n_8712, n_8713, n_8714, n_8715, n_8716, n_8717, n_8718, n_8719, n_8720, n_8721, n_8722, n_8723, n_8724, n_8725, n_8726, n_8727, n_8728, n_8729, n_8730, n_8731, n_8732, n_8733, n_8734, n_8735, n_8736, n_8737, n_8738, n_8739, n_8740, n_8741, n_8742, n_8743, n_8744, n_8745, n_8746, n_8747, n_8748, n_8749, n_8750, n_8751, n_8752, n_8753, n_8754, n_8755, n_8756, n_8757, n_8758, n_8759, n_8760, n_8761, n_8762, n_8763, n_8764, n_8765, n_8766, n_8767, n_8768, n_8769, n_8770, n_8771, n_8772, n_8773, n_8774, n_8775, n_8776, n_8777, n_8778, n_8779, n_8780, n_8781, n_8782, n_8783, n_8784, n_8785, n_8786, n_8787, n_8788, n_8789, n_8790, n_8791, n_8792, n_8793, n_8794, n_8795, n_8796, n_8797, n_8798, n_8799, n_8800, n_8801, n_8802, n_8803, n_8804, n_8805, n_8806, n_8807, n_8808, n_8809, n_8810, n_8811, n_8812, n_8813, n_8814, n_8815, n_8816, n_8817, n_8818, n_8819, n_8820, n_8821, n_8822, n_8823, n_8824, n_8825, n_8826, n_8827, n_8828, n_8829, n_8830, n_8831, n_8832, n_8833, n_8834, n_8835, n_8836, n_8837, n_8838, n_8839, n_8840, n_8841, n_8842, n_8843, n_8844, n_8845, n_8846, n_8847, n_8848, n_8849, n_8850, n_8851, n_8852, n_8853, n_8854, n_8855, n_8856, n_8857, n_8858, n_8859, n_8860, n_8861, n_8862, n_8863, n_8864, n_8865, n_8866, n_8867, n_8868, n_8869, n_8870, n_8871, n_8872, n_8873, n_8874, n_8875, n_8876, n_8877, n_8878, n_8879, n_8880, n_8881, n_8882, n_8883, n_8884, n_8885, n_8886, n_8887, n_8888, n_8889, n_8890, n_8891, n_8892, n_8893, n_8894, n_8895, n_8896, n_8897, n_8898, n_8899, n_8900, n_8901, n_8902, n_8903, n_8904, n_8905, n_8906, n_8907, n_8908, n_8909, n_8910, n_8911, n_8912, n_8913, n_8914, n_8915, n_8916, n_8917, n_8918, n_8919, n_8920, n_8921, n_8922, n_8923, n_8924, n_8925, n_8926, n_8927, n_8928, n_8929, n_8930, n_8931, n_8932, n_8933, n_8934, n_8935, n_8936, n_8937, n_8938, n_8939, n_8940, n_8941, n_8942, n_8943, n_8944, n_8945, n_8946, n_8947, n_8948, n_8949, n_8950, n_8951, n_8952, n_8953, n_8954, n_8955, n_8956, n_8957, n_8958, n_8959, n_8960, n_8961, n_8962, y13, n_8963, n_8964, n_8965, n_8966, n_8967, n_8968, n_8969, n_8970, n_8971, n_8972, n_8973, n_8974, n_8975, n_8976, n_8977, n_8978, n_8979, n_8980, n_8981, n_8982, n_8983, n_8984, n_8985, n_8986, n_8987, n_8988, n_8989, n_8990, n_8991, n_8992, n_8993, n_8994, n_8995, n_8996, n_8997, n_8998, n_8999, n_9000, n_9001, n_9002, n_9003, n_9004, n_9005, n_9006, n_9007, n_9008, n_9009, n_9010, n_9011, n_9012, n_9013, n_9014, n_9015, n_9016, n_9017, n_9018, n_9019, n_9020, n_9021, n_9022, n_9023, n_9024, n_9025, n_9026, n_9027, n_9028, n_9029, n_9030, n_9031, n_9032, n_9033, n_9034, n_9035, n_9036, n_9037, n_9038, n_9039, n_9040, n_9041, n_9042, n_9043, n_9044, n_9045, n_9046, n_9047, n_9048, n_9049, n_9050, n_9051, n_9052, n_9053, n_9054, n_9055, n_9056, n_9057, n_9058, n_9059, n_9060, n_9061, n_9062, n_9063, n_9064, n_9065, n_9066, n_9067, n_9068, n_9069, n_9070, n_9071, n_9072, n_9073, n_9074, n_9075, n_9076, n_9077, n_9078, n_9079, n_9080, n_9081, n_9082, n_9083, n_9084, n_9085, n_9086, n_9087, n_9088, n_9089, n_9090, n_9091, n_9092, n_9093, n_9094, n_9095, n_9096, n_9097, n_9098, n_9099, n_9100, n_9101, n_9102, n_9103, n_9104, n_9105, n_9106, n_9107, n_9108, n_9109, n_9110, n_9111, n_9112, n_9113, n_9114, n_9115, n_9116, n_9117, n_9118, n_9119, n_9120, n_9121, n_9122, n_9123, n_9124, n_9125, n_9126, n_9127, n_9128, n_9129, n_9130, n_9131, n_9132, n_9133, n_9134, n_9135, n_9136, n_9137, n_9138, n_9139, n_9140, n_9141, n_9142, n_9143, n_9144, n_9145, n_9146, n_9147, n_9148, n_9149, n_9150, n_9151, n_9152, n_9153, n_9154, n_9155, n_9156, n_9157, n_9158, n_9159, n_9160, n_9161, n_9162, n_9163, n_9164, n_9165, n_9166, n_9167, n_9168, n_9169, n_9170, n_9171, n_9172, n_9173, n_9174, n_9175, n_9176, n_9177, n_9178, n_9179, n_9180, n_9181, n_9182, n_9183, n_9184, n_9185, n_9186, n_9187, n_9188, n_9189, n_9190, n_9191, n_9192, n_9193, n_9194, n_9195, n_9196, n_9197, n_9198, n_9199, n_9200, n_9201, n_9202, n_9203, n_9204, n_9205, n_9206, n_9207, n_9208, n_9209, n_9210, n_9211, n_9212, n_9213, n_9214, n_9215, n_9216, n_9217, n_9218, n_9219, n_9220, n_9221, n_9222, n_9223, n_9224, n_9225, n_9226, n_9227, n_9228, n_9229, n_9230, n_9231, n_9232, n_9233, n_9234, n_9235, n_9236, n_9237, n_9238, n_9239, n_9240, n_9241, n_9242, n_9243, n_9244, n_9245, n_9246, n_9247, n_9248, n_9249, n_9250, n_9251, n_9252, n_9253, n_9254, n_9255, n_9256, n_9257, n_9258, n_9259, n_9260, n_9261, n_9262, n_9263, n_9264, n_9265, n_9266, n_9267, n_9268, n_9269, n_9270, n_9271, n_9272, n_9273, n_9274, n_9275, n_9276, n_9277, n_9278, n_9279, n_9280, n_9281, n_9282, n_9283, n_9284, n_9285, n_9286, n_9287, n_9288, n_9289, n_9290, n_9291, n_9292, n_9293, y12, n_9294, n_9295, n_9296, n_9297, n_9298, n_9299, n_9300, n_9301, n_9302, n_9303, n_9304, n_9305, n_9306, n_9307, n_9308, n_9309, n_9310, n_9311, n_9312, n_9313, n_9314, n_9315, n_9316, n_9317, n_9318, n_9319, n_9320, n_9321, n_9322, n_9323, n_9324, n_9325, n_9326, n_9327, n_9328, n_9329, n_9330, n_9331, n_9332, n_9333, n_9334, n_9335, n_9336, n_9337, n_9338, n_9339, n_9340, n_9341, n_9342, n_9343, n_9344, n_9345, n_9346, n_9347, n_9348, n_9349, n_9350, n_9351, n_9352, n_9353, n_9354, n_9355, n_9356, n_9357, n_9358, n_9359, n_9360, n_9361, n_9362, n_9363, n_9364, n_9365, n_9366, n_9367, n_9368, n_9369, n_9370, n_9371, n_9372, n_9373, n_9374, n_9375, n_9376, n_9377, n_9378, n_9379, n_9380, n_9381, n_9382, n_9383, n_9384, n_9385, n_9386, n_9387, n_9388, n_9389, n_9390, n_9391, n_9392, n_9393, n_9394, n_9395, n_9396, n_9397, n_9398, n_9399, n_9400, n_9401, n_9402, n_9403, n_9404, n_9405, n_9406, n_9407, n_9408, n_9409, n_9410, n_9411, n_9412, n_9413, n_9414, n_9415, n_9416, n_9417, n_9418, n_9419, n_9420, n_9421, n_9422, n_9423, n_9424, n_9425, n_9426, n_9427, n_9428, n_9429, n_9430, n_9431, n_9432, n_9433, n_9434, n_9435, n_9436, n_9437, n_9438, n_9439, n_9440, n_9441, n_9442, n_9443, n_9444, n_9445, n_9446, n_9447, n_9448, n_9449, n_9450, n_9451, n_9452, n_9453, n_9454, n_9455, n_9456, n_9457, n_9458, n_9459, n_9460, n_9461, n_9462, n_9463, n_9464, n_9465, n_9466, n_9467, n_9468, n_9469, n_9470, n_9471, n_9472, n_9473, n_9474, n_9475, n_9476, n_9477, n_9478, n_9479, n_9480, n_9481, n_9482, n_9483, n_9484, n_9485, n_9486, n_9487, n_9488, n_9489, n_9490, n_9491, n_9492, n_9493, n_9494, n_9495, n_9496, n_9497, n_9498, n_9499, n_9500, n_9501, n_9502, n_9503, n_9504, n_9505, n_9506, n_9507, n_9508, n_9509, n_9510, n_9511, n_9512, n_9513, n_9514, n_9515, n_9516, n_9517, n_9518, n_9519, n_9520, n_9521, n_9522, n_9523, n_9524, n_9525, n_9526, n_9527, n_9528, n_9529, n_9530, n_9531, n_9532, n_9533, n_9534, n_9535, n_9536, n_9537, n_9538, n_9539, n_9540, n_9541, n_9542, n_9543, n_9544, n_9545, n_9546, n_9547, n_9548, n_9549, n_9550, n_9551, n_9552, n_9553, n_9554, n_9555, n_9556, n_9557, n_9558, n_9559, n_9560, n_9561, n_9562, n_9563, n_9564, n_9565, n_9566, n_9567, n_9568, n_9569, n_9570, n_9571, n_9572, n_9573, n_9574, n_9575, n_9576, n_9577, n_9578, n_9579, n_9580, n_9581, n_9582, n_9583, n_9584, n_9585, n_9586, n_9587, n_9588, n_9589, n_9590, n_9591, n_9592, n_9593, n_9594, n_9595, n_9596, n_9597, n_9598, n_9599, n_9600, n_9601, n_9602, n_9603, n_9604, n_9605, n_9606, n_9607, n_9608, n_9609, n_9610, n_9611, n_9612, n_9613, n_9614, n_9615, n_9616, n_9617, n_9618, n_9619, n_9620, n_9621, n_9622, n_9623, n_9624, n_9625, n_9626, n_9627, n_9628, n_9629, n_9630, n_9631, n_9632, n_9633, n_9634, n_9635, n_9636, n_9637, n_9638, n_9639, n_9640, y11, n_9641, n_9642, n_9643, n_9644, n_9645, n_9646, n_9647, n_9648, n_9649, n_9650, n_9651, n_9652, n_9653, n_9654, n_9655, n_9656, n_9657, n_9658, n_9659, n_9660, n_9661, n_9662, n_9663, n_9664, n_9665, n_9666, n_9667, n_9668, n_9669, n_9670, n_9671, n_9672, n_9673, n_9674, n_9675, n_9676, n_9677, n_9678, n_9679, n_9680, n_9681, n_9682, n_9683, n_9684, n_9685, n_9686, n_9687, n_9688, n_9689, n_9690, n_9691, n_9692, n_9693, n_9694, n_9695, n_9696, n_9697, n_9698, n_9699, n_9700, n_9701, n_9702, n_9703, n_9704, n_9705, n_9706, n_9707, n_9708, n_9709, n_9710, n_9711, n_9712, n_9713, n_9714, n_9715, n_9716, n_9717, n_9718, n_9719, n_9720, n_9721, n_9722, n_9723, n_9724, n_9725, n_9726, n_9727, n_9728, n_9729, n_9730, n_9731, n_9732, n_9733, n_9734, n_9735, n_9736, n_9737, n_9738, n_9739, n_9740, n_9741, n_9742, n_9743, n_9744, n_9745, n_9746, n_9747, n_9748, n_9749, n_9750, n_9751, n_9752, n_9753, n_9754, n_9755, n_9756, n_9757, n_9758, n_9759, n_9760, n_9761, n_9762, n_9763, n_9764, n_9765, n_9766, n_9767, n_9768, n_9769, n_9770, n_9771, n_9772, n_9773, n_9774, n_9775, n_9776, n_9777, n_9778, n_9779, n_9780, n_9781, n_9782, n_9783, n_9784, n_9785, n_9786, n_9787, n_9788, n_9789, n_9790, n_9791, n_9792, n_9793, n_9794, n_9795, n_9796, n_9797, n_9798, n_9799, n_9800, n_9801, n_9802, n_9803, n_9804, n_9805, n_9806, n_9807, n_9808, n_9809, n_9810, n_9811, n_9812, n_9813, n_9814, n_9815, n_9816, n_9817, n_9818, n_9819, n_9820, n_9821, n_9822, n_9823, n_9824, n_9825, n_9826, n_9827, n_9828, n_9829, n_9830, n_9831, n_9832, n_9833, n_9834, n_9835, n_9836, n_9837, n_9838, n_9839, n_9840, n_9841, n_9842, n_9843, n_9844, n_9845, n_9846, n_9847, n_9848, n_9849, n_9850, n_9851, n_9852, n_9853, n_9854, n_9855, n_9856, n_9857, n_9858, n_9859, n_9860, n_9861, n_9862, n_9863, n_9864, n_9865, n_9866, n_9867, n_9868, n_9869, n_9870, n_9871, n_9872, n_9873, n_9874, n_9875, n_9876, n_9877, n_9878, n_9879, n_9880, n_9881, n_9882, n_9883, n_9884, n_9885, n_9886, n_9887, n_9888, n_9889, n_9890, n_9891, n_9892, n_9893, n_9894, n_9895, n_9896, n_9897, n_9898, n_9899, n_9900, n_9901, n_9902, n_9903, n_9904, n_9905, n_9906, n_9907, n_9908, n_9909, n_9910, n_9911, n_9912, n_9913, n_9914, n_9915, n_9916, n_9917, n_9918, n_9919, n_9920, n_9921, n_9922, n_9923, n_9924, n_9925, n_9926, n_9927, n_9928, n_9929, n_9930, n_9931, n_9932, n_9933, n_9934, n_9935, n_9936, n_9937, n_9938, n_9939, n_9940, n_9941, n_9942, n_9943, n_9944, n_9945, n_9946, n_9947, n_9948, n_9949, n_9950, n_9951, n_9952, n_9953, n_9954, n_9955, n_9956, n_9957, n_9958, n_9959, n_9960, n_9961, n_9962, n_9963, n_9964, n_9965, n_9966, n_9967, n_9968, n_9969, n_9970, n_9971, n_9972, n_9973, n_9974, n_9975, n_9976, n_9977, n_9978, n_9979, n_9980, n_9981, n_9982, n_9983, n_9984, n_9985, n_9986, n_9987, n_9988, n_9989, n_9990, n_9991, n_9992, n_9993, y10, n_9994, n_9995, n_9996, n_9997, n_9998, n_9999, n_10000, n_10001, n_10002, n_10003, n_10004, n_10005, n_10006, n_10007, n_10008, n_10009, n_10010, n_10011, n_10012, n_10013, n_10014, n_10015, n_10016, n_10017, n_10018, n_10019, n_10020, n_10021, n_10022, n_10023, n_10024, n_10025, n_10026, n_10027, n_10028, n_10029, n_10030, n_10031, n_10032, n_10033, n_10034, n_10035, n_10036, n_10037, n_10038, n_10039, n_10040, n_10041, n_10042, n_10043, n_10044, n_10045, n_10046, n_10047, n_10048, n_10049, n_10050, n_10051, n_10052, n_10053, n_10054, n_10055, n_10056, n_10057, n_10058, n_10059, n_10060, n_10061, n_10062, n_10063, n_10064, n_10065, n_10066, n_10067, n_10068, n_10069, n_10070, n_10071, n_10072, n_10073, n_10074, n_10075, n_10076, n_10077, n_10078, n_10079, n_10080, n_10081, n_10082, n_10083, n_10084, n_10085, n_10086, n_10087, n_10088, n_10089, n_10090, n_10091, n_10092, n_10093, n_10094, n_10095, n_10096, n_10097, n_10098, n_10099, n_10100, n_10101, n_10102, n_10103, n_10104, n_10105, n_10106, n_10107, n_10108, n_10109, n_10110, n_10111, n_10112, n_10113, n_10114, n_10115, n_10116, n_10117, n_10118, n_10119, n_10120, n_10121, n_10122, n_10123, n_10124, n_10125, n_10126, n_10127, n_10128, n_10129, n_10130, n_10131, n_10132, n_10133, n_10134, n_10135, n_10136, n_10137, n_10138, n_10139, n_10140, n_10141, n_10142, n_10143, n_10144, n_10145, n_10146, n_10147, n_10148, n_10149, n_10150, n_10151, n_10152, n_10153, n_10154, n_10155, n_10156, n_10157, n_10158, n_10159, n_10160, n_10161, n_10162, n_10163, n_10164, n_10165, n_10166, n_10167, n_10168, n_10169, n_10170, n_10171, n_10172, n_10173, n_10174, n_10175, n_10176, n_10177, n_10178, n_10179, n_10180, n_10181, n_10182, n_10183, n_10184, n_10185, n_10186, n_10187, n_10188, n_10189, n_10190, n_10191, n_10192, n_10193, n_10194, n_10195, n_10196, n_10197, n_10198, n_10199, n_10200, n_10201, n_10202, n_10203, n_10204, n_10205, n_10206, n_10207, n_10208, n_10209, n_10210, n_10211, n_10212, n_10213, n_10214, n_10215, n_10216, n_10217, n_10218, n_10219, n_10220, n_10221, n_10222, n_10223, n_10224, n_10225, n_10226, n_10227, n_10228, n_10229, n_10230, n_10231, n_10232, n_10233, n_10234, n_10235, n_10236, n_10237, n_10238, n_10239, n_10240, n_10241, n_10242, n_10243, n_10244, n_10245, n_10246, n_10247, n_10248, n_10249, n_10250, n_10251, n_10252, n_10253, n_10254, n_10255, n_10256, n_10257, n_10258, n_10259, n_10260, n_10261, n_10262, n_10263, n_10264, n_10265, n_10266, n_10267, n_10268, n_10269, n_10270, n_10271, n_10272, n_10273, n_10274, n_10275, n_10276, n_10277, n_10278, n_10279, n_10280, n_10281, n_10282, n_10283, n_10284, n_10285, n_10286, n_10287, n_10288, n_10289, n_10290, n_10291, n_10292, n_10293, n_10294, n_10295, n_10296, n_10297, n_10298, n_10299, n_10300, n_10301, n_10302, n_10303, n_10304, n_10305, n_10306, n_10307, n_10308, n_10309, n_10310, n_10311, n_10312, n_10313, n_10314, n_10315, n_10316, n_10317, n_10318, n_10319, n_10320, n_10321, n_10322, n_10323, n_10324, n_10325, n_10326, n_10327, n_10328, n_10329, n_10330, n_10331, n_10332, n_10333, n_10334, n_10335, n_10336, n_10337, n_10338, n_10339, n_10340, n_10341, n_10342, n_10343, n_10344, n_10345, n_10346, n_10347, n_10348, n_10349, n_10350, n_10351, n_10352, n_10353, n_10354, n_10355, n_10356, n_10357, n_10358, n_10359, n_10360, n_10361, n_10362, n_10363, n_10364, n_10365, n_10366, n_10367, n_10368, n_10369, n_10370, n_10371, n_10372, n_10373, n_10374, y9, n_10375, n_10376, n_10377, n_10378, n_10379, n_10380, n_10381, n_10382, n_10383, n_10384, n_10385, n_10386, n_10387, n_10388, n_10389, n_10390, n_10391, n_10392, n_10393, n_10394, n_10395, n_10396, n_10397, n_10398, n_10399, n_10400, n_10401, n_10402, n_10403, n_10404, n_10405, n_10406, n_10407, n_10408, n_10409, n_10410, n_10411, n_10412, n_10413, n_10414, n_10415, n_10416, n_10417, n_10418, n_10419, n_10420, n_10421, n_10422, n_10423, n_10424, n_10425, n_10426, n_10427, n_10428, n_10429, n_10430, n_10431, n_10432, n_10433, n_10434, n_10435, n_10436, n_10437, n_10438, n_10439, n_10440, n_10441, n_10442, n_10443, n_10444, n_10445, n_10446, n_10447, n_10448, n_10449, n_10450, n_10451, n_10452, n_10453, n_10454, n_10455, n_10456, n_10457, n_10458, n_10459, n_10460, n_10461, n_10462, n_10463, n_10464, n_10465, n_10466, n_10467, n_10468, n_10469, n_10470, n_10471, n_10472, n_10473, n_10474, n_10475, n_10476, n_10477, n_10478, n_10479, n_10480, n_10481, n_10482, n_10483, n_10484, n_10485, n_10486, n_10487, n_10488, n_10489, n_10490, n_10491, n_10492, n_10493, n_10494, n_10495, n_10496, n_10497, n_10498, n_10499, n_10500, n_10501, n_10502, n_10503, n_10504, n_10505, n_10506, n_10507, n_10508, n_10509, n_10510, n_10511, n_10512, n_10513, n_10514, n_10515, n_10516, n_10517, n_10518, n_10519, n_10520, n_10521, n_10522, n_10523, n_10524, n_10525, n_10526, n_10527, n_10528, n_10529, n_10530, n_10531, n_10532, n_10533, n_10534, n_10535, n_10536, n_10537, n_10538, n_10539, n_10540, n_10541, n_10542, n_10543, n_10544, n_10545, n_10546, n_10547, n_10548, n_10549, n_10550, n_10551, n_10552, n_10553, n_10554, n_10555, n_10556, n_10557, n_10558, n_10559, n_10560, n_10561, n_10562, n_10563, n_10564, n_10565, n_10566, n_10567, n_10568, n_10569, n_10570, n_10571, n_10572, n_10573, n_10574, n_10575, n_10576, n_10577, n_10578, n_10579, n_10580, n_10581, n_10582, n_10583, n_10584, n_10585, n_10586, n_10587, n_10588, n_10589, n_10590, n_10591, n_10592, n_10593, n_10594, n_10595, n_10596, n_10597, n_10598, n_10599, n_10600, n_10601, n_10602, n_10603, n_10604, n_10605, n_10606, n_10607, n_10608, n_10609, n_10610, n_10611, n_10612, n_10613, n_10614, n_10615, n_10616, n_10617, n_10618, n_10619, n_10620, n_10621, n_10622, n_10623, n_10624, n_10625, n_10626, n_10627, n_10628, n_10629, n_10630, n_10631, n_10632, n_10633, n_10634, n_10635, n_10636, n_10637, n_10638, n_10639, n_10640, n_10641, n_10642, n_10643, n_10644, n_10645, n_10646, n_10647, n_10648, n_10649, n_10650, n_10651, n_10652, n_10653, n_10654, n_10655, n_10656, n_10657, n_10658, n_10659, n_10660, n_10661, n_10662, n_10663, n_10664, n_10665, n_10666, n_10667, n_10668, n_10669, n_10670, n_10671, n_10672, n_10673, n_10674, n_10675, n_10676, n_10677, n_10678, n_10679, n_10680, n_10681, n_10682, n_10683, n_10684, n_10685, n_10686, n_10687, n_10688, n_10689, n_10690, n_10691, n_10692, n_10693, n_10694, n_10695, n_10696, n_10697, n_10698, n_10699, n_10700, n_10701, n_10702, n_10703, n_10704, n_10705, n_10706, n_10707, n_10708, n_10709, n_10710, n_10711, n_10712, n_10713, n_10714, n_10715, n_10716, n_10717, n_10718, n_10719, n_10720, n_10721, n_10722, n_10723, n_10724, n_10725, n_10726, n_10727, n_10728, n_10729, n_10730, y8, n_10731, n_10732, n_10733, n_10734, n_10735, n_10736, n_10737, n_10738, n_10739, n_10740, n_10741, n_10742, n_10743, n_10744, n_10745, n_10746, n_10747, n_10748, n_10749, n_10750, n_10751, n_10752, n_10753, n_10754, n_10755, n_10756, n_10757, n_10758, n_10759, n_10760, n_10761, n_10762, n_10763, n_10764, n_10765, n_10766, n_10767, n_10768, n_10769, n_10770, n_10771, n_10772, n_10773, n_10774, n_10775, n_10776, n_10777, n_10778, n_10779, n_10780, n_10781, n_10782, n_10783, n_10784, n_10785, n_10786, n_10787, n_10788, n_10789, n_10790, n_10791, n_10792, n_10793, n_10794, n_10795, n_10796, n_10797, n_10798, n_10799, n_10800, n_10801, n_10802, n_10803, n_10804, n_10805, n_10806, n_10807, n_10808, n_10809, n_10810, n_10811, n_10812, n_10813, n_10814, n_10815, n_10816, n_10817, n_10818, n_10819, n_10820, n_10821, n_10822, n_10823, n_10824, n_10825, n_10826, n_10827, n_10828, n_10829, n_10830, n_10831, n_10832, n_10833, n_10834, n_10835, n_10836, n_10837, n_10838, n_10839, n_10840, n_10841, n_10842, n_10843, n_10844, n_10845, n_10846, n_10847, n_10848, n_10849, n_10850, n_10851, n_10852, n_10853, n_10854, n_10855, n_10856, n_10857, n_10858, n_10859, n_10860, n_10861, n_10862, n_10863, n_10864, n_10865, n_10866, n_10867, n_10868, n_10869, n_10870, n_10871, n_10872, n_10873, n_10874, n_10875, n_10876, n_10877, n_10878, n_10879, n_10880, n_10881, n_10882, n_10883, n_10884, n_10885, n_10886, n_10887, n_10888, n_10889, n_10890, n_10891, n_10892, n_10893, n_10894, n_10895, n_10896, n_10897, n_10898, n_10899, n_10900, n_10901, n_10902, n_10903, n_10904, n_10905, n_10906, n_10907, n_10908, n_10909, n_10910, n_10911, n_10912, n_10913, n_10914, n_10915, n_10916, n_10917, n_10918, n_10919, n_10920, n_10921, n_10922, n_10923, n_10924, n_10925, n_10926, n_10927, n_10928, n_10929, n_10930, n_10931, n_10932, n_10933, n_10934, n_10935, n_10936, n_10937, n_10938, n_10939, n_10940, n_10941, n_10942, n_10943, n_10944, n_10945, n_10946, n_10947, n_10948, n_10949, n_10950, n_10951, n_10952, n_10953, n_10954, n_10955, n_10956, n_10957, n_10958, n_10959, n_10960, n_10961, n_10962, n_10963, n_10964, n_10965, n_10966, n_10967, n_10968, n_10969, n_10970, n_10971, n_10972, n_10973, n_10974, n_10975, n_10976, n_10977, n_10978, n_10979, n_10980, n_10981, n_10982, n_10983, n_10984, n_10985, n_10986, n_10987, n_10988, n_10989, n_10990, n_10991, n_10992, n_10993, n_10994, n_10995, n_10996, n_10997, n_10998, n_10999, n_11000, n_11001, n_11002, n_11003, n_11004, n_11005, n_11006, n_11007, n_11008, n_11009, n_11010, n_11011, n_11012, n_11013, n_11014, n_11015, n_11016, n_11017, n_11018, n_11019, n_11020, n_11021, n_11022, n_11023, n_11024, n_11025, n_11026, n_11027, n_11028, n_11029, n_11030, n_11031, n_11032, n_11033, n_11034, n_11035, n_11036, n_11037, n_11038, n_11039, n_11040, n_11041, n_11042, n_11043, n_11044, n_11045, n_11046, n_11047, n_11048, n_11049, n_11050, n_11051, n_11052, n_11053, n_11054, n_11055, n_11056, n_11057, n_11058, n_11059, n_11060, n_11061, n_11062, n_11063, n_11064, n_11065, n_11066, n_11067, n_11068, n_11069, n_11070, n_11071, n_11072, n_11073, n_11074, n_11075, n_11076, n_11077, n_11078, n_11079, n_11080, n_11081, n_11082, n_11083, n_11084, n_11085, n_11086, n_11087, n_11088, n_11089, n_11090, n_11091, n_11092, n_11093, n_11094, n_11095, n_11096, n_11097, n_11098, y7, n_11099, n_11100, n_11101, n_11102, n_11103, n_11104, n_11105, n_11106, n_11107, n_11108, n_11109, n_11110, n_11111, n_11112, n_11113, n_11114, n_11115, n_11116, n_11117, n_11118, n_11119, n_11120, n_11121, n_11122, n_11123, n_11124, n_11125, n_11126, n_11127, n_11128, n_11129, n_11130, n_11131, n_11132, n_11133, n_11134, n_11135, n_11136, n_11137, n_11138, n_11139, n_11140, n_11141, n_11142, n_11143, n_11144, n_11145, n_11146, n_11147, n_11148, n_11149, n_11150, n_11151, n_11152, n_11153, n_11154, n_11155, n_11156, n_11157, n_11158, n_11159, n_11160, n_11161, n_11162, n_11163, n_11164, n_11165, n_11166, n_11167, n_11168, n_11169, n_11170, n_11171, n_11172, n_11173, n_11174, n_11175, n_11176, n_11177, n_11178, n_11179, n_11180, n_11181, n_11182, n_11183, n_11184, n_11185, n_11186, n_11187, n_11188, n_11189, n_11190, n_11191, n_11192, n_11193, n_11194, n_11195, n_11196, n_11197, n_11198, n_11199, n_11200, n_11201, n_11202, n_11203, n_11204, n_11205, n_11206, n_11207, n_11208, n_11209, n_11210, n_11211, n_11212, n_11213, n_11214, n_11215, n_11216, n_11217, n_11218, n_11219, n_11220, n_11221, n_11222, n_11223, n_11224, n_11225, n_11226, n_11227, n_11228, n_11229, n_11230, n_11231, n_11232, n_11233, n_11234, n_11235, n_11236, n_11237, n_11238, n_11239, n_11240, n_11241, n_11242, n_11243, n_11244, n_11245, n_11246, n_11247, n_11248, n_11249, n_11250, n_11251, n_11252, n_11253, n_11254, n_11255, n_11256, n_11257, n_11258, n_11259, n_11260, n_11261, n_11262, n_11263, n_11264, n_11265, n_11266, n_11267, n_11268, n_11269, n_11270, n_11271, n_11272, n_11273, n_11274, n_11275, n_11276, n_11277, n_11278, n_11279, n_11280, n_11281, n_11282, n_11283, n_11284, n_11285, n_11286, n_11287, n_11288, n_11289, n_11290, n_11291, n_11292, n_11293, n_11294, n_11295, n_11296, n_11297, n_11298, n_11299, n_11300, n_11301, n_11302, n_11303, n_11304, n_11305, n_11306, n_11307, n_11308, n_11309, n_11310, n_11311, n_11312, n_11313, n_11314, n_11315, n_11316, n_11317, n_11318, n_11319, n_11320, n_11321, n_11322, n_11323, n_11324, n_11325, n_11326, n_11327, n_11328, n_11329, n_11330, n_11331, n_11332, n_11333, n_11334, n_11335, n_11336, n_11337, n_11338, n_11339, n_11340, n_11341, n_11342, n_11343, n_11344, n_11345, n_11346, n_11347, n_11348, n_11349, n_11350, n_11351, n_11352, n_11353, n_11354, n_11355, n_11356, n_11357, n_11358, n_11359, n_11360, n_11361, n_11362, n_11363, n_11364, n_11365, n_11366, n_11367, n_11368, n_11369, n_11370, n_11371, n_11372, n_11373, n_11374, n_11375, n_11376, n_11377, n_11378, n_11379, n_11380, n_11381, n_11382, n_11383, n_11384, n_11385, n_11386, n_11387, n_11388, n_11389, n_11390, n_11391, n_11392, n_11393, n_11394, n_11395, n_11396, n_11397, n_11398, n_11399, n_11400, n_11401, n_11402, n_11403, n_11404, n_11405, n_11406, n_11407, n_11408, n_11409, n_11410, n_11411, n_11412, n_11413, n_11414, n_11415, n_11416, n_11417, n_11418, n_11419, n_11420, n_11421, n_11422, n_11423, n_11424, n_11425, n_11426, n_11427, n_11428, n_11429, n_11430, n_11431, n_11432, n_11433, n_11434, n_11435, n_11436, n_11437, n_11438, n_11439, n_11440, n_11441, n_11442, n_11443, n_11444, n_11445, n_11446, n_11447, n_11448, n_11449, n_11450, n_11451, n_11452, n_11453, n_11454, n_11455, n_11456, n_11457, n_11458, n_11459, n_11460, n_11461, n_11462, n_11463, n_11464, n_11465, n_11466, n_11467, n_11468, n_11469, n_11470, n_11471, n_11472, n_11473, n_11474, n_11475, n_11476, n_11477, n_11478, n_11479, n_11480, n_11481, n_11482, n_11483, n_11484, y6, n_11485, n_11486, n_11487, n_11488, n_11489, n_11490, n_11491, n_11492, n_11493, n_11494, n_11495, n_11496, n_11497, n_11498, n_11499, n_11500, n_11501, n_11502, n_11503, n_11504, n_11505, n_11506, n_11507, n_11508, n_11509, n_11510, n_11511, n_11512, n_11513, n_11514, n_11515, n_11516, n_11517, n_11518, n_11519, n_11520, n_11521, n_11522, n_11523, n_11524, n_11525, n_11526, n_11527, n_11528, n_11529, n_11530, n_11531, n_11532, n_11533, n_11534, n_11535, n_11536, n_11537, n_11538, n_11539, n_11540, n_11541, n_11542, n_11543, n_11544, n_11545, n_11546, n_11547, n_11548, n_11549, n_11550, n_11551, n_11552, n_11553, n_11554, n_11555, n_11556, n_11557, n_11558, n_11559, n_11560, n_11561, n_11562, n_11563, n_11564, n_11565, n_11566, n_11567, n_11568, n_11569, n_11570, n_11571, n_11572, n_11573, n_11574, n_11575, n_11576, n_11577, n_11578, n_11579, n_11580, n_11581, n_11582, n_11583, n_11584, n_11585, n_11586, n_11587, n_11588, n_11589, n_11590, n_11591, n_11592, n_11593, n_11594, n_11595, n_11596, n_11597, n_11598, n_11599, n_11600, n_11601, n_11602, n_11603, n_11604, n_11605, n_11606, n_11607, n_11608, n_11609, n_11610, n_11611, n_11612, n_11613, n_11614, n_11615, n_11616, n_11617, n_11618, n_11619, n_11620, n_11621, n_11622, n_11623, n_11624, n_11625, n_11626, n_11627, n_11628, n_11629, n_11630, n_11631, n_11632, n_11633, n_11634, n_11635, n_11636, n_11637, n_11638, n_11639, n_11640, n_11641, n_11642, n_11643, n_11644, n_11645, n_11646, n_11647, n_11648, n_11649, n_11650, n_11651, n_11652, n_11653, n_11654, n_11655, n_11656, n_11657, n_11658, n_11659, n_11660, n_11661, n_11662, n_11663, n_11664, n_11665, n_11666, n_11667, n_11668, n_11669, n_11670, n_11671, n_11672, n_11673, n_11674, n_11675, n_11676, n_11677, n_11678, n_11679, n_11680, n_11681, n_11682, n_11683, n_11684, n_11685, n_11686, n_11687, n_11688, n_11689, n_11690, n_11691, n_11692, n_11693, n_11694, n_11695, n_11696, n_11697, n_11698, n_11699, n_11700, n_11701, n_11702, n_11703, n_11704, n_11705, n_11706, n_11707, n_11708, n_11709, n_11710, n_11711, n_11712, n_11713, n_11714, n_11715, n_11716, n_11717, n_11718, n_11719, n_11720, n_11721, n_11722, n_11723, n_11724, n_11725, n_11726, n_11727, n_11728, n_11729, n_11730, n_11731, n_11732, n_11733, n_11734, n_11735, n_11736, n_11737, n_11738, n_11739, n_11740, n_11741, n_11742, n_11743, n_11744, n_11745, n_11746, n_11747, n_11748, n_11749, n_11750, n_11751, n_11752, n_11753, n_11754, n_11755, n_11756, n_11757, n_11758, n_11759, n_11760, n_11761, n_11762, n_11763, n_11764, n_11765, n_11766, n_11767, n_11768, n_11769, n_11770, n_11771, n_11772, n_11773, n_11774, n_11775, n_11776, n_11777, n_11778, n_11779, n_11780, n_11781, n_11782, n_11783, n_11784, n_11785, n_11786, n_11787, n_11788, n_11789, n_11790, n_11791, n_11792, n_11793, n_11794, n_11795, n_11796, n_11797, n_11798, n_11799, n_11800, n_11801, n_11802, n_11803, n_11804, n_11805, n_11806, n_11807, n_11808, n_11809, n_11810, n_11811, n_11812, n_11813, n_11814, n_11815, n_11816, n_11817, n_11818, n_11819, n_11820, n_11821, n_11822, n_11823, n_11824, n_11825, n_11826, n_11827, n_11828, n_11829, n_11830, n_11831, n_11832, n_11833, n_11834, n_11835, n_11836, n_11837, n_11838, n_11839, n_11840, n_11841, n_11842, n_11843, n_11844, n_11845, n_11846, n_11847, n_11848, n_11849, n_11850, n_11851, n_11852, n_11853, n_11854, n_11855, n_11856, n_11857, n_11858, n_11859, n_11860, n_11861, n_11862, n_11863, y5, n_11864, n_11865, n_11866, n_11867, n_11868, n_11869, n_11870, n_11871, n_11872, n_11873, n_11874, n_11875, n_11876, n_11877, n_11878, n_11879, n_11880, n_11881, n_11882, n_11883, n_11884, n_11885, n_11886, n_11887, n_11888, n_11889, n_11890, n_11891, n_11892, n_11893, n_11894, n_11895, n_11896, n_11897, n_11898, n_11899, n_11900, n_11901, n_11902, n_11903, n_11904, n_11905, n_11906, n_11907, n_11908, n_11909, n_11910, n_11911, n_11912, n_11913, n_11914, n_11915, n_11916, n_11917, n_11918, n_11919, n_11920, n_11921, n_11922, n_11923, n_11924, n_11925, n_11926, n_11927, n_11928, n_11929, n_11930, n_11931, n_11932, n_11933, n_11934, n_11935, n_11936, n_11937, n_11938, n_11939, n_11940, n_11941, n_11942, n_11943, n_11944, n_11945, n_11946, n_11947, n_11948, n_11949, n_11950, n_11951, n_11952, n_11953, n_11954, n_11955, n_11956, n_11957, n_11958, n_11959, n_11960, n_11961, n_11962, n_11963, n_11964, n_11965, n_11966, n_11967, n_11968, n_11969, n_11970, n_11971, n_11972, n_11973, n_11974, n_11975, n_11976, n_11977, n_11978, n_11979, n_11980, n_11981, n_11982, n_11983, n_11984, n_11985, n_11986, n_11987, n_11988, n_11989, n_11990, n_11991, n_11992, n_11993, n_11994, n_11995, n_11996, n_11997, n_11998, n_11999, n_12000, n_12001, n_12002, n_12003, n_12004, n_12005, n_12006, n_12007, n_12008, n_12009, n_12010, n_12011, n_12012, n_12013, n_12014, n_12015, n_12016, n_12017, n_12018, n_12019, n_12020, n_12021, n_12022, n_12023, n_12024, n_12025, n_12026, n_12027, n_12028, n_12029, n_12030, n_12031, n_12032, n_12033, n_12034, n_12035, n_12036, n_12037, n_12038, n_12039, n_12040, n_12041, n_12042, n_12043, n_12044, n_12045, n_12046, n_12047, n_12048, n_12049, n_12050, n_12051, n_12052, n_12053, n_12054, n_12055, n_12056, n_12057, n_12058, n_12059, n_12060, n_12061, n_12062, n_12063, n_12064, n_12065, n_12066, n_12067, n_12068, n_12069, n_12070, n_12071, n_12072, n_12073, n_12074, n_12075, n_12076, n_12077, n_12078, n_12079, n_12080, n_12081, n_12082, n_12083, n_12084, n_12085, n_12086, n_12087, n_12088, n_12089, n_12090, n_12091, n_12092, n_12093, n_12094, n_12095, n_12096, n_12097, n_12098, n_12099, n_12100, n_12101, n_12102, n_12103, n_12104, n_12105, n_12106, n_12107, n_12108, n_12109, n_12110, n_12111, n_12112, n_12113, n_12114, n_12115, n_12116, n_12117, n_12118, n_12119, n_12120, n_12121, n_12122, n_12123, n_12124, n_12125, n_12126, n_12127, n_12128, n_12129, n_12130, n_12131, n_12132, n_12133, n_12134, n_12135, n_12136, n_12137, n_12138, n_12139, n_12140, n_12141, n_12142, n_12143, n_12144, n_12145, n_12146, n_12147, n_12148, n_12149, n_12150, n_12151, n_12152, n_12153, n_12154, n_12155, n_12156, n_12157, n_12158, n_12159, n_12160, n_12161, n_12162, n_12163, n_12164, n_12165, n_12166, n_12167, n_12168, n_12169, n_12170, n_12171, n_12172, n_12173, n_12174, n_12175, n_12176, n_12177, n_12178, n_12179, n_12180, n_12181, n_12182, n_12183, n_12184, n_12185, n_12186, n_12187, n_12188, n_12189, n_12190, n_12191, n_12192, n_12193, n_12194, n_12195, n_12196, n_12197, n_12198, n_12199, n_12200, n_12201, n_12202, n_12203, n_12204, n_12205, n_12206, n_12207, n_12208, n_12209, n_12210, n_12211, n_12212, n_12213, n_12214, n_12215, n_12216, n_12217, n_12218, n_12219, n_12220, n_12221, n_12222, n_12223, n_12224, n_12225, n_12226, n_12227, n_12228, n_12229, n_12230, n_12231, n_12232, n_12233, n_12234, n_12235, n_12236, n_12237, n_12238, n_12239, n_12240, n_12241, n_12242, n_12243, n_12244, n_12245, n_12246, n_12247, n_12248, n_12249, n_12250, n_12251, n_12252, n_12253, n_12254, n_12255, n_12256, n_12257, n_12258, n_12259, n_12260, n_12261, n_12262, n_12263, n_12264, n_12265, n_12266, n_12267, y4, n_12268, n_12269, n_12270, n_12271, n_12272, n_12273, n_12274, n_12275, n_12276, n_12277, n_12278, n_12279, n_12280, n_12281, n_12282, n_12283, n_12284, n_12285, n_12286, n_12287, n_12288, n_12289, n_12290, n_12291, n_12292, n_12293, n_12294, n_12295, n_12296, n_12297, n_12298, n_12299, n_12300, n_12301, n_12302, n_12303, n_12304, n_12305, n_12306, n_12307, n_12308, n_12309, n_12310, n_12311, n_12312, n_12313, n_12314, n_12315, n_12316, n_12317, n_12318, n_12319, n_12320, n_12321, n_12322, n_12323, n_12324, n_12325, n_12326, n_12327, n_12328, n_12329, n_12330, n_12331, n_12332, n_12333, n_12334, n_12335, n_12336, n_12337, n_12338, n_12339, n_12340, n_12341, n_12342, n_12343, n_12344, n_12345, n_12346, n_12347, n_12348, n_12349, n_12350, n_12351, n_12352, n_12353, n_12354, n_12355, n_12356, n_12357, n_12358, n_12359, n_12360, n_12361, n_12362, n_12363, n_12364, n_12365, n_12366, n_12367, n_12368, n_12369, n_12370, n_12371, n_12372, n_12373, n_12374, n_12375, n_12376, n_12377, n_12378, n_12379, n_12380, n_12381, n_12382, n_12383, n_12384, n_12385, n_12386, n_12387, n_12388, n_12389, n_12390, n_12391, n_12392, n_12393, n_12394, n_12395, n_12396, n_12397, n_12398, n_12399, n_12400, n_12401, n_12402, n_12403, n_12404, n_12405, n_12406, n_12407, n_12408, n_12409, n_12410, n_12411, n_12412, n_12413, n_12414, n_12415, n_12416, n_12417, n_12418, n_12419, n_12420, n_12421, n_12422, n_12423, n_12424, n_12425, n_12426, n_12427, n_12428, n_12429, n_12430, n_12431, n_12432, n_12433, n_12434, n_12435, n_12436, n_12437, n_12438, n_12439, n_12440, n_12441, n_12442, n_12443, n_12444, n_12445, n_12446, n_12447, n_12448, n_12449, n_12450, n_12451, n_12452, n_12453, n_12454, n_12455, n_12456, n_12457, n_12458, n_12459, n_12460, n_12461, n_12462, n_12463, n_12464, n_12465, n_12466, n_12467, n_12468, n_12469, n_12470, n_12471, n_12472, n_12473, n_12474, n_12475, n_12476, n_12477, n_12478, n_12479, n_12480, n_12481, n_12482, n_12483, n_12484, n_12485, n_12486, n_12487, n_12488, n_12489, n_12490, n_12491, n_12492, n_12493, n_12494, n_12495, n_12496, n_12497, n_12498, n_12499, n_12500, n_12501, n_12502, n_12503, n_12504, n_12505, n_12506, n_12507, n_12508, n_12509, n_12510, n_12511, n_12512, n_12513, n_12514, n_12515, n_12516, n_12517, n_12518, n_12519, n_12520, n_12521, n_12522, n_12523, n_12524, n_12525, n_12526, n_12527, n_12528, n_12529, n_12530, n_12531, n_12532, n_12533, n_12534, n_12535, n_12536, n_12537, n_12538, n_12539, n_12540, n_12541, n_12542, n_12543, n_12544, n_12545, n_12546, n_12547, n_12548, n_12549, n_12550, n_12551, n_12552, n_12553, n_12554, n_12555, n_12556, n_12557, n_12558, n_12559, n_12560, n_12561, n_12562, n_12563, n_12564, n_12565, n_12566, n_12567, n_12568, n_12569, n_12570, n_12571, n_12572, n_12573, n_12574, n_12575, n_12576, n_12577, n_12578, n_12579, n_12580, n_12581, n_12582, n_12583, n_12584, n_12585, n_12586, n_12587, n_12588, n_12589, n_12590, n_12591, n_12592, n_12593, n_12594, n_12595, n_12596, n_12597, n_12598, n_12599, n_12600, n_12601, n_12602, n_12603, n_12604, n_12605, n_12606, n_12607, n_12608, n_12609, n_12610, n_12611, n_12612, n_12613, n_12614, n_12615, n_12616, n_12617, n_12618, n_12619, n_12620, n_12621, n_12622, n_12623, n_12624, n_12625, n_12626, n_12627, n_12628, n_12629, n_12630, n_12631, n_12632, n_12633, n_12634, n_12635, n_12636, n_12637, n_12638, n_12639, n_12640, n_12641, n_12642, n_12643, n_12644, n_12645, n_12646, n_12647, n_12648, n_12649, n_12650, n_12651, n_12652, n_12653, n_12654, n_12655, n_12656, n_12657, n_12658, n_12659, n_12660, n_12661, n_12662, n_12663, n_12664, n_12665, n_12666, n_12667, y3, n_12668, n_12669, n_12670, n_12671, n_12672, n_12673, n_12674, n_12675, n_12676, n_12677, n_12678, n_12679, n_12680, n_12681, n_12682, n_12683, n_12684, n_12685, n_12686, n_12687, n_12688, n_12689, n_12690, n_12691, n_12692, n_12693, n_12694, n_12695, n_12696, n_12697, n_12698, n_12699, n_12700, n_12701, n_12702, n_12703, n_12704, n_12705, n_12706, n_12707, n_12708, n_12709, n_12710, n_12711, n_12712, n_12713, n_12714, n_12715, n_12716, n_12717, n_12718, n_12719, n_12720, n_12721, n_12722, n_12723, n_12724, n_12725, n_12726, n_12727, n_12728, n_12729, n_12730, n_12731, n_12732, n_12733, n_12734, n_12735, n_12736, n_12737, n_12738, n_12739, n_12740, n_12741, n_12742, n_12743, n_12744, n_12745, n_12746, n_12747, n_12748, n_12749, n_12750, n_12751, n_12752, n_12753, n_12754, n_12755, n_12756, n_12757, n_12758, n_12759, n_12760, n_12761, n_12762, n_12763, n_12764, n_12765, n_12766, n_12767, n_12768, n_12769, n_12770, n_12771, n_12772, n_12773, n_12774, n_12775, n_12776, n_12777, n_12778, n_12779, n_12780, n_12781, n_12782, n_12783, n_12784, n_12785, n_12786, n_12787, n_12788, n_12789, n_12790, n_12791, n_12792, n_12793, n_12794, n_12795, n_12796, n_12797, n_12798, n_12799, n_12800, n_12801, n_12802, n_12803, n_12804, n_12805, n_12806, n_12807, n_12808, n_12809, n_12810, n_12811, n_12812, n_12813, n_12814, n_12815, n_12816, n_12817, n_12818, n_12819, n_12820, n_12821, n_12822, n_12823, n_12824, n_12825, n_12826, n_12827, n_12828, n_12829, n_12830, n_12831, n_12832, n_12833, n_12834, n_12835, n_12836, n_12837, n_12838, n_12839, n_12840, n_12841, n_12842, n_12843, n_12844, n_12845, n_12846, n_12847, n_12848, n_12849, n_12850, n_12851, n_12852, n_12853, n_12854, n_12855, n_12856, n_12857, n_12858, n_12859, n_12860, n_12861, n_12862, n_12863, n_12864, n_12865, n_12866, n_12867, n_12868, n_12869, n_12870, n_12871, n_12872, n_12873, n_12874, n_12875, n_12876, n_12877, n_12878, n_12879, n_12880, n_12881, n_12882, n_12883, n_12884, n_12885, n_12886, n_12887, n_12888, n_12889, n_12890, n_12891, n_12892, n_12893, n_12894, n_12895, n_12896, n_12897, n_12898, n_12899, n_12900, n_12901, n_12902, n_12903, n_12904, n_12905, n_12906, n_12907, n_12908, n_12909, n_12910, n_12911, n_12912, n_12913, n_12914, n_12915, n_12916, n_12917, n_12918, n_12919, n_12920, n_12921, n_12922, n_12923, n_12924, n_12925, n_12926, n_12927, n_12928, n_12929, n_12930, n_12931, n_12932, n_12933, n_12934, n_12935, n_12936, n_12937, n_12938, n_12939, n_12940, n_12941, n_12942, n_12943, n_12944, n_12945, n_12946, n_12947, n_12948, n_12949, n_12950, n_12951, n_12952, n_12953, n_12954, n_12955, n_12956, n_12957, n_12958, n_12959, n_12960, n_12961, n_12962, n_12963, n_12964, n_12965, n_12966, n_12967, n_12968, n_12969, n_12970, n_12971, n_12972, n_12973, n_12974, n_12975, n_12976, n_12977, n_12978, n_12979, n_12980, n_12981, n_12982, n_12983, n_12984, n_12985, n_12986, n_12987, n_12988, n_12989, n_12990, n_12991, n_12992, n_12993, n_12994, n_12995, n_12996, n_12997, n_12998, n_12999, n_13000, n_13001, n_13002, n_13003, n_13004, n_13005, n_13006, n_13007, n_13008, n_13009, n_13010, n_13011, n_13012, n_13013, n_13014, n_13015, n_13016, n_13017, n_13018, n_13019, n_13020, n_13021, n_13022, n_13023, n_13024, n_13025, n_13026, n_13027, n_13028, n_13029, n_13030, n_13031, n_13032, n_13033, n_13034, n_13035, n_13036, n_13037, n_13038, n_13039, n_13040, n_13041, n_13042, n_13043, n_13044, n_13045, n_13046, n_13047, n_13048, n_13049, n_13050, n_13051, n_13052, n_13053, n_13054, n_13055, n_13056, n_13057, n_13058, n_13059, n_13060, n_13061, n_13062, n_13063, n_13064, n_13065, n_13066, n_13067, n_13068, n_13069, n_13070, n_13071, n_13072, n_13073, n_13074, n_13075, n_13076, n_13077, n_13078, n_13079, n_13080, n_13081, n_13082, n_13083, n_13084, n_13085, n_13086, n_13087, n_13088, y2, n_13089, n_13090, n_13091, n_13092, n_13093, n_13094, n_13095, n_13096, n_13097, n_13098, n_13099, n_13100, n_13101, n_13102, n_13103, n_13104, n_13105, n_13106, n_13107, n_13108, n_13109, n_13110, n_13111, n_13112, n_13113, n_13114, n_13115, n_13116, n_13117, n_13118, n_13119, n_13120, n_13121, n_13122, n_13123, n_13124, n_13125, n_13126, n_13127, n_13128, n_13129, n_13130, n_13131, n_13132, n_13133, n_13134, n_13135, n_13136, n_13137, n_13138, n_13139, n_13140, n_13141, n_13142, n_13143, n_13144, n_13145, n_13146, n_13147, n_13148, n_13149, n_13150, n_13151, n_13152, n_13153, n_13154, n_13155, n_13156, n_13157, n_13158, n_13159, n_13160, n_13161, n_13162, n_13163, n_13164, n_13165, n_13166, n_13167, n_13168, n_13169, n_13170, n_13171, n_13172, n_13173, n_13174, n_13175, n_13176, n_13177, n_13178, n_13179, n_13180, n_13181, n_13182, n_13183, n_13184, n_13185, n_13186, n_13187, n_13188, n_13189, n_13190, n_13191, n_13192, n_13193, n_13194, n_13195, n_13196, n_13197, n_13198, n_13199, n_13200, n_13201, n_13202, n_13203, n_13204, n_13205, n_13206, n_13207, n_13208, n_13209, n_13210, n_13211, n_13212, n_13213, n_13214, n_13215, n_13216, n_13217, n_13218, n_13219, n_13220, n_13221, n_13222, n_13223, n_13224, n_13225, n_13226, n_13227, n_13228, n_13229, n_13230, n_13231, n_13232, n_13233, n_13234, n_13235, n_13236, n_13237, n_13238, n_13239, n_13240, n_13241, n_13242, n_13243, n_13244, n_13245, n_13246, n_13247, n_13248, n_13249, n_13250, n_13251, n_13252, n_13253, n_13254, n_13255, n_13256, n_13257, n_13258, n_13259, n_13260, n_13261, n_13262, n_13263, n_13264, n_13265, n_13266, n_13267, n_13268, n_13269, n_13270, n_13271, n_13272, n_13273, n_13274, n_13275, n_13276, n_13277, n_13278, n_13279, n_13280, n_13281, n_13282, n_13283, n_13284, n_13285, n_13286, n_13287, n_13288, n_13289, n_13290, n_13291, n_13292, n_13293, n_13294, n_13295, n_13296, n_13297, n_13298, n_13299, n_13300, n_13301, n_13302, n_13303, n_13304, n_13305, n_13306, n_13307, n_13308, n_13309, n_13310, n_13311, n_13312, n_13313, n_13314, n_13315, n_13316, n_13317, n_13318, n_13319, n_13320, n_13321, n_13322, n_13323, n_13324, n_13325, n_13326, n_13327, n_13328, n_13329, n_13330, n_13331, n_13332, n_13333, n_13334, n_13335, n_13336, n_13337, n_13338, n_13339, n_13340, n_13341, n_13342, n_13343, n_13344, n_13345, n_13346, n_13347, n_13348, n_13349, n_13350, n_13351, n_13352, n_13353, n_13354, n_13355, n_13356, n_13357, n_13358, n_13359, n_13360, n_13361, n_13362, n_13363, n_13364, n_13365, n_13366, n_13367, n_13368, n_13369, n_13370, n_13371, n_13372, n_13373, n_13374, n_13375, n_13376, n_13377, n_13378, n_13379, n_13380, n_13381, n_13382, n_13383, n_13384, n_13385, n_13386, n_13387, n_13388, n_13389, n_13390, n_13391, n_13392, n_13393, n_13394, n_13395, n_13396, n_13397, n_13398, n_13399, n_13400, n_13401, n_13402, n_13403, n_13404, n_13405, n_13406, n_13407, n_13408, n_13409, n_13410, n_13411, n_13412, n_13413, n_13414, n_13415, n_13416, n_13417, n_13418, n_13419, n_13420, n_13421, n_13422, n_13423, n_13424, n_13425, n_13426, n_13427, n_13428, n_13429, n_13430, n_13431, n_13432, n_13433, n_13434, n_13435, n_13436, n_13437, n_13438, n_13439, n_13440, n_13441, n_13442, n_13443, n_13444, n_13445, n_13446, n_13447, n_13448, n_13449, n_13450, n_13451, n_13452, n_13453, n_13454, n_13455, n_13456, n_13457, n_13458, n_13459, n_13460, n_13461, n_13462, n_13463, n_13464, n_13465, n_13466, n_13467, n_13468, n_13469, n_13470, n_13471, n_13472, n_13473, n_13474, n_13475, n_13476, n_13477, n_13478, n_13479, n_13480, n_13481, n_13482, n_13483, n_13484, n_13485, n_13486, n_13487, n_13488, n_13489, n_13490, n_13491, y1, n_13492, n_13493, n_13494, n_13495, n_13496, n_13497, n_13498, n_13499, n_13500, n_13501, n_13502, n_13503, n_13504, n_13505, n_13506, n_13507, n_13508, n_13509, n_13510, n_13511, n_13512, n_13513, n_13514, n_13515, n_13516, n_13517, n_13518, n_13519, n_13520, n_13521, n_13522, n_13523, n_13524, n_13525, n_13526, n_13527, n_13528, n_13529, n_13530, n_13531, n_13532, n_13533, n_13534, n_13535, n_13536, n_13537, n_13538, n_13539, n_13540, n_13541, n_13542, n_13543, n_13544, n_13545, n_13546, n_13547, n_13548, n_13549, n_13550, n_13551, n_13552, n_13553, n_13554, n_13555, n_13556, n_13557, n_13558, n_13559, n_13560, n_13561, n_13562, n_13563, n_13564, n_13565, n_13566, n_13567, n_13568, n_13569, n_13570, n_13571, n_13572, n_13573, n_13574, n_13575, n_13576, n_13577, n_13578, n_13579, n_13580, n_13581, n_13582, n_13583, n_13584, n_13585, n_13586, n_13587, n_13588, n_13589, n_13590, n_13591, n_13592, n_13593, n_13594, n_13595, n_13596, n_13597, n_13598, n_13599, n_13600, n_13601, n_13602, n_13603, n_13604, n_13605, n_13606, n_13607, n_13608, n_13609, n_13610, n_13611, n_13612, n_13613, n_13614, n_13615, n_13616, n_13617, n_13618, n_13619, n_13620, n_13621, n_13622, n_13623, n_13624, n_13625, n_13626, n_13627, n_13628, n_13629, n_13630, n_13631, n_13632, n_13633, n_13634, n_13635, n_13636, n_13637, n_13638, n_13639, n_13640, n_13641, n_13642, n_13643, n_13644, n_13645, n_13646, n_13647, n_13648, n_13649, n_13650, n_13651, n_13652, n_13653, n_13654, n_13655, n_13656, n_13657, n_13658, n_13659, n_13660, n_13661, n_13662, n_13663, n_13664, n_13665, n_13666, n_13667, n_13668, n_13669, n_13670, n_13671, n_13672, n_13673, n_13674, n_13675, n_13676, n_13677, n_13678, n_13679, n_13680, n_13681, n_13682, n_13683, n_13684, n_13685, n_13686, n_13687, n_13688, n_13689, n_13690, n_13691, n_13692, n_13693, n_13694, n_13695, n_13696, n_13697, n_13698, n_13699, n_13700, n_13701, n_13702, n_13703, n_13704, n_13705, n_13706, n_13707, n_13708, n_13709, n_13710, n_13711, n_13712, n_13713, n_13714, n_13715, n_13716, n_13717, n_13718, n_13719, n_13720, n_13721, n_13722, n_13723, n_13724, n_13725, n_13726, n_13727, n_13728, n_13729, n_13730, n_13731, n_13732, n_13733, n_13734, n_13735, n_13736, n_13737, n_13738, n_13739, n_13740, n_13741, n_13742, n_13743, n_13744, n_13745, n_13746, n_13747, n_13748, n_13749, n_13750, n_13751, n_13752, n_13753, n_13754, n_13755, n_13756, n_13757, n_13758, n_13759, n_13760, n_13761, n_13762, n_13763, n_13764, n_13765, n_13766, n_13767, n_13768, n_13769, n_13770, n_13771, n_13772, n_13773, n_13774, n_13775, n_13776, n_13777, n_13778, n_13779, n_13780, n_13781, n_13782, n_13783, n_13784, n_13785, n_13786, n_13787, n_13788, n_13789, n_13790, n_13791, n_13792, n_13793, n_13794, n_13795, n_13796, n_13797, n_13798, n_13799, n_13800, n_13801, n_13802, n_13803, n_13804, n_13805, n_13806, n_13807, n_13808, n_13809, n_13810, n_13811, n_13812, n_13813, n_13814, n_13815, n_13816, n_13817, n_13818, n_13819, n_13820, n_13821, n_13822, n_13823, n_13824, n_13825, n_13826, n_13827, n_13828, n_13829, n_13830, n_13831, n_13832, n_13833, n_13834, n_13835, n_13836, n_13837, n_13838, n_13839, n_13840, n_13841, n_13842, n_13843, n_13844, n_13845, n_13846, n_13847, n_13848, n_13849, n_13850, n_13851, n_13852, n_13853, n_13854, n_13855, n_13856, n_13857, n_13858, n_13859, n_13860, n_13861, n_13862, n_13863, n_13864, n_13865, n_13866, n_13867, n_13868, n_13869, n_13870, n_13871, n_13872, n_13873, n_13874, n_13875, n_13876, n_13877, n_13878, n_13879, n_13880, n_13881, n_13882, n_13883, n_13884, n_13885, n_13886, n_13887, n_13888, n_13889, n_13890, n_13891, n_13892, n_13893, y0, n_13894, n_13895, y127, n_13896, n_13897, n_13898, n_13899, n_13900, n_13901, n_13902, n_13903, n_13904, n_13905, n_13906, n_13907, n_13908, n_13909, n_13910, n_13911, n_13912, n_13913, n_13914, n_13915, n_13916, n_13917, n_13918, n_13919, n_13920, n_13921, n_13922, n_13923, n_13924, n_13925, n_13926, n_13927, n_13928, n_13929, n_13930, n_13931, n_13932, n_13933, n_13934, n_13935, n_13936, n_13937, n_13938, n_13939, n_13940, n_13941, n_13942, n_13943, n_13944, n_13945, n_13946, n_13947, n_13948, n_13949, n_13950, n_13951, n_13952, n_13953, n_13954, n_13955, n_13956, n_13957, n_13958, y64, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y78, y79, y80, y81, y82, y83, y84, y85, y86, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y77, y87, n_13959, n_13960, n_13961, y65;
assign n_0 = ~x2 & ~x3;
assign n_1 = x8 ^ x7;
assign n_2 = ~x21 & ~x22;
assign n_3 = ~x53 & ~x54;
assign n_4 = ~x42 & x64;
assign n_5 = ~x52 & x64;
assign n_6 = ~x58 & x64;
assign n_7 = ~x54 & x64;
assign n_8 = ~x51 & x64;
assign n_9 = ~x49 & x64;
assign n_10 = ~x48 & x64;
assign n_11 = ~x46 & x64;
assign n_12 = ~x45 & x64;
assign n_13 = ~x43 & x64;
assign n_14 = ~x40 & x64;
assign n_15 = ~x37 & x64;
assign n_16 = ~x36 & x64;
assign n_17 = ~x33 & x64;
assign n_18 = x32 & x64;
assign n_19 = ~x31 & x64;
assign n_20 = ~x27 & x64;
assign n_21 = ~x25 & x64;
assign n_22 = ~x24 & x64;
assign n_23 = ~x23 & x64;
assign n_24 = ~x22 & x64;
assign n_25 = ~x20 & x64;
assign n_26 = ~x19 & x64;
assign n_27 = ~x17 & x64;
assign n_28 = ~x16 & x64;
assign n_29 = ~x14 & x64;
assign n_30 = x15 & x64;
assign n_31 = ~x13 & x64;
assign n_32 = ~x12 & x64;
assign n_33 = ~x11 & x64;
assign n_34 = ~x10 & x64;
assign n_35 = ~x9 & x64;
assign n_36 = x7 & x64;
assign n_37 = ~x5 & x64;
assign n_38 = ~x3 & x64;
assign n_39 = ~x2 & x64;
assign n_40 = ~x63 & x64;
assign n_41 = ~x63 & x65;
assign n_42 = x65 ^ x61;
assign n_43 = x61 & ~x65;
assign n_44 = ~x62 & x65;
assign n_45 = x65 ^ x60;
assign n_46 = x64 & ~x65;
assign n_47 = ~x60 & x65;
assign n_48 = x65 ^ x59;
assign n_49 = ~x59 & x65;
assign n_50 = x65 ^ x57;
assign n_51 = ~x58 & x65;
assign n_52 = ~x57 & x65;
assign n_53 = ~x56 & x65;
assign n_54 = x65 ^ x56;
assign n_55 = x65 ^ x55;
assign n_56 = ~x55 & x65;
assign n_57 = x53 & ~x65;
assign n_58 = x51 & x65;
assign n_59 = x65 ^ x50;
assign n_60 = ~x64 & x65;
assign n_61 = x64 & x65;
assign n_62 = x65 ^ x46;
assign n_63 = ~x45 & x65;
assign n_64 = ~x44 & x65;
assign n_65 = ~x43 & ~x65;
assign n_66 = ~x41 & x65;
assign n_67 = ~x40 & x65;
assign n_68 = ~x39 & x65;
assign n_69 = x65 ^ x39;
assign n_70 = ~x38 & x65;
assign n_71 = x37 & ~x65;
assign n_72 = x65 ^ x36;
assign n_73 = x65 ^ x37;
assign n_74 = ~x35 & x65;
assign n_75 = x34 & ~x65;
assign n_76 = x31 & ~x65;
assign n_77 = ~x30 & x65;
assign n_78 = x65 ^ x29;
assign n_79 = x29 & ~x65;
assign n_80 = ~x26 & x65;
assign n_81 = x25 & ~x65;
assign n_82 = ~x24 & x65;
assign n_83 = ~x21 & x65;
assign n_84 = x65 ^ x21;
assign n_85 = ~x22 & x65;
assign n_86 = ~x20 & x65;
assign n_87 = x65 ^ x19;
assign n_88 = ~x19 & x65;
assign n_89 = ~x18 & x65;
assign n_90 = x16 & ~x65;
assign n_91 = x65 ^ x16;
assign n_92 = x65 ^ x17;
assign n_93 = x17 & ~x65;
assign n_94 = ~x15 & x65;
assign n_95 = x65 ^ x64;
assign n_96 = x65 ^ x14;
assign n_97 = x14 & ~x65;
assign n_98 = ~x13 & x65;
assign n_99 = ~x12 & x65;
assign n_100 = x65 ^ x10;
assign n_101 = ~x10 & x65;
assign n_102 = ~x8 & x65;
assign n_103 = x65 ^ x8;
assign n_104 = ~x9 & x65;
assign n_105 = x7 & ~x65;
assign n_106 = x65 ^ x6;
assign n_107 = ~x4 & x65;
assign n_108 = ~x5 & x65;
assign n_109 = x65 ^ x3;
assign n_110 = x3 & ~x65;
assign n_111 = x2 & ~x65;
assign n_112 = x65 ^ x2;
assign n_113 = ~x1 & x65;
assign n_114 = x0 & ~x65;
assign n_115 = x65 ^ x0;
assign n_116 = x65 ^ x1;
assign n_117 = ~x63 & x66;
assign n_118 = ~x65 & ~x66;
assign n_119 = ~x63 & x67;
assign n_120 = x70 & ~x71;
assign n_121 = x70 & x71;
assign n_122 = ~x85 & ~x86;
assign n_123 = ~x84 & ~x87;
assign n_124 = x95 & x96;
assign n_125 = x100 & x101;
assign n_126 = ~x104 & ~x105;
assign n_127 = ~x106 & ~x107;
assign n_128 = ~x111 & ~x112;
assign n_129 = ~x113 & ~x114;
assign n_130 = x117 & x118;
assign n_131 = ~x126 & ~x127;
assign n_132 = ~x64 & n_1;
assign n_133 = n_4 ^ x65;
assign n_134 = n_5 ^ x65;
assign n_135 = n_6 ^ x65;
assign n_136 = n_8 ^ x65;
assign n_137 = ~x50 & n_8;
assign n_138 = n_9 ^ x65;
assign n_139 = n_10 ^ x65;
assign n_140 = n_11 ^ x65;
assign n_141 = n_12 ^ x65;
assign n_142 = ~x44 & n_13;
assign n_143 = n_13 ^ x65;
assign n_144 = n_14 ^ x65;
assign n_145 = x65 & n_15;
assign n_146 = ~x38 & n_15;
assign n_147 = n_15 ^ x65;
assign n_148 = n_16 ^ x65;
assign n_149 = n_17 ^ x65;
assign n_150 = n_18 ^ x64;
assign n_151 = n_19 ^ x32;
assign n_152 = ~x30 & n_19;
assign n_153 = n_21 ^ x65;
assign n_154 = ~x24 & n_21;
assign n_155 = n_22 ^ x65;
assign n_156 = ~x65 & ~n_24;
assign n_157 = n_24 ^ x65;
assign n_158 = ~x65 ^ ~n_25;
assign n_159 = n_25 ^ x65;
assign n_160 = ~x18 & n_26;
assign n_161 = ~x65 ^ ~n_27;
assign n_162 = n_27 ^ x65;
assign n_163 = ~x17 & n_28;
assign n_164 = n_28 ^ x65;
assign n_165 = ~x15 & n_28;
assign n_166 = n_29 ^ x65;
assign n_167 = ~n_29 & ~n_31;
assign n_168 = n_32 ^ x65;
assign n_169 = n_34 ^ x65;
assign n_170 = n_35 ^ x65;
assign n_171 = ~x8 & n_35;
assign n_172 = ~x6 & n_36;
assign n_173 = n_38 ^ x65;
assign n_174 = ~x65 ^ ~n_38;
assign n_175 = ~x1 & n_39;
assign n_176 = n_39 ^ x65;
assign n_177 = ~x66 & ~n_41;
assign n_178 = n_42 ^ n_43;
assign n_179 = x64 & ~n_43;
assign n_180 = n_44 ^ x65;
assign n_181 = n_46 ^ x64;
assign n_182 = n_52 ^ x56;
assign n_183 = n_52 ^ n_50;
assign n_184 = n_55 ^ n_56;
assign n_185 = n_57 ^ x65;
assign n_186 = n_60 ^ x65;
assign n_187 = x22 & n_60;
assign n_188 = ~x21 & n_60;
assign n_189 = n_26 ^ n_60;
assign n_190 = n_60 ^ n_46;
assign n_191 = x14 & n_60;
assign n_192 = n_33 ^ n_60;
assign n_193 = ~x11 & n_60;
assign n_194 = n_65 ^ x43;
assign n_195 = x64 & n_66;
assign n_196 = n_66 ^ x65;
assign n_197 = n_66 ^ x42;
assign n_198 = x64 & n_67;
assign n_199 = n_67 ^ x64;
assign n_200 = ~n_67 & ~n_68;
assign n_201 = n_68 ^ n_69;
assign n_202 = x36 & n_71;
assign n_203 = n_72 ^ n_73;
assign n_204 = x64 & n_74;
assign n_205 = n_75 ^ x65;
assign n_206 = ~n_75 & n_17;
assign n_207 = n_18 & ~n_76;
assign n_208 = n_76 ^ x31;
assign n_209 = n_78 ^ x28;
assign n_210 = n_79 ^ n_77;
assign n_211 = x64 & n_80;
assign n_212 = n_81 ^ x25;
assign n_213 = ~x64 & n_82;
assign n_214 = n_2 ^ n_83;
assign n_215 = ~x22 & n_83;
assign n_216 = n_24 & ~n_83;
assign n_217 = n_84 ^ n_85;
assign n_218 = n_87 ^ n_88;
assign n_219 = n_25 & ~n_88;
assign n_220 = n_89 ^ n_88;
assign n_221 = x15 & n_90;
assign n_222 = n_90 ^ n_91;
assign n_223 = n_92 ^ n_93;
assign n_224 = n_95 ^ n_30;
assign n_225 = n_96 ^ n_97;
assign n_226 = ~n_97 & n_31;
assign n_227 = x13 & n_97;
assign n_228 = n_29 & ~n_98;
assign n_229 = x64 & n_99;
assign n_230 = n_100 ^ n_101;
assign n_231 = ~x64 & n_101;
assign n_232 = n_101 ^ x65;
assign n_233 = x64 & n_102;
assign n_234 = x64 & ~n_105;
assign n_235 = n_105 ^ x65;
assign n_236 = n_37 & n_106;
assign n_237 = ~x64 & n_107;
assign n_238 = n_107 ^ n_108;
assign n_239 = n_109 ^ n_110;
assign n_240 = x1 & n_111;
assign n_241 = n_111 ^ n_112;
assign n_242 = x1 & ~n_114;
assign n_243 = n_115 ^ n_116;
assign n_244 = ~n_40 & n_118;
assign n_245 = n_122 & n_123;
assign n_246 = ~x108 & n_126;
assign n_247 = n_128 & n_129;
assign n_248 = ~x125 & n_131;
assign n_249 = n_132 ^ x7;
assign n_250 = n_143 & n_4;
assign n_251 = n_150 ^ x65;
assign n_252 = n_151 ^ n_150;
assign n_253 = ~n_158 ^ n_26;
assign n_254 = ~n_88 ^ ~n_160;
assign n_255 = x7 ^ n_172;
assign n_256 = ~n_174 ^ n_173;
assign n_257 = x62 & ~n_178;
assign n_258 = ~n_179 & ~n_44;
assign n_259 = x64 & ~n_180;
assign n_260 = n_181 ^ n_179;
assign n_261 = x56 & n_183;
assign n_262 = x54 & n_184;
assign n_263 = n_7 & ~n_184;
assign n_264 = n_185 ^ x53;
assign n_265 = n_189 ^ n_186;
assign n_266 = n_192 ^ n_186;
assign n_267 = x10 & n_193;
assign n_268 = x64 & ~n_194;
assign n_269 = n_199 & ~n_200;
assign n_270 = n_14 & ~n_201;
assign n_271 = x64 & ~n_201;
assign n_272 = x38 & n_201;
assign n_273 = n_202 ^ x37;
assign n_274 = n_203 ^ x65;
assign n_275 = n_207 ^ x32;
assign n_276 = n_214 ^ n_215;
assign n_277 = x18 & n_218;
assign n_278 = x64 & n_220;
assign n_279 = n_221 ^ x16;
assign n_280 = ~n_222 ^ ~n_165;
assign n_281 = n_94 ^ n_222;
assign n_282 = ~x13 & n_225;
assign n_283 = ~n_225 & ~n_226;
assign n_284 = n_227 ^ x14;
assign n_285 = x9 & n_230;
assign n_286 = n_231 ^ n_101;
assign n_287 = n_232 ^ x9;
assign n_288 = x3 & n_237;
assign n_289 = x64 & n_238;
assign n_290 = n_240 ^ x2;
assign n_291 = ~n_241 ^ ~n_175;
assign n_292 = n_113 ^ n_241;
assign n_293 = n_243 ^ x65;
assign n_294 = n_127 & n_246;
assign n_295 = ~x124 & n_248;
assign n_296 = x65 & ~n_249;
assign n_297 = x33 & n_251;
assign n_298 = n_259 ^ x65;
assign n_299 = n_260 ^ x65;
assign n_300 = n_261 ^ x57;
assign n_301 = n_262 ^ x55;
assign n_302 = n_267 ^ n_193;
assign n_303 = n_272 ^ x39;
assign n_304 = n_274 ^ x64;
assign n_305 = n_276 ^ n_217;
assign n_306 = x64 & n_276;
assign n_307 = n_277 ^ x19;
assign n_308 = n_88 ^ n_278;
assign n_309 = x64 & n_281;
assign n_310 = n_284 ^ n_225;
assign n_311 = n_285 ^ x10;
assign n_312 = n_286 ^ n_169;
assign n_313 = n_289 ^ n_108;
assign n_314 = x64 & n_292;
assign n_315 = n_293 ^ x64;
assign n_316 = ~x123 & n_295;
assign n_317 = ~x66 & ~n_298;
assign n_318 = n_300 ^ x65;
assign n_319 = n_301 ^ n_56;
assign n_320 = n_302 ^ n_231;
assign n_321 = n_303 ^ n_68;
assign n_322 = ~n_274 & ~n_304;
assign n_323 = n_305 ^ n_2;
assign n_324 = ~n_85 & ~n_306;
assign n_325 = n_222 ^ n_309;
assign n_326 = n_312 ^ n_101;
assign n_327 = n_35 ^ n_312;
assign n_328 = ~n_312 & ~n_35;
assign n_329 = n_241 ^ n_314;
assign n_330 = ~n_293 & ~n_315;
assign n_331 = ~x122 & n_316;
assign n_332 = x66 ^ n_317;
assign n_333 = x63 & n_317;
assign n_334 = n_182 ^ n_318;
assign n_335 = n_322 ^ x37;
assign n_336 = n_322 ^ n_274;
assign n_337 = ~x11 & n_326;
assign n_338 = n_327 ^ n_328;
assign n_339 = n_330 ^ x1;
assign n_340 = n_330 ^ n_293;
assign n_341 = ~x121 & n_331;
assign n_342 = n_331 ^ n_316;
assign n_343 = n_334 ^ n_300;
assign n_344 = n_335 ^ n_274;
assign n_345 = ~n_101 & n_338;
assign n_346 = n_338 ^ n_101;
assign n_347 = n_339 ^ n_293;
assign n_348 = ~x120 & n_341;
assign n_349 = n_346 ^ n_34;
assign n_350 = ~x119 & n_348;
assign n_351 = n_345 ^ n_349;
assign n_352 = ~x118 & n_350;
assign n_353 = ~x117 & n_352;
assign n_354 = n_353 & ~x116;
assign n_355 = ~x115 & n_354;
assign n_356 = n_355 & n_129;
assign n_357 = ~x114 & n_355;
assign n_358 = n_355 & n_247;
assign n_359 = ~x112 & n_356;
assign n_360 = ~x110 & n_358;
assign n_361 = ~x109 & n_360;
assign n_362 = ~x108 & n_361;
assign n_363 = n_361 & n_294;
assign n_364 = n_127 & n_362;
assign n_365 = ~x107 & n_362;
assign n_366 = ~x103 & n_363;
assign n_367 = ~x105 & n_364;
assign n_368 = ~x102 & n_366;
assign n_369 = ~x101 & n_368;
assign n_370 = ~x100 & n_369;
assign n_371 = ~x99 & n_370;
assign n_372 = ~x98 & n_371;
assign n_373 = ~x97 & n_372;
assign n_374 = ~x96 & n_373;
assign n_375 = ~x95 & n_374;
assign n_376 = ~x94 & n_375;
assign n_377 = ~x93 & n_376;
assign n_378 = ~x92 & n_377;
assign n_379 = ~x91 & n_378;
assign n_380 = ~x90 & n_379;
assign n_381 = ~x89 & n_380;
assign n_382 = ~x88 & n_381;
assign n_383 = ~x87 & n_382;
assign n_384 = n_382 & n_245;
assign n_385 = n_122 & n_383;
assign n_386 = ~x86 & n_383;
assign n_387 = ~x83 & n_384;
assign n_388 = ~x82 & n_387;
assign n_389 = ~x81 & n_388;
assign n_390 = ~x80 & n_389;
assign n_391 = ~x79 & n_390;
assign n_392 = ~x78 & n_391;
assign n_393 = ~x77 & n_392;
assign n_394 = ~x76 & n_393;
assign n_395 = ~x75 & n_394;
assign n_396 = ~x74 & n_395;
assign n_397 = ~x73 & n_396;
assign n_398 = ~x72 & n_397;
assign n_399 = ~x71 & n_398;
assign n_400 = ~x70 & n_399;
assign n_401 = ~x69 & n_400;
assign n_402 = ~x68 & n_401;
assign n_403 = ~x67 & n_402;
assign n_404 = n_402 & ~n_119;
assign n_405 = n_403 & n_177;
assign n_406 = n_403 & ~n_117;
assign n_407 = n_403 & n_244;
assign n_408 = x64 & n_405;
assign n_409 = n_257 & ~n_405;
assign y63 = n_407;
assign n_410 = n_408 ^ x62;
assign n_411 = n_178 & n_408;
assign n_412 = ~x62 & n_408;
assign n_413 = ~n_258 & ~n_409;
assign n_414 = n_410 ^ n_178;
assign n_415 = n_410 & ~n_411;
assign n_416 = n_412 ^ n_405;
assign n_417 = n_332 & ~n_413;
assign n_418 = ~n_333 & n_413;
assign n_419 = n_414 ^ n_415;
assign y62 = n_416;
assign n_420 = n_417 ^ x66;
assign n_421 = ~n_418 & n_406;
assign n_422 = n_403 & ~n_420;
assign n_423 = x61 ^ n_421;
assign n_424 = n_299 & n_421;
assign n_425 = x64 & n_421;
assign y61 = n_421;
assign n_426 = x63 & ~n_422;
assign n_427 = n_423 ^ x60;
assign n_428 = n_424 ^ n_412;
assign n_429 = n_403 & n_426;
assign n_430 = ~n_45 & n_427;
assign n_431 = n_428 ^ n_415;
assign n_432 = n_430 ^ x60;
assign n_433 = x64 & ~n_432;
assign n_434 = ~n_419 & ~n_433;
assign n_435 = x66 ^ n_434;
assign n_436 = n_431 ^ n_434;
assign n_437 = ~n_435 & ~n_436;
assign n_438 = n_437 ^ x66;
assign n_439 = n_429 & ~n_438;
assign n_440 = n_438 ^ x67;
assign n_441 = ~n_438 & n_404;
assign n_442 = n_379 ^ ~n_439;
assign n_443 = n_402 & n_440;
assign n_444 = ~n_429 & ~n_441;
assign n_445 = ~n_443 & n_426;
assign n_446 = x64 & ~n_444;
assign n_447 = x60 ^ n_444;
assign n_448 = x65 & ~n_444;
assign n_449 = ~n_435 & ~n_444;
assign y60 = ~n_444;
assign n_450 = x69 & ~n_445;
assign n_451 = ~n_446 & n_47;
assign n_452 = n_446 & ~n_447;
assign n_453 = n_447 ^ x59;
assign n_454 = n_448 ^ x61;
assign n_455 = n_449 ^ n_431;
assign n_456 = n_400 & ~n_450;
assign n_457 = n_450 ^ x69;
assign n_458 = n_425 ^ n_452;
assign n_459 = ~n_48 & ~n_453;
assign n_460 = n_458 ^ n_454;
assign n_461 = n_459 ^ x59;
assign n_462 = n_460 ^ x66;
assign n_463 = x64 & ~n_461;
assign n_464 = ~n_451 & ~n_463;
assign n_465 = n_460 ^ n_464;
assign n_466 = x66 ^ n_464;
assign n_467 = ~n_462 & ~n_465;
assign n_468 = n_467 ^ x66;
assign n_469 = n_468 ^ x67;
assign n_470 = n_455 ^ n_468;
assign n_471 = n_469 & n_470;
assign n_472 = n_471 ^ x67;
assign n_473 = n_472 ^ x68;
assign n_474 = n_472 ^ n_445;
assign n_475 = n_473 & n_445;
assign n_476 = n_473 & n_474;
assign n_477 = n_401 & n_475;
assign n_478 = n_476 ^ x68;
assign n_479 = n_445 ^ n_477;
assign n_480 = n_401 & ~n_478;
assign n_481 = n_457 ^ n_479;
assign n_482 = x64 & n_480;
assign n_483 = x65 & n_480;
assign n_484 = x65 ^ n_480;
assign n_485 = n_48 ^ n_480;
assign n_486 = ~n_466 & n_480;
assign n_487 = n_469 & n_480;
assign y59 = n_480;
assign n_488 = n_482 ^ x59;
assign n_489 = n_483 ^ x60;
assign n_490 = n_482 & n_484;
assign n_491 = x58 & ~n_485;
assign n_492 = n_486 ^ n_460;
assign n_493 = n_487 ^ n_455;
assign n_494 = n_482 & n_488;
assign n_495 = n_491 ^ n_48;
assign n_496 = n_494 ^ n_446;
assign n_497 = x64 & ~n_495;
assign n_498 = n_496 ^ n_489;
assign n_499 = n_490 ^ n_497;
assign n_500 = n_498 ^ x66;
assign n_501 = n_49 ^ n_499;
assign n_502 = n_501 ^ n_498;
assign n_503 = n_501 ^ x66;
assign n_504 = ~n_500 & n_502;
assign n_505 = n_504 ^ x66;
assign n_506 = n_505 ^ x67;
assign n_507 = n_492 ^ n_505;
assign n_508 = n_506 & n_507;
assign n_509 = n_508 ^ x67;
assign n_510 = n_509 ^ x68;
assign n_511 = n_493 ^ n_509;
assign n_512 = n_510 & ~n_511;
assign n_513 = n_512 ^ n_509;
assign n_514 = n_513 & ~n_481;
assign n_515 = n_456 & ~n_514;
assign n_516 = n_479 & ~n_515;
assign n_517 = x58 ^ n_515;
assign n_518 = x64 & n_515;
assign n_519 = n_503 & n_515;
assign n_520 = n_506 & n_515;
assign n_521 = n_510 & n_515;
assign y58 = n_515;
assign n_522 = n_135 & n_515;
assign n_523 = n_516 ^ n_439;
assign n_524 = n_517 ^ x65;
assign n_525 = n_518 ^ x58;
assign n_526 = ~n_518 & n_51;
assign n_527 = n_519 ^ n_498;
assign n_528 = n_520 ^ n_492;
assign n_529 = n_521 ^ n_493;
assign n_530 = n_488 ^ n_522;
assign n_531 = ~n_398 & n_523;
assign n_532 = x71 & ~n_523;
assign n_533 = n_523 & n_120;
assign n_534 = ~n_50 & n_524;
assign n_535 = n_530 ^ x66;
assign n_536 = n_534 ^ x57;
assign n_537 = x64 & ~n_536;
assign n_538 = ~n_537 & ~n_526;
assign n_539 = n_530 ^ n_538;
assign n_540 = x66 ^ n_538;
assign n_541 = ~n_535 & ~n_539;
assign n_542 = n_541 ^ x66;
assign n_543 = n_542 ^ x67;
assign n_544 = n_527 ^ n_542;
assign n_545 = n_543 & n_544;
assign n_546 = n_545 ^ x67;
assign n_547 = n_546 ^ x68;
assign n_548 = n_528 ^ n_546;
assign n_549 = n_547 & n_548;
assign n_550 = n_549 ^ x68;
assign n_551 = n_550 ^ x69;
assign n_552 = n_529 ^ n_550;
assign n_553 = n_551 & n_552;
assign n_554 = n_553 ^ x69;
assign n_555 = n_554 ^ x70;
assign n_556 = n_554 ^ n_523;
assign n_557 = n_554 & n_533;
assign n_558 = n_555 & ~n_556;
assign n_559 = n_558 ^ n_554;
assign n_560 = n_399 & ~n_559;
assign n_561 = n_523 & ~n_560;
assign n_562 = x65 & n_560;
assign n_563 = x64 & n_560;
assign n_564 = ~n_540 & n_560;
assign n_565 = n_543 & n_560;
assign n_566 = n_547 & n_560;
assign n_567 = n_551 & n_560;
assign y57 = n_560;
assign n_568 = ~n_300 & ~n_562;
assign n_569 = n_525 ^ n_562;
assign n_570 = n_52 & ~n_563;
assign n_571 = n_563 ^ x57;
assign n_572 = n_564 ^ n_530;
assign n_573 = n_565 ^ n_527;
assign n_574 = n_566 ^ n_528;
assign n_575 = n_567 ^ n_529;
assign n_576 = n_568 ^ n_300;
assign n_577 = n_563 & n_571;
assign n_578 = n_576 ^ n_560;
assign n_579 = n_577 ^ n_569;
assign n_580 = ~n_343 & ~n_578;
assign n_581 = n_334 ^ n_580;
assign n_582 = x64 & ~n_581;
assign n_583 = ~n_570 & ~n_582;
assign n_584 = x66 ^ n_583;
assign n_585 = n_579 ^ n_583;
assign n_586 = ~n_584 & ~n_585;
assign n_587 = n_586 ^ x66;
assign n_588 = n_587 ^ x67;
assign n_589 = n_572 ^ n_587;
assign n_590 = n_588 & n_589;
assign n_591 = n_590 ^ x67;
assign n_592 = n_591 ^ x68;
assign n_593 = n_573 ^ n_591;
assign n_594 = n_592 & n_593;
assign n_595 = n_594 ^ x68;
assign n_596 = n_595 ^ x69;
assign n_597 = n_574 ^ n_595;
assign n_598 = n_596 & n_597;
assign n_599 = n_598 ^ x69;
assign n_600 = n_599 ^ x70;
assign n_601 = n_575 ^ n_599;
assign n_602 = n_600 & ~n_601;
assign n_603 = n_602 ^ n_599;
assign n_604 = ~n_532 & ~n_603;
assign n_605 = ~n_557 ^ ~n_604;
assign n_606 = n_398 & n_605;
assign n_607 = n_561 & ~n_606;
assign n_608 = x65 ^ n_606;
assign n_609 = x64 & n_606;
assign n_610 = n_54 ^ n_606;
assign n_611 = x65 & n_606;
assign n_612 = ~n_584 & n_606;
assign n_613 = n_588 & n_606;
assign n_614 = n_592 & n_606;
assign n_615 = n_596 & n_606;
assign n_616 = n_600 & n_606;
assign y56 = n_606;
assign n_617 = ~n_439 ^ ~n_607;
assign n_618 = ~n_608 & n_609;
assign n_619 = ~x56 & n_609;
assign n_620 = x64 & ~n_610;
assign n_621 = n_612 ^ n_579;
assign n_622 = n_613 ^ n_572;
assign n_623 = n_614 ^ n_573;
assign n_624 = n_615 ^ n_574;
assign n_625 = n_616 ^ n_575;
assign n_626 = ~n_617 ^ n_561;
assign n_627 = n_398 & n_617;
assign n_628 = n_53 ^ n_618;
assign n_629 = n_611 ^ n_619;
assign n_630 = ~x55 & n_620;
assign n_631 = ~x72 ^ n_626;
assign n_632 = n_629 ^ n_571;
assign n_633 = n_628 ^ n_630;
assign n_634 = ~n_631 ^ n_561;
assign n_635 = n_633 ^ x66;
assign n_636 = n_632 ^ n_633;
assign n_637 = n_397 & n_634;
assign n_638 = n_635 & n_636;
assign n_639 = n_638 ^ x66;
assign n_640 = n_639 ^ x67;
assign n_641 = n_621 ^ n_639;
assign n_642 = n_640 & n_641;
assign n_643 = n_642 ^ x67;
assign n_644 = n_643 ^ x68;
assign n_645 = n_622 ^ n_643;
assign n_646 = n_644 & n_645;
assign n_647 = n_646 ^ x68;
assign n_648 = n_647 ^ x69;
assign n_649 = n_623 ^ n_647;
assign n_650 = n_648 & n_649;
assign n_651 = n_650 ^ x69;
assign n_652 = n_651 ^ x70;
assign n_653 = n_624 ^ n_651;
assign n_654 = n_652 & n_653;
assign n_655 = n_654 ^ x70;
assign n_656 = n_655 ^ x71;
assign n_657 = n_625 ^ n_655;
assign n_658 = n_656 & ~n_657;
assign n_659 = n_658 ^ n_655;
assign n_660 = n_637 & ~n_659;
assign n_661 = n_627 ^ n_660;
assign n_662 = n_531 & ~n_660;
assign n_663 = n_656 & n_661;
assign n_664 = ~x65 & n_661;
assign n_665 = x64 & n_661;
assign n_666 = n_635 & n_661;
assign n_667 = n_640 & n_661;
assign n_668 = n_644 & n_661;
assign n_669 = n_648 & n_661;
assign n_670 = n_652 & n_661;
assign y55 = n_661;
assign n_671 = x72 ^ n_662;
assign n_672 = x72 & ~n_662;
assign n_673 = n_663 ^ n_625;
assign n_674 = n_664 ^ x56;
assign n_675 = ~n_664 & n_263;
assign n_676 = ~x55 & n_665;
assign n_677 = n_665 ^ x55;
assign n_678 = n_665 & n_319;
assign n_679 = n_666 ^ n_632;
assign n_680 = n_667 ^ n_621;
assign n_681 = n_668 ^ n_622;
assign n_682 = n_669 ^ n_623;
assign n_683 = n_670 ^ n_624;
assign n_684 = n_671 ^ n_672;
assign n_685 = n_673 ^ x72;
assign n_686 = n_673 & n_662;
assign n_687 = n_674 ^ n_609;
assign n_688 = n_676 ^ n_661;
assign n_689 = n_56 ^ n_678;
assign n_690 = n_682 ^ x70;
assign n_691 = x70 & ~n_682;
assign n_692 = x71 & ~n_682;
assign n_693 = n_683 ^ ~n_121;
assign n_694 = n_683 ^ x71;
assign n_695 = n_684 ^ x73;
assign n_696 = n_687 ^ n_688;
assign n_697 = ~n_689 & ~n_675;
assign n_698 = n_690 ^ n_691;
assign n_699 = n_683 ^ n_691;
assign n_700 = n_696 ^ x66;
assign n_701 = n_696 ^ n_697;
assign n_702 = x66 ^ n_697;
assign n_703 = ~n_694 & n_699;
assign n_704 = ~n_700 & ~n_701;
assign n_705 = n_703 ^ x71;
assign n_706 = n_704 ^ x66;
assign n_707 = n_706 ^ x67;
assign n_708 = n_679 ^ n_706;
assign n_709 = n_707 & n_708;
assign n_710 = n_709 ^ x67;
assign n_711 = n_710 ^ x68;
assign n_712 = n_680 ^ n_710;
assign n_713 = n_711 & n_712;
assign n_714 = n_713 ^ x68;
assign n_715 = n_714 ^ x69;
assign n_716 = n_681 ^ n_714;
assign n_717 = n_715 & n_716;
assign n_718 = n_717 ^ x69;
assign n_719 = n_718 & ~n_698;
assign n_720 = n_718 ^ x70;
assign n_721 = n_718 & n_692;
assign n_722 = n_719 & n_693;
assign n_723 = ~n_691 & ~n_719;
assign n_724 = ~n_705 & ~n_721;
assign n_725 = n_723 ^ x71;
assign n_726 = ~n_722 & n_724;
assign n_727 = n_673 ^ n_726;
assign n_728 = x72 ^ n_726;
assign n_729 = n_686 & n_726;
assign n_730 = ~n_685 & ~n_727;
assign n_731 = n_730 ^ n_672;
assign n_732 = ~n_695 & ~n_731;
assign n_733 = ~n_732 & ~n_729;
assign n_734 = n_396 & ~n_733;
assign n_735 = n_662 & ~n_734;
assign n_736 = x65 ^ n_734;
assign n_737 = x64 & n_734;
assign n_738 = ~n_702 & n_734;
assign n_739 = n_707 & n_734;
assign n_740 = n_711 & n_734;
assign n_741 = n_715 & n_734;
assign n_742 = n_720 & n_734;
assign n_743 = ~n_728 & n_734;
assign y54 = n_734;
assign n_744 = ~n_725 & n_734;
assign n_745 = ~n_439 ^ ~n_735;
assign n_746 = x54 & n_737;
assign n_747 = n_737 ^ x54;
assign n_748 = n_737 & ~n_185;
assign n_749 = ~n_737 & n_3;
assign n_750 = n_738 ^ n_696;
assign n_751 = n_739 ^ n_679;
assign n_752 = n_740 ^ n_680;
assign n_753 = n_741 ^ n_681;
assign n_754 = n_742 ^ n_682;
assign n_755 = n_743 ^ n_673;
assign n_756 = n_683 ^ n_744;
assign n_757 = ~n_745 ^ x74;
assign n_758 = n_736 ^ n_746;
assign n_759 = n_748 ^ x65;
assign n_760 = ~n_264 ^ ~n_749;
assign n_761 = ~n_758 & n_734;
assign n_762 = ~n_747 & n_759;
assign n_763 = x64 & n_760;
assign n_764 = n_737 ^ n_761;
assign n_765 = ~n_763 & ~n_762;
assign n_766 = n_677 ^ n_764;
assign n_767 = x66 ^ n_765;
assign n_768 = n_766 ^ x66;
assign n_769 = n_766 ^ n_765;
assign n_770 = ~n_768 & ~n_769;
assign n_771 = n_770 ^ x66;
assign n_772 = n_771 ^ x67;
assign n_773 = n_750 ^ n_771;
assign n_774 = n_772 & n_773;
assign n_775 = n_774 ^ x67;
assign n_776 = n_775 ^ x68;
assign n_777 = n_751 ^ n_775;
assign n_778 = n_776 & n_777;
assign n_779 = n_778 ^ x68;
assign n_780 = n_779 ^ x69;
assign n_781 = n_752 ^ n_779;
assign n_782 = n_780 & n_781;
assign n_783 = n_782 ^ x69;
assign n_784 = n_783 ^ x70;
assign n_785 = n_753 ^ n_783;
assign n_786 = n_784 & n_785;
assign n_787 = n_786 ^ x70;
assign n_788 = n_787 ^ x71;
assign n_789 = n_754 ^ n_787;
assign n_790 = n_788 & n_789;
assign n_791 = n_790 ^ x71;
assign n_792 = n_791 ^ x72;
assign n_793 = n_756 ^ n_791;
assign n_794 = n_792 & n_793;
assign n_795 = n_794 ^ x72;
assign n_796 = n_795 ^ x73;
assign n_797 = n_755 ^ n_795;
assign n_798 = n_796 & ~n_797;
assign n_799 = n_798 ^ n_795;
assign n_800 = n_799 ^ x74;
assign n_801 = n_757 & n_800;
assign n_802 = x74 ^ n_801;
assign n_803 = n_395 & ~n_802;
assign n_804 = x53 ^ n_803;
assign n_805 = x64 & n_803;
assign n_806 = x65 & n_803;
assign n_807 = ~n_767 & n_803;
assign n_808 = n_772 & n_803;
assign n_809 = n_776 & n_803;
assign n_810 = n_780 & n_803;
assign n_811 = n_784 & n_803;
assign n_812 = n_788 & n_803;
assign n_813 = n_792 & n_803;
assign n_814 = n_796 & n_803;
assign n_815 = ~n_439 ^ n_803;
assign y53 = n_803;
assign n_816 = n_5 & ~n_804;
assign n_817 = n_5 ^ n_805;
assign n_818 = ~x53 & n_805;
assign n_819 = n_807 ^ n_766;
assign n_820 = n_808 ^ n_750;
assign n_821 = n_809 ^ n_751;
assign n_822 = n_810 ^ n_752;
assign n_823 = n_811 ^ n_753;
assign n_824 = n_812 ^ n_754;
assign n_825 = n_813 ^ n_756;
assign n_826 = n_814 ^ n_755;
assign n_827 = n_745 & n_815;
assign n_828 = n_816 ^ n_264;
assign n_829 = x65 & n_817;
assign n_830 = n_818 ^ n_806;
assign n_831 = n_827 ^ x75;
assign n_832 = n_828 ^ n_829;
assign n_833 = n_830 ^ n_737;
assign n_834 = n_832 ^ x66;
assign n_835 = n_833 ^ x54;
assign n_836 = n_835 ^ n_832;
assign n_837 = n_834 & n_836;
assign n_838 = n_837 ^ x66;
assign n_839 = n_838 ^ x67;
assign n_840 = n_819 ^ n_838;
assign n_841 = n_839 & n_840;
assign n_842 = n_841 ^ x67;
assign n_843 = n_842 ^ x68;
assign n_844 = n_820 ^ n_842;
assign n_845 = n_843 & n_844;
assign n_846 = n_845 ^ x68;
assign n_847 = n_846 ^ x69;
assign n_848 = n_821 ^ n_846;
assign n_849 = n_847 & n_848;
assign n_850 = n_849 ^ x69;
assign n_851 = n_850 ^ x70;
assign n_852 = n_822 ^ n_850;
assign n_853 = n_851 & n_852;
assign n_854 = n_853 ^ x70;
assign n_855 = n_854 ^ x71;
assign n_856 = n_823 ^ n_854;
assign n_857 = n_855 & n_856;
assign n_858 = n_857 ^ x71;
assign n_859 = n_858 ^ x72;
assign n_860 = n_824 ^ n_858;
assign n_861 = n_859 & n_860;
assign n_862 = n_861 ^ x72;
assign n_863 = n_862 ^ x73;
assign n_864 = n_825 ^ n_862;
assign n_865 = n_863 & n_864;
assign n_866 = n_865 ^ x73;
assign n_867 = n_866 ^ x74;
assign n_868 = n_826 ^ n_866;
assign n_869 = n_867 & n_868;
assign n_870 = n_869 ^ x74;
assign n_871 = x75 & n_870;
assign n_872 = n_870 ^ x75;
assign n_873 = n_394 & ~n_871;
assign n_874 = n_872 & ~n_831;
assign n_875 = n_827 & ~n_873;
assign n_876 = n_874 ^ x75;
assign n_877 = x75 ^ n_875;
assign n_878 = x75 & ~n_875;
assign n_879 = n_394 & ~n_876;
assign n_880 = n_877 ^ n_878;
assign n_881 = x64 & n_879;
assign n_882 = x52 ^ n_879;
assign n_883 = n_134 & n_879;
assign n_884 = n_834 & n_879;
assign n_885 = n_839 & n_879;
assign n_886 = n_843 & n_879;
assign n_887 = n_847 & n_879;
assign n_888 = n_851 & n_879;
assign n_889 = n_855 & n_879;
assign n_890 = n_859 & n_879;
assign n_891 = n_863 & n_879;
assign n_892 = n_867 & n_879;
assign y52 = n_879;
assign n_893 = n_880 ^ x76;
assign n_894 = n_882 ^ n_8;
assign n_895 = n_883 ^ n_805;
assign n_896 = n_884 ^ n_835;
assign n_897 = n_885 ^ n_819;
assign n_898 = n_886 ^ n_820;
assign n_899 = n_887 ^ n_821;
assign n_900 = n_888 ^ n_822;
assign n_901 = n_889 ^ n_823;
assign n_902 = n_890 ^ n_824;
assign n_903 = n_891 ^ n_825;
assign n_904 = n_892 ^ n_826;
assign n_905 = n_881 ^ n_894;
assign n_906 = n_895 ^ x53;
assign n_907 = n_905 ^ n_879;
assign n_908 = n_136 & n_907;
assign n_909 = n_908 ^ x65;
assign n_910 = n_909 ^ x66;
assign n_911 = n_906 ^ n_909;
assign n_912 = n_910 & n_911;
assign n_913 = n_912 ^ x66;
assign n_914 = n_913 ^ x67;
assign n_915 = n_896 ^ n_913;
assign n_916 = n_914 & n_915;
assign n_917 = n_916 ^ x67;
assign n_918 = n_917 ^ x68;
assign n_919 = n_897 ^ n_917;
assign n_920 = n_918 & n_919;
assign n_921 = n_920 ^ x68;
assign n_922 = n_921 ^ x69;
assign n_923 = n_898 ^ n_921;
assign n_924 = n_922 & n_923;
assign n_925 = n_924 ^ x69;
assign n_926 = n_925 ^ x70;
assign n_927 = n_899 ^ n_925;
assign n_928 = n_926 & n_927;
assign n_929 = n_928 ^ x70;
assign n_930 = n_929 ^ x71;
assign n_931 = n_900 ^ n_929;
assign n_932 = n_930 & n_931;
assign n_933 = n_932 ^ x71;
assign n_934 = n_933 ^ x72;
assign n_935 = n_901 ^ n_933;
assign n_936 = n_934 & n_935;
assign n_937 = n_936 ^ x72;
assign n_938 = n_937 ^ x73;
assign n_939 = n_902 ^ n_937;
assign n_940 = n_938 & n_939;
assign n_941 = n_940 ^ x73;
assign n_942 = n_941 ^ x74;
assign n_943 = n_903 ^ n_941;
assign n_944 = n_942 & n_943;
assign n_945 = n_944 ^ x74;
assign n_946 = n_945 ^ x75;
assign n_947 = n_904 ^ n_945;
assign n_948 = ~n_945 & n_875;
assign n_949 = n_946 & n_947;
assign n_950 = n_904 & n_948;
assign n_951 = n_949 ^ n_878;
assign n_952 = ~n_893 & ~n_951;
assign n_953 = ~n_952 & ~n_950;
assign n_954 = n_393 & ~n_953;
assign n_955 = n_875 & ~n_954;
assign n_956 = x64 & n_954;
assign n_957 = n_136 & n_954;
assign n_958 = n_910 & n_954;
assign n_959 = n_914 & n_954;
assign n_960 = n_918 & n_954;
assign n_961 = n_922 & n_954;
assign n_962 = n_926 & n_954;
assign n_963 = n_930 & n_954;
assign n_964 = n_934 & n_954;
assign n_965 = n_938 & n_954;
assign n_966 = n_942 & n_954;
assign n_967 = n_946 & n_954;
assign y51 = n_954;
assign n_968 = ~n_392 & n_955;
assign n_969 = ~n_439 ^ ~n_955;
assign n_970 = n_186 ^ n_956;
assign n_971 = n_957 ^ n_881;
assign n_972 = n_958 ^ n_906;
assign n_973 = n_959 ^ n_896;
assign n_974 = n_960 ^ n_897;
assign n_975 = n_961 ^ n_898;
assign n_976 = n_962 ^ n_899;
assign n_977 = n_963 ^ n_900;
assign n_978 = n_964 ^ n_901;
assign n_979 = n_965 ^ n_902;
assign n_980 = n_966 ^ n_903;
assign n_981 = n_967 ^ n_904;
assign n_982 = ~n_969 ^ x77;
assign n_983 = ~n_59 & n_970;
assign n_984 = n_971 ^ x52;
assign n_985 = n_983 ^ n_60;
assign n_986 = n_985 ^ n_137;
assign n_987 = n_58 ^ n_986;
assign n_988 = n_987 ^ x66;
assign n_989 = n_984 ^ n_987;
assign n_990 = n_988 & n_989;
assign n_991 = n_990 ^ x66;
assign n_992 = n_991 ^ x67;
assign n_993 = n_972 ^ n_991;
assign n_994 = n_992 & n_993;
assign n_995 = n_994 ^ x67;
assign n_996 = n_995 ^ x68;
assign n_997 = n_973 ^ n_995;
assign n_998 = n_996 & n_997;
assign n_999 = n_998 ^ x68;
assign n_1000 = n_999 ^ x69;
assign n_1001 = n_974 ^ n_999;
assign n_1002 = n_1000 & n_1001;
assign n_1003 = n_1002 ^ x69;
assign n_1004 = n_1003 ^ x70;
assign n_1005 = n_975 ^ n_1003;
assign n_1006 = n_1004 & n_1005;
assign n_1007 = n_1006 ^ x70;
assign n_1008 = n_1007 ^ x71;
assign n_1009 = n_976 ^ n_1007;
assign n_1010 = n_1008 & n_1009;
assign n_1011 = n_1010 ^ x71;
assign n_1012 = n_1011 ^ x72;
assign n_1013 = n_977 ^ n_1011;
assign n_1014 = n_1012 & n_1013;
assign n_1015 = n_1014 ^ x72;
assign n_1016 = n_1015 ^ x73;
assign n_1017 = n_978 ^ n_1015;
assign n_1018 = n_1016 & n_1017;
assign n_1019 = n_1018 ^ x73;
assign n_1020 = n_1019 ^ x74;
assign n_1021 = n_979 ^ n_1019;
assign n_1022 = n_1020 & n_1021;
assign n_1023 = n_1022 ^ x74;
assign n_1024 = n_1023 ^ x75;
assign n_1025 = n_980 ^ n_1023;
assign n_1026 = n_1024 & n_1025;
assign n_1027 = n_1026 ^ x75;
assign n_1028 = n_1027 ^ x76;
assign n_1029 = n_981 ^ n_1027;
assign n_1030 = n_1028 & ~n_1029;
assign n_1031 = n_1030 ^ n_1027;
assign n_1032 = n_1031 ^ ~n_969;
assign n_1033 = n_982 & ~n_1032;
assign n_1034 = x77 ^ n_1033;
assign n_1035 = n_392 & ~n_1034;
assign n_1036 = n_955 & ~n_1035;
assign n_1037 = n_60 & n_1035;
assign n_1038 = x50 ^ n_1035;
assign n_1039 = x65 & n_1035;
assign n_1040 = x64 & n_1035;
assign n_1041 = n_988 & n_1035;
assign n_1042 = n_992 & n_1035;
assign n_1043 = n_996 & n_1035;
assign n_1044 = n_1000 & n_1035;
assign n_1045 = n_1004 & n_1035;
assign n_1046 = n_1008 & n_1035;
assign n_1047 = n_1012 & n_1035;
assign n_1048 = n_1016 & n_1035;
assign n_1049 = n_1020 & n_1035;
assign n_1050 = n_1024 & n_1035;
assign n_1051 = n_1028 & n_1035;
assign y50 = n_1035;
assign n_1052 = ~n_439 ^ ~n_1036;
assign n_1053 = n_1038 ^ n_9;
assign n_1054 = n_1039 ^ n_956;
assign n_1055 = ~x50 & n_1040;
assign n_1056 = n_1041 ^ n_984;
assign n_1057 = n_1042 ^ n_972;
assign n_1058 = n_1043 ^ n_973;
assign n_1059 = n_1044 ^ n_974;
assign n_1060 = n_1045 ^ n_975;
assign n_1061 = n_1046 ^ n_976;
assign n_1062 = n_1047 ^ n_977;
assign n_1063 = n_1048 ^ n_978;
assign n_1064 = n_1049 ^ n_979;
assign n_1065 = n_1050 ^ n_980;
assign n_1066 = n_1051 ^ n_981;
assign n_1067 = ~n_1052 ^ x78;
assign n_1068 = n_392 & n_1052;
assign n_1069 = n_138 & n_1053;
assign n_1070 = n_1054 ^ n_1055;
assign n_1071 = n_391 & n_1067;
assign n_1072 = n_1069 ^ x65;
assign n_1073 = n_1070 ^ x51;
assign n_1074 = n_1037 ^ n_1072;
assign n_1075 = n_1074 ^ x66;
assign n_1076 = n_1073 ^ n_1074;
assign n_1077 = n_1075 & n_1076;
assign n_1078 = n_1077 ^ x66;
assign n_1079 = n_1078 ^ x67;
assign n_1080 = n_1056 ^ n_1078;
assign n_1081 = n_1079 & n_1080;
assign n_1082 = n_1081 ^ x67;
assign n_1083 = n_1082 ^ x68;
assign n_1084 = n_1057 ^ n_1082;
assign n_1085 = n_1083 & n_1084;
assign n_1086 = n_1085 ^ x68;
assign n_1087 = n_1086 ^ x69;
assign n_1088 = n_1058 ^ n_1086;
assign n_1089 = n_1087 & n_1088;
assign n_1090 = n_1089 ^ x69;
assign n_1091 = n_1090 ^ x70;
assign n_1092 = n_1059 ^ n_1090;
assign n_1093 = n_1091 & n_1092;
assign n_1094 = n_1093 ^ x70;
assign n_1095 = n_1094 ^ x71;
assign n_1096 = n_1060 ^ n_1094;
assign n_1097 = n_1095 & n_1096;
assign n_1098 = n_1097 ^ x71;
assign n_1099 = n_1098 ^ x72;
assign n_1100 = n_1061 ^ n_1098;
assign n_1101 = n_1099 & n_1100;
assign n_1102 = n_1101 ^ x72;
assign n_1103 = n_1102 ^ x73;
assign n_1104 = n_1062 ^ n_1102;
assign n_1105 = n_1103 & n_1104;
assign n_1106 = n_1105 ^ x73;
assign n_1107 = n_1106 ^ x74;
assign n_1108 = n_1063 ^ n_1106;
assign n_1109 = n_1107 & n_1108;
assign n_1110 = n_1109 ^ x74;
assign n_1111 = n_1110 ^ x75;
assign n_1112 = n_1064 ^ n_1110;
assign n_1113 = n_1111 & n_1112;
assign n_1114 = n_1113 ^ x75;
assign n_1115 = n_1114 ^ x76;
assign n_1116 = n_1065 ^ n_1114;
assign n_1117 = n_1115 & n_1116;
assign n_1118 = n_1117 ^ x76;
assign n_1119 = n_1118 ^ x77;
assign n_1120 = n_1066 ^ n_1118;
assign n_1121 = n_1119 & ~n_1120;
assign n_1122 = n_1121 ^ n_1118;
assign n_1123 = n_1071 & ~n_1122;
assign n_1124 = n_1068 ^ n_1123;
assign n_1125 = n_968 & ~n_1123;
assign n_1126 = n_1119 & n_1124;
assign n_1127 = x64 & n_1124;
assign n_1128 = n_138 & n_1124;
assign n_1129 = n_1075 & n_1124;
assign n_1130 = n_1079 & n_1124;
assign n_1131 = n_1083 & n_1124;
assign n_1132 = n_1087 & n_1124;
assign n_1133 = n_1091 & n_1124;
assign n_1134 = n_1095 & n_1124;
assign n_1135 = n_1099 & n_1124;
assign n_1136 = n_1103 & n_1124;
assign n_1137 = n_1107 & n_1124;
assign n_1138 = n_1111 & n_1124;
assign n_1139 = n_1115 & n_1124;
assign y49 = n_1124;
assign n_1140 = ~n_439 ^ ~n_1125;
assign n_1141 = n_1126 ^ n_1066;
assign n_1142 = n_1127 ^ x49;
assign n_1143 = n_1128 ^ n_1040;
assign n_1144 = n_1129 ^ n_1073;
assign n_1145 = n_1130 ^ n_1056;
assign n_1146 = n_1131 ^ n_1057;
assign n_1147 = n_1132 ^ n_1058;
assign n_1148 = n_1133 ^ n_1059;
assign n_1149 = n_1134 ^ n_1060;
assign n_1150 = n_1135 ^ n_1061;
assign n_1151 = n_1136 ^ n_1062;
assign n_1152 = n_1137 ^ n_1063;
assign n_1153 = n_1138 ^ n_1064;
assign n_1154 = n_1139 ^ n_1065;
assign n_1155 = ~x79 & n_1140;
assign n_1156 = n_390 & n_1140;
assign n_1157 = ~x78 ^ n_1141;
assign n_1158 = n_1142 ^ n_10;
assign n_1159 = n_1143 ^ x50;
assign n_1160 = x78 & ~n_1155;
assign n_1161 = ~n_391 & ~n_1156;
assign n_1162 = n_1157 & ~n_1155;
assign n_1163 = n_139 & n_1158;
assign n_1164 = ~n_1141 & n_1160;
assign n_1165 = n_1163 ^ x65;
assign n_1166 = ~n_1164 & ~n_1161;
assign n_1167 = n_1165 ^ x66;
assign n_1168 = n_1159 ^ n_1165;
assign n_1169 = n_1167 & n_1168;
assign n_1170 = n_1169 ^ x66;
assign n_1171 = n_1170 ^ x67;
assign n_1172 = n_1144 ^ n_1170;
assign n_1173 = n_1171 & n_1172;
assign n_1174 = n_1173 ^ x67;
assign n_1175 = n_1174 ^ x68;
assign n_1176 = n_1145 ^ n_1174;
assign n_1177 = n_1175 & n_1176;
assign n_1178 = n_1177 ^ x68;
assign n_1179 = n_1178 ^ x69;
assign n_1180 = n_1146 ^ n_1178;
assign n_1181 = n_1179 & n_1180;
assign n_1182 = n_1181 ^ x69;
assign n_1183 = n_1182 ^ x70;
assign n_1184 = n_1147 ^ n_1182;
assign n_1185 = n_1183 & n_1184;
assign n_1186 = n_1185 ^ x70;
assign n_1187 = n_1186 ^ x71;
assign n_1188 = n_1148 ^ n_1186;
assign n_1189 = n_1187 & n_1188;
assign n_1190 = n_1189 ^ x71;
assign n_1191 = n_1190 ^ x72;
assign n_1192 = n_1149 ^ n_1190;
assign n_1193 = n_1191 & n_1192;
assign n_1194 = n_1193 ^ x72;
assign n_1195 = n_1194 ^ x73;
assign n_1196 = n_1150 ^ n_1194;
assign n_1197 = n_1195 & n_1196;
assign n_1198 = n_1197 ^ x73;
assign n_1199 = n_1198 ^ x74;
assign n_1200 = n_1151 ^ n_1198;
assign n_1201 = n_1199 & n_1200;
assign n_1202 = n_1201 ^ x74;
assign n_1203 = n_1202 ^ x75;
assign n_1204 = n_1152 ^ n_1202;
assign n_1205 = n_1203 & n_1204;
assign n_1206 = n_1205 ^ x75;
assign n_1207 = n_1206 ^ x76;
assign n_1208 = n_1153 ^ n_1206;
assign n_1209 = n_1207 & n_1208;
assign n_1210 = n_1209 ^ x76;
assign n_1211 = n_1210 ^ x77;
assign n_1212 = n_1154 ^ n_1210;
assign n_1213 = n_1211 & n_1212;
assign n_1214 = n_1213 ^ x77;
assign n_1215 = n_1214 ^ x78;
assign n_1216 = n_1162 & n_1214;
assign n_1217 = ~n_1216 & n_1166;
assign n_1218 = n_1125 & ~n_1217;
assign n_1219 = n_1215 & n_1217;
assign n_1220 = n_1167 & n_1217;
assign n_1221 = x64 & n_1217;
assign n_1222 = n_10 & n_1217;
assign n_1223 = x65 & n_1217;
assign n_1224 = n_1171 & n_1217;
assign n_1225 = n_1175 & n_1217;
assign n_1226 = n_1179 & n_1217;
assign n_1227 = n_1183 & n_1217;
assign n_1228 = n_1187 & n_1217;
assign n_1229 = n_1191 & n_1217;
assign n_1230 = n_1195 & n_1217;
assign n_1231 = n_1199 & n_1217;
assign n_1232 = n_1203 & n_1217;
assign n_1233 = n_1207 & n_1217;
assign n_1234 = n_1211 & n_1217;
assign y48 = n_1217;
assign n_1235 = ~n_439 ^ ~n_1218;
assign n_1236 = ~n_389 & n_1218;
assign n_1237 = n_1219 ^ n_1141;
assign n_1238 = n_1220 ^ n_1159;
assign n_1239 = n_1221 ^ x48;
assign n_1240 = n_1221 ^ n_10;
assign n_1241 = n_1222 ^ n_1127;
assign n_1242 = n_1223 ^ x49;
assign n_1243 = n_1224 ^ n_1144;
assign n_1244 = n_1225 ^ n_1145;
assign n_1245 = n_1226 ^ n_1146;
assign n_1246 = n_1227 ^ n_1147;
assign n_1247 = n_1228 ^ n_1148;
assign n_1248 = n_1229 ^ n_1149;
assign n_1249 = n_1230 ^ n_1150;
assign n_1250 = n_1231 ^ n_1151;
assign n_1251 = n_1232 ^ n_1152;
assign n_1252 = n_1233 ^ n_1153;
assign n_1253 = n_1234 ^ n_1154;
assign n_1254 = ~n_1235 ^ x80;
assign n_1255 = ~n_1235 ^ x79;
assign n_1256 = x79 & ~n_1235;
assign n_1257 = x79 & ~n_1237;
assign n_1258 = n_1237 ^ x80;
assign n_1259 = n_1238 ^ x67;
assign n_1260 = x65 & ~n_1239;
assign n_1261 = n_1240 ^ n_61;
assign n_1262 = n_1241 ^ n_1242;
assign n_1263 = ~n_1237 & ~n_1255;
assign n_1264 = n_1257 ^ ~n_1235;
assign n_1265 = ~x47 & n_1261;
assign n_1266 = n_1263 ^ x79;
assign n_1267 = n_1254 & ~n_1264;
assign n_1268 = n_1260 ^ n_1265;
assign n_1269 = ~n_1258 & ~n_1266;
assign n_1270 = x80 ^ n_1267;
assign n_1271 = n_1268 ^ x66;
assign n_1272 = n_1262 ^ n_1268;
assign n_1273 = x80 ^ n_1269;
assign n_1274 = n_1271 & n_1272;
assign n_1275 = n_1273 ^ n_1256;
assign n_1276 = n_1274 ^ x66;
assign n_1277 = n_1276 ^ n_1238;
assign n_1278 = n_1276 ^ x67;
assign n_1279 = ~n_1259 & n_1277;
assign n_1280 = n_1279 ^ x67;
assign n_1281 = n_1280 ^ x68;
assign n_1282 = n_1243 ^ n_1280;
assign n_1283 = n_1281 & n_1282;
assign n_1284 = n_1283 ^ x68;
assign n_1285 = n_1284 ^ x69;
assign n_1286 = n_1244 ^ n_1284;
assign n_1287 = n_1285 & n_1286;
assign n_1288 = n_1287 ^ x69;
assign n_1289 = n_1288 ^ x70;
assign n_1290 = n_1245 ^ n_1288;
assign n_1291 = n_1289 & n_1290;
assign n_1292 = n_1291 ^ x70;
assign n_1293 = n_1292 ^ x71;
assign n_1294 = n_1246 ^ n_1292;
assign n_1295 = n_1293 & n_1294;
assign n_1296 = n_1295 ^ x71;
assign n_1297 = n_1296 ^ x72;
assign n_1298 = n_1247 ^ n_1296;
assign n_1299 = n_1297 & n_1298;
assign n_1300 = n_1299 ^ x72;
assign n_1301 = n_1300 ^ x73;
assign n_1302 = n_1248 ^ n_1300;
assign n_1303 = n_1301 & n_1302;
assign n_1304 = n_1303 ^ x73;
assign n_1305 = n_1304 ^ x74;
assign n_1306 = n_1249 ^ n_1304;
assign n_1307 = n_1305 & n_1306;
assign n_1308 = n_1307 ^ x74;
assign n_1309 = n_1308 ^ x75;
assign n_1310 = n_1250 ^ n_1308;
assign n_1311 = n_1309 & n_1310;
assign n_1312 = n_1311 ^ x75;
assign n_1313 = n_1312 ^ x76;
assign n_1314 = n_1251 ^ n_1312;
assign n_1315 = n_1313 & n_1314;
assign n_1316 = n_1315 ^ x76;
assign n_1317 = n_1316 ^ x77;
assign n_1318 = n_1252 ^ n_1316;
assign n_1319 = n_1317 & n_1318;
assign n_1320 = n_1319 ^ x77;
assign n_1321 = n_1320 ^ x78;
assign n_1322 = n_1253 ^ n_1320;
assign n_1323 = n_1321 & n_1322;
assign n_1324 = n_1323 ^ x78;
assign n_1325 = n_1324 ^ n_1256;
assign n_1326 = n_1324 ^ x79;
assign n_1327 = ~n_1256 ^ ~n_1325;
assign n_1328 = ~n_1327 ^ n_1256;
assign n_1329 = n_1275 & ~n_1328;
assign n_1330 = ~n_1327 ^ n_1329;
assign n_1331 = n_1330 ^ n_1256;
assign n_1332 = n_1331 ^ n_1324;
assign n_1333 = ~n_1270 & ~n_1332;
assign n_1334 = n_1270 ^ n_1333;
assign n_1335 = n_389 & ~n_1334;
assign n_1336 = ~n_439 ^ n_1335;
assign n_1337 = x64 & n_1335;
assign n_1338 = x65 & n_1335;
assign n_1339 = n_1271 & n_1335;
assign n_1340 = n_1278 & n_1335;
assign n_1341 = n_1281 & n_1335;
assign n_1342 = n_1285 & n_1335;
assign n_1343 = n_1289 & n_1335;
assign n_1344 = n_1293 & n_1335;
assign n_1345 = n_1297 & n_1335;
assign n_1346 = n_1301 & n_1335;
assign n_1347 = n_1305 & n_1335;
assign n_1348 = n_1309 & n_1335;
assign n_1349 = n_1313 & n_1335;
assign n_1350 = n_1317 & n_1335;
assign n_1351 = n_1321 & n_1335;
assign n_1352 = n_1326 & n_1335;
assign y47 = n_1335;
assign n_1353 = n_1235 & n_1336;
assign n_1354 = ~n_62 & n_1337;
assign n_1355 = ~x47 & n_1337;
assign n_1356 = n_1339 ^ n_1262;
assign n_1357 = n_1340 ^ n_1238;
assign n_1358 = n_1341 ^ n_1243;
assign n_1359 = n_1342 ^ n_1244;
assign n_1360 = n_1343 ^ n_1245;
assign n_1361 = n_1344 ^ n_1246;
assign n_1362 = n_1345 ^ n_1247;
assign n_1363 = n_1346 ^ n_1248;
assign n_1364 = n_1347 ^ n_1249;
assign n_1365 = n_1348 ^ n_1250;
assign n_1366 = n_1349 ^ n_1251;
assign n_1367 = n_1350 ^ n_1252;
assign n_1368 = n_1351 ^ n_1253;
assign n_1369 = n_1352 ^ n_1237;
assign n_1370 = n_1353 ^ x81;
assign n_1371 = n_389 & n_1353;
assign n_1372 = n_1354 ^ x47;
assign n_1373 = n_1338 ^ n_1355;
assign n_1374 = n_388 & ~n_1370;
assign n_1375 = n_1372 ^ x65;
assign n_1376 = n_1373 ^ n_1239;
assign n_1377 = n_1375 ^ n_1354;
assign n_1378 = ~n_1377 & ~n_140;
assign n_1379 = n_1378 ^ n_1372;
assign n_1380 = n_1379 ^ x66;
assign n_1381 = n_1376 ^ n_1379;
assign n_1382 = ~n_1380 & ~n_1381;
assign n_1383 = n_1382 ^ x66;
assign n_1384 = n_1383 ^ x67;
assign n_1385 = n_1356 ^ n_1383;
assign n_1386 = n_1384 & n_1385;
assign n_1387 = n_1386 ^ x67;
assign n_1388 = n_1387 ^ x68;
assign n_1389 = n_1357 ^ n_1387;
assign n_1390 = n_1388 & n_1389;
assign n_1391 = n_1390 ^ x68;
assign n_1392 = n_1391 ^ x69;
assign n_1393 = n_1358 ^ n_1391;
assign n_1394 = n_1392 & n_1393;
assign n_1395 = n_1394 ^ x69;
assign n_1396 = n_1395 ^ x70;
assign n_1397 = n_1359 ^ n_1395;
assign n_1398 = n_1396 & n_1397;
assign n_1399 = n_1398 ^ x70;
assign n_1400 = n_1399 ^ x71;
assign n_1401 = n_1360 ^ n_1399;
assign n_1402 = n_1400 & n_1401;
assign n_1403 = n_1402 ^ x71;
assign n_1404 = n_1403 ^ x72;
assign n_1405 = n_1361 ^ n_1403;
assign n_1406 = n_1404 & n_1405;
assign n_1407 = n_1406 ^ x72;
assign n_1408 = n_1407 ^ x73;
assign n_1409 = n_1362 ^ n_1407;
assign n_1410 = n_1408 & n_1409;
assign n_1411 = n_1410 ^ x73;
assign n_1412 = n_1411 ^ x74;
assign n_1413 = n_1363 ^ n_1411;
assign n_1414 = n_1412 & n_1413;
assign n_1415 = n_1414 ^ x74;
assign n_1416 = n_1415 ^ x75;
assign n_1417 = n_1364 ^ n_1415;
assign n_1418 = n_1416 & n_1417;
assign n_1419 = n_1418 ^ x75;
assign n_1420 = n_1419 ^ x76;
assign n_1421 = n_1365 ^ n_1419;
assign n_1422 = n_1420 & n_1421;
assign n_1423 = n_1422 ^ x76;
assign n_1424 = n_1423 ^ x77;
assign n_1425 = n_1366 ^ n_1423;
assign n_1426 = n_1424 & n_1425;
assign n_1427 = n_1426 ^ x77;
assign n_1428 = n_1427 ^ x78;
assign n_1429 = n_1367 ^ n_1427;
assign n_1430 = n_1428 & n_1429;
assign n_1431 = n_1430 ^ x78;
assign n_1432 = n_1431 ^ x79;
assign n_1433 = n_1368 ^ n_1431;
assign n_1434 = n_1432 & n_1433;
assign n_1435 = n_1434 ^ x79;
assign n_1436 = n_1435 ^ x80;
assign n_1437 = n_1369 ^ n_1435;
assign n_1438 = n_1436 & n_1437;
assign n_1439 = n_1438 ^ x80;
assign n_1440 = n_1374 & ~n_1439;
assign n_1441 = n_1371 ^ n_1440;
assign n_1442 = n_1236 & ~n_1440;
assign n_1443 = n_1388 & n_1441;
assign n_1444 = n_1384 & n_1441;
assign n_1445 = x64 & n_1441;
assign n_1446 = n_1441 ^ x46;
assign n_1447 = n_140 & n_1441;
assign n_1448 = ~n_1380 & n_1441;
assign n_1449 = n_1392 & n_1441;
assign n_1450 = n_1396 & n_1441;
assign n_1451 = n_1400 & n_1441;
assign n_1452 = n_1404 & n_1441;
assign n_1453 = n_1408 & n_1441;
assign n_1454 = n_1412 & n_1441;
assign n_1455 = n_1416 & n_1441;
assign n_1456 = n_1420 & n_1441;
assign n_1457 = n_1424 & n_1441;
assign n_1458 = n_1428 & n_1441;
assign n_1459 = n_1432 & n_1441;
assign n_1460 = n_1436 & n_1441;
assign y46 = n_1441;
assign n_1461 = ~n_439 ^ ~n_1442;
assign n_1462 = n_1443 ^ n_1357;
assign n_1463 = n_1444 ^ n_1356;
assign n_1464 = n_1446 ^ n_12;
assign n_1465 = n_1447 ^ n_1337;
assign n_1466 = n_1448 ^ n_1376;
assign n_1467 = n_1449 ^ n_1358;
assign n_1468 = n_1450 ^ n_1359;
assign n_1469 = n_1451 ^ n_1360;
assign n_1470 = n_1452 ^ n_1361;
assign n_1471 = n_1453 ^ n_1362;
assign n_1472 = n_1454 ^ n_1363;
assign n_1473 = n_1455 ^ n_1364;
assign n_1474 = n_1456 ^ n_1365;
assign n_1475 = n_1457 ^ n_1366;
assign n_1476 = n_1458 ^ n_1367;
assign n_1477 = n_1459 ^ n_1368;
assign n_1478 = n_1460 ^ n_1369;
assign n_1479 = ~n_1461 ^ x82;
assign n_1480 = ~x69 ^ n_1462;
assign n_1481 = n_1462 ^ x69;
assign n_1482 = n_1463 ^ x68;
assign n_1483 = x68 & ~n_1463;
assign n_1484 = n_1445 ^ n_1464;
assign n_1485 = n_1465 ^ x47;
assign n_1486 = n_1482 ^ n_1483;
assign n_1487 = n_1483 ^ n_1462;
assign n_1488 = n_1484 ^ n_1441;
assign n_1489 = n_1480 & ~n_1486;
assign n_1490 = ~n_1481 & n_1487;
assign n_1491 = n_141 & n_1488;
assign n_1492 = n_1490 ^ x69;
assign n_1493 = n_1491 ^ x65;
assign n_1494 = n_1493 ^ x66;
assign n_1495 = n_1485 ^ n_1493;
assign n_1496 = n_1494 & n_1495;
assign n_1497 = n_1496 ^ x66;
assign n_1498 = n_1497 ^ x67;
assign n_1499 = n_1466 ^ n_1497;
assign n_1500 = n_1498 & n_1499;
assign n_1501 = n_1500 ^ x67;
assign n_1502 = n_1501 ^ x68;
assign n_1503 = n_1501 ^ n_1463;
assign n_1504 = n_1489 & n_1501;
assign n_1505 = n_1502 & n_1503;
assign n_1506 = ~n_1492 & ~n_1504;
assign n_1507 = n_1505 ^ x68;
assign n_1508 = x70 ^ n_1506;
assign n_1509 = n_1467 ^ n_1506;
assign n_1510 = n_1507 ^ x69;
assign n_1511 = ~n_1508 & ~n_1509;
assign n_1512 = n_1511 ^ x70;
assign n_1513 = n_1512 ^ x71;
assign n_1514 = n_1468 ^ n_1512;
assign n_1515 = n_1513 & n_1514;
assign n_1516 = n_1515 ^ x71;
assign n_1517 = n_1516 ^ x72;
assign n_1518 = n_1469 ^ n_1516;
assign n_1519 = n_1517 & n_1518;
assign n_1520 = n_1519 ^ x72;
assign n_1521 = n_1520 ^ x73;
assign n_1522 = n_1470 ^ n_1520;
assign n_1523 = n_1521 & n_1522;
assign n_1524 = n_1523 ^ x73;
assign n_1525 = n_1524 ^ x74;
assign n_1526 = n_1471 ^ n_1524;
assign n_1527 = n_1525 & n_1526;
assign n_1528 = n_1527 ^ x74;
assign n_1529 = n_1528 ^ x75;
assign n_1530 = n_1472 ^ n_1528;
assign n_1531 = n_1529 & n_1530;
assign n_1532 = n_1531 ^ x75;
assign n_1533 = n_1532 ^ x76;
assign n_1534 = n_1473 ^ n_1532;
assign n_1535 = n_1533 & n_1534;
assign n_1536 = n_1535 ^ x76;
assign n_1537 = n_1536 ^ x77;
assign n_1538 = n_1474 ^ n_1536;
assign n_1539 = n_1537 & n_1538;
assign n_1540 = n_1539 ^ x77;
assign n_1541 = n_1540 ^ x78;
assign n_1542 = n_1475 ^ n_1540;
assign n_1543 = n_1541 & n_1542;
assign n_1544 = n_1543 ^ x78;
assign n_1545 = n_1544 ^ x79;
assign n_1546 = n_1476 ^ n_1544;
assign n_1547 = n_1545 & n_1546;
assign n_1548 = n_1547 ^ x79;
assign n_1549 = n_1548 ^ x80;
assign n_1550 = n_1477 ^ n_1548;
assign n_1551 = n_1549 & n_1550;
assign n_1552 = n_1551 ^ x80;
assign n_1553 = n_1552 ^ x81;
assign n_1554 = n_1478 ^ n_1552;
assign n_1555 = n_1553 & ~n_1554;
assign n_1556 = n_1555 ^ n_1552;
assign n_1557 = n_1556 ^ ~n_1461;
assign n_1558 = n_1479 & ~n_1557;
assign n_1559 = x82 ^ n_1558;
assign n_1560 = n_387 & ~n_1559;
assign n_1561 = n_1442 & ~n_1560;
assign n_1562 = x65 & n_1560;
assign n_1563 = n_12 & n_1560;
assign n_1564 = x64 & n_1560;
assign n_1565 = n_1494 & n_1560;
assign n_1566 = n_1498 & n_1560;
assign n_1567 = n_1502 & n_1560;
assign n_1568 = ~n_1508 & n_1560;
assign n_1569 = n_1513 & n_1560;
assign n_1570 = n_1517 & n_1560;
assign n_1571 = n_1521 & n_1560;
assign n_1572 = n_1525 & n_1560;
assign n_1573 = n_1529 & n_1560;
assign n_1574 = n_1533 & n_1560;
assign n_1575 = n_1537 & n_1560;
assign n_1576 = n_1541 & n_1560;
assign n_1577 = n_1545 & n_1560;
assign n_1578 = n_1549 & n_1560;
assign n_1579 = n_1553 & n_1560;
assign y45 = n_1560;
assign n_1580 = n_1510 & n_1560;
assign n_1581 = ~n_439 ^ ~n_1561;
assign n_1582 = n_64 ^ n_1562;
assign n_1583 = n_1562 ^ n_1563;
assign n_1584 = n_1564 ^ n_12;
assign n_1585 = n_1565 ^ n_1485;
assign n_1586 = n_1566 ^ n_1466;
assign n_1587 = n_1567 ^ n_1463;
assign n_1588 = n_1568 ^ n_1467;
assign n_1589 = n_1569 ^ n_1468;
assign n_1590 = n_1570 ^ n_1469;
assign n_1591 = n_1571 ^ n_1470;
assign n_1592 = n_1572 ^ n_1471;
assign n_1593 = n_1573 ^ n_1472;
assign n_1594 = n_1574 ^ n_1473;
assign n_1595 = n_1575 ^ n_1474;
assign n_1596 = n_1576 ^ n_1475;
assign n_1597 = n_1577 ^ n_1476;
assign n_1598 = n_1578 ^ n_1477;
assign n_1599 = n_1579 ^ n_1478;
assign n_1600 = n_1462 ^ n_1580;
assign n_1601 = ~n_1581 ^ x83;
assign n_1602 = x64 & n_1582;
assign n_1603 = n_1583 ^ n_1445;
assign n_1604 = ~x44 & n_1584;
assign n_1605 = n_1603 ^ x46;
assign n_1606 = n_1604 ^ n_1602;
assign n_1607 = n_1605 ^ x66;
assign n_1608 = n_63 ^ n_1606;
assign n_1609 = n_1608 ^ n_1605;
assign n_1610 = n_1608 ^ x66;
assign n_1611 = ~n_1607 & n_1609;
assign n_1612 = n_1611 ^ x66;
assign n_1613 = n_1612 ^ x67;
assign n_1614 = n_1585 ^ n_1612;
assign n_1615 = n_1613 & n_1614;
assign n_1616 = n_1615 ^ x67;
assign n_1617 = n_1616 ^ x68;
assign n_1618 = n_1586 ^ n_1616;
assign n_1619 = n_1617 & n_1618;
assign n_1620 = n_1619 ^ x68;
assign n_1621 = n_1620 ^ x69;
assign n_1622 = n_1587 ^ n_1620;
assign n_1623 = n_1621 & n_1622;
assign n_1624 = n_1623 ^ x69;
assign n_1625 = n_1624 ^ x70;
assign n_1626 = n_1600 ^ n_1624;
assign n_1627 = n_1625 & n_1626;
assign n_1628 = n_1627 ^ x70;
assign n_1629 = n_1628 ^ x71;
assign n_1630 = n_1588 ^ n_1628;
assign n_1631 = n_1629 & n_1630;
assign n_1632 = n_1631 ^ x71;
assign n_1633 = n_1632 ^ x72;
assign n_1634 = n_1589 ^ n_1632;
assign n_1635 = n_1633 & n_1634;
assign n_1636 = n_1635 ^ x72;
assign n_1637 = n_1636 ^ x73;
assign n_1638 = n_1590 ^ n_1636;
assign n_1639 = n_1637 & n_1638;
assign n_1640 = n_1639 ^ x73;
assign n_1641 = n_1640 ^ x74;
assign n_1642 = n_1591 ^ n_1640;
assign n_1643 = n_1641 & n_1642;
assign n_1644 = n_1643 ^ x74;
assign n_1645 = n_1644 ^ x75;
assign n_1646 = n_1592 ^ n_1644;
assign n_1647 = n_1645 & n_1646;
assign n_1648 = n_1647 ^ x75;
assign n_1649 = n_1648 ^ x76;
assign n_1650 = n_1593 ^ n_1648;
assign n_1651 = n_1649 & n_1650;
assign n_1652 = n_1651 ^ x76;
assign n_1653 = n_1652 ^ x77;
assign n_1654 = n_1594 ^ n_1652;
assign n_1655 = n_1653 & n_1654;
assign n_1656 = n_1655 ^ x77;
assign n_1657 = n_1656 ^ x78;
assign n_1658 = n_1595 ^ n_1656;
assign n_1659 = n_1657 & n_1658;
assign n_1660 = n_1659 ^ x78;
assign n_1661 = n_1660 ^ x79;
assign n_1662 = n_1596 ^ n_1660;
assign n_1663 = n_1661 & n_1662;
assign n_1664 = n_1663 ^ x79;
assign n_1665 = n_1664 ^ x80;
assign n_1666 = n_1597 ^ n_1664;
assign n_1667 = n_1665 & n_1666;
assign n_1668 = n_1667 ^ x80;
assign n_1669 = n_1668 ^ x81;
assign n_1670 = n_1598 ^ n_1668;
assign n_1671 = n_1669 & n_1670;
assign n_1672 = n_1671 ^ x81;
assign n_1673 = n_1672 ^ x82;
assign n_1674 = n_1599 ^ n_1672;
assign n_1675 = n_1673 & ~n_1674;
assign n_1676 = n_1675 ^ n_1672;
assign n_1677 = n_1676 ^ ~n_1581;
assign n_1678 = n_1601 & ~n_1677;
assign n_1679 = x83 ^ n_1678;
assign n_1680 = ~n_1679 & n_384;
assign n_1681 = n_1610 & n_1680;
assign n_1682 = x64 & n_1680;
assign n_1683 = x65 & n_1680;
assign n_1684 = n_1613 & n_1680;
assign n_1685 = n_1617 & n_1680;
assign n_1686 = n_1621 & n_1680;
assign n_1687 = n_1625 & n_1680;
assign n_1688 = n_1629 & n_1680;
assign n_1689 = n_1633 & n_1680;
assign n_1690 = n_1637 & n_1680;
assign n_1691 = n_1641 & n_1680;
assign n_1692 = n_1645 & n_1680;
assign n_1693 = n_1649 & n_1680;
assign n_1694 = n_1653 & n_1680;
assign n_1695 = n_1657 & n_1680;
assign n_1696 = n_1661 & n_1680;
assign n_1697 = n_1665 & n_1680;
assign n_1698 = n_1669 & n_1680;
assign n_1699 = n_1673 & n_1680;
assign n_1700 = ~n_439 ^ n_1680;
assign y44 = n_1680;
assign n_1701 = n_1681 ^ n_1605;
assign n_1702 = x65 & n_1682;
assign n_1703 = ~x43 & n_1682;
assign n_1704 = n_1682 ^ x44;
assign n_1705 = n_1684 ^ n_1585;
assign n_1706 = n_1685 ^ n_1586;
assign n_1707 = n_1686 ^ n_1587;
assign n_1708 = n_1687 ^ n_1600;
assign n_1709 = n_1688 ^ n_1588;
assign n_1710 = n_1689 ^ n_1589;
assign n_1711 = n_1690 ^ n_1590;
assign n_1712 = n_1691 ^ n_1591;
assign n_1713 = n_1692 ^ n_1592;
assign n_1714 = n_1693 ^ n_1593;
assign n_1715 = n_1694 ^ n_1594;
assign n_1716 = n_1695 ^ n_1595;
assign n_1717 = n_1696 ^ n_1596;
assign n_1718 = n_1697 ^ n_1597;
assign n_1719 = n_1698 ^ n_1598;
assign n_1720 = n_1699 ^ n_1599;
assign n_1721 = n_1581 & n_1700;
assign n_1722 = n_1701 ^ x67;
assign n_1723 = n_1702 ^ n_64;
assign n_1724 = n_1703 ^ n_142;
assign n_1725 = n_1682 & n_1704;
assign n_1726 = n_1724 ^ n_268;
assign n_1727 = n_1725 ^ n_1564;
assign n_1728 = n_1723 ^ n_1726;
assign n_1729 = n_1683 ^ n_1727;
assign n_1730 = n_1728 ^ x66;
assign n_1731 = n_1729 ^ x45;
assign n_1732 = n_1731 ^ n_1728;
assign n_1733 = n_1730 & n_1732;
assign n_1734 = n_1733 ^ x66;
assign n_1735 = n_1734 ^ n_1701;
assign n_1736 = n_1734 ^ x67;
assign n_1737 = ~n_1722 & n_1735;
assign n_1738 = n_1737 ^ x67;
assign n_1739 = n_1738 ^ x68;
assign n_1740 = n_1705 ^ n_1738;
assign n_1741 = n_1739 & n_1740;
assign n_1742 = n_1741 ^ x68;
assign n_1743 = n_1742 ^ x69;
assign n_1744 = n_1706 ^ n_1742;
assign n_1745 = n_1743 & n_1744;
assign n_1746 = n_1745 ^ x69;
assign n_1747 = n_1746 ^ x70;
assign n_1748 = n_1707 ^ n_1746;
assign n_1749 = n_1747 & n_1748;
assign n_1750 = n_1749 ^ x70;
assign n_1751 = n_1750 ^ x71;
assign n_1752 = n_1708 ^ n_1750;
assign n_1753 = n_1751 & n_1752;
assign n_1754 = n_1753 ^ x71;
assign n_1755 = n_1754 ^ x72;
assign n_1756 = n_1709 ^ n_1754;
assign n_1757 = n_1755 & n_1756;
assign n_1758 = n_1757 ^ x72;
assign n_1759 = n_1758 ^ x73;
assign n_1760 = n_1710 ^ n_1758;
assign n_1761 = n_1759 & n_1760;
assign n_1762 = n_1761 ^ x73;
assign n_1763 = n_1762 ^ x74;
assign n_1764 = n_1711 ^ n_1762;
assign n_1765 = n_1763 & n_1764;
assign n_1766 = n_1765 ^ x74;
assign n_1767 = n_1766 ^ x75;
assign n_1768 = n_1712 ^ n_1766;
assign n_1769 = n_1767 & n_1768;
assign n_1770 = n_1769 ^ x75;
assign n_1771 = n_1770 ^ x76;
assign n_1772 = n_1713 ^ n_1770;
assign n_1773 = n_1771 & n_1772;
assign n_1774 = n_1773 ^ x76;
assign n_1775 = n_1774 ^ x77;
assign n_1776 = n_1714 ^ n_1774;
assign n_1777 = n_1775 & n_1776;
assign n_1778 = n_1777 ^ x77;
assign n_1779 = n_1778 ^ x78;
assign n_1780 = n_1715 ^ n_1778;
assign n_1781 = n_1779 & n_1780;
assign n_1782 = n_1781 ^ x78;
assign n_1783 = n_1782 ^ x79;
assign n_1784 = n_1716 ^ n_1782;
assign n_1785 = n_1783 & n_1784;
assign n_1786 = n_1785 ^ x79;
assign n_1787 = n_1786 ^ x80;
assign n_1788 = n_1717 ^ n_1786;
assign n_1789 = n_1787 & n_1788;
assign n_1790 = n_1789 ^ x80;
assign n_1791 = n_1790 ^ x81;
assign n_1792 = n_1718 ^ n_1790;
assign n_1793 = n_1791 & n_1792;
assign n_1794 = n_1793 ^ x81;
assign n_1795 = n_1794 ^ x82;
assign n_1796 = n_1719 ^ n_1794;
assign n_1797 = n_1795 & n_1796;
assign n_1798 = n_1797 ^ x82;
assign n_1799 = n_1798 ^ x83;
assign n_1800 = n_1720 ^ n_1798;
assign n_1801 = n_1799 & n_1800;
assign n_1802 = n_1801 ^ x83;
assign n_1803 = n_1802 ^ x84;
assign n_1804 = n_1721 ^ n_1802;
assign n_1805 = x84 & n_1802;
assign n_1806 = n_1803 & n_1804;
assign n_1807 = n_385 & ~n_1805;
assign n_1808 = n_1806 ^ x84;
assign n_1809 = n_1721 & ~n_1807;
assign n_1810 = n_385 & ~n_1808;
assign n_1811 = n_1721 ^ n_1809;
assign n_1812 = x64 & n_1810;
assign n_1813 = n_1767 & n_1810;
assign n_1814 = n_1763 & n_1810;
assign n_1815 = n_143 & n_1810;
assign n_1816 = x65 ^ n_1810;
assign n_1817 = n_1730 & n_1810;
assign n_1818 = n_1736 & n_1810;
assign n_1819 = n_1739 & n_1810;
assign n_1820 = n_1743 & n_1810;
assign n_1821 = n_1747 & n_1810;
assign n_1822 = n_1751 & n_1810;
assign n_1823 = n_1755 & n_1810;
assign n_1824 = n_1759 & n_1810;
assign n_1825 = n_1771 & n_1810;
assign n_1826 = n_1775 & n_1810;
assign n_1827 = n_1779 & n_1810;
assign n_1828 = n_1783 & n_1810;
assign n_1829 = n_1787 & n_1810;
assign n_1830 = n_1791 & n_1810;
assign n_1831 = n_1795 & n_1810;
assign n_1832 = n_1799 & n_1810;
assign y43 = n_1810;
assign n_1833 = n_4 ^ n_1812;
assign n_1834 = ~n_1812 & n_4;
assign n_1835 = n_1813 ^ n_1712;
assign n_1836 = n_1814 ^ n_1711;
assign n_1837 = n_1815 ^ n_1704;
assign n_1838 = n_1812 & n_1816;
assign n_1839 = n_1817 ^ n_1731;
assign n_1840 = n_1818 ^ n_1701;
assign n_1841 = n_1819 ^ n_1705;
assign n_1842 = n_1820 ^ n_1706;
assign n_1843 = n_1821 ^ n_1707;
assign n_1844 = n_1822 ^ n_1708;
assign n_1845 = n_1823 ^ n_1709;
assign n_1846 = n_1824 ^ n_1710;
assign n_1847 = n_1825 ^ n_1713;
assign n_1848 = n_1826 ^ n_1714;
assign n_1849 = n_1827 ^ n_1715;
assign n_1850 = n_1828 ^ n_1716;
assign n_1851 = n_1829 ^ n_1717;
assign n_1852 = n_1830 ^ n_1718;
assign n_1853 = n_1831 ^ n_1719;
assign n_1854 = n_1832 ^ n_1720;
assign n_1855 = n_1833 ^ n_1834;
assign n_1856 = n_1835 ^ x76;
assign n_1857 = n_1836 ^ x75;
assign n_1858 = n_1837 ^ x66;
assign n_1859 = n_1855 ^ x43;
assign n_1860 = n_1855 ^ n_250;
assign n_1861 = n_1860 ^ n_1838;
assign n_1862 = n_1861 ^ n_194;
assign n_1863 = n_1862 ^ n_1837;
assign n_1864 = n_1862 ^ x66;
assign n_1865 = ~n_1858 & ~n_1863;
assign n_1866 = n_1865 ^ x66;
assign n_1867 = n_1866 ^ x67;
assign n_1868 = n_1839 ^ n_1866;
assign n_1869 = n_1867 & n_1868;
assign n_1870 = n_1869 ^ x67;
assign n_1871 = n_1870 ^ x68;
assign n_1872 = n_1840 ^ n_1870;
assign n_1873 = n_1871 & n_1872;
assign n_1874 = n_1873 ^ x68;
assign n_1875 = n_1874 ^ x69;
assign n_1876 = n_1841 ^ n_1874;
assign n_1877 = n_1875 & n_1876;
assign n_1878 = n_1877 ^ x69;
assign n_1879 = n_1878 ^ x70;
assign n_1880 = n_1842 ^ n_1878;
assign n_1881 = n_1879 & n_1880;
assign n_1882 = n_1881 ^ x70;
assign n_1883 = n_1882 ^ x71;
assign n_1884 = n_1843 ^ n_1882;
assign n_1885 = n_1883 & n_1884;
assign n_1886 = n_1885 ^ x71;
assign n_1887 = n_1886 ^ x72;
assign n_1888 = n_1844 ^ n_1886;
assign n_1889 = n_1887 & n_1888;
assign n_1890 = n_1889 ^ x72;
assign n_1891 = n_1890 ^ x73;
assign n_1892 = n_1845 ^ n_1890;
assign n_1893 = n_1891 & n_1892;
assign n_1894 = n_1893 ^ x73;
assign n_1895 = n_1894 ^ x74;
assign n_1896 = n_1846 ^ n_1894;
assign n_1897 = n_1895 & n_1896;
assign n_1898 = n_1897 ^ x74;
assign n_1899 = n_1898 ^ n_1836;
assign n_1900 = n_1898 ^ x75;
assign n_1901 = ~n_1857 & n_1899;
assign n_1902 = n_1901 ^ x75;
assign n_1903 = n_1902 ^ n_1835;
assign n_1904 = n_1902 ^ x76;
assign n_1905 = ~n_1856 & n_1903;
assign n_1906 = n_1905 ^ x76;
assign n_1907 = n_1906 ^ x77;
assign n_1908 = n_1847 ^ n_1906;
assign n_1909 = n_1907 & n_1908;
assign n_1910 = n_1909 ^ x77;
assign n_1911 = n_1910 ^ x78;
assign n_1912 = n_1848 ^ n_1910;
assign n_1913 = n_1911 & n_1912;
assign n_1914 = n_1913 ^ x78;
assign n_1915 = n_1914 ^ x79;
assign n_1916 = n_1849 ^ n_1914;
assign n_1917 = n_1915 & n_1916;
assign n_1918 = n_1917 ^ x79;
assign n_1919 = n_1918 ^ x80;
assign n_1920 = n_1850 ^ n_1918;
assign n_1921 = n_1919 & n_1920;
assign n_1922 = n_1921 ^ x80;
assign n_1923 = n_1922 ^ x81;
assign n_1924 = n_1851 ^ n_1922;
assign n_1925 = n_1923 & n_1924;
assign n_1926 = n_1925 ^ x81;
assign n_1927 = n_1926 ^ x82;
assign n_1928 = n_1852 ^ n_1926;
assign n_1929 = n_1927 & n_1928;
assign n_1930 = n_1929 ^ x82;
assign n_1931 = n_1930 ^ x83;
assign n_1932 = n_1853 ^ n_1930;
assign n_1933 = n_1931 & n_1932;
assign n_1934 = n_1933 ^ x83;
assign n_1935 = n_1934 ^ x84;
assign n_1936 = n_1854 ^ n_1934;
assign n_1937 = n_1935 & n_1936;
assign n_1938 = n_1937 ^ x84;
assign n_1939 = n_1938 ^ x85;
assign n_1940 = n_1938 ^ ~n_1811;
assign n_1941 = ~n_1940 ^ n_1721;
assign n_1942 = n_1939 & n_1941;
assign n_1943 = n_1942 ^ x85;
assign n_1944 = ~n_1943 & n_386;
assign n_1945 = n_133 & ~n_1944;
assign n_1946 = x64 & n_1944;
assign n_1947 = ~n_1864 & n_1944;
assign n_1948 = n_1919 & n_1944;
assign n_1949 = n_1915 & n_1944;
assign n_1950 = n_1867 & n_1944;
assign n_1951 = n_1871 & n_1944;
assign n_1952 = n_1875 & n_1944;
assign n_1953 = n_1879 & n_1944;
assign n_1954 = n_1883 & n_1944;
assign n_1955 = n_1887 & n_1944;
assign n_1956 = n_1891 & n_1944;
assign n_1957 = n_1895 & n_1944;
assign n_1958 = n_1900 & n_1944;
assign n_1959 = n_1904 & n_1944;
assign n_1960 = n_1907 & n_1944;
assign n_1961 = n_1911 & n_1944;
assign n_1962 = n_1923 & n_1944;
assign n_1963 = n_1927 & n_1944;
assign n_1964 = n_1931 & n_1944;
assign n_1965 = n_1935 & n_1944;
assign n_1966 = n_1809 & ~n_1944;
assign y42 = n_1944;
assign n_1967 = n_1945 ^ x65;
assign n_1968 = n_1946 ^ x42;
assign n_1969 = n_1946 ^ n_4;
assign n_1970 = n_1947 ^ n_1837;
assign n_1971 = n_1948 ^ n_1850;
assign n_1972 = n_1949 ^ n_1849;
assign n_1973 = n_1950 ^ n_1839;
assign n_1974 = n_1951 ^ n_1840;
assign n_1975 = n_1952 ^ n_1841;
assign n_1976 = n_1953 ^ n_1842;
assign n_1977 = n_1954 ^ n_1843;
assign n_1978 = n_1955 ^ n_1844;
assign n_1979 = n_1956 ^ n_1845;
assign n_1980 = n_1957 ^ n_1846;
assign n_1981 = n_1958 ^ n_1836;
assign n_1982 = n_1959 ^ n_1835;
assign n_1983 = n_1960 ^ n_1847;
assign n_1984 = n_1961 ^ n_1848;
assign n_1985 = n_1962 ^ n_1851;
assign n_1986 = n_1963 ^ n_1852;
assign n_1987 = n_1964 ^ n_1853;
assign n_1988 = n_1965 ^ n_1854;
assign n_1989 = ~n_439 ^ ~n_1966;
assign n_1990 = n_1967 ^ n_1834;
assign n_1991 = ~x65 & ~n_1968;
assign n_1992 = x41 & n_1969;
assign n_1993 = n_1971 ^ x81;
assign n_1994 = n_1972 ^ x80;
assign n_1995 = n_1987 ^ x84;
assign n_1996 = ~x84 & n_1987;
assign n_1997 = n_1988 ^ x85;
assign n_1998 = x85 & ~n_1988;
assign n_1999 = x86 ^ ~n_1989;
assign n_2000 = n_386 & n_1989;
assign n_2001 = n_1859 ^ n_1990;
assign n_2002 = n_1991 ^ x42;
assign n_2003 = n_1992 ^ n_4;
assign n_2004 = n_1995 ^ n_1996;
assign n_2005 = n_1997 ^ n_1998;
assign n_2006 = n_383 & n_1999;
assign n_2007 = n_2001 ^ x66;
assign n_2008 = n_2003 ^ n_195;
assign n_2009 = ~n_1996 & ~n_2005;
assign n_2010 = ~n_1998 & n_2006;
assign n_2011 = n_2002 ^ n_2008;
assign n_2012 = n_2011 ^ n_2001;
assign n_2013 = n_2011 ^ x66;
assign n_2014 = ~n_2007 & ~n_2012;
assign n_2015 = n_2014 ^ x66;
assign n_2016 = n_2015 ^ x67;
assign n_2017 = n_1970 ^ n_2015;
assign n_2018 = n_2016 & n_2017;
assign n_2019 = n_2018 ^ x67;
assign n_2020 = n_2019 ^ x68;
assign n_2021 = n_1973 ^ n_2019;
assign n_2022 = n_2020 & n_2021;
assign n_2023 = n_2022 ^ x68;
assign n_2024 = n_2023 ^ x69;
assign n_2025 = n_1974 ^ n_2023;
assign n_2026 = n_2024 & n_2025;
assign n_2027 = n_2026 ^ x69;
assign n_2028 = n_2027 ^ x70;
assign n_2029 = n_1975 ^ n_2027;
assign n_2030 = n_2028 & n_2029;
assign n_2031 = n_2030 ^ x70;
assign n_2032 = n_2031 ^ x71;
assign n_2033 = n_1976 ^ n_2031;
assign n_2034 = n_2032 & n_2033;
assign n_2035 = n_2034 ^ x71;
assign n_2036 = n_2035 ^ x72;
assign n_2037 = n_1977 ^ n_2035;
assign n_2038 = n_2036 & n_2037;
assign n_2039 = n_2038 ^ x72;
assign n_2040 = n_2039 ^ x73;
assign n_2041 = n_1978 ^ n_2039;
assign n_2042 = n_2040 & n_2041;
assign n_2043 = n_2042 ^ x73;
assign n_2044 = n_2043 ^ x74;
assign n_2045 = n_1979 ^ n_2043;
assign n_2046 = n_2044 & n_2045;
assign n_2047 = n_2046 ^ x74;
assign n_2048 = n_2047 ^ x75;
assign n_2049 = n_1980 ^ n_2047;
assign n_2050 = n_2048 & n_2049;
assign n_2051 = n_2050 ^ x75;
assign n_2052 = n_2051 ^ x76;
assign n_2053 = n_1981 ^ n_2051;
assign n_2054 = n_2052 & n_2053;
assign n_2055 = n_2054 ^ x76;
assign n_2056 = n_2055 ^ x77;
assign n_2057 = n_1982 ^ n_2055;
assign n_2058 = n_2056 & n_2057;
assign n_2059 = n_2058 ^ x77;
assign n_2060 = n_2059 ^ x78;
assign n_2061 = n_1983 ^ n_2059;
assign n_2062 = n_2060 & n_2061;
assign n_2063 = n_2062 ^ x78;
assign n_2064 = n_2063 ^ x79;
assign n_2065 = n_1984 ^ n_2063;
assign n_2066 = n_2064 & n_2065;
assign n_2067 = n_2066 ^ x79;
assign n_2068 = n_2067 ^ n_1972;
assign n_2069 = n_2067 ^ x80;
assign n_2070 = ~n_1994 & n_2068;
assign n_2071 = n_2070 ^ x80;
assign n_2072 = n_2071 ^ n_1971;
assign n_2073 = n_2071 ^ x81;
assign n_2074 = ~n_1993 & n_2072;
assign n_2075 = n_2074 ^ x81;
assign n_2076 = n_2075 ^ x82;
assign n_2077 = n_1985 ^ n_2075;
assign n_2078 = n_2076 & n_2077;
assign n_2079 = n_2078 ^ x82;
assign n_2080 = n_2079 ^ x83;
assign n_2081 = n_1986 ^ n_2079;
assign n_2082 = n_2080 & n_2081;
assign n_2083 = n_2082 ^ x83;
assign n_2084 = ~n_2083 & ~n_2004;
assign n_2085 = n_2083 ^ x84;
assign n_2086 = ~n_1996 & ~n_2084;
assign n_2087 = ~n_2084 & n_2009;
assign n_2088 = n_2086 ^ x85;
assign n_2089 = ~n_2087 & n_2010;
assign n_2090 = ~n_2000 ^ ~n_2089;
assign n_2091 = n_2020 & n_2090;
assign n_2092 = n_2016 & n_2090;
assign n_2093 = x65 & ~n_2090;
assign n_2094 = x64 & n_2090;
assign n_2095 = n_2090 & ~n_2013;
assign n_2096 = n_2024 & n_2090;
assign n_2097 = n_2028 & n_2090;
assign n_2098 = n_2032 & n_2090;
assign n_2099 = n_2036 & n_2090;
assign n_2100 = n_2040 & n_2090;
assign n_2101 = n_2044 & n_2090;
assign n_2102 = n_2048 & n_2090;
assign n_2103 = n_2052 & n_2090;
assign n_2104 = n_2056 & n_2090;
assign n_2105 = n_2060 & n_2090;
assign n_2106 = n_2064 & n_2090;
assign n_2107 = n_2090 & n_2069;
assign n_2108 = n_2090 & n_2073;
assign n_2109 = n_2076 & n_2090;
assign n_2110 = n_2080 & n_2090;
assign n_2111 = n_2090 & n_2085;
assign n_2112 = ~n_439 ^ n_2090;
assign y41 = n_2090;
assign n_2113 = n_2090 & n_2088;
assign n_2114 = n_2091 ^ n_1973;
assign n_2115 = n_2092 ^ n_1970;
assign n_2116 = n_196 ^ n_2093;
assign n_2117 = ~x41 & n_2094;
assign n_2118 = n_2094 ^ x41;
assign n_2119 = n_2095 ^ n_2001;
assign n_2120 = n_2096 ^ n_1974;
assign n_2121 = n_2097 ^ n_1975;
assign n_2122 = n_2098 ^ n_1976;
assign n_2123 = n_2099 ^ n_1977;
assign n_2124 = n_2100 ^ n_1978;
assign n_2125 = n_2101 ^ n_1979;
assign n_2126 = n_2102 ^ n_1980;
assign n_2127 = n_2103 ^ n_1981;
assign n_2128 = n_2104 ^ n_1982;
assign n_2129 = n_2105 ^ n_1983;
assign n_2130 = n_2106 ^ n_1984;
assign n_2131 = n_2107 ^ n_1972;
assign n_2132 = n_2108 ^ n_1971;
assign n_2133 = n_2109 ^ n_1985;
assign n_2134 = n_2110 ^ n_1986;
assign n_2135 = n_2111 ^ n_1987;
assign n_2136 = n_1989 & n_2112;
assign n_2137 = n_1988 ^ n_2113;
assign n_2138 = n_2114 ^ x69;
assign n_2139 = n_2115 ^ x68;
assign n_2140 = n_2116 ^ n_2117;
assign n_2141 = n_144 & ~n_2118;
assign n_2142 = ~n_383 & n_2136;
assign n_2143 = x88 & ~n_2136;
assign n_2144 = n_2140 ^ n_1946;
assign n_2145 = n_198 ^ n_2141;
assign n_2146 = n_381 & ~n_2143;
assign n_2147 = n_2144 ^ n_197;
assign n_2148 = n_2145 ^ x66;
assign n_2149 = n_2147 ^ x66;
assign n_2150 = n_2145 ^ n_2147;
assign n_2151 = ~n_2149 & n_2150;
assign n_2152 = n_2151 ^ x66;
assign n_2153 = n_2152 ^ x67;
assign n_2154 = n_2119 ^ n_2152;
assign n_2155 = n_2153 & n_2154;
assign n_2156 = n_2155 ^ x67;
assign n_2157 = n_2156 ^ n_2115;
assign n_2158 = n_2156 ^ x68;
assign n_2159 = ~n_2139 & n_2157;
assign n_2160 = n_2159 ^ x68;
assign n_2161 = n_2160 ^ n_2114;
assign n_2162 = n_2160 ^ n_2138;
assign n_2163 = ~n_2138 & n_2161;
assign n_2164 = n_2162 ^ n_2114;
assign n_2165 = n_2163 ^ x69;
assign n_2166 = n_2165 ^ x70;
assign n_2167 = n_2120 ^ n_2165;
assign n_2168 = n_2166 & n_2167;
assign n_2169 = n_2168 ^ x70;
assign n_2170 = n_2169 ^ x71;
assign n_2171 = n_2121 ^ n_2169;
assign n_2172 = n_2170 & n_2171;
assign n_2173 = n_2172 ^ x71;
assign n_2174 = n_2173 ^ x72;
assign n_2175 = n_2122 ^ n_2173;
assign n_2176 = n_2174 & n_2175;
assign n_2177 = n_2176 ^ x72;
assign n_2178 = n_2177 ^ x73;
assign n_2179 = n_2123 ^ n_2177;
assign n_2180 = n_2178 & n_2179;
assign n_2181 = n_2180 ^ x73;
assign n_2182 = n_2181 ^ x74;
assign n_2183 = n_2124 ^ n_2181;
assign n_2184 = n_2182 & n_2183;
assign n_2185 = n_2184 ^ x74;
assign n_2186 = n_2185 ^ x75;
assign n_2187 = n_2125 ^ n_2185;
assign n_2188 = n_2186 & n_2187;
assign n_2189 = n_2188 ^ x75;
assign n_2190 = n_2189 ^ x76;
assign n_2191 = n_2126 ^ n_2189;
assign n_2192 = n_2190 & n_2191;
assign n_2193 = n_2192 ^ x76;
assign n_2194 = n_2193 ^ x77;
assign n_2195 = n_2127 ^ n_2193;
assign n_2196 = n_2194 & n_2195;
assign n_2197 = n_2196 ^ x77;
assign n_2198 = n_2197 ^ x78;
assign n_2199 = n_2128 ^ n_2197;
assign n_2200 = n_2198 & n_2199;
assign n_2201 = n_2200 ^ x78;
assign n_2202 = n_2201 ^ x79;
assign n_2203 = n_2129 ^ n_2201;
assign n_2204 = n_2202 & n_2203;
assign n_2205 = n_2204 ^ x79;
assign n_2206 = n_2205 ^ x80;
assign n_2207 = n_2130 ^ n_2205;
assign n_2208 = n_2206 & n_2207;
assign n_2209 = n_2208 ^ x80;
assign n_2210 = n_2209 ^ x81;
assign n_2211 = n_2131 ^ n_2209;
assign n_2212 = n_2210 & n_2211;
assign n_2213 = n_2212 ^ x81;
assign n_2214 = n_2213 ^ x82;
assign n_2215 = n_2132 ^ n_2213;
assign n_2216 = n_2214 & n_2215;
assign n_2217 = n_2216 ^ x82;
assign n_2218 = n_2217 ^ x83;
assign n_2219 = n_2133 ^ n_2217;
assign n_2220 = n_2218 & n_2219;
assign n_2221 = n_2220 ^ x83;
assign n_2222 = n_2221 ^ x84;
assign n_2223 = n_2134 ^ n_2221;
assign n_2224 = n_2222 & n_2223;
assign n_2225 = n_2224 ^ x84;
assign n_2226 = n_2225 ^ x85;
assign n_2227 = n_2135 ^ n_2225;
assign n_2228 = n_2226 & n_2227;
assign n_2229 = n_2228 ^ x85;
assign n_2230 = n_2229 ^ x86;
assign n_2231 = n_2137 ^ n_2229;
assign n_2232 = n_2230 & n_2231;
assign n_2233 = n_2232 ^ x86;
assign n_2234 = n_382 & ~n_2233;
assign n_2235 = n_2233 ^ x87;
assign n_2236 = n_2136 ^ n_2233;
assign n_2237 = ~n_2234 & n_2142;
assign n_2238 = n_2235 & n_2236;
assign n_2239 = ~x88 ^ n_2237;
assign n_2240 = n_2238 ^ x87;
assign n_2241 = n_382 & ~n_2240;
assign n_2242 = n_2178 & n_2241;
assign n_2243 = n_2174 & n_2241;
assign n_2244 = n_144 & n_2241;
assign n_2245 = x64 & n_2241;
assign n_2246 = n_2148 & n_2241;
assign n_2247 = n_2153 & n_2241;
assign n_2248 = n_2158 & n_2241;
assign n_2249 = n_2164 & n_2241;
assign n_2250 = n_2166 & n_2241;
assign n_2251 = n_2170 & n_2241;
assign n_2252 = n_2182 & n_2241;
assign n_2253 = n_2186 & n_2241;
assign n_2254 = n_2190 & n_2241;
assign n_2255 = n_2194 & n_2241;
assign n_2256 = n_2198 & n_2241;
assign n_2257 = n_2202 & n_2241;
assign n_2258 = n_2206 & n_2241;
assign n_2259 = n_2210 & n_2241;
assign n_2260 = n_2214 & n_2241;
assign n_2261 = n_2218 & n_2241;
assign n_2262 = n_2222 & n_2241;
assign n_2263 = n_2226 & n_2241;
assign n_2264 = n_2230 & n_2241;
assign y40 = n_2241;
assign n_2265 = n_2242 ^ n_2123;
assign n_2266 = n_2243 ^ n_2122;
assign n_2267 = n_2244 ^ n_2094;
assign n_2268 = ~n_69 & n_2245;
assign n_2269 = n_2246 ^ n_2147;
assign n_2270 = n_2247 ^ n_2119;
assign n_2271 = n_2248 ^ n_2115;
assign n_2272 = n_2249 ^ n_2114;
assign n_2273 = n_2250 ^ n_2120;
assign n_2274 = n_2251 ^ n_2121;
assign n_2275 = n_2252 ^ n_2124;
assign n_2276 = n_2253 ^ n_2125;
assign n_2277 = n_2254 ^ n_2126;
assign n_2278 = n_2255 ^ n_2127;
assign n_2279 = n_2256 ^ n_2128;
assign n_2280 = n_2257 ^ n_2129;
assign n_2281 = n_2258 ^ n_2130;
assign n_2282 = n_2259 ^ n_2131;
assign n_2283 = n_2260 ^ n_2132;
assign n_2284 = n_2261 ^ n_2133;
assign n_2285 = n_2262 ^ n_2134;
assign n_2286 = n_2263 ^ n_2135;
assign n_2287 = n_2264 ^ n_2137;
assign n_2288 = n_2265 ^ x74;
assign n_2289 = n_2266 ^ x73;
assign n_2290 = n_2267 ^ x41;
assign n_2291 = n_2268 ^ n_269;
assign n_2292 = n_2290 ^ x66;
assign n_2293 = n_270 ^ n_2291;
assign n_2294 = n_2293 ^ n_2290;
assign n_2295 = n_2293 ^ x66;
assign n_2296 = ~n_2292 & n_2294;
assign n_2297 = n_2296 ^ x66;
assign n_2298 = n_2297 ^ x67;
assign n_2299 = n_2269 ^ n_2297;
assign n_2300 = n_2298 & n_2299;
assign n_2301 = n_2300 ^ x67;
assign n_2302 = n_2301 ^ x68;
assign n_2303 = n_2270 ^ n_2301;
assign n_2304 = n_2302 & n_2303;
assign n_2305 = n_2304 ^ x68;
assign n_2306 = n_2305 ^ x69;
assign n_2307 = n_2271 ^ n_2305;
assign n_2308 = n_2306 & n_2307;
assign n_2309 = n_2308 ^ x69;
assign n_2310 = n_2309 ^ x70;
assign n_2311 = n_2272 ^ n_2309;
assign n_2312 = n_2310 & n_2311;
assign n_2313 = n_2312 ^ x70;
assign n_2314 = n_2313 ^ x71;
assign n_2315 = n_2273 ^ n_2313;
assign n_2316 = n_2314 & n_2315;
assign n_2317 = n_2316 ^ x71;
assign n_2318 = n_2317 ^ x72;
assign n_2319 = n_2274 ^ n_2317;
assign n_2320 = n_2318 & n_2319;
assign n_2321 = n_2320 ^ x72;
assign n_2322 = n_2321 ^ n_2266;
assign n_2323 = n_2321 ^ x73;
assign n_2324 = ~n_2289 & n_2322;
assign n_2325 = n_2324 ^ x73;
assign n_2326 = n_2325 ^ n_2265;
assign n_2327 = n_2325 ^ x74;
assign n_2328 = ~n_2288 & n_2326;
assign n_2329 = n_2328 ^ x74;
assign n_2330 = n_2329 ^ x75;
assign n_2331 = n_2275 ^ n_2329;
assign n_2332 = n_2330 & n_2331;
assign n_2333 = n_2332 ^ x75;
assign n_2334 = n_2333 ^ x76;
assign n_2335 = n_2276 ^ n_2333;
assign n_2336 = n_2334 & n_2335;
assign n_2337 = n_2336 ^ x76;
assign n_2338 = n_2337 ^ x77;
assign n_2339 = n_2277 ^ n_2337;
assign n_2340 = n_2338 & n_2339;
assign n_2341 = n_2340 ^ x77;
assign n_2342 = n_2341 ^ x78;
assign n_2343 = n_2278 ^ n_2341;
assign n_2344 = n_2342 & n_2343;
assign n_2345 = n_2344 ^ x78;
assign n_2346 = n_2345 ^ x79;
assign n_2347 = n_2279 ^ n_2345;
assign n_2348 = n_2346 & n_2347;
assign n_2349 = n_2348 ^ x79;
assign n_2350 = n_2349 ^ x80;
assign n_2351 = n_2280 ^ n_2349;
assign n_2352 = n_2350 & n_2351;
assign n_2353 = n_2352 ^ x80;
assign n_2354 = n_2353 ^ x81;
assign n_2355 = n_2281 ^ n_2353;
assign n_2356 = n_2354 & n_2355;
assign n_2357 = n_2356 ^ x81;
assign n_2358 = n_2357 ^ x82;
assign n_2359 = n_2282 ^ n_2357;
assign n_2360 = n_2358 & n_2359;
assign n_2361 = n_2360 ^ x82;
assign n_2362 = n_2361 ^ x83;
assign n_2363 = n_2283 ^ n_2361;
assign n_2364 = n_2362 & n_2363;
assign n_2365 = n_2364 ^ x83;
assign n_2366 = n_2365 ^ x84;
assign n_2367 = n_2284 ^ n_2365;
assign n_2368 = n_2366 & n_2367;
assign n_2369 = n_2368 ^ x84;
assign n_2370 = n_2369 ^ x85;
assign n_2371 = n_2285 ^ n_2369;
assign n_2372 = n_2370 & n_2371;
assign n_2373 = n_2372 ^ x85;
assign n_2374 = n_2373 ^ x86;
assign n_2375 = n_2286 ^ n_2373;
assign n_2376 = n_2374 & n_2375;
assign n_2377 = n_2376 ^ x86;
assign n_2378 = n_2377 ^ x87;
assign n_2379 = n_2287 ^ n_2377;
assign n_2380 = n_2378 & ~n_2379;
assign n_2381 = n_2380 ^ n_2377;
assign n_2382 = n_2239 & n_2381;
assign n_2383 = n_2146 & ~n_2382;
assign n_2384 = n_2237 & ~n_2383;
assign n_2385 = x65 & n_2383;
assign n_2386 = x64 & n_2383;
assign n_2387 = ~x38 & ~n_2383;
assign n_2388 = n_2295 & n_2383;
assign n_2389 = n_2298 & n_2383;
assign n_2390 = n_2302 & n_2383;
assign n_2391 = n_2306 & n_2383;
assign n_2392 = n_2378 & n_2383;
assign n_2393 = n_2374 & n_2383;
assign n_2394 = n_2310 & n_2383;
assign n_2395 = n_2314 & n_2383;
assign n_2396 = n_2318 & n_2383;
assign n_2397 = n_2323 & n_2383;
assign n_2398 = n_2327 & n_2383;
assign n_2399 = n_2330 & n_2383;
assign n_2400 = n_2334 & n_2383;
assign n_2401 = n_2338 & n_2383;
assign n_2402 = n_2342 & n_2383;
assign n_2403 = n_2346 & n_2383;
assign n_2404 = n_2350 & n_2383;
assign n_2405 = n_2354 & n_2383;
assign n_2406 = n_2358 & n_2383;
assign n_2407 = n_2362 & n_2383;
assign n_2408 = n_2366 & n_2383;
assign n_2409 = n_2370 & n_2383;
assign y39 = n_2383;
assign n_2410 = ~n_439 ^ ~n_2384;
assign n_2411 = ~x39 & n_2386;
assign n_2412 = n_2386 & n_321;
assign n_2413 = ~n_2387 & ~n_70;
assign n_2414 = n_2388 ^ n_2290;
assign n_2415 = n_2389 ^ n_2269;
assign n_2416 = n_2390 ^ n_2270;
assign n_2417 = n_2391 ^ n_2271;
assign n_2418 = n_2392 ^ n_2287;
assign n_2419 = n_2393 ^ n_2286;
assign n_2420 = n_2394 ^ n_2272;
assign n_2421 = n_2395 ^ n_2273;
assign n_2422 = n_2396 ^ n_2274;
assign n_2423 = n_2397 ^ n_2266;
assign n_2424 = n_2398 ^ n_2265;
assign n_2425 = n_2399 ^ n_2275;
assign n_2426 = n_2400 ^ n_2276;
assign n_2427 = n_2401 ^ n_2277;
assign n_2428 = n_2402 ^ n_2278;
assign n_2429 = n_2403 ^ n_2279;
assign n_2430 = n_2404 ^ n_2280;
assign n_2431 = n_2405 ^ n_2281;
assign n_2432 = n_2406 ^ n_2282;
assign n_2433 = n_2407 ^ n_2283;
assign n_2434 = n_2408 ^ n_2284;
assign n_2435 = n_2409 ^ n_2285;
assign n_2436 = n_2411 ^ n_2245;
assign n_2437 = n_68 ^ n_2412;
assign n_2438 = n_271 & ~n_2413;
assign n_2439 = n_2418 ^ x88;
assign n_2440 = n_2419 ^ x87;
assign n_2441 = n_2385 ^ n_2436;
assign n_2442 = ~n_2437 & ~n_2438;
assign n_2443 = n_2441 ^ x40;
assign n_2444 = x66 ^ n_2442;
assign n_2445 = n_2443 ^ x66;
assign n_2446 = n_2443 ^ n_2442;
assign n_2447 = ~n_2445 & ~n_2446;
assign n_2448 = n_2447 ^ x66;
assign n_2449 = n_2448 ^ x67;
assign n_2450 = n_2414 ^ n_2448;
assign n_2451 = n_2449 & n_2450;
assign n_2452 = n_2451 ^ x67;
assign n_2453 = n_2452 ^ x68;
assign n_2454 = n_2415 ^ n_2452;
assign n_2455 = n_2453 & n_2454;
assign n_2456 = n_2455 ^ x68;
assign n_2457 = n_2456 ^ x69;
assign n_2458 = n_2416 ^ n_2456;
assign n_2459 = n_2457 & n_2458;
assign n_2460 = n_2459 ^ x69;
assign n_2461 = n_2460 ^ x70;
assign n_2462 = n_2417 ^ n_2460;
assign n_2463 = n_2461 & n_2462;
assign n_2464 = n_2463 ^ x70;
assign n_2465 = n_2464 ^ x71;
assign n_2466 = n_2420 ^ n_2464;
assign n_2467 = n_2465 & n_2466;
assign n_2468 = n_2467 ^ x71;
assign n_2469 = n_2468 ^ x72;
assign n_2470 = n_2421 ^ n_2468;
assign n_2471 = n_2469 & n_2470;
assign n_2472 = n_2471 ^ x72;
assign n_2473 = n_2472 ^ x73;
assign n_2474 = n_2422 ^ n_2472;
assign n_2475 = n_2473 & n_2474;
assign n_2476 = n_2475 ^ x73;
assign n_2477 = n_2476 ^ x74;
assign n_2478 = n_2423 ^ n_2476;
assign n_2479 = n_2477 & n_2478;
assign n_2480 = n_2479 ^ x74;
assign n_2481 = n_2480 ^ x75;
assign n_2482 = n_2424 ^ n_2480;
assign n_2483 = n_2481 & n_2482;
assign n_2484 = n_2483 ^ x75;
assign n_2485 = n_2484 ^ x76;
assign n_2486 = n_2425 ^ n_2484;
assign n_2487 = n_2485 & n_2486;
assign n_2488 = n_2487 ^ x76;
assign n_2489 = n_2488 ^ x77;
assign n_2490 = n_2426 ^ n_2488;
assign n_2491 = n_2489 & n_2490;
assign n_2492 = n_2491 ^ x77;
assign n_2493 = n_2492 ^ x78;
assign n_2494 = n_2427 ^ n_2492;
assign n_2495 = n_2493 & n_2494;
assign n_2496 = n_2495 ^ x78;
assign n_2497 = n_2496 ^ x79;
assign n_2498 = n_2428 ^ n_2496;
assign n_2499 = n_2497 & n_2498;
assign n_2500 = n_2499 ^ x79;
assign n_2501 = n_2500 ^ x80;
assign n_2502 = n_2429 ^ n_2500;
assign n_2503 = n_2501 & n_2502;
assign n_2504 = n_2503 ^ x80;
assign n_2505 = n_2504 ^ x81;
assign n_2506 = n_2430 ^ n_2504;
assign n_2507 = n_2505 & n_2506;
assign n_2508 = n_2507 ^ x81;
assign n_2509 = n_2508 ^ x82;
assign n_2510 = n_2431 ^ n_2508;
assign n_2511 = n_2509 & n_2510;
assign n_2512 = n_2511 ^ x82;
assign n_2513 = n_2512 ^ x83;
assign n_2514 = n_2432 ^ n_2512;
assign n_2515 = n_2513 & n_2514;
assign n_2516 = n_2515 ^ x83;
assign n_2517 = n_2516 ^ x84;
assign n_2518 = n_2433 ^ n_2516;
assign n_2519 = n_2517 & n_2518;
assign n_2520 = n_2519 ^ x84;
assign n_2521 = n_2520 ^ x85;
assign n_2522 = n_2434 ^ n_2520;
assign n_2523 = n_2521 & n_2522;
assign n_2524 = n_2523 ^ x85;
assign n_2525 = n_2524 ^ x86;
assign n_2526 = n_2435 ^ n_2524;
assign n_2527 = n_2525 & n_2526;
assign n_2528 = n_2527 ^ x86;
assign n_2529 = n_2528 ^ n_2419;
assign n_2530 = n_2528 ^ x87;
assign n_2531 = ~n_2440 & n_2529;
assign n_2532 = n_2531 ^ x87;
assign n_2533 = n_2532 ^ n_2418;
assign n_2534 = n_2532 ^ x88;
assign n_2535 = ~n_2439 & n_2533;
assign n_2536 = n_2535 ^ x88;
assign n_2537 = n_2536 ^ x89;
assign n_2538 = n_2536 ^ ~n_2410;
assign n_2539 = n_2537 & ~n_2538;
assign n_2540 = n_2539 ^ x89;
assign n_2541 = n_380 & ~n_2540;
assign n_2542 = ~x90 ^ ~n_2540;
assign n_2543 = n_2465 & n_2541;
assign n_2544 = n_2461 & n_2541;
assign n_2545 = x65 & n_2541;
assign n_2546 = x64 & n_2541;
assign n_2547 = n_2541 & ~n_2444;
assign n_2548 = n_2449 & n_2541;
assign n_2549 = n_2453 & n_2541;
assign n_2550 = n_2457 & n_2541;
assign n_2551 = n_2469 & n_2541;
assign n_2552 = n_2473 & n_2541;
assign n_2553 = n_2477 & n_2541;
assign n_2554 = n_2481 & n_2541;
assign n_2555 = n_2485 & n_2541;
assign n_2556 = n_2489 & n_2541;
assign n_2557 = n_2493 & n_2541;
assign n_2558 = n_2497 & n_2541;
assign n_2559 = n_2501 & n_2541;
assign n_2560 = n_2505 & n_2541;
assign n_2561 = n_2509 & n_2541;
assign n_2562 = n_2513 & n_2541;
assign n_2563 = n_2517 & n_2541;
assign n_2564 = n_2521 & n_2541;
assign n_2565 = n_2525 & n_2541;
assign n_2566 = n_2541 & n_2530;
assign n_2567 = n_2541 & n_2534;
assign y38 = n_2541;
assign n_2568 = ~n_2541 & n_145;
assign n_2569 = n_2410 & n_2542;
assign n_2570 = n_2543 ^ n_2420;
assign n_2571 = n_2544 ^ n_2417;
assign n_2572 = x38 & n_2546;
assign n_2573 = n_2546 ^ n_2386;
assign n_2574 = n_2546 & ~n_71;
assign n_2575 = n_2546 ^ x38;
assign n_2576 = n_2547 ^ n_2443;
assign n_2577 = n_2548 ^ n_2414;
assign n_2578 = n_2549 ^ n_2415;
assign n_2579 = n_2550 ^ n_2416;
assign n_2580 = n_2551 ^ n_2421;
assign n_2581 = n_2552 ^ n_2422;
assign n_2582 = n_2553 ^ n_2423;
assign n_2583 = n_2554 ^ n_2424;
assign n_2584 = n_2555 ^ n_2425;
assign n_2585 = n_2556 ^ n_2426;
assign n_2586 = n_2557 ^ n_2427;
assign n_2587 = n_2558 ^ n_2428;
assign n_2588 = n_2559 ^ n_2429;
assign n_2589 = n_2560 ^ n_2430;
assign n_2590 = n_2561 ^ n_2431;
assign n_2591 = n_2562 ^ n_2432;
assign n_2592 = n_2563 ^ n_2433;
assign n_2593 = n_2564 ^ n_2434;
assign n_2594 = n_2565 ^ n_2435;
assign n_2595 = n_2566 ^ n_2419;
assign n_2596 = n_2567 ^ n_2418;
assign n_2597 = ~n_439 ^ ~n_2569;
assign n_2598 = ~x72 ^ n_2570;
assign n_2599 = n_2570 ^ x72;
assign n_2600 = n_2571 ^ x71;
assign n_2601 = x71 & ~n_2571;
assign n_2602 = n_2572 ^ n_2573;
assign n_2603 = n_2574 ^ n_146;
assign n_2604 = n_2600 ^ n_2601;
assign n_2605 = n_2601 ^ n_2570;
assign n_2606 = n_2545 ^ n_2602;
assign n_2607 = n_2603 ^ n_70;
assign n_2608 = n_2598 & ~n_2604;
assign n_2609 = ~n_2599 & n_2605;
assign n_2610 = n_2606 ^ x39;
assign n_2611 = n_2607 ^ n_2568;
assign n_2612 = n_2609 ^ x72;
assign n_2613 = n_2610 ^ x66;
assign n_2614 = n_2611 ^ n_2610;
assign n_2615 = n_2611 ^ x66;
assign n_2616 = ~n_2613 & n_2614;
assign n_2617 = n_2616 ^ x66;
assign n_2618 = n_2617 ^ x67;
assign n_2619 = n_2576 ^ n_2617;
assign n_2620 = n_2618 & n_2619;
assign n_2621 = n_2620 ^ x67;
assign n_2622 = n_2621 ^ x68;
assign n_2623 = n_2577 ^ n_2621;
assign n_2624 = n_2622 & n_2623;
assign n_2625 = n_2624 ^ x68;
assign n_2626 = n_2625 ^ x69;
assign n_2627 = n_2578 ^ n_2625;
assign n_2628 = n_2626 & n_2627;
assign n_2629 = n_2628 ^ x69;
assign n_2630 = n_2629 ^ x70;
assign n_2631 = n_2579 ^ n_2629;
assign n_2632 = n_2630 & n_2631;
assign n_2633 = n_2632 ^ x70;
assign n_2634 = n_2633 ^ x71;
assign n_2635 = n_2633 ^ n_2571;
assign n_2636 = n_2608 & n_2633;
assign n_2637 = n_2634 & n_2635;
assign n_2638 = ~n_2612 & ~n_2636;
assign n_2639 = n_2637 ^ x71;
assign n_2640 = x73 ^ n_2638;
assign n_2641 = n_2580 ^ n_2638;
assign n_2642 = n_2639 ^ x72;
assign n_2643 = ~n_2640 & ~n_2641;
assign n_2644 = n_2643 ^ x73;
assign n_2645 = n_2644 ^ x74;
assign n_2646 = n_2581 ^ n_2644;
assign n_2647 = n_2645 & n_2646;
assign n_2648 = n_2647 ^ x74;
assign n_2649 = n_2648 ^ x75;
assign n_2650 = n_2582 ^ n_2648;
assign n_2651 = n_2649 & n_2650;
assign n_2652 = n_2651 ^ x75;
assign n_2653 = n_2652 ^ x76;
assign n_2654 = n_2583 ^ n_2652;
assign n_2655 = n_2653 & n_2654;
assign n_2656 = n_2655 ^ x76;
assign n_2657 = n_2656 ^ x77;
assign n_2658 = n_2584 ^ n_2656;
assign n_2659 = n_2657 & n_2658;
assign n_2660 = n_2659 ^ x77;
assign n_2661 = n_2660 ^ x78;
assign n_2662 = n_2585 ^ n_2660;
assign n_2663 = n_2661 & n_2662;
assign n_2664 = n_2663 ^ x78;
assign n_2665 = n_2664 ^ x79;
assign n_2666 = n_2586 ^ n_2664;
assign n_2667 = n_2665 & n_2666;
assign n_2668 = n_2667 ^ x79;
assign n_2669 = n_2668 ^ x80;
assign n_2670 = n_2587 ^ n_2668;
assign n_2671 = n_2669 & n_2670;
assign n_2672 = n_2671 ^ x80;
assign n_2673 = n_2672 ^ x81;
assign n_2674 = n_2588 ^ n_2672;
assign n_2675 = n_2673 & n_2674;
assign n_2676 = n_2675 ^ x81;
assign n_2677 = n_2676 ^ x82;
assign n_2678 = n_2589 ^ n_2676;
assign n_2679 = n_2677 & n_2678;
assign n_2680 = n_2679 ^ x82;
assign n_2681 = n_2680 ^ x83;
assign n_2682 = n_2590 ^ n_2680;
assign n_2683 = n_2681 & n_2682;
assign n_2684 = n_2683 ^ x83;
assign n_2685 = n_2684 ^ x84;
assign n_2686 = n_2591 ^ n_2684;
assign n_2687 = n_2685 & n_2686;
assign n_2688 = n_2687 ^ x84;
assign n_2689 = n_2688 ^ x85;
assign n_2690 = n_2592 ^ n_2688;
assign n_2691 = n_2689 & n_2690;
assign n_2692 = n_2691 ^ x85;
assign n_2693 = n_2692 ^ x86;
assign n_2694 = n_2593 ^ n_2692;
assign n_2695 = n_2693 & n_2694;
assign n_2696 = n_2695 ^ x86;
assign n_2697 = n_2696 ^ x87;
assign n_2698 = n_2594 ^ n_2696;
assign n_2699 = n_2697 & n_2698;
assign n_2700 = n_2699 ^ x87;
assign n_2701 = n_2700 ^ x88;
assign n_2702 = n_2595 ^ n_2700;
assign n_2703 = n_2701 & n_2702;
assign n_2704 = n_2703 ^ x88;
assign n_2705 = n_2704 ^ x89;
assign n_2706 = n_2596 ^ n_2704;
assign n_2707 = n_2705 & n_2706;
assign n_2708 = n_2707 ^ x89;
assign n_2709 = x90 & n_2708;
assign n_2710 = n_2708 ^ x90;
assign n_2711 = ~n_2597 ^ n_2708;
assign n_2712 = ~n_2709 & ~n_442;
assign n_2713 = n_2710 & ~n_2711;
assign n_2714 = n_2410 & ~n_2712;
assign n_2715 = x90 ^ n_2713;
assign n_2716 = n_379 & ~n_2715;
assign n_2717 = n_2705 & n_2716;
assign n_2718 = n_2701 & n_2716;
assign n_2719 = n_2669 & n_2716;
assign n_2720 = n_2665 & n_2716;
assign n_2721 = n_147 & n_2716;
assign n_2722 = x64 & n_2716;
assign n_2723 = ~n_336 & ~n_2716;
assign n_2724 = n_2615 & n_2716;
assign n_2725 = n_2618 & n_2716;
assign n_2726 = n_2622 & n_2716;
assign n_2727 = n_2626 & n_2716;
assign n_2728 = n_2630 & n_2716;
assign n_2729 = n_2634 & n_2716;
assign n_2730 = ~n_2640 & n_2716;
assign n_2731 = n_2645 & n_2716;
assign n_2732 = n_2649 & n_2716;
assign n_2733 = n_2653 & n_2716;
assign n_2734 = n_2657 & n_2716;
assign n_2735 = n_2661 & n_2716;
assign n_2736 = n_2673 & n_2716;
assign n_2737 = n_2677 & n_2716;
assign n_2738 = n_2681 & n_2716;
assign n_2739 = n_2685 & n_2716;
assign n_2740 = n_2689 & n_2716;
assign n_2741 = n_2693 & n_2716;
assign n_2742 = n_2697 & n_2716;
assign y37 = n_2716;
assign n_2743 = n_2642 & n_2716;
assign n_2744 = n_2717 ^ n_2596;
assign n_2745 = n_2718 ^ n_2595;
assign n_2746 = n_2719 ^ n_2587;
assign n_2747 = n_2720 ^ n_2586;
assign n_2748 = n_2575 ^ n_2721;
assign n_2749 = n_2722 ^ x37;
assign n_2750 = n_2722 & n_273;
assign n_2751 = n_2723 ^ x65;
assign n_2752 = n_2724 ^ n_2610;
assign n_2753 = n_2725 ^ n_2576;
assign n_2754 = n_2726 ^ n_2577;
assign n_2755 = n_2727 ^ n_2578;
assign n_2756 = n_2728 ^ n_2579;
assign n_2757 = n_2729 ^ n_2571;
assign n_2758 = n_2730 ^ n_2580;
assign n_2759 = n_2731 ^ n_2581;
assign n_2760 = n_2732 ^ n_2582;
assign n_2761 = n_2733 ^ n_2583;
assign n_2762 = n_2734 ^ n_2584;
assign n_2763 = n_2735 ^ n_2585;
assign n_2764 = n_2736 ^ n_2588;
assign n_2765 = n_2737 ^ n_2589;
assign n_2766 = n_2738 ^ n_2590;
assign n_2767 = n_2739 ^ n_2591;
assign n_2768 = n_2740 ^ n_2592;
assign n_2769 = n_2741 ^ n_2593;
assign n_2770 = n_2742 ^ n_2594;
assign n_2771 = n_2570 ^ n_2743;
assign n_2772 = n_2744 ^ x90;
assign n_2773 = n_2745 ^ x89;
assign n_2774 = n_2746 ^ x81;
assign n_2775 = n_2747 ^ x80;
assign n_2776 = n_2748 ^ x66;
assign n_2777 = ~n_344 & n_2751;
assign n_2778 = x65 ^ n_2777;
assign n_2779 = n_2778 ^ x65;
assign n_2780 = n_2779 ^ x65;
assign n_2781 = ~n_2780 & ~n_2750;
assign n_2782 = n_2748 ^ n_2781;
assign n_2783 = x66 ^ n_2781;
assign n_2784 = ~n_2776 & ~n_2782;
assign n_2785 = n_2784 ^ x66;
assign n_2786 = n_2785 ^ x67;
assign n_2787 = n_2752 ^ n_2785;
assign n_2788 = n_2786 & n_2787;
assign n_2789 = n_2788 ^ x67;
assign n_2790 = n_2789 ^ x68;
assign n_2791 = n_2753 ^ n_2789;
assign n_2792 = n_2790 & n_2791;
assign n_2793 = n_2792 ^ x68;
assign n_2794 = n_2793 ^ x69;
assign n_2795 = n_2754 ^ n_2793;
assign n_2796 = n_2794 & n_2795;
assign n_2797 = n_2796 ^ x69;
assign n_2798 = n_2797 ^ x70;
assign n_2799 = n_2755 ^ n_2797;
assign n_2800 = n_2798 & n_2799;
assign n_2801 = n_2800 ^ x70;
assign n_2802 = n_2801 ^ x71;
assign n_2803 = n_2756 ^ n_2801;
assign n_2804 = n_2802 & n_2803;
assign n_2805 = n_2804 ^ x71;
assign n_2806 = n_2805 ^ x72;
assign n_2807 = n_2757 ^ n_2805;
assign n_2808 = n_2806 & n_2807;
assign n_2809 = n_2808 ^ x72;
assign n_2810 = n_2809 ^ x73;
assign n_2811 = n_2771 ^ n_2809;
assign n_2812 = n_2810 & n_2811;
assign n_2813 = n_2812 ^ x73;
assign n_2814 = n_2813 ^ x74;
assign n_2815 = n_2758 ^ n_2813;
assign n_2816 = n_2814 & n_2815;
assign n_2817 = n_2816 ^ x74;
assign n_2818 = n_2817 ^ x75;
assign n_2819 = n_2759 ^ n_2817;
assign n_2820 = n_2818 & n_2819;
assign n_2821 = n_2820 ^ x75;
assign n_2822 = n_2821 ^ x76;
assign n_2823 = n_2760 ^ n_2821;
assign n_2824 = n_2822 & n_2823;
assign n_2825 = n_2824 ^ x76;
assign n_2826 = n_2825 ^ x77;
assign n_2827 = n_2761 ^ n_2825;
assign n_2828 = n_2826 & n_2827;
assign n_2829 = n_2828 ^ x77;
assign n_2830 = n_2829 ^ x78;
assign n_2831 = n_2762 ^ n_2829;
assign n_2832 = n_2830 & n_2831;
assign n_2833 = n_2832 ^ x78;
assign n_2834 = n_2833 ^ x79;
assign n_2835 = n_2763 ^ n_2833;
assign n_2836 = n_2834 & n_2835;
assign n_2837 = n_2836 ^ x79;
assign n_2838 = n_2837 ^ n_2747;
assign n_2839 = n_2837 ^ x80;
assign n_2840 = ~n_2775 & n_2838;
assign n_2841 = n_2840 ^ x80;
assign n_2842 = n_2841 ^ n_2746;
assign n_2843 = n_2841 ^ x81;
assign n_2844 = ~n_2774 & n_2842;
assign n_2845 = n_2844 ^ x81;
assign n_2846 = n_2845 ^ x82;
assign n_2847 = n_2764 ^ n_2845;
assign n_2848 = n_2846 & n_2847;
assign n_2849 = n_2848 ^ x82;
assign n_2850 = n_2849 ^ x83;
assign n_2851 = n_2765 ^ n_2849;
assign n_2852 = n_2850 & n_2851;
assign n_2853 = n_2852 ^ x83;
assign n_2854 = n_2853 ^ x84;
assign n_2855 = n_2766 ^ n_2853;
assign n_2856 = n_2854 & n_2855;
assign n_2857 = n_2856 ^ x84;
assign n_2858 = n_2857 ^ x85;
assign n_2859 = n_2767 ^ n_2857;
assign n_2860 = n_2858 & n_2859;
assign n_2861 = n_2860 ^ x85;
assign n_2862 = n_2861 ^ x86;
assign n_2863 = n_2768 ^ n_2861;
assign n_2864 = n_2862 & n_2863;
assign n_2865 = n_2864 ^ x86;
assign n_2866 = n_2865 ^ x87;
assign n_2867 = n_2769 ^ n_2865;
assign n_2868 = n_2866 & n_2867;
assign n_2869 = n_2868 ^ x87;
assign n_2870 = n_2869 ^ x88;
assign n_2871 = n_2770 ^ n_2869;
assign n_2872 = n_2870 & n_2871;
assign n_2873 = n_2872 ^ x88;
assign n_2874 = n_2873 ^ n_2745;
assign n_2875 = n_2873 ^ x89;
assign n_2876 = ~n_2773 & n_2874;
assign n_2877 = n_2876 ^ x89;
assign n_2878 = n_2877 ^ n_2744;
assign n_2879 = n_2877 ^ x90;
assign n_2880 = ~n_2772 & n_2878;
assign n_2881 = n_2880 ^ x90;
assign n_2882 = n_2881 ^ x91;
assign n_2883 = n_2881 ^ n_2714;
assign n_2884 = n_2882 & n_2883;
assign n_2885 = n_2884 ^ x91;
assign n_2886 = n_378 & ~n_2885;
assign n_2887 = n_2714 & ~n_2886;
assign n_2888 = n_2879 & n_2886;
assign n_2889 = n_2875 & n_2886;
assign n_2890 = n_2870 & n_2886;
assign n_2891 = n_2866 & n_2886;
assign n_2892 = n_2862 & n_2886;
assign n_2893 = n_2790 & n_2886;
assign n_2894 = n_2786 & n_2886;
assign n_2895 = x64 & n_2886;
assign n_2896 = n_148 & n_2886;
assign n_2897 = ~n_2783 & n_2886;
assign n_2898 = n_2794 & n_2886;
assign n_2899 = n_2798 & n_2886;
assign n_2900 = n_2802 & n_2886;
assign n_2901 = n_2806 & n_2886;
assign n_2902 = n_2810 & n_2886;
assign n_2903 = n_2814 & n_2886;
assign n_2904 = n_2818 & n_2886;
assign n_2905 = n_2822 & n_2886;
assign n_2906 = n_2826 & n_2886;
assign n_2907 = n_2830 & n_2886;
assign n_2908 = n_2834 & n_2886;
assign n_2909 = n_2839 & n_2886;
assign n_2910 = n_2843 & n_2886;
assign n_2911 = n_2846 & n_2886;
assign n_2912 = n_2850 & n_2886;
assign n_2913 = n_2854 & n_2886;
assign n_2914 = n_2858 & n_2886;
assign y36 = n_2886;
assign n_2915 = ~n_439 ^ ~n_2887;
assign n_2916 = n_2888 ^ n_2744;
assign n_2917 = n_2889 ^ n_2745;
assign n_2918 = n_2890 ^ n_2770;
assign n_2919 = n_2891 ^ n_2769;
assign n_2920 = n_2892 ^ n_2768;
assign n_2921 = n_2893 ^ n_2753;
assign n_2922 = n_2894 ^ n_2752;
assign n_2923 = n_16 ^ n_2895;
assign n_2924 = n_2895 ^ x36;
assign n_2925 = n_2749 ^ n_2896;
assign n_2926 = n_2897 ^ n_2748;
assign n_2927 = n_2898 ^ n_2754;
assign n_2928 = n_2899 ^ n_2755;
assign n_2929 = n_2900 ^ n_2756;
assign n_2930 = n_2901 ^ n_2757;
assign n_2931 = n_2902 ^ n_2771;
assign n_2932 = n_2903 ^ n_2758;
assign n_2933 = n_2904 ^ n_2759;
assign n_2934 = n_2905 ^ n_2760;
assign n_2935 = n_2906 ^ n_2761;
assign n_2936 = n_2907 ^ n_2762;
assign n_2937 = n_2908 ^ n_2763;
assign n_2938 = n_2909 ^ n_2747;
assign n_2939 = n_2910 ^ n_2746;
assign n_2940 = n_2911 ^ n_2764;
assign n_2941 = n_2912 ^ n_2765;
assign n_2942 = n_2913 ^ n_2766;
assign n_2943 = n_2914 ^ n_2767;
assign n_2944 = ~x92 ^ n_2915;
assign n_2945 = ~n_2915 ^ x92;
assign n_2946 = n_2916 ^ x91;
assign n_2947 = x91 & ~n_2916;
assign n_2948 = n_2917 ^ x90;
assign n_2949 = n_2918 ^ x89;
assign n_2950 = ~x88 ^ n_2919;
assign n_2951 = n_2919 ^ x88;
assign n_2952 = n_2920 ^ x87;
assign n_2953 = x87 & ~n_2920;
assign n_2954 = ~x69 ^ n_2921;
assign n_2955 = n_2921 ^ x69;
assign n_2956 = n_2922 ^ x68;
assign n_2957 = x68 & ~n_2922;
assign n_2958 = ~x35 & n_2923;
assign n_2959 = x65 & ~n_2924;
assign n_2960 = n_2946 ^ n_2947;
assign n_2961 = n_2947 ^ x92;
assign n_2962 = n_2952 ^ n_2953;
assign n_2963 = n_2953 ^ n_2919;
assign n_2964 = n_2956 ^ n_2957;
assign n_2965 = n_2957 ^ n_2921;
assign n_2966 = n_2958 ^ n_204;
assign n_2967 = n_2944 ^ ~n_2960;
assign n_2968 = n_2945 & n_2961;
assign n_2969 = n_2950 & ~n_2962;
assign n_2970 = ~n_2951 & n_2963;
assign n_2971 = n_2954 & ~n_2964;
assign n_2972 = ~n_2955 & n_2965;
assign n_2973 = n_2966 ^ n_2959;
assign n_2974 = n_2968 ^ x92;
assign n_2975 = n_2970 ^ x88;
assign n_2976 = n_2972 ^ x69;
assign n_2977 = n_2973 ^ x66;
assign n_2978 = n_2925 ^ n_2973;
assign n_2979 = n_377 & ~n_2974;
assign n_2980 = n_2977 & n_2978;
assign n_2981 = n_2980 ^ x66;
assign n_2982 = n_2981 ^ x67;
assign n_2983 = n_2926 ^ n_2981;
assign n_2984 = n_2982 & n_2983;
assign n_2985 = n_2984 ^ x67;
assign n_2986 = n_2985 ^ x68;
assign n_2987 = n_2985 ^ n_2922;
assign n_2988 = n_2971 & n_2985;
assign n_2989 = n_2986 & n_2987;
assign n_2990 = ~n_2976 & ~n_2988;
assign n_2991 = n_2989 ^ x68;
assign n_2992 = x70 ^ n_2990;
assign n_2993 = n_2927 ^ n_2990;
assign n_2994 = n_2991 ^ x69;
assign n_2995 = ~n_2992 & ~n_2993;
assign n_2996 = n_2995 ^ x70;
assign n_2997 = n_2996 ^ x71;
assign n_2998 = n_2928 ^ n_2996;
assign n_2999 = n_2997 & n_2998;
assign n_3000 = n_2999 ^ x71;
assign n_3001 = n_3000 ^ x72;
assign n_3002 = n_2929 ^ n_3000;
assign n_3003 = n_3001 & n_3002;
assign n_3004 = n_3003 ^ x72;
assign n_3005 = n_3004 ^ x73;
assign n_3006 = n_2930 ^ n_3004;
assign n_3007 = n_3005 & n_3006;
assign n_3008 = n_3007 ^ x73;
assign n_3009 = n_3008 ^ x74;
assign n_3010 = n_2931 ^ n_3008;
assign n_3011 = n_3009 & n_3010;
assign n_3012 = n_3011 ^ x74;
assign n_3013 = n_3012 ^ x75;
assign n_3014 = n_2932 ^ n_3012;
assign n_3015 = n_3013 & n_3014;
assign n_3016 = n_3015 ^ x75;
assign n_3017 = n_3016 ^ x76;
assign n_3018 = n_2933 ^ n_3016;
assign n_3019 = n_3017 & n_3018;
assign n_3020 = n_3019 ^ x76;
assign n_3021 = n_3020 ^ x77;
assign n_3022 = n_2934 ^ n_3020;
assign n_3023 = n_3021 & n_3022;
assign n_3024 = n_3023 ^ x77;
assign n_3025 = n_3024 ^ x78;
assign n_3026 = n_2935 ^ n_3024;
assign n_3027 = n_3025 & n_3026;
assign n_3028 = n_3027 ^ x78;
assign n_3029 = n_3028 ^ x79;
assign n_3030 = n_2936 ^ n_3028;
assign n_3031 = n_3029 & n_3030;
assign n_3032 = n_3031 ^ x79;
assign n_3033 = n_3032 ^ x80;
assign n_3034 = n_2937 ^ n_3032;
assign n_3035 = n_3033 & n_3034;
assign n_3036 = n_3035 ^ x80;
assign n_3037 = n_3036 ^ x81;
assign n_3038 = n_2938 ^ n_3036;
assign n_3039 = n_3037 & n_3038;
assign n_3040 = n_3039 ^ x81;
assign n_3041 = n_3040 ^ x82;
assign n_3042 = n_2939 ^ n_3040;
assign n_3043 = n_3041 & n_3042;
assign n_3044 = n_3043 ^ x82;
assign n_3045 = n_3044 ^ x83;
assign n_3046 = n_2940 ^ n_3044;
assign n_3047 = n_3045 & n_3046;
assign n_3048 = n_3047 ^ x83;
assign n_3049 = n_3048 ^ x84;
assign n_3050 = n_2941 ^ n_3048;
assign n_3051 = n_3049 & n_3050;
assign n_3052 = n_3051 ^ x84;
assign n_3053 = n_3052 ^ x85;
assign n_3054 = n_2942 ^ n_3052;
assign n_3055 = n_3053 & n_3054;
assign n_3056 = n_3055 ^ x85;
assign n_3057 = n_3056 ^ x86;
assign n_3058 = n_2943 ^ n_3056;
assign n_3059 = n_3057 & n_3058;
assign n_3060 = n_3059 ^ x86;
assign n_3061 = n_3060 ^ x87;
assign n_3062 = n_3060 ^ n_2920;
assign n_3063 = n_2969 & n_3060;
assign n_3064 = n_3061 & n_3062;
assign n_3065 = ~n_2975 & ~n_3063;
assign n_3066 = n_3064 ^ x87;
assign n_3067 = n_2918 ^ n_3065;
assign n_3068 = x89 ^ n_3065;
assign n_3069 = n_3066 ^ x88;
assign n_3070 = ~n_2949 & ~n_3067;
assign n_3071 = n_3070 ^ x89;
assign n_3072 = n_3071 ^ n_2917;
assign n_3073 = n_3071 ^ x90;
assign n_3074 = ~n_2948 & n_3072;
assign n_3075 = n_3074 ^ x90;
assign n_3076 = ~n_2967 & n_3075;
assign n_3077 = n_3075 ^ x91;
assign n_3078 = ~n_3076 & n_2979;
assign n_3079 = n_3073 & n_3078;
assign n_3080 = ~n_3068 & n_3078;
assign n_3081 = n_3017 & n_3078;
assign n_3082 = n_3013 & n_3078;
assign n_3083 = x35 ^ n_3078;
assign n_3084 = x64 & n_3078;
assign n_3085 = x65 & n_3078;
assign n_3086 = n_2977 & n_3078;
assign n_3087 = n_2982 & n_3078;
assign n_3088 = n_2986 & n_3078;
assign n_3089 = ~n_2992 & n_3078;
assign n_3090 = n_2997 & n_3078;
assign n_3091 = n_3001 & n_3078;
assign n_3092 = n_3005 & n_3078;
assign n_3093 = n_3009 & n_3078;
assign n_3094 = n_3021 & n_3078;
assign n_3095 = n_3025 & n_3078;
assign n_3096 = n_3029 & n_3078;
assign n_3097 = n_3033 & n_3078;
assign n_3098 = n_3037 & n_3078;
assign n_3099 = n_3041 & n_3078;
assign n_3100 = n_3045 & n_3078;
assign n_3101 = n_3049 & n_3078;
assign n_3102 = n_3053 & n_3078;
assign n_3103 = n_3057 & n_3078;
assign n_3104 = n_3061 & n_3078;
assign n_3105 = n_3077 & n_3078;
assign n_3106 = n_2915 & ~n_3078;
assign y35 = n_3078;
assign n_3107 = n_2994 & n_3078;
assign n_3108 = n_3069 & n_3078;
assign n_3109 = n_3079 ^ n_2917;
assign n_3110 = n_3080 ^ n_2918;
assign n_3111 = n_3081 ^ n_2933;
assign n_3112 = n_3082 ^ n_2932;
assign n_3113 = ~x34 & n_3083;
assign n_3114 = x65 & n_3084;
assign n_3115 = n_3084 & n_3083;
assign n_3116 = n_3084 ^ x35;
assign n_3117 = n_3086 ^ n_2925;
assign n_3118 = n_3087 ^ n_2926;
assign n_3119 = n_3088 ^ n_2922;
assign n_3120 = n_3089 ^ n_2927;
assign n_3121 = n_3090 ^ n_2928;
assign n_3122 = n_3091 ^ n_2929;
assign n_3123 = n_3092 ^ n_2930;
assign n_3124 = n_3093 ^ n_2931;
assign n_3125 = n_3094 ^ n_2934;
assign n_3126 = n_3095 ^ n_2935;
assign n_3127 = n_3096 ^ n_2936;
assign n_3128 = n_3097 ^ n_2937;
assign n_3129 = n_3098 ^ n_2938;
assign n_3130 = n_3099 ^ n_2939;
assign n_3131 = n_3100 ^ n_2940;
assign n_3132 = n_3101 ^ n_2941;
assign n_3133 = n_3102 ^ n_2942;
assign n_3134 = n_3103 ^ n_2943;
assign n_3135 = n_3104 ^ n_2920;
assign n_3136 = n_3105 ^ n_2916;
assign n_3137 = ~n_439 & ~n_3106;
assign n_3138 = n_2921 ^ n_3107;
assign n_3139 = n_2919 ^ n_3108;
assign n_3140 = ~x91 ^ n_3109;
assign n_3141 = n_3109 ^ x91;
assign n_3142 = n_3110 ^ x90;
assign n_3143 = x90 & ~n_3110;
assign n_3144 = ~x77 ^ n_3111;
assign n_3145 = n_3111 ^ x77;
assign n_3146 = n_3112 ^ x76;
assign n_3147 = x76 & ~n_3112;
assign n_3148 = n_3113 ^ n_205;
assign n_3149 = n_3115 ^ n_3085;
assign n_3150 = ~n_377 & ~n_3137;
assign n_3151 = x93 ^ n_3137;
assign n_3152 = n_375 & ~n_3137;
assign n_3153 = n_3142 ^ n_3143;
assign n_3154 = n_3143 ^ n_3109;
assign n_3155 = n_3146 ^ n_3147;
assign n_3156 = n_3147 ^ n_3111;
assign n_3157 = x64 & ~n_3148;
assign n_3158 = n_3149 ^ n_2895;
assign n_3159 = ~n_376 & ~n_3152;
assign n_3160 = n_3140 & ~n_3153;
assign n_3161 = ~n_3141 & n_3154;
assign n_3162 = n_3144 & ~n_3155;
assign n_3163 = ~n_3145 & n_3156;
assign n_3164 = n_3114 ^ n_3157;
assign n_3165 = n_3158 ^ x36;
assign n_3166 = n_3161 ^ x91;
assign n_3167 = n_3163 ^ x77;
assign n_3168 = n_3164 ^ n_74;
assign n_3169 = n_3168 ^ x66;
assign n_3170 = n_3165 ^ n_3168;
assign n_3171 = n_3169 & n_3170;
assign n_3172 = n_3171 ^ x66;
assign n_3173 = n_3172 ^ x67;
assign n_3174 = n_3117 ^ n_3172;
assign n_3175 = n_3173 & n_3174;
assign n_3176 = n_3175 ^ x67;
assign n_3177 = n_3176 ^ x68;
assign n_3178 = n_3118 ^ n_3176;
assign n_3179 = n_3177 & n_3178;
assign n_3180 = n_3179 ^ x68;
assign n_3181 = n_3180 ^ x69;
assign n_3182 = n_3119 ^ n_3180;
assign n_3183 = n_3181 & n_3182;
assign n_3184 = n_3183 ^ x69;
assign n_3185 = n_3184 ^ x70;
assign n_3186 = n_3138 ^ n_3184;
assign n_3187 = n_3185 & n_3186;
assign n_3188 = n_3187 ^ x70;
assign n_3189 = n_3188 ^ x71;
assign n_3190 = n_3120 ^ n_3188;
assign n_3191 = n_3189 & n_3190;
assign n_3192 = n_3191 ^ x71;
assign n_3193 = n_3192 ^ x72;
assign n_3194 = n_3121 ^ n_3192;
assign n_3195 = n_3193 & n_3194;
assign n_3196 = n_3195 ^ x72;
assign n_3197 = n_3196 ^ x73;
assign n_3198 = n_3122 ^ n_3196;
assign n_3199 = n_3197 & n_3198;
assign n_3200 = n_3199 ^ x73;
assign n_3201 = n_3200 ^ x74;
assign n_3202 = n_3123 ^ n_3200;
assign n_3203 = n_3201 & n_3202;
assign n_3204 = n_3203 ^ x74;
assign n_3205 = n_3204 ^ x75;
assign n_3206 = n_3124 ^ n_3204;
assign n_3207 = n_3205 & n_3206;
assign n_3208 = n_3207 ^ x75;
assign n_3209 = n_3208 ^ x76;
assign n_3210 = n_3208 ^ n_3112;
assign n_3211 = n_3162 & n_3208;
assign n_3212 = n_3209 & n_3210;
assign n_3213 = ~n_3167 & ~n_3211;
assign n_3214 = n_3212 ^ x76;
assign n_3215 = x78 ^ n_3213;
assign n_3216 = n_3125 ^ n_3213;
assign n_3217 = n_3214 ^ x77;
assign n_3218 = ~n_3215 & ~n_3216;
assign n_3219 = n_3218 ^ x78;
assign n_3220 = n_3219 ^ x79;
assign n_3221 = n_3126 ^ n_3219;
assign n_3222 = n_3220 & n_3221;
assign n_3223 = n_3222 ^ x79;
assign n_3224 = n_3223 ^ x80;
assign n_3225 = n_3127 ^ n_3223;
assign n_3226 = n_3224 & n_3225;
assign n_3227 = n_3226 ^ x80;
assign n_3228 = n_3227 ^ x81;
assign n_3229 = n_3128 ^ n_3227;
assign n_3230 = n_3228 & n_3229;
assign n_3231 = n_3230 ^ x81;
assign n_3232 = n_3231 ^ x82;
assign n_3233 = n_3129 ^ n_3231;
assign n_3234 = n_3232 & n_3233;
assign n_3235 = n_3234 ^ x82;
assign n_3236 = n_3235 ^ x83;
assign n_3237 = n_3130 ^ n_3235;
assign n_3238 = n_3236 & n_3237;
assign n_3239 = n_3238 ^ x83;
assign n_3240 = n_3239 ^ x84;
assign n_3241 = n_3131 ^ n_3239;
assign n_3242 = n_3240 & n_3241;
assign n_3243 = n_3242 ^ x84;
assign n_3244 = n_3243 ^ x85;
assign n_3245 = n_3132 ^ n_3243;
assign n_3246 = n_3244 & n_3245;
assign n_3247 = n_3246 ^ x85;
assign n_3248 = n_3247 ^ x86;
assign n_3249 = n_3133 ^ n_3247;
assign n_3250 = n_3248 & n_3249;
assign n_3251 = n_3250 ^ x86;
assign n_3252 = n_3251 ^ x87;
assign n_3253 = n_3134 ^ n_3251;
assign n_3254 = n_3252 & n_3253;
assign n_3255 = n_3254 ^ x87;
assign n_3256 = n_3255 ^ x88;
assign n_3257 = n_3135 ^ n_3255;
assign n_3258 = n_3256 & n_3257;
assign n_3259 = n_3258 ^ x88;
assign n_3260 = n_3259 ^ x89;
assign n_3261 = n_3139 ^ n_3259;
assign n_3262 = n_3260 & n_3261;
assign n_3263 = n_3262 ^ x89;
assign n_3264 = n_3263 ^ x90;
assign n_3265 = n_3263 ^ n_3110;
assign n_3266 = n_3160 & n_3263;
assign n_3267 = n_3264 & n_3265;
assign n_3268 = ~n_3166 & ~n_3266;
assign n_3269 = n_3267 ^ x90;
assign n_3270 = x92 ^ n_3268;
assign n_3271 = n_3136 ^ n_3268;
assign n_3272 = n_3269 ^ x91;
assign n_3273 = ~n_3270 & ~n_3271;
assign n_3274 = n_3273 ^ x92;
assign n_3275 = n_376 & ~n_3274;
assign n_3276 = n_3274 ^ x93;
assign n_3277 = ~n_3275 & n_3150;
assign n_3278 = n_3151 & n_3276;
assign n_3279 = ~x94 & n_3277;
assign n_3280 = n_3278 ^ x93;
assign n_3281 = x93 ^ ~n_3279;
assign n_3282 = n_376 & ~n_3280;
assign n_3283 = ~n_3270 & n_3282;
assign n_3284 = n_3236 & n_3282;
assign n_3285 = n_3232 & n_3282;
assign n_3286 = x65 & n_3282;
assign n_3287 = x64 & n_3282;
assign n_3288 = n_3169 & n_3282;
assign n_3289 = n_3173 & n_3282;
assign n_3290 = n_3177 & n_3282;
assign n_3291 = n_3181 & n_3282;
assign n_3292 = n_3185 & n_3282;
assign n_3293 = n_3189 & n_3282;
assign n_3294 = n_3193 & n_3282;
assign n_3295 = n_3197 & n_3282;
assign n_3296 = n_3201 & n_3282;
assign n_3297 = n_3205 & n_3282;
assign n_3298 = n_3209 & n_3282;
assign n_3299 = ~n_3215 & n_3282;
assign n_3300 = n_3220 & n_3282;
assign n_3301 = n_3224 & n_3282;
assign n_3302 = n_3228 & n_3282;
assign n_3303 = n_3240 & n_3282;
assign n_3304 = n_3244 & n_3282;
assign n_3305 = n_3248 & n_3282;
assign n_3306 = n_3252 & n_3282;
assign n_3307 = n_3256 & n_3282;
assign n_3308 = n_3260 & n_3282;
assign n_3309 = n_3264 & n_3282;
assign y34 = n_3282;
assign n_3310 = n_3217 & n_3282;
assign n_3311 = n_3272 & n_3282;
assign n_3312 = n_3283 ^ n_3136;
assign n_3313 = n_3284 ^ n_3130;
assign n_3314 = n_3285 ^ n_3129;
assign n_3315 = n_3286 ^ n_3282;
assign n_3316 = n_3116 ^ n_3286;
assign n_3317 = n_3287 ^ x33;
assign n_3318 = n_3287 ^ x34;
assign n_3319 = n_3288 ^ n_3165;
assign n_3320 = n_3289 ^ n_3117;
assign n_3321 = n_3290 ^ n_3118;
assign n_3322 = n_3291 ^ n_3119;
assign n_3323 = n_3292 ^ n_3138;
assign n_3324 = n_3293 ^ n_3120;
assign n_3325 = n_3294 ^ n_3121;
assign n_3326 = n_3295 ^ n_3122;
assign n_3327 = n_3296 ^ n_3123;
assign n_3328 = n_3297 ^ n_3124;
assign n_3329 = n_3298 ^ n_3112;
assign n_3330 = n_3299 ^ n_3125;
assign n_3331 = n_3300 ^ n_3126;
assign n_3332 = n_3301 ^ n_3127;
assign n_3333 = n_3302 ^ n_3128;
assign n_3334 = n_3303 ^ n_3131;
assign n_3335 = n_3304 ^ n_3132;
assign n_3336 = n_3305 ^ n_3133;
assign n_3337 = n_3306 ^ n_3134;
assign n_3338 = n_3307 ^ n_3135;
assign n_3339 = n_3308 ^ n_3139;
assign n_3340 = n_3309 ^ n_3110;
assign n_3341 = n_3111 ^ n_3310;
assign n_3342 = n_3109 ^ n_3311;
assign n_3343 = ~x93 ^ n_3312;
assign n_3344 = ~n_3312 & ~n_3281;
assign n_3345 = ~x84 ^ n_3313;
assign n_3346 = n_3313 ^ x84;
assign n_3347 = n_3314 ^ x83;
assign n_3348 = x83 & ~n_3314;
assign n_3349 = n_206 & ~n_3315;
assign n_3350 = n_3287 & n_3318;
assign n_3351 = n_3343 & ~n_3279;
assign n_3352 = ~n_3344 & ~n_3159;
assign n_3353 = n_3347 ^ n_3348;
assign n_3354 = n_3348 ^ n_3313;
assign n_3355 = n_3350 ^ n_3287;
assign n_3356 = n_3316 ^ n_3350;
assign n_3357 = n_3345 & ~n_3353;
assign n_3358 = ~n_3346 & n_3354;
assign n_3359 = ~n_3317 & n_3355;
assign n_3360 = n_3358 ^ x84;
assign n_3361 = n_3359 ^ n_3350;
assign n_3362 = n_3361 ^ n_3287;
assign n_3363 = n_3362 ^ n_3318;
assign n_3364 = ~x65 & ~n_3363;
assign n_3365 = n_3318 ^ n_3364;
assign n_3366 = n_3365 & ~n_3349;
assign n_3367 = x66 ^ n_3366;
assign n_3368 = n_3356 ^ n_3366;
assign n_3369 = ~n_3367 & ~n_3368;
assign n_3370 = n_3369 ^ x66;
assign n_3371 = n_3370 ^ x67;
assign n_3372 = n_3319 ^ n_3370;
assign n_3373 = n_3371 & n_3372;
assign n_3374 = n_3373 ^ x67;
assign n_3375 = n_3374 ^ x68;
assign n_3376 = n_3320 ^ n_3374;
assign n_3377 = n_3375 & n_3376;
assign n_3378 = n_3377 ^ x68;
assign n_3379 = n_3378 ^ x69;
assign n_3380 = n_3321 ^ n_3378;
assign n_3381 = n_3379 & n_3380;
assign n_3382 = n_3381 ^ x69;
assign n_3383 = n_3382 ^ x70;
assign n_3384 = n_3322 ^ n_3382;
assign n_3385 = n_3383 & n_3384;
assign n_3386 = n_3385 ^ x70;
assign n_3387 = n_3386 ^ x71;
assign n_3388 = n_3323 ^ n_3386;
assign n_3389 = n_3387 & n_3388;
assign n_3390 = n_3389 ^ x71;
assign n_3391 = n_3390 ^ x72;
assign n_3392 = n_3324 ^ n_3390;
assign n_3393 = n_3391 & n_3392;
assign n_3394 = n_3393 ^ x72;
assign n_3395 = n_3394 ^ x73;
assign n_3396 = n_3325 ^ n_3394;
assign n_3397 = n_3395 & n_3396;
assign n_3398 = n_3397 ^ x73;
assign n_3399 = n_3398 ^ x74;
assign n_3400 = n_3326 ^ n_3398;
assign n_3401 = n_3399 & n_3400;
assign n_3402 = n_3401 ^ x74;
assign n_3403 = n_3402 ^ x75;
assign n_3404 = n_3327 ^ n_3402;
assign n_3405 = n_3403 & n_3404;
assign n_3406 = n_3405 ^ x75;
assign n_3407 = n_3406 ^ x76;
assign n_3408 = n_3328 ^ n_3406;
assign n_3409 = n_3407 & n_3408;
assign n_3410 = n_3409 ^ x76;
assign n_3411 = n_3410 ^ x77;
assign n_3412 = n_3329 ^ n_3410;
assign n_3413 = n_3411 & n_3412;
assign n_3414 = n_3413 ^ x77;
assign n_3415 = n_3414 ^ x78;
assign n_3416 = n_3341 ^ n_3414;
assign n_3417 = n_3415 & n_3416;
assign n_3418 = n_3417 ^ x78;
assign n_3419 = n_3418 ^ x79;
assign n_3420 = n_3330 ^ n_3418;
assign n_3421 = n_3419 & n_3420;
assign n_3422 = n_3421 ^ x79;
assign n_3423 = n_3422 ^ x80;
assign n_3424 = n_3331 ^ n_3422;
assign n_3425 = n_3423 & n_3424;
assign n_3426 = n_3425 ^ x80;
assign n_3427 = n_3426 ^ x81;
assign n_3428 = n_3332 ^ n_3426;
assign n_3429 = n_3427 & n_3428;
assign n_3430 = n_3429 ^ x81;
assign n_3431 = n_3430 ^ x82;
assign n_3432 = n_3333 ^ n_3430;
assign n_3433 = n_3431 & n_3432;
assign n_3434 = n_3433 ^ x82;
assign n_3435 = n_3434 ^ x83;
assign n_3436 = n_3434 ^ n_3314;
assign n_3437 = n_3357 & n_3434;
assign n_3438 = n_3435 & n_3436;
assign n_3439 = ~n_3360 & ~n_3437;
assign n_3440 = n_3438 ^ x83;
assign n_3441 = x85 ^ n_3439;
assign n_3442 = n_3334 ^ n_3439;
assign n_3443 = n_3440 ^ x84;
assign n_3444 = ~n_3441 & ~n_3442;
assign n_3445 = n_3444 ^ x85;
assign n_3446 = n_3445 ^ x86;
assign n_3447 = n_3335 ^ n_3445;
assign n_3448 = n_3446 & n_3447;
assign n_3449 = n_3448 ^ x86;
assign n_3450 = n_3449 ^ x87;
assign n_3451 = n_3336 ^ n_3449;
assign n_3452 = n_3450 & n_3451;
assign n_3453 = n_3452 ^ x87;
assign n_3454 = n_3453 ^ x88;
assign n_3455 = n_3337 ^ n_3453;
assign n_3456 = n_3454 & n_3455;
assign n_3457 = n_3456 ^ x88;
assign n_3458 = n_3457 ^ x89;
assign n_3459 = n_3338 ^ n_3457;
assign n_3460 = n_3458 & n_3459;
assign n_3461 = n_3460 ^ x89;
assign n_3462 = n_3461 ^ x90;
assign n_3463 = n_3339 ^ n_3461;
assign n_3464 = n_3462 & n_3463;
assign n_3465 = n_3464 ^ x90;
assign n_3466 = n_3465 ^ x91;
assign n_3467 = n_3340 ^ n_3465;
assign n_3468 = n_3466 & n_3467;
assign n_3469 = n_3468 ^ x91;
assign n_3470 = n_3469 ^ x92;
assign n_3471 = n_3342 ^ n_3469;
assign n_3472 = n_3470 & n_3471;
assign n_3473 = n_3472 ^ x92;
assign n_3474 = n_3473 ^ x93;
assign n_3475 = n_3351 & n_3473;
assign n_3476 = ~n_3475 & n_3352;
assign n_3477 = n_3277 & ~n_3476;
assign n_3478 = ~n_3441 & n_3476;
assign n_3479 = n_149 & n_3476;
assign n_3480 = x64 & n_3476;
assign n_3481 = ~n_3367 & n_3476;
assign n_3482 = n_3371 & n_3476;
assign n_3483 = n_3375 & n_3476;
assign n_3484 = n_3379 & n_3476;
assign n_3485 = n_3383 & n_3476;
assign n_3486 = n_3387 & n_3476;
assign n_3487 = n_3391 & n_3476;
assign n_3488 = n_3395 & n_3476;
assign n_3489 = n_3399 & n_3476;
assign n_3490 = n_3403 & n_3476;
assign n_3491 = n_3407 & n_3476;
assign n_3492 = n_3411 & n_3476;
assign n_3493 = n_3415 & n_3476;
assign n_3494 = n_3419 & n_3476;
assign n_3495 = n_3423 & n_3476;
assign n_3496 = n_3427 & n_3476;
assign n_3497 = n_3431 & n_3476;
assign n_3498 = n_3435 & n_3476;
assign n_3499 = n_3446 & n_3476;
assign n_3500 = n_3450 & n_3476;
assign n_3501 = n_3454 & n_3476;
assign n_3502 = n_3458 & n_3476;
assign n_3503 = n_3462 & n_3476;
assign n_3504 = n_3466 & n_3476;
assign n_3505 = n_3470 & n_3476;
assign n_3506 = n_3474 & n_3476;
assign y33 = n_3476;
assign n_3507 = n_3443 & n_3476;
assign n_3508 = ~n_439 ^ ~n_3477;
assign n_3509 = n_3478 ^ n_3334;
assign n_3510 = n_3479 ^ n_3287;
assign n_3511 = n_3480 ^ x32;
assign n_3512 = n_3480 ^ n_46;
assign n_3513 = n_3481 ^ n_3356;
assign n_3514 = n_3482 ^ n_3319;
assign n_3515 = n_3483 ^ n_3320;
assign n_3516 = n_3484 ^ n_3321;
assign n_3517 = n_3485 ^ n_3322;
assign n_3518 = n_3486 ^ n_3323;
assign n_3519 = n_3487 ^ n_3324;
assign n_3520 = n_3488 ^ n_3325;
assign n_3521 = n_3489 ^ n_3326;
assign n_3522 = n_3490 ^ n_3327;
assign n_3523 = n_3491 ^ n_3328;
assign n_3524 = n_3492 ^ n_3329;
assign n_3525 = n_3493 ^ n_3341;
assign n_3526 = n_3494 ^ n_3330;
assign n_3527 = n_3495 ^ n_3331;
assign n_3528 = n_3496 ^ n_3332;
assign n_3529 = n_3497 ^ n_3333;
assign n_3530 = n_3498 ^ n_3314;
assign n_3531 = n_3499 ^ n_3335;
assign n_3532 = n_3500 ^ n_3336;
assign n_3533 = n_3501 ^ n_3337;
assign n_3534 = n_3502 ^ n_3338;
assign n_3535 = n_3503 ^ n_3339;
assign n_3536 = n_3504 ^ n_3340;
assign n_3537 = n_3505 ^ n_3342;
assign n_3538 = n_3506 ^ n_3312;
assign n_3539 = n_3313 ^ n_3507;
assign n_3540 = ~n_3508 ^ x95;
assign n_3541 = ~x86 ^ n_3509;
assign n_3542 = n_3509 ^ x86;
assign n_3543 = n_3510 ^ x34;
assign n_3544 = ~n_3511 & n_3512;
assign n_3545 = n_3539 ^ x85;
assign n_3546 = x85 & ~n_3539;
assign n_3547 = n_3543 ^ x66;
assign n_3548 = n_3544 ^ x65;
assign n_3549 = n_3545 ^ n_3546;
assign n_3550 = n_3546 ^ n_3509;
assign n_3551 = n_3548 ^ n_297;
assign n_3552 = n_3541 & ~n_3549;
assign n_3553 = ~n_3542 & n_3550;
assign n_3554 = n_3551 ^ n_3543;
assign n_3555 = n_3551 ^ x66;
assign n_3556 = n_3553 ^ x86;
assign n_3557 = ~n_3547 & n_3554;
assign n_3558 = n_3557 ^ x66;
assign n_3559 = n_3558 ^ x67;
assign n_3560 = n_3513 ^ n_3558;
assign n_3561 = n_3559 & n_3560;
assign n_3562 = n_3561 ^ x67;
assign n_3563 = n_3562 ^ x68;
assign n_3564 = n_3514 ^ n_3562;
assign n_3565 = n_3563 & n_3564;
assign n_3566 = n_3565 ^ x68;
assign n_3567 = n_3566 ^ x69;
assign n_3568 = n_3515 ^ n_3566;
assign n_3569 = n_3567 & n_3568;
assign n_3570 = n_3569 ^ x69;
assign n_3571 = n_3570 ^ x70;
assign n_3572 = n_3516 ^ n_3570;
assign n_3573 = n_3571 & n_3572;
assign n_3574 = n_3573 ^ x70;
assign n_3575 = n_3574 ^ x71;
assign n_3576 = n_3517 ^ n_3574;
assign n_3577 = n_3575 & n_3576;
assign n_3578 = n_3577 ^ x71;
assign n_3579 = n_3578 ^ x72;
assign n_3580 = n_3518 ^ n_3578;
assign n_3581 = n_3579 & n_3580;
assign n_3582 = n_3581 ^ x72;
assign n_3583 = n_3582 ^ x73;
assign n_3584 = n_3519 ^ n_3582;
assign n_3585 = n_3583 & n_3584;
assign n_3586 = n_3585 ^ x73;
assign n_3587 = n_3586 ^ x74;
assign n_3588 = n_3520 ^ n_3586;
assign n_3589 = n_3587 & n_3588;
assign n_3590 = n_3589 ^ x74;
assign n_3591 = n_3590 ^ x75;
assign n_3592 = n_3521 ^ n_3590;
assign n_3593 = n_3591 & n_3592;
assign n_3594 = n_3593 ^ x75;
assign n_3595 = n_3594 ^ x76;
assign n_3596 = n_3522 ^ n_3594;
assign n_3597 = n_3595 & n_3596;
assign n_3598 = n_3597 ^ x76;
assign n_3599 = n_3598 ^ x77;
assign n_3600 = n_3523 ^ n_3598;
assign n_3601 = n_3599 & n_3600;
assign n_3602 = n_3601 ^ x77;
assign n_3603 = n_3602 ^ x78;
assign n_3604 = n_3524 ^ n_3602;
assign n_3605 = n_3603 & n_3604;
assign n_3606 = n_3605 ^ x78;
assign n_3607 = n_3606 ^ x79;
assign n_3608 = n_3525 ^ n_3606;
assign n_3609 = n_3607 & n_3608;
assign n_3610 = n_3609 ^ x79;
assign n_3611 = n_3610 ^ x80;
assign n_3612 = n_3526 ^ n_3610;
assign n_3613 = n_3611 & n_3612;
assign n_3614 = n_3613 ^ x80;
assign n_3615 = n_3614 ^ x81;
assign n_3616 = n_3527 ^ n_3614;
assign n_3617 = n_3615 & n_3616;
assign n_3618 = n_3617 ^ x81;
assign n_3619 = n_3618 ^ x82;
assign n_3620 = n_3528 ^ n_3618;
assign n_3621 = n_3619 & n_3620;
assign n_3622 = n_3621 ^ x82;
assign n_3623 = n_3622 ^ x83;
assign n_3624 = n_3529 ^ n_3622;
assign n_3625 = n_3623 & n_3624;
assign n_3626 = n_3625 ^ x83;
assign n_3627 = n_3626 ^ x84;
assign n_3628 = n_3530 ^ n_3626;
assign n_3629 = n_3627 & n_3628;
assign n_3630 = n_3629 ^ x84;
assign n_3631 = n_3630 ^ x85;
assign n_3632 = n_3630 ^ n_3539;
assign n_3633 = n_3552 & n_3630;
assign n_3634 = n_3631 & n_3632;
assign n_3635 = ~n_3556 & ~n_3633;
assign n_3636 = n_3634 ^ x85;
assign n_3637 = x87 ^ n_3635;
assign n_3638 = n_3531 ^ n_3635;
assign n_3639 = n_3636 ^ x86;
assign n_3640 = ~n_3637 & ~n_3638;
assign n_3641 = n_3640 ^ x87;
assign n_3642 = n_3641 ^ x88;
assign n_3643 = n_3532 ^ n_3641;
assign n_3644 = n_3642 & n_3643;
assign n_3645 = n_3644 ^ x88;
assign n_3646 = n_3645 ^ x89;
assign n_3647 = n_3533 ^ n_3645;
assign n_3648 = n_3646 & n_3647;
assign n_3649 = n_3648 ^ x89;
assign n_3650 = n_3649 ^ x90;
assign n_3651 = n_3534 ^ n_3649;
assign n_3652 = n_3650 & n_3651;
assign n_3653 = n_3652 ^ x90;
assign n_3654 = n_3653 ^ x91;
assign n_3655 = n_3535 ^ n_3653;
assign n_3656 = n_3654 & n_3655;
assign n_3657 = n_3656 ^ x91;
assign n_3658 = n_3657 ^ x92;
assign n_3659 = n_3536 ^ n_3657;
assign n_3660 = n_3658 & n_3659;
assign n_3661 = n_3660 ^ x92;
assign n_3662 = n_3661 ^ x93;
assign n_3663 = n_3537 ^ n_3661;
assign n_3664 = n_3662 & n_3663;
assign n_3665 = n_3664 ^ x93;
assign n_3666 = n_3665 ^ x94;
assign n_3667 = n_3538 ^ n_3665;
assign n_3668 = n_3666 & ~n_3667;
assign n_3669 = n_3668 ^ n_3665;
assign n_3670 = n_3669 ^ x95;
assign n_3671 = n_3540 & n_3670;
assign n_3672 = x95 ^ n_3671;
assign n_3673 = n_374 & ~n_3672;
assign n_3674 = n_3508 & ~n_3673;
assign n_3675 = n_3607 & n_3673;
assign n_3676 = n_3603 & n_3673;
assign n_3677 = n_251 & n_3673;
assign n_3678 = x65 ^ n_3673;
assign n_3679 = n_3555 & n_3673;
assign n_3680 = n_3559 & n_3673;
assign n_3681 = n_3563 & n_3673;
assign n_3682 = n_3567 & n_3673;
assign n_3683 = n_3571 & n_3673;
assign n_3684 = n_3575 & n_3673;
assign n_3685 = n_3579 & n_3673;
assign n_3686 = n_3583 & n_3673;
assign n_3687 = n_3587 & n_3673;
assign n_3688 = n_3591 & n_3673;
assign n_3689 = n_3595 & n_3673;
assign n_3690 = n_3599 & n_3673;
assign n_3691 = n_3611 & n_3673;
assign n_3692 = n_3615 & n_3673;
assign n_3693 = n_3619 & n_3673;
assign n_3694 = n_3623 & n_3673;
assign n_3695 = n_3627 & n_3673;
assign n_3696 = n_3631 & n_3673;
assign n_3697 = ~n_3637 & n_3673;
assign n_3698 = n_3642 & n_3673;
assign n_3699 = n_3646 & n_3673;
assign n_3700 = n_3650 & n_3673;
assign n_3701 = n_3654 & n_3673;
assign n_3702 = n_3658 & n_3673;
assign n_3703 = n_3662 & n_3673;
assign n_3704 = n_3666 & n_3673;
assign n_3705 = x64 & ~n_3673;
assign y32 = n_3673;
assign n_3706 = ~n_275 & n_3673;
assign n_3707 = n_3639 & n_3673;
assign n_3708 = ~n_439 ^ ~n_3674;
assign n_3709 = n_3675 ^ n_3525;
assign n_3710 = n_3676 ^ n_3524;
assign n_3711 = n_3677 ^ n_3480;
assign n_3712 = n_19 & ~n_3678;
assign n_3713 = n_3679 ^ n_3543;
assign n_3714 = n_3680 ^ n_3513;
assign n_3715 = n_3681 ^ n_3514;
assign n_3716 = n_3682 ^ n_3515;
assign n_3717 = n_3683 ^ n_3516;
assign n_3718 = n_3684 ^ n_3517;
assign n_3719 = n_3685 ^ n_3518;
assign n_3720 = n_3686 ^ n_3519;
assign n_3721 = n_3687 ^ n_3520;
assign n_3722 = n_3688 ^ n_3521;
assign n_3723 = n_3689 ^ n_3522;
assign n_3724 = n_3690 ^ n_3523;
assign n_3725 = n_3691 ^ n_3526;
assign n_3726 = n_3692 ^ n_3527;
assign n_3727 = n_3693 ^ n_3528;
assign n_3728 = n_3694 ^ n_3529;
assign n_3729 = n_3695 ^ n_3530;
assign n_3730 = n_3696 ^ n_3539;
assign n_3731 = n_3697 ^ n_3531;
assign n_3732 = n_3698 ^ n_3532;
assign n_3733 = n_3699 ^ n_3533;
assign n_3734 = n_3700 ^ n_3534;
assign n_3735 = n_3701 ^ n_3535;
assign n_3736 = n_3702 ^ n_3536;
assign n_3737 = n_3703 ^ n_3537;
assign n_3738 = n_3704 ^ n_3538;
assign n_3739 = x32 ^ n_3706;
assign n_3740 = n_3509 ^ n_3707;
assign n_3741 = ~n_3708 ^ x96;
assign n_3742 = x96 & ~n_3708;
assign n_3743 = x97 & ~n_3708;
assign n_3744 = ~x80 ^ n_3709;
assign n_3745 = n_3709 ^ x80;
assign n_3746 = n_3710 ^ x79;
assign n_3747 = x79 & ~n_3710;
assign n_3748 = n_3711 ^ x33;
assign n_3749 = n_3712 ^ n_3673;
assign n_3750 = ~x95 & n_3738;
assign n_3751 = ~n_3738 & n_124;
assign n_3752 = n_3739 ^ x65;
assign n_3753 = n_3741 ^ n_3742;
assign n_3754 = n_373 & ~n_3742;
assign n_3755 = n_3743 ^ x97;
assign n_3756 = n_372 & ~n_3743;
assign n_3757 = n_3746 ^ n_3747;
assign n_3758 = n_3747 ^ n_3709;
assign n_3759 = n_3748 ^ x66;
assign n_3760 = n_252 ^ n_3749;
assign n_3761 = x96 & ~n_3750;
assign n_3762 = n_373 & ~n_3751;
assign n_3763 = ~n_3750 & n_3753;
assign n_3764 = x95 & n_3753;
assign n_3765 = n_3744 & ~n_3757;
assign n_3766 = ~n_3745 & n_3758;
assign n_3767 = n_3739 & n_3760;
assign n_3768 = ~n_3738 & n_3764;
assign n_3769 = n_3766 ^ x80;
assign n_3770 = n_3767 ^ n_3749;
assign n_3771 = n_3754 & ~n_3768;
assign n_3772 = ~n_3752 & n_3770;
assign n_3773 = x65 ^ n_3772;
assign n_3774 = n_3773 ^ n_3748;
assign n_3775 = n_3773 ^ x66;
assign n_3776 = ~n_3759 & n_3774;
assign n_3777 = n_3776 ^ x66;
assign n_3778 = n_3777 ^ x67;
assign n_3779 = n_3713 ^ n_3777;
assign n_3780 = n_3778 & n_3779;
assign n_3781 = n_3780 ^ x67;
assign n_3782 = n_3781 ^ x68;
assign n_3783 = n_3714 ^ n_3781;
assign n_3784 = n_3782 & n_3783;
assign n_3785 = n_3784 ^ x68;
assign n_3786 = n_3785 ^ x69;
assign n_3787 = n_3715 ^ n_3785;
assign n_3788 = n_3786 & n_3787;
assign n_3789 = n_3788 ^ x69;
assign n_3790 = n_3789 ^ x70;
assign n_3791 = n_3716 ^ n_3789;
assign n_3792 = n_3790 & n_3791;
assign n_3793 = n_3792 ^ x70;
assign n_3794 = n_3793 ^ x71;
assign n_3795 = n_3717 ^ n_3793;
assign n_3796 = n_3794 & n_3795;
assign n_3797 = n_3796 ^ x71;
assign n_3798 = n_3797 ^ x72;
assign n_3799 = n_3718 ^ n_3797;
assign n_3800 = n_3798 & n_3799;
assign n_3801 = n_3800 ^ x72;
assign n_3802 = n_3801 ^ x73;
assign n_3803 = n_3719 ^ n_3801;
assign n_3804 = n_3802 & n_3803;
assign n_3805 = n_3804 ^ x73;
assign n_3806 = n_3805 ^ x74;
assign n_3807 = n_3720 ^ n_3805;
assign n_3808 = n_3806 & n_3807;
assign n_3809 = n_3808 ^ x74;
assign n_3810 = n_3809 ^ x75;
assign n_3811 = n_3721 ^ n_3809;
assign n_3812 = n_3810 & n_3811;
assign n_3813 = n_3812 ^ x75;
assign n_3814 = n_3813 ^ x76;
assign n_3815 = n_3722 ^ n_3813;
assign n_3816 = n_3814 & n_3815;
assign n_3817 = n_3816 ^ x76;
assign n_3818 = n_3817 ^ x77;
assign n_3819 = n_3723 ^ n_3817;
assign n_3820 = n_3818 & n_3819;
assign n_3821 = n_3820 ^ x77;
assign n_3822 = n_3821 ^ x78;
assign n_3823 = n_3724 ^ n_3821;
assign n_3824 = n_3822 & n_3823;
assign n_3825 = n_3824 ^ x78;
assign n_3826 = n_3825 ^ x79;
assign n_3827 = n_3825 ^ n_3710;
assign n_3828 = n_3765 & n_3825;
assign n_3829 = n_3826 & n_3827;
assign n_3830 = ~n_3769 & ~n_3828;
assign n_3831 = n_3829 ^ x79;
assign n_3832 = x81 ^ n_3830;
assign n_3833 = n_3725 ^ n_3830;
assign n_3834 = n_3831 ^ x80;
assign n_3835 = ~n_3832 & ~n_3833;
assign n_3836 = n_3835 ^ x81;
assign n_3837 = n_3836 ^ x82;
assign n_3838 = n_3726 ^ n_3836;
assign n_3839 = n_3837 & n_3838;
assign n_3840 = n_3839 ^ x82;
assign n_3841 = n_3840 ^ x83;
assign n_3842 = n_3727 ^ n_3840;
assign n_3843 = n_3841 & n_3842;
assign n_3844 = n_3843 ^ x83;
assign n_3845 = n_3844 ^ x84;
assign n_3846 = n_3728 ^ n_3844;
assign n_3847 = n_3845 & n_3846;
assign n_3848 = n_3847 ^ x84;
assign n_3849 = n_3848 ^ x85;
assign n_3850 = n_3729 ^ n_3848;
assign n_3851 = n_3849 & n_3850;
assign n_3852 = n_3851 ^ x85;
assign n_3853 = n_3852 ^ x86;
assign n_3854 = n_3730 ^ n_3852;
assign n_3855 = n_3853 & n_3854;
assign n_3856 = n_3855 ^ x86;
assign n_3857 = n_3856 ^ x87;
assign n_3858 = n_3740 ^ n_3856;
assign n_3859 = n_3857 & n_3858;
assign n_3860 = n_3859 ^ x87;
assign n_3861 = n_3860 ^ x88;
assign n_3862 = n_3731 ^ n_3860;
assign n_3863 = n_3861 & n_3862;
assign n_3864 = n_3863 ^ x88;
assign n_3865 = n_3864 ^ x89;
assign n_3866 = n_3732 ^ n_3864;
assign n_3867 = n_3865 & n_3866;
assign n_3868 = n_3867 ^ x89;
assign n_3869 = n_3868 ^ x90;
assign n_3870 = n_3733 ^ n_3868;
assign n_3871 = n_3869 & n_3870;
assign n_3872 = n_3871 ^ x90;
assign n_3873 = n_3872 ^ x91;
assign n_3874 = n_3734 ^ n_3872;
assign n_3875 = n_3873 & n_3874;
assign n_3876 = n_3875 ^ x91;
assign n_3877 = n_3876 ^ x92;
assign n_3878 = n_3735 ^ n_3876;
assign n_3879 = n_3877 & n_3878;
assign n_3880 = n_3879 ^ x92;
assign n_3881 = n_3880 ^ x93;
assign n_3882 = n_3736 ^ n_3880;
assign n_3883 = n_3881 & n_3882;
assign n_3884 = n_3883 ^ x93;
assign n_3885 = n_3884 ^ x94;
assign n_3886 = n_3737 ^ n_3884;
assign n_3887 = n_3885 & n_3886;
assign n_3888 = n_3887 ^ x94;
assign n_3889 = n_3888 ^ x95;
assign n_3890 = n_3888 & n_3761;
assign n_3891 = n_3888 & n_3763;
assign n_3892 = ~n_3890 & n_3762;
assign n_3893 = ~n_3891 & n_3771;
assign n_3894 = n_3708 & ~n_3892;
assign n_3895 = x64 ^ n_3893;
assign n_3896 = ~x65 & n_3893;
assign n_3897 = x64 & n_3893;
assign n_3898 = ~x30 & n_3893;
assign n_3899 = n_3775 & n_3893;
assign n_3900 = n_3778 & n_3893;
assign n_3901 = n_3782 & n_3893;
assign n_3902 = n_3786 & n_3893;
assign n_3903 = n_3790 & n_3893;
assign n_3904 = n_3794 & n_3893;
assign n_3905 = n_3798 & n_3893;
assign n_3906 = n_3802 & n_3893;
assign n_3907 = n_3806 & n_3893;
assign n_3908 = n_3810 & n_3893;
assign n_3909 = n_3814 & n_3893;
assign n_3910 = n_3818 & n_3893;
assign n_3911 = n_3822 & n_3893;
assign n_3912 = n_3826 & n_3893;
assign n_3913 = ~n_3832 & n_3893;
assign n_3914 = n_3837 & n_3893;
assign n_3915 = n_3841 & n_3893;
assign n_3916 = n_3845 & n_3893;
assign n_3917 = n_3849 & n_3893;
assign n_3918 = n_3853 & n_3893;
assign n_3919 = n_3857 & n_3893;
assign n_3920 = n_3861 & n_3893;
assign n_3921 = n_3865 & n_3893;
assign n_3922 = n_3869 & n_3893;
assign n_3923 = n_3873 & n_3893;
assign n_3924 = n_3877 & n_3893;
assign n_3925 = n_3881 & n_3893;
assign n_3926 = n_3885 & n_3893;
assign n_3927 = n_3889 & n_3893;
assign y31 = n_3893;
assign n_3928 = n_3834 & n_3893;
assign n_3929 = ~n_439 ^ ~n_3894;
assign n_3930 = ~n_19 & ~n_3895;
assign n_3931 = ~x30 & n_3895;
assign n_3932 = x65 & ~n_3897;
assign n_3933 = n_3897 ^ x31;
assign n_3934 = n_77 ^ n_3898;
assign n_3935 = n_3898 ^ x65;
assign n_3936 = n_3899 ^ n_3748;
assign n_3937 = n_3900 ^ n_3713;
assign n_3938 = n_3901 ^ n_3714;
assign n_3939 = n_3902 ^ n_3715;
assign n_3940 = n_3903 ^ n_3716;
assign n_3941 = n_3904 ^ n_3717;
assign n_3942 = n_3905 ^ n_3718;
assign n_3943 = n_3906 ^ n_3719;
assign n_3944 = n_3907 ^ n_3720;
assign n_3945 = n_3908 ^ n_3721;
assign n_3946 = n_3909 ^ n_3722;
assign n_3947 = n_3910 ^ n_3723;
assign n_3948 = n_3911 ^ n_3724;
assign n_3949 = n_3912 ^ n_3710;
assign n_3950 = n_3913 ^ n_3725;
assign n_3951 = n_3914 ^ n_3726;
assign n_3952 = n_3915 ^ n_3727;
assign n_3953 = n_3916 ^ n_3728;
assign n_3954 = n_3917 ^ n_3729;
assign n_3955 = n_3918 ^ n_3730;
assign n_3956 = n_3919 ^ n_3740;
assign n_3957 = n_3920 ^ n_3731;
assign n_3958 = n_3921 ^ n_3732;
assign n_3959 = n_3922 ^ n_3733;
assign n_3960 = n_3923 ^ n_3734;
assign n_3961 = n_3924 ^ n_3735;
assign n_3962 = n_3925 ^ n_3736;
assign n_3963 = n_3926 ^ n_3737;
assign n_3964 = n_3927 ^ n_3738;
assign n_3965 = n_3709 ^ n_3928;
assign n_3966 = ~n_3929 ^ x98;
assign n_3967 = ~x98 & n_3929;
assign n_3968 = n_3755 ^ ~n_3929;
assign n_3969 = n_3930 ^ n_3705;
assign n_3970 = n_208 ^ n_3932;
assign n_3971 = x64 & n_3934;
assign n_3972 = n_3931 ^ n_3935;
assign n_3973 = n_3966 ^ n_3967;
assign n_3974 = n_3969 ^ n_3896;
assign n_3975 = n_152 ^ n_3971;
assign n_3976 = n_371 & n_3973;
assign n_3977 = n_3974 ^ x32;
assign n_3978 = n_3970 ^ n_3975;
assign n_3979 = n_3977 ^ x66;
assign n_3980 = n_3978 ^ n_3977;
assign n_3981 = n_3978 ^ x66;
assign n_3982 = n_3979 & ~n_3980;
assign n_3983 = n_3982 ^ x66;
assign n_3984 = n_3983 ^ x67;
assign n_3985 = n_3936 ^ n_3983;
assign n_3986 = n_3984 & n_3985;
assign n_3987 = n_3986 ^ x67;
assign n_3988 = n_3987 ^ x68;
assign n_3989 = n_3937 ^ n_3987;
assign n_3990 = n_3988 & n_3989;
assign n_3991 = n_3990 ^ x68;
assign n_3992 = n_3991 ^ x69;
assign n_3993 = n_3938 ^ n_3991;
assign n_3994 = n_3992 & n_3993;
assign n_3995 = n_3994 ^ x69;
assign n_3996 = n_3995 ^ x70;
assign n_3997 = n_3939 ^ n_3995;
assign n_3998 = n_3996 & n_3997;
assign n_3999 = n_3998 ^ x70;
assign n_4000 = n_3999 ^ x71;
assign n_4001 = n_3940 ^ n_3999;
assign n_4002 = n_4000 & n_4001;
assign n_4003 = n_4002 ^ x71;
assign n_4004 = n_4003 ^ x72;
assign n_4005 = n_3941 ^ n_4003;
assign n_4006 = n_4004 & n_4005;
assign n_4007 = n_4006 ^ x72;
assign n_4008 = n_4007 ^ x73;
assign n_4009 = n_3942 ^ n_4007;
assign n_4010 = n_4008 & n_4009;
assign n_4011 = n_4010 ^ x73;
assign n_4012 = n_4011 ^ x74;
assign n_4013 = n_3943 ^ n_4011;
assign n_4014 = n_4012 & n_4013;
assign n_4015 = n_4014 ^ x74;
assign n_4016 = n_4015 ^ x75;
assign n_4017 = n_3944 ^ n_4015;
assign n_4018 = n_4016 & n_4017;
assign n_4019 = n_4018 ^ x75;
assign n_4020 = n_4019 ^ x76;
assign n_4021 = n_3945 ^ n_4019;
assign n_4022 = n_4020 & n_4021;
assign n_4023 = n_4022 ^ x76;
assign n_4024 = n_4023 ^ x77;
assign n_4025 = n_3946 ^ n_4023;
assign n_4026 = n_4024 & n_4025;
assign n_4027 = n_4026 ^ x77;
assign n_4028 = n_4027 ^ x78;
assign n_4029 = n_3947 ^ n_4027;
assign n_4030 = n_4028 & n_4029;
assign n_4031 = n_4030 ^ x78;
assign n_4032 = n_4031 ^ x79;
assign n_4033 = n_3948 ^ n_4031;
assign n_4034 = n_4032 & n_4033;
assign n_4035 = n_4034 ^ x79;
assign n_4036 = n_4035 ^ x80;
assign n_4037 = n_3949 ^ n_4035;
assign n_4038 = n_4036 & n_4037;
assign n_4039 = n_4038 ^ x80;
assign n_4040 = n_4039 ^ x81;
assign n_4041 = n_3965 ^ n_4039;
assign n_4042 = n_4040 & n_4041;
assign n_4043 = n_4042 ^ x81;
assign n_4044 = n_4043 ^ x82;
assign n_4045 = n_3950 ^ n_4043;
assign n_4046 = n_4044 & n_4045;
assign n_4047 = n_4046 ^ x82;
assign n_4048 = n_4047 ^ x83;
assign n_4049 = n_3951 ^ n_4047;
assign n_4050 = n_4048 & n_4049;
assign n_4051 = n_4050 ^ x83;
assign n_4052 = n_4051 ^ x84;
assign n_4053 = n_3952 ^ n_4051;
assign n_4054 = n_4052 & n_4053;
assign n_4055 = n_4054 ^ x84;
assign n_4056 = n_4055 ^ x85;
assign n_4057 = n_3953 ^ n_4055;
assign n_4058 = n_4056 & n_4057;
assign n_4059 = n_4058 ^ x85;
assign n_4060 = n_4059 ^ x86;
assign n_4061 = n_3954 ^ n_4059;
assign n_4062 = n_4060 & n_4061;
assign n_4063 = n_4062 ^ x86;
assign n_4064 = n_4063 ^ x87;
assign n_4065 = n_3955 ^ n_4063;
assign n_4066 = n_4064 & n_4065;
assign n_4067 = n_4066 ^ x87;
assign n_4068 = n_4067 ^ x88;
assign n_4069 = n_3956 ^ n_4067;
assign n_4070 = n_4068 & n_4069;
assign n_4071 = n_4070 ^ x88;
assign n_4072 = n_4071 ^ x89;
assign n_4073 = n_3957 ^ n_4071;
assign n_4074 = n_4072 & n_4073;
assign n_4075 = n_4074 ^ x89;
assign n_4076 = n_4075 ^ x90;
assign n_4077 = n_3958 ^ n_4075;
assign n_4078 = n_4076 & n_4077;
assign n_4079 = n_4078 ^ x90;
assign n_4080 = n_4079 ^ x91;
assign n_4081 = n_3959 ^ n_4079;
assign n_4082 = n_4080 & n_4081;
assign n_4083 = n_4082 ^ x91;
assign n_4084 = n_4083 ^ x92;
assign n_4085 = n_3960 ^ n_4083;
assign n_4086 = n_4084 & n_4085;
assign n_4087 = n_4086 ^ x92;
assign n_4088 = n_4087 ^ x93;
assign n_4089 = n_3961 ^ n_4087;
assign n_4090 = n_4088 & n_4089;
assign n_4091 = n_4090 ^ x93;
assign n_4092 = n_4091 ^ x94;
assign n_4093 = n_3962 ^ n_4091;
assign n_4094 = n_4092 & n_4093;
assign n_4095 = n_4094 ^ x94;
assign n_4096 = n_4095 ^ x95;
assign n_4097 = n_3963 ^ n_4095;
assign n_4098 = n_4096 & n_4097;
assign n_4099 = n_4098 ^ x95;
assign n_4100 = n_4099 ^ x96;
assign n_4101 = n_3964 ^ n_4099;
assign n_4102 = n_4100 & ~n_4101;
assign n_4103 = n_4102 ^ n_4099;
assign n_4104 = n_4103 & n_3968;
assign n_4105 = ~n_439 ^ ~n_4104;
assign n_4106 = n_3756 & ~n_4104;
assign n_4107 = n_3967 & n_4105;
assign n_4108 = n_3988 & n_4106;
assign n_4109 = n_3984 & n_4106;
assign n_4110 = x30 ^ n_4106;
assign n_4111 = n_3981 & n_4106;
assign n_4112 = n_3992 & n_4106;
assign n_4113 = n_3996 & n_4106;
assign n_4114 = n_4000 & n_4106;
assign n_4115 = n_4004 & n_4106;
assign n_4116 = n_4008 & n_4106;
assign n_4117 = n_4012 & n_4106;
assign n_4118 = n_4016 & n_4106;
assign n_4119 = n_4020 & n_4106;
assign n_4120 = n_4024 & n_4106;
assign n_4121 = n_4028 & n_4106;
assign n_4122 = n_4032 & n_4106;
assign n_4123 = n_4036 & n_4106;
assign n_4124 = n_4040 & n_4106;
assign n_4125 = n_4044 & n_4106;
assign n_4126 = n_4048 & n_4106;
assign n_4127 = n_4052 & n_4106;
assign n_4128 = n_4056 & n_4106;
assign n_4129 = n_4060 & n_4106;
assign n_4130 = n_4064 & n_4106;
assign n_4131 = n_4068 & n_4106;
assign n_4132 = n_4072 & n_4106;
assign n_4133 = n_4076 & n_4106;
assign n_4134 = n_4080 & n_4106;
assign n_4135 = n_4084 & n_4106;
assign n_4136 = n_4088 & n_4106;
assign n_4137 = n_4092 & n_4106;
assign n_4138 = n_4096 & n_4106;
assign n_4139 = n_4100 & n_4106;
assign n_4140 = x64 & n_4106;
assign n_4141 = n_3894 & ~n_4106;
assign y30 = n_4106;
assign n_4142 = n_3972 & n_4106;
assign n_4143 = n_4108 ^ n_3937;
assign n_4144 = n_4109 ^ n_3936;
assign n_4145 = ~n_78 & n_4110;
assign n_4146 = n_4111 ^ n_3977;
assign n_4147 = n_4112 ^ n_3938;
assign n_4148 = n_4113 ^ n_3939;
assign n_4149 = n_4114 ^ n_3940;
assign n_4150 = n_4115 ^ n_3941;
assign n_4151 = n_4116 ^ n_3942;
assign n_4152 = n_4117 ^ n_3943;
assign n_4153 = n_4118 ^ n_3944;
assign n_4154 = n_4119 ^ n_3945;
assign n_4155 = n_4120 ^ n_3946;
assign n_4156 = n_4121 ^ n_3947;
assign n_4157 = n_4122 ^ n_3948;
assign n_4158 = n_4123 ^ n_3949;
assign n_4159 = n_4124 ^ n_3965;
assign n_4160 = n_4125 ^ n_3950;
assign n_4161 = n_4126 ^ n_3951;
assign n_4162 = n_4127 ^ n_3952;
assign n_4163 = n_4128 ^ n_3953;
assign n_4164 = n_4129 ^ n_3954;
assign n_4165 = n_4130 ^ n_3955;
assign n_4166 = n_4131 ^ n_3956;
assign n_4167 = n_4132 ^ n_3957;
assign n_4168 = n_4133 ^ n_3958;
assign n_4169 = n_4134 ^ n_3959;
assign n_4170 = n_4135 ^ n_3960;
assign n_4171 = n_4136 ^ n_3961;
assign n_4172 = n_4137 ^ n_3962;
assign n_4173 = n_4138 ^ n_3963;
assign n_4174 = n_4139 ^ n_3964;
assign n_4175 = n_3933 ^ n_4142;
assign n_4176 = n_4143 ^ x69;
assign n_4177 = n_4144 ^ x68;
assign n_4178 = n_4145 ^ n_210;
assign n_4179 = x64 & ~n_4178;
assign n_4180 = n_77 ^ n_4179;
assign n_4181 = n_4180 ^ x66;
assign n_4182 = n_4175 ^ n_4180;
assign n_4183 = n_4181 & n_4182;
assign n_4184 = n_4183 ^ x66;
assign n_4185 = n_4184 ^ x67;
assign n_4186 = n_4146 ^ n_4184;
assign n_4187 = n_4185 & ~n_4186;
assign n_4188 = n_4187 ^ x67;
assign n_4189 = n_4188 ^ n_4144;
assign n_4190 = n_4188 ^ x68;
assign n_4191 = ~n_4177 & n_4189;
assign n_4192 = n_4191 ^ x68;
assign n_4193 = n_4192 ^ n_4143;
assign n_4194 = n_4192 ^ x69;
assign n_4195 = ~n_4176 & n_4193;
assign n_4196 = n_4195 ^ x69;
assign n_4197 = n_4196 ^ x70;
assign n_4198 = n_4147 ^ n_4196;
assign n_4199 = n_4197 & n_4198;
assign n_4200 = n_4199 ^ x70;
assign n_4201 = n_4200 ^ x71;
assign n_4202 = n_4148 ^ n_4200;
assign n_4203 = n_4201 & n_4202;
assign n_4204 = n_4203 ^ x71;
assign n_4205 = n_4204 ^ x72;
assign n_4206 = n_4149 ^ n_4204;
assign n_4207 = n_4205 & n_4206;
assign n_4208 = n_4207 ^ x72;
assign n_4209 = n_4208 ^ x73;
assign n_4210 = n_4150 ^ n_4208;
assign n_4211 = n_4209 & n_4210;
assign n_4212 = n_4211 ^ x73;
assign n_4213 = n_4212 ^ x74;
assign n_4214 = n_4151 ^ n_4212;
assign n_4215 = n_4213 & n_4214;
assign n_4216 = n_4215 ^ x74;
assign n_4217 = n_4216 ^ x75;
assign n_4218 = n_4152 ^ n_4216;
assign n_4219 = n_4217 & n_4218;
assign n_4220 = n_4219 ^ x75;
assign n_4221 = n_4220 ^ x76;
assign n_4222 = n_4153 ^ n_4220;
assign n_4223 = n_4221 & n_4222;
assign n_4224 = n_4223 ^ x76;
assign n_4225 = n_4224 ^ x77;
assign n_4226 = n_4154 ^ n_4224;
assign n_4227 = n_4225 & n_4226;
assign n_4228 = n_4227 ^ x77;
assign n_4229 = n_4228 ^ x78;
assign n_4230 = n_4155 ^ n_4228;
assign n_4231 = n_4229 & n_4230;
assign n_4232 = n_4231 ^ x78;
assign n_4233 = n_4232 ^ x79;
assign n_4234 = n_4156 ^ n_4232;
assign n_4235 = n_4233 & n_4234;
assign n_4236 = n_4235 ^ x79;
assign n_4237 = n_4236 ^ x80;
assign n_4238 = n_4157 ^ n_4236;
assign n_4239 = n_4237 & n_4238;
assign n_4240 = n_4239 ^ x80;
assign n_4241 = n_4240 ^ x81;
assign n_4242 = n_4158 ^ n_4240;
assign n_4243 = n_4241 & n_4242;
assign n_4244 = n_4243 ^ x81;
assign n_4245 = n_4244 ^ x82;
assign n_4246 = n_4159 ^ n_4244;
assign n_4247 = n_4245 & n_4246;
assign n_4248 = n_4247 ^ x82;
assign n_4249 = n_4248 ^ x83;
assign n_4250 = n_4160 ^ n_4248;
assign n_4251 = n_4249 & n_4250;
assign n_4252 = n_4251 ^ x83;
assign n_4253 = n_4252 ^ x84;
assign n_4254 = n_4161 ^ n_4252;
assign n_4255 = n_4253 & n_4254;
assign n_4256 = n_4255 ^ x84;
assign n_4257 = n_4256 ^ x85;
assign n_4258 = n_4162 ^ n_4256;
assign n_4259 = n_4257 & n_4258;
assign n_4260 = n_4259 ^ x85;
assign n_4261 = n_4260 ^ x86;
assign n_4262 = n_4163 ^ n_4260;
assign n_4263 = n_4261 & n_4262;
assign n_4264 = n_4263 ^ x86;
assign n_4265 = n_4264 ^ x87;
assign n_4266 = n_4164 ^ n_4264;
assign n_4267 = n_4265 & n_4266;
assign n_4268 = n_4267 ^ x87;
assign n_4269 = n_4268 ^ x88;
assign n_4270 = n_4165 ^ n_4268;
assign n_4271 = n_4269 & n_4270;
assign n_4272 = n_4271 ^ x88;
assign n_4273 = n_4272 ^ x89;
assign n_4274 = n_4166 ^ n_4272;
assign n_4275 = n_4273 & n_4274;
assign n_4276 = n_4275 ^ x89;
assign n_4277 = n_4276 ^ x90;
assign n_4278 = n_4167 ^ n_4276;
assign n_4279 = n_4277 & n_4278;
assign n_4280 = n_4279 ^ x90;
assign n_4281 = n_4280 ^ x91;
assign n_4282 = n_4168 ^ n_4280;
assign n_4283 = n_4281 & n_4282;
assign n_4284 = n_4283 ^ x91;
assign n_4285 = n_4284 ^ x92;
assign n_4286 = n_4169 ^ n_4284;
assign n_4287 = n_4285 & n_4286;
assign n_4288 = n_4287 ^ x92;
assign n_4289 = n_4288 ^ x93;
assign n_4290 = n_4170 ^ n_4288;
assign n_4291 = n_4289 & n_4290;
assign n_4292 = n_4291 ^ x93;
assign n_4293 = n_4292 ^ x94;
assign n_4294 = n_4171 ^ n_4292;
assign n_4295 = n_4293 & n_4294;
assign n_4296 = n_4295 ^ x94;
assign n_4297 = n_4296 ^ x95;
assign n_4298 = n_4172 ^ n_4296;
assign n_4299 = n_4297 & n_4298;
assign n_4300 = n_4299 ^ x95;
assign n_4301 = n_4300 ^ x96;
assign n_4302 = n_4173 ^ n_4300;
assign n_4303 = n_4301 & n_4302;
assign n_4304 = n_4303 ^ x96;
assign n_4305 = n_4304 ^ x97;
assign n_4306 = n_4174 ^ n_4304;
assign n_4307 = n_4305 & ~n_4306;
assign n_4308 = n_4307 ^ n_4304;
assign n_4309 = ~n_4107 & n_4308;
assign n_4310 = n_3976 & ~n_4309;
assign n_4311 = n_4194 & n_4310;
assign n_4312 = n_4190 & n_4310;
assign n_4313 = x28 ^ n_4310;
assign n_4314 = x64 & n_4310;
assign n_4315 = x65 & n_4310;
assign n_4316 = n_4181 & n_4310;
assign n_4317 = n_4185 & n_4310;
assign n_4318 = n_4197 & n_4310;
assign n_4319 = n_4201 & n_4310;
assign n_4320 = n_4205 & n_4310;
assign n_4321 = n_4209 & n_4310;
assign n_4322 = n_4213 & n_4310;
assign n_4323 = n_4217 & n_4310;
assign n_4324 = n_4221 & n_4310;
assign n_4325 = n_4225 & n_4310;
assign n_4326 = n_4229 & n_4310;
assign n_4327 = n_4233 & n_4310;
assign n_4328 = n_4237 & n_4310;
assign n_4329 = n_4241 & n_4310;
assign n_4330 = n_4245 & n_4310;
assign n_4331 = n_4249 & n_4310;
assign n_4332 = n_4253 & n_4310;
assign n_4333 = n_4257 & n_4310;
assign n_4334 = n_4261 & n_4310;
assign n_4335 = n_4265 & n_4310;
assign n_4336 = n_4269 & n_4310;
assign n_4337 = n_4273 & n_4310;
assign n_4338 = n_4277 & n_4310;
assign n_4339 = n_4305 & n_4310;
assign n_4340 = n_4301 & n_4310;
assign n_4341 = n_4289 & n_4310;
assign n_4342 = n_4285 & n_4310;
assign n_4343 = n_4281 & n_4310;
assign n_4344 = n_4293 & n_4310;
assign n_4345 = n_4297 & n_4310;
assign y29 = n_4310;
assign n_4346 = n_4141 & ~n_4310;
assign n_4347 = n_4311 ^ n_4143;
assign n_4348 = n_4312 ^ n_4144;
assign n_4349 = n_209 & ~n_4313;
assign n_4350 = ~x29 & n_4314;
assign n_4351 = n_4316 ^ n_4175;
assign n_4352 = n_4317 ^ n_4146;
assign n_4353 = n_4318 ^ n_4147;
assign n_4354 = n_4319 ^ n_4148;
assign n_4355 = n_4320 ^ n_4149;
assign n_4356 = n_4321 ^ n_4150;
assign n_4357 = n_4322 ^ n_4151;
assign n_4358 = n_4323 ^ n_4152;
assign n_4359 = n_4324 ^ n_4153;
assign n_4360 = n_4325 ^ n_4154;
assign n_4361 = n_4326 ^ n_4155;
assign n_4362 = n_4327 ^ n_4156;
assign n_4363 = n_4328 ^ n_4157;
assign n_4364 = n_4329 ^ n_4158;
assign n_4365 = n_4330 ^ n_4159;
assign n_4366 = n_4331 ^ n_4160;
assign n_4367 = n_4332 ^ n_4161;
assign n_4368 = n_4333 ^ n_4162;
assign n_4369 = n_4334 ^ n_4163;
assign n_4370 = n_4335 ^ n_4164;
assign n_4371 = n_4336 ^ n_4165;
assign n_4372 = n_4337 ^ n_4166;
assign n_4373 = n_4338 ^ n_4167;
assign n_4374 = n_4339 ^ n_4174;
assign n_4375 = n_4340 ^ n_4173;
assign n_4376 = n_4341 ^ n_4170;
assign n_4377 = n_4342 ^ n_4169;
assign n_4378 = n_4343 ^ n_4168;
assign n_4379 = n_4344 ^ n_4171;
assign n_4380 = n_4345 ^ n_4172;
assign n_4381 = ~n_439 ^ ~n_4346;
assign n_4382 = ~x70 ^ n_4347;
assign n_4383 = n_4347 ^ x70;
assign n_4384 = n_4348 ^ x69;
assign n_4385 = x69 & ~n_4348;
assign n_4386 = n_4349 ^ x28;
assign n_4387 = n_4350 ^ n_79;
assign n_4388 = n_4140 ^ n_4350;
assign n_4389 = ~x98 ^ n_4374;
assign n_4390 = n_4374 ^ x98;
assign n_4391 = n_4375 ^ x97;
assign n_4392 = x97 & ~n_4375;
assign n_4393 = ~x94 ^ n_4376;
assign n_4394 = n_4376 ^ x94;
assign n_4395 = n_4377 ^ x93;
assign n_4396 = x93 & ~n_4377;
assign n_4397 = n_4384 ^ n_4385;
assign n_4398 = n_4385 ^ n_4347;
assign n_4399 = x64 & ~n_4386;
assign n_4400 = n_4315 ^ n_4388;
assign n_4401 = n_4391 ^ n_4392;
assign n_4402 = n_4392 ^ n_4374;
assign n_4403 = n_4395 ^ n_4396;
assign n_4404 = n_4396 ^ n_4376;
assign n_4405 = n_4382 & ~n_4397;
assign n_4406 = ~n_4383 & n_4398;
assign n_4407 = n_78 ^ n_4399;
assign n_4408 = n_4400 ^ x30;
assign n_4409 = n_4389 & ~n_4401;
assign n_4410 = ~n_4390 & n_4402;
assign n_4411 = n_4393 & ~n_4403;
assign n_4412 = ~n_4394 & n_4404;
assign n_4413 = n_4406 ^ x70;
assign n_4414 = n_4407 ^ n_4387;
assign n_4415 = n_4410 ^ x98;
assign n_4416 = n_4412 ^ x94;
assign n_4417 = n_4414 ^ x66;
assign n_4418 = n_4408 ^ n_4414;
assign n_4419 = n_4417 & n_4418;
assign n_4420 = n_4419 ^ x66;
assign n_4421 = n_4420 ^ x67;
assign n_4422 = n_4351 ^ n_4420;
assign n_4423 = n_4421 & n_4422;
assign n_4424 = n_4423 ^ x67;
assign n_4425 = n_4424 ^ x68;
assign n_4426 = n_4352 ^ n_4424;
assign n_4427 = n_4425 & ~n_4426;
assign n_4428 = n_4427 ^ x68;
assign n_4429 = n_4428 ^ x69;
assign n_4430 = n_4428 ^ n_4348;
assign n_4431 = n_4405 & n_4428;
assign n_4432 = n_4429 & n_4430;
assign n_4433 = ~n_4413 & ~n_4431;
assign n_4434 = n_4432 ^ x69;
assign n_4435 = x71 ^ n_4433;
assign n_4436 = n_4353 ^ n_4433;
assign n_4437 = n_4434 ^ x70;
assign n_4438 = ~n_4435 & ~n_4436;
assign n_4439 = n_4438 ^ x71;
assign n_4440 = n_4439 ^ x72;
assign n_4441 = n_4354 ^ n_4439;
assign n_4442 = n_4440 & n_4441;
assign n_4443 = n_4442 ^ x72;
assign n_4444 = n_4443 ^ x73;
assign n_4445 = n_4355 ^ n_4443;
assign n_4446 = n_4444 & n_4445;
assign n_4447 = n_4446 ^ x73;
assign n_4448 = n_4447 ^ x74;
assign n_4449 = n_4356 ^ n_4447;
assign n_4450 = n_4448 & n_4449;
assign n_4451 = n_4450 ^ x74;
assign n_4452 = n_4451 ^ x75;
assign n_4453 = n_4357 ^ n_4451;
assign n_4454 = n_4452 & n_4453;
assign n_4455 = n_4454 ^ x75;
assign n_4456 = n_4455 ^ x76;
assign n_4457 = n_4358 ^ n_4455;
assign n_4458 = n_4456 & n_4457;
assign n_4459 = n_4458 ^ x76;
assign n_4460 = n_4459 ^ x77;
assign n_4461 = n_4359 ^ n_4459;
assign n_4462 = n_4460 & n_4461;
assign n_4463 = n_4462 ^ x77;
assign n_4464 = n_4463 ^ x78;
assign n_4465 = n_4360 ^ n_4463;
assign n_4466 = n_4464 & n_4465;
assign n_4467 = n_4466 ^ x78;
assign n_4468 = n_4467 ^ x79;
assign n_4469 = n_4361 ^ n_4467;
assign n_4470 = n_4468 & n_4469;
assign n_4471 = n_4470 ^ x79;
assign n_4472 = n_4471 ^ x80;
assign n_4473 = n_4362 ^ n_4471;
assign n_4474 = n_4472 & n_4473;
assign n_4475 = n_4474 ^ x80;
assign n_4476 = n_4475 ^ x81;
assign n_4477 = n_4363 ^ n_4475;
assign n_4478 = n_4476 & n_4477;
assign n_4479 = n_4478 ^ x81;
assign n_4480 = n_4479 ^ x82;
assign n_4481 = n_4364 ^ n_4479;
assign n_4482 = n_4480 & n_4481;
assign n_4483 = n_4482 ^ x82;
assign n_4484 = n_4483 ^ x83;
assign n_4485 = n_4365 ^ n_4483;
assign n_4486 = n_4484 & n_4485;
assign n_4487 = n_4486 ^ x83;
assign n_4488 = n_4487 ^ x84;
assign n_4489 = n_4366 ^ n_4487;
assign n_4490 = n_4488 & n_4489;
assign n_4491 = n_4490 ^ x84;
assign n_4492 = n_4491 ^ x85;
assign n_4493 = n_4367 ^ n_4491;
assign n_4494 = n_4492 & n_4493;
assign n_4495 = n_4494 ^ x85;
assign n_4496 = n_4495 ^ x86;
assign n_4497 = n_4368 ^ n_4495;
assign n_4498 = n_4496 & n_4497;
assign n_4499 = n_4498 ^ x86;
assign n_4500 = n_4499 ^ x87;
assign n_4501 = n_4369 ^ n_4499;
assign n_4502 = n_4500 & n_4501;
assign n_4503 = n_4502 ^ x87;
assign n_4504 = n_4503 ^ x88;
assign n_4505 = n_4370 ^ n_4503;
assign n_4506 = n_4504 & n_4505;
assign n_4507 = n_4506 ^ x88;
assign n_4508 = n_4507 ^ x89;
assign n_4509 = n_4371 ^ n_4507;
assign n_4510 = n_4508 & n_4509;
assign n_4511 = n_4510 ^ x89;
assign n_4512 = n_4511 ^ x90;
assign n_4513 = n_4372 ^ n_4511;
assign n_4514 = n_4512 & n_4513;
assign n_4515 = n_4514 ^ x90;
assign n_4516 = n_4515 ^ x91;
assign n_4517 = n_4373 ^ n_4515;
assign n_4518 = n_4516 & n_4517;
assign n_4519 = n_4518 ^ x91;
assign n_4520 = n_4519 ^ x92;
assign n_4521 = n_4378 ^ n_4519;
assign n_4522 = n_4520 & n_4521;
assign n_4523 = n_4522 ^ x92;
assign n_4524 = n_4523 ^ x93;
assign n_4525 = n_4523 ^ n_4377;
assign n_4526 = n_4411 & n_4523;
assign n_4527 = n_4524 & n_4525;
assign n_4528 = ~n_4416 & ~n_4526;
assign n_4529 = n_4527 ^ x93;
assign n_4530 = x95 ^ n_4528;
assign n_4531 = n_4379 ^ n_4528;
assign n_4532 = n_4529 ^ x94;
assign n_4533 = ~n_4530 & ~n_4531;
assign n_4534 = n_4533 ^ x95;
assign n_4535 = n_4534 ^ x96;
assign n_4536 = n_4380 ^ n_4534;
assign n_4537 = n_4535 & n_4536;
assign n_4538 = n_4537 ^ x96;
assign n_4539 = n_4538 ^ x97;
assign n_4540 = n_4538 ^ n_4375;
assign n_4541 = n_4409 & n_4538;
assign n_4542 = n_4539 & n_4540;
assign n_4543 = ~n_4415 & ~n_4541;
assign n_4544 = n_4542 ^ x97;
assign n_4545 = x99 ^ n_4543;
assign n_4546 = ~n_4381 ^ n_4543;
assign n_4547 = n_4544 ^ x98;
assign n_4548 = ~n_4545 & ~n_4546;
assign n_4549 = n_4548 ^ n_4543;
assign n_4550 = n_370 & n_4549;
assign n_4551 = n_4520 & n_4550;
assign n_4552 = n_4516 & n_4550;
assign n_4553 = n_4500 & n_4550;
assign n_4554 = n_4496 & n_4550;
assign n_4555 = n_4476 & n_4550;
assign n_4556 = n_4472 & n_4550;
assign n_4557 = n_4460 & n_4550;
assign n_4558 = n_4456 & n_4550;
assign n_4559 = x65 & n_4550;
assign n_4560 = x64 & n_4550;
assign n_4561 = x65 ^ n_4550;
assign n_4562 = n_4417 & n_4550;
assign n_4563 = n_4421 & n_4550;
assign n_4564 = n_4425 & n_4550;
assign n_4565 = n_4429 & n_4550;
assign n_4566 = ~n_4435 & n_4550;
assign n_4567 = n_4440 & n_4550;
assign n_4568 = n_4444 & n_4550;
assign n_4569 = n_4448 & n_4550;
assign n_4570 = n_4452 & n_4550;
assign n_4571 = n_4464 & n_4550;
assign n_4572 = n_4468 & n_4550;
assign n_4573 = n_4484 & n_4550;
assign n_4574 = n_4480 & n_4550;
assign n_4575 = n_4488 & n_4550;
assign n_4576 = n_4492 & n_4550;
assign n_4577 = n_4504 & n_4550;
assign n_4578 = n_4508 & n_4550;
assign n_4579 = n_4512 & n_4550;
assign n_4580 = n_4524 & n_4550;
assign n_4581 = ~n_4530 & n_4550;
assign n_4582 = n_4535 & n_4550;
assign n_4583 = n_4539 & n_4550;
assign n_4584 = n_4381 & ~n_4550;
assign y28 = n_4550;
assign n_4585 = n_4437 & n_4550;
assign n_4586 = n_4532 & n_4550;
assign n_4587 = n_4547 & n_4550;
assign n_4588 = n_4551 ^ n_4378;
assign n_4589 = n_4552 ^ n_4373;
assign n_4590 = n_4553 ^ n_4369;
assign n_4591 = n_4554 ^ n_4368;
assign n_4592 = n_4555 ^ n_4363;
assign n_4593 = n_4556 ^ n_4362;
assign n_4594 = n_4557 ^ n_4359;
assign n_4595 = n_4558 ^ n_4358;
assign n_4596 = ~x28 & n_4560;
assign n_4597 = n_4560 ^ x28;
assign n_4598 = n_4561 ^ x28;
assign n_4599 = n_4562 ^ n_4408;
assign n_4600 = n_4563 ^ n_4351;
assign n_4601 = n_4564 ^ n_4352;
assign n_4602 = n_4565 ^ n_4348;
assign n_4603 = n_4566 ^ n_4353;
assign n_4604 = n_4567 ^ n_4354;
assign n_4605 = n_4568 ^ n_4355;
assign n_4606 = n_4569 ^ n_4356;
assign n_4607 = n_4570 ^ n_4357;
assign n_4608 = n_4571 ^ n_4360;
assign n_4609 = n_4572 ^ n_4361;
assign n_4610 = n_4573 ^ n_4365;
assign n_4611 = n_4574 ^ n_4364;
assign n_4612 = n_4575 ^ n_4366;
assign n_4613 = n_4576 ^ n_4367;
assign n_4614 = n_4577 ^ n_4370;
assign n_4615 = n_4578 ^ n_4371;
assign n_4616 = n_4579 ^ n_4372;
assign n_4617 = n_4580 ^ n_4377;
assign n_4618 = n_4581 ^ n_4379;
assign n_4619 = n_4582 ^ n_4380;
assign n_4620 = n_4583 ^ n_4375;
assign n_4621 = ~n_439 & ~n_4584;
assign n_4622 = n_4347 ^ n_4585;
assign n_4623 = n_4376 ^ n_4586;
assign n_4624 = n_4374 ^ n_4587;
assign n_4625 = ~x93 ^ n_4588;
assign n_4626 = n_4588 ^ x93;
assign n_4627 = n_4589 ^ x92;
assign n_4628 = x92 & ~n_4589;
assign n_4629 = ~x88 ^ n_4590;
assign n_4630 = n_4590 ^ x88;
assign n_4631 = n_4591 ^ x87;
assign n_4632 = x87 & ~n_4591;
assign n_4633 = ~x82 ^ n_4592;
assign n_4634 = n_4592 ^ x82;
assign n_4635 = n_4593 ^ x81;
assign n_4636 = x81 & ~n_4593;
assign n_4637 = n_4594 ^ x78;
assign n_4638 = n_4595 ^ x77;
assign n_4639 = n_4559 ^ n_4596;
assign n_4640 = x65 & ~n_4597;
assign n_4641 = x64 & ~n_4598;
assign n_4642 = ~x84 ^ n_4610;
assign n_4643 = n_4610 ^ x84;
assign n_4644 = n_4611 ^ x83;
assign n_4645 = x83 & ~n_4611;
assign n_4646 = n_4621 ^ x100;
assign n_4647 = n_4627 ^ n_4628;
assign n_4648 = n_4628 ^ n_4588;
assign n_4649 = n_4631 ^ n_4632;
assign n_4650 = n_4632 ^ n_4590;
assign n_4651 = n_4635 ^ n_4636;
assign n_4652 = n_4636 ^ n_4592;
assign n_4653 = n_4639 ^ n_4314;
assign n_4654 = ~x27 & n_4641;
assign n_4655 = n_4644 ^ n_4645;
assign n_4656 = n_4645 ^ n_4610;
assign n_4657 = n_4625 & ~n_4647;
assign n_4658 = ~n_4626 & n_4648;
assign n_4659 = n_4629 & ~n_4649;
assign n_4660 = ~n_4630 & n_4650;
assign n_4661 = n_4633 & ~n_4651;
assign n_4662 = ~n_4634 & n_4652;
assign n_4663 = n_4653 ^ x29;
assign n_4664 = n_4640 ^ n_4654;
assign n_4665 = n_4642 & ~n_4655;
assign n_4666 = ~n_4643 & n_4656;
assign n_4667 = n_4658 ^ x93;
assign n_4668 = n_4660 ^ x88;
assign n_4669 = n_4662 ^ x82;
assign n_4670 = n_4663 ^ x66;
assign n_4671 = n_4664 ^ n_4663;
assign n_4672 = n_4664 ^ x66;
assign n_4673 = n_4666 ^ x84;
assign n_4674 = ~n_4670 & n_4671;
assign n_4675 = n_4674 ^ x66;
assign n_4676 = n_4675 ^ x67;
assign n_4677 = n_4599 ^ n_4675;
assign n_4678 = n_4676 & n_4677;
assign n_4679 = n_4678 ^ x67;
assign n_4680 = n_4679 ^ x68;
assign n_4681 = n_4600 ^ n_4679;
assign n_4682 = n_4680 & n_4681;
assign n_4683 = n_4682 ^ x68;
assign n_4684 = n_4683 ^ x69;
assign n_4685 = n_4601 ^ n_4683;
assign n_4686 = n_4684 & ~n_4685;
assign n_4687 = n_4686 ^ x69;
assign n_4688 = n_4687 ^ x70;
assign n_4689 = n_4602 ^ n_4687;
assign n_4690 = n_4688 & n_4689;
assign n_4691 = n_4690 ^ x70;
assign n_4692 = n_4691 ^ x71;
assign n_4693 = n_4622 ^ n_4691;
assign n_4694 = n_4692 & n_4693;
assign n_4695 = n_4694 ^ x71;
assign n_4696 = n_4695 ^ x72;
assign n_4697 = n_4603 ^ n_4695;
assign n_4698 = n_4696 & n_4697;
assign n_4699 = n_4698 ^ x72;
assign n_4700 = n_4699 ^ x73;
assign n_4701 = n_4604 ^ n_4699;
assign n_4702 = n_4700 & n_4701;
assign n_4703 = n_4702 ^ x73;
assign n_4704 = n_4703 ^ x74;
assign n_4705 = n_4605 ^ n_4703;
assign n_4706 = n_4704 & n_4705;
assign n_4707 = n_4706 ^ x74;
assign n_4708 = n_4707 ^ x75;
assign n_4709 = n_4606 ^ n_4707;
assign n_4710 = n_4708 & n_4709;
assign n_4711 = n_4710 ^ x75;
assign n_4712 = n_4711 ^ x76;
assign n_4713 = n_4607 ^ n_4711;
assign n_4714 = n_4712 & n_4713;
assign n_4715 = n_4714 ^ x76;
assign n_4716 = n_4715 ^ n_4595;
assign n_4717 = n_4715 ^ x77;
assign n_4718 = ~n_4638 & n_4716;
assign n_4719 = n_4718 ^ x77;
assign n_4720 = n_4719 ^ n_4594;
assign n_4721 = n_4719 ^ x78;
assign n_4722 = ~n_4637 & n_4720;
assign n_4723 = n_4722 ^ x78;
assign n_4724 = n_4723 ^ x79;
assign n_4725 = n_4608 ^ n_4723;
assign n_4726 = n_4724 & n_4725;
assign n_4727 = n_4726 ^ x79;
assign n_4728 = n_4727 ^ x80;
assign n_4729 = n_4609 ^ n_4727;
assign n_4730 = n_4728 & n_4729;
assign n_4731 = n_4730 ^ x80;
assign n_4732 = n_4731 ^ x81;
assign n_4733 = n_4731 ^ n_4593;
assign n_4734 = n_4661 & n_4731;
assign n_4735 = n_4732 & n_4733;
assign n_4736 = ~n_4669 & ~n_4734;
assign n_4737 = n_4735 ^ x81;
assign n_4738 = x83 ^ n_4736;
assign n_4739 = n_4611 ^ n_4736;
assign n_4740 = n_4665 & ~n_4736;
assign n_4741 = n_4737 ^ x82;
assign n_4742 = ~n_4738 & ~n_4739;
assign n_4743 = ~n_4673 & ~n_4740;
assign n_4744 = n_4742 ^ x83;
assign n_4745 = x85 ^ n_4743;
assign n_4746 = n_4612 ^ n_4743;
assign n_4747 = n_4744 ^ x84;
assign n_4748 = ~n_4745 & ~n_4746;
assign n_4749 = n_4748 ^ x85;
assign n_4750 = n_4749 ^ x86;
assign n_4751 = n_4613 ^ n_4749;
assign n_4752 = n_4750 & n_4751;
assign n_4753 = n_4752 ^ x86;
assign n_4754 = n_4753 ^ x87;
assign n_4755 = n_4753 ^ n_4591;
assign n_4756 = n_4659 & n_4753;
assign n_4757 = n_4754 & n_4755;
assign n_4758 = ~n_4668 & ~n_4756;
assign n_4759 = n_4757 ^ x87;
assign n_4760 = x89 ^ n_4758;
assign n_4761 = n_4614 ^ n_4758;
assign n_4762 = n_4759 ^ x88;
assign n_4763 = ~n_4760 & ~n_4761;
assign n_4764 = n_4763 ^ x89;
assign n_4765 = n_4764 ^ x90;
assign n_4766 = n_4615 ^ n_4764;
assign n_4767 = n_4765 & n_4766;
assign n_4768 = n_4767 ^ x90;
assign n_4769 = n_4768 ^ x91;
assign n_4770 = n_4616 ^ n_4768;
assign n_4771 = n_4769 & n_4770;
assign n_4772 = n_4771 ^ x91;
assign n_4773 = n_4772 ^ x92;
assign n_4774 = n_4772 ^ n_4589;
assign n_4775 = n_4657 & n_4772;
assign n_4776 = n_4773 & n_4774;
assign n_4777 = ~n_4667 & ~n_4775;
assign n_4778 = n_4776 ^ x92;
assign n_4779 = x94 ^ n_4777;
assign n_4780 = n_4617 ^ n_4777;
assign n_4781 = n_4778 ^ x93;
assign n_4782 = ~n_4779 & ~n_4780;
assign n_4783 = n_4782 ^ x94;
assign n_4784 = n_4783 ^ x95;
assign n_4785 = n_4623 ^ n_4783;
assign n_4786 = n_4784 & n_4785;
assign n_4787 = n_4786 ^ x95;
assign n_4788 = n_4787 ^ x96;
assign n_4789 = n_4618 ^ n_4787;
assign n_4790 = n_4788 & n_4789;
assign n_4791 = n_4790 ^ x96;
assign n_4792 = n_4791 ^ x97;
assign n_4793 = n_4619 ^ n_4791;
assign n_4794 = n_4792 & n_4793;
assign n_4795 = n_4794 ^ x97;
assign n_4796 = n_4795 ^ x98;
assign n_4797 = n_4620 ^ n_4795;
assign n_4798 = n_4796 & n_4797;
assign n_4799 = n_4798 ^ x98;
assign n_4800 = n_4799 ^ x99;
assign n_4801 = n_4624 ^ n_4799;
assign n_4802 = n_4800 & ~n_4801;
assign n_4803 = n_4802 ^ n_4799;
assign n_4804 = n_4803 ^ x100;
assign n_4805 = n_4646 & n_4804;
assign n_4806 = x100 ^ n_4805;
assign n_4807 = n_369 & ~n_4806;
assign n_4808 = n_4800 & n_4807;
assign n_4809 = n_4584 & ~n_4807;
assign n_4810 = n_4788 & n_4807;
assign n_4811 = n_4784 & n_4807;
assign n_4812 = n_4773 & n_4807;
assign n_4813 = ~n_4760 & n_4807;
assign n_4814 = n_4717 & n_4807;
assign n_4815 = n_4712 & n_4807;
assign n_4816 = n_20 & n_4807;
assign n_4817 = x65 & n_4807;
assign n_4818 = x64 & n_4807;
assign n_4819 = n_4672 & n_4807;
assign n_4820 = n_4676 & n_4807;
assign n_4821 = n_4680 & n_4807;
assign n_4822 = n_4684 & n_4807;
assign n_4823 = n_4688 & n_4807;
assign n_4824 = n_4692 & n_4807;
assign n_4825 = n_4696 & n_4807;
assign n_4826 = n_4700 & n_4807;
assign n_4827 = n_4704 & n_4807;
assign n_4828 = n_4708 & n_4807;
assign n_4829 = n_4721 & n_4807;
assign n_4830 = n_4724 & n_4807;
assign n_4831 = n_4728 & n_4807;
assign n_4832 = n_4732 & n_4807;
assign n_4833 = ~n_4738 & n_4807;
assign n_4834 = ~n_4745 & n_4807;
assign n_4835 = n_4750 & n_4807;
assign n_4836 = n_4754 & n_4807;
assign n_4837 = n_4765 & n_4807;
assign n_4838 = n_4769 & n_4807;
assign n_4839 = ~n_4779 & n_4807;
assign n_4840 = n_4792 & n_4807;
assign n_4841 = n_4796 & n_4807;
assign y27 = n_4807;
assign n_4842 = n_4781 & n_4807;
assign n_4843 = n_4762 & n_4807;
assign n_4844 = n_4741 & n_4807;
assign n_4845 = n_4747 & n_4807;
assign n_4846 = n_4808 ^ n_4624;
assign n_4847 = ~n_439 ^ ~n_4809;
assign n_4848 = ~n_368 & n_4809;
assign n_4849 = n_4810 ^ n_4618;
assign n_4850 = n_4811 ^ n_4623;
assign n_4851 = n_4812 ^ n_4589;
assign n_4852 = n_4813 ^ n_4614;
assign n_4853 = n_4814 ^ n_4595;
assign n_4854 = n_4815 ^ n_4607;
assign n_4855 = n_4816 ^ n_4560;
assign n_4856 = n_4817 ^ x28;
assign n_4857 = n_4818 ^ n_20;
assign n_4858 = n_4818 ^ x27;
assign n_4859 = n_4819 ^ n_4663;
assign n_4860 = n_4820 ^ n_4599;
assign n_4861 = n_4821 ^ n_4600;
assign n_4862 = n_4822 ^ n_4601;
assign n_4863 = n_4823 ^ n_4602;
assign n_4864 = n_4824 ^ n_4622;
assign n_4865 = n_4825 ^ n_4603;
assign n_4866 = n_4826 ^ n_4604;
assign n_4867 = n_4827 ^ n_4605;
assign n_4868 = n_4828 ^ n_4606;
assign n_4869 = n_4829 ^ n_4594;
assign n_4870 = n_4830 ^ n_4608;
assign n_4871 = n_4831 ^ n_4609;
assign n_4872 = n_4832 ^ n_4593;
assign n_4873 = n_4833 ^ n_4611;
assign n_4874 = n_4834 ^ n_4612;
assign n_4875 = n_4835 ^ n_4613;
assign n_4876 = n_4836 ^ n_4591;
assign n_4877 = n_4837 ^ n_4615;
assign n_4878 = n_4838 ^ n_4616;
assign n_4879 = n_4839 ^ n_4617;
assign n_4880 = n_4840 ^ n_4619;
assign n_4881 = n_4841 ^ n_4620;
assign n_4882 = n_4588 ^ n_4842;
assign n_4883 = n_4590 ^ n_4843;
assign n_4884 = n_4592 ^ n_4844;
assign n_4885 = n_4610 ^ n_4845;
assign n_4886 = ~n_4847 ^ x101;
assign n_4887 = x101 & ~n_4847;
assign n_4888 = x100 & ~n_4847;
assign n_4889 = n_4847 & n_363;
assign n_4890 = ~x97 ^ n_4849;
assign n_4891 = n_4849 ^ x97;
assign n_4892 = n_4850 ^ x96;
assign n_4893 = x96 & ~n_4850;
assign n_4894 = n_4851 ^ x93;
assign n_4895 = ~x90 ^ n_4852;
assign n_4896 = n_4852 ^ x90;
assign n_4897 = ~x78 ^ n_4853;
assign n_4898 = n_4853 ^ x78;
assign n_4899 = n_4854 ^ x77;
assign n_4900 = x77 & ~n_4854;
assign n_4901 = n_4855 ^ n_4856;
assign n_4902 = ~x26 & n_4857;
assign n_4903 = x65 & ~n_4858;
assign n_4904 = n_4882 ^ x94;
assign n_4905 = n_4883 ^ x89;
assign n_4906 = x89 & ~n_4883;
assign n_4907 = n_4886 ^ n_4887;
assign n_4908 = n_368 & ~n_4887;
assign n_4909 = ~n_366 & ~n_4889;
assign n_4910 = n_4892 ^ n_4893;
assign n_4911 = n_4893 ^ n_4849;
assign n_4912 = n_4899 ^ n_4900;
assign n_4913 = n_4900 ^ n_4853;
assign n_4914 = n_4901 ^ x66;
assign n_4915 = n_4902 ^ n_211;
assign n_4916 = n_4905 ^ n_4906;
assign n_4917 = n_4906 ^ n_4852;
assign n_4918 = ~n_4846 & n_4907;
assign n_4919 = n_4890 & ~n_4910;
assign n_4920 = ~n_4891 & n_4911;
assign n_4921 = n_4897 & ~n_4912;
assign n_4922 = ~n_4898 & n_4913;
assign n_4923 = n_4915 ^ n_4903;
assign n_4924 = n_4895 & ~n_4916;
assign n_4925 = ~n_4896 & n_4917;
assign n_4926 = ~n_4918 ^ ~n_125;
assign n_4927 = x100 & n_4918;
assign n_4928 = n_4920 ^ x97;
assign n_4929 = n_4922 ^ x78;
assign n_4930 = n_4923 ^ n_4901;
assign n_4931 = n_4923 ^ x66;
assign n_4932 = n_4925 ^ x90;
assign n_4933 = ~n_4927 & n_4908;
assign n_4934 = ~n_4914 & n_4930;
assign n_4935 = n_4934 ^ x66;
assign n_4936 = n_4935 ^ x67;
assign n_4937 = n_4859 ^ n_4935;
assign n_4938 = n_4936 & n_4937;
assign n_4939 = n_4938 ^ x67;
assign n_4940 = n_4939 ^ x68;
assign n_4941 = n_4860 ^ n_4939;
assign n_4942 = n_4940 & n_4941;
assign n_4943 = n_4942 ^ x68;
assign n_4944 = n_4943 ^ x69;
assign n_4945 = n_4861 ^ n_4943;
assign n_4946 = n_4944 & n_4945;
assign n_4947 = n_4946 ^ x69;
assign n_4948 = n_4947 ^ x70;
assign n_4949 = n_4862 ^ n_4947;
assign n_4950 = n_4948 & ~n_4949;
assign n_4951 = n_4950 ^ x70;
assign n_4952 = n_4951 ^ x71;
assign n_4953 = n_4863 ^ n_4951;
assign n_4954 = n_4952 & n_4953;
assign n_4955 = n_4954 ^ x71;
assign n_4956 = n_4955 ^ x72;
assign n_4957 = n_4864 ^ n_4955;
assign n_4958 = n_4956 & n_4957;
assign n_4959 = n_4958 ^ x72;
assign n_4960 = n_4959 ^ x73;
assign n_4961 = n_4865 ^ n_4959;
assign n_4962 = n_4960 & n_4961;
assign n_4963 = n_4962 ^ x73;
assign n_4964 = n_4963 ^ x74;
assign n_4965 = n_4866 ^ n_4963;
assign n_4966 = n_4964 & n_4965;
assign n_4967 = n_4966 ^ x74;
assign n_4968 = n_4967 ^ x75;
assign n_4969 = n_4867 ^ n_4967;
assign n_4970 = n_4968 & n_4969;
assign n_4971 = n_4970 ^ x75;
assign n_4972 = n_4971 ^ x76;
assign n_4973 = n_4868 ^ n_4971;
assign n_4974 = n_4972 & n_4973;
assign n_4975 = n_4974 ^ x76;
assign n_4976 = n_4975 ^ x77;
assign n_4977 = n_4975 ^ n_4854;
assign n_4978 = n_4921 & n_4975;
assign n_4979 = n_4976 & n_4977;
assign n_4980 = ~n_4929 & ~n_4978;
assign n_4981 = n_4979 ^ x77;
assign n_4982 = x79 ^ n_4980;
assign n_4983 = n_4869 ^ n_4980;
assign n_4984 = n_4981 ^ x78;
assign n_4985 = ~n_4982 & ~n_4983;
assign n_4986 = n_4985 ^ x79;
assign n_4987 = n_4986 ^ x80;
assign n_4988 = n_4870 ^ n_4986;
assign n_4989 = n_4987 & n_4988;
assign n_4990 = n_4989 ^ x80;
assign n_4991 = n_4990 ^ x81;
assign n_4992 = n_4871 ^ n_4990;
assign n_4993 = n_4991 & n_4992;
assign n_4994 = n_4993 ^ x81;
assign n_4995 = n_4994 ^ x82;
assign n_4996 = n_4872 ^ n_4994;
assign n_4997 = n_4995 & n_4996;
assign n_4998 = n_4997 ^ x82;
assign n_4999 = n_4998 ^ x83;
assign n_5000 = n_4884 ^ n_4998;
assign n_5001 = n_4999 & n_5000;
assign n_5002 = n_5001 ^ x83;
assign n_5003 = n_5002 ^ x84;
assign n_5004 = n_4873 ^ n_5002;
assign n_5005 = n_5003 & n_5004;
assign n_5006 = n_5005 ^ x84;
assign n_5007 = n_5006 ^ x85;
assign n_5008 = n_4885 ^ n_5006;
assign n_5009 = n_5007 & n_5008;
assign n_5010 = n_5009 ^ x85;
assign n_5011 = n_5010 ^ x86;
assign n_5012 = n_4874 ^ n_5010;
assign n_5013 = n_5011 & n_5012;
assign n_5014 = n_5013 ^ x86;
assign n_5015 = n_5014 ^ x87;
assign n_5016 = n_4875 ^ n_5014;
assign n_5017 = n_5015 & n_5016;
assign n_5018 = n_5017 ^ x87;
assign n_5019 = n_5018 ^ x88;
assign n_5020 = n_4876 ^ n_5018;
assign n_5021 = n_5019 & n_5020;
assign n_5022 = n_5021 ^ x88;
assign n_5023 = n_5022 ^ x89;
assign n_5024 = n_5022 ^ n_4883;
assign n_5025 = n_4924 & n_5022;
assign n_5026 = n_5023 & n_5024;
assign n_5027 = ~n_4932 & ~n_5025;
assign n_5028 = n_5026 ^ x89;
assign n_5029 = x91 ^ n_5027;
assign n_5030 = n_4877 ^ n_5027;
assign n_5031 = n_5028 ^ x90;
assign n_5032 = ~n_5029 & ~n_5030;
assign n_5033 = n_5032 ^ x91;
assign n_5034 = n_5033 ^ x92;
assign n_5035 = n_4878 ^ n_5033;
assign n_5036 = n_5034 & n_5035;
assign n_5037 = n_5036 ^ x92;
assign n_5038 = n_5037 ^ n_4851;
assign n_5039 = n_5037 ^ x93;
assign n_5040 = ~n_4894 & n_5038;
assign n_5041 = n_5040 ^ x93;
assign n_5042 = n_5041 ^ n_4882;
assign n_5043 = n_5041 ^ x94;
assign n_5044 = ~n_4904 & n_5042;
assign n_5045 = n_5044 ^ x94;
assign n_5046 = n_5045 ^ x95;
assign n_5047 = n_4879 ^ n_5045;
assign n_5048 = n_5046 & n_5047;
assign n_5049 = n_5048 ^ x95;
assign n_5050 = n_5049 ^ x96;
assign n_5051 = n_5049 ^ n_4850;
assign n_5052 = n_4919 & n_5049;
assign n_5053 = n_5050 & n_5051;
assign n_5054 = ~n_4928 & ~n_5052;
assign n_5055 = n_5053 ^ x96;
assign n_5056 = x98 ^ n_5054;
assign n_5057 = n_4880 ^ n_5054;
assign n_5058 = n_5055 ^ x97;
assign n_5059 = ~n_5056 & ~n_5057;
assign n_5060 = n_5059 ^ x98;
assign n_5061 = n_5060 ^ x99;
assign n_5062 = n_4881 ^ n_5060;
assign n_5063 = n_5061 & n_5062;
assign n_5064 = n_5063 ^ x99;
assign n_5065 = n_5064 ^ x100;
assign n_5066 = n_4926 & n_5064;
assign n_5067 = n_5064 & n_4888;
assign n_5068 = ~n_5066 & n_4933;
assign n_5069 = n_5065 & n_5068;
assign n_5070 = ~n_439 & n_5068;
assign n_5071 = n_5068 & ~n_5067;
assign n_5072 = n_5069 ^ n_4846;
assign n_5073 = n_4847 & ~n_5070;
assign n_5074 = n_5023 & n_5071;
assign n_5075 = x65 & n_5071;
assign n_5076 = x64 & n_5071;
assign n_5077 = x65 ^ n_5071;
assign n_5078 = n_4931 & n_5071;
assign n_5079 = n_4936 & n_5071;
assign n_5080 = n_4940 & n_5071;
assign n_5081 = n_4944 & n_5071;
assign n_5082 = n_4948 & n_5071;
assign n_5083 = n_4952 & n_5071;
assign n_5084 = n_4956 & n_5071;
assign n_5085 = n_4960 & n_5071;
assign n_5086 = n_4964 & n_5071;
assign n_5087 = n_4968 & n_5071;
assign n_5088 = n_4972 & n_5071;
assign n_5089 = n_4976 & n_5071;
assign n_5090 = ~n_4982 & n_5071;
assign n_5091 = n_4987 & n_5071;
assign n_5092 = n_4991 & n_5071;
assign n_5093 = n_4995 & n_5071;
assign n_5094 = n_4999 & n_5071;
assign n_5095 = n_5003 & n_5071;
assign n_5096 = n_5007 & n_5071;
assign n_5097 = n_5011 & n_5071;
assign n_5098 = n_5015 & n_5071;
assign n_5099 = n_5019 & n_5071;
assign n_5100 = n_5034 & n_5071;
assign n_5101 = ~n_5029 & n_5071;
assign n_5102 = n_5039 & n_5071;
assign n_5103 = n_5043 & n_5071;
assign n_5104 = n_5046 & n_5071;
assign n_5105 = n_5050 & n_5071;
assign n_5106 = ~n_5056 & n_5071;
assign n_5107 = n_5061 & n_5071;
assign y26 = n_5071;
assign n_5108 = n_5031 & n_5071;
assign n_5109 = n_4984 & n_5071;
assign n_5110 = n_5058 & n_5071;
assign n_5111 = x102 ^ n_5073;
assign n_5112 = n_5074 ^ n_4883;
assign n_5113 = n_5075 ^ n_4818;
assign n_5114 = ~x26 & n_5076;
assign n_5115 = n_5076 & n_212;
assign n_5116 = n_5077 ^ n_5075;
assign n_5117 = n_5078 ^ n_4901;
assign n_5118 = n_5079 ^ n_4859;
assign n_5119 = n_5080 ^ n_4860;
assign n_5120 = n_5081 ^ n_4861;
assign n_5121 = n_5082 ^ n_4862;
assign n_5122 = n_5083 ^ n_4863;
assign n_5123 = n_5084 ^ n_4864;
assign n_5124 = n_5085 ^ n_4865;
assign n_5125 = n_5086 ^ n_4866;
assign n_5126 = n_5087 ^ n_4867;
assign n_5127 = n_5088 ^ n_4868;
assign n_5128 = n_5089 ^ n_4854;
assign n_5129 = n_5090 ^ n_4869;
assign n_5130 = n_5091 ^ n_4870;
assign n_5131 = n_5092 ^ n_4871;
assign n_5132 = n_5093 ^ n_4872;
assign n_5133 = n_5094 ^ n_4884;
assign n_5134 = n_5095 ^ n_4873;
assign n_5135 = n_5096 ^ n_4885;
assign n_5136 = n_5097 ^ n_4874;
assign n_5137 = n_5098 ^ n_4875;
assign n_5138 = n_5099 ^ n_4876;
assign n_5139 = n_5100 ^ n_4878;
assign n_5140 = n_5101 ^ n_4877;
assign n_5141 = n_5102 ^ n_4851;
assign n_5142 = n_5103 ^ n_4882;
assign n_5143 = n_5104 ^ n_4879;
assign n_5144 = n_5105 ^ n_4850;
assign n_5145 = n_5106 ^ n_4880;
assign n_5146 = n_5107 ^ n_4881;
assign n_5147 = n_4852 ^ n_5108;
assign n_5148 = n_4853 ^ n_5109;
assign n_5149 = n_4849 ^ n_5110;
assign n_5150 = n_5112 ^ x90;
assign n_5151 = x90 & ~n_5112;
assign n_5152 = n_5113 ^ n_5114;
assign n_5153 = n_5115 ^ n_80;
assign n_5154 = n_5116 ^ x26;
assign n_5155 = ~x93 ^ n_5139;
assign n_5156 = n_5139 ^ x93;
assign n_5157 = n_5140 ^ x92;
assign n_5158 = x92 & ~n_5140;
assign n_5159 = ~x91 ^ n_5147;
assign n_5160 = n_5147 ^ x91;
assign n_5161 = n_5150 ^ n_5151;
assign n_5162 = n_5151 ^ n_5147;
assign n_5163 = n_5152 ^ x27;
assign n_5164 = n_21 & ~n_5154;
assign n_5165 = n_5157 ^ n_5158;
assign n_5166 = n_5158 ^ n_5139;
assign n_5167 = n_5159 & ~n_5161;
assign n_5168 = ~n_5160 & n_5162;
assign n_5169 = n_5163 ^ x66;
assign n_5170 = n_5153 ^ n_5164;
assign n_5171 = n_5155 & ~n_5165;
assign n_5172 = ~n_5156 & n_5166;
assign n_5173 = n_5168 ^ x91;
assign n_5174 = n_5170 ^ n_5163;
assign n_5175 = n_5170 ^ x66;
assign n_5176 = n_5172 ^ x93;
assign n_5177 = ~n_5169 & n_5174;
assign n_5178 = n_5177 ^ x66;
assign n_5179 = n_5178 ^ x67;
assign n_5180 = n_5117 ^ n_5178;
assign n_5181 = n_5179 & n_5180;
assign n_5182 = n_5181 ^ x67;
assign n_5183 = n_5182 ^ x68;
assign n_5184 = n_5118 ^ n_5182;
assign n_5185 = n_5183 & n_5184;
assign n_5186 = n_5185 ^ x68;
assign n_5187 = n_5186 ^ x69;
assign n_5188 = n_5119 ^ n_5186;
assign n_5189 = n_5187 & n_5188;
assign n_5190 = n_5189 ^ x69;
assign n_5191 = n_5190 ^ x70;
assign n_5192 = n_5120 ^ n_5190;
assign n_5193 = n_5191 & n_5192;
assign n_5194 = n_5193 ^ x70;
assign n_5195 = n_5194 ^ x71;
assign n_5196 = n_5121 ^ n_5194;
assign n_5197 = n_5195 & ~n_5196;
assign n_5198 = n_5197 ^ x71;
assign n_5199 = n_5198 ^ x72;
assign n_5200 = n_5122 ^ n_5198;
assign n_5201 = n_5199 & n_5200;
assign n_5202 = n_5201 ^ x72;
assign n_5203 = n_5202 ^ x73;
assign n_5204 = n_5123 ^ n_5202;
assign n_5205 = n_5203 & n_5204;
assign n_5206 = n_5205 ^ x73;
assign n_5207 = n_5206 ^ x74;
assign n_5208 = n_5124 ^ n_5206;
assign n_5209 = n_5207 & n_5208;
assign n_5210 = n_5209 ^ x74;
assign n_5211 = n_5210 ^ x75;
assign n_5212 = n_5125 ^ n_5210;
assign n_5213 = n_5211 & n_5212;
assign n_5214 = n_5213 ^ x75;
assign n_5215 = n_5214 ^ x76;
assign n_5216 = n_5126 ^ n_5214;
assign n_5217 = n_5215 & n_5216;
assign n_5218 = n_5217 ^ x76;
assign n_5219 = n_5218 ^ x77;
assign n_5220 = n_5127 ^ n_5218;
assign n_5221 = n_5219 & n_5220;
assign n_5222 = n_5221 ^ x77;
assign n_5223 = n_5222 ^ x78;
assign n_5224 = n_5128 ^ n_5222;
assign n_5225 = n_5223 & n_5224;
assign n_5226 = n_5225 ^ x78;
assign n_5227 = n_5226 ^ x79;
assign n_5228 = n_5148 ^ n_5226;
assign n_5229 = n_5227 & n_5228;
assign n_5230 = n_5229 ^ x79;
assign n_5231 = n_5230 ^ x80;
assign n_5232 = n_5129 ^ n_5230;
assign n_5233 = n_5231 & n_5232;
assign n_5234 = n_5233 ^ x80;
assign n_5235 = n_5234 ^ x81;
assign n_5236 = n_5130 ^ n_5234;
assign n_5237 = n_5235 & n_5236;
assign n_5238 = n_5237 ^ x81;
assign n_5239 = n_5238 ^ x82;
assign n_5240 = n_5131 ^ n_5238;
assign n_5241 = n_5239 & n_5240;
assign n_5242 = n_5241 ^ x82;
assign n_5243 = n_5242 ^ x83;
assign n_5244 = n_5132 ^ n_5242;
assign n_5245 = n_5243 & n_5244;
assign n_5246 = n_5245 ^ x83;
assign n_5247 = n_5246 ^ x84;
assign n_5248 = n_5133 ^ n_5246;
assign n_5249 = n_5247 & n_5248;
assign n_5250 = n_5249 ^ x84;
assign n_5251 = n_5250 ^ x85;
assign n_5252 = n_5134 ^ n_5250;
assign n_5253 = n_5251 & n_5252;
assign n_5254 = n_5253 ^ x85;
assign n_5255 = n_5254 ^ x86;
assign n_5256 = n_5135 ^ n_5254;
assign n_5257 = n_5255 & n_5256;
assign n_5258 = n_5257 ^ x86;
assign n_5259 = n_5258 ^ x87;
assign n_5260 = n_5136 ^ n_5258;
assign n_5261 = n_5259 & n_5260;
assign n_5262 = n_5261 ^ x87;
assign n_5263 = n_5262 ^ x88;
assign n_5264 = n_5137 ^ n_5262;
assign n_5265 = n_5263 & n_5264;
assign n_5266 = n_5265 ^ x88;
assign n_5267 = n_5266 ^ x89;
assign n_5268 = n_5138 ^ n_5266;
assign n_5269 = n_5267 & n_5268;
assign n_5270 = n_5269 ^ x89;
assign n_5271 = n_5270 ^ x90;
assign n_5272 = n_5270 ^ n_5112;
assign n_5273 = n_5167 & n_5270;
assign n_5274 = n_5271 & n_5272;
assign n_5275 = ~n_5173 & ~n_5273;
assign n_5276 = n_5274 ^ x90;
assign n_5277 = x92 ^ n_5275;
assign n_5278 = n_5140 ^ n_5275;
assign n_5279 = n_5171 & ~n_5275;
assign n_5280 = n_5276 ^ x91;
assign n_5281 = ~n_5277 & ~n_5278;
assign n_5282 = ~n_5176 & ~n_5279;
assign n_5283 = n_5281 ^ x92;
assign n_5284 = x94 ^ n_5282;
assign n_5285 = n_5141 ^ n_5282;
assign n_5286 = n_5283 ^ x93;
assign n_5287 = ~n_5284 & ~n_5285;
assign n_5288 = n_5287 ^ x94;
assign n_5289 = n_5288 ^ x95;
assign n_5290 = n_5142 ^ n_5288;
assign n_5291 = n_5289 & n_5290;
assign n_5292 = n_5291 ^ x95;
assign n_5293 = n_5292 ^ x96;
assign n_5294 = n_5143 ^ n_5292;
assign n_5295 = n_5293 & n_5294;
assign n_5296 = n_5295 ^ x96;
assign n_5297 = n_5296 ^ x97;
assign n_5298 = n_5144 ^ n_5296;
assign n_5299 = n_5297 & n_5298;
assign n_5300 = n_5299 ^ x97;
assign n_5301 = n_5300 ^ x98;
assign n_5302 = n_5149 ^ n_5300;
assign n_5303 = n_5301 & n_5302;
assign n_5304 = n_5303 ^ x98;
assign n_5305 = n_5304 ^ x99;
assign n_5306 = n_5145 ^ n_5304;
assign n_5307 = n_5305 & n_5306;
assign n_5308 = n_5307 ^ x99;
assign n_5309 = n_5308 ^ x100;
assign n_5310 = n_5146 ^ n_5308;
assign n_5311 = n_5309 & n_5310;
assign n_5312 = n_5311 ^ x100;
assign n_5313 = n_5312 ^ x101;
assign n_5314 = n_5072 ^ n_5312;
assign n_5315 = n_5313 & n_5314;
assign n_5316 = n_5315 ^ x101;
assign n_5317 = n_366 & ~n_5316;
assign n_5318 = n_5316 ^ x102;
assign n_5319 = ~n_5317 & n_4848;
assign n_5320 = ~n_5111 & n_5318;
assign n_5321 = ~n_439 ^ ~n_5319;
assign n_5322 = x102 ^ n_5320;
assign n_5323 = ~x103 & n_5321;
assign n_5324 = n_366 & ~n_5322;
assign n_5325 = x102 & ~n_5323;
assign n_5326 = n_5313 & n_5324;
assign n_5327 = n_5297 & n_5324;
assign n_5328 = n_5293 & n_5324;
assign n_5329 = n_5195 & n_5324;
assign n_5330 = n_5191 & n_5324;
assign n_5331 = n_153 & n_5324;
assign n_5332 = x64 & n_5324;
assign n_5333 = n_5175 & n_5324;
assign n_5334 = n_5179 & n_5324;
assign n_5335 = n_5183 & n_5324;
assign n_5336 = n_5187 & n_5324;
assign n_5337 = n_5199 & n_5324;
assign n_5338 = n_5203 & n_5324;
assign n_5339 = n_5207 & n_5324;
assign n_5340 = n_5211 & n_5324;
assign n_5341 = n_5215 & n_5324;
assign n_5342 = n_5219 & n_5324;
assign n_5343 = n_5223 & n_5324;
assign n_5344 = n_5227 & n_5324;
assign n_5345 = n_5231 & n_5324;
assign n_5346 = n_5235 & n_5324;
assign n_5347 = n_5239 & n_5324;
assign n_5348 = n_5243 & n_5324;
assign n_5349 = n_5247 & n_5324;
assign n_5350 = n_5251 & n_5324;
assign n_5351 = n_5255 & n_5324;
assign n_5352 = n_5259 & n_5324;
assign n_5353 = n_5263 & n_5324;
assign n_5354 = n_5267 & n_5324;
assign n_5355 = n_5271 & n_5324;
assign n_5356 = ~n_5277 & n_5324;
assign n_5357 = ~n_5284 & n_5324;
assign n_5358 = n_5289 & n_5324;
assign n_5359 = n_5301 & n_5324;
assign n_5360 = n_5305 & n_5324;
assign n_5361 = n_5309 & n_5324;
assign y25 = n_5324;
assign n_5362 = n_5280 & n_5324;
assign n_5363 = n_5286 & n_5324;
assign n_5364 = n_5326 ^ n_5072;
assign n_5365 = n_5327 ^ n_5144;
assign n_5366 = n_5328 ^ n_5143;
assign n_5367 = n_5329 ^ n_5121;
assign n_5368 = n_5330 ^ n_5120;
assign n_5369 = n_5331 ^ n_5076;
assign n_5370 = n_5332 ^ x24;
assign n_5371 = n_5332 ^ x65;
assign n_5372 = n_5333 ^ n_5163;
assign n_5373 = n_5334 ^ n_5117;
assign n_5374 = n_5335 ^ n_5118;
assign n_5375 = n_5336 ^ n_5119;
assign n_5376 = n_5337 ^ n_5122;
assign n_5377 = n_5338 ^ n_5123;
assign n_5378 = n_5339 ^ n_5124;
assign n_5379 = n_5340 ^ n_5125;
assign n_5380 = n_5341 ^ n_5126;
assign n_5381 = n_5342 ^ n_5127;
assign n_5382 = n_5343 ^ n_5128;
assign n_5383 = n_5344 ^ n_5148;
assign n_5384 = n_5345 ^ n_5129;
assign n_5385 = n_5346 ^ n_5130;
assign n_5386 = n_5347 ^ n_5131;
assign n_5387 = n_5348 ^ n_5132;
assign n_5388 = n_5349 ^ n_5133;
assign n_5389 = n_5350 ^ n_5134;
assign n_5390 = n_5351 ^ n_5135;
assign n_5391 = n_5352 ^ n_5136;
assign n_5392 = n_5353 ^ n_5137;
assign n_5393 = n_5354 ^ n_5138;
assign n_5394 = n_5355 ^ n_5112;
assign n_5395 = n_5356 ^ n_5140;
assign n_5396 = n_5357 ^ n_5141;
assign n_5397 = n_5358 ^ n_5142;
assign n_5398 = n_5359 ^ n_5149;
assign n_5399 = n_5360 ^ n_5145;
assign n_5400 = n_5361 ^ n_5146;
assign n_5401 = n_5147 ^ n_5362;
assign n_5402 = n_5139 ^ n_5363;
assign n_5403 = ~x102 ^ n_5364;
assign n_5404 = ~n_5364 & n_5325;
assign n_5405 = n_5365 ^ x98;
assign n_5406 = n_5366 ^ x97;
assign n_5407 = ~x72 ^ ~n_5367;
assign n_5408 = n_5367 ^ x72;
assign n_5409 = n_5368 ^ x71;
assign n_5410 = x71 & ~n_5368;
assign n_5411 = n_5369 ^ x26;
assign n_5412 = n_5370 & n_5371;
assign n_5413 = n_5403 & ~n_5323;
assign n_5414 = ~n_5404 & ~n_4909;
assign n_5415 = n_5409 ^ n_5410;
assign n_5416 = n_5410 ^ n_5367;
assign n_5417 = n_5411 ^ x66;
assign n_5418 = n_213 ^ n_5412;
assign n_5419 = n_5407 & ~n_5415;
assign n_5420 = n_5408 & ~n_5416;
assign n_5421 = n_154 ^ n_5418;
assign n_5422 = n_5420 ^ x72;
assign n_5423 = n_5421 ^ n_212;
assign n_5424 = n_5423 ^ n_5411;
assign n_5425 = n_5423 ^ x66;
assign n_5426 = ~n_5417 & n_5424;
assign n_5427 = n_5426 ^ x66;
assign n_5428 = n_5427 ^ x67;
assign n_5429 = n_5372 ^ n_5427;
assign n_5430 = n_5428 & n_5429;
assign n_5431 = n_5430 ^ x67;
assign n_5432 = n_5431 ^ x68;
assign n_5433 = n_5373 ^ n_5431;
assign n_5434 = n_5432 & n_5433;
assign n_5435 = n_5434 ^ x68;
assign n_5436 = n_5435 ^ x69;
assign n_5437 = n_5374 ^ n_5435;
assign n_5438 = n_5436 & n_5437;
assign n_5439 = n_5438 ^ x69;
assign n_5440 = n_5439 ^ x70;
assign n_5441 = n_5375 ^ n_5439;
assign n_5442 = n_5440 & n_5441;
assign n_5443 = n_5442 ^ x70;
assign n_5444 = n_5443 ^ x71;
assign n_5445 = n_5443 ^ n_5368;
assign n_5446 = n_5419 & n_5443;
assign n_5447 = n_5444 & n_5445;
assign n_5448 = ~n_5422 & ~n_5446;
assign n_5449 = n_5447 ^ x71;
assign n_5450 = x73 ^ n_5448;
assign n_5451 = n_5376 ^ n_5448;
assign n_5452 = n_5449 ^ x72;
assign n_5453 = ~n_5450 & ~n_5451;
assign n_5454 = n_5453 ^ x73;
assign n_5455 = n_5454 ^ x74;
assign n_5456 = n_5377 ^ n_5454;
assign n_5457 = n_5455 & n_5456;
assign n_5458 = n_5457 ^ x74;
assign n_5459 = n_5458 ^ x75;
assign n_5460 = n_5378 ^ n_5458;
assign n_5461 = n_5459 & n_5460;
assign n_5462 = n_5461 ^ x75;
assign n_5463 = n_5462 ^ x76;
assign n_5464 = n_5379 ^ n_5462;
assign n_5465 = n_5463 & n_5464;
assign n_5466 = n_5465 ^ x76;
assign n_5467 = n_5466 ^ x77;
assign n_5468 = n_5380 ^ n_5466;
assign n_5469 = n_5467 & n_5468;
assign n_5470 = n_5469 ^ x77;
assign n_5471 = n_5470 ^ x78;
assign n_5472 = n_5381 ^ n_5470;
assign n_5473 = n_5471 & n_5472;
assign n_5474 = n_5473 ^ x78;
assign n_5475 = n_5474 ^ x79;
assign n_5476 = n_5382 ^ n_5474;
assign n_5477 = n_5475 & n_5476;
assign n_5478 = n_5477 ^ x79;
assign n_5479 = n_5478 ^ x80;
assign n_5480 = n_5383 ^ n_5478;
assign n_5481 = n_5479 & n_5480;
assign n_5482 = n_5481 ^ x80;
assign n_5483 = n_5482 ^ x81;
assign n_5484 = n_5384 ^ n_5482;
assign n_5485 = n_5483 & n_5484;
assign n_5486 = n_5485 ^ x81;
assign n_5487 = n_5486 ^ x82;
assign n_5488 = n_5385 ^ n_5486;
assign n_5489 = n_5487 & n_5488;
assign n_5490 = n_5489 ^ x82;
assign n_5491 = n_5490 ^ x83;
assign n_5492 = n_5386 ^ n_5490;
assign n_5493 = n_5491 & n_5492;
assign n_5494 = n_5493 ^ x83;
assign n_5495 = n_5494 ^ x84;
assign n_5496 = n_5387 ^ n_5494;
assign n_5497 = n_5495 & n_5496;
assign n_5498 = n_5497 ^ x84;
assign n_5499 = n_5498 ^ x85;
assign n_5500 = n_5388 ^ n_5498;
assign n_5501 = n_5499 & n_5500;
assign n_5502 = n_5501 ^ x85;
assign n_5503 = n_5502 ^ x86;
assign n_5504 = n_5389 ^ n_5502;
assign n_5505 = n_5503 & n_5504;
assign n_5506 = n_5505 ^ x86;
assign n_5507 = n_5506 ^ x87;
assign n_5508 = n_5390 ^ n_5506;
assign n_5509 = n_5507 & n_5508;
assign n_5510 = n_5509 ^ x87;
assign n_5511 = n_5510 ^ x88;
assign n_5512 = n_5391 ^ n_5510;
assign n_5513 = n_5511 & n_5512;
assign n_5514 = n_5513 ^ x88;
assign n_5515 = n_5514 ^ x89;
assign n_5516 = n_5392 ^ n_5514;
assign n_5517 = n_5515 & n_5516;
assign n_5518 = n_5517 ^ x89;
assign n_5519 = n_5518 ^ x90;
assign n_5520 = n_5393 ^ n_5518;
assign n_5521 = n_5519 & n_5520;
assign n_5522 = n_5521 ^ x90;
assign n_5523 = n_5522 ^ x91;
assign n_5524 = n_5394 ^ n_5522;
assign n_5525 = n_5523 & n_5524;
assign n_5526 = n_5525 ^ x91;
assign n_5527 = n_5526 ^ x92;
assign n_5528 = n_5401 ^ n_5526;
assign n_5529 = n_5527 & n_5528;
assign n_5530 = n_5529 ^ x92;
assign n_5531 = n_5530 ^ x93;
assign n_5532 = n_5395 ^ n_5530;
assign n_5533 = n_5531 & n_5532;
assign n_5534 = n_5533 ^ x93;
assign n_5535 = n_5534 ^ x94;
assign n_5536 = n_5402 ^ n_5534;
assign n_5537 = n_5535 & n_5536;
assign n_5538 = n_5537 ^ x94;
assign n_5539 = n_5538 ^ x95;
assign n_5540 = n_5396 ^ n_5538;
assign n_5541 = n_5539 & n_5540;
assign n_5542 = n_5541 ^ x95;
assign n_5543 = n_5542 ^ x96;
assign n_5544 = n_5397 ^ n_5542;
assign n_5545 = n_5543 & n_5544;
assign n_5546 = n_5545 ^ x96;
assign n_5547 = n_5546 ^ n_5366;
assign n_5548 = n_5546 ^ x97;
assign n_5549 = ~n_5406 & n_5547;
assign n_5550 = n_5549 ^ x97;
assign n_5551 = n_5550 ^ n_5365;
assign n_5552 = n_5550 ^ x98;
assign n_5553 = ~n_5405 & n_5551;
assign n_5554 = n_5553 ^ x98;
assign n_5555 = n_5554 ^ x99;
assign n_5556 = n_5398 ^ n_5554;
assign n_5557 = n_5555 & n_5556;
assign n_5558 = n_5557 ^ x99;
assign n_5559 = n_5558 ^ x100;
assign n_5560 = n_5399 ^ n_5558;
assign n_5561 = n_5559 & n_5560;
assign n_5562 = n_5561 ^ x100;
assign n_5563 = n_5562 ^ x101;
assign n_5564 = n_5400 ^ n_5562;
assign n_5565 = n_5563 & n_5564;
assign n_5566 = n_5565 ^ x101;
assign n_5567 = n_5566 ^ x102;
assign n_5568 = n_5413 & n_5566;
assign n_5569 = ~n_5568 & n_5414;
assign n_5570 = n_5319 & ~n_5569;
assign n_5571 = n_5567 & n_5569;
assign n_5572 = n_5543 & n_5569;
assign n_5573 = n_5539 & n_5569;
assign n_5574 = n_5527 & n_5569;
assign n_5575 = n_5523 & n_5569;
assign n_5576 = n_5503 & n_5569;
assign n_5577 = n_5499 & n_5569;
assign n_5578 = x64 & n_5569;
assign n_5579 = x65 ^ n_5569;
assign n_5580 = n_5425 & n_5569;
assign n_5581 = n_5428 & n_5569;
assign n_5582 = n_5432 & n_5569;
assign n_5583 = n_5436 & n_5569;
assign n_5584 = n_5440 & n_5569;
assign n_5585 = n_5444 & n_5569;
assign n_5586 = ~n_5450 & n_5569;
assign n_5587 = n_5455 & n_5569;
assign n_5588 = n_5459 & n_5569;
assign n_5589 = n_5463 & n_5569;
assign n_5590 = n_5467 & n_5569;
assign n_5591 = n_5471 & n_5569;
assign n_5592 = n_5475 & n_5569;
assign n_5593 = n_5479 & n_5569;
assign n_5594 = n_5483 & n_5569;
assign n_5595 = n_5487 & n_5569;
assign n_5596 = n_5491 & n_5569;
assign n_5597 = n_5495 & n_5569;
assign n_5598 = n_5511 & n_5569;
assign n_5599 = n_5507 & n_5569;
assign n_5600 = n_5515 & n_5569;
assign n_5601 = n_5519 & n_5569;
assign n_5602 = n_5531 & n_5569;
assign n_5603 = n_5535 & n_5569;
assign n_5604 = n_5548 & n_5569;
assign n_5605 = n_5552 & n_5569;
assign n_5606 = n_5555 & n_5569;
assign n_5607 = n_5559 & n_5569;
assign n_5608 = n_5563 & n_5569;
assign n_5609 = n_23 ^ n_5569;
assign y24 = n_5569;
assign n_5610 = n_155 & n_5569;
assign n_5611 = n_5452 & n_5569;
assign n_5612 = ~n_439 ^ ~n_5570;
assign n_5613 = n_5571 ^ n_5364;
assign n_5614 = n_5572 ^ n_5397;
assign n_5615 = n_5573 ^ n_5396;
assign n_5616 = n_5574 ^ n_5401;
assign n_5617 = n_5575 ^ n_5394;
assign n_5618 = n_5576 ^ n_5389;
assign n_5619 = n_5577 ^ n_5388;
assign n_5620 = x65 & n_5578;
assign n_5621 = n_5578 ^ x24;
assign n_5622 = n_5579 ^ x24;
assign n_5623 = n_5580 ^ n_5411;
assign n_5624 = n_5581 ^ n_5372;
assign n_5625 = n_5582 ^ n_5373;
assign n_5626 = n_5583 ^ n_5374;
assign n_5627 = n_5584 ^ n_5375;
assign n_5628 = n_5585 ^ n_5368;
assign n_5629 = n_5586 ^ n_5376;
assign n_5630 = n_5587 ^ n_5377;
assign n_5631 = n_5588 ^ n_5378;
assign n_5632 = n_5589 ^ n_5379;
assign n_5633 = n_5590 ^ n_5380;
assign n_5634 = n_5591 ^ n_5381;
assign n_5635 = n_5592 ^ n_5382;
assign n_5636 = n_5593 ^ n_5383;
assign n_5637 = n_5594 ^ n_5384;
assign n_5638 = n_5595 ^ n_5385;
assign n_5639 = n_5596 ^ n_5386;
assign n_5640 = n_5597 ^ n_5387;
assign n_5641 = n_5598 ^ n_5391;
assign n_5642 = n_5599 ^ n_5390;
assign n_5643 = n_5600 ^ n_5392;
assign n_5644 = n_5601 ^ n_5393;
assign n_5645 = n_5602 ^ n_5395;
assign n_5646 = n_5603 ^ n_5402;
assign n_5647 = n_5604 ^ n_5366;
assign n_5648 = n_5605 ^ n_5365;
assign n_5649 = n_5606 ^ n_5398;
assign n_5650 = n_5607 ^ n_5399;
assign n_5651 = n_5608 ^ n_5400;
assign n_5652 = n_5609 ^ n_5579;
assign n_5653 = n_5332 ^ n_5610;
assign n_5654 = n_5367 ^ n_5611;
assign n_5655 = ~n_5612 ^ x104;
assign n_5656 = n_5613 ^ x103;
assign n_5657 = n_5614 ^ x97;
assign n_5658 = n_5615 ^ x96;
assign n_5659 = ~x93 ^ n_5616;
assign n_5660 = n_5616 ^ x93;
assign n_5661 = n_5617 ^ x92;
assign n_5662 = x92 & ~n_5617;
assign n_5663 = ~x87 ^ n_5618;
assign n_5664 = n_5618 ^ x87;
assign n_5665 = n_5619 ^ x86;
assign n_5666 = x86 & ~n_5619;
assign n_5667 = n_5620 ^ n_82;
assign n_5668 = n_23 & ~n_5622;
assign n_5669 = ~x89 ^ n_5641;
assign n_5670 = n_5641 ^ x89;
assign n_5671 = n_5642 ^ x88;
assign n_5672 = x88 & ~n_5642;
assign n_5673 = n_5653 ^ x25;
assign n_5674 = n_5661 ^ n_5662;
assign n_5675 = n_5662 ^ n_5616;
assign n_5676 = n_5665 ^ n_5666;
assign n_5677 = n_5666 ^ n_5618;
assign n_5678 = n_5667 ^ n_5668;
assign n_5679 = n_5671 ^ n_5672;
assign n_5680 = n_5672 ^ n_5641;
assign n_5681 = n_5673 ^ x66;
assign n_5682 = n_5659 & ~n_5674;
assign n_5683 = ~n_5660 & n_5675;
assign n_5684 = n_5663 & ~n_5676;
assign n_5685 = ~n_5664 & n_5677;
assign n_5686 = n_5678 ^ n_5673;
assign n_5687 = n_5678 ^ x66;
assign n_5688 = n_5669 & ~n_5679;
assign n_5689 = ~n_5670 & n_5680;
assign n_5690 = n_5683 ^ x93;
assign n_5691 = n_5685 ^ x87;
assign n_5692 = ~n_5681 & n_5686;
assign n_5693 = n_5689 ^ x89;
assign n_5694 = n_5692 ^ x66;
assign n_5695 = n_5694 ^ x67;
assign n_5696 = n_5623 ^ n_5694;
assign n_5697 = n_5695 & n_5696;
assign n_5698 = n_5697 ^ x67;
assign n_5699 = n_5698 ^ x68;
assign n_5700 = n_5624 ^ n_5698;
assign n_5701 = n_5699 & n_5700;
assign n_5702 = n_5701 ^ x68;
assign n_5703 = n_5702 ^ x69;
assign n_5704 = n_5625 ^ n_5702;
assign n_5705 = n_5703 & n_5704;
assign n_5706 = n_5705 ^ x69;
assign n_5707 = n_5706 ^ x70;
assign n_5708 = n_5626 ^ n_5706;
assign n_5709 = n_5707 & n_5708;
assign n_5710 = n_5709 ^ x70;
assign n_5711 = n_5710 ^ x71;
assign n_5712 = n_5627 ^ n_5710;
assign n_5713 = n_5711 & n_5712;
assign n_5714 = n_5713 ^ x71;
assign n_5715 = n_5714 ^ x72;
assign n_5716 = n_5628 ^ n_5714;
assign n_5717 = n_5715 & n_5716;
assign n_5718 = n_5717 ^ x72;
assign n_5719 = n_5718 ^ x73;
assign n_5720 = n_5654 ^ n_5718;
assign n_5721 = n_5719 & ~n_5720;
assign n_5722 = n_5721 ^ x73;
assign n_5723 = n_5722 ^ x74;
assign n_5724 = n_5629 ^ n_5722;
assign n_5725 = n_5723 & n_5724;
assign n_5726 = n_5725 ^ x74;
assign n_5727 = n_5726 ^ x75;
assign n_5728 = n_5630 ^ n_5726;
assign n_5729 = n_5727 & n_5728;
assign n_5730 = n_5729 ^ x75;
assign n_5731 = n_5730 ^ x76;
assign n_5732 = n_5631 ^ n_5730;
assign n_5733 = n_5731 & n_5732;
assign n_5734 = n_5733 ^ x76;
assign n_5735 = n_5734 ^ x77;
assign n_5736 = n_5632 ^ n_5734;
assign n_5737 = n_5735 & n_5736;
assign n_5738 = n_5737 ^ x77;
assign n_5739 = n_5738 ^ x78;
assign n_5740 = n_5633 ^ n_5738;
assign n_5741 = n_5739 & n_5740;
assign n_5742 = n_5741 ^ x78;
assign n_5743 = n_5742 ^ x79;
assign n_5744 = n_5634 ^ n_5742;
assign n_5745 = n_5743 & n_5744;
assign n_5746 = n_5745 ^ x79;
assign n_5747 = n_5746 ^ x80;
assign n_5748 = n_5635 ^ n_5746;
assign n_5749 = n_5747 & n_5748;
assign n_5750 = n_5749 ^ x80;
assign n_5751 = n_5750 ^ x81;
assign n_5752 = n_5636 ^ n_5750;
assign n_5753 = n_5751 & n_5752;
assign n_5754 = n_5753 ^ x81;
assign n_5755 = n_5754 ^ x82;
assign n_5756 = n_5637 ^ n_5754;
assign n_5757 = n_5755 & n_5756;
assign n_5758 = n_5757 ^ x82;
assign n_5759 = n_5758 ^ x83;
assign n_5760 = n_5638 ^ n_5758;
assign n_5761 = n_5759 & n_5760;
assign n_5762 = n_5761 ^ x83;
assign n_5763 = n_5762 ^ x84;
assign n_5764 = n_5639 ^ n_5762;
assign n_5765 = n_5763 & n_5764;
assign n_5766 = n_5765 ^ x84;
assign n_5767 = n_5766 ^ x85;
assign n_5768 = n_5640 ^ n_5766;
assign n_5769 = n_5767 & n_5768;
assign n_5770 = n_5769 ^ x85;
assign n_5771 = n_5770 ^ x86;
assign n_5772 = n_5770 ^ n_5619;
assign n_5773 = n_5684 & n_5770;
assign n_5774 = n_5771 & n_5772;
assign n_5775 = ~n_5691 & ~n_5773;
assign n_5776 = n_5774 ^ x86;
assign n_5777 = x88 ^ n_5775;
assign n_5778 = n_5642 ^ n_5775;
assign n_5779 = n_5688 & ~n_5775;
assign n_5780 = n_5776 ^ x87;
assign n_5781 = ~n_5777 & ~n_5778;
assign n_5782 = ~n_5693 & ~n_5779;
assign n_5783 = n_5781 ^ x88;
assign n_5784 = x90 ^ n_5782;
assign n_5785 = n_5643 ^ n_5782;
assign n_5786 = n_5783 ^ x89;
assign n_5787 = ~n_5784 & ~n_5785;
assign n_5788 = n_5787 ^ x90;
assign n_5789 = n_5788 ^ x91;
assign n_5790 = n_5644 ^ n_5788;
assign n_5791 = n_5789 & n_5790;
assign n_5792 = n_5791 ^ x91;
assign n_5793 = n_5792 ^ x92;
assign n_5794 = n_5792 ^ n_5617;
assign n_5795 = n_5682 & n_5792;
assign n_5796 = n_5793 & n_5794;
assign n_5797 = ~n_5690 & ~n_5795;
assign n_5798 = n_5796 ^ x92;
assign n_5799 = x94 ^ n_5797;
assign n_5800 = n_5645 ^ n_5797;
assign n_5801 = n_5798 ^ x93;
assign n_5802 = ~n_5799 & ~n_5800;
assign n_5803 = n_5802 ^ x94;
assign n_5804 = n_5803 ^ x95;
assign n_5805 = n_5646 ^ n_5803;
assign n_5806 = n_5804 & n_5805;
assign n_5807 = n_5806 ^ x95;
assign n_5808 = n_5807 ^ n_5615;
assign n_5809 = n_5807 ^ x96;
assign n_5810 = ~n_5658 & n_5808;
assign n_5811 = n_5810 ^ x96;
assign n_5812 = n_5811 ^ n_5614;
assign n_5813 = n_5811 ^ x97;
assign n_5814 = ~n_5657 & n_5812;
assign n_5815 = n_5814 ^ x97;
assign n_5816 = n_5815 ^ x98;
assign n_5817 = n_5647 ^ n_5815;
assign n_5818 = n_5816 & n_5817;
assign n_5819 = n_5818 ^ x98;
assign n_5820 = n_5819 ^ x99;
assign n_5821 = n_5648 ^ n_5819;
assign n_5822 = n_5820 & n_5821;
assign n_5823 = n_5822 ^ x99;
assign n_5824 = n_5823 ^ x100;
assign n_5825 = n_5649 ^ n_5823;
assign n_5826 = n_5824 & n_5825;
assign n_5827 = n_5826 ^ x100;
assign n_5828 = n_5827 ^ x101;
assign n_5829 = n_5650 ^ n_5827;
assign n_5830 = n_5828 & n_5829;
assign n_5831 = n_5830 ^ x101;
assign n_5832 = n_5831 ^ x102;
assign n_5833 = n_5651 ^ n_5831;
assign n_5834 = n_5832 & n_5833;
assign n_5835 = n_5834 ^ x102;
assign n_5836 = n_5835 ^ n_5613;
assign n_5837 = n_5835 ^ x103;
assign n_5838 = ~n_5656 & n_5836;
assign n_5839 = n_5838 ^ x103;
assign n_5840 = n_5839 ^ ~n_5612;
assign n_5841 = n_5655 & ~n_5840;
assign n_5842 = x104 ^ n_5841;
assign n_5843 = n_367 & ~n_5842;
assign n_5844 = n_5570 & ~n_5843;
assign n_5845 = n_5816 & n_5843;
assign n_5846 = n_5711 & n_5843;
assign n_5847 = n_5707 & n_5843;
assign n_5848 = n_5652 & n_5843;
assign n_5849 = x64 & n_5843;
assign n_5850 = n_5687 & n_5843;
assign n_5851 = n_5695 & n_5843;
assign n_5852 = n_5699 & n_5843;
assign n_5853 = n_5703 & n_5843;
assign n_5854 = n_5715 & n_5843;
assign n_5855 = n_5719 & n_5843;
assign n_5856 = n_5723 & n_5843;
assign n_5857 = n_5727 & n_5843;
assign n_5858 = n_5731 & n_5843;
assign n_5859 = n_5735 & n_5843;
assign n_5860 = n_5739 & n_5843;
assign n_5861 = n_5743 & n_5843;
assign n_5862 = n_5747 & n_5843;
assign n_5863 = n_5751 & n_5843;
assign n_5864 = n_5755 & n_5843;
assign n_5865 = n_5759 & n_5843;
assign n_5866 = n_5763 & n_5843;
assign n_5867 = n_5767 & n_5843;
assign n_5868 = n_5771 & n_5843;
assign n_5869 = ~n_5777 & n_5843;
assign n_5870 = ~n_5784 & n_5843;
assign n_5871 = n_5789 & n_5843;
assign n_5872 = n_5793 & n_5843;
assign n_5873 = ~n_5799 & n_5843;
assign n_5874 = n_5804 & n_5843;
assign n_5875 = n_5809 & n_5843;
assign n_5876 = n_5813 & n_5843;
assign n_5877 = n_5820 & n_5843;
assign n_5878 = n_5824 & n_5843;
assign n_5879 = n_5828 & n_5843;
assign n_5880 = n_5832 & n_5843;
assign n_5881 = n_5837 & n_5843;
assign y23 = n_5843;
assign n_5882 = n_5780 & n_5843;
assign n_5883 = n_5786 & n_5843;
assign n_5884 = n_5801 & n_5843;
assign n_5885 = ~n_439 ^ ~n_5844;
assign n_5886 = n_5845 ^ n_5647;
assign n_5887 = n_5846 ^ n_5627;
assign n_5888 = n_5847 ^ n_5626;
assign n_5889 = n_5848 ^ n_5621;
assign n_5890 = n_5849 ^ x23;
assign n_5891 = n_5850 ^ n_5673;
assign n_5892 = n_5851 ^ n_5623;
assign n_5893 = n_5852 ^ n_5624;
assign n_5894 = n_5853 ^ n_5625;
assign n_5895 = n_5854 ^ n_5628;
assign n_5896 = n_5855 ^ n_5654;
assign n_5897 = n_5856 ^ n_5629;
assign n_5898 = n_5857 ^ n_5630;
assign n_5899 = n_5858 ^ n_5631;
assign n_5900 = n_5859 ^ n_5632;
assign n_5901 = n_5860 ^ n_5633;
assign n_5902 = n_5861 ^ n_5634;
assign n_5903 = n_5862 ^ n_5635;
assign n_5904 = n_5863 ^ n_5636;
assign n_5905 = n_5864 ^ n_5637;
assign n_5906 = n_5865 ^ n_5638;
assign n_5907 = n_5866 ^ n_5639;
assign n_5908 = n_5867 ^ n_5640;
assign n_5909 = n_5868 ^ n_5619;
assign n_5910 = n_5869 ^ n_5642;
assign n_5911 = n_5870 ^ n_5643;
assign n_5912 = n_5871 ^ n_5644;
assign n_5913 = n_5872 ^ n_5617;
assign n_5914 = n_5873 ^ n_5645;
assign n_5915 = n_5874 ^ n_5646;
assign n_5916 = n_5875 ^ n_5615;
assign n_5917 = n_5876 ^ n_5614;
assign n_5918 = n_5877 ^ n_5648;
assign n_5919 = n_5878 ^ n_5649;
assign n_5920 = n_5879 ^ n_5650;
assign n_5921 = n_5880 ^ n_5651;
assign n_5922 = n_5881 ^ n_5613;
assign n_5923 = n_5618 ^ n_5882;
assign n_5924 = n_5641 ^ n_5883;
assign n_5925 = n_5616 ^ n_5884;
assign n_5926 = ~n_5885 ^ x105;
assign n_5927 = ~n_5885 ^ x106;
assign n_5928 = x107 & ~n_5885;
assign n_5929 = n_361 & n_5885;
assign n_5930 = x109 & ~n_5885;
assign n_5931 = n_5886 ^ x99;
assign n_5932 = n_5886 ^ x98;
assign n_5933 = ~x72 ^ n_5887;
assign n_5934 = n_5887 ^ x72;
assign n_5935 = n_5888 ^ x71;
assign n_5936 = x71 & ~n_5888;
assign n_5937 = n_5889 ^ x66;
assign n_5938 = n_5890 ^ x65;
assign n_5939 = n_24 ^ n_5890;
assign n_5940 = ~n_5890 & n_187;
assign n_5941 = n_5928 ^ x107;
assign n_5942 = n_362 & ~n_5928;
assign n_5943 = n_360 & ~n_5930;
assign n_5944 = n_5935 ^ n_5936;
assign n_5945 = n_5936 ^ n_5887;
assign n_5946 = ~n_5938 & ~n_305;
assign n_5947 = ~n_5938 & n_216;
assign n_5948 = ~n_5938 & n_5939;
assign n_5949 = n_5933 & ~n_5944;
assign n_5950 = ~n_5934 & n_5945;
assign n_5951 = ~n_5947 ^ ~n_5940;
assign n_5952 = n_5948 ^ x65;
assign n_5953 = n_5950 ^ x72;
assign n_5954 = n_5952 ^ n_5889;
assign n_5955 = n_5952 ^ x66;
assign n_5956 = ~n_5937 & n_5954;
assign n_5957 = n_5956 ^ x66;
assign n_5958 = n_5957 ^ x67;
assign n_5959 = n_5891 ^ n_5957;
assign n_5960 = n_5958 & n_5959;
assign n_5961 = n_5960 ^ x67;
assign n_5962 = n_5961 ^ x68;
assign n_5963 = n_5892 ^ n_5961;
assign n_5964 = n_5962 & n_5963;
assign n_5965 = n_5964 ^ x68;
assign n_5966 = n_5965 ^ x69;
assign n_5967 = n_5893 ^ n_5965;
assign n_5968 = n_5966 & n_5967;
assign n_5969 = n_5968 ^ x69;
assign n_5970 = n_5969 ^ x70;
assign n_5971 = n_5894 ^ n_5969;
assign n_5972 = n_5970 & n_5971;
assign n_5973 = n_5972 ^ x70;
assign n_5974 = n_5973 ^ x71;
assign n_5975 = n_5973 ^ n_5888;
assign n_5976 = n_5949 & n_5973;
assign n_5977 = n_5974 & n_5975;
assign n_5978 = ~n_5953 & ~n_5976;
assign n_5979 = n_5977 ^ x71;
assign n_5980 = x73 ^ n_5978;
assign n_5981 = n_5895 ^ n_5978;
assign n_5982 = n_5979 ^ x72;
assign n_5983 = ~n_5980 & ~n_5981;
assign n_5984 = n_5983 ^ x73;
assign n_5985 = n_5984 ^ x74;
assign n_5986 = n_5896 ^ n_5984;
assign n_5987 = n_5985 & ~n_5986;
assign n_5988 = n_5987 ^ x74;
assign n_5989 = n_5988 ^ x75;
assign n_5990 = n_5897 ^ n_5988;
assign n_5991 = n_5989 & n_5990;
assign n_5992 = n_5991 ^ x75;
assign n_5993 = n_5992 ^ x76;
assign n_5994 = n_5898 ^ n_5992;
assign n_5995 = n_5993 & n_5994;
assign n_5996 = n_5995 ^ x76;
assign n_5997 = n_5996 ^ x77;
assign n_5998 = n_5899 ^ n_5996;
assign n_5999 = n_5997 & n_5998;
assign n_6000 = n_5999 ^ x77;
assign n_6001 = n_6000 ^ x78;
assign n_6002 = n_5900 ^ n_6000;
assign n_6003 = n_6001 & n_6002;
assign n_6004 = n_6003 ^ x78;
assign n_6005 = n_6004 ^ x79;
assign n_6006 = n_5901 ^ n_6004;
assign n_6007 = n_6005 & n_6006;
assign n_6008 = n_6007 ^ x79;
assign n_6009 = n_6008 ^ x80;
assign n_6010 = n_5902 ^ n_6008;
assign n_6011 = n_6009 & n_6010;
assign n_6012 = n_6011 ^ x80;
assign n_6013 = n_6012 ^ x81;
assign n_6014 = n_5903 ^ n_6012;
assign n_6015 = n_6013 & n_6014;
assign n_6016 = n_6015 ^ x81;
assign n_6017 = n_6016 ^ x82;
assign n_6018 = n_5904 ^ n_6016;
assign n_6019 = n_6017 & n_6018;
assign n_6020 = n_6019 ^ x82;
assign n_6021 = n_6020 ^ x83;
assign n_6022 = n_5905 ^ n_6020;
assign n_6023 = n_6021 & n_6022;
assign n_6024 = n_6023 ^ x83;
assign n_6025 = n_6024 ^ x84;
assign n_6026 = n_5906 ^ n_6024;
assign n_6027 = n_6025 & n_6026;
assign n_6028 = n_6027 ^ x84;
assign n_6029 = n_6028 ^ x85;
assign n_6030 = n_5907 ^ n_6028;
assign n_6031 = n_6029 & n_6030;
assign n_6032 = n_6031 ^ x85;
assign n_6033 = n_6032 ^ x86;
assign n_6034 = n_5908 ^ n_6032;
assign n_6035 = n_6033 & n_6034;
assign n_6036 = n_6035 ^ x86;
assign n_6037 = n_6036 ^ x87;
assign n_6038 = n_5909 ^ n_6036;
assign n_6039 = n_6037 & n_6038;
assign n_6040 = n_6039 ^ x87;
assign n_6041 = n_6040 ^ x88;
assign n_6042 = n_5923 ^ n_6040;
assign n_6043 = n_6041 & n_6042;
assign n_6044 = n_6043 ^ x88;
assign n_6045 = n_6044 ^ x89;
assign n_6046 = n_5910 ^ n_6044;
assign n_6047 = n_6045 & n_6046;
assign n_6048 = n_6047 ^ x89;
assign n_6049 = n_6048 ^ x90;
assign n_6050 = n_5924 ^ n_6048;
assign n_6051 = n_6049 & n_6050;
assign n_6052 = n_6051 ^ x90;
assign n_6053 = n_6052 ^ x91;
assign n_6054 = n_5911 ^ n_6052;
assign n_6055 = n_6053 & n_6054;
assign n_6056 = n_6055 ^ x91;
assign n_6057 = n_6056 ^ x92;
assign n_6058 = n_5912 ^ n_6056;
assign n_6059 = n_6057 & n_6058;
assign n_6060 = n_6059 ^ x92;
assign n_6061 = n_6060 ^ x93;
assign n_6062 = n_5913 ^ n_6060;
assign n_6063 = n_6061 & n_6062;
assign n_6064 = n_6063 ^ x93;
assign n_6065 = n_6064 ^ x94;
assign n_6066 = n_5925 ^ n_6064;
assign n_6067 = n_6065 & n_6066;
assign n_6068 = n_6067 ^ x94;
assign n_6069 = n_6068 ^ x95;
assign n_6070 = n_5914 ^ n_6068;
assign n_6071 = n_6069 & n_6070;
assign n_6072 = n_6071 ^ x95;
assign n_6073 = n_6072 ^ x96;
assign n_6074 = n_5915 ^ n_6072;
assign n_6075 = n_6073 & n_6074;
assign n_6076 = n_6075 ^ x96;
assign n_6077 = n_6076 ^ x97;
assign n_6078 = n_5916 ^ n_6076;
assign n_6079 = n_6077 & n_6078;
assign n_6080 = n_6079 ^ x97;
assign n_6081 = n_6080 ^ x98;
assign n_6082 = n_5917 ^ n_6080;
assign n_6083 = n_6081 & n_6082;
assign n_6084 = n_5932 ^ n_6083;
assign n_6085 = n_6083 ^ x98;
assign n_6086 = ~n_5931 & n_6084;
assign n_6087 = n_6085 ^ x99;
assign n_6088 = n_6086 ^ x99;
assign n_6089 = n_6088 ^ x100;
assign n_6090 = n_5918 ^ n_6088;
assign n_6091 = n_6089 & n_6090;
assign n_6092 = n_6091 ^ x100;
assign n_6093 = n_6092 ^ x101;
assign n_6094 = n_5919 ^ n_6092;
assign n_6095 = n_6093 & n_6094;
assign n_6096 = n_6095 ^ x101;
assign n_6097 = n_6096 ^ x102;
assign n_6098 = n_5920 ^ n_6096;
assign n_6099 = n_6097 & n_6098;
assign n_6100 = n_6099 ^ x102;
assign n_6101 = n_6100 ^ x103;
assign n_6102 = n_5921 ^ n_6100;
assign n_6103 = n_6101 & n_6102;
assign n_6104 = n_6103 ^ x103;
assign n_6105 = n_6104 ^ x104;
assign n_6106 = n_5922 ^ n_6104;
assign n_6107 = n_6105 & n_6106;
assign n_6108 = n_6107 ^ x104;
assign n_6109 = n_6108 ^ x105;
assign n_6110 = n_6109 & n_5926;
assign n_6111 = n_5927 ^ n_6109;
assign n_6112 = n_6110 ^ x105;
assign n_6113 = n_6109 & ~n_6111;
assign n_6114 = n_364 & ~n_6112;
assign n_6115 = n_6113 ^ n_6109;
assign n_6116 = n_6087 & n_6114;
assign n_6117 = n_6081 & n_6114;
assign n_6118 = n_6057 & n_6114;
assign n_6119 = n_6053 & n_6114;
assign n_6120 = x64 & n_6114;
assign n_6121 = n_215 ^ n_6114;
assign n_6122 = n_5890 ^ n_6114;
assign n_6123 = n_5955 & n_6114;
assign n_6124 = n_5958 & n_6114;
assign n_6125 = n_5962 & n_6114;
assign n_6126 = n_5966 & n_6114;
assign n_6127 = n_5970 & n_6114;
assign n_6128 = n_5974 & n_6114;
assign n_6129 = ~n_5980 & n_6114;
assign n_6130 = n_5985 & n_6114;
assign n_6131 = n_5989 & n_6114;
assign n_6132 = n_5993 & n_6114;
assign n_6133 = n_5997 & n_6114;
assign n_6134 = n_6001 & n_6114;
assign n_6135 = n_6005 & n_6114;
assign n_6136 = n_6009 & n_6114;
assign n_6137 = n_6013 & n_6114;
assign n_6138 = n_6017 & n_6114;
assign n_6139 = n_6021 & n_6114;
assign n_6140 = n_6025 & n_6114;
assign n_6141 = n_6029 & n_6114;
assign n_6142 = n_6033 & n_6114;
assign n_6143 = n_6037 & n_6114;
assign n_6144 = n_6041 & n_6114;
assign n_6145 = n_6045 & n_6114;
assign n_6146 = n_6049 & n_6114;
assign n_6147 = n_6065 & n_6114;
assign n_6148 = n_6061 & n_6114;
assign n_6149 = n_6069 & n_6114;
assign n_6150 = n_6073 & n_6114;
assign n_6151 = n_6077 & n_6114;
assign n_6152 = n_6093 & n_6114;
assign n_6153 = n_6089 & n_6114;
assign n_6154 = n_6097 & n_6114;
assign n_6155 = n_6101 & n_6114;
assign n_6156 = n_6105 & n_6114;
assign n_6157 = n_157 & n_6114;
assign n_6158 = ~n_323 & ~n_6114;
assign y22 = n_6114;
assign n_6159 = n_5951 & n_6114;
assign n_6160 = n_5982 & n_6114;
assign n_6161 = n_6116 ^ n_5886;
assign n_6162 = n_6117 ^ n_5917;
assign n_6163 = n_6118 ^ n_5912;
assign n_6164 = n_6119 ^ n_5911;
assign n_6165 = ~n_6120 & n_85;
assign n_6166 = ~x21 & n_6120;
assign n_6167 = n_6120 & n_5946;
assign n_6168 = ~n_6122 & n_6114;
assign n_6169 = ~n_6122 & ~n_156;
assign n_6170 = n_6123 ^ n_5889;
assign n_6171 = n_6124 ^ n_5891;
assign n_6172 = n_6125 ^ n_5892;
assign n_6173 = n_6126 ^ n_5893;
assign n_6174 = n_6127 ^ n_5894;
assign n_6175 = n_6128 ^ n_5888;
assign n_6176 = n_6129 ^ n_5895;
assign n_6177 = n_6130 ^ n_5896;
assign n_6178 = n_6131 ^ n_5897;
assign n_6179 = n_6132 ^ n_5898;
assign n_6180 = n_6133 ^ n_5899;
assign n_6181 = n_6134 ^ n_5900;
assign n_6182 = n_6135 ^ n_5901;
assign n_6183 = n_6136 ^ n_5902;
assign n_6184 = n_6137 ^ n_5903;
assign n_6185 = n_6138 ^ n_5904;
assign n_6186 = n_6139 ^ n_5905;
assign n_6187 = n_6140 ^ n_5906;
assign n_6188 = n_6141 ^ n_5907;
assign n_6189 = n_6142 ^ n_5908;
assign n_6190 = n_6143 ^ n_5909;
assign n_6191 = n_6144 ^ n_5923;
assign n_6192 = n_6145 ^ n_5910;
assign n_6193 = n_6146 ^ n_5924;
assign n_6194 = n_6147 ^ n_5925;
assign n_6195 = n_6148 ^ n_5913;
assign n_6196 = n_6149 ^ n_5914;
assign n_6197 = n_6150 ^ n_5915;
assign n_6198 = n_6151 ^ n_5916;
assign n_6199 = n_6152 ^ n_5919;
assign n_6200 = n_6153 ^ n_5918;
assign n_6201 = n_6154 ^ n_5920;
assign n_6202 = n_6155 ^ n_5921;
assign n_6203 = n_6156 ^ n_5922;
assign n_6204 = n_6157 ^ n_5890;
assign n_6205 = n_6158 ^ n_305;
assign n_6206 = n_5887 ^ n_6160;
assign n_6207 = x100 ^ ~n_6161;
assign n_6208 = n_6161 ^ x100;
assign n_6209 = n_6162 ^ x99;
assign n_6210 = ~x99 & n_6162;
assign n_6211 = ~x93 ^ n_6163;
assign n_6212 = n_6163 ^ x93;
assign n_6213 = n_6164 ^ x92;
assign n_6214 = x92 & ~n_6164;
assign n_6215 = ~n_6122 & n_6165;
assign n_6216 = n_324 ^ ~n_6166;
assign n_6217 = ~x66 & ~n_6167;
assign n_6218 = n_6168 ^ n_6114;
assign n_6219 = n_5890 & ~n_6169;
assign n_6220 = ~x95 ^ n_6194;
assign n_6221 = n_6194 ^ x95;
assign n_6222 = n_6195 ^ x94;
assign n_6223 = x94 & ~n_6195;
assign n_6224 = ~x102 ^ n_6199;
assign n_6225 = n_6199 ^ x102;
assign n_6226 = n_6200 ^ x101;
assign n_6227 = x101 & ~n_6200;
assign n_6228 = ~n_83 & n_6205;
assign n_6229 = n_6209 ^ n_6210;
assign n_6230 = n_6210 ^ n_6161;
assign n_6231 = n_6213 ^ n_6214;
assign n_6232 = n_6214 ^ n_6163;
assign n_6233 = ~n_6121 & n_6218;
assign n_6234 = ~n_6216 & n_6219;
assign n_6235 = n_6222 ^ n_6223;
assign n_6236 = n_6223 ^ n_6194;
assign n_6237 = n_6226 ^ n_6227;
assign n_6238 = n_6227 ^ n_6199;
assign n_6239 = x64 & ~n_6228;
assign n_6240 = n_6207 & ~n_6229;
assign n_6241 = ~n_6208 & ~n_6230;
assign n_6242 = n_6211 & ~n_6231;
assign n_6243 = ~n_6212 & n_6232;
assign n_6244 = n_6233 ^ n_6168;
assign n_6245 = ~n_6234 ^ ~n_6159;
assign n_6246 = n_6220 & ~n_6235;
assign n_6247 = ~n_6221 & n_6236;
assign n_6248 = n_6224 & ~n_6237;
assign n_6249 = ~n_6225 & n_6238;
assign n_6250 = ~n_6165 & ~n_6239;
assign n_6251 = n_6241 ^ x100;
assign n_6252 = n_6243 ^ x93;
assign n_6253 = n_6244 ^ n_6114;
assign n_6254 = n_6247 ^ x95;
assign n_6255 = n_6249 ^ x102;
assign n_6256 = x66 ^ n_6250;
assign n_6257 = n_6253 ^ n_5890;
assign n_6258 = n_306 & ~n_6257;
assign n_6259 = n_6217 & ~n_6258;
assign n_6260 = ~n_6215 & n_6259;
assign n_6261 = ~n_6245 & ~n_6260;
assign n_6262 = x67 ^ n_6261;
assign n_6263 = n_6170 ^ n_6261;
assign n_6264 = n_6262 & n_6263;
assign n_6265 = n_6264 ^ x67;
assign n_6266 = n_6265 ^ x68;
assign n_6267 = n_6171 ^ n_6265;
assign n_6268 = n_6266 & n_6267;
assign n_6269 = n_6268 ^ x68;
assign n_6270 = n_6269 ^ x69;
assign n_6271 = n_6172 ^ n_6269;
assign n_6272 = n_6270 & n_6271;
assign n_6273 = n_6272 ^ x69;
assign n_6274 = n_6273 ^ x70;
assign n_6275 = n_6173 ^ n_6273;
assign n_6276 = n_6274 & n_6275;
assign n_6277 = n_6276 ^ x70;
assign n_6278 = n_6277 ^ x71;
assign n_6279 = n_6174 ^ n_6277;
assign n_6280 = n_6278 & n_6279;
assign n_6281 = n_6280 ^ x71;
assign n_6282 = n_6281 ^ x72;
assign n_6283 = n_6175 ^ n_6281;
assign n_6284 = n_6282 & n_6283;
assign n_6285 = n_6284 ^ x72;
assign n_6286 = n_6285 ^ x73;
assign n_6287 = n_6206 ^ n_6285;
assign n_6288 = n_6286 & n_6287;
assign n_6289 = n_6288 ^ x73;
assign n_6290 = n_6289 ^ x74;
assign n_6291 = n_6176 ^ n_6289;
assign n_6292 = n_6290 & n_6291;
assign n_6293 = n_6292 ^ x74;
assign n_6294 = n_6293 ^ x75;
assign n_6295 = n_6177 ^ n_6293;
assign n_6296 = n_6294 & ~n_6295;
assign n_6297 = n_6296 ^ x75;
assign n_6298 = n_6297 ^ x76;
assign n_6299 = n_6178 ^ n_6297;
assign n_6300 = n_6298 & n_6299;
assign n_6301 = n_6300 ^ x76;
assign n_6302 = n_6301 ^ x77;
assign n_6303 = n_6179 ^ n_6301;
assign n_6304 = n_6302 & n_6303;
assign n_6305 = n_6304 ^ x77;
assign n_6306 = n_6305 ^ x78;
assign n_6307 = n_6180 ^ n_6305;
assign n_6308 = n_6306 & n_6307;
assign n_6309 = n_6308 ^ x78;
assign n_6310 = n_6309 ^ x79;
assign n_6311 = n_6181 ^ n_6309;
assign n_6312 = n_6310 & n_6311;
assign n_6313 = n_6312 ^ x79;
assign n_6314 = n_6313 ^ x80;
assign n_6315 = n_6182 ^ n_6313;
assign n_6316 = n_6314 & n_6315;
assign n_6317 = n_6316 ^ x80;
assign n_6318 = n_6317 ^ x81;
assign n_6319 = n_6183 ^ n_6317;
assign n_6320 = n_6318 & n_6319;
assign n_6321 = n_6320 ^ x81;
assign n_6322 = n_6321 ^ x82;
assign n_6323 = n_6184 ^ n_6321;
assign n_6324 = n_6322 & n_6323;
assign n_6325 = n_6324 ^ x82;
assign n_6326 = n_6325 ^ x83;
assign n_6327 = n_6185 ^ n_6325;
assign n_6328 = n_6326 & n_6327;
assign n_6329 = n_6328 ^ x83;
assign n_6330 = n_6329 ^ x84;
assign n_6331 = n_6186 ^ n_6329;
assign n_6332 = n_6330 & n_6331;
assign n_6333 = n_6332 ^ x84;
assign n_6334 = n_6333 ^ x85;
assign n_6335 = n_6187 ^ n_6333;
assign n_6336 = n_6334 & n_6335;
assign n_6337 = n_6336 ^ x85;
assign n_6338 = n_6337 ^ x86;
assign n_6339 = n_6188 ^ n_6337;
assign n_6340 = n_6338 & n_6339;
assign n_6341 = n_6340 ^ x86;
assign n_6342 = n_6341 ^ x87;
assign n_6343 = n_6189 ^ n_6341;
assign n_6344 = n_6342 & n_6343;
assign n_6345 = n_6344 ^ x87;
assign n_6346 = n_6345 ^ x88;
assign n_6347 = n_6190 ^ n_6345;
assign n_6348 = n_6346 & n_6347;
assign n_6349 = n_6348 ^ x88;
assign n_6350 = n_6349 ^ x89;
assign n_6351 = n_6191 ^ n_6349;
assign n_6352 = n_6350 & n_6351;
assign n_6353 = n_6352 ^ x89;
assign n_6354 = n_6353 ^ x90;
assign n_6355 = n_6192 ^ n_6353;
assign n_6356 = n_6354 & n_6355;
assign n_6357 = n_6356 ^ x90;
assign n_6358 = n_6357 ^ x91;
assign n_6359 = n_6193 ^ n_6357;
assign n_6360 = n_6358 & n_6359;
assign n_6361 = n_6360 ^ x91;
assign n_6362 = n_6361 ^ x92;
assign n_6363 = n_6361 ^ n_6164;
assign n_6364 = n_6242 & n_6361;
assign n_6365 = n_6362 & n_6363;
assign n_6366 = ~n_6252 & ~n_6364;
assign n_6367 = n_6365 ^ x92;
assign n_6368 = x94 ^ n_6366;
assign n_6369 = n_6195 ^ n_6366;
assign n_6370 = n_6246 & ~n_6366;
assign n_6371 = n_6367 ^ x93;
assign n_6372 = ~n_6368 & ~n_6369;
assign n_6373 = ~n_6254 & ~n_6370;
assign n_6374 = n_6372 ^ x94;
assign n_6375 = x96 ^ n_6373;
assign n_6376 = n_6196 ^ n_6373;
assign n_6377 = n_6374 ^ x95;
assign n_6378 = ~n_6375 & ~n_6376;
assign n_6379 = n_6378 ^ x96;
assign n_6380 = n_6379 ^ x97;
assign n_6381 = n_6197 ^ n_6379;
assign n_6382 = n_6380 & n_6381;
assign n_6383 = n_6382 ^ x97;
assign n_6384 = n_6383 ^ x98;
assign n_6385 = n_6198 ^ n_6383;
assign n_6386 = n_6384 & n_6385;
assign n_6387 = n_6386 ^ x98;
assign n_6388 = n_6387 ^ x99;
assign n_6389 = n_6387 ^ n_6162;
assign n_6390 = n_6240 & ~n_6387;
assign n_6391 = n_6388 & n_6389;
assign n_6392 = n_6251 & ~n_6390;
assign n_6393 = n_6391 ^ x99;
assign n_6394 = x101 ^ n_6392;
assign n_6395 = n_6200 ^ n_6392;
assign n_6396 = n_6248 & n_6392;
assign n_6397 = n_6393 ^ x100;
assign n_6398 = n_6394 & n_6395;
assign n_6399 = ~n_6255 & ~n_6396;
assign n_6400 = n_6398 ^ x101;
assign n_6401 = x103 ^ n_6399;
assign n_6402 = n_6201 ^ n_6399;
assign n_6403 = n_6400 ^ x102;
assign n_6404 = ~n_6401 & ~n_6402;
assign n_6405 = n_6404 ^ x103;
assign n_6406 = n_6405 ^ x104;
assign n_6407 = n_6202 ^ n_6405;
assign n_6408 = n_6406 & n_6407;
assign n_6409 = n_6408 ^ x104;
assign n_6410 = n_6409 ^ x105;
assign n_6411 = n_6203 ^ n_6409;
assign n_6412 = n_6410 & n_6411;
assign n_6413 = n_6412 ^ x105;
assign n_6414 = n_6413 ^ x106;
assign n_6415 = n_6109 & ~n_6413;
assign n_6416 = n_6413 ^ ~n_5885;
assign n_6417 = n_6413 ^ n_6109;
assign n_6418 = ~n_6414 & ~n_6415;
assign n_6419 = n_6417 & n_6115;
assign n_6420 = n_365 & ~n_6418;
assign n_6421 = n_6419 ^ n_6113;
assign n_6422 = n_5885 & ~n_6420;
assign n_6423 = n_6421 ^ n_6109;
assign n_6424 = n_5941 ^ n_6422;
assign n_6425 = n_6423 ^ n_5927;
assign n_6426 = n_6416 & ~n_6425;
assign n_6427 = n_6413 ^ n_6426;
assign n_6428 = n_365 & ~n_6427;
assign n_6429 = n_6406 & n_6428;
assign n_6430 = ~n_6401 & n_6428;
assign n_6431 = n_6394 & n_6428;
assign n_6432 = n_6384 & n_6428;
assign n_6433 = n_6380 & n_6428;
assign n_6434 = n_6318 & n_6428;
assign n_6435 = n_6314 & n_6428;
assign n_6436 = n_6274 & n_6428;
assign n_6437 = n_6270 & n_6428;
assign n_6438 = ~x64 & n_6428;
assign n_6439 = n_6262 & n_6428;
assign n_6440 = n_6266 & n_6428;
assign n_6441 = n_6278 & n_6428;
assign n_6442 = n_6282 & n_6428;
assign n_6443 = n_6286 & n_6428;
assign n_6444 = n_6290 & n_6428;
assign n_6445 = n_6294 & n_6428;
assign n_6446 = n_6298 & n_6428;
assign n_6447 = n_6302 & n_6428;
assign n_6448 = n_6306 & n_6428;
assign n_6449 = n_6310 & n_6428;
assign n_6450 = n_6322 & n_6428;
assign n_6451 = n_6326 & n_6428;
assign n_6452 = n_6330 & n_6428;
assign n_6453 = n_6334 & n_6428;
assign n_6454 = n_6338 & n_6428;
assign n_6455 = n_6342 & n_6428;
assign n_6456 = n_6346 & n_6428;
assign n_6457 = n_6350 & n_6428;
assign n_6458 = n_6354 & n_6428;
assign n_6459 = n_6358 & n_6428;
assign n_6460 = n_6362 & n_6428;
assign n_6461 = ~n_6368 & n_6428;
assign n_6462 = ~n_6375 & n_6428;
assign n_6463 = n_6388 & n_6428;
assign n_6464 = n_6410 & n_6428;
assign y21 = n_6428;
assign n_6465 = n_6403 & n_6428;
assign n_6466 = ~n_6256 & n_6428;
assign n_6467 = n_6371 & n_6428;
assign n_6468 = n_6377 & n_6428;
assign n_6469 = n_6397 & n_6428;
assign n_6470 = n_6429 ^ n_6202;
assign n_6471 = n_6430 ^ n_6201;
assign n_6472 = n_6431 ^ n_6200;
assign n_6473 = n_6432 ^ n_6198;
assign n_6474 = n_6433 ^ n_6197;
assign n_6475 = n_6434 ^ n_6183;
assign n_6476 = n_6435 ^ n_6182;
assign n_6477 = n_6436 ^ n_6173;
assign n_6478 = n_6437 ^ n_6172;
assign n_6479 = n_6438 ^ n_6428;
assign n_6480 = x65 & n_6438;
assign n_6481 = n_6439 ^ n_6170;
assign n_6482 = n_6440 ^ n_6171;
assign n_6483 = n_6441 ^ n_6174;
assign n_6484 = n_6442 ^ n_6175;
assign n_6485 = n_6443 ^ n_6206;
assign n_6486 = n_6444 ^ n_6176;
assign n_6487 = n_6445 ^ n_6177;
assign n_6488 = n_6446 ^ n_6178;
assign n_6489 = n_6447 ^ n_6179;
assign n_6490 = n_6448 ^ n_6180;
assign n_6491 = n_6449 ^ n_6181;
assign n_6492 = n_6450 ^ n_6184;
assign n_6493 = n_6451 ^ n_6185;
assign n_6494 = n_6452 ^ n_6186;
assign n_6495 = n_6453 ^ n_6187;
assign n_6496 = n_6454 ^ n_6188;
assign n_6497 = n_6455 ^ n_6189;
assign n_6498 = n_6456 ^ n_6190;
assign n_6499 = n_6457 ^ n_6191;
assign n_6500 = n_6458 ^ n_6192;
assign n_6501 = n_6459 ^ n_6193;
assign n_6502 = n_6460 ^ n_6164;
assign n_6503 = n_6461 ^ n_6195;
assign n_6504 = n_6462 ^ n_6196;
assign n_6505 = n_6463 ^ n_6162;
assign n_6506 = n_6464 ^ n_6203;
assign n_6507 = n_6199 ^ n_6465;
assign n_6508 = n_6204 ^ n_6466;
assign n_6509 = n_6163 ^ n_6467;
assign n_6510 = n_6194 ^ n_6468;
assign n_6511 = n_6161 ^ n_6469;
assign n_6512 = n_6470 ^ x105;
assign n_6513 = n_6471 ^ x104;
assign n_6514 = n_6472 ^ x102;
assign n_6515 = ~x99 ^ n_6473;
assign n_6516 = n_6473 ^ x99;
assign n_6517 = n_6474 ^ x98;
assign n_6518 = x98 & ~n_6474;
assign n_6519 = ~x82 ^ n_6475;
assign n_6520 = n_6475 ^ x82;
assign n_6521 = n_6476 ^ x81;
assign n_6522 = x81 & ~n_6476;
assign n_6523 = n_6477 ^ x71;
assign n_6524 = n_6478 ^ x70;
assign n_6525 = n_6479 ^ x21;
assign n_6526 = ~n_84 & n_6479;
assign n_6527 = n_6507 ^ x103;
assign n_6528 = n_6517 ^ n_6518;
assign n_6529 = n_6518 ^ n_6473;
assign n_6530 = n_6521 ^ n_6522;
assign n_6531 = n_6522 ^ n_6475;
assign n_6532 = n_6525 ^ x65;
assign n_6533 = n_25 ^ n_6525;
assign n_6534 = n_6525 & ~n_86;
assign n_6535 = n_6526 ^ n_6480;
assign n_6536 = n_6515 & ~n_6528;
assign n_6537 = ~n_6516 & n_6529;
assign n_6538 = n_6519 & ~n_6530;
assign n_6539 = ~n_6520 & n_6531;
assign n_6540 = ~n_6532 ^ ~n_218;
assign n_6541 = ~n_6532 & n_219;
assign n_6542 = ~n_6532 & n_6533;
assign n_6543 = n_6535 ^ n_6120;
assign n_6544 = n_6537 ^ x99;
assign n_6545 = n_6539 ^ x82;
assign n_6546 = n_6542 ^ x65;
assign n_6547 = n_6543 ^ x22;
assign n_6548 = n_6546 ^ x66;
assign n_6549 = n_6547 ^ n_6546;
assign n_6550 = n_6548 & n_6549;
assign n_6551 = n_6550 ^ x66;
assign n_6552 = n_6551 ^ x67;
assign n_6553 = n_6508 ^ n_6551;
assign n_6554 = n_6552 & n_6553;
assign n_6555 = n_6554 ^ x67;
assign n_6556 = n_6555 ^ x68;
assign n_6557 = n_6481 ^ n_6555;
assign n_6558 = n_6556 & n_6557;
assign n_6559 = n_6558 ^ x68;
assign n_6560 = n_6559 ^ x69;
assign n_6561 = n_6482 ^ n_6559;
assign n_6562 = n_6560 & n_6561;
assign n_6563 = n_6562 ^ x69;
assign n_6564 = n_6563 ^ n_6478;
assign n_6565 = n_6563 ^ x70;
assign n_6566 = ~n_6524 & n_6564;
assign n_6567 = n_6566 ^ x70;
assign n_6568 = n_6567 ^ n_6477;
assign n_6569 = n_6567 ^ x71;
assign n_6570 = ~n_6523 & n_6568;
assign n_6571 = n_6570 ^ x71;
assign n_6572 = n_6571 ^ x72;
assign n_6573 = n_6483 ^ n_6571;
assign n_6574 = n_6572 & n_6573;
assign n_6575 = n_6574 ^ x72;
assign n_6576 = n_6575 ^ x73;
assign n_6577 = n_6484 ^ n_6575;
assign n_6578 = n_6576 & n_6577;
assign n_6579 = n_6578 ^ x73;
assign n_6580 = n_6579 ^ x74;
assign n_6581 = n_6485 ^ n_6579;
assign n_6582 = n_6580 & n_6581;
assign n_6583 = n_6582 ^ x74;
assign n_6584 = n_6583 ^ x75;
assign n_6585 = n_6486 ^ n_6583;
assign n_6586 = n_6584 & n_6585;
assign n_6587 = n_6586 ^ x75;
assign n_6588 = n_6587 ^ x76;
assign n_6589 = n_6487 ^ n_6587;
assign n_6590 = n_6588 & ~n_6589;
assign n_6591 = n_6590 ^ x76;
assign n_6592 = n_6591 ^ x77;
assign n_6593 = n_6488 ^ n_6591;
assign n_6594 = n_6592 & n_6593;
assign n_6595 = n_6594 ^ x77;
assign n_6596 = n_6595 ^ x78;
assign n_6597 = n_6489 ^ n_6595;
assign n_6598 = n_6596 & n_6597;
assign n_6599 = n_6598 ^ x78;
assign n_6600 = n_6599 ^ x79;
assign n_6601 = n_6490 ^ n_6599;
assign n_6602 = n_6600 & n_6601;
assign n_6603 = n_6602 ^ x79;
assign n_6604 = n_6603 ^ x80;
assign n_6605 = n_6491 ^ n_6603;
assign n_6606 = n_6604 & n_6605;
assign n_6607 = n_6606 ^ x80;
assign n_6608 = n_6607 ^ x81;
assign n_6609 = n_6607 ^ n_6476;
assign n_6610 = n_6538 & n_6607;
assign n_6611 = n_6608 & n_6609;
assign n_6612 = ~n_6545 & ~n_6610;
assign n_6613 = n_6611 ^ x81;
assign n_6614 = x83 ^ n_6612;
assign n_6615 = n_6492 ^ n_6612;
assign n_6616 = n_6613 ^ x82;
assign n_6617 = ~n_6614 & ~n_6615;
assign n_6618 = n_6617 ^ x83;
assign n_6619 = n_6618 ^ x84;
assign n_6620 = n_6493 ^ n_6618;
assign n_6621 = n_6619 & n_6620;
assign n_6622 = n_6621 ^ x84;
assign n_6623 = n_6622 ^ x85;
assign n_6624 = n_6494 ^ n_6622;
assign n_6625 = n_6623 & n_6624;
assign n_6626 = n_6625 ^ x85;
assign n_6627 = n_6626 ^ x86;
assign n_6628 = n_6495 ^ n_6626;
assign n_6629 = n_6627 & n_6628;
assign n_6630 = n_6629 ^ x86;
assign n_6631 = n_6630 ^ x87;
assign n_6632 = n_6496 ^ n_6630;
assign n_6633 = n_6631 & n_6632;
assign n_6634 = n_6633 ^ x87;
assign n_6635 = n_6634 ^ x88;
assign n_6636 = n_6497 ^ n_6634;
assign n_6637 = n_6635 & n_6636;
assign n_6638 = n_6637 ^ x88;
assign n_6639 = n_6638 ^ x89;
assign n_6640 = n_6498 ^ n_6638;
assign n_6641 = n_6639 & n_6640;
assign n_6642 = n_6641 ^ x89;
assign n_6643 = n_6642 ^ x90;
assign n_6644 = n_6499 ^ n_6642;
assign n_6645 = n_6643 & n_6644;
assign n_6646 = n_6645 ^ x90;
assign n_6647 = n_6646 ^ x91;
assign n_6648 = n_6500 ^ n_6646;
assign n_6649 = n_6647 & n_6648;
assign n_6650 = n_6649 ^ x91;
assign n_6651 = n_6650 ^ x92;
assign n_6652 = n_6501 ^ n_6650;
assign n_6653 = n_6651 & n_6652;
assign n_6654 = n_6653 ^ x92;
assign n_6655 = n_6654 ^ x93;
assign n_6656 = n_6502 ^ n_6654;
assign n_6657 = n_6655 & n_6656;
assign n_6658 = n_6657 ^ x93;
assign n_6659 = n_6658 ^ x94;
assign n_6660 = n_6509 ^ n_6658;
assign n_6661 = n_6659 & n_6660;
assign n_6662 = n_6661 ^ x94;
assign n_6663 = n_6662 ^ x95;
assign n_6664 = n_6503 ^ n_6662;
assign n_6665 = n_6663 & n_6664;
assign n_6666 = n_6665 ^ x95;
assign n_6667 = n_6666 ^ x96;
assign n_6668 = n_6510 ^ n_6666;
assign n_6669 = n_6667 & n_6668;
assign n_6670 = n_6669 ^ x96;
assign n_6671 = n_6670 ^ x97;
assign n_6672 = n_6504 ^ n_6670;
assign n_6673 = n_6671 & n_6672;
assign n_6674 = n_6673 ^ x97;
assign n_6675 = n_6674 ^ x98;
assign n_6676 = n_6674 ^ n_6474;
assign n_6677 = n_6536 & n_6674;
assign n_6678 = n_6675 & n_6676;
assign n_6679 = ~n_6544 & ~n_6677;
assign n_6680 = n_6678 ^ x98;
assign n_6681 = x100 ^ n_6679;
assign n_6682 = n_6505 ^ n_6679;
assign n_6683 = n_6680 ^ x99;
assign n_6684 = ~n_6681 & ~n_6682;
assign n_6685 = n_6684 ^ x100;
assign n_6686 = n_6685 ^ x101;
assign n_6687 = n_6511 ^ n_6685;
assign n_6688 = n_6686 & n_6687;
assign n_6689 = n_6688 ^ x101;
assign n_6690 = n_6689 ^ n_6472;
assign n_6691 = n_6689 ^ x102;
assign n_6692 = ~n_6514 & n_6690;
assign n_6693 = n_6692 ^ x102;
assign n_6694 = n_6693 ^ n_6507;
assign n_6695 = n_6693 ^ x103;
assign n_6696 = ~n_6527 & n_6694;
assign n_6697 = n_6696 ^ x103;
assign n_6698 = n_6697 ^ n_6471;
assign n_6699 = n_6697 ^ x104;
assign n_6700 = ~n_6513 & n_6698;
assign n_6701 = n_6700 ^ x104;
assign n_6702 = n_6701 ^ n_6470;
assign n_6703 = n_6701 ^ x105;
assign n_6704 = ~n_6512 & n_6702;
assign n_6705 = n_6704 ^ x105;
assign n_6706 = n_6705 ^ x106;
assign n_6707 = n_6506 ^ n_6705;
assign n_6708 = n_6706 & n_6707;
assign n_6709 = n_6708 ^ x106;
assign n_6710 = n_6709 & ~n_6424;
assign n_6711 = n_6709 ^ x107;
assign n_6712 = ~n_6710 & n_5942;
assign n_6713 = ~x108 & ~n_6711;
assign n_6714 = n_6706 & n_6712;
assign n_6715 = x64 & n_6712;
assign n_6716 = n_6525 ^ n_6712;
assign n_6717 = x20 & n_6712;
assign n_6718 = x20 ^ n_6712;
assign n_6719 = x19 ^ n_6712;
assign n_6720 = n_26 ^ n_6712;
assign n_6721 = n_6548 & n_6712;
assign n_6722 = n_6552 & n_6712;
assign n_6723 = n_6556 & n_6712;
assign n_6724 = n_6560 & n_6712;
assign n_6725 = n_6565 & n_6712;
assign n_6726 = n_6569 & n_6712;
assign n_6727 = n_6572 & n_6712;
assign n_6728 = n_6576 & n_6712;
assign n_6729 = n_6580 & n_6712;
assign n_6730 = n_6584 & n_6712;
assign n_6731 = n_6588 & n_6712;
assign n_6732 = n_6592 & n_6712;
assign n_6733 = n_6596 & n_6712;
assign n_6734 = n_6600 & n_6712;
assign n_6735 = n_6604 & n_6712;
assign n_6736 = n_6608 & n_6712;
assign n_6737 = ~n_6614 & n_6712;
assign n_6738 = n_6619 & n_6712;
assign n_6739 = n_6623 & n_6712;
assign n_6740 = n_6627 & n_6712;
assign n_6741 = n_6631 & n_6712;
assign n_6742 = n_6635 & n_6712;
assign n_6743 = n_6639 & n_6712;
assign n_6744 = n_6643 & n_6712;
assign n_6745 = n_6647 & n_6712;
assign n_6746 = n_6651 & n_6712;
assign n_6747 = n_6655 & n_6712;
assign n_6748 = n_6659 & n_6712;
assign n_6749 = n_6663 & n_6712;
assign n_6750 = n_6667 & n_6712;
assign n_6751 = n_6671 & n_6712;
assign n_6752 = n_6675 & n_6712;
assign n_6753 = ~n_6681 & n_6712;
assign n_6754 = n_6686 & n_6712;
assign n_6755 = n_6691 & n_6712;
assign n_6756 = n_6695 & n_6712;
assign n_6757 = n_6699 & n_6712;
assign n_6758 = n_6703 & n_6712;
assign n_6759 = n_159 & n_6712;
assign y20 = n_6712;
assign n_6760 = n_6616 & n_6712;
assign n_6761 = n_6683 & n_6712;
assign n_6762 = n_6713 ^ x108;
assign n_6763 = n_6713 & ~n_6420;
assign n_6764 = n_6714 ^ n_6506;
assign n_6765 = ~n_6715 & n_86;
assign n_6766 = n_6715 & n_6541;
assign n_6767 = n_6717 & ~n_218;
assign n_6768 = n_6717 & n_188;
assign n_6769 = n_6719 & ~n_6712;
assign n_6770 = n_6720 & n_253;
assign n_6771 = n_6721 ^ n_6547;
assign n_6772 = n_6722 ^ n_6508;
assign n_6773 = n_6723 ^ n_6481;
assign n_6774 = n_6724 ^ n_6482;
assign n_6775 = n_6725 ^ n_6478;
assign n_6776 = n_6726 ^ n_6477;
assign n_6777 = n_6727 ^ n_6483;
assign n_6778 = n_6728 ^ n_6484;
assign n_6779 = n_6729 ^ n_6485;
assign n_6780 = n_6730 ^ n_6486;
assign n_6781 = n_6731 ^ n_6487;
assign n_6782 = n_6732 ^ n_6488;
assign n_6783 = n_6733 ^ n_6489;
assign n_6784 = n_6734 ^ n_6490;
assign n_6785 = n_6735 ^ n_6491;
assign n_6786 = n_6736 ^ n_6476;
assign n_6787 = n_6737 ^ n_6492;
assign n_6788 = n_6738 ^ n_6493;
assign n_6789 = n_6739 ^ n_6494;
assign n_6790 = n_6740 ^ n_6495;
assign n_6791 = n_6741 ^ n_6496;
assign n_6792 = n_6742 ^ n_6497;
assign n_6793 = n_6743 ^ n_6498;
assign n_6794 = n_6744 ^ n_6499;
assign n_6795 = n_6745 ^ n_6500;
assign n_6796 = n_6746 ^ n_6501;
assign n_6797 = n_6747 ^ n_6502;
assign n_6798 = n_6748 ^ n_6509;
assign n_6799 = n_6749 ^ n_6503;
assign n_6800 = n_6750 ^ n_6510;
assign n_6801 = n_6751 ^ n_6504;
assign n_6802 = n_6752 ^ n_6474;
assign n_6803 = n_6753 ^ n_6505;
assign n_6804 = n_6754 ^ n_6511;
assign n_6805 = n_6755 ^ n_6472;
assign n_6806 = n_6756 ^ n_6507;
assign n_6807 = n_6757 ^ n_6471;
assign n_6808 = n_6758 ^ n_6470;
assign n_6809 = n_6759 ^ n_6525;
assign n_6810 = n_6475 ^ n_6760;
assign n_6811 = n_6473 ^ n_6761;
assign n_6812 = ~x107 & n_6764;
assign n_6813 = n_6764 ^ x107;
assign n_6814 = n_6765 & ~n_6716;
assign n_6815 = ~n_6768 ^ ~n_6766;
assign n_6816 = n_6769 ^ n_6712;
assign n_6817 = n_6770 ^ n_6712;
assign n_6818 = ~n_6812 ^ ~n_6763;
assign n_6819 = n_6813 ^ n_6812;
assign n_6820 = ~x66 & ~n_6814;
assign n_6821 = n_6718 & ~n_6816;
assign n_6822 = n_6534 & ~n_6817;
assign n_6823 = n_6821 ^ n_6769;
assign n_6824 = ~n_6815 ^ ~n_6822;
assign n_6825 = n_6823 ^ n_6712;
assign n_6826 = n_6825 ^ x19;
assign n_6827 = ~x65 & n_6826;
assign n_6828 = x19 ^ n_6827;
assign n_6829 = ~n_6525 & ~n_6828;
assign n_6830 = n_6828 & ~n_6767;
assign n_6831 = ~n_6540 ^ n_6829;
assign n_6832 = x64 & ~n_6830;
assign n_6833 = n_6717 & n_6831;
assign n_6834 = ~n_6765 & ~n_6832;
assign n_6835 = n_6833 ^ n_6829;
assign n_6836 = x66 ^ n_6834;
assign n_6837 = x64 & n_6835;
assign n_6838 = n_6820 & ~n_6837;
assign n_6839 = ~n_6824 & ~n_6838;
assign n_6840 = x67 ^ n_6839;
assign n_6841 = n_6771 ^ n_6839;
assign n_6842 = n_6840 & n_6841;
assign n_6843 = n_6842 ^ x67;
assign n_6844 = n_6843 ^ x68;
assign n_6845 = n_6772 ^ n_6843;
assign n_6846 = n_6844 & n_6845;
assign n_6847 = n_6846 ^ x68;
assign n_6848 = n_6847 ^ x69;
assign n_6849 = n_6773 ^ n_6847;
assign n_6850 = n_6848 & n_6849;
assign n_6851 = n_6850 ^ x69;
assign n_6852 = n_6851 ^ x70;
assign n_6853 = n_6774 ^ n_6851;
assign n_6854 = n_6852 & n_6853;
assign n_6855 = n_6854 ^ x70;
assign n_6856 = n_6855 ^ x71;
assign n_6857 = n_6775 ^ n_6855;
assign n_6858 = n_6856 & n_6857;
assign n_6859 = n_6858 ^ x71;
assign n_6860 = n_6859 ^ x72;
assign n_6861 = n_6776 ^ n_6859;
assign n_6862 = n_6860 & n_6861;
assign n_6863 = n_6862 ^ x72;
assign n_6864 = n_6863 ^ x73;
assign n_6865 = n_6777 ^ n_6863;
assign n_6866 = n_6864 & n_6865;
assign n_6867 = n_6866 ^ x73;
assign n_6868 = n_6867 ^ x74;
assign n_6869 = n_6778 ^ n_6867;
assign n_6870 = n_6868 & n_6869;
assign n_6871 = n_6870 ^ x74;
assign n_6872 = n_6871 ^ x75;
assign n_6873 = n_6779 ^ n_6871;
assign n_6874 = n_6872 & n_6873;
assign n_6875 = n_6874 ^ x75;
assign n_6876 = n_6875 ^ x76;
assign n_6877 = n_6780 ^ n_6875;
assign n_6878 = n_6876 & n_6877;
assign n_6879 = n_6878 ^ x76;
assign n_6880 = n_6879 ^ x77;
assign n_6881 = n_6781 ^ n_6879;
assign n_6882 = n_6880 & ~n_6881;
assign n_6883 = n_6882 ^ x77;
assign n_6884 = n_6883 ^ x78;
assign n_6885 = n_6782 ^ n_6883;
assign n_6886 = n_6884 & n_6885;
assign n_6887 = n_6886 ^ x78;
assign n_6888 = n_6887 ^ x79;
assign n_6889 = n_6783 ^ n_6887;
assign n_6890 = n_6888 & n_6889;
assign n_6891 = n_6890 ^ x79;
assign n_6892 = n_6891 ^ x80;
assign n_6893 = n_6784 ^ n_6891;
assign n_6894 = n_6892 & n_6893;
assign n_6895 = n_6894 ^ x80;
assign n_6896 = n_6895 ^ x81;
assign n_6897 = n_6785 ^ n_6895;
assign n_6898 = n_6896 & n_6897;
assign n_6899 = n_6898 ^ x81;
assign n_6900 = n_6899 ^ x82;
assign n_6901 = n_6786 ^ n_6899;
assign n_6902 = n_6900 & n_6901;
assign n_6903 = n_6902 ^ x82;
assign n_6904 = n_6903 ^ x83;
assign n_6905 = n_6810 ^ n_6903;
assign n_6906 = n_6904 & n_6905;
assign n_6907 = n_6906 ^ x83;
assign n_6908 = n_6907 ^ x84;
assign n_6909 = n_6787 ^ n_6907;
assign n_6910 = n_6908 & n_6909;
assign n_6911 = n_6910 ^ x84;
assign n_6912 = n_6911 ^ x85;
assign n_6913 = n_6788 ^ n_6911;
assign n_6914 = n_6912 & n_6913;
assign n_6915 = n_6914 ^ x85;
assign n_6916 = n_6915 ^ x86;
assign n_6917 = n_6789 ^ n_6915;
assign n_6918 = n_6916 & n_6917;
assign n_6919 = n_6918 ^ x86;
assign n_6920 = n_6919 ^ x87;
assign n_6921 = n_6790 ^ n_6919;
assign n_6922 = n_6920 & n_6921;
assign n_6923 = n_6922 ^ x87;
assign n_6924 = n_6923 ^ x88;
assign n_6925 = n_6791 ^ n_6923;
assign n_6926 = n_6924 & n_6925;
assign n_6927 = n_6926 ^ x88;
assign n_6928 = n_6927 ^ x89;
assign n_6929 = n_6792 ^ n_6927;
assign n_6930 = n_6928 & n_6929;
assign n_6931 = n_6930 ^ x89;
assign n_6932 = n_6931 ^ x90;
assign n_6933 = n_6793 ^ n_6931;
assign n_6934 = n_6932 & n_6933;
assign n_6935 = n_6934 ^ x90;
assign n_6936 = n_6935 ^ x91;
assign n_6937 = n_6794 ^ n_6935;
assign n_6938 = n_6936 & n_6937;
assign n_6939 = n_6938 ^ x91;
assign n_6940 = n_6939 ^ x92;
assign n_6941 = n_6795 ^ n_6939;
assign n_6942 = n_6940 & n_6941;
assign n_6943 = n_6942 ^ x92;
assign n_6944 = n_6943 ^ x93;
assign n_6945 = n_6796 ^ n_6943;
assign n_6946 = n_6944 & n_6945;
assign n_6947 = n_6946 ^ x93;
assign n_6948 = n_6947 ^ x94;
assign n_6949 = n_6797 ^ n_6947;
assign n_6950 = n_6948 & n_6949;
assign n_6951 = n_6950 ^ x94;
assign n_6952 = n_6951 ^ x95;
assign n_6953 = n_6798 ^ n_6951;
assign n_6954 = n_6952 & n_6953;
assign n_6955 = n_6954 ^ x95;
assign n_6956 = n_6955 ^ x96;
assign n_6957 = n_6799 ^ n_6955;
assign n_6958 = n_6956 & n_6957;
assign n_6959 = n_6958 ^ x96;
assign n_6960 = n_6959 ^ x97;
assign n_6961 = n_6800 ^ n_6959;
assign n_6962 = n_6960 & n_6961;
assign n_6963 = n_6962 ^ x97;
assign n_6964 = n_6963 ^ x98;
assign n_6965 = n_6801 ^ n_6963;
assign n_6966 = n_6964 & n_6965;
assign n_6967 = n_6966 ^ x98;
assign n_6968 = n_6967 ^ x99;
assign n_6969 = n_6802 ^ n_6967;
assign n_6970 = n_6968 & n_6969;
assign n_6971 = n_6970 ^ x99;
assign n_6972 = n_6971 ^ x100;
assign n_6973 = n_6811 ^ n_6971;
assign n_6974 = n_6972 & n_6973;
assign n_6975 = n_6974 ^ x100;
assign n_6976 = n_6975 ^ x101;
assign n_6977 = n_6803 ^ n_6975;
assign n_6978 = n_6976 & n_6977;
assign n_6979 = n_6978 ^ x101;
assign n_6980 = n_6979 ^ x102;
assign n_6981 = n_6804 ^ n_6979;
assign n_6982 = n_6980 & n_6981;
assign n_6983 = n_6982 ^ x102;
assign n_6984 = n_6983 ^ x103;
assign n_6985 = n_6805 ^ n_6983;
assign n_6986 = n_6984 & n_6985;
assign n_6987 = n_6986 ^ x103;
assign n_6988 = n_6987 ^ x104;
assign n_6989 = n_6806 ^ n_6987;
assign n_6990 = n_6988 & n_6989;
assign n_6991 = n_6990 ^ x104;
assign n_6992 = n_6991 ^ x105;
assign n_6993 = n_6807 ^ n_6991;
assign n_6994 = n_6992 & n_6993;
assign n_6995 = n_6994 ^ x105;
assign n_6996 = n_6995 ^ x106;
assign n_6997 = n_6808 ^ n_6995;
assign n_6998 = n_6996 & n_6997;
assign n_6999 = n_6998 ^ x106;
assign n_7000 = ~n_6999 & ~n_6819;
assign n_7001 = n_6999 ^ x107;
assign n_7002 = ~n_6812 & ~n_7000;
assign n_7003 = ~n_7000 & ~n_6818;
assign n_7004 = ~n_7002 & n_6762;
assign n_7005 = n_362 & ~n_7002;
assign n_7006 = n_5929 & ~n_7003;
assign n_7007 = n_7004 ^ x108;
assign n_7008 = ~n_7005 & ~n_7006;
assign n_7009 = n_361 & ~n_7007;
assign n_7010 = n_6996 & ~n_7008;
assign n_7011 = n_6992 & ~n_7008;
assign n_7012 = n_6960 & ~n_7008;
assign n_7013 = n_6956 & ~n_7008;
assign n_7014 = n_6892 & ~n_7008;
assign n_7015 = n_6888 & ~n_7008;
assign n_7016 = n_265 & ~n_7008;
assign n_7017 = x64 & ~n_7008;
assign n_7018 = n_6840 & ~n_7008;
assign n_7019 = n_6844 & ~n_7008;
assign n_7020 = n_6848 & ~n_7008;
assign n_7021 = n_6852 & ~n_7008;
assign n_7022 = n_6856 & ~n_7008;
assign n_7023 = n_6860 & ~n_7008;
assign n_7024 = n_6864 & ~n_7008;
assign n_7025 = n_6868 & ~n_7008;
assign n_7026 = n_6872 & ~n_7008;
assign n_7027 = n_6876 & ~n_7008;
assign n_7028 = n_6880 & ~n_7008;
assign n_7029 = n_6884 & ~n_7008;
assign n_7030 = n_6896 & ~n_7008;
assign n_7031 = n_6900 & ~n_7008;
assign n_7032 = n_6904 & ~n_7008;
assign n_7033 = n_6908 & ~n_7008;
assign n_7034 = n_6912 & ~n_7008;
assign n_7035 = n_6916 & ~n_7008;
assign n_7036 = n_6920 & ~n_7008;
assign n_7037 = n_6924 & ~n_7008;
assign n_7038 = n_6928 & ~n_7008;
assign n_7039 = n_6932 & ~n_7008;
assign n_7040 = n_6936 & ~n_7008;
assign n_7041 = n_6940 & ~n_7008;
assign n_7042 = n_6944 & ~n_7008;
assign n_7043 = n_6948 & ~n_7008;
assign n_7044 = n_6952 & ~n_7008;
assign n_7045 = n_6968 & ~n_7008;
assign n_7046 = n_6964 & ~n_7008;
assign n_7047 = n_6972 & ~n_7008;
assign n_7048 = n_6976 & ~n_7008;
assign n_7049 = n_6980 & ~n_7008;
assign n_7050 = n_6984 & ~n_7008;
assign n_7051 = n_6988 & ~n_7008;
assign n_7052 = n_7001 & ~n_7008;
assign y19 = ~n_7008;
assign n_7053 = n_254 & n_7008;
assign n_7054 = ~n_6836 & ~n_7008;
assign n_7055 = n_6422 & ~n_7009;
assign n_7056 = n_7010 ^ n_6808;
assign n_7057 = n_7011 ^ n_6807;
assign n_7058 = n_7012 ^ n_6800;
assign n_7059 = n_7013 ^ n_6799;
assign n_7060 = n_7014 ^ n_6784;
assign n_7061 = n_7015 ^ n_6783;
assign n_7062 = n_7016 ^ n_6715;
assign n_7063 = n_7017 & n_307;
assign n_7064 = n_7018 ^ n_6771;
assign n_7065 = n_7019 ^ n_6772;
assign n_7066 = n_7020 ^ n_6773;
assign n_7067 = n_7021 ^ n_6774;
assign n_7068 = n_7022 ^ n_6775;
assign n_7069 = n_7023 ^ n_6776;
assign n_7070 = n_7024 ^ n_6777;
assign n_7071 = n_7025 ^ n_6778;
assign n_7072 = n_7026 ^ n_6779;
assign n_7073 = n_7027 ^ n_6780;
assign n_7074 = n_7028 ^ n_6781;
assign n_7075 = n_7029 ^ n_6782;
assign n_7076 = n_7030 ^ n_6785;
assign n_7077 = n_7031 ^ n_6786;
assign n_7078 = n_7032 ^ n_6810;
assign n_7079 = n_7033 ^ n_6787;
assign n_7080 = n_7034 ^ n_6788;
assign n_7081 = n_7035 ^ n_6789;
assign n_7082 = n_7036 ^ n_6790;
assign n_7083 = n_7037 ^ n_6791;
assign n_7084 = n_7038 ^ n_6792;
assign n_7085 = n_7039 ^ n_6793;
assign n_7086 = n_7040 ^ n_6794;
assign n_7087 = n_7041 ^ n_6795;
assign n_7088 = n_7042 ^ n_6796;
assign n_7089 = n_7043 ^ n_6797;
assign n_7090 = n_7044 ^ n_6798;
assign n_7091 = n_7045 ^ n_6802;
assign n_7092 = n_7046 ^ n_6801;
assign n_7093 = n_7047 ^ n_6811;
assign n_7094 = n_7048 ^ n_6803;
assign n_7095 = n_7049 ^ n_6804;
assign n_7096 = n_7050 ^ n_6805;
assign n_7097 = n_7051 ^ n_6806;
assign n_7098 = n_7052 ^ n_6764;
assign n_7099 = ~n_308 & ~n_7053;
assign n_7100 = n_6809 ^ n_7054;
assign n_7101 = ~x109 ^ n_7055;
assign n_7102 = ~x107 ^ n_7056;
assign n_7103 = n_7056 ^ x107;
assign n_7104 = n_7057 ^ x106;
assign n_7105 = x106 & ~n_7057;
assign n_7106 = x98 ^ ~n_7058;
assign n_7107 = n_7058 ^ x98;
assign n_7108 = n_7059 ^ x97;
assign n_7109 = ~x97 & n_7059;
assign n_7110 = x81 ^ ~n_7060;
assign n_7111 = n_7060 ^ x81;
assign n_7112 = n_7061 ^ x80;
assign n_7113 = ~x80 & n_7061;
assign n_7114 = n_7062 ^ x20;
assign n_7115 = ~x100 ^ n_7091;
assign n_7116 = n_7091 ^ x100;
assign n_7117 = n_7092 ^ x99;
assign n_7118 = x99 & ~n_7092;
assign n_7119 = ~n_7063 & n_7099;
assign n_7120 = n_7104 ^ n_7105;
assign n_7121 = n_7105 ^ n_7056;
assign n_7122 = n_7108 ^ n_7109;
assign n_7123 = n_7109 ^ n_7058;
assign n_7124 = n_7112 ^ n_7113;
assign n_7125 = n_7113 ^ n_7060;
assign n_7126 = n_7114 ^ x66;
assign n_7127 = n_7117 ^ n_7118;
assign n_7128 = n_7118 ^ n_7091;
assign n_7129 = n_7114 ^ n_7119;
assign n_7130 = x66 ^ n_7119;
assign n_7131 = n_7102 & ~n_7120;
assign n_7132 = ~n_7103 & n_7121;
assign n_7133 = n_7106 & ~n_7122;
assign n_7134 = ~n_7107 & ~n_7123;
assign n_7135 = n_7110 & ~n_7124;
assign n_7136 = ~n_7111 & ~n_7125;
assign n_7137 = n_7115 & ~n_7127;
assign n_7138 = ~n_7116 & n_7128;
assign n_7139 = ~n_7126 & ~n_7129;
assign n_7140 = n_7132 ^ x107;
assign n_7141 = n_7134 ^ x98;
assign n_7142 = n_7136 ^ x81;
assign n_7143 = n_7138 ^ x100;
assign n_7144 = n_7139 ^ x66;
assign n_7145 = n_7144 ^ x67;
assign n_7146 = n_7100 ^ n_7144;
assign n_7147 = n_7145 & n_7146;
assign n_7148 = n_7147 ^ x67;
assign n_7149 = n_7148 ^ x68;
assign n_7150 = n_7064 ^ n_7148;
assign n_7151 = n_7149 & n_7150;
assign n_7152 = n_7151 ^ x68;
assign n_7153 = n_7152 ^ x69;
assign n_7154 = n_7065 ^ n_7152;
assign n_7155 = n_7153 & n_7154;
assign n_7156 = n_7155 ^ x69;
assign n_7157 = n_7156 ^ x70;
assign n_7158 = n_7066 ^ n_7156;
assign n_7159 = n_7157 & n_7158;
assign n_7160 = n_7159 ^ x70;
assign n_7161 = n_7160 ^ x71;
assign n_7162 = n_7067 ^ n_7160;
assign n_7163 = n_7161 & n_7162;
assign n_7164 = n_7163 ^ x71;
assign n_7165 = n_7164 ^ x72;
assign n_7166 = n_7068 ^ n_7164;
assign n_7167 = n_7165 & n_7166;
assign n_7168 = n_7167 ^ x72;
assign n_7169 = n_7168 ^ x73;
assign n_7170 = n_7069 ^ n_7168;
assign n_7171 = n_7169 & n_7170;
assign n_7172 = n_7171 ^ x73;
assign n_7173 = n_7172 ^ x74;
assign n_7174 = n_7070 ^ n_7172;
assign n_7175 = n_7173 & n_7174;
assign n_7176 = n_7175 ^ x74;
assign n_7177 = n_7176 ^ x75;
assign n_7178 = n_7071 ^ n_7176;
assign n_7179 = n_7177 & n_7178;
assign n_7180 = n_7179 ^ x75;
assign n_7181 = n_7180 ^ x76;
assign n_7182 = n_7072 ^ n_7180;
assign n_7183 = n_7181 & n_7182;
assign n_7184 = n_7183 ^ x76;
assign n_7185 = n_7184 ^ x77;
assign n_7186 = n_7073 ^ n_7184;
assign n_7187 = n_7185 & n_7186;
assign n_7188 = n_7187 ^ x77;
assign n_7189 = n_7188 ^ x78;
assign n_7190 = n_7074 ^ n_7188;
assign n_7191 = n_7189 & ~n_7190;
assign n_7192 = n_7191 ^ x78;
assign n_7193 = n_7192 ^ x79;
assign n_7194 = n_7075 ^ n_7192;
assign n_7195 = n_7193 & n_7194;
assign n_7196 = n_7195 ^ x79;
assign n_7197 = n_7196 ^ x80;
assign n_7198 = n_7196 ^ n_7061;
assign n_7199 = n_7135 & ~n_7196;
assign n_7200 = n_7197 & n_7198;
assign n_7201 = n_7142 & ~n_7199;
assign n_7202 = n_7200 ^ x80;
assign n_7203 = x82 ^ n_7201;
assign n_7204 = n_7076 ^ n_7201;
assign n_7205 = n_7202 ^ x81;
assign n_7206 = n_7203 & n_7204;
assign n_7207 = n_7206 ^ x82;
assign n_7208 = n_7207 ^ x83;
assign n_7209 = n_7077 ^ n_7207;
assign n_7210 = n_7208 & n_7209;
assign n_7211 = n_7210 ^ x83;
assign n_7212 = n_7211 ^ x84;
assign n_7213 = n_7078 ^ n_7211;
assign n_7214 = n_7212 & n_7213;
assign n_7215 = n_7214 ^ x84;
assign n_7216 = n_7215 ^ x85;
assign n_7217 = n_7079 ^ n_7215;
assign n_7218 = n_7216 & n_7217;
assign n_7219 = n_7218 ^ x85;
assign n_7220 = n_7219 ^ x86;
assign n_7221 = n_7080 ^ n_7219;
assign n_7222 = n_7220 & n_7221;
assign n_7223 = n_7222 ^ x86;
assign n_7224 = n_7223 ^ x87;
assign n_7225 = n_7081 ^ n_7223;
assign n_7226 = n_7224 & n_7225;
assign n_7227 = n_7226 ^ x87;
assign n_7228 = n_7227 ^ x88;
assign n_7229 = n_7082 ^ n_7227;
assign n_7230 = n_7228 & n_7229;
assign n_7231 = n_7230 ^ x88;
assign n_7232 = n_7231 ^ x89;
assign n_7233 = n_7083 ^ n_7231;
assign n_7234 = n_7232 & n_7233;
assign n_7235 = n_7234 ^ x89;
assign n_7236 = n_7235 ^ x90;
assign n_7237 = n_7084 ^ n_7235;
assign n_7238 = n_7236 & n_7237;
assign n_7239 = n_7238 ^ x90;
assign n_7240 = n_7239 ^ x91;
assign n_7241 = n_7085 ^ n_7239;
assign n_7242 = n_7240 & n_7241;
assign n_7243 = n_7242 ^ x91;
assign n_7244 = n_7243 ^ x92;
assign n_7245 = n_7086 ^ n_7243;
assign n_7246 = n_7244 & n_7245;
assign n_7247 = n_7246 ^ x92;
assign n_7248 = n_7247 ^ x93;
assign n_7249 = n_7087 ^ n_7247;
assign n_7250 = n_7248 & n_7249;
assign n_7251 = n_7250 ^ x93;
assign n_7252 = n_7251 ^ x94;
assign n_7253 = n_7088 ^ n_7251;
assign n_7254 = n_7252 & n_7253;
assign n_7255 = n_7254 ^ x94;
assign n_7256 = n_7255 ^ x95;
assign n_7257 = n_7089 ^ n_7255;
assign n_7258 = n_7256 & n_7257;
assign n_7259 = n_7258 ^ x95;
assign n_7260 = n_7259 ^ x96;
assign n_7261 = n_7090 ^ n_7259;
assign n_7262 = n_7260 & n_7261;
assign n_7263 = n_7262 ^ x96;
assign n_7264 = n_7263 ^ x97;
assign n_7265 = n_7263 ^ n_7059;
assign n_7266 = n_7133 & ~n_7263;
assign n_7267 = n_7264 & n_7265;
assign n_7268 = n_7141 & ~n_7266;
assign n_7269 = n_7267 ^ x97;
assign n_7270 = x99 ^ n_7268;
assign n_7271 = n_7092 ^ n_7268;
assign n_7272 = n_7137 & n_7268;
assign n_7273 = n_7269 ^ x98;
assign n_7274 = n_7270 & n_7271;
assign n_7275 = ~n_7143 & ~n_7272;
assign n_7276 = n_7274 ^ x99;
assign n_7277 = x101 ^ n_7275;
assign n_7278 = n_7093 ^ n_7275;
assign n_7279 = n_7276 ^ x100;
assign n_7280 = ~n_7277 & ~n_7278;
assign n_7281 = n_7280 ^ x101;
assign n_7282 = n_7281 ^ x102;
assign n_7283 = n_7094 ^ n_7281;
assign n_7284 = n_7282 & n_7283;
assign n_7285 = n_7284 ^ x102;
assign n_7286 = n_7285 ^ x103;
assign n_7287 = n_7095 ^ n_7285;
assign n_7288 = n_7286 & n_7287;
assign n_7289 = n_7288 ^ x103;
assign n_7290 = n_7289 ^ x104;
assign n_7291 = n_7096 ^ n_7289;
assign n_7292 = n_7290 & n_7291;
assign n_7293 = n_7292 ^ x104;
assign n_7294 = n_7293 ^ x105;
assign n_7295 = n_7097 ^ n_7293;
assign n_7296 = n_7294 & n_7295;
assign n_7297 = n_7296 ^ x105;
assign n_7298 = n_7297 ^ x106;
assign n_7299 = n_7297 ^ n_7057;
assign n_7300 = n_7131 & n_7297;
assign n_7301 = n_7298 & n_7299;
assign n_7302 = ~n_7140 & ~n_7300;
assign n_7303 = n_7301 ^ x106;
assign n_7304 = x108 ^ n_7302;
assign n_7305 = n_7098 ^ n_7302;
assign n_7306 = n_7303 ^ x107;
assign n_7307 = ~n_7304 & ~n_7305;
assign n_7308 = n_7307 ^ x108;
assign n_7309 = n_7308 ^ x109;
assign n_7310 = n_7308 & n_7101;
assign n_7311 = n_360 & n_7309;
assign n_7312 = ~n_7310 & n_5943;
assign n_7313 = ~n_7311 & n_7055;
assign n_7314 = n_7216 & n_7312;
assign n_7315 = n_7212 & n_7312;
assign n_7316 = x65 & n_7312;
assign n_7317 = x64 & n_7312;
assign n_7318 = ~n_7130 & n_7312;
assign n_7319 = n_7145 & n_7312;
assign n_7320 = n_7149 & n_7312;
assign n_7321 = n_7153 & n_7312;
assign n_7322 = n_7157 & n_7312;
assign n_7323 = n_7161 & n_7312;
assign n_7324 = n_7165 & n_7312;
assign n_7325 = n_7169 & n_7312;
assign n_7326 = n_7173 & n_7312;
assign n_7327 = n_7177 & n_7312;
assign n_7328 = n_7181 & n_7312;
assign n_7329 = n_7185 & n_7312;
assign n_7330 = n_7189 & n_7312;
assign n_7331 = n_7193 & n_7312;
assign n_7332 = n_7197 & n_7312;
assign n_7333 = n_7203 & n_7312;
assign n_7334 = n_7208 & n_7312;
assign n_7335 = n_7220 & n_7312;
assign n_7336 = n_7224 & n_7312;
assign n_7337 = n_7228 & n_7312;
assign n_7338 = n_7232 & n_7312;
assign n_7339 = n_7236 & n_7312;
assign n_7340 = n_7240 & n_7312;
assign n_7341 = n_7244 & n_7312;
assign n_7342 = n_7248 & n_7312;
assign n_7343 = n_7252 & n_7312;
assign n_7344 = n_7256 & n_7312;
assign n_7345 = n_7260 & n_7312;
assign n_7346 = n_7264 & n_7312;
assign n_7347 = n_7270 & n_7312;
assign n_7348 = ~n_7277 & n_7312;
assign n_7349 = n_7282 & n_7312;
assign n_7350 = n_7286 & n_7312;
assign n_7351 = n_7290 & n_7312;
assign n_7352 = n_7294 & n_7312;
assign n_7353 = n_7298 & n_7312;
assign n_7354 = ~n_7304 & n_7312;
assign y18 = n_7312;
assign n_7355 = n_7205 & n_7312;
assign n_7356 = n_7273 & n_7312;
assign n_7357 = n_7279 & n_7312;
assign n_7358 = n_7306 & n_7312;
assign n_7359 = x110 ^ n_7313;
assign n_7360 = n_7314 ^ n_7079;
assign n_7361 = n_7315 ^ n_7078;
assign n_7362 = n_7317 ^ x18;
assign n_7363 = n_7318 ^ n_7114;
assign n_7364 = n_7319 ^ n_7100;
assign n_7365 = n_7320 ^ n_7064;
assign n_7366 = n_7321 ^ n_7065;
assign n_7367 = n_7322 ^ n_7066;
assign n_7368 = n_7323 ^ n_7067;
assign n_7369 = n_7324 ^ n_7068;
assign n_7370 = n_7325 ^ n_7069;
assign n_7371 = n_7326 ^ n_7070;
assign n_7372 = n_7327 ^ n_7071;
assign n_7373 = n_7328 ^ n_7072;
assign n_7374 = n_7329 ^ n_7073;
assign n_7375 = n_7330 ^ n_7074;
assign n_7376 = n_7331 ^ n_7075;
assign n_7377 = n_7332 ^ n_7061;
assign n_7378 = n_7333 ^ n_7076;
assign n_7379 = n_7334 ^ n_7077;
assign n_7380 = n_7335 ^ n_7080;
assign n_7381 = n_7336 ^ n_7081;
assign n_7382 = n_7337 ^ n_7082;
assign n_7383 = n_7338 ^ n_7083;
assign n_7384 = n_7339 ^ n_7084;
assign n_7385 = n_7340 ^ n_7085;
assign n_7386 = n_7341 ^ n_7086;
assign n_7387 = n_7342 ^ n_7087;
assign n_7388 = n_7343 ^ n_7088;
assign n_7389 = n_7344 ^ n_7089;
assign n_7390 = n_7345 ^ n_7090;
assign n_7391 = n_7346 ^ n_7059;
assign n_7392 = n_7347 ^ n_7092;
assign n_7393 = n_7348 ^ n_7093;
assign n_7394 = n_7349 ^ n_7094;
assign n_7395 = n_7350 ^ n_7095;
assign n_7396 = n_7351 ^ n_7096;
assign n_7397 = n_7352 ^ n_7097;
assign n_7398 = n_7353 ^ n_7057;
assign n_7399 = n_7354 ^ n_7098;
assign n_7400 = n_7060 ^ n_7355;
assign n_7401 = n_7058 ^ n_7356;
assign n_7402 = n_7091 ^ n_7357;
assign n_7403 = n_7056 ^ n_7358;
assign n_7404 = ~x86 ^ n_7360;
assign n_7405 = n_7360 ^ x86;
assign n_7406 = n_7361 ^ x85;
assign n_7407 = x85 & ~n_7361;
assign n_7408 = n_7317 & n_7362;
assign n_7409 = n_7362 ^ x65;
assign n_7410 = n_27 ^ n_7362;
assign n_7411 = ~n_7362 & n_222;
assign n_7412 = n_7362 & ~n_223;
assign n_7413 = ~n_7362 & n_163;
assign n_7414 = n_7406 ^ n_7407;
assign n_7415 = n_7407 ^ n_7360;
assign n_7416 = n_7408 ^ n_7017;
assign n_7417 = x17 & n_7409;
assign n_7418 = ~n_7409 & n_7410;
assign n_7419 = n_7411 ^ n_222;
assign n_7420 = ~x66 & ~n_7413;
assign n_7421 = n_7404 & ~n_7414;
assign n_7422 = ~n_7405 & n_7415;
assign n_7423 = n_7316 ^ n_7416;
assign n_7424 = n_60 & n_7417;
assign n_7425 = n_7418 ^ x65;
assign n_7426 = n_7419 ^ n_7409;
assign n_7427 = n_7422 ^ x86;
assign n_7428 = n_7423 ^ x19;
assign n_7429 = n_7425 ^ x66;
assign n_7430 = n_27 & ~n_7426;
assign n_7431 = n_7428 ^ x66;
assign n_7432 = n_7425 ^ n_7428;
assign n_7433 = n_7430 ^ n_7424;
assign n_7434 = ~n_7431 & n_7432;
assign n_7435 = n_7434 ^ x66;
assign n_7436 = n_7435 ^ x67;
assign n_7437 = n_7363 ^ n_7435;
assign n_7438 = n_7436 & n_7437;
assign n_7439 = n_7438 ^ x67;
assign n_7440 = n_7439 ^ x68;
assign n_7441 = n_7364 ^ n_7439;
assign n_7442 = n_7440 & n_7441;
assign n_7443 = n_7442 ^ x68;
assign n_7444 = n_7443 ^ x69;
assign n_7445 = n_7365 ^ n_7443;
assign n_7446 = n_7444 & n_7445;
assign n_7447 = n_7446 ^ x69;
assign n_7448 = n_7447 ^ x70;
assign n_7449 = n_7366 ^ n_7447;
assign n_7450 = n_7448 & n_7449;
assign n_7451 = n_7450 ^ x70;
assign n_7452 = n_7451 ^ x71;
assign n_7453 = n_7367 ^ n_7451;
assign n_7454 = n_7452 & n_7453;
assign n_7455 = n_7454 ^ x71;
assign n_7456 = n_7455 ^ x72;
assign n_7457 = n_7368 ^ n_7455;
assign n_7458 = n_7456 & n_7457;
assign n_7459 = n_7458 ^ x72;
assign n_7460 = n_7459 ^ x73;
assign n_7461 = n_7369 ^ n_7459;
assign n_7462 = n_7460 & n_7461;
assign n_7463 = n_7462 ^ x73;
assign n_7464 = n_7463 ^ x74;
assign n_7465 = n_7370 ^ n_7463;
assign n_7466 = n_7464 & n_7465;
assign n_7467 = n_7466 ^ x74;
assign n_7468 = n_7467 ^ x75;
assign n_7469 = n_7371 ^ n_7467;
assign n_7470 = n_7468 & n_7469;
assign n_7471 = n_7470 ^ x75;
assign n_7472 = n_7471 ^ x76;
assign n_7473 = n_7372 ^ n_7471;
assign n_7474 = n_7472 & n_7473;
assign n_7475 = n_7474 ^ x76;
assign n_7476 = n_7475 ^ x77;
assign n_7477 = n_7373 ^ n_7475;
assign n_7478 = n_7476 & n_7477;
assign n_7479 = n_7478 ^ x77;
assign n_7480 = n_7479 ^ x78;
assign n_7481 = n_7374 ^ n_7479;
assign n_7482 = n_7480 & n_7481;
assign n_7483 = n_7482 ^ x78;
assign n_7484 = n_7483 ^ x79;
assign n_7485 = n_7375 ^ n_7483;
assign n_7486 = n_7484 & ~n_7485;
assign n_7487 = n_7486 ^ x79;
assign n_7488 = n_7487 ^ x80;
assign n_7489 = n_7376 ^ n_7487;
assign n_7490 = n_7488 & n_7489;
assign n_7491 = n_7490 ^ x80;
assign n_7492 = n_7491 ^ x81;
assign n_7493 = n_7377 ^ n_7491;
assign n_7494 = n_7492 & n_7493;
assign n_7495 = n_7494 ^ x81;
assign n_7496 = n_7495 ^ x82;
assign n_7497 = n_7400 ^ n_7495;
assign n_7498 = n_7496 & n_7497;
assign n_7499 = n_7498 ^ x82;
assign n_7500 = n_7499 ^ x83;
assign n_7501 = n_7378 ^ n_7499;
assign n_7502 = n_7500 & n_7501;
assign n_7503 = n_7502 ^ x83;
assign n_7504 = n_7503 ^ x84;
assign n_7505 = n_7379 ^ n_7503;
assign n_7506 = n_7504 & n_7505;
assign n_7507 = n_7506 ^ x84;
assign n_7508 = n_7507 ^ x85;
assign n_7509 = n_7507 ^ n_7361;
assign n_7510 = n_7421 & n_7507;
assign n_7511 = n_7508 & n_7509;
assign n_7512 = ~n_7427 & ~n_7510;
assign n_7513 = n_7511 ^ x85;
assign n_7514 = x87 ^ n_7512;
assign n_7515 = n_7380 ^ n_7512;
assign n_7516 = n_7513 ^ x86;
assign n_7517 = ~n_7514 & ~n_7515;
assign n_7518 = n_7517 ^ x87;
assign n_7519 = n_7518 ^ x88;
assign n_7520 = n_7381 ^ n_7518;
assign n_7521 = n_7519 & n_7520;
assign n_7522 = n_7521 ^ x88;
assign n_7523 = n_7522 ^ x89;
assign n_7524 = n_7382 ^ n_7522;
assign n_7525 = n_7523 & n_7524;
assign n_7526 = n_7525 ^ x89;
assign n_7527 = n_7526 ^ x90;
assign n_7528 = n_7383 ^ n_7526;
assign n_7529 = n_7527 & n_7528;
assign n_7530 = n_7529 ^ x90;
assign n_7531 = n_7530 ^ x91;
assign n_7532 = n_7384 ^ n_7530;
assign n_7533 = n_7531 & n_7532;
assign n_7534 = n_7533 ^ x91;
assign n_7535 = n_7534 ^ x92;
assign n_7536 = n_7385 ^ n_7534;
assign n_7537 = n_7535 & n_7536;
assign n_7538 = n_7537 ^ x92;
assign n_7539 = n_7538 ^ x93;
assign n_7540 = n_7386 ^ n_7538;
assign n_7541 = n_7539 & n_7540;
assign n_7542 = n_7541 ^ x93;
assign n_7543 = n_7542 ^ x94;
assign n_7544 = n_7387 ^ n_7542;
assign n_7545 = n_7543 & n_7544;
assign n_7546 = n_7545 ^ x94;
assign n_7547 = n_7546 ^ x95;
assign n_7548 = n_7388 ^ n_7546;
assign n_7549 = n_7547 & n_7548;
assign n_7550 = n_7549 ^ x95;
assign n_7551 = n_7550 ^ x96;
assign n_7552 = n_7389 ^ n_7550;
assign n_7553 = n_7551 & n_7552;
assign n_7554 = n_7553 ^ x96;
assign n_7555 = n_7554 ^ x97;
assign n_7556 = n_7390 ^ n_7554;
assign n_7557 = n_7555 & n_7556;
assign n_7558 = n_7557 ^ x97;
assign n_7559 = n_7558 ^ x98;
assign n_7560 = n_7391 ^ n_7558;
assign n_7561 = n_7559 & n_7560;
assign n_7562 = n_7561 ^ x98;
assign n_7563 = n_7562 ^ x99;
assign n_7564 = n_7401 ^ n_7562;
assign n_7565 = n_7563 & n_7564;
assign n_7566 = n_7565 ^ x99;
assign n_7567 = n_7566 ^ x100;
assign n_7568 = n_7392 ^ n_7566;
assign n_7569 = n_7567 & n_7568;
assign n_7570 = n_7569 ^ x100;
assign n_7571 = n_7570 ^ x101;
assign n_7572 = n_7402 ^ n_7570;
assign n_7573 = n_7571 & n_7572;
assign n_7574 = n_7573 ^ x101;
assign n_7575 = n_7574 ^ x102;
assign n_7576 = n_7393 ^ n_7574;
assign n_7577 = n_7575 & n_7576;
assign n_7578 = n_7577 ^ x102;
assign n_7579 = n_7578 ^ x103;
assign n_7580 = n_7394 ^ n_7578;
assign n_7581 = n_7579 & n_7580;
assign n_7582 = n_7581 ^ x103;
assign n_7583 = n_7582 ^ x104;
assign n_7584 = n_7395 ^ n_7582;
assign n_7585 = n_7583 & n_7584;
assign n_7586 = n_7585 ^ x104;
assign n_7587 = n_7586 ^ x105;
assign n_7588 = n_7396 ^ n_7586;
assign n_7589 = n_7587 & n_7588;
assign n_7590 = n_7589 ^ x105;
assign n_7591 = n_7590 ^ x106;
assign n_7592 = n_7397 ^ n_7590;
assign n_7593 = n_7591 & n_7592;
assign n_7594 = n_7593 ^ x106;
assign n_7595 = n_7594 ^ x107;
assign n_7596 = n_7398 ^ n_7594;
assign n_7597 = n_7595 & n_7596;
assign n_7598 = n_7597 ^ x107;
assign n_7599 = n_7598 ^ x108;
assign n_7600 = n_7403 ^ n_7598;
assign n_7601 = n_7599 & n_7600;
assign n_7602 = n_7601 ^ x108;
assign n_7603 = n_7602 ^ x109;
assign n_7604 = n_7399 ^ n_7602;
assign n_7605 = n_7603 & n_7604;
assign n_7606 = n_7605 ^ x109;
assign n_7607 = ~n_7606 & n_358;
assign n_7608 = n_7606 ^ x110;
assign n_7609 = n_7607 ^ n_360;
assign n_7610 = n_7608 & ~n_7359;
assign n_7611 = ~n_7609 & n_7313;
assign n_7612 = n_7610 ^ x110;
assign n_7613 = n_7313 ^ n_7611;
assign n_7614 = ~n_7612 & n_358;
assign n_7615 = n_7603 & n_7614;
assign n_7616 = n_7591 & n_7614;
assign n_7617 = n_7587 & n_7614;
assign n_7618 = n_7567 & n_7614;
assign n_7619 = n_7563 & n_7614;
assign n_7620 = n_7543 & n_7614;
assign n_7621 = n_7539 & n_7614;
assign n_7622 = n_7444 & n_7614;
assign n_7623 = n_7440 & n_7614;
assign n_7624 = x17 & n_7614;
assign n_7625 = n_7411 & ~n_7614;
assign n_7626 = x64 & n_7614;
assign n_7627 = n_7362 ^ n_7614;
assign n_7628 = ~x65 & n_7614;
assign n_7629 = n_93 ^ ~n_7614;
assign n_7630 = n_161 & n_7614;
assign n_7631 = n_7429 & n_7614;
assign n_7632 = n_7436 & n_7614;
assign n_7633 = n_7448 & n_7614;
assign n_7634 = n_7452 & n_7614;
assign n_7635 = n_7456 & n_7614;
assign n_7636 = n_7460 & n_7614;
assign n_7637 = n_7464 & n_7614;
assign n_7638 = n_7468 & n_7614;
assign n_7639 = n_7472 & n_7614;
assign n_7640 = n_7476 & n_7614;
assign n_7641 = n_7480 & n_7614;
assign n_7642 = n_7484 & n_7614;
assign n_7643 = n_7488 & n_7614;
assign n_7644 = n_7492 & n_7614;
assign n_7645 = n_7496 & n_7614;
assign n_7646 = n_7500 & n_7614;
assign n_7647 = n_7504 & n_7614;
assign n_7648 = n_7508 & n_7614;
assign n_7649 = ~n_7514 & n_7614;
assign n_7650 = n_7519 & n_7614;
assign n_7651 = n_7523 & n_7614;
assign n_7652 = n_7527 & n_7614;
assign n_7653 = n_7531 & n_7614;
assign n_7654 = n_7535 & n_7614;
assign n_7655 = n_7547 & n_7614;
assign n_7656 = n_7551 & n_7614;
assign n_7657 = n_7555 & n_7614;
assign n_7658 = n_7559 & n_7614;
assign n_7659 = n_7571 & n_7614;
assign n_7660 = n_7575 & n_7614;
assign n_7661 = n_7579 & n_7614;
assign n_7662 = n_7583 & n_7614;
assign n_7663 = n_7595 & n_7614;
assign n_7664 = n_7599 & n_7614;
assign n_7665 = n_162 & n_7614;
assign y17 = n_7614;
assign n_7666 = n_7433 & n_7614;
assign n_7667 = n_7516 & n_7614;
assign n_7668 = n_7615 ^ n_7399;
assign n_7669 = n_7616 ^ n_7397;
assign n_7670 = n_7617 ^ n_7396;
assign n_7671 = n_7618 ^ n_7392;
assign n_7672 = n_7619 ^ n_7401;
assign n_7673 = n_7620 ^ n_7387;
assign n_7674 = n_7621 ^ n_7386;
assign n_7675 = n_7622 ^ n_7365;
assign n_7676 = n_7623 ^ n_7364;
assign n_7677 = ~n_90 & n_7624;
assign n_7678 = ~n_7626 & n_223;
assign n_7679 = ~x16 & ~n_7628;
assign n_7680 = n_28 & n_7629;
assign n_7681 = ~n_7630 & n_7412;
assign n_7682 = n_7631 ^ n_7428;
assign n_7683 = n_7632 ^ n_7363;
assign n_7684 = n_7633 ^ n_7366;
assign n_7685 = n_7634 ^ n_7367;
assign n_7686 = n_7635 ^ n_7368;
assign n_7687 = n_7636 ^ n_7369;
assign n_7688 = n_7637 ^ n_7370;
assign n_7689 = n_7638 ^ n_7371;
assign n_7690 = n_7639 ^ n_7372;
assign n_7691 = n_7640 ^ n_7373;
assign n_7692 = n_7641 ^ n_7374;
assign n_7693 = n_7642 ^ n_7375;
assign n_7694 = n_7643 ^ n_7376;
assign n_7695 = n_7644 ^ n_7377;
assign n_7696 = n_7645 ^ n_7400;
assign n_7697 = n_7646 ^ n_7378;
assign n_7698 = n_7647 ^ n_7379;
assign n_7699 = n_7648 ^ n_7361;
assign n_7700 = n_7649 ^ n_7380;
assign n_7701 = n_7650 ^ n_7381;
assign n_7702 = n_7651 ^ n_7382;
assign n_7703 = n_7652 ^ n_7383;
assign n_7704 = n_7653 ^ n_7384;
assign n_7705 = n_7654 ^ n_7385;
assign n_7706 = n_7655 ^ n_7388;
assign n_7707 = n_7656 ^ n_7389;
assign n_7708 = n_7657 ^ n_7390;
assign n_7709 = n_7658 ^ n_7391;
assign n_7710 = n_7659 ^ n_7402;
assign n_7711 = n_7660 ^ n_7393;
assign n_7712 = n_7661 ^ n_7394;
assign n_7713 = n_7662 ^ n_7395;
assign n_7714 = n_7663 ^ n_7398;
assign n_7715 = n_7664 ^ n_7403;
assign n_7716 = n_7665 ^ n_7362;
assign n_7717 = n_7360 ^ n_7667;
assign n_7718 = n_7668 ^ x110;
assign n_7719 = n_7669 ^ x107;
assign n_7720 = n_7670 ^ x106;
assign n_7721 = n_7671 ^ x101;
assign n_7722 = n_7672 ^ x100;
assign n_7723 = n_7673 ^ x95;
assign n_7724 = n_7674 ^ x94;
assign n_7725 = n_7675 ^ x70;
assign n_7726 = n_7676 ^ x69;
assign n_7727 = ~n_7409 & n_7677;
assign n_7728 = n_7678 & ~n_7627;
assign n_7729 = ~n_93 & n_7679;
assign n_7730 = ~n_7680 & n_7681;
assign n_7731 = n_7727 ^ n_7625;
assign n_7732 = ~n_7728 & n_7420;
assign n_7733 = ~n_7677 & ~n_7729;
assign n_7734 = ~n_7730 ^ ~n_7666;
assign n_7735 = x64 & n_7731;
assign n_7736 = x64 & ~n_7733;
assign n_7737 = ~n_7735 & n_7732;
assign n_7738 = ~n_7678 & ~n_7736;
assign n_7739 = ~n_7734 & ~n_7737;
assign n_7740 = x66 ^ n_7738;
assign n_7741 = x67 ^ n_7739;
assign n_7742 = n_7682 ^ n_7739;
assign n_7743 = n_7741 & n_7742;
assign n_7744 = n_7743 ^ x67;
assign n_7745 = n_7744 ^ x68;
assign n_7746 = n_7683 ^ n_7744;
assign n_7747 = n_7745 & n_7746;
assign n_7748 = n_7747 ^ x68;
assign n_7749 = n_7748 ^ n_7676;
assign n_7750 = n_7748 ^ x69;
assign n_7751 = ~n_7726 & n_7749;
assign n_7752 = n_7751 ^ x69;
assign n_7753 = n_7752 ^ n_7675;
assign n_7754 = n_7752 ^ x70;
assign n_7755 = ~n_7725 & n_7753;
assign n_7756 = n_7755 ^ x70;
assign n_7757 = n_7756 ^ x71;
assign n_7758 = n_7684 ^ n_7756;
assign n_7759 = n_7757 & n_7758;
assign n_7760 = n_7759 ^ x71;
assign n_7761 = n_7760 ^ x72;
assign n_7762 = n_7685 ^ n_7760;
assign n_7763 = n_7761 & n_7762;
assign n_7764 = n_7763 ^ x72;
assign n_7765 = n_7764 ^ x73;
assign n_7766 = n_7686 ^ n_7764;
assign n_7767 = n_7765 & n_7766;
assign n_7768 = n_7767 ^ x73;
assign n_7769 = n_7768 ^ x74;
assign n_7770 = n_7687 ^ n_7768;
assign n_7771 = n_7769 & n_7770;
assign n_7772 = n_7771 ^ x74;
assign n_7773 = n_7772 ^ x75;
assign n_7774 = n_7688 ^ n_7772;
assign n_7775 = n_7773 & n_7774;
assign n_7776 = n_7775 ^ x75;
assign n_7777 = n_7776 ^ x76;
assign n_7778 = n_7689 ^ n_7776;
assign n_7779 = n_7777 & n_7778;
assign n_7780 = n_7779 ^ x76;
assign n_7781 = n_7780 ^ x77;
assign n_7782 = n_7690 ^ n_7780;
assign n_7783 = n_7781 & n_7782;
assign n_7784 = n_7783 ^ x77;
assign n_7785 = n_7784 ^ x78;
assign n_7786 = n_7691 ^ n_7784;
assign n_7787 = n_7785 & n_7786;
assign n_7788 = n_7787 ^ x78;
assign n_7789 = n_7788 ^ x79;
assign n_7790 = n_7692 ^ n_7788;
assign n_7791 = n_7789 & n_7790;
assign n_7792 = n_7791 ^ x79;
assign n_7793 = n_7792 ^ x80;
assign n_7794 = n_7693 ^ n_7792;
assign n_7795 = n_7793 & ~n_7794;
assign n_7796 = n_7795 ^ x80;
assign n_7797 = n_7796 ^ x81;
assign n_7798 = n_7694 ^ n_7796;
assign n_7799 = n_7797 & n_7798;
assign n_7800 = n_7799 ^ x81;
assign n_7801 = n_7800 ^ x82;
assign n_7802 = n_7695 ^ n_7800;
assign n_7803 = n_7801 & n_7802;
assign n_7804 = n_7803 ^ x82;
assign n_7805 = n_7804 ^ x83;
assign n_7806 = n_7696 ^ n_7804;
assign n_7807 = n_7805 & n_7806;
assign n_7808 = n_7807 ^ x83;
assign n_7809 = n_7808 ^ x84;
assign n_7810 = n_7697 ^ n_7808;
assign n_7811 = n_7809 & n_7810;
assign n_7812 = n_7811 ^ x84;
assign n_7813 = n_7812 ^ x85;
assign n_7814 = n_7698 ^ n_7812;
assign n_7815 = n_7813 & n_7814;
assign n_7816 = n_7815 ^ x85;
assign n_7817 = n_7816 ^ x86;
assign n_7818 = n_7699 ^ n_7816;
assign n_7819 = n_7817 & n_7818;
assign n_7820 = n_7819 ^ x86;
assign n_7821 = n_7820 ^ x87;
assign n_7822 = n_7717 ^ n_7820;
assign n_7823 = n_7821 & n_7822;
assign n_7824 = n_7823 ^ x87;
assign n_7825 = n_7824 ^ x88;
assign n_7826 = n_7700 ^ n_7824;
assign n_7827 = n_7825 & n_7826;
assign n_7828 = n_7827 ^ x88;
assign n_7829 = n_7828 ^ x89;
assign n_7830 = n_7701 ^ n_7828;
assign n_7831 = n_7829 & n_7830;
assign n_7832 = n_7831 ^ x89;
assign n_7833 = n_7832 ^ x90;
assign n_7834 = n_7702 ^ n_7832;
assign n_7835 = n_7833 & n_7834;
assign n_7836 = n_7835 ^ x90;
assign n_7837 = n_7836 ^ x91;
assign n_7838 = n_7703 ^ n_7836;
assign n_7839 = n_7837 & n_7838;
assign n_7840 = n_7839 ^ x91;
assign n_7841 = n_7840 ^ x92;
assign n_7842 = n_7704 ^ n_7840;
assign n_7843 = n_7841 & n_7842;
assign n_7844 = n_7843 ^ x92;
assign n_7845 = n_7844 ^ x93;
assign n_7846 = n_7705 ^ n_7844;
assign n_7847 = n_7845 & n_7846;
assign n_7848 = n_7847 ^ x93;
assign n_7849 = n_7848 ^ n_7674;
assign n_7850 = n_7848 ^ x94;
assign n_7851 = ~n_7724 & n_7849;
assign n_7852 = n_7851 ^ x94;
assign n_7853 = n_7852 ^ n_7673;
assign n_7854 = n_7852 ^ x95;
assign n_7855 = ~n_7723 & n_7853;
assign n_7856 = n_7855 ^ x95;
assign n_7857 = n_7856 ^ x96;
assign n_7858 = n_7706 ^ n_7856;
assign n_7859 = n_7857 & n_7858;
assign n_7860 = n_7859 ^ x96;
assign n_7861 = n_7860 ^ x97;
assign n_7862 = n_7707 ^ n_7860;
assign n_7863 = n_7861 & n_7862;
assign n_7864 = n_7863 ^ x97;
assign n_7865 = n_7864 ^ x98;
assign n_7866 = n_7708 ^ n_7864;
assign n_7867 = n_7865 & n_7866;
assign n_7868 = n_7867 ^ x98;
assign n_7869 = n_7868 ^ x99;
assign n_7870 = n_7709 ^ n_7868;
assign n_7871 = n_7869 & n_7870;
assign n_7872 = n_7871 ^ x99;
assign n_7873 = n_7872 ^ n_7672;
assign n_7874 = n_7872 ^ x100;
assign n_7875 = ~n_7722 & n_7873;
assign n_7876 = n_7875 ^ x100;
assign n_7877 = n_7876 ^ n_7671;
assign n_7878 = n_7876 ^ x101;
assign n_7879 = ~n_7721 & n_7877;
assign n_7880 = n_7879 ^ x101;
assign n_7881 = n_7880 ^ x102;
assign n_7882 = n_7710 ^ n_7880;
assign n_7883 = n_7881 & n_7882;
assign n_7884 = n_7883 ^ x102;
assign n_7885 = n_7884 ^ x103;
assign n_7886 = n_7711 ^ n_7884;
assign n_7887 = n_7885 & n_7886;
assign n_7888 = n_7887 ^ x103;
assign n_7889 = n_7888 ^ x104;
assign n_7890 = n_7712 ^ n_7888;
assign n_7891 = n_7889 & n_7890;
assign n_7892 = n_7891 ^ x104;
assign n_7893 = n_7892 ^ x105;
assign n_7894 = n_7713 ^ n_7892;
assign n_7895 = n_7893 & n_7894;
assign n_7896 = n_7895 ^ x105;
assign n_7897 = n_7896 ^ n_7670;
assign n_7898 = n_7896 ^ x106;
assign n_7899 = ~n_7720 & n_7897;
assign n_7900 = n_7899 ^ x106;
assign n_7901 = n_7900 ^ n_7669;
assign n_7902 = n_7900 ^ x107;
assign n_7903 = ~n_7719 & n_7901;
assign n_7904 = n_7903 ^ x107;
assign n_7905 = n_7904 ^ x108;
assign n_7906 = n_7714 ^ n_7904;
assign n_7907 = n_7905 & n_7906;
assign n_7908 = n_7907 ^ x108;
assign n_7909 = n_7908 ^ x109;
assign n_7910 = n_7715 ^ n_7908;
assign n_7911 = n_7909 & n_7910;
assign n_7912 = n_7911 ^ x109;
assign n_7913 = n_7912 ^ n_7668;
assign n_7914 = n_7912 ^ x110;
assign n_7915 = ~n_7718 & n_7913;
assign n_7916 = n_7915 ^ x110;
assign n_7917 = n_7916 ^ x111;
assign n_7918 = n_7916 ^ ~n_7613;
assign n_7919 = ~n_7918 ^ n_7313;
assign n_7920 = n_7917 & n_7919;
assign n_7921 = n_7920 ^ x111;
assign n_7922 = n_359 & ~n_7921;
assign n_7923 = n_7909 & n_7922;
assign n_7924 = n_7905 & n_7922;
assign n_7925 = n_7889 & n_7922;
assign n_7926 = n_7885 & n_7922;
assign n_7927 = n_7797 & n_7922;
assign n_7928 = n_7793 & n_7922;
assign n_7929 = n_164 & n_7922;
assign n_7930 = x64 & n_7922;
assign n_7931 = n_7741 & n_7922;
assign n_7932 = n_7745 & n_7922;
assign n_7933 = n_7750 & n_7922;
assign n_7934 = n_7754 & n_7922;
assign n_7935 = n_7757 & n_7922;
assign n_7936 = n_7761 & n_7922;
assign n_7937 = n_7765 & n_7922;
assign n_7938 = n_7769 & n_7922;
assign n_7939 = n_7773 & n_7922;
assign n_7940 = n_7777 & n_7922;
assign n_7941 = n_7781 & n_7922;
assign n_7942 = n_7785 & n_7922;
assign n_7943 = n_7789 & n_7922;
assign n_7944 = n_7801 & n_7922;
assign n_7945 = n_7805 & n_7922;
assign n_7946 = n_7809 & n_7922;
assign n_7947 = n_7813 & n_7922;
assign n_7948 = n_7817 & n_7922;
assign n_7949 = n_7821 & n_7922;
assign n_7950 = n_7825 & n_7922;
assign n_7951 = n_7829 & n_7922;
assign n_7952 = n_7833 & n_7922;
assign n_7953 = n_7837 & n_7922;
assign n_7954 = n_7841 & n_7922;
assign n_7955 = n_7845 & n_7922;
assign n_7956 = n_7850 & n_7922;
assign n_7957 = n_7854 & n_7922;
assign n_7958 = n_7857 & n_7922;
assign n_7959 = n_7861 & n_7922;
assign n_7960 = n_7865 & n_7922;
assign n_7961 = n_7869 & n_7922;
assign n_7962 = n_7874 & n_7922;
assign n_7963 = n_7878 & n_7922;
assign n_7964 = n_7881 & n_7922;
assign n_7965 = n_7893 & n_7922;
assign n_7966 = n_7898 & n_7922;
assign n_7967 = n_7902 & n_7922;
assign n_7968 = n_7914 & n_7922;
assign y16 = n_7922;
assign n_7969 = n_280 & ~n_7922;
assign n_7970 = ~n_7740 & n_7922;
assign n_7971 = n_7923 ^ n_7715;
assign n_7972 = n_7924 ^ n_7714;
assign n_7973 = n_7925 ^ n_7712;
assign n_7974 = n_7926 ^ n_7711;
assign n_7975 = n_7927 ^ n_7694;
assign n_7976 = n_7928 ^ n_7693;
assign n_7977 = n_7929 ^ n_7626;
assign n_7978 = n_7930 & n_279;
assign n_7979 = n_7931 ^ n_7682;
assign n_7980 = n_7932 ^ n_7683;
assign n_7981 = n_7933 ^ n_7676;
assign n_7982 = n_7934 ^ n_7675;
assign n_7983 = n_7935 ^ n_7684;
assign n_7984 = n_7936 ^ n_7685;
assign n_7985 = n_7937 ^ n_7686;
assign n_7986 = n_7938 ^ n_7687;
assign n_7987 = n_7939 ^ n_7688;
assign n_7988 = n_7940 ^ n_7689;
assign n_7989 = n_7941 ^ n_7690;
assign n_7990 = n_7942 ^ n_7691;
assign n_7991 = n_7943 ^ n_7692;
assign n_7992 = n_7944 ^ n_7695;
assign n_7993 = n_7945 ^ n_7696;
assign n_7994 = n_7946 ^ n_7697;
assign n_7995 = n_7947 ^ n_7698;
assign n_7996 = n_7948 ^ n_7699;
assign n_7997 = n_7949 ^ n_7717;
assign n_7998 = n_7950 ^ n_7700;
assign n_7999 = n_7951 ^ n_7701;
assign n_8000 = n_7952 ^ n_7702;
assign n_8001 = n_7953 ^ n_7703;
assign n_8002 = n_7954 ^ n_7704;
assign n_8003 = n_7955 ^ n_7705;
assign n_8004 = n_7956 ^ n_7674;
assign n_8005 = n_7957 ^ n_7673;
assign n_8006 = n_7958 ^ n_7706;
assign n_8007 = n_7959 ^ n_7707;
assign n_8008 = n_7960 ^ n_7708;
assign n_8009 = n_7961 ^ n_7709;
assign n_8010 = n_7962 ^ n_7672;
assign n_8011 = n_7963 ^ n_7671;
assign n_8012 = n_7964 ^ n_7710;
assign n_8013 = n_7965 ^ n_7713;
assign n_8014 = n_7966 ^ n_7670;
assign n_8015 = n_7967 ^ n_7669;
assign n_8016 = n_7968 ^ n_7668;
assign n_8017 = ~n_325 & ~n_7969;
assign n_8018 = n_7716 ^ n_7970;
assign n_8019 = n_7971 ^ x110;
assign n_8020 = n_7972 ^ x109;
assign n_8021 = ~x105 ^ n_7973;
assign n_8022 = n_7973 ^ x105;
assign n_8023 = n_7974 ^ x104;
assign n_8024 = x104 & ~n_7974;
assign n_8025 = ~x82 ^ n_7975;
assign n_8026 = n_7975 ^ x82;
assign n_8027 = n_7976 ^ x81;
assign n_8028 = x81 & n_7976;
assign n_8029 = n_7977 ^ x17;
assign n_8030 = ~n_7978 & n_8017;
assign n_8031 = n_8023 ^ n_8024;
assign n_8032 = n_8024 ^ n_7973;
assign n_8033 = n_8027 ^ n_8028;
assign n_8034 = n_8028 ^ n_7975;
assign n_8035 = n_8029 ^ x66;
assign n_8036 = n_8029 ^ n_8030;
assign n_8037 = x66 ^ n_8030;
assign n_8038 = n_8021 & ~n_8031;
assign n_8039 = ~n_8022 & n_8032;
assign n_8040 = n_8025 & n_8033;
assign n_8041 = ~n_8026 & n_8034;
assign n_8042 = ~n_8035 & ~n_8036;
assign n_8043 = n_8039 ^ x105;
assign n_8044 = n_8041 ^ x82;
assign n_8045 = n_8042 ^ x66;
assign n_8046 = n_8045 ^ x67;
assign n_8047 = n_8018 ^ n_8045;
assign n_8048 = n_8046 & n_8047;
assign n_8049 = n_8048 ^ x67;
assign n_8050 = n_8049 ^ x68;
assign n_8051 = n_7979 ^ n_8049;
assign n_8052 = n_8050 & n_8051;
assign n_8053 = n_8052 ^ x68;
assign n_8054 = n_8053 ^ x69;
assign n_8055 = n_7980 ^ n_8053;
assign n_8056 = n_8054 & n_8055;
assign n_8057 = n_8056 ^ x69;
assign n_8058 = n_8057 ^ x70;
assign n_8059 = n_7981 ^ n_8057;
assign n_8060 = n_8058 & n_8059;
assign n_8061 = n_8060 ^ x70;
assign n_8062 = n_8061 ^ x71;
assign n_8063 = n_7982 ^ n_8061;
assign n_8064 = n_8062 & n_8063;
assign n_8065 = n_8064 ^ x71;
assign n_8066 = n_8065 ^ x72;
assign n_8067 = n_7983 ^ n_8065;
assign n_8068 = n_8066 & n_8067;
assign n_8069 = n_8068 ^ x72;
assign n_8070 = n_8069 ^ x73;
assign n_8071 = n_7984 ^ n_8069;
assign n_8072 = n_8070 & n_8071;
assign n_8073 = n_8072 ^ x73;
assign n_8074 = n_8073 ^ x74;
assign n_8075 = n_7985 ^ n_8073;
assign n_8076 = n_8074 & n_8075;
assign n_8077 = n_8076 ^ x74;
assign n_8078 = n_8077 ^ x75;
assign n_8079 = n_7986 ^ n_8077;
assign n_8080 = n_8078 & n_8079;
assign n_8081 = n_8080 ^ x75;
assign n_8082 = n_8081 ^ x76;
assign n_8083 = n_7987 ^ n_8081;
assign n_8084 = n_8082 & n_8083;
assign n_8085 = n_8084 ^ x76;
assign n_8086 = n_8085 ^ x77;
assign n_8087 = n_7988 ^ n_8085;
assign n_8088 = n_8086 & n_8087;
assign n_8089 = n_8088 ^ x77;
assign n_8090 = n_8089 ^ x78;
assign n_8091 = n_7989 ^ n_8089;
assign n_8092 = n_8090 & n_8091;
assign n_8093 = n_8092 ^ x78;
assign n_8094 = n_8093 ^ x79;
assign n_8095 = n_7990 ^ n_8093;
assign n_8096 = n_8094 & n_8095;
assign n_8097 = n_8096 ^ x79;
assign n_8098 = n_8097 ^ x80;
assign n_8099 = n_7991 ^ n_8097;
assign n_8100 = n_8098 & n_8099;
assign n_8101 = n_8100 ^ x80;
assign n_8102 = n_8101 ^ x81;
assign n_8103 = n_8101 ^ n_7976;
assign n_8104 = n_8040 & n_8101;
assign n_8105 = n_8102 & ~n_8103;
assign n_8106 = ~n_8044 & ~n_8104;
assign n_8107 = n_8105 ^ x81;
assign n_8108 = x83 ^ n_8106;
assign n_8109 = n_7992 ^ n_8106;
assign n_8110 = n_8107 ^ x82;
assign n_8111 = ~n_8108 & ~n_8109;
assign n_8112 = n_8111 ^ x83;
assign n_8113 = n_8112 ^ x84;
assign n_8114 = n_7993 ^ n_8112;
assign n_8115 = n_8113 & n_8114;
assign n_8116 = n_8115 ^ x84;
assign n_8117 = n_8116 ^ x85;
assign n_8118 = n_7994 ^ n_8116;
assign n_8119 = n_8117 & n_8118;
assign n_8120 = n_8119 ^ x85;
assign n_8121 = n_8120 ^ x86;
assign n_8122 = n_7995 ^ n_8120;
assign n_8123 = n_8121 & n_8122;
assign n_8124 = n_8123 ^ x86;
assign n_8125 = n_8124 ^ x87;
assign n_8126 = n_7996 ^ n_8124;
assign n_8127 = n_8125 & n_8126;
assign n_8128 = n_8127 ^ x87;
assign n_8129 = n_8128 ^ x88;
assign n_8130 = n_7997 ^ n_8128;
assign n_8131 = n_8129 & n_8130;
assign n_8132 = n_8131 ^ x88;
assign n_8133 = n_8132 ^ x89;
assign n_8134 = n_7998 ^ n_8132;
assign n_8135 = n_8133 & n_8134;
assign n_8136 = n_8135 ^ x89;
assign n_8137 = n_8136 ^ x90;
assign n_8138 = n_7999 ^ n_8136;
assign n_8139 = n_8137 & n_8138;
assign n_8140 = n_8139 ^ x90;
assign n_8141 = n_8140 ^ x91;
assign n_8142 = n_8000 ^ n_8140;
assign n_8143 = n_8141 & n_8142;
assign n_8144 = n_8143 ^ x91;
assign n_8145 = n_8144 ^ x92;
assign n_8146 = n_8001 ^ n_8144;
assign n_8147 = n_8145 & n_8146;
assign n_8148 = n_8147 ^ x92;
assign n_8149 = n_8148 ^ x93;
assign n_8150 = n_8002 ^ n_8148;
assign n_8151 = n_8149 & n_8150;
assign n_8152 = n_8151 ^ x93;
assign n_8153 = n_8152 ^ x94;
assign n_8154 = n_8003 ^ n_8152;
assign n_8155 = n_8153 & n_8154;
assign n_8156 = n_8155 ^ x94;
assign n_8157 = n_8156 ^ x95;
assign n_8158 = n_8004 ^ n_8156;
assign n_8159 = n_8157 & n_8158;
assign n_8160 = n_8159 ^ x95;
assign n_8161 = n_8160 ^ x96;
assign n_8162 = n_8005 ^ n_8160;
assign n_8163 = n_8161 & n_8162;
assign n_8164 = n_8163 ^ x96;
assign n_8165 = n_8164 ^ x97;
assign n_8166 = n_8006 ^ n_8164;
assign n_8167 = n_8165 & n_8166;
assign n_8168 = n_8167 ^ x97;
assign n_8169 = n_8168 ^ x98;
assign n_8170 = n_8007 ^ n_8168;
assign n_8171 = n_8169 & n_8170;
assign n_8172 = n_8171 ^ x98;
assign n_8173 = n_8172 ^ x99;
assign n_8174 = n_8008 ^ n_8172;
assign n_8175 = n_8173 & n_8174;
assign n_8176 = n_8175 ^ x99;
assign n_8177 = n_8176 ^ x100;
assign n_8178 = n_8009 ^ n_8176;
assign n_8179 = n_8177 & n_8178;
assign n_8180 = n_8179 ^ x100;
assign n_8181 = n_8180 ^ x101;
assign n_8182 = n_8010 ^ n_8180;
assign n_8183 = n_8181 & n_8182;
assign n_8184 = n_8183 ^ x101;
assign n_8185 = n_8184 ^ x102;
assign n_8186 = n_8011 ^ n_8184;
assign n_8187 = n_8185 & n_8186;
assign n_8188 = n_8187 ^ x102;
assign n_8189 = n_8188 ^ x103;
assign n_8190 = n_8012 ^ n_8188;
assign n_8191 = n_8189 & n_8190;
assign n_8192 = n_8191 ^ x103;
assign n_8193 = n_8192 ^ x104;
assign n_8194 = n_8192 ^ n_7974;
assign n_8195 = n_8038 & n_8192;
assign n_8196 = n_8193 & n_8194;
assign n_8197 = ~n_8043 & ~n_8195;
assign n_8198 = n_8196 ^ x104;
assign n_8199 = x106 ^ n_8197;
assign n_8200 = n_8013 ^ n_8197;
assign n_8201 = n_8198 ^ x105;
assign n_8202 = ~n_8199 & ~n_8200;
assign n_8203 = n_8202 ^ x106;
assign n_8204 = n_8203 ^ x107;
assign n_8205 = n_8014 ^ n_8203;
assign n_8206 = n_8204 & n_8205;
assign n_8207 = n_8206 ^ x107;
assign n_8208 = n_8207 ^ x108;
assign n_8209 = n_8015 ^ n_8207;
assign n_8210 = n_8208 & n_8209;
assign n_8211 = n_8210 ^ x108;
assign n_8212 = n_8211 ^ n_7972;
assign n_8213 = n_8211 ^ x109;
assign n_8214 = ~n_8020 & n_8212;
assign n_8215 = n_8214 ^ x109;
assign n_8216 = n_8215 ^ n_7971;
assign n_8217 = n_8215 ^ x110;
assign n_8218 = ~n_8019 & n_8216;
assign n_8219 = n_8218 ^ x110;
assign n_8220 = n_8219 ^ n_8016;
assign n_8221 = n_8016 & ~n_8219;
assign n_8222 = n_8219 ^ x111;
assign n_8223 = n_8220 ^ n_8221;
assign n_8224 = ~x111 & ~n_8223;
assign n_8225 = ~n_7916 & n_8224;
assign n_8226 = ~n_8221 & ~n_8224;
assign n_8227 = n_8224 ^ x111;
assign n_8228 = n_8225 ^ n_8226;
assign n_8229 = n_8226 & n_7611;
assign n_8230 = n_7916 & n_8226;
assign n_8231 = n_8226 ^ n_7055;
assign n_8232 = n_356 & ~n_8226;
assign n_8233 = n_8226 ^ n_359;
assign n_8234 = n_8227 ^ n_8226;
assign n_8235 = ~x112 & n_8228;
assign n_8236 = n_8232 ^ n_8233;
assign n_8237 = n_8234 ^ n_8230;
assign n_8238 = n_8226 ^ n_8235;
assign n_8239 = ~n_8231 & n_8236;
assign n_8240 = ~n_8237 & n_7922;
assign n_8241 = n_356 & ~n_8238;
assign n_8242 = n_8239 ^ n_8232;
assign n_8243 = n_8229 ^ n_8240;
assign n_8244 = n_7611 & ~n_8241;
assign n_8245 = n_8243 ^ n_8242;
assign n_8246 = n_7313 ^ n_8244;
assign n_8247 = n_8129 & n_8245;
assign n_8248 = n_8125 & n_8245;
assign n_8249 = n_8117 & n_8245;
assign n_8250 = n_8113 & n_8245;
assign n_8251 = n_8082 & n_8245;
assign n_8252 = n_8078 & n_8245;
assign n_8253 = x64 & n_8245;
assign n_8254 = n_8245 & ~n_8037;
assign n_8255 = n_8046 & n_8245;
assign n_8256 = n_8050 & n_8245;
assign n_8257 = n_8054 & n_8245;
assign n_8258 = n_8058 & n_8245;
assign n_8259 = n_8062 & n_8245;
assign n_8260 = n_8066 & n_8245;
assign n_8261 = n_8070 & n_8245;
assign n_8262 = n_8074 & n_8245;
assign n_8263 = n_8086 & n_8245;
assign n_8264 = n_8090 & n_8245;
assign n_8265 = n_8094 & n_8245;
assign n_8266 = n_8098 & n_8245;
assign n_8267 = n_8245 & n_8102;
assign n_8268 = ~n_8108 & n_8245;
assign n_8269 = n_8121 & n_8245;
assign n_8270 = n_8137 & n_8245;
assign n_8271 = n_8133 & n_8245;
assign n_8272 = n_8141 & n_8245;
assign n_8273 = n_8145 & n_8245;
assign n_8274 = n_8149 & n_8245;
assign n_8275 = n_8153 & n_8245;
assign n_8276 = n_8157 & n_8245;
assign n_8277 = n_8161 & n_8245;
assign n_8278 = n_8165 & n_8245;
assign n_8279 = n_8169 & n_8245;
assign n_8280 = n_8173 & n_8245;
assign n_8281 = n_8177 & n_8245;
assign n_8282 = n_8181 & n_8245;
assign n_8283 = n_8185 & n_8245;
assign n_8284 = n_8189 & n_8245;
assign n_8285 = n_8245 & n_8193;
assign n_8286 = ~n_8199 & n_8245;
assign n_8287 = n_8204 & n_8245;
assign n_8288 = n_8208 & n_8245;
assign n_8289 = n_8245 & n_8213;
assign n_8290 = n_8245 & n_8217;
assign n_8291 = n_8245 & n_8222;
assign y15 = n_8245;
assign n_8292 = n_8245 & n_224;
assign n_8293 = n_8245 & n_8110;
assign n_8294 = n_8245 & n_8201;
assign n_8295 = n_8247 ^ n_7997;
assign n_8296 = n_8248 ^ n_7996;
assign n_8297 = n_8249 ^ n_7994;
assign n_8298 = n_8250 ^ n_7993;
assign n_8299 = n_8251 ^ n_7987;
assign n_8300 = n_8252 ^ n_7986;
assign n_8301 = n_8253 ^ x15;
assign n_8302 = n_8254 ^ n_8029;
assign n_8303 = n_8255 ^ n_8018;
assign n_8304 = n_8256 ^ n_7979;
assign n_8305 = n_8257 ^ n_7980;
assign n_8306 = n_8258 ^ n_7981;
assign n_8307 = n_8259 ^ n_7982;
assign n_8308 = n_8260 ^ n_7983;
assign n_8309 = n_8261 ^ n_7984;
assign n_8310 = n_8262 ^ n_7985;
assign n_8311 = n_8263 ^ n_7988;
assign n_8312 = n_8264 ^ n_7989;
assign n_8313 = n_8265 ^ n_7990;
assign n_8314 = n_8266 ^ n_7991;
assign n_8315 = n_8267 ^ n_7976;
assign n_8316 = n_8268 ^ n_7992;
assign n_8317 = n_8269 ^ n_7995;
assign n_8318 = n_8270 ^ n_7999;
assign n_8319 = n_8271 ^ n_7998;
assign n_8320 = n_8272 ^ n_8000;
assign n_8321 = n_8273 ^ n_8001;
assign n_8322 = n_8274 ^ n_8002;
assign n_8323 = n_8275 ^ n_8003;
assign n_8324 = n_8276 ^ n_8004;
assign n_8325 = n_8277 ^ n_8005;
assign n_8326 = n_8278 ^ n_8006;
assign n_8327 = n_8279 ^ n_8007;
assign n_8328 = n_8280 ^ n_8008;
assign n_8329 = n_8281 ^ n_8009;
assign n_8330 = n_8282 ^ n_8010;
assign n_8331 = n_8283 ^ n_8011;
assign n_8332 = n_8284 ^ n_8012;
assign n_8333 = n_8285 ^ n_7974;
assign n_8334 = n_8286 ^ n_8013;
assign n_8335 = n_8287 ^ n_8014;
assign n_8336 = n_8288 ^ n_8015;
assign n_8337 = n_8289 ^ n_7972;
assign n_8338 = n_8290 ^ n_7971;
assign n_8339 = n_8291 ^ n_8016;
assign n_8340 = n_95 ^ n_8292;
assign n_8341 = n_7975 ^ n_8293;
assign n_8342 = n_7973 ^ n_8294;
assign n_8343 = ~x89 ^ n_8295;
assign n_8344 = n_8295 ^ x89;
assign n_8345 = n_8296 ^ x88;
assign n_8346 = x88 & ~n_8296;
assign n_8347 = n_8297 ^ x86;
assign n_8348 = n_8298 ^ x85;
assign n_8349 = ~x77 ^ n_8299;
assign n_8350 = n_8299 ^ x77;
assign n_8351 = n_8300 ^ x76;
assign n_8352 = x76 & ~n_8300;
assign n_8353 = n_8301 ^ x65;
assign n_8354 = n_29 ^ n_8301;
assign n_8355 = ~n_8301 & n_191;
assign n_8356 = n_8301 & n_283;
assign n_8357 = ~x91 ^ n_8318;
assign n_8358 = n_8318 ^ x91;
assign n_8359 = n_8319 ^ x90;
assign n_8360 = x90 & ~n_8319;
assign n_8361 = n_190 ^ n_8340;
assign n_8362 = n_8345 ^ n_8346;
assign n_8363 = n_8346 ^ n_8295;
assign n_8364 = n_8351 ^ n_8352;
assign n_8365 = n_8352 ^ n_8299;
assign n_8366 = ~n_8353 & n_228;
assign n_8367 = ~n_8353 & n_8354;
assign n_8368 = n_8359 ^ n_8360;
assign n_8369 = n_8360 ^ n_8318;
assign n_8370 = n_8361 ^ n_7930;
assign n_8371 = n_8343 & ~n_8362;
assign n_8372 = ~n_8344 & n_8363;
assign n_8373 = n_8349 & ~n_8364;
assign n_8374 = ~n_8350 & n_8365;
assign n_8375 = ~n_8366 ^ ~n_8355;
assign n_8376 = n_8367 ^ x65;
assign n_8377 = n_8357 & ~n_8368;
assign n_8378 = ~n_8358 & n_8369;
assign n_8379 = n_8370 ^ x16;
assign n_8380 = n_8372 ^ x89;
assign n_8381 = n_8374 ^ x77;
assign n_8382 = ~n_8375 ^ n_8356;
assign n_8383 = n_8376 ^ x66;
assign n_8384 = n_8378 ^ x91;
assign n_8385 = n_8379 ^ n_8376;
assign n_8386 = n_8383 & n_8385;
assign n_8387 = n_8386 ^ x66;
assign n_8388 = n_8387 ^ x67;
assign n_8389 = n_8302 ^ n_8387;
assign n_8390 = n_8388 & n_8389;
assign n_8391 = n_8390 ^ x67;
assign n_8392 = n_8391 ^ x68;
assign n_8393 = n_8303 ^ n_8391;
assign n_8394 = n_8392 & n_8393;
assign n_8395 = n_8394 ^ x68;
assign n_8396 = n_8395 ^ x69;
assign n_8397 = n_8304 ^ n_8395;
assign n_8398 = n_8396 & n_8397;
assign n_8399 = n_8398 ^ x69;
assign n_8400 = n_8399 ^ x70;
assign n_8401 = n_8305 ^ n_8399;
assign n_8402 = n_8400 & n_8401;
assign n_8403 = n_8402 ^ x70;
assign n_8404 = n_8403 ^ x71;
assign n_8405 = n_8306 ^ n_8403;
assign n_8406 = n_8404 & n_8405;
assign n_8407 = n_8406 ^ x71;
assign n_8408 = n_8407 ^ x72;
assign n_8409 = n_8307 ^ n_8407;
assign n_8410 = n_8408 & n_8409;
assign n_8411 = n_8410 ^ x72;
assign n_8412 = n_8411 ^ x73;
assign n_8413 = n_8308 ^ n_8411;
assign n_8414 = n_8412 & n_8413;
assign n_8415 = n_8414 ^ x73;
assign n_8416 = n_8415 ^ x74;
assign n_8417 = n_8309 ^ n_8415;
assign n_8418 = n_8416 & n_8417;
assign n_8419 = n_8418 ^ x74;
assign n_8420 = n_8419 ^ x75;
assign n_8421 = n_8310 ^ n_8419;
assign n_8422 = n_8420 & n_8421;
assign n_8423 = n_8422 ^ x75;
assign n_8424 = n_8423 ^ x76;
assign n_8425 = n_8423 ^ n_8300;
assign n_8426 = n_8373 & n_8423;
assign n_8427 = n_8424 & n_8425;
assign n_8428 = ~n_8381 & ~n_8426;
assign n_8429 = n_8427 ^ x76;
assign n_8430 = x78 ^ n_8428;
assign n_8431 = n_8311 ^ n_8428;
assign n_8432 = n_8429 ^ x77;
assign n_8433 = ~n_8430 & ~n_8431;
assign n_8434 = n_8433 ^ x78;
assign n_8435 = n_8434 ^ x79;
assign n_8436 = n_8312 ^ n_8434;
assign n_8437 = n_8435 & n_8436;
assign n_8438 = n_8437 ^ x79;
assign n_8439 = n_8438 ^ x80;
assign n_8440 = n_8313 ^ n_8438;
assign n_8441 = n_8439 & n_8440;
assign n_8442 = n_8441 ^ x80;
assign n_8443 = n_8442 ^ x81;
assign n_8444 = n_8314 ^ n_8442;
assign n_8445 = n_8443 & n_8444;
assign n_8446 = n_8445 ^ x81;
assign n_8447 = n_8446 ^ x82;
assign n_8448 = n_8315 ^ n_8446;
assign n_8449 = n_8447 & ~n_8448;
assign n_8450 = n_8449 ^ x82;
assign n_8451 = n_8450 ^ x83;
assign n_8452 = n_8341 ^ n_8450;
assign n_8453 = n_8451 & n_8452;
assign n_8454 = n_8453 ^ x83;
assign n_8455 = n_8454 ^ x84;
assign n_8456 = n_8316 ^ n_8454;
assign n_8457 = n_8455 & n_8456;
assign n_8458 = n_8457 ^ x84;
assign n_8459 = n_8458 ^ n_8298;
assign n_8460 = n_8458 ^ x85;
assign n_8461 = ~n_8348 & n_8459;
assign n_8462 = n_8461 ^ x85;
assign n_8463 = n_8462 ^ n_8297;
assign n_8464 = n_8462 ^ x86;
assign n_8465 = ~n_8347 & n_8463;
assign n_8466 = n_8465 ^ x86;
assign n_8467 = n_8466 ^ x87;
assign n_8468 = n_8317 ^ n_8466;
assign n_8469 = n_8467 & n_8468;
assign n_8470 = n_8469 ^ x87;
assign n_8471 = n_8470 ^ x88;
assign n_8472 = n_8470 ^ n_8296;
assign n_8473 = n_8371 & n_8470;
assign n_8474 = n_8471 & n_8472;
assign n_8475 = ~n_8380 & ~n_8473;
assign n_8476 = n_8474 ^ x88;
assign n_8477 = x90 ^ n_8475;
assign n_8478 = n_8319 ^ n_8475;
assign n_8479 = n_8377 & ~n_8475;
assign n_8480 = n_8476 ^ x89;
assign n_8481 = ~n_8477 & ~n_8478;
assign n_8482 = ~n_8384 & ~n_8479;
assign n_8483 = n_8481 ^ x90;
assign n_8484 = x92 ^ n_8482;
assign n_8485 = n_8320 ^ n_8482;
assign n_8486 = n_8483 ^ x91;
assign n_8487 = ~n_8484 & ~n_8485;
assign n_8488 = n_8487 ^ x92;
assign n_8489 = n_8488 ^ x93;
assign n_8490 = n_8321 ^ n_8488;
assign n_8491 = n_8489 & n_8490;
assign n_8492 = n_8491 ^ x93;
assign n_8493 = n_8492 ^ x94;
assign n_8494 = n_8322 ^ n_8492;
assign n_8495 = n_8493 & n_8494;
assign n_8496 = n_8495 ^ x94;
assign n_8497 = n_8496 ^ x95;
assign n_8498 = n_8323 ^ n_8496;
assign n_8499 = n_8497 & n_8498;
assign n_8500 = n_8499 ^ x95;
assign n_8501 = n_8500 ^ x96;
assign n_8502 = n_8324 ^ n_8500;
assign n_8503 = n_8501 & n_8502;
assign n_8504 = n_8503 ^ x96;
assign n_8505 = n_8504 ^ x97;
assign n_8506 = n_8325 ^ n_8504;
assign n_8507 = n_8505 & n_8506;
assign n_8508 = n_8507 ^ x97;
assign n_8509 = n_8508 ^ x98;
assign n_8510 = n_8326 ^ n_8508;
assign n_8511 = n_8509 & n_8510;
assign n_8512 = n_8511 ^ x98;
assign n_8513 = n_8512 ^ x99;
assign n_8514 = n_8327 ^ n_8512;
assign n_8515 = n_8513 & n_8514;
assign n_8516 = n_8515 ^ x99;
assign n_8517 = n_8516 ^ x100;
assign n_8518 = n_8328 ^ n_8516;
assign n_8519 = n_8517 & n_8518;
assign n_8520 = n_8519 ^ x100;
assign n_8521 = n_8520 ^ x101;
assign n_8522 = n_8329 ^ n_8520;
assign n_8523 = n_8521 & n_8522;
assign n_8524 = n_8523 ^ x101;
assign n_8525 = n_8524 ^ x102;
assign n_8526 = n_8330 ^ n_8524;
assign n_8527 = n_8525 & n_8526;
assign n_8528 = n_8527 ^ x102;
assign n_8529 = n_8528 ^ x103;
assign n_8530 = n_8331 ^ n_8528;
assign n_8531 = n_8529 & n_8530;
assign n_8532 = n_8531 ^ x103;
assign n_8533 = n_8532 ^ x104;
assign n_8534 = n_8332 ^ n_8532;
assign n_8535 = n_8533 & n_8534;
assign n_8536 = n_8535 ^ x104;
assign n_8537 = n_8536 ^ x105;
assign n_8538 = n_8333 ^ n_8536;
assign n_8539 = n_8537 & n_8538;
assign n_8540 = n_8539 ^ x105;
assign n_8541 = n_8540 ^ x106;
assign n_8542 = n_8342 ^ n_8540;
assign n_8543 = n_8541 & n_8542;
assign n_8544 = n_8543 ^ x106;
assign n_8545 = n_8544 ^ x107;
assign n_8546 = n_8334 ^ n_8544;
assign n_8547 = n_8545 & n_8546;
assign n_8548 = n_8547 ^ x107;
assign n_8549 = n_8548 ^ x108;
assign n_8550 = n_8335 ^ n_8548;
assign n_8551 = n_8549 & n_8550;
assign n_8552 = n_8551 ^ x108;
assign n_8553 = n_8552 ^ x109;
assign n_8554 = n_8336 ^ n_8552;
assign n_8555 = n_8553 & n_8554;
assign n_8556 = n_8555 ^ x109;
assign n_8557 = n_8556 ^ x110;
assign n_8558 = n_8337 ^ n_8556;
assign n_8559 = n_8557 & n_8558;
assign n_8560 = n_8559 ^ x110;
assign n_8561 = n_8560 ^ x111;
assign n_8562 = n_8338 ^ n_8560;
assign n_8563 = n_8561 & n_8562;
assign n_8564 = n_8563 ^ x111;
assign n_8565 = n_8564 ^ x112;
assign n_8566 = n_8339 ^ n_8564;
assign n_8567 = n_8565 & n_8566;
assign n_8568 = n_8567 ^ x112;
assign n_8569 = n_8568 ^ x113;
assign n_8570 = n_8568 ^ ~n_8246;
assign n_8571 = n_357 & n_8569;
assign n_8572 = ~n_8570 ^ n_7313;
assign n_8573 = ~n_8571 & n_8244;
assign n_8574 = n_8569 & n_8572;
assign n_8575 = n_8574 ^ x113;
assign n_8576 = n_357 & ~n_8575;
assign n_8577 = n_8541 & n_8576;
assign n_8578 = n_8537 & n_8576;
assign n_8579 = n_8501 & n_8576;
assign n_8580 = n_8497 & n_8576;
assign n_8581 = n_8455 & n_8576;
assign n_8582 = n_8451 & n_8576;
assign n_8583 = x64 & n_8576;
assign n_8584 = n_8301 ^ n_8576;
assign n_8585 = ~n_8301 & ~n_8576;
assign n_8586 = n_284 & n_8576;
assign n_8587 = ~x65 & n_8576;
assign n_8588 = n_8383 & n_8576;
assign n_8589 = n_8388 & n_8576;
assign n_8590 = n_8392 & n_8576;
assign n_8591 = n_8396 & n_8576;
assign n_8592 = n_8400 & n_8576;
assign n_8593 = n_8404 & n_8576;
assign n_8594 = n_8408 & n_8576;
assign n_8595 = n_8412 & n_8576;
assign n_8596 = n_8416 & n_8576;
assign n_8597 = n_8420 & n_8576;
assign n_8598 = n_8424 & n_8576;
assign n_8599 = ~n_8430 & n_8576;
assign n_8600 = n_8435 & n_8576;
assign n_8601 = n_8439 & n_8576;
assign n_8602 = n_8443 & n_8576;
assign n_8603 = n_8447 & n_8576;
assign n_8604 = n_8460 & n_8576;
assign n_8605 = n_8464 & n_8576;
assign n_8606 = n_8467 & n_8576;
assign n_8607 = n_8471 & n_8576;
assign n_8608 = ~n_8477 & n_8576;
assign n_8609 = ~n_8484 & n_8576;
assign n_8610 = n_8489 & n_8576;
assign n_8611 = n_8493 & n_8576;
assign n_8612 = n_8505 & n_8576;
assign n_8613 = n_8509 & n_8576;
assign n_8614 = n_8513 & n_8576;
assign n_8615 = n_8517 & n_8576;
assign n_8616 = n_8521 & n_8576;
assign n_8617 = n_8525 & n_8576;
assign n_8618 = n_8529 & n_8576;
assign n_8619 = n_8533 & n_8576;
assign n_8620 = n_8545 & n_8576;
assign n_8621 = n_8549 & n_8576;
assign n_8622 = n_8553 & n_8576;
assign n_8623 = n_8557 & n_8576;
assign n_8624 = n_8561 & n_8576;
assign n_8625 = n_8565 & n_8576;
assign n_8626 = n_166 & n_8576;
assign y14 = n_8576;
assign n_8627 = n_8432 & n_8576;
assign n_8628 = n_8480 & n_8576;
assign n_8629 = n_8486 & n_8576;
assign n_8630 = n_8577 ^ n_8342;
assign n_8631 = n_8578 ^ n_8333;
assign n_8632 = n_8579 ^ n_8324;
assign n_8633 = n_8580 ^ n_8323;
assign n_8634 = n_8581 ^ n_8316;
assign n_8635 = n_8582 ^ n_8341;
assign n_8636 = ~n_8583 & n_225;
assign n_8637 = n_8583 & n_310;
assign n_8638 = n_8585 & n_226;
assign n_8639 = n_282 ^ n_8586;
assign n_8640 = n_226 & ~n_8587;
assign n_8641 = n_8587 & n_167;
assign n_8642 = n_8588 ^ n_8379;
assign n_8643 = n_8589 ^ n_8302;
assign n_8644 = n_8590 ^ n_8303;
assign n_8645 = n_8591 ^ n_8304;
assign n_8646 = n_8592 ^ n_8305;
assign n_8647 = n_8593 ^ n_8306;
assign n_8648 = n_8594 ^ n_8307;
assign n_8649 = n_8595 ^ n_8308;
assign n_8650 = n_8596 ^ n_8309;
assign n_8651 = n_8597 ^ n_8310;
assign n_8652 = n_8598 ^ n_8300;
assign n_8653 = n_8599 ^ n_8311;
assign n_8654 = n_8600 ^ n_8312;
assign n_8655 = n_8601 ^ n_8313;
assign n_8656 = n_8602 ^ n_8314;
assign n_8657 = n_8603 ^ n_8315;
assign n_8658 = n_8604 ^ n_8298;
assign n_8659 = n_8605 ^ n_8297;
assign n_8660 = n_8606 ^ n_8317;
assign n_8661 = n_8607 ^ n_8296;
assign n_8662 = n_8608 ^ n_8319;
assign n_8663 = n_8609 ^ n_8320;
assign n_8664 = n_8610 ^ n_8321;
assign n_8665 = n_8611 ^ n_8322;
assign n_8666 = n_8612 ^ n_8325;
assign n_8667 = n_8613 ^ n_8326;
assign n_8668 = n_8614 ^ n_8327;
assign n_8669 = n_8615 ^ n_8328;
assign n_8670 = n_8616 ^ n_8329;
assign n_8671 = n_8617 ^ n_8330;
assign n_8672 = n_8618 ^ n_8331;
assign n_8673 = n_8619 ^ n_8332;
assign n_8674 = n_8620 ^ n_8334;
assign n_8675 = n_8621 ^ n_8335;
assign n_8676 = n_8622 ^ n_8336;
assign n_8677 = n_8623 ^ n_8337;
assign n_8678 = n_8624 ^ n_8338;
assign n_8679 = n_8625 ^ n_8339;
assign n_8680 = n_8626 ^ n_8301;
assign n_8681 = n_8299 ^ n_8627;
assign n_8682 = n_8295 ^ n_8628;
assign n_8683 = n_8318 ^ n_8629;
assign n_8684 = ~x107 ^ n_8630;
assign n_8685 = n_8630 ^ x107;
assign n_8686 = n_8631 ^ x106;
assign n_8687 = x106 & ~n_8631;
assign n_8688 = n_8632 ^ x97;
assign n_8689 = n_8633 ^ x96;
assign n_8690 = ~x85 ^ n_8634;
assign n_8691 = n_8634 ^ x85;
assign n_8692 = n_8635 ^ x84;
assign n_8693 = x84 & ~n_8635;
assign n_8694 = n_8636 & ~n_8584;
assign n_8695 = n_8637 ^ n_225;
assign n_8696 = ~x66 & ~n_8638;
assign n_8697 = ~n_8353 & n_8639;
assign n_8698 = ~n_8375 ^ n_8641;
assign n_8699 = n_8686 ^ n_8687;
assign n_8700 = n_8687 ^ n_8630;
assign n_8701 = n_8692 ^ n_8693;
assign n_8702 = n_8693 ^ n_8634;
assign n_8703 = ~n_8640 & ~n_8695;
assign n_8704 = ~n_8694 & n_8696;
assign n_8705 = n_282 ^ n_8697;
assign n_8706 = n_8698 ^ ~n_8375;
assign n_8707 = n_8684 & ~n_8699;
assign n_8708 = ~n_8685 & n_8700;
assign n_8709 = n_8690 & ~n_8701;
assign n_8710 = ~n_8691 & n_8702;
assign n_8711 = x66 ^ n_8703;
assign n_8712 = x64 & n_8705;
assign n_8713 = n_8706 ^ n_8576;
assign n_8714 = n_8708 ^ x107;
assign n_8715 = n_8710 ^ x85;
assign n_8716 = n_8704 & ~n_8712;
assign n_8717 = ~n_8382 & n_8713;
assign n_8718 = n_8356 ^ n_8717;
assign n_8719 = ~n_8718 & ~n_8716;
assign n_8720 = x67 ^ n_8719;
assign n_8721 = n_8642 ^ n_8719;
assign n_8722 = n_8720 & n_8721;
assign n_8723 = n_8722 ^ x67;
assign n_8724 = n_8723 ^ x68;
assign n_8725 = n_8643 ^ n_8723;
assign n_8726 = n_8724 & n_8725;
assign n_8727 = n_8726 ^ x68;
assign n_8728 = n_8727 ^ x69;
assign n_8729 = n_8644 ^ n_8727;
assign n_8730 = n_8728 & n_8729;
assign n_8731 = n_8730 ^ x69;
assign n_8732 = n_8731 ^ x70;
assign n_8733 = n_8645 ^ n_8731;
assign n_8734 = n_8732 & n_8733;
assign n_8735 = n_8734 ^ x70;
assign n_8736 = n_8735 ^ x71;
assign n_8737 = n_8646 ^ n_8735;
assign n_8738 = n_8736 & n_8737;
assign n_8739 = n_8738 ^ x71;
assign n_8740 = n_8739 ^ x72;
assign n_8741 = n_8647 ^ n_8739;
assign n_8742 = n_8740 & n_8741;
assign n_8743 = n_8742 ^ x72;
assign n_8744 = n_8743 ^ x73;
assign n_8745 = n_8648 ^ n_8743;
assign n_8746 = n_8744 & n_8745;
assign n_8747 = n_8746 ^ x73;
assign n_8748 = n_8747 ^ x74;
assign n_8749 = n_8649 ^ n_8747;
assign n_8750 = n_8748 & n_8749;
assign n_8751 = n_8750 ^ x74;
assign n_8752 = n_8751 ^ x75;
assign n_8753 = n_8650 ^ n_8751;
assign n_8754 = n_8752 & n_8753;
assign n_8755 = n_8754 ^ x75;
assign n_8756 = n_8755 ^ x76;
assign n_8757 = n_8651 ^ n_8755;
assign n_8758 = n_8756 & n_8757;
assign n_8759 = n_8758 ^ x76;
assign n_8760 = n_8759 ^ x77;
assign n_8761 = n_8652 ^ n_8759;
assign n_8762 = n_8760 & n_8761;
assign n_8763 = n_8762 ^ x77;
assign n_8764 = n_8763 ^ x78;
assign n_8765 = n_8681 ^ n_8763;
assign n_8766 = n_8764 & n_8765;
assign n_8767 = n_8766 ^ x78;
assign n_8768 = n_8767 ^ x79;
assign n_8769 = n_8653 ^ n_8767;
assign n_8770 = n_8768 & n_8769;
assign n_8771 = n_8770 ^ x79;
assign n_8772 = n_8771 ^ x80;
assign n_8773 = n_8654 ^ n_8771;
assign n_8774 = n_8772 & n_8773;
assign n_8775 = n_8774 ^ x80;
assign n_8776 = n_8775 ^ x81;
assign n_8777 = n_8655 ^ n_8775;
assign n_8778 = n_8776 & n_8777;
assign n_8779 = n_8778 ^ x81;
assign n_8780 = n_8779 ^ x82;
assign n_8781 = n_8656 ^ n_8779;
assign n_8782 = n_8780 & n_8781;
assign n_8783 = n_8782 ^ x82;
assign n_8784 = n_8783 ^ x83;
assign n_8785 = n_8657 ^ n_8783;
assign n_8786 = n_8784 & ~n_8785;
assign n_8787 = n_8786 ^ x83;
assign n_8788 = n_8787 ^ x84;
assign n_8789 = n_8787 ^ n_8635;
assign n_8790 = n_8709 & n_8787;
assign n_8791 = n_8788 & n_8789;
assign n_8792 = ~n_8715 & ~n_8790;
assign n_8793 = n_8791 ^ x84;
assign n_8794 = x86 ^ n_8792;
assign n_8795 = n_8658 ^ n_8792;
assign n_8796 = n_8793 ^ x85;
assign n_8797 = ~n_8794 & ~n_8795;
assign n_8798 = n_8797 ^ x86;
assign n_8799 = n_8798 ^ x87;
assign n_8800 = n_8659 ^ n_8798;
assign n_8801 = n_8799 & n_8800;
assign n_8802 = n_8801 ^ x87;
assign n_8803 = n_8802 ^ x88;
assign n_8804 = n_8660 ^ n_8802;
assign n_8805 = n_8803 & n_8804;
assign n_8806 = n_8805 ^ x88;
assign n_8807 = n_8806 ^ x89;
assign n_8808 = n_8661 ^ n_8806;
assign n_8809 = n_8807 & n_8808;
assign n_8810 = n_8809 ^ x89;
assign n_8811 = n_8810 ^ x90;
assign n_8812 = n_8682 ^ n_8810;
assign n_8813 = n_8811 & n_8812;
assign n_8814 = n_8813 ^ x90;
assign n_8815 = n_8814 ^ x91;
assign n_8816 = n_8662 ^ n_8814;
assign n_8817 = n_8815 & n_8816;
assign n_8818 = n_8817 ^ x91;
assign n_8819 = n_8818 ^ x92;
assign n_8820 = n_8683 ^ n_8818;
assign n_8821 = n_8819 & n_8820;
assign n_8822 = n_8821 ^ x92;
assign n_8823 = n_8822 ^ x93;
assign n_8824 = n_8663 ^ n_8822;
assign n_8825 = n_8823 & n_8824;
assign n_8826 = n_8825 ^ x93;
assign n_8827 = n_8826 ^ x94;
assign n_8828 = n_8664 ^ n_8826;
assign n_8829 = n_8827 & n_8828;
assign n_8830 = n_8829 ^ x94;
assign n_8831 = n_8830 ^ x95;
assign n_8832 = n_8665 ^ n_8830;
assign n_8833 = n_8831 & n_8832;
assign n_8834 = n_8833 ^ x95;
assign n_8835 = n_8834 ^ n_8633;
assign n_8836 = n_8834 ^ x96;
assign n_8837 = ~n_8689 & n_8835;
assign n_8838 = n_8837 ^ x96;
assign n_8839 = n_8838 ^ n_8632;
assign n_8840 = n_8838 ^ x97;
assign n_8841 = ~n_8688 & n_8839;
assign n_8842 = n_8841 ^ x97;
assign n_8843 = n_8842 ^ x98;
assign n_8844 = n_8666 ^ n_8842;
assign n_8845 = n_8843 & n_8844;
assign n_8846 = n_8845 ^ x98;
assign n_8847 = n_8846 ^ x99;
assign n_8848 = n_8667 ^ n_8846;
assign n_8849 = n_8847 & n_8848;
assign n_8850 = n_8849 ^ x99;
assign n_8851 = n_8850 ^ x100;
assign n_8852 = n_8668 ^ n_8850;
assign n_8853 = n_8851 & n_8852;
assign n_8854 = n_8853 ^ x100;
assign n_8855 = n_8854 ^ x101;
assign n_8856 = n_8669 ^ n_8854;
assign n_8857 = n_8855 & n_8856;
assign n_8858 = n_8857 ^ x101;
assign n_8859 = n_8858 ^ x102;
assign n_8860 = n_8670 ^ n_8858;
assign n_8861 = n_8859 & n_8860;
assign n_8862 = n_8861 ^ x102;
assign n_8863 = n_8862 ^ x103;
assign n_8864 = n_8671 ^ n_8862;
assign n_8865 = n_8863 & n_8864;
assign n_8866 = n_8865 ^ x103;
assign n_8867 = n_8866 ^ x104;
assign n_8868 = n_8672 ^ n_8866;
assign n_8869 = n_8867 & n_8868;
assign n_8870 = n_8869 ^ x104;
assign n_8871 = n_8870 ^ x105;
assign n_8872 = n_8673 ^ n_8870;
assign n_8873 = n_8871 & n_8872;
assign n_8874 = n_8873 ^ x105;
assign n_8875 = n_8874 ^ x106;
assign n_8876 = n_8874 ^ n_8631;
assign n_8877 = n_8707 & n_8874;
assign n_8878 = n_8875 & n_8876;
assign n_8879 = ~n_8714 & ~n_8877;
assign n_8880 = n_8878 ^ x106;
assign n_8881 = x108 ^ n_8879;
assign n_8882 = n_8674 ^ n_8879;
assign n_8883 = n_8880 ^ x107;
assign n_8884 = ~n_8881 & ~n_8882;
assign n_8885 = n_8884 ^ x108;
assign n_8886 = n_8885 ^ x109;
assign n_8887 = n_8675 ^ n_8885;
assign n_8888 = n_8886 & n_8887;
assign n_8889 = n_8888 ^ x109;
assign n_8890 = n_8889 ^ x110;
assign n_8891 = n_8676 ^ n_8889;
assign n_8892 = n_8890 & n_8891;
assign n_8893 = n_8892 ^ x110;
assign n_8894 = n_8893 ^ x111;
assign n_8895 = n_8677 ^ n_8893;
assign n_8896 = n_8894 & n_8895;
assign n_8897 = n_8896 ^ x111;
assign n_8898 = n_8897 ^ x112;
assign n_8899 = n_8678 ^ n_8897;
assign n_8900 = n_8898 & n_8899;
assign n_8901 = n_8900 ^ x112;
assign n_8902 = n_8901 ^ x113;
assign n_8903 = n_8679 ^ n_8901;
assign n_8904 = n_8902 & n_8903;
assign n_8905 = n_8904 ^ x113;
assign n_8906 = n_8905 ^ x114;
assign n_8907 = n_8905 ^ n_8573;
assign n_8908 = n_355 & n_8906;
assign n_8909 = n_8906 & n_8907;
assign n_8910 = ~n_8908 & n_8573;
assign n_8911 = n_8909 ^ x114;
assign n_8912 = ~x115 ^ n_8910;
assign n_8913 = x115 ^ n_8910;
assign n_8914 = n_355 & ~n_8911;
assign n_8915 = n_8902 & n_8914;
assign n_8916 = n_8851 & n_8914;
assign n_8917 = n_8847 & n_8914;
assign n_8918 = n_8752 & n_8914;
assign n_8919 = n_8748 & n_8914;
assign n_8920 = n_31 & n_8914;
assign n_8921 = x65 & n_8914;
assign n_8922 = x64 & n_8914;
assign n_8923 = n_8720 & n_8914;
assign n_8924 = n_8724 & n_8914;
assign n_8925 = n_8728 & n_8914;
assign n_8926 = n_8732 & n_8914;
assign n_8927 = n_8736 & n_8914;
assign n_8928 = n_8740 & n_8914;
assign n_8929 = n_8744 & n_8914;
assign n_8930 = n_8756 & n_8914;
assign n_8931 = n_8760 & n_8914;
assign n_8932 = n_8764 & n_8914;
assign n_8933 = n_8768 & n_8914;
assign n_8934 = n_8772 & n_8914;
assign n_8935 = n_8776 & n_8914;
assign n_8936 = n_8780 & n_8914;
assign n_8937 = n_8784 & n_8914;
assign n_8938 = n_8788 & n_8914;
assign n_8939 = ~n_8794 & n_8914;
assign n_8940 = n_8799 & n_8914;
assign n_8941 = n_8803 & n_8914;
assign n_8942 = n_8807 & n_8914;
assign n_8943 = n_8811 & n_8914;
assign n_8944 = n_8815 & n_8914;
assign n_8945 = n_8819 & n_8914;
assign n_8946 = n_8823 & n_8914;
assign n_8947 = n_8827 & n_8914;
assign n_8948 = n_8831 & n_8914;
assign n_8949 = n_8836 & n_8914;
assign n_8950 = n_8840 & n_8914;
assign n_8951 = n_8843 & n_8914;
assign n_8952 = n_8855 & n_8914;
assign n_8953 = n_8859 & n_8914;
assign n_8954 = n_8863 & n_8914;
assign n_8955 = n_8867 & n_8914;
assign n_8956 = n_8871 & n_8914;
assign n_8957 = n_8875 & n_8914;
assign n_8958 = ~n_8881 & n_8914;
assign n_8959 = n_8886 & n_8914;
assign n_8960 = n_8890 & n_8914;
assign n_8961 = n_8894 & n_8914;
assign n_8962 = n_8898 & n_8914;
assign y13 = n_8914;
assign n_8963 = ~n_8711 & n_8914;
assign n_8964 = n_8796 & n_8914;
assign n_8965 = n_8883 & n_8914;
assign n_8966 = n_8915 ^ n_8679;
assign n_8967 = n_8916 ^ n_8668;
assign n_8968 = n_8917 ^ n_8667;
assign n_8969 = n_8918 ^ n_8650;
assign n_8970 = n_8919 ^ n_8649;
assign n_8971 = n_8920 ^ n_8583;
assign n_8972 = n_8921 ^ x14;
assign n_8973 = x65 & n_8922;
assign n_8974 = n_8922 ^ n_31;
assign n_8975 = n_8923 ^ n_8642;
assign n_8976 = n_8924 ^ n_8643;
assign n_8977 = n_8925 ^ n_8644;
assign n_8978 = n_8926 ^ n_8645;
assign n_8979 = n_8927 ^ n_8646;
assign n_8980 = n_8928 ^ n_8647;
assign n_8981 = n_8929 ^ n_8648;
assign n_8982 = n_8930 ^ n_8651;
assign n_8983 = n_8931 ^ n_8652;
assign n_8984 = n_8932 ^ n_8681;
assign n_8985 = n_8933 ^ n_8653;
assign n_8986 = n_8934 ^ n_8654;
assign n_8987 = n_8935 ^ n_8655;
assign n_8988 = n_8936 ^ n_8656;
assign n_8989 = n_8937 ^ n_8657;
assign n_8990 = n_8938 ^ n_8635;
assign n_8991 = n_8939 ^ n_8658;
assign n_8992 = n_8940 ^ n_8659;
assign n_8993 = n_8941 ^ n_8660;
assign n_8994 = n_8942 ^ n_8661;
assign n_8995 = n_8943 ^ n_8682;
assign n_8996 = n_8944 ^ n_8662;
assign n_8997 = n_8945 ^ n_8683;
assign n_8998 = n_8946 ^ n_8663;
assign n_8999 = n_8947 ^ n_8664;
assign n_9000 = n_8948 ^ n_8665;
assign n_9001 = n_8949 ^ n_8633;
assign n_9002 = n_8950 ^ n_8632;
assign n_9003 = n_8951 ^ n_8666;
assign n_9004 = n_8952 ^ n_8669;
assign n_9005 = n_8953 ^ n_8670;
assign n_9006 = n_8954 ^ n_8671;
assign n_9007 = n_8955 ^ n_8672;
assign n_9008 = n_8956 ^ n_8673;
assign n_9009 = n_8957 ^ n_8631;
assign n_9010 = n_8958 ^ n_8674;
assign n_9011 = n_8959 ^ n_8675;
assign n_9012 = n_8960 ^ n_8676;
assign n_9013 = n_8961 ^ n_8677;
assign n_9014 = n_8962 ^ n_8678;
assign n_9015 = n_8680 ^ n_8963;
assign n_9016 = n_8634 ^ n_8964;
assign n_9017 = n_8630 ^ n_8965;
assign n_9018 = n_8966 ^ x114;
assign n_9019 = x114 & ~n_8966;
assign n_9020 = ~x101 ^ n_8967;
assign n_9021 = n_8967 ^ x101;
assign n_9022 = n_8968 ^ x100;
assign n_9023 = x100 & ~n_8968;
assign n_9024 = ~x76 ^ n_8969;
assign n_9025 = n_8969 ^ x76;
assign n_9026 = n_8970 ^ x75;
assign n_9027 = x75 & ~n_8970;
assign n_9028 = n_8971 ^ n_8972;
assign n_9029 = n_229 ^ n_8973;
assign n_9030 = ~x12 & n_8974;
assign n_9031 = n_9018 ^ n_9019;
assign n_9032 = n_9019 ^ x115;
assign n_9033 = n_9022 ^ n_9023;
assign n_9034 = n_9023 ^ n_8967;
assign n_9035 = n_9026 ^ n_9027;
assign n_9036 = n_9027 ^ n_8969;
assign n_9037 = n_9028 ^ x66;
assign n_9038 = n_9029 ^ n_9030;
assign n_9039 = n_8912 & ~n_9031;
assign n_9040 = ~n_8913 & n_9032;
assign n_9041 = n_9020 & ~n_9033;
assign n_9042 = ~n_9021 & n_9034;
assign n_9043 = n_9024 & ~n_9035;
assign n_9044 = ~n_9025 & n_9036;
assign n_9045 = n_9038 ^ n_98;
assign n_9046 = n_9040 ^ x115;
assign n_9047 = n_9042 ^ x101;
assign n_9048 = n_9044 ^ x76;
assign n_9049 = n_9045 ^ n_9028;
assign n_9050 = n_9045 ^ x66;
assign n_9051 = ~n_9046 & n_354;
assign n_9052 = ~n_9037 & n_9049;
assign n_9053 = n_9052 ^ x66;
assign n_9054 = n_9053 ^ x67;
assign n_9055 = n_9015 ^ n_9053;
assign n_9056 = n_9054 & n_9055;
assign n_9057 = n_9056 ^ x67;
assign n_9058 = n_9057 ^ x68;
assign n_9059 = n_8975 ^ n_9057;
assign n_9060 = n_9058 & n_9059;
assign n_9061 = n_9060 ^ x68;
assign n_9062 = n_9061 ^ x69;
assign n_9063 = n_8976 ^ n_9061;
assign n_9064 = n_9062 & n_9063;
assign n_9065 = n_9064 ^ x69;
assign n_9066 = n_9065 ^ x70;
assign n_9067 = n_8977 ^ n_9065;
assign n_9068 = n_9066 & n_9067;
assign n_9069 = n_9068 ^ x70;
assign n_9070 = n_9069 ^ x71;
assign n_9071 = n_8978 ^ n_9069;
assign n_9072 = n_9070 & n_9071;
assign n_9073 = n_9072 ^ x71;
assign n_9074 = n_9073 ^ x72;
assign n_9075 = n_8979 ^ n_9073;
assign n_9076 = n_9074 & n_9075;
assign n_9077 = n_9076 ^ x72;
assign n_9078 = n_9077 ^ x73;
assign n_9079 = n_8980 ^ n_9077;
assign n_9080 = n_9078 & n_9079;
assign n_9081 = n_9080 ^ x73;
assign n_9082 = n_9081 ^ x74;
assign n_9083 = n_8981 ^ n_9081;
assign n_9084 = n_9082 & n_9083;
assign n_9085 = n_9084 ^ x74;
assign n_9086 = n_9085 ^ x75;
assign n_9087 = n_9085 ^ n_8970;
assign n_9088 = n_9043 & n_9085;
assign n_9089 = n_9086 & n_9087;
assign n_9090 = ~n_9048 & ~n_9088;
assign n_9091 = n_9089 ^ x75;
assign n_9092 = x77 ^ n_9090;
assign n_9093 = n_8982 ^ n_9090;
assign n_9094 = n_9091 ^ x76;
assign n_9095 = ~n_9092 & ~n_9093;
assign n_9096 = n_9095 ^ x77;
assign n_9097 = n_9096 ^ x78;
assign n_9098 = n_8983 ^ n_9096;
assign n_9099 = n_9097 & n_9098;
assign n_9100 = n_9099 ^ x78;
assign n_9101 = n_9100 ^ x79;
assign n_9102 = n_8984 ^ n_9100;
assign n_9103 = n_9101 & n_9102;
assign n_9104 = n_9103 ^ x79;
assign n_9105 = n_9104 ^ x80;
assign n_9106 = n_8985 ^ n_9104;
assign n_9107 = n_9105 & n_9106;
assign n_9108 = n_9107 ^ x80;
assign n_9109 = n_9108 ^ x81;
assign n_9110 = n_8986 ^ n_9108;
assign n_9111 = n_9109 & n_9110;
assign n_9112 = n_9111 ^ x81;
assign n_9113 = n_9112 ^ x82;
assign n_9114 = n_8987 ^ n_9112;
assign n_9115 = n_9113 & n_9114;
assign n_9116 = n_9115 ^ x82;
assign n_9117 = n_9116 ^ x83;
assign n_9118 = n_8988 ^ n_9116;
assign n_9119 = n_9117 & n_9118;
assign n_9120 = n_9119 ^ x83;
assign n_9121 = n_9120 ^ x84;
assign n_9122 = n_8989 ^ n_9120;
assign n_9123 = n_9121 & ~n_9122;
assign n_9124 = n_9123 ^ x84;
assign n_9125 = n_9124 ^ x85;
assign n_9126 = n_8990 ^ n_9124;
assign n_9127 = n_9125 & n_9126;
assign n_9128 = n_9127 ^ x85;
assign n_9129 = n_9128 ^ x86;
assign n_9130 = n_9016 ^ n_9128;
assign n_9131 = n_9129 & n_9130;
assign n_9132 = n_9131 ^ x86;
assign n_9133 = n_9132 ^ x87;
assign n_9134 = n_8991 ^ n_9132;
assign n_9135 = n_9133 & n_9134;
assign n_9136 = n_9135 ^ x87;
assign n_9137 = n_9136 ^ x88;
assign n_9138 = n_8992 ^ n_9136;
assign n_9139 = n_9137 & n_9138;
assign n_9140 = n_9139 ^ x88;
assign n_9141 = n_9140 ^ x89;
assign n_9142 = n_8993 ^ n_9140;
assign n_9143 = n_9141 & n_9142;
assign n_9144 = n_9143 ^ x89;
assign n_9145 = n_9144 ^ x90;
assign n_9146 = n_8994 ^ n_9144;
assign n_9147 = n_9145 & n_9146;
assign n_9148 = n_9147 ^ x90;
assign n_9149 = n_9148 ^ x91;
assign n_9150 = n_8995 ^ n_9148;
assign n_9151 = n_9149 & n_9150;
assign n_9152 = n_9151 ^ x91;
assign n_9153 = n_9152 ^ x92;
assign n_9154 = n_8996 ^ n_9152;
assign n_9155 = n_9153 & n_9154;
assign n_9156 = n_9155 ^ x92;
assign n_9157 = n_9156 ^ x93;
assign n_9158 = n_8997 ^ n_9156;
assign n_9159 = n_9157 & n_9158;
assign n_9160 = n_9159 ^ x93;
assign n_9161 = n_9160 ^ x94;
assign n_9162 = n_8998 ^ n_9160;
assign n_9163 = n_9161 & n_9162;
assign n_9164 = n_9163 ^ x94;
assign n_9165 = n_9164 ^ x95;
assign n_9166 = n_8999 ^ n_9164;
assign n_9167 = n_9165 & n_9166;
assign n_9168 = n_9167 ^ x95;
assign n_9169 = n_9168 ^ x96;
assign n_9170 = n_9000 ^ n_9168;
assign n_9171 = n_9169 & n_9170;
assign n_9172 = n_9171 ^ x96;
assign n_9173 = n_9172 ^ x97;
assign n_9174 = n_9001 ^ n_9172;
assign n_9175 = n_9173 & n_9174;
assign n_9176 = n_9175 ^ x97;
assign n_9177 = n_9176 ^ x98;
assign n_9178 = n_9002 ^ n_9176;
assign n_9179 = n_9177 & n_9178;
assign n_9180 = n_9179 ^ x98;
assign n_9181 = n_9180 ^ x99;
assign n_9182 = n_9003 ^ n_9180;
assign n_9183 = n_9181 & n_9182;
assign n_9184 = n_9183 ^ x99;
assign n_9185 = n_9184 ^ x100;
assign n_9186 = n_9184 ^ n_8968;
assign n_9187 = n_9041 & n_9184;
assign n_9188 = n_9185 & n_9186;
assign n_9189 = ~n_9047 & ~n_9187;
assign n_9190 = n_9188 ^ x100;
assign n_9191 = x102 ^ n_9189;
assign n_9192 = n_9004 ^ n_9189;
assign n_9193 = n_9190 ^ x101;
assign n_9194 = ~n_9191 & ~n_9192;
assign n_9195 = n_9194 ^ x102;
assign n_9196 = n_9195 ^ x103;
assign n_9197 = n_9005 ^ n_9195;
assign n_9198 = n_9196 & n_9197;
assign n_9199 = n_9198 ^ x103;
assign n_9200 = n_9199 ^ x104;
assign n_9201 = n_9006 ^ n_9199;
assign n_9202 = n_9200 & n_9201;
assign n_9203 = n_9202 ^ x104;
assign n_9204 = n_9203 ^ x105;
assign n_9205 = n_9007 ^ n_9203;
assign n_9206 = n_9204 & n_9205;
assign n_9207 = n_9206 ^ x105;
assign n_9208 = n_9207 ^ x106;
assign n_9209 = n_9008 ^ n_9207;
assign n_9210 = n_9208 & n_9209;
assign n_9211 = n_9210 ^ x106;
assign n_9212 = n_9211 ^ x107;
assign n_9213 = n_9009 ^ n_9211;
assign n_9214 = n_9212 & n_9213;
assign n_9215 = n_9214 ^ x107;
assign n_9216 = n_9215 ^ x108;
assign n_9217 = n_9017 ^ n_9215;
assign n_9218 = n_9216 & n_9217;
assign n_9219 = n_9218 ^ x108;
assign n_9220 = n_9219 ^ x109;
assign n_9221 = n_9010 ^ n_9219;
assign n_9222 = n_9220 & n_9221;
assign n_9223 = n_9222 ^ x109;
assign n_9224 = n_9223 ^ x110;
assign n_9225 = n_9011 ^ n_9223;
assign n_9226 = n_9224 & n_9225;
assign n_9227 = n_9226 ^ x110;
assign n_9228 = n_9227 ^ x111;
assign n_9229 = n_9012 ^ n_9227;
assign n_9230 = n_9228 & n_9229;
assign n_9231 = n_9230 ^ x111;
assign n_9232 = n_9231 ^ x112;
assign n_9233 = n_9013 ^ n_9231;
assign n_9234 = n_9232 & n_9233;
assign n_9235 = n_9234 ^ x112;
assign n_9236 = n_9235 ^ x113;
assign n_9237 = n_9014 ^ n_9235;
assign n_9238 = n_9236 & n_9237;
assign n_9239 = n_9238 ^ x113;
assign n_9240 = n_9239 ^ x114;
assign n_9241 = n_9239 ^ n_8966;
assign n_9242 = n_9039 & n_9239;
assign n_9243 = n_9240 & n_9241;
assign n_9244 = ~n_9242 & n_9051;
assign n_9245 = n_9243 ^ x114;
assign n_9246 = n_9185 & n_9244;
assign n_9247 = n_9181 & n_9244;
assign n_9248 = n_9097 & n_9244;
assign n_9249 = ~n_9092 & n_9244;
assign n_9250 = n_9074 & n_9244;
assign n_9251 = n_9070 & n_9244;
assign n_9252 = x65 ^ n_9244;
assign n_9253 = n_9050 & n_9244;
assign n_9254 = n_9054 & n_9244;
assign n_9255 = n_9058 & n_9244;
assign n_9256 = n_9062 & n_9244;
assign n_9257 = n_9066 & n_9244;
assign n_9258 = n_9078 & n_9244;
assign n_9259 = n_9082 & n_9244;
assign n_9260 = n_9086 & n_9244;
assign n_9261 = n_9101 & n_9244;
assign n_9262 = n_9105 & n_9244;
assign n_9263 = n_9109 & n_9244;
assign n_9264 = n_9113 & n_9244;
assign n_9265 = n_9117 & n_9244;
assign n_9266 = n_9121 & n_9244;
assign n_9267 = n_9125 & n_9244;
assign n_9268 = n_9129 & n_9244;
assign n_9269 = n_9133 & n_9244;
assign n_9270 = n_9137 & n_9244;
assign n_9271 = n_9141 & n_9244;
assign n_9272 = n_9145 & n_9244;
assign n_9273 = n_9149 & n_9244;
assign n_9274 = n_9153 & n_9244;
assign n_9275 = n_9157 & n_9244;
assign n_9276 = n_9161 & n_9244;
assign n_9277 = n_9165 & n_9244;
assign n_9278 = n_9169 & n_9244;
assign n_9279 = n_9173 & n_9244;
assign n_9280 = n_9177 & n_9244;
assign n_9281 = ~n_9191 & n_9244;
assign n_9282 = n_9196 & n_9244;
assign n_9283 = n_9200 & n_9244;
assign n_9284 = n_9204 & n_9244;
assign n_9285 = n_9208 & n_9244;
assign n_9286 = n_9212 & n_9244;
assign n_9287 = n_9216 & n_9244;
assign n_9288 = n_9220 & n_9244;
assign n_9289 = n_9224 & n_9244;
assign n_9290 = n_9228 & n_9244;
assign n_9291 = n_9232 & n_9244;
assign n_9292 = n_9236 & n_9244;
assign n_9293 = n_9240 & n_9244;
assign y12 = n_9244;
assign n_9294 = n_168 & n_9244;
assign n_9295 = n_9094 & n_9244;
assign n_9296 = n_9193 & n_9244;
assign n_9297 = n_9245 ^ x115;
assign n_9298 = n_9246 ^ n_8968;
assign n_9299 = n_9247 ^ n_9003;
assign n_9300 = n_9248 ^ n_8983;
assign n_9301 = n_9249 ^ n_8982;
assign n_9302 = n_9250 ^ n_8979;
assign n_9303 = n_9251 ^ n_8978;
assign n_9304 = x64 & n_9252;
assign n_9305 = n_9252 ^ x12;
assign n_9306 = n_9253 ^ n_9028;
assign n_9307 = n_9254 ^ n_9015;
assign n_9308 = n_9255 ^ n_8975;
assign n_9309 = n_9256 ^ n_8976;
assign n_9310 = n_9257 ^ n_8977;
assign n_9311 = n_9258 ^ n_8980;
assign n_9312 = n_9259 ^ n_8981;
assign n_9313 = n_9260 ^ n_8970;
assign n_9314 = n_9261 ^ n_8984;
assign n_9315 = n_9262 ^ n_8985;
assign n_9316 = n_9263 ^ n_8986;
assign n_9317 = n_9264 ^ n_8987;
assign n_9318 = n_9265 ^ n_8988;
assign n_9319 = n_9266 ^ n_8989;
assign n_9320 = n_9267 ^ n_8990;
assign n_9321 = n_9268 ^ n_9016;
assign n_9322 = n_9269 ^ n_8991;
assign n_9323 = n_9270 ^ n_8992;
assign n_9324 = n_9271 ^ n_8993;
assign n_9325 = n_9272 ^ n_8994;
assign n_9326 = n_9273 ^ n_8995;
assign n_9327 = n_9274 ^ n_8996;
assign n_9328 = n_9275 ^ n_8997;
assign n_9329 = n_9276 ^ n_8998;
assign n_9330 = n_9277 ^ n_8999;
assign n_9331 = n_9278 ^ n_9000;
assign n_9332 = n_9279 ^ n_9001;
assign n_9333 = n_9280 ^ n_9002;
assign n_9334 = n_9281 ^ n_9004;
assign n_9335 = n_9282 ^ n_9005;
assign n_9336 = n_9283 ^ n_9006;
assign n_9337 = n_9284 ^ n_9007;
assign n_9338 = n_9285 ^ n_9008;
assign n_9339 = n_9286 ^ n_9009;
assign n_9340 = n_9287 ^ n_9017;
assign n_9341 = n_9288 ^ n_9010;
assign n_9342 = n_9289 ^ n_9011;
assign n_9343 = n_9290 ^ n_9012;
assign n_9344 = n_9291 ^ n_9013;
assign n_9345 = n_9292 ^ n_9014;
assign n_9346 = n_9293 ^ n_8966;
assign n_9347 = n_8922 ^ n_9294;
assign n_9348 = n_8969 ^ n_9295;
assign n_9349 = n_8967 ^ n_9296;
assign n_9350 = ~n_9297 & n_8910;
assign n_9351 = ~x101 ^ n_9298;
assign n_9352 = n_9298 ^ x101;
assign n_9353 = n_9299 ^ x100;
assign n_9354 = x100 & ~n_9299;
assign n_9355 = ~x79 ^ n_9300;
assign n_9356 = n_9300 ^ x79;
assign n_9357 = n_9301 ^ x78;
assign n_9358 = x78 & ~n_9301;
assign n_9359 = n_9302 ^ x73;
assign n_9360 = n_9303 ^ x72;
assign n_9361 = n_9304 ^ x64;
assign n_9362 = n_9304 ^ n_186;
assign n_9363 = n_33 & ~n_9305;
assign n_9364 = n_9346 ^ x115;
assign n_9365 = ~x115 & n_9346;
assign n_9366 = n_9347 ^ x13;
assign n_9367 = n_9348 ^ x77;
assign n_9368 = n_9353 ^ n_9354;
assign n_9369 = n_9354 ^ n_9298;
assign n_9370 = n_9357 ^ n_9358;
assign n_9371 = n_9358 ^ n_9300;
assign n_9372 = n_9361 & n_9244;
assign n_9373 = n_9364 ^ n_9365;
assign n_9374 = ~n_9365 ^ ~n_9350;
assign n_9375 = n_9366 ^ x66;
assign n_9376 = n_9351 & ~n_9368;
assign n_9377 = ~n_9352 & n_9369;
assign n_9378 = n_9355 & ~n_9370;
assign n_9379 = ~n_9356 & n_9371;
assign n_9380 = n_9372 ^ n_99;
assign n_9381 = n_9377 ^ x101;
assign n_9382 = n_9379 ^ x79;
assign n_9383 = n_9380 ^ n_9363;
assign n_9384 = n_9383 ^ n_9366;
assign n_9385 = n_9383 ^ x66;
assign n_9386 = ~n_9375 & n_9384;
assign n_9387 = n_9386 ^ x66;
assign n_9388 = n_9387 ^ x67;
assign n_9389 = n_9306 ^ n_9387;
assign n_9390 = n_9388 & n_9389;
assign n_9391 = n_9390 ^ x67;
assign n_9392 = n_9391 ^ x68;
assign n_9393 = n_9307 ^ n_9391;
assign n_9394 = n_9392 & n_9393;
assign n_9395 = n_9394 ^ x68;
assign n_9396 = n_9395 ^ x69;
assign n_9397 = n_9308 ^ n_9395;
assign n_9398 = n_9396 & n_9397;
assign n_9399 = n_9398 ^ x69;
assign n_9400 = n_9399 ^ x70;
assign n_9401 = n_9309 ^ n_9399;
assign n_9402 = n_9400 & n_9401;
assign n_9403 = n_9402 ^ x70;
assign n_9404 = n_9403 ^ x71;
assign n_9405 = n_9310 ^ n_9403;
assign n_9406 = n_9404 & n_9405;
assign n_9407 = n_9406 ^ x71;
assign n_9408 = n_9407 ^ n_9303;
assign n_9409 = n_9407 ^ x72;
assign n_9410 = ~n_9360 & n_9408;
assign n_9411 = n_9410 ^ x72;
assign n_9412 = n_9411 ^ n_9302;
assign n_9413 = n_9411 ^ x73;
assign n_9414 = ~n_9359 & n_9412;
assign n_9415 = n_9414 ^ x73;
assign n_9416 = n_9415 ^ x74;
assign n_9417 = n_9311 ^ n_9415;
assign n_9418 = n_9416 & n_9417;
assign n_9419 = n_9418 ^ x74;
assign n_9420 = n_9419 ^ x75;
assign n_9421 = n_9312 ^ n_9419;
assign n_9422 = n_9420 & n_9421;
assign n_9423 = n_9422 ^ x75;
assign n_9424 = n_9423 ^ x76;
assign n_9425 = n_9313 ^ n_9423;
assign n_9426 = n_9424 & n_9425;
assign n_9427 = n_9426 ^ x76;
assign n_9428 = n_9427 ^ n_9348;
assign n_9429 = n_9427 ^ x77;
assign n_9430 = n_9428 & ~n_9367;
assign n_9431 = n_9430 ^ x77;
assign n_9432 = n_9431 ^ x78;
assign n_9433 = n_9431 ^ n_9301;
assign n_9434 = n_9378 & n_9431;
assign n_9435 = n_9432 & n_9433;
assign n_9436 = ~n_9382 & ~n_9434;
assign n_9437 = n_9435 ^ x78;
assign n_9438 = x80 ^ n_9436;
assign n_9439 = n_9314 ^ n_9436;
assign n_9440 = n_9437 ^ x79;
assign n_9441 = ~n_9438 & ~n_9439;
assign n_9442 = n_9441 ^ x80;
assign n_9443 = n_9442 ^ x81;
assign n_9444 = n_9315 ^ n_9442;
assign n_9445 = n_9443 & n_9444;
assign n_9446 = n_9445 ^ x81;
assign n_9447 = n_9446 ^ x82;
assign n_9448 = n_9316 ^ n_9446;
assign n_9449 = n_9447 & n_9448;
assign n_9450 = n_9449 ^ x82;
assign n_9451 = n_9450 ^ x83;
assign n_9452 = n_9317 ^ n_9450;
assign n_9453 = n_9451 & n_9452;
assign n_9454 = n_9453 ^ x83;
assign n_9455 = n_9454 ^ x84;
assign n_9456 = n_9318 ^ n_9454;
assign n_9457 = n_9455 & n_9456;
assign n_9458 = n_9457 ^ x84;
assign n_9459 = n_9458 ^ x85;
assign n_9460 = n_9319 ^ n_9458;
assign n_9461 = n_9459 & ~n_9460;
assign n_9462 = n_9461 ^ x85;
assign n_9463 = n_9462 ^ x86;
assign n_9464 = n_9320 ^ n_9462;
assign n_9465 = n_9463 & n_9464;
assign n_9466 = n_9465 ^ x86;
assign n_9467 = n_9466 ^ x87;
assign n_9468 = n_9321 ^ n_9466;
assign n_9469 = n_9467 & n_9468;
assign n_9470 = n_9469 ^ x87;
assign n_9471 = n_9470 ^ x88;
assign n_9472 = n_9322 ^ n_9470;
assign n_9473 = n_9471 & n_9472;
assign n_9474 = n_9473 ^ x88;
assign n_9475 = n_9474 ^ x89;
assign n_9476 = n_9323 ^ n_9474;
assign n_9477 = n_9475 & n_9476;
assign n_9478 = n_9477 ^ x89;
assign n_9479 = n_9478 ^ x90;
assign n_9480 = n_9324 ^ n_9478;
assign n_9481 = n_9479 & n_9480;
assign n_9482 = n_9481 ^ x90;
assign n_9483 = n_9482 ^ x91;
assign n_9484 = n_9325 ^ n_9482;
assign n_9485 = n_9483 & n_9484;
assign n_9486 = n_9485 ^ x91;
assign n_9487 = n_9486 ^ x92;
assign n_9488 = n_9326 ^ n_9486;
assign n_9489 = n_9487 & n_9488;
assign n_9490 = n_9489 ^ x92;
assign n_9491 = n_9490 ^ x93;
assign n_9492 = n_9327 ^ n_9490;
assign n_9493 = n_9491 & n_9492;
assign n_9494 = n_9493 ^ x93;
assign n_9495 = n_9494 ^ x94;
assign n_9496 = n_9328 ^ n_9494;
assign n_9497 = n_9495 & n_9496;
assign n_9498 = n_9497 ^ x94;
assign n_9499 = n_9498 ^ x95;
assign n_9500 = n_9329 ^ n_9498;
assign n_9501 = n_9499 & n_9500;
assign n_9502 = n_9501 ^ x95;
assign n_9503 = n_9502 ^ x96;
assign n_9504 = n_9330 ^ n_9502;
assign n_9505 = n_9503 & n_9504;
assign n_9506 = n_9505 ^ x96;
assign n_9507 = n_9506 ^ x97;
assign n_9508 = n_9331 ^ n_9506;
assign n_9509 = n_9507 & n_9508;
assign n_9510 = n_9509 ^ x97;
assign n_9511 = n_9510 ^ x98;
assign n_9512 = n_9332 ^ n_9510;
assign n_9513 = n_9511 & n_9512;
assign n_9514 = n_9513 ^ x98;
assign n_9515 = n_9514 ^ x99;
assign n_9516 = n_9333 ^ n_9514;
assign n_9517 = n_9515 & n_9516;
assign n_9518 = n_9517 ^ x99;
assign n_9519 = n_9518 ^ x100;
assign n_9520 = n_9518 ^ n_9299;
assign n_9521 = n_9376 & n_9518;
assign n_9522 = n_9519 & n_9520;
assign n_9523 = ~n_9381 & ~n_9521;
assign n_9524 = n_9522 ^ x100;
assign n_9525 = x102 ^ n_9523;
assign n_9526 = n_9349 ^ n_9523;
assign n_9527 = n_9524 ^ x101;
assign n_9528 = ~n_9525 & ~n_9526;
assign n_9529 = n_9528 ^ x102;
assign n_9530 = n_9529 ^ x103;
assign n_9531 = n_9334 ^ n_9529;
assign n_9532 = n_9530 & n_9531;
assign n_9533 = n_9532 ^ x103;
assign n_9534 = n_9533 ^ x104;
assign n_9535 = n_9335 ^ n_9533;
assign n_9536 = n_9534 & n_9535;
assign n_9537 = n_9536 ^ x104;
assign n_9538 = n_9537 ^ x105;
assign n_9539 = n_9336 ^ n_9537;
assign n_9540 = n_9538 & n_9539;
assign n_9541 = n_9540 ^ x105;
assign n_9542 = n_9541 ^ x106;
assign n_9543 = n_9337 ^ n_9541;
assign n_9544 = n_9542 & n_9543;
assign n_9545 = n_9544 ^ x106;
assign n_9546 = n_9545 ^ x107;
assign n_9547 = n_9338 ^ n_9545;
assign n_9548 = n_9546 & n_9547;
assign n_9549 = n_9548 ^ x107;
assign n_9550 = n_9549 ^ x108;
assign n_9551 = n_9339 ^ n_9549;
assign n_9552 = n_9550 & n_9551;
assign n_9553 = n_9552 ^ x108;
assign n_9554 = n_9553 ^ x109;
assign n_9555 = n_9340 ^ n_9553;
assign n_9556 = n_9554 & n_9555;
assign n_9557 = n_9556 ^ x109;
assign n_9558 = n_9557 ^ x110;
assign n_9559 = n_9341 ^ n_9557;
assign n_9560 = n_9558 & n_9559;
assign n_9561 = n_9560 ^ x110;
assign n_9562 = n_9561 ^ x111;
assign n_9563 = n_9342 ^ n_9561;
assign n_9564 = n_9562 & n_9563;
assign n_9565 = n_9564 ^ x111;
assign n_9566 = n_9565 ^ x112;
assign n_9567 = n_9343 ^ n_9565;
assign n_9568 = n_9566 & n_9567;
assign n_9569 = n_9568 ^ x112;
assign n_9570 = n_9569 ^ x113;
assign n_9571 = n_9344 ^ n_9569;
assign n_9572 = n_9570 & n_9571;
assign n_9573 = n_9572 ^ x113;
assign n_9574 = n_9573 ^ x114;
assign n_9575 = n_9345 ^ n_9573;
assign n_9576 = n_9574 & n_9575;
assign n_9577 = n_9576 ^ x114;
assign n_9578 = ~n_9577 & ~n_9373;
assign n_9579 = n_9577 ^ x115;
assign n_9580 = ~n_9365 & ~n_9578;
assign n_9581 = ~n_9578 & ~n_9374;
assign n_9582 = ~n_9580 & n_8910;
assign n_9583 = n_9580 ^ x116;
assign n_9584 = n_9297 & ~n_9580;
assign n_9585 = ~x116 & ~n_9581;
assign n_9586 = ~n_9583 & n_9584;
assign n_9587 = ~n_9582 & ~n_9585;
assign n_9588 = n_9583 ^ n_9586;
assign n_9589 = n_353 & ~n_9587;
assign n_9590 = n_353 & n_9588;
assign n_9591 = x64 & n_9589;
assign n_9592 = n_9566 & n_9589;
assign n_9593 = n_9562 & n_9589;
assign n_9594 = n_9424 & n_9589;
assign n_9595 = n_9420 & n_9589;
assign n_9596 = n_9396 & n_9589;
assign n_9597 = n_9392 & n_9589;
assign n_9598 = n_266 & n_9589;
assign n_9599 = n_9385 & n_9589;
assign n_9600 = n_9388 & n_9589;
assign n_9601 = n_9400 & n_9589;
assign n_9602 = n_9404 & n_9589;
assign n_9603 = n_9409 & n_9589;
assign n_9604 = n_9413 & n_9589;
assign n_9605 = n_9416 & n_9589;
assign n_9606 = n_9429 & n_9589;
assign n_9607 = n_9432 & n_9589;
assign n_9608 = ~n_9438 & n_9589;
assign n_9609 = n_9443 & n_9589;
assign n_9610 = n_9447 & n_9589;
assign n_9611 = n_9451 & n_9589;
assign n_9612 = n_9455 & n_9589;
assign n_9613 = n_9459 & n_9589;
assign n_9614 = n_9463 & n_9589;
assign n_9615 = n_9467 & n_9589;
assign n_9616 = n_9471 & n_9589;
assign n_9617 = n_9475 & n_9589;
assign n_9618 = n_9479 & n_9589;
assign n_9619 = n_9483 & n_9589;
assign n_9620 = n_9487 & n_9589;
assign n_9621 = n_9491 & n_9589;
assign n_9622 = n_9495 & n_9589;
assign n_9623 = n_9499 & n_9589;
assign n_9624 = n_9503 & n_9589;
assign n_9625 = n_9507 & n_9589;
assign n_9626 = n_9511 & n_9589;
assign n_9627 = n_9515 & n_9589;
assign n_9628 = n_9519 & n_9589;
assign n_9629 = ~n_9525 & n_9589;
assign n_9630 = n_9530 & n_9589;
assign n_9631 = n_9534 & n_9589;
assign n_9632 = n_9538 & n_9589;
assign n_9633 = n_9542 & n_9589;
assign n_9634 = n_9546 & n_9589;
assign n_9635 = n_9550 & n_9589;
assign n_9636 = n_9554 & n_9589;
assign n_9637 = n_9558 & n_9589;
assign n_9638 = n_9570 & n_9589;
assign n_9639 = n_9574 & n_9589;
assign n_9640 = n_9579 & n_9589;
assign y11 = n_9589;
assign n_9641 = n_9440 & n_9589;
assign n_9642 = n_9527 & n_9589;
assign n_9643 = n_8910 & ~n_9590;
assign n_9644 = n_9591 ^ x11;
assign n_9645 = n_326 & n_9591;
assign n_9646 = n_9592 ^ n_9343;
assign n_9647 = n_9593 ^ n_9342;
assign n_9648 = n_9594 ^ n_9313;
assign n_9649 = n_9595 ^ n_9312;
assign n_9650 = n_9596 ^ n_9308;
assign n_9651 = n_9597 ^ n_9307;
assign n_9652 = n_9598 ^ n_9362;
assign n_9653 = n_9599 ^ n_9366;
assign n_9654 = n_9600 ^ n_9306;
assign n_9655 = n_9601 ^ n_9309;
assign n_9656 = n_9602 ^ n_9310;
assign n_9657 = n_9603 ^ n_9303;
assign n_9658 = n_9604 ^ n_9302;
assign n_9659 = n_9605 ^ n_9311;
assign n_9660 = n_9606 ^ n_9348;
assign n_9661 = n_9607 ^ n_9301;
assign n_9662 = n_9608 ^ n_9314;
assign n_9663 = n_9609 ^ n_9315;
assign n_9664 = n_9610 ^ n_9316;
assign n_9665 = n_9611 ^ n_9317;
assign n_9666 = n_9612 ^ n_9318;
assign n_9667 = n_9613 ^ n_9319;
assign n_9668 = n_9614 ^ n_9320;
assign n_9669 = n_9615 ^ n_9321;
assign n_9670 = n_9616 ^ n_9322;
assign n_9671 = n_9617 ^ n_9323;
assign n_9672 = n_9618 ^ n_9324;
assign n_9673 = n_9619 ^ n_9325;
assign n_9674 = n_9620 ^ n_9326;
assign n_9675 = n_9621 ^ n_9327;
assign n_9676 = n_9622 ^ n_9328;
assign n_9677 = n_9623 ^ n_9329;
assign n_9678 = n_9624 ^ n_9330;
assign n_9679 = n_9625 ^ n_9331;
assign n_9680 = n_9626 ^ n_9332;
assign n_9681 = n_9627 ^ n_9333;
assign n_9682 = n_9628 ^ n_9299;
assign n_9683 = n_9629 ^ n_9349;
assign n_9684 = n_9630 ^ n_9334;
assign n_9685 = n_9631 ^ n_9335;
assign n_9686 = n_9632 ^ n_9336;
assign n_9687 = n_9633 ^ n_9337;
assign n_9688 = n_9634 ^ n_9338;
assign n_9689 = n_9635 ^ n_9339;
assign n_9690 = n_9636 ^ n_9340;
assign n_9691 = n_9637 ^ n_9341;
assign n_9692 = n_9638 ^ n_9344;
assign n_9693 = n_9639 ^ n_9345;
assign n_9694 = n_9640 ^ n_9346;
assign n_9695 = n_9300 ^ n_9641;
assign n_9696 = n_9298 ^ n_9642;
assign n_9697 = x117 ^ n_9643;
assign n_9698 = x119 & ~n_9643;
assign n_9699 = n_9644 ^ x65;
assign n_9700 = n_9644 & ~n_287;
assign n_9701 = n_9644 & n_345;
assign n_9702 = n_9645 ^ n_101;
assign n_9703 = ~x113 ^ n_9646;
assign n_9704 = n_9646 ^ x113;
assign n_9705 = n_9647 ^ x112;
assign n_9706 = x112 & ~n_9647;
assign n_9707 = ~x77 ^ n_9648;
assign n_9708 = n_9648 ^ x77;
assign n_9709 = n_9649 ^ x76;
assign n_9710 = x76 & ~n_9649;
assign n_9711 = n_9650 ^ x70;
assign n_9712 = n_9651 ^ x69;
assign n_9713 = n_9652 ^ x12;
assign n_9714 = n_348 & ~n_9698;
assign n_9715 = ~n_311 & n_9699;
assign n_9716 = ~n_9699 & n_351;
assign n_9717 = n_9700 ^ x9;
assign n_9718 = n_320 ^ n_9702;
assign n_9719 = n_9705 ^ n_9706;
assign n_9720 = n_9706 ^ n_9646;
assign n_9721 = n_9709 ^ n_9710;
assign n_9722 = n_9710 ^ n_9648;
assign n_9723 = n_9713 ^ x66;
assign n_9724 = n_9716 ^ n_267;
assign n_9725 = n_9718 ^ n_337;
assign n_9726 = n_9703 & ~n_9719;
assign n_9727 = ~n_9704 & n_9720;
assign n_9728 = n_9707 & ~n_9721;
assign n_9729 = ~n_9708 & n_9722;
assign n_9730 = n_9701 ^ n_9724;
assign n_9731 = n_9725 ^ n_9713;
assign n_9732 = n_9725 ^ x66;
assign n_9733 = n_9727 ^ x113;
assign n_9734 = n_9729 ^ x77;
assign n_9735 = ~n_9723 & n_9731;
assign n_9736 = n_9735 ^ x66;
assign n_9737 = n_9736 ^ x67;
assign n_9738 = n_9653 ^ n_9736;
assign n_9739 = n_9737 & n_9738;
assign n_9740 = n_9739 ^ x67;
assign n_9741 = n_9740 ^ x68;
assign n_9742 = n_9654 ^ n_9740;
assign n_9743 = n_9741 & n_9742;
assign n_9744 = n_9743 ^ x68;
assign n_9745 = n_9744 ^ n_9651;
assign n_9746 = n_9744 ^ x69;
assign n_9747 = ~n_9712 & n_9745;
assign n_9748 = n_9747 ^ x69;
assign n_9749 = n_9748 ^ n_9650;
assign n_9750 = n_9748 ^ x70;
assign n_9751 = ~n_9711 & n_9749;
assign n_9752 = n_9751 ^ x70;
assign n_9753 = n_9752 ^ x71;
assign n_9754 = n_9655 ^ n_9752;
assign n_9755 = n_9753 & n_9754;
assign n_9756 = n_9755 ^ x71;
assign n_9757 = n_9756 ^ x72;
assign n_9758 = n_9656 ^ n_9756;
assign n_9759 = n_9757 & n_9758;
assign n_9760 = n_9759 ^ x72;
assign n_9761 = n_9760 ^ x73;
assign n_9762 = n_9657 ^ n_9760;
assign n_9763 = n_9761 & n_9762;
assign n_9764 = n_9763 ^ x73;
assign n_9765 = n_9764 ^ x74;
assign n_9766 = n_9658 ^ n_9764;
assign n_9767 = n_9765 & n_9766;
assign n_9768 = n_9767 ^ x74;
assign n_9769 = n_9768 ^ x75;
assign n_9770 = n_9659 ^ n_9768;
assign n_9771 = n_9769 & n_9770;
assign n_9772 = n_9771 ^ x75;
assign n_9773 = n_9772 ^ x76;
assign n_9774 = n_9772 ^ n_9649;
assign n_9775 = n_9728 & n_9772;
assign n_9776 = n_9773 & n_9774;
assign n_9777 = ~n_9734 & ~n_9775;
assign n_9778 = n_9776 ^ x76;
assign n_9779 = x78 ^ n_9777;
assign n_9780 = n_9660 ^ n_9777;
assign n_9781 = n_9778 ^ x77;
assign n_9782 = ~n_9779 & ~n_9780;
assign n_9783 = n_9782 ^ x78;
assign n_9784 = n_9783 ^ x79;
assign n_9785 = n_9661 ^ n_9783;
assign n_9786 = n_9784 & n_9785;
assign n_9787 = n_9786 ^ x79;
assign n_9788 = n_9787 ^ x80;
assign n_9789 = n_9695 ^ n_9787;
assign n_9790 = n_9788 & n_9789;
assign n_9791 = n_9790 ^ x80;
assign n_9792 = n_9791 ^ x81;
assign n_9793 = n_9662 ^ n_9791;
assign n_9794 = n_9792 & n_9793;
assign n_9795 = n_9794 ^ x81;
assign n_9796 = n_9795 ^ x82;
assign n_9797 = n_9663 ^ n_9795;
assign n_9798 = n_9796 & n_9797;
assign n_9799 = n_9798 ^ x82;
assign n_9800 = n_9799 ^ x83;
assign n_9801 = n_9664 ^ n_9799;
assign n_9802 = n_9800 & n_9801;
assign n_9803 = n_9802 ^ x83;
assign n_9804 = n_9803 ^ x84;
assign n_9805 = n_9665 ^ n_9803;
assign n_9806 = n_9804 & n_9805;
assign n_9807 = n_9806 ^ x84;
assign n_9808 = n_9807 ^ x85;
assign n_9809 = n_9666 ^ n_9807;
assign n_9810 = n_9808 & n_9809;
assign n_9811 = n_9810 ^ x85;
assign n_9812 = n_9811 ^ x86;
assign n_9813 = n_9667 ^ n_9811;
assign n_9814 = n_9812 & ~n_9813;
assign n_9815 = n_9814 ^ x86;
assign n_9816 = n_9815 ^ x87;
assign n_9817 = n_9668 ^ n_9815;
assign n_9818 = n_9816 & n_9817;
assign n_9819 = n_9818 ^ x87;
assign n_9820 = n_9819 ^ x88;
assign n_9821 = n_9669 ^ n_9819;
assign n_9822 = n_9820 & n_9821;
assign n_9823 = n_9822 ^ x88;
assign n_9824 = n_9823 ^ x89;
assign n_9825 = n_9670 ^ n_9823;
assign n_9826 = n_9824 & n_9825;
assign n_9827 = n_9826 ^ x89;
assign n_9828 = n_9827 ^ x90;
assign n_9829 = n_9671 ^ n_9827;
assign n_9830 = n_9828 & n_9829;
assign n_9831 = n_9830 ^ x90;
assign n_9832 = n_9831 ^ x91;
assign n_9833 = n_9672 ^ n_9831;
assign n_9834 = n_9832 & n_9833;
assign n_9835 = n_9834 ^ x91;
assign n_9836 = n_9835 ^ x92;
assign n_9837 = n_9673 ^ n_9835;
assign n_9838 = n_9836 & n_9837;
assign n_9839 = n_9838 ^ x92;
assign n_9840 = n_9839 ^ x93;
assign n_9841 = n_9674 ^ n_9839;
assign n_9842 = n_9840 & n_9841;
assign n_9843 = n_9842 ^ x93;
assign n_9844 = n_9843 ^ x94;
assign n_9845 = n_9675 ^ n_9843;
assign n_9846 = n_9844 & n_9845;
assign n_9847 = n_9846 ^ x94;
assign n_9848 = n_9847 ^ x95;
assign n_9849 = n_9676 ^ n_9847;
assign n_9850 = n_9848 & n_9849;
assign n_9851 = n_9850 ^ x95;
assign n_9852 = n_9851 ^ x96;
assign n_9853 = n_9677 ^ n_9851;
assign n_9854 = n_9852 & n_9853;
assign n_9855 = n_9854 ^ x96;
assign n_9856 = n_9855 ^ x97;
assign n_9857 = n_9678 ^ n_9855;
assign n_9858 = n_9856 & n_9857;
assign n_9859 = n_9858 ^ x97;
assign n_9860 = n_9859 ^ x98;
assign n_9861 = n_9679 ^ n_9859;
assign n_9862 = n_9860 & n_9861;
assign n_9863 = n_9862 ^ x98;
assign n_9864 = n_9863 ^ x99;
assign n_9865 = n_9680 ^ n_9863;
assign n_9866 = n_9864 & n_9865;
assign n_9867 = n_9866 ^ x99;
assign n_9868 = n_9867 ^ x100;
assign n_9869 = n_9681 ^ n_9867;
assign n_9870 = n_9868 & n_9869;
assign n_9871 = n_9870 ^ x100;
assign n_9872 = n_9871 ^ x101;
assign n_9873 = n_9682 ^ n_9871;
assign n_9874 = n_9872 & n_9873;
assign n_9875 = n_9874 ^ x101;
assign n_9876 = n_9875 ^ x102;
assign n_9877 = n_9696 ^ n_9875;
assign n_9878 = n_9876 & n_9877;
assign n_9879 = n_9878 ^ x102;
assign n_9880 = n_9879 ^ x103;
assign n_9881 = n_9683 ^ n_9879;
assign n_9882 = n_9880 & n_9881;
assign n_9883 = n_9882 ^ x103;
assign n_9884 = n_9883 ^ x104;
assign n_9885 = n_9684 ^ n_9883;
assign n_9886 = n_9884 & n_9885;
assign n_9887 = n_9886 ^ x104;
assign n_9888 = n_9887 ^ x105;
assign n_9889 = n_9685 ^ n_9887;
assign n_9890 = n_9888 & n_9889;
assign n_9891 = n_9890 ^ x105;
assign n_9892 = n_9891 ^ x106;
assign n_9893 = n_9686 ^ n_9891;
assign n_9894 = n_9892 & n_9893;
assign n_9895 = n_9894 ^ x106;
assign n_9896 = n_9895 ^ x107;
assign n_9897 = n_9687 ^ n_9895;
assign n_9898 = n_9896 & n_9897;
assign n_9899 = n_9898 ^ x107;
assign n_9900 = n_9899 ^ x108;
assign n_9901 = n_9688 ^ n_9899;
assign n_9902 = n_9900 & n_9901;
assign n_9903 = n_9902 ^ x108;
assign n_9904 = n_9903 ^ x109;
assign n_9905 = n_9689 ^ n_9903;
assign n_9906 = n_9904 & n_9905;
assign n_9907 = n_9906 ^ x109;
assign n_9908 = n_9907 ^ x110;
assign n_9909 = n_9690 ^ n_9907;
assign n_9910 = n_9908 & n_9909;
assign n_9911 = n_9910 ^ x110;
assign n_9912 = n_9911 ^ x111;
assign n_9913 = n_9691 ^ n_9911;
assign n_9914 = n_9912 & n_9913;
assign n_9915 = n_9914 ^ x111;
assign n_9916 = n_9915 ^ x112;
assign n_9917 = n_9915 ^ n_9647;
assign n_9918 = n_9726 & n_9915;
assign n_9919 = n_9916 & n_9917;
assign n_9920 = ~n_9733 & ~n_9918;
assign n_9921 = n_9919 ^ x112;
assign n_9922 = x114 ^ n_9920;
assign n_9923 = n_9692 ^ n_9920;
assign n_9924 = n_9921 ^ x113;
assign n_9925 = ~n_9922 & ~n_9923;
assign n_9926 = n_9925 ^ x114;
assign n_9927 = n_9926 ^ x115;
assign n_9928 = n_9693 ^ n_9926;
assign n_9929 = n_9927 & n_9928;
assign n_9930 = n_9929 ^ x115;
assign n_9931 = n_9930 ^ x116;
assign n_9932 = n_9694 ^ n_9930;
assign n_9933 = n_9931 & n_9932;
assign n_9934 = n_9933 ^ x116;
assign n_9935 = n_9934 ^ x117;
assign n_9936 = n_9935 & ~n_9697;
assign n_9937 = n_9936 ^ x117;
assign n_9938 = n_352 & ~n_9937;
assign n_9939 = n_311 ^ n_9938;
assign n_9940 = x64 & n_9938;
assign n_9941 = n_9644 ^ n_9938;
assign n_9942 = n_328 & n_9938;
assign n_9943 = n_9732 & n_9938;
assign n_9944 = n_9737 & n_9938;
assign n_9945 = n_9741 & n_9938;
assign n_9946 = n_9750 & n_9938;
assign n_9947 = n_9746 & n_9938;
assign n_9948 = n_9753 & n_9938;
assign n_9949 = n_9757 & n_9938;
assign n_9950 = n_9761 & n_9938;
assign n_9951 = n_9765 & n_9938;
assign n_9952 = n_9769 & n_9938;
assign n_9953 = n_9773 & n_9938;
assign n_9954 = ~n_9779 & n_9938;
assign n_9955 = n_9784 & n_9938;
assign n_9956 = n_9788 & n_9938;
assign n_9957 = n_9792 & n_9938;
assign n_9958 = n_9796 & n_9938;
assign n_9959 = n_9800 & n_9938;
assign n_9960 = n_9804 & n_9938;
assign n_9961 = n_9808 & n_9938;
assign n_9962 = n_9812 & n_9938;
assign n_9963 = n_9816 & n_9938;
assign n_9964 = n_9820 & n_9938;
assign n_9965 = n_9824 & n_9938;
assign n_9966 = n_9828 & n_9938;
assign n_9967 = n_9832 & n_9938;
assign n_9968 = n_9916 & n_9938;
assign n_9969 = n_9896 & n_9938;
assign n_9970 = n_9892 & n_9938;
assign n_9971 = n_9836 & n_9938;
assign n_9972 = n_9840 & n_9938;
assign n_9973 = n_9844 & n_9938;
assign n_9974 = n_9848 & n_9938;
assign n_9975 = n_9852 & n_9938;
assign n_9976 = n_9856 & n_9938;
assign n_9977 = n_9860 & n_9938;
assign n_9978 = n_9864 & n_9938;
assign n_9979 = n_9868 & n_9938;
assign n_9980 = n_9872 & n_9938;
assign n_9981 = n_9876 & n_9938;
assign n_9982 = n_9880 & n_9938;
assign n_9983 = n_9884 & n_9938;
assign n_9984 = n_9888 & n_9938;
assign n_9985 = n_9900 & n_9938;
assign n_9986 = n_9904 & n_9938;
assign n_9987 = n_9908 & n_9938;
assign n_9988 = n_9912 & n_9938;
assign n_9989 = n_9927 & n_9938;
assign n_9990 = ~n_9922 & n_9938;
assign n_9991 = n_9935 & n_9938;
assign n_9992 = n_9931 & n_9938;
assign n_9993 = n_169 & n_9938;
assign y10 = n_9938;
assign n_9994 = n_9781 & n_9938;
assign n_9995 = n_9924 & n_9938;
assign n_9996 = n_9699 ^ n_9939;
assign n_9997 = n_101 & ~n_9940;
assign n_9998 = n_338 ^ n_9940;
assign n_9999 = ~n_311 & n_9940;
assign n_10000 = n_9942 ^ n_9724;
assign n_10001 = n_9943 ^ n_9713;
assign n_10002 = n_9944 ^ n_9653;
assign n_10003 = n_9945 ^ n_9654;
assign n_10004 = n_9946 ^ n_9650;
assign n_10005 = n_9947 ^ n_9651;
assign n_10006 = n_9948 ^ n_9655;
assign n_10007 = n_9949 ^ n_9656;
assign n_10008 = n_9950 ^ n_9657;
assign n_10009 = n_9951 ^ n_9658;
assign n_10010 = n_9952 ^ n_9659;
assign n_10011 = n_9953 ^ n_9649;
assign n_10012 = n_9954 ^ n_9660;
assign n_10013 = n_9955 ^ n_9661;
assign n_10014 = n_9956 ^ n_9695;
assign n_10015 = n_9957 ^ n_9662;
assign n_10016 = n_9958 ^ n_9663;
assign n_10017 = n_9959 ^ n_9664;
assign n_10018 = n_9960 ^ n_9665;
assign n_10019 = n_9961 ^ n_9666;
assign n_10020 = n_9962 ^ n_9667;
assign n_10021 = n_9963 ^ n_9668;
assign n_10022 = n_9964 ^ n_9669;
assign n_10023 = n_9965 ^ n_9670;
assign n_10024 = n_9966 ^ n_9671;
assign n_10025 = n_9967 ^ n_9672;
assign n_10026 = n_9968 ^ n_9647;
assign n_10027 = n_9969 ^ n_9687;
assign n_10028 = n_9970 ^ n_9686;
assign n_10029 = n_9971 ^ n_9673;
assign n_10030 = n_9972 ^ n_9674;
assign n_10031 = n_9973 ^ n_9675;
assign n_10032 = n_9974 ^ n_9676;
assign n_10033 = n_9975 ^ n_9677;
assign n_10034 = n_9976 ^ n_9678;
assign n_10035 = n_9977 ^ n_9679;
assign n_10036 = n_9978 ^ n_9680;
assign n_10037 = n_9979 ^ n_9681;
assign n_10038 = n_9980 ^ n_9682;
assign n_10039 = n_9981 ^ n_9696;
assign n_10040 = n_9982 ^ n_9683;
assign n_10041 = n_9983 ^ n_9684;
assign n_10042 = n_9984 ^ n_9685;
assign n_10043 = n_9985 ^ n_9688;
assign n_10044 = n_9986 ^ n_9689;
assign n_10045 = n_9987 ^ n_9690;
assign n_10046 = n_9988 ^ n_9691;
assign n_10047 = n_9989 ^ n_9693;
assign n_10048 = n_9990 ^ n_9692;
assign n_10049 = n_9991 ^ n_9643;
assign n_10050 = n_9992 ^ n_9694;
assign n_10051 = n_9993 ^ n_9644;
assign n_10052 = n_9648 ^ n_9994;
assign n_10053 = n_9646 ^ n_9995;
assign n_10054 = n_9996 & ~n_9715;
assign n_10055 = n_9997 & ~n_9941;
assign n_10056 = n_346 & n_9998;
assign n_10057 = n_9999 ^ x66;
assign n_10058 = n_10000 ^ n_9724;
assign n_10059 = n_10004 ^ x71;
assign n_10060 = n_10004 ^ x70;
assign n_10061 = n_10005 ^ n_10004;
assign n_10062 = n_10026 ^ x113;
assign n_10063 = x113 & ~n_10026;
assign n_10064 = ~x108 ^ n_10027;
assign n_10065 = n_10027 ^ x108;
assign n_10066 = n_10028 ^ x107;
assign n_10067 = x107 & ~n_10028;
assign n_10068 = ~x116 ^ n_10047;
assign n_10069 = n_10047 ^ x116;
assign n_10070 = n_10048 ^ x115;
assign n_10071 = x115 & ~n_10048;
assign n_10072 = n_10049 ^ x118;
assign n_10073 = x118 & ~n_10049;
assign n_10074 = x120 & ~n_10049;
assign n_10075 = ~x114 ^ n_10053;
assign n_10076 = n_10053 ^ x114;
assign n_10077 = ~n_9717 & ~n_10054;
assign n_10078 = ~x66 & ~n_10055;
assign n_10079 = n_10056 ^ n_10057;
assign n_10080 = n_10058 ^ n_9938;
assign n_10081 = n_10004 & n_10061;
assign n_10082 = n_10062 ^ n_10063;
assign n_10083 = n_10063 ^ n_10053;
assign n_10084 = n_10066 ^ n_10067;
assign n_10085 = n_10067 ^ n_10027;
assign n_10086 = n_10070 ^ n_10071;
assign n_10087 = n_10071 ^ n_10047;
assign n_10088 = n_10072 ^ n_10073;
assign n_10089 = n_350 & ~n_10073;
assign n_10090 = n_341 & ~n_10074;
assign n_10091 = x64 & n_10077;
assign n_10092 = n_9730 & n_10080;
assign n_10093 = n_10081 ^ n_10005;
assign n_10094 = n_10060 ^ n_10081;
assign n_10095 = n_10075 & ~n_10082;
assign n_10096 = ~n_10076 & n_10083;
assign n_10097 = n_10064 & ~n_10084;
assign n_10098 = ~n_10065 & n_10085;
assign n_10099 = n_10068 & ~n_10086;
assign n_10100 = ~n_10069 & n_10087;
assign n_10101 = ~n_10050 & ~n_10088;
assign n_10102 = ~n_10091 & n_10078;
assign n_10103 = n_9701 ^ n_10092;
assign n_10104 = n_10094 ^ n_10004;
assign n_10105 = n_10096 ^ x114;
assign n_10106 = n_10098 ^ x108;
assign n_10107 = n_10100 ^ x116;
assign n_10108 = ~n_10101 ^ ~n_130;
assign n_10109 = x117 & n_10101;
assign n_10110 = ~n_10103 & ~n_10102;
assign n_10111 = ~n_10109 & n_10089;
assign n_10112 = x67 ^ n_10110;
assign n_10113 = n_10001 ^ n_10110;
assign n_10114 = n_10112 & n_10113;
assign n_10115 = n_10114 ^ x67;
assign n_10116 = n_10115 ^ x68;
assign n_10117 = n_10002 ^ n_10115;
assign n_10118 = n_10116 & n_10117;
assign n_10119 = n_10118 ^ x68;
assign n_10120 = n_10119 ^ x69;
assign n_10121 = n_10003 ^ n_10119;
assign n_10122 = n_10120 & n_10121;
assign n_10123 = n_10122 ^ x69;
assign n_10124 = ~x70 ^ ~n_10123;
assign n_10125 = n_10123 ^ x70;
assign n_10126 = n_10005 ^ n_10123;
assign n_10127 = n_10124 & ~n_10093;
assign n_10128 = n_10125 ^ n_10059;
assign n_10129 = n_10125 & n_10126;
assign n_10130 = ~n_10128 & n_10104;
assign n_10131 = n_10129 ^ x70;
assign n_10132 = n_10130 ^ n_10081;
assign n_10133 = n_10131 ^ x71;
assign n_10134 = n_10132 ^ n_10004;
assign n_10135 = ~n_10059 & n_10134;
assign n_10136 = x71 ^ n_10135;
assign n_10137 = ~n_10127 & ~n_10136;
assign n_10138 = x72 ^ n_10137;
assign n_10139 = n_10006 ^ n_10137;
assign n_10140 = ~n_10138 & ~n_10139;
assign n_10141 = n_10140 ^ x72;
assign n_10142 = n_10141 ^ x73;
assign n_10143 = n_10007 ^ n_10141;
assign n_10144 = n_10142 & n_10143;
assign n_10145 = n_10144 ^ x73;
assign n_10146 = n_10145 ^ x74;
assign n_10147 = n_10008 ^ n_10145;
assign n_10148 = n_10146 & n_10147;
assign n_10149 = n_10148 ^ x74;
assign n_10150 = n_10149 ^ x75;
assign n_10151 = n_10009 ^ n_10149;
assign n_10152 = n_10150 & n_10151;
assign n_10153 = n_10152 ^ x75;
assign n_10154 = n_10153 ^ x76;
assign n_10155 = n_10010 ^ n_10153;
assign n_10156 = n_10154 & n_10155;
assign n_10157 = n_10156 ^ x76;
assign n_10158 = n_10157 ^ x77;
assign n_10159 = n_10011 ^ n_10157;
assign n_10160 = n_10158 & n_10159;
assign n_10161 = n_10160 ^ x77;
assign n_10162 = n_10161 ^ x78;
assign n_10163 = n_10052 ^ n_10161;
assign n_10164 = n_10162 & n_10163;
assign n_10165 = n_10164 ^ x78;
assign n_10166 = n_10165 ^ x79;
assign n_10167 = n_10012 ^ n_10165;
assign n_10168 = n_10166 & n_10167;
assign n_10169 = n_10168 ^ x79;
assign n_10170 = n_10169 ^ x80;
assign n_10171 = n_10013 ^ n_10169;
assign n_10172 = n_10170 & n_10171;
assign n_10173 = n_10172 ^ x80;
assign n_10174 = n_10173 ^ x81;
assign n_10175 = n_10014 ^ n_10173;
assign n_10176 = n_10174 & n_10175;
assign n_10177 = n_10176 ^ x81;
assign n_10178 = n_10177 ^ x82;
assign n_10179 = n_10015 ^ n_10177;
assign n_10180 = n_10178 & n_10179;
assign n_10181 = n_10180 ^ x82;
assign n_10182 = n_10181 ^ x83;
assign n_10183 = n_10016 ^ n_10181;
assign n_10184 = n_10182 & n_10183;
assign n_10185 = n_10184 ^ x83;
assign n_10186 = n_10185 ^ x84;
assign n_10187 = n_10017 ^ n_10185;
assign n_10188 = n_10186 & n_10187;
assign n_10189 = n_10188 ^ x84;
assign n_10190 = n_10189 ^ x85;
assign n_10191 = n_10018 ^ n_10189;
assign n_10192 = n_10190 & n_10191;
assign n_10193 = n_10192 ^ x85;
assign n_10194 = n_10193 ^ x86;
assign n_10195 = n_10019 ^ n_10193;
assign n_10196 = n_10194 & n_10195;
assign n_10197 = n_10196 ^ x86;
assign n_10198 = n_10197 ^ x87;
assign n_10199 = n_10020 ^ n_10197;
assign n_10200 = n_10198 & ~n_10199;
assign n_10201 = n_10200 ^ x87;
assign n_10202 = n_10201 ^ x88;
assign n_10203 = n_10021 ^ n_10201;
assign n_10204 = n_10202 & n_10203;
assign n_10205 = n_10204 ^ x88;
assign n_10206 = n_10205 ^ x89;
assign n_10207 = n_10022 ^ n_10205;
assign n_10208 = n_10206 & n_10207;
assign n_10209 = n_10208 ^ x89;
assign n_10210 = n_10209 ^ x90;
assign n_10211 = n_10023 ^ n_10209;
assign n_10212 = n_10210 & n_10211;
assign n_10213 = n_10212 ^ x90;
assign n_10214 = n_10213 ^ x91;
assign n_10215 = n_10024 ^ n_10213;
assign n_10216 = n_10214 & n_10215;
assign n_10217 = n_10216 ^ x91;
assign n_10218 = n_10217 ^ x92;
assign n_10219 = n_10025 ^ n_10217;
assign n_10220 = n_10218 & n_10219;
assign n_10221 = n_10220 ^ x92;
assign n_10222 = n_10221 ^ x93;
assign n_10223 = n_10029 ^ n_10221;
assign n_10224 = n_10222 & n_10223;
assign n_10225 = n_10224 ^ x93;
assign n_10226 = n_10225 ^ x94;
assign n_10227 = n_10030 ^ n_10225;
assign n_10228 = n_10226 & n_10227;
assign n_10229 = n_10228 ^ x94;
assign n_10230 = n_10229 ^ x95;
assign n_10231 = n_10031 ^ n_10229;
assign n_10232 = n_10230 & n_10231;
assign n_10233 = n_10232 ^ x95;
assign n_10234 = n_10233 ^ x96;
assign n_10235 = n_10032 ^ n_10233;
assign n_10236 = n_10234 & n_10235;
assign n_10237 = n_10236 ^ x96;
assign n_10238 = n_10237 ^ x97;
assign n_10239 = n_10033 ^ n_10237;
assign n_10240 = n_10238 & n_10239;
assign n_10241 = n_10240 ^ x97;
assign n_10242 = n_10241 ^ x98;
assign n_10243 = n_10034 ^ n_10241;
assign n_10244 = n_10242 & n_10243;
assign n_10245 = n_10244 ^ x98;
assign n_10246 = n_10245 ^ x99;
assign n_10247 = n_10035 ^ n_10245;
assign n_10248 = n_10246 & n_10247;
assign n_10249 = n_10248 ^ x99;
assign n_10250 = n_10249 ^ x100;
assign n_10251 = n_10036 ^ n_10249;
assign n_10252 = n_10250 & n_10251;
assign n_10253 = n_10252 ^ x100;
assign n_10254 = n_10253 ^ x101;
assign n_10255 = n_10037 ^ n_10253;
assign n_10256 = n_10254 & n_10255;
assign n_10257 = n_10256 ^ x101;
assign n_10258 = n_10257 ^ x102;
assign n_10259 = n_10038 ^ n_10257;
assign n_10260 = n_10258 & n_10259;
assign n_10261 = n_10260 ^ x102;
assign n_10262 = n_10261 ^ x103;
assign n_10263 = n_10039 ^ n_10261;
assign n_10264 = n_10262 & n_10263;
assign n_10265 = n_10264 ^ x103;
assign n_10266 = n_10265 ^ x104;
assign n_10267 = n_10040 ^ n_10265;
assign n_10268 = n_10266 & n_10267;
assign n_10269 = n_10268 ^ x104;
assign n_10270 = n_10269 ^ x105;
assign n_10271 = n_10041 ^ n_10269;
assign n_10272 = n_10270 & n_10271;
assign n_10273 = n_10272 ^ x105;
assign n_10274 = n_10273 ^ x106;
assign n_10275 = n_10042 ^ n_10273;
assign n_10276 = n_10274 & n_10275;
assign n_10277 = n_10276 ^ x106;
assign n_10278 = n_10277 ^ x107;
assign n_10279 = n_10277 ^ n_10028;
assign n_10280 = n_10097 & n_10277;
assign n_10281 = n_10278 & n_10279;
assign n_10282 = ~n_10106 & ~n_10280;
assign n_10283 = n_10281 ^ x107;
assign n_10284 = x109 ^ n_10282;
assign n_10285 = n_10043 ^ n_10282;
assign n_10286 = n_10283 ^ x108;
assign n_10287 = ~n_10284 & ~n_10285;
assign n_10288 = n_10287 ^ x109;
assign n_10289 = n_10288 ^ x110;
assign n_10290 = n_10044 ^ n_10288;
assign n_10291 = n_10289 & n_10290;
assign n_10292 = n_10291 ^ x110;
assign n_10293 = n_10292 ^ x111;
assign n_10294 = n_10045 ^ n_10292;
assign n_10295 = n_10293 & n_10294;
assign n_10296 = n_10295 ^ x111;
assign n_10297 = n_10296 ^ x112;
assign n_10298 = n_10046 ^ n_10296;
assign n_10299 = n_10297 & n_10298;
assign n_10300 = n_10299 ^ x112;
assign n_10301 = n_10300 ^ x113;
assign n_10302 = n_10300 ^ n_10026;
assign n_10303 = n_10095 & n_10300;
assign n_10304 = n_10301 & n_10302;
assign n_10305 = ~n_10105 & ~n_10303;
assign n_10306 = n_10304 ^ x113;
assign n_10307 = x115 ^ n_10305;
assign n_10308 = n_10048 ^ n_10305;
assign n_10309 = n_10099 & ~n_10305;
assign n_10310 = n_10306 ^ x114;
assign n_10311 = ~n_10307 & ~n_10308;
assign n_10312 = ~n_10107 & ~n_10309;
assign n_10313 = n_10311 ^ x115;
assign n_10314 = x117 & ~n_10312;
assign n_10315 = x117 ^ n_10312;
assign n_10316 = n_10050 ^ n_10312;
assign n_10317 = n_10108 & ~n_10312;
assign n_10318 = n_10313 ^ x116;
assign n_10319 = n_10314 & ~n_10049;
assign n_10320 = ~n_10315 & ~n_10316;
assign n_10321 = ~n_10317 & n_10111;
assign n_10322 = n_10320 ^ x117;
assign n_10323 = ~n_10315 & n_10321;
assign n_10324 = ~n_10319 & n_10321;
assign n_10325 = n_10322 ^ x118;
assign n_10326 = n_10323 ^ n_10050;
assign n_10327 = n_10222 & n_10324;
assign n_10328 = n_10218 & n_10324;
assign n_10329 = n_170 & n_10324;
assign n_10330 = x64 & n_10324;
assign n_10331 = n_10112 & n_10324;
assign n_10332 = n_10116 & n_10324;
assign n_10333 = n_10120 & n_10324;
assign n_10334 = n_10125 & n_10324;
assign n_10335 = ~n_10138 & n_10324;
assign n_10336 = n_10142 & n_10324;
assign n_10337 = n_10146 & n_10324;
assign n_10338 = n_10150 & n_10324;
assign n_10339 = n_10154 & n_10324;
assign n_10340 = n_10158 & n_10324;
assign n_10341 = n_10162 & n_10324;
assign n_10342 = n_10166 & n_10324;
assign n_10343 = n_10170 & n_10324;
assign n_10344 = n_10174 & n_10324;
assign n_10345 = n_10178 & n_10324;
assign n_10346 = n_10182 & n_10324;
assign n_10347 = n_10186 & n_10324;
assign n_10348 = n_10190 & n_10324;
assign n_10349 = n_10194 & n_10324;
assign n_10350 = n_10198 & n_10324;
assign n_10351 = n_10202 & n_10324;
assign n_10352 = n_10206 & n_10324;
assign n_10353 = n_10210 & n_10324;
assign n_10354 = n_10214 & n_10324;
assign n_10355 = n_10226 & n_10324;
assign n_10356 = n_10230 & n_10324;
assign n_10357 = n_10234 & n_10324;
assign n_10358 = n_10238 & n_10324;
assign n_10359 = n_10242 & n_10324;
assign n_10360 = n_10246 & n_10324;
assign n_10361 = n_10250 & n_10324;
assign n_10362 = n_10254 & n_10324;
assign n_10363 = n_10258 & n_10324;
assign n_10364 = n_10262 & n_10324;
assign n_10365 = n_10266 & n_10324;
assign n_10366 = n_10270 & n_10324;
assign n_10367 = n_10274 & n_10324;
assign n_10368 = n_10278 & n_10324;
assign n_10369 = ~n_10284 & n_10324;
assign n_10370 = n_10289 & n_10324;
assign n_10371 = n_10293 & n_10324;
assign n_10372 = n_10297 & n_10324;
assign n_10373 = n_10301 & n_10324;
assign n_10374 = ~n_10307 & n_10324;
assign y9 = n_10324;
assign n_10375 = ~n_10079 & n_10324;
assign n_10376 = n_10133 & n_10324;
assign n_10377 = n_10318 & n_10324;
assign n_10378 = n_10286 & n_10324;
assign n_10379 = n_10310 & n_10324;
assign n_10380 = n_350 & n_10325;
assign n_10381 = ~x118 ^ n_10326;
assign n_10382 = n_10326 ^ x118;
assign n_10383 = n_10327 ^ n_10029;
assign n_10384 = n_10328 ^ n_10025;
assign n_10385 = n_10329 ^ n_9940;
assign n_10386 = n_10330 & ~n_103;
assign n_10387 = n_10331 ^ n_10001;
assign n_10388 = n_10332 ^ n_10002;
assign n_10389 = n_10333 ^ n_10003;
assign n_10390 = n_10334 ^ n_10005;
assign n_10391 = n_10335 ^ n_10006;
assign n_10392 = n_10336 ^ n_10007;
assign n_10393 = n_10337 ^ n_10008;
assign n_10394 = n_10338 ^ n_10009;
assign n_10395 = n_10339 ^ n_10010;
assign n_10396 = n_10340 ^ n_10011;
assign n_10397 = n_10341 ^ n_10052;
assign n_10398 = n_10342 ^ n_10012;
assign n_10399 = n_10343 ^ n_10013;
assign n_10400 = n_10344 ^ n_10014;
assign n_10401 = n_10345 ^ n_10015;
assign n_10402 = n_10346 ^ n_10016;
assign n_10403 = n_10347 ^ n_10017;
assign n_10404 = n_10348 ^ n_10018;
assign n_10405 = n_10349 ^ n_10019;
assign n_10406 = n_10350 ^ n_10020;
assign n_10407 = n_10351 ^ n_10021;
assign n_10408 = n_10352 ^ n_10022;
assign n_10409 = n_10353 ^ n_10023;
assign n_10410 = n_10354 ^ n_10024;
assign n_10411 = n_10355 ^ n_10030;
assign n_10412 = n_10356 ^ n_10031;
assign n_10413 = n_10357 ^ n_10032;
assign n_10414 = n_10358 ^ n_10033;
assign n_10415 = n_10359 ^ n_10034;
assign n_10416 = n_10360 ^ n_10035;
assign n_10417 = n_10361 ^ n_10036;
assign n_10418 = n_10362 ^ n_10037;
assign n_10419 = n_10363 ^ n_10038;
assign n_10420 = n_10364 ^ n_10039;
assign n_10421 = n_10365 ^ n_10040;
assign n_10422 = n_10366 ^ n_10041;
assign n_10423 = n_10367 ^ n_10042;
assign n_10424 = n_10368 ^ n_10028;
assign n_10425 = n_10369 ^ n_10043;
assign n_10426 = n_10370 ^ n_10044;
assign n_10427 = n_10371 ^ n_10045;
assign n_10428 = n_10372 ^ n_10046;
assign n_10429 = n_10373 ^ n_10026;
assign n_10430 = n_10374 ^ n_10048;
assign n_10431 = n_10051 ^ n_10375;
assign n_10432 = n_10004 ^ n_10376;
assign n_10433 = n_10047 ^ n_10377;
assign n_10434 = n_10027 ^ n_10378;
assign n_10435 = n_10053 ^ n_10379;
assign n_10436 = n_10049 & ~n_10380;
assign n_10437 = ~x94 ^ n_10383;
assign n_10438 = n_10383 ^ x94;
assign n_10439 = n_10384 ^ x93;
assign n_10440 = x93 & ~n_10384;
assign n_10441 = n_10385 ^ x10;
assign n_10442 = n_233 ^ n_10386;
assign n_10443 = n_10433 ^ x117;
assign n_10444 = x117 & ~n_10433;
assign n_10445 = n_350 & n_10436;
assign n_10446 = x121 & ~n_10436;
assign n_10447 = n_10439 ^ n_10440;
assign n_10448 = n_10440 ^ n_10383;
assign n_10449 = n_10441 ^ x66;
assign n_10450 = n_171 ^ n_10442;
assign n_10451 = n_10443 ^ n_10444;
assign n_10452 = n_10444 ^ n_10326;
assign n_10453 = n_331 & ~n_10446;
assign n_10454 = n_10437 & ~n_10447;
assign n_10455 = ~n_10438 & n_10448;
assign n_10456 = n_10450 ^ n_104;
assign n_10457 = n_10381 & ~n_10451;
assign n_10458 = ~n_10382 & n_10452;
assign n_10459 = n_10455 ^ x94;
assign n_10460 = n_10456 ^ n_10441;
assign n_10461 = n_10456 ^ x66;
assign n_10462 = n_10458 ^ x118;
assign n_10463 = ~n_10449 & n_10460;
assign n_10464 = n_10463 ^ x66;
assign n_10465 = n_10464 ^ x67;
assign n_10466 = n_10431 ^ n_10464;
assign n_10467 = n_10465 & n_10466;
assign n_10468 = n_10467 ^ x67;
assign n_10469 = n_10468 ^ x68;
assign n_10470 = n_10387 ^ n_10468;
assign n_10471 = n_10469 & n_10470;
assign n_10472 = n_10471 ^ x68;
assign n_10473 = n_10472 ^ x69;
assign n_10474 = n_10388 ^ n_10472;
assign n_10475 = n_10473 & n_10474;
assign n_10476 = n_10475 ^ x69;
assign n_10477 = n_10476 ^ x70;
assign n_10478 = n_10389 ^ n_10476;
assign n_10479 = n_10477 & n_10478;
assign n_10480 = n_10479 ^ x70;
assign n_10481 = n_10480 ^ x71;
assign n_10482 = n_10390 ^ n_10480;
assign n_10483 = n_10481 & n_10482;
assign n_10484 = n_10483 ^ x71;
assign n_10485 = n_10484 ^ x72;
assign n_10486 = n_10432 ^ n_10484;
assign n_10487 = n_10485 & n_10486;
assign n_10488 = n_10487 ^ x72;
assign n_10489 = n_10488 ^ x73;
assign n_10490 = n_10391 ^ n_10488;
assign n_10491 = n_10489 & n_10490;
assign n_10492 = n_10491 ^ x73;
assign n_10493 = n_10492 ^ x74;
assign n_10494 = n_10392 ^ n_10492;
assign n_10495 = n_10493 & n_10494;
assign n_10496 = n_10495 ^ x74;
assign n_10497 = n_10496 ^ x75;
assign n_10498 = n_10393 ^ n_10496;
assign n_10499 = n_10497 & n_10498;
assign n_10500 = n_10499 ^ x75;
assign n_10501 = n_10500 ^ x76;
assign n_10502 = n_10394 ^ n_10500;
assign n_10503 = n_10501 & n_10502;
assign n_10504 = n_10503 ^ x76;
assign n_10505 = n_10504 ^ x77;
assign n_10506 = n_10395 ^ n_10504;
assign n_10507 = n_10505 & n_10506;
assign n_10508 = n_10507 ^ x77;
assign n_10509 = n_10508 ^ x78;
assign n_10510 = n_10396 ^ n_10508;
assign n_10511 = n_10509 & n_10510;
assign n_10512 = n_10511 ^ x78;
assign n_10513 = n_10512 ^ x79;
assign n_10514 = n_10397 ^ n_10512;
assign n_10515 = n_10513 & n_10514;
assign n_10516 = n_10515 ^ x79;
assign n_10517 = n_10516 ^ x80;
assign n_10518 = n_10398 ^ n_10516;
assign n_10519 = n_10517 & n_10518;
assign n_10520 = n_10519 ^ x80;
assign n_10521 = n_10520 ^ x81;
assign n_10522 = n_10399 ^ n_10520;
assign n_10523 = n_10521 & n_10522;
assign n_10524 = n_10523 ^ x81;
assign n_10525 = n_10524 ^ x82;
assign n_10526 = n_10400 ^ n_10524;
assign n_10527 = n_10525 & n_10526;
assign n_10528 = n_10527 ^ x82;
assign n_10529 = n_10528 ^ x83;
assign n_10530 = n_10401 ^ n_10528;
assign n_10531 = n_10529 & n_10530;
assign n_10532 = n_10531 ^ x83;
assign n_10533 = n_10532 ^ x84;
assign n_10534 = n_10402 ^ n_10532;
assign n_10535 = n_10533 & n_10534;
assign n_10536 = n_10535 ^ x84;
assign n_10537 = n_10536 ^ x85;
assign n_10538 = n_10403 ^ n_10536;
assign n_10539 = n_10537 & n_10538;
assign n_10540 = n_10539 ^ x85;
assign n_10541 = n_10540 ^ x86;
assign n_10542 = n_10404 ^ n_10540;
assign n_10543 = n_10541 & n_10542;
assign n_10544 = n_10543 ^ x86;
assign n_10545 = n_10544 ^ x87;
assign n_10546 = n_10405 ^ n_10544;
assign n_10547 = n_10545 & n_10546;
assign n_10548 = n_10547 ^ x87;
assign n_10549 = n_10548 ^ x88;
assign n_10550 = n_10406 ^ n_10548;
assign n_10551 = n_10549 & ~n_10550;
assign n_10552 = n_10551 ^ x88;
assign n_10553 = n_10552 ^ x89;
assign n_10554 = n_10407 ^ n_10552;
assign n_10555 = n_10553 & n_10554;
assign n_10556 = n_10555 ^ x89;
assign n_10557 = n_10556 ^ x90;
assign n_10558 = n_10408 ^ n_10556;
assign n_10559 = n_10557 & n_10558;
assign n_10560 = n_10559 ^ x90;
assign n_10561 = n_10560 ^ x91;
assign n_10562 = n_10409 ^ n_10560;
assign n_10563 = n_10561 & n_10562;
assign n_10564 = n_10563 ^ x91;
assign n_10565 = n_10564 ^ x92;
assign n_10566 = n_10410 ^ n_10564;
assign n_10567 = n_10565 & n_10566;
assign n_10568 = n_10567 ^ x92;
assign n_10569 = n_10568 ^ x93;
assign n_10570 = n_10568 ^ n_10384;
assign n_10571 = n_10454 & n_10568;
assign n_10572 = n_10569 & n_10570;
assign n_10573 = ~n_10459 & ~n_10571;
assign n_10574 = n_10572 ^ x93;
assign n_10575 = x95 ^ n_10573;
assign n_10576 = n_10411 ^ n_10573;
assign n_10577 = n_10574 ^ x94;
assign n_10578 = ~n_10575 & ~n_10576;
assign n_10579 = n_10578 ^ x95;
assign n_10580 = n_10579 ^ x96;
assign n_10581 = n_10412 ^ n_10579;
assign n_10582 = n_10580 & n_10581;
assign n_10583 = n_10582 ^ x96;
assign n_10584 = n_10583 ^ x97;
assign n_10585 = n_10413 ^ n_10583;
assign n_10586 = n_10584 & n_10585;
assign n_10587 = n_10586 ^ x97;
assign n_10588 = n_10587 ^ x98;
assign n_10589 = n_10414 ^ n_10587;
assign n_10590 = n_10588 & n_10589;
assign n_10591 = n_10590 ^ x98;
assign n_10592 = n_10591 ^ x99;
assign n_10593 = n_10415 ^ n_10591;
assign n_10594 = n_10592 & n_10593;
assign n_10595 = n_10594 ^ x99;
assign n_10596 = n_10595 ^ x100;
assign n_10597 = n_10416 ^ n_10595;
assign n_10598 = n_10596 & n_10597;
assign n_10599 = n_10598 ^ x100;
assign n_10600 = n_10599 ^ x101;
assign n_10601 = n_10417 ^ n_10599;
assign n_10602 = n_10600 & n_10601;
assign n_10603 = n_10602 ^ x101;
assign n_10604 = n_10603 ^ x102;
assign n_10605 = n_10418 ^ n_10603;
assign n_10606 = n_10604 & n_10605;
assign n_10607 = n_10606 ^ x102;
assign n_10608 = n_10607 ^ x103;
assign n_10609 = n_10419 ^ n_10607;
assign n_10610 = n_10608 & n_10609;
assign n_10611 = n_10610 ^ x103;
assign n_10612 = n_10611 ^ x104;
assign n_10613 = n_10420 ^ n_10611;
assign n_10614 = n_10612 & n_10613;
assign n_10615 = n_10614 ^ x104;
assign n_10616 = n_10615 ^ x105;
assign n_10617 = n_10421 ^ n_10615;
assign n_10618 = n_10616 & n_10617;
assign n_10619 = n_10618 ^ x105;
assign n_10620 = n_10619 ^ x106;
assign n_10621 = n_10422 ^ n_10619;
assign n_10622 = n_10620 & n_10621;
assign n_10623 = n_10622 ^ x106;
assign n_10624 = n_10623 ^ x107;
assign n_10625 = n_10423 ^ n_10623;
assign n_10626 = n_10624 & n_10625;
assign n_10627 = n_10626 ^ x107;
assign n_10628 = n_10627 ^ x108;
assign n_10629 = n_10424 ^ n_10627;
assign n_10630 = n_10628 & n_10629;
assign n_10631 = n_10630 ^ x108;
assign n_10632 = n_10631 ^ x109;
assign n_10633 = n_10434 ^ n_10631;
assign n_10634 = n_10632 & n_10633;
assign n_10635 = n_10634 ^ x109;
assign n_10636 = n_10635 ^ x110;
assign n_10637 = n_10425 ^ n_10635;
assign n_10638 = n_10636 & n_10637;
assign n_10639 = n_10638 ^ x110;
assign n_10640 = n_10639 ^ x111;
assign n_10641 = n_10426 ^ n_10639;
assign n_10642 = n_10640 & n_10641;
assign n_10643 = n_10642 ^ x111;
assign n_10644 = n_10643 ^ x112;
assign n_10645 = n_10427 ^ n_10643;
assign n_10646 = n_10644 & n_10645;
assign n_10647 = n_10646 ^ x112;
assign n_10648 = n_10647 ^ x113;
assign n_10649 = n_10428 ^ n_10647;
assign n_10650 = n_10648 & n_10649;
assign n_10651 = n_10650 ^ x113;
assign n_10652 = n_10651 ^ x114;
assign n_10653 = n_10429 ^ n_10651;
assign n_10654 = n_10652 & n_10653;
assign n_10655 = n_10654 ^ x114;
assign n_10656 = n_10655 ^ x115;
assign n_10657 = n_10435 ^ n_10655;
assign n_10658 = n_10656 & n_10657;
assign n_10659 = n_10658 ^ x115;
assign n_10660 = n_10659 ^ x116;
assign n_10661 = n_10430 ^ n_10659;
assign n_10662 = n_10660 & n_10661;
assign n_10663 = n_10662 ^ x116;
assign n_10664 = n_10663 ^ x117;
assign n_10665 = n_10663 ^ n_10433;
assign n_10666 = n_10457 & n_10663;
assign n_10667 = n_10664 & n_10665;
assign n_10668 = ~n_10462 & ~n_10666;
assign n_10669 = n_10667 ^ x117;
assign n_10670 = x119 ^ n_10668;
assign n_10671 = n_10668 & n_9714;
assign n_10672 = n_10669 ^ x118;
assign n_10673 = n_348 & ~n_10670;
assign n_10674 = ~n_10445 & ~n_10671;
assign n_10675 = ~n_10673 & n_10436;
assign n_10676 = n_10624 & ~n_10674;
assign n_10677 = n_10620 & ~n_10674;
assign n_10678 = n_10584 & ~n_10674;
assign n_10679 = n_10580 & ~n_10674;
assign n_10680 = n_10513 & ~n_10674;
assign n_10681 = n_10509 & ~n_10674;
assign n_10682 = n_10485 & ~n_10674;
assign n_10683 = n_10481 & ~n_10674;
assign n_10684 = x64 ^ n_10674;
assign n_10685 = x64 & ~n_10674;
assign n_10686 = x8 ^ n_10674;
assign n_10687 = x65 & ~n_10674;
assign n_10688 = n_10461 & ~n_10674;
assign n_10689 = n_10465 & ~n_10674;
assign n_10690 = n_10469 & ~n_10674;
assign n_10691 = n_10473 & ~n_10674;
assign n_10692 = n_10477 & ~n_10674;
assign n_10693 = n_10489 & ~n_10674;
assign n_10694 = n_10493 & ~n_10674;
assign n_10695 = n_10497 & ~n_10674;
assign n_10696 = n_10501 & ~n_10674;
assign n_10697 = n_10505 & ~n_10674;
assign n_10698 = n_10517 & ~n_10674;
assign n_10699 = n_10521 & ~n_10674;
assign n_10700 = n_10525 & ~n_10674;
assign n_10701 = n_10529 & ~n_10674;
assign n_10702 = n_10533 & ~n_10674;
assign n_10703 = n_10537 & ~n_10674;
assign n_10704 = n_10541 & ~n_10674;
assign n_10705 = n_10545 & ~n_10674;
assign n_10706 = n_10549 & ~n_10674;
assign n_10707 = n_10553 & ~n_10674;
assign n_10708 = n_10557 & ~n_10674;
assign n_10709 = n_10561 & ~n_10674;
assign n_10710 = n_10565 & ~n_10674;
assign n_10711 = n_10569 & ~n_10674;
assign n_10712 = ~n_10575 & ~n_10674;
assign n_10713 = n_10588 & ~n_10674;
assign n_10714 = n_10592 & ~n_10674;
assign n_10715 = n_10596 & ~n_10674;
assign n_10716 = n_10600 & ~n_10674;
assign n_10717 = n_10604 & ~n_10674;
assign n_10718 = n_10608 & ~n_10674;
assign n_10719 = n_10612 & ~n_10674;
assign n_10720 = n_10616 & ~n_10674;
assign n_10721 = n_10628 & ~n_10674;
assign n_10722 = n_10632 & ~n_10674;
assign n_10723 = n_10636 & ~n_10674;
assign n_10724 = n_10664 & ~n_10674;
assign n_10725 = n_10640 & ~n_10674;
assign n_10726 = n_10644 & ~n_10674;
assign n_10727 = n_10648 & ~n_10674;
assign n_10728 = n_10652 & ~n_10674;
assign n_10729 = n_10656 & ~n_10674;
assign n_10730 = n_10660 & ~n_10674;
assign y8 = ~n_10674;
assign n_10731 = n_10577 & ~n_10674;
assign n_10732 = n_10672 & ~n_10674;
assign n_10733 = ~x120 ^ n_10675;
assign n_10734 = x122 & ~n_10675;
assign n_10735 = n_10676 ^ n_10423;
assign n_10736 = n_10677 ^ n_10422;
assign n_10737 = n_10678 ^ n_10413;
assign n_10738 = n_10679 ^ n_10412;
assign n_10739 = n_10680 ^ n_10397;
assign n_10740 = n_10681 ^ n_10396;
assign n_10741 = n_10682 ^ n_10432;
assign n_10742 = n_10683 ^ n_10390;
assign n_10743 = n_10684 ^ n_10685;
assign n_10744 = ~x8 & n_10685;
assign n_10745 = n_234 & n_10686;
assign n_10746 = n_10688 ^ n_10441;
assign n_10747 = n_10689 ^ n_10431;
assign n_10748 = n_10690 ^ n_10387;
assign n_10749 = n_10691 ^ n_10388;
assign n_10750 = n_10692 ^ n_10389;
assign n_10751 = n_10693 ^ n_10391;
assign n_10752 = n_10694 ^ n_10392;
assign n_10753 = n_10695 ^ n_10393;
assign n_10754 = n_10696 ^ n_10394;
assign n_10755 = n_10697 ^ n_10395;
assign n_10756 = n_10698 ^ n_10398;
assign n_10757 = n_10699 ^ n_10399;
assign n_10758 = n_10700 ^ n_10400;
assign n_10759 = n_10701 ^ n_10401;
assign n_10760 = n_10702 ^ n_10402;
assign n_10761 = n_10703 ^ n_10403;
assign n_10762 = n_10704 ^ n_10404;
assign n_10763 = n_10705 ^ n_10405;
assign n_10764 = n_10706 ^ n_10406;
assign n_10765 = n_10707 ^ n_10407;
assign n_10766 = n_10708 ^ n_10408;
assign n_10767 = n_10709 ^ n_10409;
assign n_10768 = n_10710 ^ n_10410;
assign n_10769 = n_10711 ^ n_10384;
assign n_10770 = n_10712 ^ n_10411;
assign n_10771 = n_10713 ^ n_10414;
assign n_10772 = n_10714 ^ n_10415;
assign n_10773 = n_10715 ^ n_10416;
assign n_10774 = n_10716 ^ n_10417;
assign n_10775 = n_10717 ^ n_10418;
assign n_10776 = n_10718 ^ n_10419;
assign n_10777 = n_10719 ^ n_10420;
assign n_10778 = n_10720 ^ n_10421;
assign n_10779 = n_10721 ^ n_10424;
assign n_10780 = n_10722 ^ n_10434;
assign n_10781 = n_10723 ^ n_10425;
assign n_10782 = n_10724 ^ n_10433;
assign n_10783 = n_10725 ^ n_10426;
assign n_10784 = n_10726 ^ n_10427;
assign n_10785 = n_10727 ^ n_10428;
assign n_10786 = n_10728 ^ n_10429;
assign n_10787 = n_10729 ^ n_10435;
assign n_10788 = n_10730 ^ n_10430;
assign n_10789 = n_10383 ^ n_10731;
assign n_10790 = n_10326 ^ n_10732;
assign n_10791 = n_316 & ~n_10734;
assign n_10792 = ~x108 ^ n_10735;
assign n_10793 = n_10735 ^ x108;
assign n_10794 = n_10736 ^ x107;
assign n_10795 = x107 & ~n_10736;
assign n_10796 = n_10737 ^ x98;
assign n_10797 = n_10738 ^ x97;
assign n_10798 = ~x80 ^ n_10739;
assign n_10799 = n_10739 ^ x80;
assign n_10800 = n_10740 ^ x79;
assign n_10801 = x79 & ~n_10740;
assign n_10802 = n_10741 ^ x73;
assign n_10803 = n_10742 ^ x72;
assign n_10804 = n_102 & n_10743;
assign n_10805 = n_10687 ^ n_10744;
assign n_10806 = n_10782 ^ x118;
assign n_10807 = x118 & ~n_10782;
assign n_10808 = ~x119 ^ n_10790;
assign n_10809 = n_10790 ^ x119;
assign n_10810 = n_10794 ^ n_10795;
assign n_10811 = n_10795 ^ n_10735;
assign n_10812 = n_10800 ^ n_10801;
assign n_10813 = n_10801 ^ n_10739;
assign n_10814 = n_10804 ^ n_10745;
assign n_10815 = n_10805 ^ n_10330;
assign n_10816 = n_10806 ^ n_10807;
assign n_10817 = n_10807 ^ n_10790;
assign n_10818 = n_10792 & ~n_10810;
assign n_10819 = ~n_10793 & n_10811;
assign n_10820 = n_10798 & ~n_10812;
assign n_10821 = ~n_10799 & n_10813;
assign n_10822 = ~n_10814 & ~n_296;
assign n_10823 = n_10815 ^ x9;
assign n_10824 = n_10808 & ~n_10816;
assign n_10825 = ~n_10809 & n_10817;
assign n_10826 = n_10819 ^ x108;
assign n_10827 = n_10821 ^ x80;
assign n_10828 = x66 ^ n_10822;
assign n_10829 = n_10823 ^ n_10822;
assign n_10830 = n_10825 ^ x119;
assign n_10831 = ~n_10828 & ~n_10829;
assign n_10832 = n_10831 ^ x66;
assign n_10833 = n_10832 ^ x67;
assign n_10834 = n_10746 ^ n_10832;
assign n_10835 = n_10833 & n_10834;
assign n_10836 = n_10835 ^ x67;
assign n_10837 = n_10836 ^ x68;
assign n_10838 = n_10747 ^ n_10836;
assign n_10839 = n_10837 & n_10838;
assign n_10840 = n_10839 ^ x68;
assign n_10841 = n_10840 ^ x69;
assign n_10842 = n_10748 ^ n_10840;
assign n_10843 = n_10841 & n_10842;
assign n_10844 = n_10843 ^ x69;
assign n_10845 = n_10844 ^ x70;
assign n_10846 = n_10749 ^ n_10844;
assign n_10847 = n_10845 & n_10846;
assign n_10848 = n_10847 ^ x70;
assign n_10849 = n_10848 ^ x71;
assign n_10850 = n_10750 ^ n_10848;
assign n_10851 = n_10849 & n_10850;
assign n_10852 = n_10851 ^ x71;
assign n_10853 = n_10852 ^ n_10742;
assign n_10854 = n_10852 ^ x72;
assign n_10855 = ~n_10803 & n_10853;
assign n_10856 = n_10855 ^ x72;
assign n_10857 = n_10856 ^ n_10741;
assign n_10858 = n_10856 ^ x73;
assign n_10859 = ~n_10802 & n_10857;
assign n_10860 = n_10859 ^ x73;
assign n_10861 = n_10860 ^ x74;
assign n_10862 = n_10751 ^ n_10860;
assign n_10863 = n_10861 & n_10862;
assign n_10864 = n_10863 ^ x74;
assign n_10865 = n_10864 ^ x75;
assign n_10866 = n_10752 ^ n_10864;
assign n_10867 = n_10865 & n_10866;
assign n_10868 = n_10867 ^ x75;
assign n_10869 = n_10868 ^ x76;
assign n_10870 = n_10753 ^ n_10868;
assign n_10871 = n_10869 & n_10870;
assign n_10872 = n_10871 ^ x76;
assign n_10873 = n_10872 ^ x77;
assign n_10874 = n_10754 ^ n_10872;
assign n_10875 = n_10873 & n_10874;
assign n_10876 = n_10875 ^ x77;
assign n_10877 = n_10876 ^ x78;
assign n_10878 = n_10755 ^ n_10876;
assign n_10879 = n_10877 & n_10878;
assign n_10880 = n_10879 ^ x78;
assign n_10881 = n_10880 ^ x79;
assign n_10882 = n_10880 ^ n_10740;
assign n_10883 = n_10820 & n_10880;
assign n_10884 = n_10881 & n_10882;
assign n_10885 = ~n_10827 & ~n_10883;
assign n_10886 = n_10884 ^ x79;
assign n_10887 = x81 ^ n_10885;
assign n_10888 = n_10756 ^ n_10885;
assign n_10889 = n_10886 ^ x80;
assign n_10890 = ~n_10887 & ~n_10888;
assign n_10891 = n_10890 ^ x81;
assign n_10892 = n_10891 ^ x82;
assign n_10893 = n_10757 ^ n_10891;
assign n_10894 = n_10892 & n_10893;
assign n_10895 = n_10894 ^ x82;
assign n_10896 = n_10895 ^ x83;
assign n_10897 = n_10758 ^ n_10895;
assign n_10898 = n_10896 & n_10897;
assign n_10899 = n_10898 ^ x83;
assign n_10900 = n_10899 ^ x84;
assign n_10901 = n_10759 ^ n_10899;
assign n_10902 = n_10900 & n_10901;
assign n_10903 = n_10902 ^ x84;
assign n_10904 = n_10903 ^ x85;
assign n_10905 = n_10760 ^ n_10903;
assign n_10906 = n_10904 & n_10905;
assign n_10907 = n_10906 ^ x85;
assign n_10908 = n_10907 ^ x86;
assign n_10909 = n_10761 ^ n_10907;
assign n_10910 = n_10908 & n_10909;
assign n_10911 = n_10910 ^ x86;
assign n_10912 = n_10911 ^ x87;
assign n_10913 = n_10762 ^ n_10911;
assign n_10914 = n_10912 & n_10913;
assign n_10915 = n_10914 ^ x87;
assign n_10916 = n_10915 ^ x88;
assign n_10917 = n_10763 ^ n_10915;
assign n_10918 = n_10916 & n_10917;
assign n_10919 = n_10918 ^ x88;
assign n_10920 = n_10919 ^ x89;
assign n_10921 = n_10764 ^ n_10919;
assign n_10922 = n_10920 & ~n_10921;
assign n_10923 = n_10922 ^ x89;
assign n_10924 = n_10923 ^ x90;
assign n_10925 = n_10765 ^ n_10923;
assign n_10926 = n_10924 & n_10925;
assign n_10927 = n_10926 ^ x90;
assign n_10928 = n_10927 ^ x91;
assign n_10929 = n_10766 ^ n_10927;
assign n_10930 = n_10928 & n_10929;
assign n_10931 = n_10930 ^ x91;
assign n_10932 = n_10931 ^ x92;
assign n_10933 = n_10767 ^ n_10931;
assign n_10934 = n_10932 & n_10933;
assign n_10935 = n_10934 ^ x92;
assign n_10936 = n_10935 ^ x93;
assign n_10937 = n_10768 ^ n_10935;
assign n_10938 = n_10936 & n_10937;
assign n_10939 = n_10938 ^ x93;
assign n_10940 = n_10939 ^ x94;
assign n_10941 = n_10769 ^ n_10939;
assign n_10942 = n_10940 & n_10941;
assign n_10943 = n_10942 ^ x94;
assign n_10944 = n_10943 ^ x95;
assign n_10945 = n_10789 ^ n_10943;
assign n_10946 = n_10944 & n_10945;
assign n_10947 = n_10946 ^ x95;
assign n_10948 = n_10947 ^ x96;
assign n_10949 = n_10770 ^ n_10947;
assign n_10950 = n_10948 & n_10949;
assign n_10951 = n_10950 ^ x96;
assign n_10952 = n_10951 ^ n_10738;
assign n_10953 = n_10951 ^ x97;
assign n_10954 = ~n_10797 & n_10952;
assign n_10955 = n_10954 ^ x97;
assign n_10956 = n_10955 ^ n_10737;
assign n_10957 = n_10955 ^ x98;
assign n_10958 = ~n_10796 & n_10956;
assign n_10959 = n_10958 ^ x98;
assign n_10960 = n_10959 ^ x99;
assign n_10961 = n_10771 ^ n_10959;
assign n_10962 = n_10960 & n_10961;
assign n_10963 = n_10962 ^ x99;
assign n_10964 = n_10963 ^ x100;
assign n_10965 = n_10772 ^ n_10963;
assign n_10966 = n_10964 & n_10965;
assign n_10967 = n_10966 ^ x100;
assign n_10968 = n_10967 ^ x101;
assign n_10969 = n_10773 ^ n_10967;
assign n_10970 = n_10968 & n_10969;
assign n_10971 = n_10970 ^ x101;
assign n_10972 = n_10971 ^ x102;
assign n_10973 = n_10774 ^ n_10971;
assign n_10974 = n_10972 & n_10973;
assign n_10975 = n_10974 ^ x102;
assign n_10976 = n_10975 ^ x103;
assign n_10977 = n_10775 ^ n_10975;
assign n_10978 = n_10976 & n_10977;
assign n_10979 = n_10978 ^ x103;
assign n_10980 = n_10979 ^ x104;
assign n_10981 = n_10776 ^ n_10979;
assign n_10982 = n_10980 & n_10981;
assign n_10983 = n_10982 ^ x104;
assign n_10984 = n_10983 ^ x105;
assign n_10985 = n_10777 ^ n_10983;
assign n_10986 = n_10984 & n_10985;
assign n_10987 = n_10986 ^ x105;
assign n_10988 = n_10987 ^ x106;
assign n_10989 = n_10778 ^ n_10987;
assign n_10990 = n_10988 & n_10989;
assign n_10991 = n_10990 ^ x106;
assign n_10992 = n_10991 ^ x107;
assign n_10993 = n_10991 ^ n_10736;
assign n_10994 = n_10818 & n_10991;
assign n_10995 = n_10992 & n_10993;
assign n_10996 = ~n_10826 & ~n_10994;
assign n_10997 = n_10995 ^ x107;
assign n_10998 = x109 ^ n_10996;
assign n_10999 = n_10779 ^ n_10996;
assign n_11000 = n_10997 ^ x108;
assign n_11001 = ~n_10998 & ~n_10999;
assign n_11002 = n_11001 ^ x109;
assign n_11003 = n_11002 ^ x110;
assign n_11004 = n_10780 ^ n_11002;
assign n_11005 = n_11003 & n_11004;
assign n_11006 = n_11005 ^ x110;
assign n_11007 = n_11006 ^ x111;
assign n_11008 = n_10781 ^ n_11006;
assign n_11009 = n_11007 & n_11008;
assign n_11010 = n_11009 ^ x111;
assign n_11011 = n_11010 ^ x112;
assign n_11012 = n_10783 ^ n_11010;
assign n_11013 = n_11011 & n_11012;
assign n_11014 = n_11013 ^ x112;
assign n_11015 = n_11014 ^ x113;
assign n_11016 = n_10784 ^ n_11014;
assign n_11017 = n_11015 & n_11016;
assign n_11018 = n_11017 ^ x113;
assign n_11019 = n_11018 ^ x114;
assign n_11020 = n_10785 ^ n_11018;
assign n_11021 = n_11019 & n_11020;
assign n_11022 = n_11021 ^ x114;
assign n_11023 = n_11022 ^ x115;
assign n_11024 = n_10786 ^ n_11022;
assign n_11025 = n_11023 & n_11024;
assign n_11026 = n_11025 ^ x115;
assign n_11027 = n_11026 ^ x116;
assign n_11028 = n_10787 ^ n_11026;
assign n_11029 = n_11027 & n_11028;
assign n_11030 = n_11029 ^ x116;
assign n_11031 = n_11030 ^ x117;
assign n_11032 = n_10788 ^ n_11030;
assign n_11033 = n_11031 & n_11032;
assign n_11034 = n_11033 ^ x117;
assign n_11035 = n_11034 ^ x118;
assign n_11036 = n_11034 ^ n_10782;
assign n_11037 = n_10824 & n_11034;
assign n_11038 = n_11035 & n_11036;
assign n_11039 = ~n_10830 & ~n_11037;
assign n_11040 = n_11038 ^ x118;
assign n_11041 = n_10733 & ~n_11039;
assign n_11042 = x120 ^ n_11039;
assign n_11043 = n_11040 ^ x119;
assign n_11044 = ~n_11041 & n_10090;
assign n_11045 = n_341 & ~n_11042;
assign n_11046 = n_11011 & n_11044;
assign n_11047 = n_11007 & n_11044;
assign n_11048 = n_10992 & n_11044;
assign n_11049 = n_10960 & n_11044;
assign n_11050 = n_10957 & n_11044;
assign n_11051 = n_10944 & n_11044;
assign n_11052 = n_10940 & n_11044;
assign n_11053 = n_10920 & n_11044;
assign n_11054 = n_10916 & n_11044;
assign n_11055 = n_10869 & n_11044;
assign n_11056 = n_10865 & n_11044;
assign n_11057 = x65 & n_11044;
assign n_11058 = x64 & n_11044;
assign n_11059 = ~n_10828 & n_11044;
assign n_11060 = n_10833 & n_11044;
assign n_11061 = n_10837 & n_11044;
assign n_11062 = n_10841 & n_11044;
assign n_11063 = n_10845 & n_11044;
assign n_11064 = n_10849 & n_11044;
assign n_11065 = n_10854 & n_11044;
assign n_11066 = n_10858 & n_11044;
assign n_11067 = n_10861 & n_11044;
assign n_11068 = n_10873 & n_11044;
assign n_11069 = n_10877 & n_11044;
assign n_11070 = n_10881 & n_11044;
assign n_11071 = ~n_10887 & n_11044;
assign n_11072 = n_10892 & n_11044;
assign n_11073 = n_10896 & n_11044;
assign n_11074 = n_10900 & n_11044;
assign n_11075 = n_10904 & n_11044;
assign n_11076 = n_10908 & n_11044;
assign n_11077 = n_10912 & n_11044;
assign n_11078 = n_10924 & n_11044;
assign n_11079 = n_10928 & n_11044;
assign n_11080 = n_10932 & n_11044;
assign n_11081 = n_10936 & n_11044;
assign n_11082 = n_10948 & n_11044;
assign n_11083 = n_10953 & n_11044;
assign n_11084 = n_10964 & n_11044;
assign n_11085 = n_10968 & n_11044;
assign n_11086 = n_10972 & n_11044;
assign n_11087 = n_10976 & n_11044;
assign n_11088 = n_10980 & n_11044;
assign n_11089 = n_10984 & n_11044;
assign n_11090 = n_10988 & n_11044;
assign n_11091 = ~n_10998 & n_11044;
assign n_11092 = n_11003 & n_11044;
assign n_11093 = n_11015 & n_11044;
assign n_11094 = n_11019 & n_11044;
assign n_11095 = n_11023 & n_11044;
assign n_11096 = n_11027 & n_11044;
assign n_11097 = n_11031 & n_11044;
assign n_11098 = n_11035 & n_11044;
assign y7 = n_11044;
assign n_11099 = n_11000 & n_11044;
assign n_11100 = n_10889 & n_11044;
assign n_11101 = n_11043 & n_11044;
assign n_11102 = ~n_11045 & n_10675;
assign n_11103 = n_11046 ^ n_10783;
assign n_11104 = n_11047 ^ n_10781;
assign n_11105 = n_11048 ^ n_10736;
assign n_11106 = n_11049 ^ n_10771;
assign n_11107 = n_11050 ^ n_10737;
assign n_11108 = n_11051 ^ n_10789;
assign n_11109 = n_11052 ^ n_10769;
assign n_11110 = n_11053 ^ n_10764;
assign n_11111 = n_11054 ^ n_10763;
assign n_11112 = n_11055 ^ n_10753;
assign n_11113 = n_11056 ^ n_10752;
assign n_11114 = n_11057 ^ n_10685;
assign n_11115 = n_11058 ^ x7;
assign n_11116 = n_11058 ^ x6;
assign n_11117 = n_11058 ^ n_46;
assign n_11118 = n_11059 ^ n_10823;
assign n_11119 = n_11060 ^ n_10746;
assign n_11120 = n_11061 ^ n_10747;
assign n_11121 = n_11062 ^ n_10748;
assign n_11122 = n_11063 ^ n_10749;
assign n_11123 = n_11064 ^ n_10750;
assign n_11124 = n_11065 ^ n_10742;
assign n_11125 = n_11066 ^ n_10741;
assign n_11126 = n_11067 ^ n_10751;
assign n_11127 = n_11068 ^ n_10754;
assign n_11128 = n_11069 ^ n_10755;
assign n_11129 = n_11070 ^ n_10740;
assign n_11130 = n_11071 ^ n_10756;
assign n_11131 = n_11072 ^ n_10757;
assign n_11132 = n_11073 ^ n_10758;
assign n_11133 = n_11074 ^ n_10759;
assign n_11134 = n_11075 ^ n_10760;
assign n_11135 = n_11076 ^ n_10761;
assign n_11136 = n_11077 ^ n_10762;
assign n_11137 = n_11078 ^ n_10765;
assign n_11138 = n_11079 ^ n_10766;
assign n_11139 = n_11080 ^ n_10767;
assign n_11140 = n_11081 ^ n_10768;
assign n_11141 = n_11082 ^ n_10770;
assign n_11142 = n_11083 ^ n_10738;
assign n_11143 = n_11084 ^ n_10772;
assign n_11144 = n_11085 ^ n_10773;
assign n_11145 = n_11086 ^ n_10774;
assign n_11146 = n_11087 ^ n_10775;
assign n_11147 = n_11088 ^ n_10776;
assign n_11148 = n_11089 ^ n_10777;
assign n_11149 = n_11090 ^ n_10778;
assign n_11150 = n_11091 ^ n_10779;
assign n_11151 = n_11092 ^ n_10780;
assign n_11152 = n_11093 ^ n_10784;
assign n_11153 = n_11094 ^ n_10785;
assign n_11154 = n_11095 ^ n_10786;
assign n_11155 = n_11096 ^ n_10787;
assign n_11156 = n_11097 ^ n_10788;
assign n_11157 = n_11098 ^ n_10782;
assign n_11158 = n_10735 ^ n_11099;
assign n_11159 = n_10739 ^ n_11100;
assign n_11160 = n_10790 ^ n_11101;
assign n_11161 = ~x121 & n_11102;
assign n_11162 = ~n_331 & n_11102;
assign n_11163 = x124 & ~n_11102;
assign n_11164 = ~x113 ^ n_11103;
assign n_11165 = n_11103 ^ x113;
assign n_11166 = n_11104 ^ x112;
assign n_11167 = x112 & ~n_11104;
assign n_11168 = n_11105 ^ x108;
assign n_11169 = x108 & ~n_11105;
assign n_11170 = n_11106 ^ x100;
assign n_11171 = n_11107 ^ x99;
assign n_11172 = n_11108 ^ x96;
assign n_11173 = n_11109 ^ x95;
assign n_11174 = n_11110 ^ x90;
assign n_11175 = n_11111 ^ x89;
assign n_11176 = ~x77 ^ n_11112;
assign n_11177 = n_11112 ^ x77;
assign n_11178 = n_11113 ^ x76;
assign n_11179 = x76 & ~n_11113;
assign n_11180 = n_11058 & n_11115;
assign n_11181 = ~n_11116 & n_11117;
assign n_11182 = ~x109 ^ n_11158;
assign n_11183 = n_11158 ^ x109;
assign n_11184 = n_248 & ~n_11163;
assign n_11185 = n_11166 ^ n_11167;
assign n_11186 = n_11167 ^ n_11103;
assign n_11187 = n_11168 ^ n_11169;
assign n_11188 = n_11169 ^ n_11158;
assign n_11189 = n_11178 ^ n_11179;
assign n_11190 = n_11179 ^ n_11112;
assign n_11191 = n_11114 ^ n_11180;
assign n_11192 = n_11181 ^ n_255;
assign n_11193 = n_11164 & ~n_11185;
assign n_11194 = ~n_11165 & n_11186;
assign n_11195 = n_11182 & ~n_11187;
assign n_11196 = ~n_11183 & n_11188;
assign n_11197 = n_11176 & ~n_11189;
assign n_11198 = ~n_11177 & n_11190;
assign n_11199 = n_11191 ^ x8;
assign n_11200 = n_11192 ^ n_235;
assign n_11201 = n_11194 ^ x113;
assign n_11202 = n_11196 ^ x109;
assign n_11203 = n_11198 ^ x77;
assign n_11204 = n_11199 ^ x66;
assign n_11205 = n_11200 ^ n_11199;
assign n_11206 = n_11200 ^ x66;
assign n_11207 = ~n_11204 & n_11205;
assign n_11208 = n_11207 ^ x66;
assign n_11209 = n_11208 ^ x67;
assign n_11210 = n_11118 ^ n_11208;
assign n_11211 = n_11209 & n_11210;
assign n_11212 = n_11211 ^ x67;
assign n_11213 = n_11212 ^ x68;
assign n_11214 = n_11119 ^ n_11212;
assign n_11215 = n_11213 & n_11214;
assign n_11216 = n_11215 ^ x68;
assign n_11217 = n_11216 ^ x69;
assign n_11218 = n_11120 ^ n_11216;
assign n_11219 = n_11217 & n_11218;
assign n_11220 = n_11219 ^ x69;
assign n_11221 = n_11220 ^ x70;
assign n_11222 = n_11121 ^ n_11220;
assign n_11223 = n_11221 & n_11222;
assign n_11224 = n_11223 ^ x70;
assign n_11225 = n_11224 ^ x71;
assign n_11226 = n_11122 ^ n_11224;
assign n_11227 = n_11225 & n_11226;
assign n_11228 = n_11227 ^ x71;
assign n_11229 = n_11228 ^ x72;
assign n_11230 = n_11123 ^ n_11228;
assign n_11231 = n_11229 & n_11230;
assign n_11232 = n_11231 ^ x72;
assign n_11233 = n_11232 ^ x73;
assign n_11234 = n_11124 ^ n_11232;
assign n_11235 = n_11233 & n_11234;
assign n_11236 = n_11235 ^ x73;
assign n_11237 = n_11236 ^ x74;
assign n_11238 = n_11125 ^ n_11236;
assign n_11239 = n_11237 & n_11238;
assign n_11240 = n_11239 ^ x74;
assign n_11241 = n_11240 ^ x75;
assign n_11242 = n_11126 ^ n_11240;
assign n_11243 = n_11241 & n_11242;
assign n_11244 = n_11243 ^ x75;
assign n_11245 = n_11244 ^ x76;
assign n_11246 = n_11244 ^ n_11113;
assign n_11247 = n_11197 & n_11244;
assign n_11248 = n_11245 & n_11246;
assign n_11249 = ~n_11203 & ~n_11247;
assign n_11250 = n_11248 ^ x76;
assign n_11251 = x78 ^ n_11249;
assign n_11252 = n_11127 ^ n_11249;
assign n_11253 = n_11250 ^ x77;
assign n_11254 = ~n_11251 & ~n_11252;
assign n_11255 = n_11254 ^ x78;
assign n_11256 = n_11255 ^ x79;
assign n_11257 = n_11128 ^ n_11255;
assign n_11258 = n_11256 & n_11257;
assign n_11259 = n_11258 ^ x79;
assign n_11260 = n_11259 ^ x80;
assign n_11261 = n_11129 ^ n_11259;
assign n_11262 = n_11260 & n_11261;
assign n_11263 = n_11262 ^ x80;
assign n_11264 = n_11263 ^ x81;
assign n_11265 = n_11159 ^ n_11263;
assign n_11266 = n_11264 & n_11265;
assign n_11267 = n_11266 ^ x81;
assign n_11268 = n_11267 ^ x82;
assign n_11269 = n_11130 ^ n_11267;
assign n_11270 = n_11268 & n_11269;
assign n_11271 = n_11270 ^ x82;
assign n_11272 = n_11271 ^ x83;
assign n_11273 = n_11131 ^ n_11271;
assign n_11274 = n_11272 & n_11273;
assign n_11275 = n_11274 ^ x83;
assign n_11276 = n_11275 ^ x84;
assign n_11277 = n_11132 ^ n_11275;
assign n_11278 = n_11276 & n_11277;
assign n_11279 = n_11278 ^ x84;
assign n_11280 = n_11279 ^ x85;
assign n_11281 = n_11133 ^ n_11279;
assign n_11282 = n_11280 & n_11281;
assign n_11283 = n_11282 ^ x85;
assign n_11284 = n_11283 ^ x86;
assign n_11285 = n_11134 ^ n_11283;
assign n_11286 = n_11284 & n_11285;
assign n_11287 = n_11286 ^ x86;
assign n_11288 = n_11287 ^ x87;
assign n_11289 = n_11135 ^ n_11287;
assign n_11290 = n_11288 & n_11289;
assign n_11291 = n_11290 ^ x87;
assign n_11292 = n_11291 ^ x88;
assign n_11293 = n_11136 ^ n_11291;
assign n_11294 = n_11292 & n_11293;
assign n_11295 = n_11294 ^ x88;
assign n_11296 = n_11295 ^ n_11111;
assign n_11297 = n_11295 ^ x89;
assign n_11298 = ~n_11175 & n_11296;
assign n_11299 = n_11298 ^ x89;
assign n_11300 = n_11299 ^ n_11110;
assign n_11301 = n_11299 ^ x90;
assign n_11302 = n_11174 & ~n_11300;
assign n_11303 = n_11302 ^ x90;
assign n_11304 = n_11303 ^ x91;
assign n_11305 = n_11137 ^ n_11303;
assign n_11306 = n_11304 & n_11305;
assign n_11307 = n_11306 ^ x91;
assign n_11308 = n_11307 ^ x92;
assign n_11309 = n_11138 ^ n_11307;
assign n_11310 = n_11308 & n_11309;
assign n_11311 = n_11310 ^ x92;
assign n_11312 = n_11311 ^ x93;
assign n_11313 = n_11139 ^ n_11311;
assign n_11314 = n_11312 & n_11313;
assign n_11315 = n_11314 ^ x93;
assign n_11316 = n_11315 ^ x94;
assign n_11317 = n_11140 ^ n_11315;
assign n_11318 = n_11316 & n_11317;
assign n_11319 = n_11318 ^ x94;
assign n_11320 = n_11319 ^ n_11109;
assign n_11321 = n_11319 ^ x95;
assign n_11322 = ~n_11173 & n_11320;
assign n_11323 = n_11322 ^ x95;
assign n_11324 = n_11323 ^ n_11108;
assign n_11325 = n_11323 ^ x96;
assign n_11326 = ~n_11172 & n_11324;
assign n_11327 = n_11326 ^ x96;
assign n_11328 = n_11327 ^ x97;
assign n_11329 = n_11141 ^ n_11327;
assign n_11330 = n_11328 & n_11329;
assign n_11331 = n_11330 ^ x97;
assign n_11332 = n_11331 ^ x98;
assign n_11333 = n_11142 ^ n_11331;
assign n_11334 = n_11332 & n_11333;
assign n_11335 = n_11334 ^ x98;
assign n_11336 = n_11335 ^ n_11107;
assign n_11337 = n_11335 ^ x99;
assign n_11338 = ~n_11171 & n_11336;
assign n_11339 = n_11338 ^ x99;
assign n_11340 = n_11339 ^ n_11106;
assign n_11341 = n_11339 ^ x100;
assign n_11342 = ~n_11170 & n_11340;
assign n_11343 = n_11342 ^ x100;
assign n_11344 = n_11343 ^ x101;
assign n_11345 = n_11143 ^ n_11343;
assign n_11346 = n_11344 & n_11345;
assign n_11347 = n_11346 ^ x101;
assign n_11348 = n_11347 ^ x102;
assign n_11349 = n_11144 ^ n_11347;
assign n_11350 = n_11348 & n_11349;
assign n_11351 = n_11350 ^ x102;
assign n_11352 = n_11351 ^ x103;
assign n_11353 = n_11145 ^ n_11351;
assign n_11354 = n_11352 & n_11353;
assign n_11355 = n_11354 ^ x103;
assign n_11356 = n_11355 ^ x104;
assign n_11357 = n_11146 ^ n_11355;
assign n_11358 = n_11356 & n_11357;
assign n_11359 = n_11358 ^ x104;
assign n_11360 = n_11359 ^ x105;
assign n_11361 = n_11147 ^ n_11359;
assign n_11362 = n_11360 & n_11361;
assign n_11363 = n_11362 ^ x105;
assign n_11364 = n_11363 ^ x106;
assign n_11365 = n_11148 ^ n_11363;
assign n_11366 = n_11364 & n_11365;
assign n_11367 = n_11366 ^ x106;
assign n_11368 = n_11367 ^ x107;
assign n_11369 = n_11149 ^ n_11367;
assign n_11370 = n_11368 & n_11369;
assign n_11371 = n_11370 ^ x107;
assign n_11372 = n_11371 ^ x108;
assign n_11373 = n_11371 ^ n_11105;
assign n_11374 = n_11195 & n_11371;
assign n_11375 = n_11372 & n_11373;
assign n_11376 = ~n_11202 & ~n_11374;
assign n_11377 = n_11375 ^ x108;
assign n_11378 = x110 ^ n_11376;
assign n_11379 = n_11150 ^ n_11376;
assign n_11380 = n_11377 ^ x109;
assign n_11381 = ~n_11378 & ~n_11379;
assign n_11382 = n_11381 ^ x110;
assign n_11383 = n_11382 ^ x111;
assign n_11384 = n_11151 ^ n_11382;
assign n_11385 = n_11383 & n_11384;
assign n_11386 = n_11385 ^ x111;
assign n_11387 = n_11386 ^ x112;
assign n_11388 = n_11386 ^ n_11104;
assign n_11389 = n_11193 & n_11386;
assign n_11390 = n_11387 & n_11388;
assign n_11391 = ~n_11201 & ~n_11389;
assign n_11392 = n_11390 ^ x112;
assign n_11393 = x114 ^ n_11391;
assign n_11394 = n_11152 ^ n_11391;
assign n_11395 = n_11392 ^ x113;
assign n_11396 = ~n_11393 & ~n_11394;
assign n_11397 = n_11396 ^ x114;
assign n_11398 = n_11397 ^ x115;
assign n_11399 = n_11153 ^ n_11397;
assign n_11400 = n_11398 & n_11399;
assign n_11401 = n_11400 ^ x115;
assign n_11402 = n_11401 ^ x116;
assign n_11403 = n_11154 ^ n_11401;
assign n_11404 = n_11402 & n_11403;
assign n_11405 = n_11404 ^ x116;
assign n_11406 = n_11405 ^ x117;
assign n_11407 = n_11155 ^ n_11405;
assign n_11408 = n_11406 & n_11407;
assign n_11409 = n_11408 ^ x117;
assign n_11410 = n_11409 ^ x118;
assign n_11411 = n_11156 ^ n_11409;
assign n_11412 = n_11410 & n_11411;
assign n_11413 = n_11412 ^ x118;
assign n_11414 = n_11413 ^ x119;
assign n_11415 = n_11157 ^ n_11413;
assign n_11416 = n_11414 & n_11415;
assign n_11417 = n_11416 ^ x119;
assign n_11418 = n_11417 ^ x120;
assign n_11419 = n_11160 ^ n_11417;
assign n_11420 = n_11418 & n_11419;
assign n_11421 = n_11420 ^ x120;
assign n_11422 = n_11421 ^ n_11161;
assign n_11423 = n_11161 & ~n_11421;
assign n_11424 = n_11421 ^ x121;
assign n_11425 = n_11422 ^ n_11423;
assign n_11426 = ~n_11423 & ~n_11162;
assign n_11427 = ~n_11424 & n_11102;
assign n_11428 = ~n_11425 & n_10453;
assign n_11429 = n_331 & n_11427;
assign n_11430 = n_11414 & n_11428;
assign n_11431 = n_11410 & n_11428;
assign n_11432 = n_11406 & n_11428;
assign n_11433 = ~n_11393 & n_11428;
assign n_11434 = n_11368 & n_11428;
assign n_11435 = n_11364 & n_11428;
assign n_11436 = n_11312 & n_11428;
assign n_11437 = n_11308 & n_11428;
assign n_11438 = n_11288 & n_11428;
assign n_11439 = n_11284 & n_11428;
assign n_11440 = n_11245 & n_11428;
assign n_11441 = n_11241 & n_11428;
assign n_11442 = x65 & n_11428;
assign n_11443 = x64 & n_11428;
assign n_11444 = n_11206 & n_11428;
assign n_11445 = n_11209 & n_11428;
assign n_11446 = n_11213 & n_11428;
assign n_11447 = n_11217 & n_11428;
assign n_11448 = n_11221 & n_11428;
assign n_11449 = n_11225 & n_11428;
assign n_11450 = n_11229 & n_11428;
assign n_11451 = n_11233 & n_11428;
assign n_11452 = n_11237 & n_11428;
assign n_11453 = ~n_11251 & n_11428;
assign n_11454 = n_11256 & n_11428;
assign n_11455 = n_11260 & n_11428;
assign n_11456 = n_11264 & n_11428;
assign n_11457 = n_11268 & n_11428;
assign n_11458 = n_11272 & n_11428;
assign n_11459 = n_11276 & n_11428;
assign n_11460 = n_11280 & n_11428;
assign n_11461 = n_11292 & n_11428;
assign n_11462 = n_11297 & n_11428;
assign n_11463 = n_11301 & n_11428;
assign n_11464 = n_11304 & n_11428;
assign n_11465 = n_11316 & n_11428;
assign n_11466 = n_11321 & n_11428;
assign n_11467 = n_11325 & n_11428;
assign n_11468 = n_11328 & n_11428;
assign n_11469 = n_11332 & n_11428;
assign n_11470 = n_11337 & n_11428;
assign n_11471 = n_11341 & n_11428;
assign n_11472 = n_11344 & n_11428;
assign n_11473 = n_11348 & n_11428;
assign n_11474 = n_11352 & n_11428;
assign n_11475 = n_11356 & n_11428;
assign n_11476 = n_11360 & n_11428;
assign n_11477 = n_11372 & n_11428;
assign n_11478 = ~n_11378 & n_11428;
assign n_11479 = n_11383 & n_11428;
assign n_11480 = n_11387 & n_11428;
assign n_11481 = n_11398 & n_11428;
assign n_11482 = n_11402 & n_11428;
assign n_11483 = n_11418 & n_11428;
assign n_11484 = x65 ^ n_11428;
assign y6 = n_11428;
assign n_11485 = n_11395 & n_11428;
assign n_11486 = n_11253 & n_11428;
assign n_11487 = n_11380 & n_11428;
assign n_11488 = n_11430 ^ n_11157;
assign n_11489 = n_11431 ^ n_11156;
assign n_11490 = n_11432 ^ n_11155;
assign n_11491 = n_11433 ^ n_11152;
assign n_11492 = n_11434 ^ n_11149;
assign n_11493 = n_11435 ^ n_11148;
assign n_11494 = n_11436 ^ n_11139;
assign n_11495 = n_11437 ^ n_11138;
assign n_11496 = n_11438 ^ n_11135;
assign n_11497 = n_11439 ^ n_11134;
assign n_11498 = n_11440 ^ n_11113;
assign n_11499 = n_11441 ^ n_11126;
assign n_11500 = ~x6 & n_11443;
assign n_11501 = n_11443 ^ x6;
assign n_11502 = x5 & n_11443;
assign n_11503 = n_37 ^ n_11443;
assign n_11504 = n_11444 ^ n_11199;
assign n_11505 = n_11445 ^ n_11118;
assign n_11506 = n_11446 ^ n_11119;
assign n_11507 = n_11447 ^ n_11120;
assign n_11508 = n_11448 ^ n_11121;
assign n_11509 = n_11449 ^ n_11122;
assign n_11510 = n_11450 ^ n_11123;
assign n_11511 = n_11451 ^ n_11124;
assign n_11512 = n_11452 ^ n_11125;
assign n_11513 = n_11453 ^ n_11127;
assign n_11514 = n_11454 ^ n_11128;
assign n_11515 = n_11455 ^ n_11129;
assign n_11516 = n_11456 ^ n_11159;
assign n_11517 = n_11457 ^ n_11130;
assign n_11518 = n_11458 ^ n_11131;
assign n_11519 = n_11459 ^ n_11132;
assign n_11520 = n_11460 ^ n_11133;
assign n_11521 = n_11461 ^ n_11136;
assign n_11522 = n_11462 ^ n_11111;
assign n_11523 = n_11463 ^ n_11110;
assign n_11524 = n_11464 ^ n_11137;
assign n_11525 = n_11465 ^ n_11140;
assign n_11526 = n_11466 ^ n_11109;
assign n_11527 = n_11467 ^ n_11108;
assign n_11528 = n_11468 ^ n_11141;
assign n_11529 = n_11469 ^ n_11142;
assign n_11530 = n_11470 ^ n_11107;
assign n_11531 = n_11471 ^ n_11106;
assign n_11532 = n_11472 ^ n_11143;
assign n_11533 = n_11473 ^ n_11144;
assign n_11534 = n_11474 ^ n_11145;
assign n_11535 = n_11475 ^ n_11146;
assign n_11536 = n_11476 ^ n_11147;
assign n_11537 = n_11477 ^ n_11105;
assign n_11538 = n_11478 ^ n_11150;
assign n_11539 = n_11479 ^ n_11151;
assign n_11540 = n_11480 ^ n_11104;
assign n_11541 = n_11481 ^ n_11153;
assign n_11542 = n_11482 ^ n_11154;
assign n_11543 = n_11483 ^ n_11160;
assign n_11544 = n_11103 ^ n_11485;
assign n_11545 = n_11112 ^ n_11486;
assign n_11546 = n_11158 ^ n_11487;
assign n_11547 = n_11488 ^ x120;
assign n_11548 = n_11489 ^ x119;
assign n_11549 = n_11490 ^ x118;
assign n_11550 = n_11491 ^ x115;
assign n_11551 = ~x108 ^ n_11492;
assign n_11552 = n_11492 ^ x108;
assign n_11553 = n_11493 ^ x107;
assign n_11554 = x107 & ~n_11493;
assign n_11555 = n_11494 ^ x94;
assign n_11556 = n_11495 ^ x93;
assign n_11557 = n_11496 ^ x88;
assign n_11558 = n_11497 ^ x87;
assign n_11559 = n_11498 ^ x77;
assign n_11560 = n_11499 ^ x76;
assign n_11561 = n_11442 ^ n_11500;
assign n_11562 = x65 & ~n_11501;
assign n_11563 = n_106 ^ n_11502;
assign n_11564 = n_11502 ^ n_11503;
assign n_11565 = n_11544 ^ x114;
assign n_11566 = n_11553 ^ n_11554;
assign n_11567 = n_11554 ^ n_11492;
assign n_11568 = n_11561 ^ n_11115;
assign n_11569 = n_236 ^ n_11564;
assign n_11570 = n_11551 & ~n_11566;
assign n_11571 = ~n_11552 & n_11567;
assign n_11572 = n_11568 ^ x66;
assign n_11573 = n_11562 ^ n_11569;
assign n_11574 = n_11571 ^ x108;
assign n_11575 = n_11573 ^ n_11568;
assign n_11576 = n_11573 ^ x66;
assign n_11577 = ~n_11572 & n_11575;
assign n_11578 = n_11577 ^ x66;
assign n_11579 = n_11578 ^ x67;
assign n_11580 = n_11504 ^ n_11578;
assign n_11581 = n_11579 & n_11580;
assign n_11582 = n_11581 ^ x67;
assign n_11583 = n_11582 ^ x68;
assign n_11584 = n_11505 ^ n_11582;
assign n_11585 = n_11583 & n_11584;
assign n_11586 = n_11585 ^ x68;
assign n_11587 = n_11586 ^ x69;
assign n_11588 = n_11506 ^ n_11586;
assign n_11589 = n_11587 & n_11588;
assign n_11590 = n_11589 ^ x69;
assign n_11591 = n_11590 ^ x70;
assign n_11592 = n_11507 ^ n_11590;
assign n_11593 = n_11591 & n_11592;
assign n_11594 = n_11593 ^ x70;
assign n_11595 = n_11594 ^ x71;
assign n_11596 = n_11508 ^ n_11594;
assign n_11597 = n_11595 & n_11596;
assign n_11598 = n_11597 ^ x71;
assign n_11599 = n_11598 ^ x72;
assign n_11600 = n_11509 ^ n_11598;
assign n_11601 = n_11599 & n_11600;
assign n_11602 = n_11601 ^ x72;
assign n_11603 = n_11602 ^ x73;
assign n_11604 = n_11510 ^ n_11602;
assign n_11605 = n_11603 & n_11604;
assign n_11606 = n_11605 ^ x73;
assign n_11607 = n_11606 ^ x74;
assign n_11608 = n_11511 ^ n_11606;
assign n_11609 = n_11607 & n_11608;
assign n_11610 = n_11609 ^ x74;
assign n_11611 = n_11610 ^ x75;
assign n_11612 = n_11512 ^ n_11610;
assign n_11613 = n_11611 & n_11612;
assign n_11614 = n_11613 ^ x75;
assign n_11615 = n_11614 ^ n_11499;
assign n_11616 = n_11614 ^ x76;
assign n_11617 = ~n_11560 & n_11615;
assign n_11618 = n_11617 ^ x76;
assign n_11619 = n_11618 ^ n_11498;
assign n_11620 = n_11618 ^ x77;
assign n_11621 = ~n_11559 & n_11619;
assign n_11622 = n_11621 ^ x77;
assign n_11623 = n_11622 ^ x78;
assign n_11624 = n_11545 ^ n_11622;
assign n_11625 = n_11623 & n_11624;
assign n_11626 = n_11625 ^ x78;
assign n_11627 = n_11626 ^ x79;
assign n_11628 = n_11513 ^ n_11626;
assign n_11629 = n_11627 & n_11628;
assign n_11630 = n_11629 ^ x79;
assign n_11631 = n_11630 ^ x80;
assign n_11632 = n_11514 ^ n_11630;
assign n_11633 = n_11631 & n_11632;
assign n_11634 = n_11633 ^ x80;
assign n_11635 = n_11634 ^ x81;
assign n_11636 = n_11515 ^ n_11634;
assign n_11637 = n_11635 & n_11636;
assign n_11638 = n_11637 ^ x81;
assign n_11639 = n_11638 ^ x82;
assign n_11640 = n_11516 ^ n_11638;
assign n_11641 = n_11639 & n_11640;
assign n_11642 = n_11641 ^ x82;
assign n_11643 = n_11642 ^ x83;
assign n_11644 = n_11517 ^ n_11642;
assign n_11645 = n_11643 & n_11644;
assign n_11646 = n_11645 ^ x83;
assign n_11647 = n_11646 ^ x84;
assign n_11648 = n_11518 ^ n_11646;
assign n_11649 = n_11647 & n_11648;
assign n_11650 = n_11649 ^ x84;
assign n_11651 = n_11650 ^ x85;
assign n_11652 = n_11519 ^ n_11650;
assign n_11653 = n_11651 & n_11652;
assign n_11654 = n_11653 ^ x85;
assign n_11655 = n_11654 ^ x86;
assign n_11656 = n_11520 ^ n_11654;
assign n_11657 = n_11655 & n_11656;
assign n_11658 = n_11657 ^ x86;
assign n_11659 = n_11658 ^ n_11497;
assign n_11660 = n_11658 ^ x87;
assign n_11661 = ~n_11558 & n_11659;
assign n_11662 = n_11661 ^ x87;
assign n_11663 = n_11662 ^ n_11496;
assign n_11664 = n_11662 ^ x88;
assign n_11665 = ~n_11557 & n_11663;
assign n_11666 = n_11665 ^ x88;
assign n_11667 = n_11666 ^ x89;
assign n_11668 = n_11521 ^ n_11666;
assign n_11669 = n_11667 & n_11668;
assign n_11670 = n_11669 ^ x89;
assign n_11671 = n_11670 ^ x90;
assign n_11672 = n_11522 ^ n_11670;
assign n_11673 = n_11671 & n_11672;
assign n_11674 = n_11673 ^ x90;
assign n_11675 = n_11674 ^ x91;
assign n_11676 = n_11523 ^ n_11674;
assign n_11677 = n_11675 & ~n_11676;
assign n_11678 = n_11677 ^ x91;
assign n_11679 = n_11678 ^ x92;
assign n_11680 = n_11524 ^ n_11678;
assign n_11681 = n_11679 & n_11680;
assign n_11682 = n_11681 ^ x92;
assign n_11683 = n_11682 ^ n_11495;
assign n_11684 = n_11682 ^ x93;
assign n_11685 = ~n_11556 & n_11683;
assign n_11686 = n_11685 ^ x93;
assign n_11687 = n_11686 ^ n_11494;
assign n_11688 = n_11686 ^ x94;
assign n_11689 = ~n_11555 & n_11687;
assign n_11690 = n_11689 ^ x94;
assign n_11691 = n_11690 ^ x95;
assign n_11692 = n_11525 ^ n_11690;
assign n_11693 = n_11691 & n_11692;
assign n_11694 = n_11693 ^ x95;
assign n_11695 = n_11694 ^ x96;
assign n_11696 = n_11526 ^ n_11694;
assign n_11697 = n_11695 & n_11696;
assign n_11698 = n_11697 ^ x96;
assign n_11699 = n_11698 ^ x97;
assign n_11700 = n_11527 ^ n_11698;
assign n_11701 = n_11699 & n_11700;
assign n_11702 = n_11701 ^ x97;
assign n_11703 = n_11702 ^ x98;
assign n_11704 = n_11528 ^ n_11702;
assign n_11705 = n_11703 & n_11704;
assign n_11706 = n_11705 ^ x98;
assign n_11707 = n_11706 ^ x99;
assign n_11708 = n_11529 ^ n_11706;
assign n_11709 = n_11707 & n_11708;
assign n_11710 = n_11709 ^ x99;
assign n_11711 = n_11710 ^ x100;
assign n_11712 = n_11530 ^ n_11710;
assign n_11713 = n_11711 & n_11712;
assign n_11714 = n_11713 ^ x100;
assign n_11715 = n_11714 ^ x101;
assign n_11716 = n_11531 ^ n_11714;
assign n_11717 = n_11715 & n_11716;
assign n_11718 = n_11717 ^ x101;
assign n_11719 = n_11718 ^ x102;
assign n_11720 = n_11532 ^ n_11718;
assign n_11721 = n_11719 & n_11720;
assign n_11722 = n_11721 ^ x102;
assign n_11723 = n_11722 ^ x103;
assign n_11724 = n_11533 ^ n_11722;
assign n_11725 = n_11723 & n_11724;
assign n_11726 = n_11725 ^ x103;
assign n_11727 = n_11726 ^ x104;
assign n_11728 = n_11534 ^ n_11726;
assign n_11729 = n_11727 & n_11728;
assign n_11730 = n_11729 ^ x104;
assign n_11731 = n_11730 ^ x105;
assign n_11732 = n_11535 ^ n_11730;
assign n_11733 = n_11731 & n_11732;
assign n_11734 = n_11733 ^ x105;
assign n_11735 = n_11734 ^ x106;
assign n_11736 = n_11536 ^ n_11734;
assign n_11737 = n_11735 & n_11736;
assign n_11738 = n_11737 ^ x106;
assign n_11739 = n_11738 ^ x107;
assign n_11740 = n_11738 ^ n_11493;
assign n_11741 = n_11570 & n_11738;
assign n_11742 = n_11739 & n_11740;
assign n_11743 = ~n_11574 & ~n_11741;
assign n_11744 = n_11742 ^ x107;
assign n_11745 = x109 ^ n_11743;
assign n_11746 = n_11537 ^ n_11743;
assign n_11747 = n_11744 ^ x108;
assign n_11748 = ~n_11745 & ~n_11746;
assign n_11749 = n_11748 ^ x109;
assign n_11750 = n_11749 ^ x110;
assign n_11751 = n_11546 ^ n_11749;
assign n_11752 = n_11750 & n_11751;
assign n_11753 = n_11752 ^ x110;
assign n_11754 = n_11753 ^ x111;
assign n_11755 = n_11538 ^ n_11753;
assign n_11756 = n_11754 & n_11755;
assign n_11757 = n_11756 ^ x111;
assign n_11758 = n_11757 ^ x112;
assign n_11759 = n_11539 ^ n_11757;
assign n_11760 = n_11758 & n_11759;
assign n_11761 = n_11760 ^ x112;
assign n_11762 = n_11761 ^ x113;
assign n_11763 = n_11540 ^ n_11761;
assign n_11764 = n_11762 & n_11763;
assign n_11765 = n_11764 ^ x113;
assign n_11766 = n_11765 ^ n_11544;
assign n_11767 = n_11765 ^ x114;
assign n_11768 = ~n_11565 & n_11766;
assign n_11769 = n_11768 ^ x114;
assign n_11770 = n_11769 ^ n_11491;
assign n_11771 = n_11769 ^ x115;
assign n_11772 = ~n_11550 & n_11770;
assign n_11773 = n_11772 ^ x115;
assign n_11774 = n_11773 ^ x116;
assign n_11775 = n_11541 ^ n_11773;
assign n_11776 = n_11774 & n_11775;
assign n_11777 = n_11776 ^ x116;
assign n_11778 = n_11777 ^ x117;
assign n_11779 = n_11542 ^ n_11777;
assign n_11780 = n_11778 & n_11779;
assign n_11781 = n_11780 ^ x117;
assign n_11782 = n_11781 ^ n_11490;
assign n_11783 = n_11781 ^ x118;
assign n_11784 = ~n_11549 & n_11782;
assign n_11785 = n_11784 ^ x118;
assign n_11786 = n_11785 ^ n_11489;
assign n_11787 = n_11785 ^ x119;
assign n_11788 = ~n_11548 & n_11786;
assign n_11789 = n_11788 ^ x119;
assign n_11790 = n_11789 ^ n_11488;
assign n_11791 = n_11789 ^ x120;
assign n_11792 = ~n_11547 & n_11790;
assign n_11793 = n_11792 ^ x120;
assign n_11794 = n_11793 ^ x121;
assign n_11795 = n_11543 ^ n_11793;
assign n_11796 = n_11794 & n_11795;
assign n_11797 = n_11796 ^ x121;
assign n_11798 = ~n_11797 & n_342;
assign n_11799 = ~n_11797 & n_10791;
assign n_11800 = ~n_11798 & ~n_11426;
assign n_11801 = ~n_11799 & ~n_11429;
assign n_11802 = x127 & ~n_11800;
assign n_11803 = n_11794 & ~n_11801;
assign n_11804 = n_11767 & ~n_11801;
assign n_11805 = n_11762 & ~n_11801;
assign n_11806 = n_11739 & ~n_11801;
assign n_11807 = n_11711 & ~n_11801;
assign n_11808 = n_11707 & ~n_11801;
assign n_11809 = n_11675 & ~n_11801;
assign n_11810 = n_11671 & ~n_11801;
assign n_11811 = n_11639 & ~n_11801;
assign n_11812 = n_11635 & ~n_11801;
assign n_11813 = n_11631 & ~n_11801;
assign n_11814 = n_11627 & ~n_11801;
assign n_11815 = n_11603 & ~n_11801;
assign n_11816 = n_11599 & ~n_11801;
assign n_11817 = n_37 ^ n_11801;
assign n_11818 = n_11428 ^ n_11801;
assign n_11819 = n_11484 & n_11801;
assign n_11820 = x5 ^ n_11801;
assign n_11821 = x4 ^ n_11801;
assign n_11822 = n_11576 & ~n_11801;
assign n_11823 = n_11579 & ~n_11801;
assign n_11824 = n_11583 & ~n_11801;
assign n_11825 = n_11587 & ~n_11801;
assign n_11826 = n_11591 & ~n_11801;
assign n_11827 = n_11595 & ~n_11801;
assign n_11828 = n_11607 & ~n_11801;
assign n_11829 = n_11611 & ~n_11801;
assign n_11830 = n_11616 & ~n_11801;
assign n_11831 = n_11620 & ~n_11801;
assign n_11832 = n_11623 & ~n_11801;
assign n_11833 = n_11647 & ~n_11801;
assign n_11834 = n_11643 & ~n_11801;
assign n_11835 = n_11651 & ~n_11801;
assign n_11836 = n_11655 & ~n_11801;
assign n_11837 = n_11660 & ~n_11801;
assign n_11838 = n_11664 & ~n_11801;
assign n_11839 = n_11667 & ~n_11801;
assign n_11840 = n_11679 & ~n_11801;
assign n_11841 = n_11684 & ~n_11801;
assign n_11842 = n_11688 & ~n_11801;
assign n_11843 = n_11691 & ~n_11801;
assign n_11844 = n_11695 & ~n_11801;
assign n_11845 = n_11699 & ~n_11801;
assign n_11846 = n_11703 & ~n_11801;
assign n_11847 = n_11715 & ~n_11801;
assign n_11848 = n_11719 & ~n_11801;
assign n_11849 = n_11723 & ~n_11801;
assign n_11850 = n_11727 & ~n_11801;
assign n_11851 = n_11731 & ~n_11801;
assign n_11852 = n_11735 & ~n_11801;
assign n_11853 = ~n_11745 & ~n_11801;
assign n_11854 = n_11750 & ~n_11801;
assign n_11855 = n_11754 & ~n_11801;
assign n_11856 = n_11758 & ~n_11801;
assign n_11857 = n_11771 & ~n_11801;
assign n_11858 = n_11774 & ~n_11801;
assign n_11859 = n_11778 & ~n_11801;
assign n_11860 = n_11783 & ~n_11801;
assign n_11861 = n_11787 & ~n_11801;
assign n_11862 = n_11791 & ~n_11801;
assign n_11863 = x64 & n_11801;
assign y5 = ~n_11801;
assign n_11864 = n_11747 & ~n_11801;
assign n_11865 = n_11803 ^ n_11543;
assign n_11866 = n_11804 ^ n_11544;
assign n_11867 = n_11805 ^ n_11540;
assign n_11868 = n_11806 ^ n_11493;
assign n_11869 = n_11807 ^ n_11530;
assign n_11870 = n_11808 ^ n_11529;
assign n_11871 = n_11809 ^ n_11523;
assign n_11872 = n_11810 ^ n_11522;
assign n_11873 = n_11811 ^ n_11516;
assign n_11874 = n_11812 ^ n_11515;
assign n_11875 = n_11813 ^ n_11514;
assign n_11876 = n_11814 ^ n_11513;
assign n_11877 = n_11815 ^ n_11510;
assign n_11878 = n_11816 ^ n_11509;
assign n_11879 = n_11817 & ~n_11818;
assign n_11880 = n_11820 ^ n_95;
assign n_11881 = x64 & n_11821;
assign n_11882 = n_11822 ^ n_11568;
assign n_11883 = n_11823 ^ n_11504;
assign n_11884 = n_11824 ^ n_11505;
assign n_11885 = n_11825 ^ n_11506;
assign n_11886 = n_11826 ^ n_11507;
assign n_11887 = n_11827 ^ n_11508;
assign n_11888 = n_11828 ^ n_11511;
assign n_11889 = n_11829 ^ n_11512;
assign n_11890 = n_11830 ^ n_11499;
assign n_11891 = n_11831 ^ n_11498;
assign n_11892 = n_11832 ^ n_11545;
assign n_11893 = n_11833 ^ n_11518;
assign n_11894 = n_11834 ^ n_11517;
assign n_11895 = n_11835 ^ n_11519;
assign n_11896 = n_11836 ^ n_11520;
assign n_11897 = n_11837 ^ n_11497;
assign n_11898 = n_11838 ^ n_11496;
assign n_11899 = n_11839 ^ n_11521;
assign n_11900 = n_11840 ^ n_11524;
assign n_11901 = n_11841 ^ n_11495;
assign n_11902 = n_11842 ^ n_11494;
assign n_11903 = n_11843 ^ n_11525;
assign n_11904 = n_11844 ^ n_11526;
assign n_11905 = n_11845 ^ n_11527;
assign n_11906 = n_11846 ^ n_11528;
assign n_11907 = n_11847 ^ n_11531;
assign n_11908 = n_11848 ^ n_11532;
assign n_11909 = n_11849 ^ n_11533;
assign n_11910 = n_11850 ^ n_11534;
assign n_11911 = n_11851 ^ n_11535;
assign n_11912 = n_11852 ^ n_11536;
assign n_11913 = n_11853 ^ n_11537;
assign n_11914 = n_11854 ^ n_11546;
assign n_11915 = n_11855 ^ n_11538;
assign n_11916 = n_11856 ^ n_11539;
assign n_11917 = n_11857 ^ n_11491;
assign n_11918 = n_11858 ^ n_11541;
assign n_11919 = n_11859 ^ n_11542;
assign n_11920 = n_11860 ^ n_11490;
assign n_11921 = n_11861 ^ n_11489;
assign n_11922 = n_11862 ^ n_11488;
assign n_11923 = n_11492 ^ n_11864;
assign n_11924 = n_11865 ^ x122;
assign n_11925 = n_11866 ^ x115;
assign n_11926 = n_11867 ^ x114;
assign n_11927 = n_11868 ^ x108;
assign n_11928 = x108 & ~n_11868;
assign n_11929 = n_11869 ^ x101;
assign n_11930 = n_11870 ^ x100;
assign n_11931 = ~x92 ^ ~n_11871;
assign n_11932 = n_11871 ^ x92;
assign n_11933 = n_11872 ^ x91;
assign n_11934 = x91 & ~n_11872;
assign n_11935 = ~x83 ^ n_11873;
assign n_11936 = n_11873 ^ x83;
assign n_11937 = n_11874 ^ x82;
assign n_11938 = x82 & ~n_11874;
assign n_11939 = n_11875 ^ x81;
assign n_11940 = n_11876 ^ x80;
assign n_11941 = n_11877 ^ x74;
assign n_11942 = n_11878 ^ x73;
assign n_11943 = n_11879 ^ n_11819;
assign n_11944 = n_11881 ^ n_11801;
assign n_11945 = ~x85 ^ n_11893;
assign n_11946 = n_11893 ^ x85;
assign n_11947 = n_11894 ^ x84;
assign n_11948 = x84 & ~n_11894;
assign n_11949 = ~x109 ^ n_11923;
assign n_11950 = n_11923 ^ x109;
assign n_11951 = n_11927 ^ n_11928;
assign n_11952 = n_11928 ^ n_11923;
assign n_11953 = n_11933 ^ n_11934;
assign n_11954 = n_11934 ^ n_11871;
assign n_11955 = n_11937 ^ n_11938;
assign n_11956 = n_11938 ^ n_11873;
assign n_11957 = n_11943 ^ n_11563;
assign n_11958 = n_11880 & n_11944;
assign n_11959 = n_11947 ^ n_11948;
assign n_11960 = n_11948 ^ n_11893;
assign n_11961 = n_11949 & ~n_11951;
assign n_11962 = ~n_11950 & n_11952;
assign n_11963 = n_11931 & ~n_11953;
assign n_11964 = n_11932 & ~n_11954;
assign n_11965 = n_11935 & ~n_11955;
assign n_11966 = ~n_11936 & n_11956;
assign n_11967 = n_11957 ^ x66;
assign n_11968 = n_11958 ^ n_11881;
assign n_11969 = n_11945 & ~n_11959;
assign n_11970 = ~n_11946 & n_11960;
assign n_11971 = n_11962 ^ x109;
assign n_11972 = n_11964 ^ x92;
assign n_11973 = n_11966 ^ x83;
assign n_11974 = n_11968 ^ n_11801;
assign n_11975 = n_11970 ^ x85;
assign n_11976 = n_11974 ^ x64;
assign n_11977 = n_11820 & n_11976;
assign n_11978 = ~n_313 & ~n_11977;
assign n_11979 = n_11957 ^ n_11978;
assign n_11980 = x66 ^ n_11978;
assign n_11981 = ~n_11967 & ~n_11979;
assign n_11982 = n_11981 ^ x66;
assign n_11983 = n_11982 ^ x67;
assign n_11984 = n_11882 ^ n_11982;
assign n_11985 = n_11983 & n_11984;
assign n_11986 = n_11985 ^ x67;
assign n_11987 = n_11986 ^ x68;
assign n_11988 = n_11883 ^ n_11986;
assign n_11989 = n_11987 & n_11988;
assign n_11990 = n_11989 ^ x68;
assign n_11991 = n_11990 ^ x69;
assign n_11992 = n_11884 ^ n_11990;
assign n_11993 = n_11991 & n_11992;
assign n_11994 = n_11993 ^ x69;
assign n_11995 = n_11994 ^ x70;
assign n_11996 = n_11885 ^ n_11994;
assign n_11997 = n_11995 & n_11996;
assign n_11998 = n_11997 ^ x70;
assign n_11999 = n_11998 ^ x71;
assign n_12000 = n_11886 ^ n_11998;
assign n_12001 = n_11999 & n_12000;
assign n_12002 = n_12001 ^ x71;
assign n_12003 = n_12002 ^ x72;
assign n_12004 = n_11887 ^ n_12002;
assign n_12005 = n_12003 & n_12004;
assign n_12006 = n_12005 ^ x72;
assign n_12007 = n_12006 ^ n_11878;
assign n_12008 = n_12006 ^ x73;
assign n_12009 = ~n_11942 & n_12007;
assign n_12010 = n_12009 ^ x73;
assign n_12011 = n_12010 ^ n_11877;
assign n_12012 = n_12010 ^ x74;
assign n_12013 = ~n_11941 & n_12011;
assign n_12014 = n_12013 ^ x74;
assign n_12015 = n_12014 ^ x75;
assign n_12016 = n_11888 ^ n_12014;
assign n_12017 = n_12015 & n_12016;
assign n_12018 = n_12017 ^ x75;
assign n_12019 = n_12018 ^ x76;
assign n_12020 = n_11889 ^ n_12018;
assign n_12021 = n_12019 & n_12020;
assign n_12022 = n_12021 ^ x76;
assign n_12023 = n_12022 ^ x77;
assign n_12024 = n_11890 ^ n_12022;
assign n_12025 = n_12023 & n_12024;
assign n_12026 = n_12025 ^ x77;
assign n_12027 = n_12026 ^ x78;
assign n_12028 = n_11891 ^ n_12026;
assign n_12029 = n_12027 & n_12028;
assign n_12030 = n_12029 ^ x78;
assign n_12031 = n_12030 ^ x79;
assign n_12032 = n_11892 ^ n_12030;
assign n_12033 = n_12031 & n_12032;
assign n_12034 = n_12033 ^ x79;
assign n_12035 = n_12034 ^ n_11876;
assign n_12036 = n_12034 ^ x80;
assign n_12037 = ~n_11940 & n_12035;
assign n_12038 = n_12037 ^ x80;
assign n_12039 = n_12038 ^ n_11875;
assign n_12040 = n_12038 ^ x81;
assign n_12041 = ~n_11939 & n_12039;
assign n_12042 = n_12041 ^ x81;
assign n_12043 = n_12042 ^ x82;
assign n_12044 = n_12042 ^ n_11874;
assign n_12045 = n_11965 & n_12042;
assign n_12046 = n_12043 & n_12044;
assign n_12047 = ~n_11973 & ~n_12045;
assign n_12048 = n_12046 ^ x82;
assign n_12049 = x84 ^ n_12047;
assign n_12050 = n_11894 ^ n_12047;
assign n_12051 = n_11969 & ~n_12047;
assign n_12052 = n_12048 ^ x83;
assign n_12053 = ~n_12049 & ~n_12050;
assign n_12054 = ~n_11975 & ~n_12051;
assign n_12055 = n_12053 ^ x84;
assign n_12056 = x86 ^ n_12054;
assign n_12057 = n_11895 ^ n_12054;
assign n_12058 = n_12055 ^ x85;
assign n_12059 = ~n_12056 & ~n_12057;
assign n_12060 = n_12059 ^ x86;
assign n_12061 = n_12060 ^ x87;
assign n_12062 = n_11896 ^ n_12060;
assign n_12063 = n_12061 & n_12062;
assign n_12064 = n_12063 ^ x87;
assign n_12065 = n_12064 ^ x88;
assign n_12066 = n_11897 ^ n_12064;
assign n_12067 = n_12065 & n_12066;
assign n_12068 = n_12067 ^ x88;
assign n_12069 = n_12068 ^ x89;
assign n_12070 = n_11898 ^ n_12068;
assign n_12071 = n_12069 & n_12070;
assign n_12072 = n_12071 ^ x89;
assign n_12073 = n_12072 ^ x90;
assign n_12074 = n_11899 ^ n_12072;
assign n_12075 = n_12073 & n_12074;
assign n_12076 = n_12075 ^ x90;
assign n_12077 = n_12076 ^ x91;
assign n_12078 = n_12076 ^ n_11872;
assign n_12079 = n_11963 & n_12076;
assign n_12080 = n_12077 & n_12078;
assign n_12081 = ~n_11972 & ~n_12079;
assign n_12082 = n_12080 ^ x91;
assign n_12083 = x93 ^ n_12081;
assign n_12084 = n_11900 ^ n_12081;
assign n_12085 = n_12082 ^ x92;
assign n_12086 = ~n_12083 & ~n_12084;
assign n_12087 = n_12086 ^ x93;
assign n_12088 = n_12087 ^ x94;
assign n_12089 = n_11901 ^ n_12087;
assign n_12090 = n_12088 & n_12089;
assign n_12091 = n_12090 ^ x94;
assign n_12092 = n_12091 ^ x95;
assign n_12093 = n_11902 ^ n_12091;
assign n_12094 = n_12092 & n_12093;
assign n_12095 = n_12094 ^ x95;
assign n_12096 = n_12095 ^ x96;
assign n_12097 = n_11903 ^ n_12095;
assign n_12098 = n_12096 & n_12097;
assign n_12099 = n_12098 ^ x96;
assign n_12100 = n_12099 ^ x97;
assign n_12101 = n_11904 ^ n_12099;
assign n_12102 = n_12100 & n_12101;
assign n_12103 = n_12102 ^ x97;
assign n_12104 = n_12103 ^ x98;
assign n_12105 = n_11905 ^ n_12103;
assign n_12106 = n_12104 & n_12105;
assign n_12107 = n_12106 ^ x98;
assign n_12108 = n_12107 ^ x99;
assign n_12109 = n_11906 ^ n_12107;
assign n_12110 = n_12108 & n_12109;
assign n_12111 = n_12110 ^ x99;
assign n_12112 = n_12111 ^ n_11870;
assign n_12113 = n_12111 ^ x100;
assign n_12114 = ~n_11930 & n_12112;
assign n_12115 = n_12114 ^ x100;
assign n_12116 = n_12115 ^ n_11869;
assign n_12117 = n_12115 ^ x101;
assign n_12118 = ~n_11929 & n_12116;
assign n_12119 = n_12118 ^ x101;
assign n_12120 = n_12119 ^ x102;
assign n_12121 = n_11907 ^ n_12119;
assign n_12122 = n_12120 & n_12121;
assign n_12123 = n_12122 ^ x102;
assign n_12124 = n_12123 ^ x103;
assign n_12125 = n_11908 ^ n_12123;
assign n_12126 = n_12124 & n_12125;
assign n_12127 = n_12126 ^ x103;
assign n_12128 = n_12127 ^ x104;
assign n_12129 = n_11909 ^ n_12127;
assign n_12130 = n_12128 & n_12129;
assign n_12131 = n_12130 ^ x104;
assign n_12132 = n_12131 ^ x105;
assign n_12133 = n_11910 ^ n_12131;
assign n_12134 = n_12132 & n_12133;
assign n_12135 = n_12134 ^ x105;
assign n_12136 = n_12135 ^ x106;
assign n_12137 = n_11911 ^ n_12135;
assign n_12138 = n_12136 & n_12137;
assign n_12139 = n_12138 ^ x106;
assign n_12140 = n_12139 ^ x107;
assign n_12141 = n_11912 ^ n_12139;
assign n_12142 = n_12140 & n_12141;
assign n_12143 = n_12142 ^ x107;
assign n_12144 = n_12143 ^ x108;
assign n_12145 = n_12143 ^ n_11868;
assign n_12146 = n_11961 & n_12143;
assign n_12147 = n_12144 & n_12145;
assign n_12148 = ~n_11971 & ~n_12146;
assign n_12149 = n_12147 ^ x108;
assign n_12150 = x110 ^ n_12148;
assign n_12151 = n_11913 ^ n_12148;
assign n_12152 = n_12149 ^ x109;
assign n_12153 = ~n_12150 & ~n_12151;
assign n_12154 = n_12153 ^ x110;
assign n_12155 = n_12154 ^ x111;
assign n_12156 = n_11914 ^ n_12154;
assign n_12157 = n_12155 & n_12156;
assign n_12158 = n_12157 ^ x111;
assign n_12159 = n_12158 ^ x112;
assign n_12160 = n_11915 ^ n_12158;
assign n_12161 = n_12159 & n_12160;
assign n_12162 = n_12161 ^ x112;
assign n_12163 = n_12162 ^ x113;
assign n_12164 = n_11916 ^ n_12162;
assign n_12165 = n_12163 & n_12164;
assign n_12166 = n_12165 ^ x113;
assign n_12167 = n_12166 ^ n_11867;
assign n_12168 = n_12166 ^ x114;
assign n_12169 = ~n_11926 & n_12167;
assign n_12170 = n_12169 ^ x114;
assign n_12171 = n_12170 ^ n_11866;
assign n_12172 = n_12170 ^ x115;
assign n_12173 = ~n_11925 & n_12171;
assign n_12174 = n_12173 ^ x115;
assign n_12175 = n_12174 ^ x116;
assign n_12176 = n_11917 ^ n_12174;
assign n_12177 = n_12175 & n_12176;
assign n_12178 = n_12177 ^ x116;
assign n_12179 = n_12178 ^ x117;
assign n_12180 = n_11918 ^ n_12178;
assign n_12181 = n_12179 & n_12180;
assign n_12182 = n_12181 ^ x117;
assign n_12183 = n_12182 ^ x118;
assign n_12184 = n_11919 ^ n_12182;
assign n_12185 = n_12183 & n_12184;
assign n_12186 = n_12185 ^ x118;
assign n_12187 = n_12186 ^ x119;
assign n_12188 = n_11920 ^ n_12186;
assign n_12189 = n_12187 & n_12188;
assign n_12190 = n_12189 ^ x119;
assign n_12191 = n_12190 ^ x120;
assign n_12192 = n_11921 ^ n_12190;
assign n_12193 = n_12191 & n_12192;
assign n_12194 = n_12193 ^ x120;
assign n_12195 = n_12194 ^ x121;
assign n_12196 = n_11922 ^ n_12194;
assign n_12197 = n_12195 & n_12196;
assign n_12198 = n_12197 ^ x121;
assign n_12199 = n_12198 ^ n_11865;
assign n_12200 = n_12198 ^ x122;
assign n_12201 = ~n_11924 & n_12199;
assign n_12202 = n_12201 ^ x122;
assign n_12203 = n_12202 ^ x123;
assign n_12204 = n_12203 & n_11800;
assign n_12205 = ~x123 & ~n_12203;
assign n_12206 = n_295 & n_12204;
assign n_12207 = n_12205 ^ n_12204;
assign n_12208 = n_12206 ^ n_11800;
assign n_12209 = n_295 & n_12207;
assign n_12210 = ~x124 ^ n_12208;
assign n_12211 = n_12159 & n_12209;
assign n_12212 = n_12155 & n_12209;
assign n_12213 = n_12092 & n_12209;
assign n_12214 = n_12088 & n_12209;
assign n_12215 = n_12065 & n_12209;
assign n_12216 = n_12061 & n_12209;
assign n_12217 = n_12012 & n_12209;
assign n_12218 = n_12008 & n_12209;
assign n_12219 = x64 ^ n_12209;
assign n_12220 = ~x64 & ~n_12209;
assign n_12221 = x4 & n_12209;
assign n_12222 = ~n_60 & n_12209;
assign n_12223 = ~n_11980 & n_12209;
assign n_12224 = n_11983 & n_12209;
assign n_12225 = n_11987 & n_12209;
assign n_12226 = n_11991 & n_12209;
assign n_12227 = n_11995 & n_12209;
assign n_12228 = n_11999 & n_12209;
assign n_12229 = n_12003 & n_12209;
assign n_12230 = n_12015 & n_12209;
assign n_12231 = n_12019 & n_12209;
assign n_12232 = n_12023 & n_12209;
assign n_12233 = n_12027 & n_12209;
assign n_12234 = n_12031 & n_12209;
assign n_12235 = n_12036 & n_12209;
assign n_12236 = n_12040 & n_12209;
assign n_12237 = n_12043 & n_12209;
assign n_12238 = ~n_12049 & n_12209;
assign n_12239 = ~n_12056 & n_12209;
assign n_12240 = n_12069 & n_12209;
assign n_12241 = n_12073 & n_12209;
assign n_12242 = n_12077 & n_12209;
assign n_12243 = ~n_12083 & n_12209;
assign n_12244 = n_12096 & n_12209;
assign n_12245 = n_12100 & n_12209;
assign n_12246 = n_12104 & n_12209;
assign n_12247 = n_12108 & n_12209;
assign n_12248 = n_12113 & n_12209;
assign n_12249 = n_12117 & n_12209;
assign n_12250 = n_12120 & n_12209;
assign n_12251 = n_12124 & n_12209;
assign n_12252 = n_12128 & n_12209;
assign n_12253 = n_12132 & n_12209;
assign n_12254 = n_12136 & n_12209;
assign n_12255 = n_12140 & n_12209;
assign n_12256 = n_12144 & n_12209;
assign n_12257 = ~n_12150 & n_12209;
assign n_12258 = n_12163 & n_12209;
assign n_12259 = n_12168 & n_12209;
assign n_12260 = n_12172 & n_12209;
assign n_12261 = n_12175 & n_12209;
assign n_12262 = n_12179 & n_12209;
assign n_12263 = n_12183 & n_12209;
assign n_12264 = n_12187 & n_12209;
assign n_12265 = n_12191 & n_12209;
assign n_12266 = n_12195 & n_12209;
assign n_12267 = n_12200 & n_12209;
assign y4 = n_12209;
assign n_12268 = n_12052 & n_12209;
assign n_12269 = n_12058 & n_12209;
assign n_12270 = n_12085 & n_12209;
assign n_12271 = n_12152 & n_12209;
assign n_12272 = n_12211 ^ n_11915;
assign n_12273 = n_12212 ^ n_11914;
assign n_12274 = n_12213 ^ n_11902;
assign n_12275 = n_12214 ^ n_11901;
assign n_12276 = n_12215 ^ n_11897;
assign n_12277 = n_12216 ^ n_11896;
assign n_12278 = n_12217 ^ n_11877;
assign n_12279 = n_12218 ^ n_11878;
assign n_12280 = n_12219 ^ n_12220;
assign n_12281 = n_11863 ^ n_12220;
assign n_12282 = n_46 & n_12221;
assign n_12283 = ~n_107 & n_12222;
assign n_12284 = n_12223 ^ n_11957;
assign n_12285 = n_12224 ^ n_11882;
assign n_12286 = n_12225 ^ n_11883;
assign n_12287 = n_12226 ^ n_11884;
assign n_12288 = n_12227 ^ n_11885;
assign n_12289 = n_12228 ^ n_11886;
assign n_12290 = n_12229 ^ n_11887;
assign n_12291 = n_12230 ^ n_11888;
assign n_12292 = n_12231 ^ n_11889;
assign n_12293 = n_12232 ^ n_11890;
assign n_12294 = n_12233 ^ n_11891;
assign n_12295 = n_12234 ^ n_11892;
assign n_12296 = n_12235 ^ n_11876;
assign n_12297 = n_12236 ^ n_11875;
assign n_12298 = n_12237 ^ n_11874;
assign n_12299 = n_12238 ^ n_11894;
assign n_12300 = n_12239 ^ n_11895;
assign n_12301 = n_12240 ^ n_11898;
assign n_12302 = n_12241 ^ n_11899;
assign n_12303 = n_12242 ^ n_11872;
assign n_12304 = n_12243 ^ n_11900;
assign n_12305 = n_12244 ^ n_11903;
assign n_12306 = n_12245 ^ n_11904;
assign n_12307 = n_12246 ^ n_11905;
assign n_12308 = n_12247 ^ n_11906;
assign n_12309 = n_12248 ^ n_11870;
assign n_12310 = n_12249 ^ n_11869;
assign n_12311 = n_12250 ^ n_11907;
assign n_12312 = n_12251 ^ n_11908;
assign n_12313 = n_12252 ^ n_11909;
assign n_12314 = n_12253 ^ n_11910;
assign n_12315 = n_12254 ^ n_11911;
assign n_12316 = n_12255 ^ n_11912;
assign n_12317 = n_12256 ^ n_11868;
assign n_12318 = n_12257 ^ n_11913;
assign n_12319 = n_12258 ^ n_11916;
assign n_12320 = n_12259 ^ n_11867;
assign n_12321 = n_12260 ^ n_11866;
assign n_12322 = n_12261 ^ n_11917;
assign n_12323 = n_12262 ^ n_11918;
assign n_12324 = n_12263 ^ n_11919;
assign n_12325 = n_12264 ^ n_11920;
assign n_12326 = n_12265 ^ n_11921;
assign n_12327 = n_12266 ^ n_11922;
assign n_12328 = n_12267 ^ n_11865;
assign n_12329 = n_11873 ^ n_12268;
assign n_12330 = n_11893 ^ n_12269;
assign n_12331 = n_11871 ^ n_12270;
assign n_12332 = n_11923 ^ n_12271;
assign n_12333 = n_12272 ^ x113;
assign n_12334 = n_12273 ^ x112;
assign n_12335 = ~x96 ^ n_12274;
assign n_12336 = n_12274 ^ x96;
assign n_12337 = n_12275 ^ x95;
assign n_12338 = x95 & ~n_12275;
assign n_12339 = ~x89 ^ n_12276;
assign n_12340 = n_12276 ^ x89;
assign n_12341 = n_12277 ^ x88;
assign n_12342 = x88 & ~n_12277;
assign n_12343 = ~x75 ^ n_12278;
assign n_12344 = n_12278 ^ x75;
assign n_12345 = n_12279 ^ x74;
assign n_12346 = x74 & ~n_12279;
assign n_12347 = n_12280 ^ x4;
assign n_12348 = n_12281 ^ n_12283;
assign n_12349 = n_12337 ^ n_12338;
assign n_12350 = n_12338 ^ n_12274;
assign n_12351 = n_12341 ^ n_12342;
assign n_12352 = n_12342 ^ n_12276;
assign n_12353 = n_12345 ^ n_12346;
assign n_12354 = n_12346 ^ n_12278;
assign n_12355 = n_12347 ^ n_38;
assign n_12356 = n_12347 ^ x65;
assign n_12357 = ~n_12347 & ~n_239;
assign n_12358 = n_12348 ^ n_12282;
assign n_12359 = n_12335 & ~n_12349;
assign n_12360 = ~n_12336 & n_12350;
assign n_12361 = n_12339 & ~n_12351;
assign n_12362 = ~n_12340 & n_12352;
assign n_12363 = n_12343 & ~n_12353;
assign n_12364 = ~n_12344 & n_12354;
assign n_12365 = n_173 & ~n_12355;
assign n_12366 = ~n_111 ^ n_12356;
assign n_12367 = n_38 & n_12356;
assign n_12368 = n_12358 ^ x5;
assign n_12369 = n_12360 ^ x96;
assign n_12370 = n_12362 ^ x89;
assign n_12371 = n_12364 ^ x75;
assign n_12372 = n_12365 ^ x65;
assign n_12373 = ~n_241 & n_12367;
assign n_12374 = n_12372 ^ x66;
assign n_12375 = n_12368 ^ n_12372;
assign n_12376 = n_288 ^ n_12373;
assign n_12377 = n_12374 & ~n_12375;
assign n_12378 = n_12377 ^ x66;
assign n_12379 = n_12378 ^ x67;
assign n_12380 = n_12284 ^ n_12378;
assign n_12381 = n_12379 & n_12380;
assign n_12382 = n_12381 ^ x67;
assign n_12383 = n_12382 ^ x68;
assign n_12384 = n_12285 ^ n_12382;
assign n_12385 = n_12383 & n_12384;
assign n_12386 = n_12385 ^ x68;
assign n_12387 = n_12386 ^ x69;
assign n_12388 = n_12286 ^ n_12386;
assign n_12389 = n_12387 & n_12388;
assign n_12390 = n_12389 ^ x69;
assign n_12391 = n_12390 ^ x70;
assign n_12392 = n_12287 ^ n_12390;
assign n_12393 = n_12391 & n_12392;
assign n_12394 = n_12393 ^ x70;
assign n_12395 = n_12394 ^ x71;
assign n_12396 = n_12288 ^ n_12394;
assign n_12397 = n_12395 & n_12396;
assign n_12398 = n_12397 ^ x71;
assign n_12399 = n_12398 ^ x72;
assign n_12400 = n_12289 ^ n_12398;
assign n_12401 = n_12399 & n_12400;
assign n_12402 = n_12401 ^ x72;
assign n_12403 = n_12402 ^ x73;
assign n_12404 = n_12290 ^ n_12402;
assign n_12405 = n_12403 & n_12404;
assign n_12406 = n_12405 ^ x73;
assign n_12407 = n_12406 ^ x74;
assign n_12408 = n_12406 ^ n_12279;
assign n_12409 = n_12363 & n_12406;
assign n_12410 = n_12407 & n_12408;
assign n_12411 = ~n_12371 & ~n_12409;
assign n_12412 = n_12410 ^ x74;
assign n_12413 = x76 ^ n_12411;
assign n_12414 = n_12291 ^ n_12411;
assign n_12415 = n_12412 ^ x75;
assign n_12416 = ~n_12413 & ~n_12414;
assign n_12417 = n_12416 ^ x76;
assign n_12418 = n_12417 ^ x77;
assign n_12419 = n_12292 ^ n_12417;
assign n_12420 = n_12418 & n_12419;
assign n_12421 = n_12420 ^ x77;
assign n_12422 = n_12421 ^ x78;
assign n_12423 = n_12293 ^ n_12421;
assign n_12424 = n_12422 & n_12423;
assign n_12425 = n_12424 ^ x78;
assign n_12426 = n_12425 ^ x79;
assign n_12427 = n_12294 ^ n_12425;
assign n_12428 = n_12426 & n_12427;
assign n_12429 = n_12428 ^ x79;
assign n_12430 = n_12429 ^ x80;
assign n_12431 = n_12295 ^ n_12429;
assign n_12432 = n_12430 & n_12431;
assign n_12433 = n_12432 ^ x80;
assign n_12434 = n_12433 ^ x81;
assign n_12435 = n_12296 ^ n_12433;
assign n_12436 = n_12434 & n_12435;
assign n_12437 = n_12436 ^ x81;
assign n_12438 = n_12437 ^ x82;
assign n_12439 = n_12297 ^ n_12437;
assign n_12440 = n_12438 & n_12439;
assign n_12441 = n_12440 ^ x82;
assign n_12442 = n_12441 ^ x83;
assign n_12443 = n_12298 ^ n_12441;
assign n_12444 = n_12442 & n_12443;
assign n_12445 = n_12444 ^ x83;
assign n_12446 = n_12445 ^ x84;
assign n_12447 = n_12329 ^ n_12445;
assign n_12448 = n_12446 & n_12447;
assign n_12449 = n_12448 ^ x84;
assign n_12450 = n_12449 ^ x85;
assign n_12451 = n_12299 ^ n_12449;
assign n_12452 = n_12450 & n_12451;
assign n_12453 = n_12452 ^ x85;
assign n_12454 = n_12453 ^ x86;
assign n_12455 = n_12330 ^ n_12453;
assign n_12456 = n_12454 & n_12455;
assign n_12457 = n_12456 ^ x86;
assign n_12458 = n_12457 ^ x87;
assign n_12459 = n_12300 ^ n_12457;
assign n_12460 = n_12458 & n_12459;
assign n_12461 = n_12460 ^ x87;
assign n_12462 = n_12461 ^ x88;
assign n_12463 = n_12461 ^ n_12277;
assign n_12464 = n_12361 & n_12461;
assign n_12465 = n_12462 & n_12463;
assign n_12466 = ~n_12370 & ~n_12464;
assign n_12467 = n_12465 ^ x88;
assign n_12468 = x90 ^ n_12466;
assign n_12469 = n_12301 ^ n_12466;
assign n_12470 = n_12467 ^ x89;
assign n_12471 = ~n_12468 & ~n_12469;
assign n_12472 = n_12471 ^ x90;
assign n_12473 = n_12472 ^ x91;
assign n_12474 = n_12302 ^ n_12472;
assign n_12475 = n_12473 & n_12474;
assign n_12476 = n_12475 ^ x91;
assign n_12477 = n_12476 ^ x92;
assign n_12478 = n_12303 ^ n_12476;
assign n_12479 = n_12477 & n_12478;
assign n_12480 = n_12479 ^ x92;
assign n_12481 = n_12480 ^ x93;
assign n_12482 = n_12331 ^ n_12480;
assign n_12483 = n_12481 & ~n_12482;
assign n_12484 = n_12483 ^ x93;
assign n_12485 = n_12484 ^ x94;
assign n_12486 = n_12304 ^ n_12484;
assign n_12487 = n_12485 & n_12486;
assign n_12488 = n_12487 ^ x94;
assign n_12489 = n_12488 ^ x95;
assign n_12490 = n_12488 ^ n_12275;
assign n_12491 = n_12359 & n_12488;
assign n_12492 = n_12489 & n_12490;
assign n_12493 = ~n_12369 & ~n_12491;
assign n_12494 = n_12492 ^ x95;
assign n_12495 = x97 ^ n_12493;
assign n_12496 = n_12305 ^ n_12493;
assign n_12497 = n_12494 ^ x96;
assign n_12498 = ~n_12495 & ~n_12496;
assign n_12499 = n_12498 ^ x97;
assign n_12500 = n_12499 ^ x98;
assign n_12501 = n_12306 ^ n_12499;
assign n_12502 = n_12500 & n_12501;
assign n_12503 = n_12502 ^ x98;
assign n_12504 = n_12503 ^ x99;
assign n_12505 = n_12307 ^ n_12503;
assign n_12506 = n_12504 & n_12505;
assign n_12507 = n_12506 ^ x99;
assign n_12508 = n_12507 ^ x100;
assign n_12509 = n_12308 ^ n_12507;
assign n_12510 = n_12508 & n_12509;
assign n_12511 = n_12510 ^ x100;
assign n_12512 = n_12511 ^ x101;
assign n_12513 = n_12309 ^ n_12511;
assign n_12514 = n_12512 & n_12513;
assign n_12515 = n_12514 ^ x101;
assign n_12516 = n_12515 ^ x102;
assign n_12517 = n_12310 ^ n_12515;
assign n_12518 = n_12516 & n_12517;
assign n_12519 = n_12518 ^ x102;
assign n_12520 = n_12519 ^ x103;
assign n_12521 = n_12311 ^ n_12519;
assign n_12522 = n_12520 & n_12521;
assign n_12523 = n_12522 ^ x103;
assign n_12524 = n_12523 ^ x104;
assign n_12525 = n_12312 ^ n_12523;
assign n_12526 = n_12524 & n_12525;
assign n_12527 = n_12526 ^ x104;
assign n_12528 = n_12527 ^ x105;
assign n_12529 = n_12313 ^ n_12527;
assign n_12530 = n_12528 & n_12529;
assign n_12531 = n_12530 ^ x105;
assign n_12532 = n_12531 ^ x106;
assign n_12533 = n_12314 ^ n_12531;
assign n_12534 = n_12532 & n_12533;
assign n_12535 = n_12534 ^ x106;
assign n_12536 = n_12535 ^ x107;
assign n_12537 = n_12315 ^ n_12535;
assign n_12538 = n_12536 & n_12537;
assign n_12539 = n_12538 ^ x107;
assign n_12540 = n_12539 ^ x108;
assign n_12541 = n_12316 ^ n_12539;
assign n_12542 = n_12540 & n_12541;
assign n_12543 = n_12542 ^ x108;
assign n_12544 = n_12543 ^ x109;
assign n_12545 = n_12317 ^ n_12543;
assign n_12546 = n_12544 & n_12545;
assign n_12547 = n_12546 ^ x109;
assign n_12548 = n_12547 ^ x110;
assign n_12549 = n_12332 ^ n_12547;
assign n_12550 = n_12548 & n_12549;
assign n_12551 = n_12550 ^ x110;
assign n_12552 = n_12551 ^ x111;
assign n_12553 = n_12318 ^ n_12551;
assign n_12554 = n_12552 & n_12553;
assign n_12555 = n_12554 ^ x111;
assign n_12556 = n_12555 ^ n_12273;
assign n_12557 = n_12555 ^ x112;
assign n_12558 = ~n_12334 & n_12556;
assign n_12559 = n_12558 ^ x112;
assign n_12560 = n_12559 ^ n_12272;
assign n_12561 = n_12559 ^ x113;
assign n_12562 = ~n_12333 & n_12560;
assign n_12563 = n_12562 ^ x113;
assign n_12564 = n_12563 ^ x114;
assign n_12565 = n_12319 ^ n_12563;
assign n_12566 = n_12564 & n_12565;
assign n_12567 = n_12566 ^ x114;
assign n_12568 = n_12567 ^ x115;
assign n_12569 = n_12320 ^ n_12567;
assign n_12570 = n_12568 & n_12569;
assign n_12571 = n_12570 ^ x115;
assign n_12572 = n_12571 ^ x116;
assign n_12573 = n_12321 ^ n_12571;
assign n_12574 = n_12572 & n_12573;
assign n_12575 = n_12574 ^ x116;
assign n_12576 = n_12575 ^ x117;
assign n_12577 = n_12322 ^ n_12575;
assign n_12578 = n_12576 & n_12577;
assign n_12579 = n_12578 ^ x117;
assign n_12580 = n_12579 ^ x118;
assign n_12581 = n_12323 ^ n_12579;
assign n_12582 = n_12580 & n_12581;
assign n_12583 = n_12582 ^ x118;
assign n_12584 = n_12583 ^ x119;
assign n_12585 = n_12324 ^ n_12583;
assign n_12586 = n_12584 & n_12585;
assign n_12587 = n_12586 ^ x119;
assign n_12588 = n_12587 ^ x120;
assign n_12589 = n_12325 ^ n_12587;
assign n_12590 = n_12588 & n_12589;
assign n_12591 = n_12590 ^ x120;
assign n_12592 = n_12591 ^ x121;
assign n_12593 = n_12326 ^ n_12591;
assign n_12594 = n_12592 & n_12593;
assign n_12595 = n_12594 ^ x121;
assign n_12596 = n_12595 ^ x122;
assign n_12597 = n_12327 ^ n_12595;
assign n_12598 = n_12596 & n_12597;
assign n_12599 = n_12598 ^ x122;
assign n_12600 = n_12599 ^ x123;
assign n_12601 = n_12328 ^ n_12599;
assign n_12602 = n_12600 & n_12601;
assign n_12603 = n_12602 ^ x123;
assign n_12604 = n_12210 & n_12603;
assign n_12605 = n_12603 ^ x124;
assign n_12606 = ~n_12604 & n_11184;
assign n_12607 = n_12208 & n_12605;
assign n_12608 = x64 & n_12606;
assign n_12609 = n_12347 ^ n_12606;
assign n_12610 = x3 & n_12606;
assign n_12611 = n_110 ^ ~n_12606;
assign n_12612 = n_174 & n_12606;
assign n_12613 = n_12374 & n_12606;
assign n_12614 = n_12568 & n_12606;
assign n_12615 = n_12564 & n_12606;
assign n_12616 = n_12516 & n_12606;
assign n_12617 = n_12512 & n_12606;
assign n_12618 = n_12504 & n_12606;
assign n_12619 = n_12500 & n_12606;
assign n_12620 = n_12481 & n_12606;
assign n_12621 = n_12477 & n_12606;
assign n_12622 = n_12387 & n_12606;
assign n_12623 = n_12379 & n_12606;
assign n_12624 = n_12383 & n_12606;
assign n_12625 = n_12391 & n_12606;
assign n_12626 = n_12395 & n_12606;
assign n_12627 = n_12399 & n_12606;
assign n_12628 = n_12403 & n_12606;
assign n_12629 = n_12407 & n_12606;
assign n_12630 = ~n_12413 & n_12606;
assign n_12631 = n_12418 & n_12606;
assign n_12632 = n_12422 & n_12606;
assign n_12633 = n_12426 & n_12606;
assign n_12634 = n_12430 & n_12606;
assign n_12635 = n_12434 & n_12606;
assign n_12636 = n_12438 & n_12606;
assign n_12637 = n_12442 & n_12606;
assign n_12638 = n_12446 & n_12606;
assign n_12639 = n_12450 & n_12606;
assign n_12640 = n_12454 & n_12606;
assign n_12641 = n_12458 & n_12606;
assign n_12642 = n_12462 & n_12606;
assign n_12643 = ~n_12468 & n_12606;
assign n_12644 = n_12473 & n_12606;
assign n_12645 = n_12485 & n_12606;
assign n_12646 = n_12489 & n_12606;
assign n_12647 = ~n_12495 & n_12606;
assign n_12648 = n_12508 & n_12606;
assign n_12649 = n_12520 & n_12606;
assign n_12650 = n_12524 & n_12606;
assign n_12651 = n_12528 & n_12606;
assign n_12652 = n_12532 & n_12606;
assign n_12653 = n_12536 & n_12606;
assign n_12654 = n_12540 & n_12606;
assign n_12655 = n_12544 & n_12606;
assign n_12656 = n_12548 & n_12606;
assign n_12657 = n_12552 & n_12606;
assign n_12658 = n_12557 & n_12606;
assign n_12659 = n_12561 & n_12606;
assign n_12660 = n_12572 & n_12606;
assign n_12661 = n_12576 & n_12606;
assign n_12662 = n_12580 & n_12606;
assign n_12663 = n_12584 & n_12606;
assign n_12664 = n_12588 & n_12606;
assign n_12665 = n_12592 & n_12606;
assign n_12666 = n_12596 & n_12606;
assign n_12667 = n_12600 & n_12606;
assign y3 = n_12606;
assign n_12668 = n_0 & ~n_12606;
assign n_12669 = n_12376 & n_12606;
assign n_12670 = n_12415 & n_12606;
assign n_12671 = n_12470 & n_12606;
assign n_12672 = n_12497 & n_12606;
assign n_12673 = n_248 & n_12607;
assign n_12674 = ~n_12608 & n_239;
assign n_12675 = n_12610 & ~n_111;
assign n_12676 = n_12611 & n_39;
assign n_12677 = n_12612 ^ n_256;
assign n_12678 = ~n_12612 & n_12357;
assign n_12679 = n_12613 ^ n_12368;
assign n_12680 = n_12614 ^ n_12320;
assign n_12681 = n_12615 ^ n_12319;
assign n_12682 = n_12616 ^ n_12310;
assign n_12683 = n_12617 ^ n_12309;
assign n_12684 = n_12618 ^ n_12307;
assign n_12685 = n_12619 ^ n_12306;
assign n_12686 = n_12620 ^ n_12331;
assign n_12687 = n_12621 ^ n_12303;
assign n_12688 = n_12622 ^ n_12286;
assign n_12689 = n_12623 ^ n_12284;
assign n_12690 = n_12624 ^ n_12285;
assign n_12691 = n_12625 ^ n_12287;
assign n_12692 = n_12626 ^ n_12288;
assign n_12693 = n_12627 ^ n_12289;
assign n_12694 = n_12628 ^ n_12290;
assign n_12695 = n_12629 ^ n_12279;
assign n_12696 = n_12630 ^ n_12291;
assign n_12697 = n_12631 ^ n_12292;
assign n_12698 = n_12632 ^ n_12293;
assign n_12699 = n_12633 ^ n_12294;
assign n_12700 = n_12634 ^ n_12295;
assign n_12701 = n_12635 ^ n_12296;
assign n_12702 = n_12636 ^ n_12297;
assign n_12703 = n_12637 ^ n_12298;
assign n_12704 = n_12638 ^ n_12329;
assign n_12705 = n_12639 ^ n_12299;
assign n_12706 = n_12640 ^ n_12330;
assign n_12707 = n_12641 ^ n_12300;
assign n_12708 = n_12642 ^ n_12277;
assign n_12709 = n_12643 ^ n_12301;
assign n_12710 = n_12644 ^ n_12302;
assign n_12711 = n_12645 ^ n_12304;
assign n_12712 = n_12646 ^ n_12275;
assign n_12713 = n_12647 ^ n_12305;
assign n_12714 = n_12648 ^ n_12308;
assign n_12715 = n_12649 ^ n_12311;
assign n_12716 = n_12650 ^ n_12312;
assign n_12717 = n_12651 ^ n_12313;
assign n_12718 = n_12652 ^ n_12314;
assign n_12719 = n_12653 ^ n_12315;
assign n_12720 = n_12654 ^ n_12316;
assign n_12721 = n_12655 ^ n_12317;
assign n_12722 = n_12656 ^ n_12332;
assign n_12723 = n_12657 ^ n_12318;
assign n_12724 = n_12658 ^ n_12273;
assign n_12725 = n_12659 ^ n_12272;
assign n_12726 = n_12660 ^ n_12321;
assign n_12727 = n_12661 ^ n_12322;
assign n_12728 = n_12662 ^ n_12323;
assign n_12729 = n_12663 ^ n_12324;
assign n_12730 = n_12664 ^ n_12325;
assign n_12731 = n_12665 ^ n_12326;
assign n_12732 = n_12666 ^ n_12327;
assign n_12733 = n_12667 ^ n_12328;
assign n_12734 = ~n_241 & ~n_12668;
assign n_12735 = n_12278 ^ n_12670;
assign n_12736 = n_12276 ^ n_12671;
assign n_12737 = n_12274 ^ n_12672;
assign n_12738 = n_12208 ^ n_12673;
assign n_12739 = n_12674 & n_12609;
assign n_12740 = ~n_12677 ^ n_12347;
assign n_12741 = ~n_12676 & n_12678;
assign n_12742 = ~x116 ^ n_12680;
assign n_12743 = n_12680 ^ x116;
assign n_12744 = n_12681 ^ x115;
assign n_12745 = x115 & ~n_12681;
assign n_12746 = ~x103 ^ n_12682;
assign n_12747 = n_12682 ^ x103;
assign n_12748 = n_12683 ^ x102;
assign n_12749 = x102 & ~n_12683;
assign n_12750 = ~x100 ^ n_12684;
assign n_12751 = n_12684 ^ x100;
assign n_12752 = n_12685 ^ x99;
assign n_12753 = x99 & ~n_12685;
assign n_12754 = n_12686 ^ x94;
assign n_12755 = n_12687 ^ x93;
assign n_12756 = x70 & ~n_12688;
assign n_12757 = ~n_121 ^ n_12691;
assign n_12758 = n_12691 ^ x71;
assign n_12759 = n_12347 & ~n_12734;
assign n_12760 = ~n_12675 & n_12734;
assign n_12761 = n_12738 ^ n_11102;
assign n_12762 = ~x66 & ~n_12739;
assign n_12763 = ~n_12741 ^ ~n_12669;
assign n_12764 = n_12744 ^ n_12745;
assign n_12765 = n_12745 ^ n_12680;
assign n_12766 = n_12748 ^ n_12749;
assign n_12767 = n_12749 ^ n_12682;
assign n_12768 = n_12752 ^ n_12753;
assign n_12769 = n_12753 ^ n_12684;
assign n_12770 = n_12756 ^ n_12691;
assign n_12771 = ~n_12366 ^ n_12759;
assign n_12772 = x64 & ~n_12760;
assign n_12773 = n_12742 & ~n_12764;
assign n_12774 = ~n_12743 & n_12765;
assign n_12775 = n_12746 & ~n_12766;
assign n_12776 = ~n_12747 & n_12767;
assign n_12777 = n_12750 & ~n_12768;
assign n_12778 = ~n_12751 & n_12769;
assign n_12779 = ~n_12758 & n_12770;
assign n_12780 = n_12610 & n_12771;
assign n_12781 = ~n_12674 & ~n_12772;
assign n_12782 = n_12774 ^ x116;
assign n_12783 = n_12776 ^ x103;
assign n_12784 = n_12778 ^ x100;
assign n_12785 = n_12779 ^ x71;
assign n_12786 = n_12780 ^ n_12759;
assign n_12787 = x66 ^ n_12781;
assign n_12788 = x64 & n_12786;
assign n_12789 = n_12762 & ~n_12788;
assign n_12790 = ~n_12763 & ~n_12789;
assign n_12791 = x67 ^ n_12790;
assign n_12792 = n_12679 ^ n_12790;
assign n_12793 = n_12791 & ~n_12792;
assign n_12794 = n_12793 ^ x67;
assign n_12795 = n_12794 ^ x68;
assign n_12796 = n_12689 ^ n_12794;
assign n_12797 = n_12795 & n_12796;
assign n_12798 = n_12797 ^ x68;
assign n_12799 = n_12798 ^ x69;
assign n_12800 = n_12690 ^ n_12798;
assign n_12801 = n_12799 & n_12800;
assign n_12802 = n_12801 ^ x69;
assign n_12803 = ~n_12688 & n_12802;
assign n_12804 = x70 & n_12802;
assign n_12805 = n_12802 ^ x70;
assign n_12806 = x71 & n_12803;
assign n_12807 = n_12756 ^ n_12803;
assign n_12808 = ~n_12803 ^ ~n_12804;
assign n_12809 = ~n_12806 & ~n_12785;
assign n_12810 = n_12807 ^ n_12804;
assign n_12811 = n_12808 & n_12757;
assign n_12812 = n_12810 ^ x71;
assign n_12813 = ~n_12811 & n_12809;
assign n_12814 = x72 ^ n_12813;
assign n_12815 = n_12692 ^ n_12813;
assign n_12816 = ~n_12814 & ~n_12815;
assign n_12817 = n_12816 ^ x72;
assign n_12818 = n_12817 ^ x73;
assign n_12819 = n_12693 ^ n_12817;
assign n_12820 = n_12818 & n_12819;
assign n_12821 = n_12820 ^ x73;
assign n_12822 = n_12821 ^ x74;
assign n_12823 = n_12694 ^ n_12821;
assign n_12824 = n_12822 & n_12823;
assign n_12825 = n_12824 ^ x74;
assign n_12826 = n_12825 ^ x75;
assign n_12827 = n_12695 ^ n_12825;
assign n_12828 = n_12826 & n_12827;
assign n_12829 = n_12828 ^ x75;
assign n_12830 = n_12829 ^ x76;
assign n_12831 = n_12735 ^ n_12829;
assign n_12832 = n_12830 & n_12831;
assign n_12833 = n_12832 ^ x76;
assign n_12834 = n_12833 ^ x77;
assign n_12835 = n_12696 ^ n_12833;
assign n_12836 = n_12834 & n_12835;
assign n_12837 = n_12836 ^ x77;
assign n_12838 = n_12837 ^ x78;
assign n_12839 = n_12697 ^ n_12837;
assign n_12840 = n_12838 & n_12839;
assign n_12841 = n_12840 ^ x78;
assign n_12842 = n_12841 ^ x79;
assign n_12843 = n_12698 ^ n_12841;
assign n_12844 = n_12842 & n_12843;
assign n_12845 = n_12844 ^ x79;
assign n_12846 = n_12845 ^ x80;
assign n_12847 = n_12699 ^ n_12845;
assign n_12848 = n_12846 & n_12847;
assign n_12849 = n_12848 ^ x80;
assign n_12850 = n_12849 ^ x81;
assign n_12851 = n_12700 ^ n_12849;
assign n_12852 = n_12850 & n_12851;
assign n_12853 = n_12852 ^ x81;
assign n_12854 = n_12853 ^ x82;
assign n_12855 = n_12701 ^ n_12853;
assign n_12856 = n_12854 & n_12855;
assign n_12857 = n_12856 ^ x82;
assign n_12858 = n_12857 ^ x83;
assign n_12859 = n_12702 ^ n_12857;
assign n_12860 = n_12858 & n_12859;
assign n_12861 = n_12860 ^ x83;
assign n_12862 = n_12861 ^ x84;
assign n_12863 = n_12703 ^ n_12861;
assign n_12864 = n_12862 & n_12863;
assign n_12865 = n_12864 ^ x84;
assign n_12866 = n_12865 ^ x85;
assign n_12867 = n_12704 ^ n_12865;
assign n_12868 = n_12866 & n_12867;
assign n_12869 = n_12868 ^ x85;
assign n_12870 = n_12869 ^ x86;
assign n_12871 = n_12705 ^ n_12869;
assign n_12872 = n_12870 & n_12871;
assign n_12873 = n_12872 ^ x86;
assign n_12874 = n_12873 ^ x87;
assign n_12875 = n_12706 ^ n_12873;
assign n_12876 = n_12874 & n_12875;
assign n_12877 = n_12876 ^ x87;
assign n_12878 = n_12877 ^ x88;
assign n_12879 = n_12707 ^ n_12877;
assign n_12880 = n_12878 & n_12879;
assign n_12881 = n_12880 ^ x88;
assign n_12882 = n_12881 ^ x89;
assign n_12883 = n_12708 ^ n_12881;
assign n_12884 = n_12882 & n_12883;
assign n_12885 = n_12884 ^ x89;
assign n_12886 = n_12885 ^ x90;
assign n_12887 = n_12736 ^ n_12885;
assign n_12888 = n_12886 & n_12887;
assign n_12889 = n_12888 ^ x90;
assign n_12890 = n_12889 ^ x91;
assign n_12891 = n_12709 ^ n_12889;
assign n_12892 = n_12890 & n_12891;
assign n_12893 = n_12892 ^ x91;
assign n_12894 = n_12893 ^ x92;
assign n_12895 = n_12710 ^ n_12893;
assign n_12896 = n_12894 & n_12895;
assign n_12897 = n_12896 ^ x92;
assign n_12898 = n_12897 ^ n_12687;
assign n_12899 = n_12897 ^ x93;
assign n_12900 = ~n_12755 & n_12898;
assign n_12901 = n_12900 ^ x93;
assign n_12902 = n_12901 ^ n_12686;
assign n_12903 = n_12901 ^ x94;
assign n_12904 = n_12754 & ~n_12902;
assign n_12905 = n_12904 ^ x94;
assign n_12906 = n_12905 ^ x95;
assign n_12907 = n_12711 ^ n_12905;
assign n_12908 = n_12906 & n_12907;
assign n_12909 = n_12908 ^ x95;
assign n_12910 = n_12909 ^ x96;
assign n_12911 = n_12712 ^ n_12909;
assign n_12912 = n_12910 & n_12911;
assign n_12913 = n_12912 ^ x96;
assign n_12914 = n_12913 ^ x97;
assign n_12915 = n_12737 ^ n_12913;
assign n_12916 = n_12914 & n_12915;
assign n_12917 = n_12916 ^ x97;
assign n_12918 = n_12917 ^ x98;
assign n_12919 = n_12713 ^ n_12917;
assign n_12920 = n_12918 & n_12919;
assign n_12921 = n_12920 ^ x98;
assign n_12922 = n_12921 ^ x99;
assign n_12923 = n_12921 ^ n_12685;
assign n_12924 = n_12777 & n_12921;
assign n_12925 = n_12922 & n_12923;
assign n_12926 = ~n_12784 & ~n_12924;
assign n_12927 = n_12925 ^ x99;
assign n_12928 = x101 ^ n_12926;
assign n_12929 = n_12714 ^ n_12926;
assign n_12930 = n_12927 ^ x100;
assign n_12931 = ~n_12928 & ~n_12929;
assign n_12932 = n_12931 ^ x101;
assign n_12933 = n_12932 ^ x102;
assign n_12934 = n_12932 ^ n_12683;
assign n_12935 = n_12775 & n_12932;
assign n_12936 = n_12933 & n_12934;
assign n_12937 = ~n_12783 & ~n_12935;
assign n_12938 = n_12936 ^ x102;
assign n_12939 = x104 ^ n_12937;
assign n_12940 = n_12715 ^ n_12937;
assign n_12941 = n_12938 ^ x103;
assign n_12942 = ~n_12939 & ~n_12940;
assign n_12943 = n_12942 ^ x104;
assign n_12944 = n_12943 ^ x105;
assign n_12945 = n_12716 ^ n_12943;
assign n_12946 = n_12944 & n_12945;
assign n_12947 = n_12946 ^ x105;
assign n_12948 = n_12947 ^ x106;
assign n_12949 = n_12717 ^ n_12947;
assign n_12950 = n_12948 & n_12949;
assign n_12951 = n_12950 ^ x106;
assign n_12952 = n_12951 ^ x107;
assign n_12953 = n_12718 ^ n_12951;
assign n_12954 = n_12952 & n_12953;
assign n_12955 = n_12954 ^ x107;
assign n_12956 = n_12955 ^ x108;
assign n_12957 = n_12719 ^ n_12955;
assign n_12958 = n_12956 & n_12957;
assign n_12959 = n_12958 ^ x108;
assign n_12960 = n_12959 ^ x109;
assign n_12961 = n_12720 ^ n_12959;
assign n_12962 = n_12960 & n_12961;
assign n_12963 = n_12962 ^ x109;
assign n_12964 = n_12963 ^ x110;
assign n_12965 = n_12721 ^ n_12963;
assign n_12966 = n_12964 & n_12965;
assign n_12967 = n_12966 ^ x110;
assign n_12968 = n_12967 ^ x111;
assign n_12969 = n_12722 ^ n_12967;
assign n_12970 = n_12968 & n_12969;
assign n_12971 = n_12970 ^ x111;
assign n_12972 = n_12971 ^ x112;
assign n_12973 = n_12723 ^ n_12971;
assign n_12974 = n_12972 & n_12973;
assign n_12975 = n_12974 ^ x112;
assign n_12976 = n_12975 ^ x113;
assign n_12977 = n_12724 ^ n_12975;
assign n_12978 = n_12976 & n_12977;
assign n_12979 = n_12978 ^ x113;
assign n_12980 = n_12979 ^ x114;
assign n_12981 = n_12725 ^ n_12979;
assign n_12982 = n_12980 & n_12981;
assign n_12983 = n_12982 ^ x114;
assign n_12984 = n_12983 ^ x115;
assign n_12985 = n_12983 ^ n_12681;
assign n_12986 = n_12773 & n_12983;
assign n_12987 = n_12984 & n_12985;
assign n_12988 = ~n_12782 & ~n_12986;
assign n_12989 = n_12987 ^ x115;
assign n_12990 = x117 ^ n_12988;
assign n_12991 = n_12726 ^ n_12988;
assign n_12992 = n_12989 ^ x116;
assign n_12993 = ~n_12990 & ~n_12991;
assign n_12994 = n_12993 ^ x117;
assign n_12995 = n_12994 ^ x118;
assign n_12996 = n_12727 ^ n_12994;
assign n_12997 = n_12995 & n_12996;
assign n_12998 = n_12997 ^ x118;
assign n_12999 = n_12998 ^ x119;
assign n_13000 = n_12728 ^ n_12998;
assign n_13001 = n_12999 & n_13000;
assign n_13002 = n_13001 ^ x119;
assign n_13003 = n_13002 ^ x120;
assign n_13004 = n_12729 ^ n_13002;
assign n_13005 = n_13003 & n_13004;
assign n_13006 = n_13005 ^ x120;
assign n_13007 = n_13006 ^ x121;
assign n_13008 = n_12730 ^ n_13006;
assign n_13009 = n_13007 & n_13008;
assign n_13010 = n_13009 ^ x121;
assign n_13011 = n_13010 ^ x122;
assign n_13012 = n_12731 ^ n_13010;
assign n_13013 = n_13011 & n_13012;
assign n_13014 = n_13013 ^ x122;
assign n_13015 = n_13014 ^ x123;
assign n_13016 = n_12732 ^ n_13014;
assign n_13017 = n_13015 & n_13016;
assign n_13018 = n_13017 ^ x123;
assign n_13019 = n_13018 ^ x124;
assign n_13020 = n_12733 ^ n_13018;
assign n_13021 = n_13019 & n_13020;
assign n_13022 = n_13021 ^ x124;
assign n_13023 = n_13022 ^ x125;
assign n_13024 = n_13022 ^ ~n_12761;
assign n_13025 = n_13023 & n_12738;
assign n_13026 = ~n_13024 ^ n_11102;
assign n_13027 = n_131 & n_13025;
assign n_13028 = n_13023 & n_13026;
assign n_13029 = n_12738 ^ n_13027;
assign n_13030 = n_13028 ^ x125;
assign n_13031 = n_131 & ~n_13030;
assign n_13032 = n_12795 & n_13031;
assign n_13033 = n_12791 & n_13031;
assign n_13034 = x64 & n_13031;
assign n_13035 = n_176 & n_13031;
assign n_13036 = n_12799 & n_13031;
assign n_13037 = n_12805 & n_13031;
assign n_13038 = n_12812 & n_13031;
assign n_13039 = ~n_12814 & n_13031;
assign n_13040 = n_12818 & n_13031;
assign n_13041 = n_12822 & n_13031;
assign n_13042 = n_12826 & n_13031;
assign n_13043 = n_12830 & n_13031;
assign n_13044 = n_12834 & n_13031;
assign n_13045 = n_12838 & n_13031;
assign n_13046 = n_12842 & n_13031;
assign n_13047 = n_12846 & n_13031;
assign n_13048 = n_12850 & n_13031;
assign n_13049 = n_12854 & n_13031;
assign n_13050 = n_12858 & n_13031;
assign n_13051 = n_12862 & n_13031;
assign n_13052 = n_12995 & n_13031;
assign n_13053 = ~n_12990 & n_13031;
assign n_13054 = n_12976 & n_13031;
assign n_13055 = n_12972 & n_13031;
assign n_13056 = n_12933 & n_13031;
assign n_13057 = n_12866 & n_13031;
assign n_13058 = n_12870 & n_13031;
assign n_13059 = n_12874 & n_13031;
assign n_13060 = n_12878 & n_13031;
assign n_13061 = n_12882 & n_13031;
assign n_13062 = n_12886 & n_13031;
assign n_13063 = n_12890 & n_13031;
assign n_13064 = n_12894 & n_13031;
assign n_13065 = n_12899 & n_13031;
assign n_13066 = n_12903 & n_13031;
assign n_13067 = n_12906 & n_13031;
assign n_13068 = n_12910 & n_13031;
assign n_13069 = n_12914 & n_13031;
assign n_13070 = n_12918 & n_13031;
assign n_13071 = n_12922 & n_13031;
assign n_13072 = ~n_12928 & n_13031;
assign n_13073 = ~n_12939 & n_13031;
assign n_13074 = n_12944 & n_13031;
assign n_13075 = n_12948 & n_13031;
assign n_13076 = n_12952 & n_13031;
assign n_13077 = n_12956 & n_13031;
assign n_13078 = n_12960 & n_13031;
assign n_13079 = n_12964 & n_13031;
assign n_13080 = n_12968 & n_13031;
assign n_13081 = n_12980 & n_13031;
assign n_13082 = n_12984 & n_13031;
assign n_13083 = n_12999 & n_13031;
assign n_13084 = n_13003 & n_13031;
assign n_13085 = n_13007 & n_13031;
assign n_13086 = n_13011 & n_13031;
assign n_13087 = n_13015 & n_13031;
assign n_13088 = n_13019 & n_13031;
assign y2 = n_13031;
assign n_13089 = n_291 & ~n_13031;
assign n_13090 = ~n_12787 & n_13031;
assign n_13091 = n_12941 & n_13031;
assign n_13092 = n_12930 & n_13031;
assign n_13093 = n_12992 & n_13031;
assign n_13094 = n_13032 ^ n_12689;
assign n_13095 = n_13033 ^ n_12679;
assign n_13096 = n_13034 & n_290;
assign n_13097 = n_13035 ^ n_12608;
assign n_13098 = n_13036 ^ n_12690;
assign n_13099 = n_13037 ^ n_12688;
assign n_13100 = n_13038 ^ n_12691;
assign n_13101 = n_13039 ^ n_12692;
assign n_13102 = n_13040 ^ n_12693;
assign n_13103 = n_13041 ^ n_12694;
assign n_13104 = n_13042 ^ n_12695;
assign n_13105 = n_13043 ^ n_12735;
assign n_13106 = n_13044 ^ n_12696;
assign n_13107 = n_13045 ^ n_12697;
assign n_13108 = n_13046 ^ n_12698;
assign n_13109 = n_13047 ^ n_12699;
assign n_13110 = n_13048 ^ n_12700;
assign n_13111 = n_13049 ^ n_12701;
assign n_13112 = n_13050 ^ n_12702;
assign n_13113 = n_13051 ^ n_12703;
assign n_13114 = n_13052 ^ n_12727;
assign n_13115 = n_13053 ^ n_12726;
assign n_13116 = n_13054 ^ n_12724;
assign n_13117 = n_13055 ^ n_12723;
assign n_13118 = n_13056 ^ n_12683;
assign n_13119 = n_13057 ^ n_12704;
assign n_13120 = n_13058 ^ n_12705;
assign n_13121 = n_13059 ^ n_12706;
assign n_13122 = n_13060 ^ n_12707;
assign n_13123 = n_13061 ^ n_12708;
assign n_13124 = n_13062 ^ n_12736;
assign n_13125 = n_13063 ^ n_12709;
assign n_13126 = n_13064 ^ n_12710;
assign n_13127 = n_13065 ^ n_12687;
assign n_13128 = n_13066 ^ n_12686;
assign n_13129 = n_13067 ^ n_12711;
assign n_13130 = n_13068 ^ n_12712;
assign n_13131 = n_13069 ^ n_12737;
assign n_13132 = n_13070 ^ n_12713;
assign n_13133 = n_13071 ^ n_12685;
assign n_13134 = n_13072 ^ n_12714;
assign n_13135 = n_13073 ^ n_12715;
assign n_13136 = n_13074 ^ n_12716;
assign n_13137 = n_13075 ^ n_12717;
assign n_13138 = n_13076 ^ n_12718;
assign n_13139 = n_13077 ^ n_12719;
assign n_13140 = n_13078 ^ n_12720;
assign n_13141 = n_13079 ^ n_12721;
assign n_13142 = n_13080 ^ n_12722;
assign n_13143 = n_13081 ^ n_12725;
assign n_13144 = n_13082 ^ n_12681;
assign n_13145 = n_13083 ^ n_12728;
assign n_13146 = n_13084 ^ n_12729;
assign n_13147 = n_13085 ^ n_12730;
assign n_13148 = n_13086 ^ n_12731;
assign n_13149 = n_13087 ^ n_12732;
assign n_13150 = n_13088 ^ n_12733;
assign n_13151 = ~n_329 & ~n_13089;
assign n_13152 = n_12740 ^ n_13090;
assign n_13153 = n_12682 ^ n_13091;
assign n_13154 = n_12684 ^ n_13092;
assign n_13155 = n_12680 ^ n_13093;
assign n_13156 = ~x69 ^ n_13094;
assign n_13157 = n_13094 ^ x69;
assign n_13158 = n_13095 ^ x68;
assign n_13159 = x68 & n_13095;
assign n_13160 = n_13097 ^ x3;
assign n_13161 = ~x119 ^ n_13114;
assign n_13162 = n_13114 ^ x119;
assign n_13163 = n_13115 ^ x118;
assign n_13164 = x118 & ~n_13115;
assign n_13165 = ~x114 ^ n_13116;
assign n_13166 = n_13116 ^ x114;
assign n_13167 = n_13117 ^ x113;
assign n_13168 = x113 & ~n_13117;
assign n_13169 = n_13118 ^ x103;
assign n_13170 = ~n_13096 & n_13151;
assign n_13171 = n_13153 ^ x104;
assign n_13172 = n_13158 ^ n_13159;
assign n_13173 = n_13159 ^ n_13094;
assign n_13174 = n_13163 ^ n_13164;
assign n_13175 = n_13164 ^ n_13114;
assign n_13176 = n_13167 ^ n_13168;
assign n_13177 = n_13168 ^ n_13116;
assign n_13178 = x66 ^ n_13170;
assign n_13179 = n_13160 ^ n_13170;
assign n_13180 = n_13156 & n_13172;
assign n_13181 = ~n_13157 & n_13173;
assign n_13182 = n_13161 & ~n_13174;
assign n_13183 = ~n_13162 & n_13175;
assign n_13184 = n_13165 & ~n_13176;
assign n_13185 = ~n_13166 & n_13177;
assign n_13186 = ~n_13178 & ~n_13179;
assign n_13187 = n_13181 ^ x69;
assign n_13188 = n_13183 ^ x119;
assign n_13189 = n_13185 ^ x114;
assign n_13190 = n_13186 ^ x66;
assign n_13191 = n_13190 ^ x67;
assign n_13192 = n_13152 ^ n_13190;
assign n_13193 = n_13191 & ~n_13192;
assign n_13194 = n_13193 ^ x67;
assign n_13195 = n_13194 ^ x68;
assign n_13196 = n_13194 ^ n_13095;
assign n_13197 = n_13180 & n_13194;
assign n_13198 = n_13195 & ~n_13196;
assign n_13199 = ~n_13187 & ~n_13197;
assign n_13200 = n_13198 ^ x68;
assign n_13201 = x70 ^ n_13199;
assign n_13202 = n_13098 ^ n_13199;
assign n_13203 = n_13200 ^ x69;
assign n_13204 = ~n_13201 & ~n_13202;
assign n_13205 = n_13204 ^ x70;
assign n_13206 = n_13205 ^ x71;
assign n_13207 = n_13099 ^ n_13205;
assign n_13208 = n_13206 & n_13207;
assign n_13209 = n_13208 ^ x71;
assign n_13210 = n_13209 ^ x72;
assign n_13211 = n_13100 ^ n_13209;
assign n_13212 = n_13210 & n_13211;
assign n_13213 = n_13212 ^ x72;
assign n_13214 = n_13213 ^ x73;
assign n_13215 = n_13101 ^ n_13213;
assign n_13216 = n_13214 & n_13215;
assign n_13217 = n_13216 ^ x73;
assign n_13218 = n_13217 ^ x74;
assign n_13219 = n_13102 ^ n_13217;
assign n_13220 = n_13218 & n_13219;
assign n_13221 = n_13220 ^ x74;
assign n_13222 = n_13221 ^ x75;
assign n_13223 = n_13103 ^ n_13221;
assign n_13224 = n_13222 & n_13223;
assign n_13225 = n_13224 ^ x75;
assign n_13226 = n_13225 ^ x76;
assign n_13227 = n_13104 ^ n_13225;
assign n_13228 = n_13226 & n_13227;
assign n_13229 = n_13228 ^ x76;
assign n_13230 = n_13229 ^ x77;
assign n_13231 = n_13105 ^ n_13229;
assign n_13232 = n_13230 & n_13231;
assign n_13233 = n_13232 ^ x77;
assign n_13234 = n_13233 ^ x78;
assign n_13235 = n_13106 ^ n_13233;
assign n_13236 = n_13234 & n_13235;
assign n_13237 = n_13236 ^ x78;
assign n_13238 = n_13237 ^ x79;
assign n_13239 = n_13107 ^ n_13237;
assign n_13240 = n_13238 & n_13239;
assign n_13241 = n_13240 ^ x79;
assign n_13242 = n_13241 ^ x80;
assign n_13243 = n_13108 ^ n_13241;
assign n_13244 = n_13242 & n_13243;
assign n_13245 = n_13244 ^ x80;
assign n_13246 = n_13245 ^ x81;
assign n_13247 = n_13109 ^ n_13245;
assign n_13248 = n_13246 & n_13247;
assign n_13249 = n_13248 ^ x81;
assign n_13250 = n_13249 ^ x82;
assign n_13251 = n_13110 ^ n_13249;
assign n_13252 = n_13250 & n_13251;
assign n_13253 = n_13252 ^ x82;
assign n_13254 = n_13253 ^ x83;
assign n_13255 = n_13111 ^ n_13253;
assign n_13256 = n_13254 & n_13255;
assign n_13257 = n_13256 ^ x83;
assign n_13258 = n_13257 ^ x84;
assign n_13259 = n_13112 ^ n_13257;
assign n_13260 = n_13258 & n_13259;
assign n_13261 = n_13260 ^ x84;
assign n_13262 = n_13261 ^ x85;
assign n_13263 = n_13113 ^ n_13261;
assign n_13264 = n_13262 & n_13263;
assign n_13265 = n_13264 ^ x85;
assign n_13266 = n_13265 ^ x86;
assign n_13267 = n_13119 ^ n_13265;
assign n_13268 = n_13266 & n_13267;
assign n_13269 = n_13268 ^ x86;
assign n_13270 = n_13269 ^ x87;
assign n_13271 = n_13120 ^ n_13269;
assign n_13272 = n_13270 & n_13271;
assign n_13273 = n_13272 ^ x87;
assign n_13274 = n_13273 ^ x88;
assign n_13275 = n_13121 ^ n_13273;
assign n_13276 = n_13274 & n_13275;
assign n_13277 = n_13276 ^ x88;
assign n_13278 = n_13277 ^ x89;
assign n_13279 = n_13122 ^ n_13277;
assign n_13280 = n_13278 & n_13279;
assign n_13281 = n_13280 ^ x89;
assign n_13282 = n_13281 ^ x90;
assign n_13283 = n_13123 ^ n_13281;
assign n_13284 = n_13282 & n_13283;
assign n_13285 = n_13284 ^ x90;
assign n_13286 = n_13285 ^ x91;
assign n_13287 = n_13124 ^ n_13285;
assign n_13288 = n_13286 & n_13287;
assign n_13289 = n_13288 ^ x91;
assign n_13290 = n_13289 ^ x92;
assign n_13291 = n_13125 ^ n_13289;
assign n_13292 = n_13290 & n_13291;
assign n_13293 = n_13292 ^ x92;
assign n_13294 = n_13293 ^ x93;
assign n_13295 = n_13126 ^ n_13293;
assign n_13296 = n_13294 & n_13295;
assign n_13297 = n_13296 ^ x93;
assign n_13298 = n_13297 ^ x94;
assign n_13299 = n_13127 ^ n_13297;
assign n_13300 = n_13298 & n_13299;
assign n_13301 = n_13300 ^ x94;
assign n_13302 = n_13301 ^ x95;
assign n_13303 = n_13128 ^ n_13301;
assign n_13304 = n_13302 & ~n_13303;
assign n_13305 = n_13304 ^ x95;
assign n_13306 = n_13305 ^ x96;
assign n_13307 = n_13129 ^ n_13305;
assign n_13308 = n_13306 & n_13307;
assign n_13309 = n_13308 ^ x96;
assign n_13310 = n_13309 ^ x97;
assign n_13311 = n_13130 ^ n_13309;
assign n_13312 = n_13310 & n_13311;
assign n_13313 = n_13312 ^ x97;
assign n_13314 = n_13313 ^ x98;
assign n_13315 = n_13131 ^ n_13313;
assign n_13316 = n_13314 & n_13315;
assign n_13317 = n_13316 ^ x98;
assign n_13318 = n_13317 ^ x99;
assign n_13319 = n_13132 ^ n_13317;
assign n_13320 = n_13318 & n_13319;
assign n_13321 = n_13320 ^ x99;
assign n_13322 = n_13321 ^ x100;
assign n_13323 = n_13133 ^ n_13321;
assign n_13324 = n_13322 & n_13323;
assign n_13325 = n_13324 ^ x100;
assign n_13326 = n_13325 ^ x101;
assign n_13327 = n_13154 ^ n_13325;
assign n_13328 = n_13326 & n_13327;
assign n_13329 = n_13328 ^ x101;
assign n_13330 = n_13329 ^ x102;
assign n_13331 = n_13134 ^ n_13329;
assign n_13332 = n_13330 & n_13331;
assign n_13333 = n_13332 ^ x102;
assign n_13334 = n_13333 ^ n_13118;
assign n_13335 = n_13333 ^ x103;
assign n_13336 = ~n_13169 & n_13334;
assign n_13337 = n_13336 ^ x103;
assign n_13338 = n_13337 ^ n_13153;
assign n_13339 = n_13337 ^ x104;
assign n_13340 = ~n_13171 & n_13338;
assign n_13341 = n_13340 ^ x104;
assign n_13342 = n_13341 ^ x105;
assign n_13343 = n_13135 ^ n_13341;
assign n_13344 = n_13342 & n_13343;
assign n_13345 = n_13344 ^ x105;
assign n_13346 = n_13345 ^ x106;
assign n_13347 = n_13136 ^ n_13345;
assign n_13348 = n_13346 & n_13347;
assign n_13349 = n_13348 ^ x106;
assign n_13350 = n_13349 ^ x107;
assign n_13351 = n_13137 ^ n_13349;
assign n_13352 = n_13350 & n_13351;
assign n_13353 = n_13352 ^ x107;
assign n_13354 = n_13353 ^ x108;
assign n_13355 = n_13138 ^ n_13353;
assign n_13356 = n_13354 & n_13355;
assign n_13357 = n_13356 ^ x108;
assign n_13358 = n_13357 ^ x109;
assign n_13359 = n_13139 ^ n_13357;
assign n_13360 = n_13358 & n_13359;
assign n_13361 = n_13360 ^ x109;
assign n_13362 = n_13361 ^ x110;
assign n_13363 = n_13140 ^ n_13361;
assign n_13364 = n_13362 & n_13363;
assign n_13365 = n_13364 ^ x110;
assign n_13366 = n_13365 ^ x111;
assign n_13367 = n_13141 ^ n_13365;
assign n_13368 = n_13366 & n_13367;
assign n_13369 = n_13368 ^ x111;
assign n_13370 = n_13369 ^ x112;
assign n_13371 = n_13142 ^ n_13369;
assign n_13372 = n_13370 & n_13371;
assign n_13373 = n_13372 ^ x112;
assign n_13374 = n_13373 ^ x113;
assign n_13375 = n_13373 ^ n_13117;
assign n_13376 = n_13184 & n_13373;
assign n_13377 = n_13374 & n_13375;
assign n_13378 = ~n_13189 & ~n_13376;
assign n_13379 = n_13377 ^ x113;
assign n_13380 = x115 ^ n_13378;
assign n_13381 = n_13143 ^ n_13378;
assign n_13382 = n_13379 ^ x114;
assign n_13383 = ~n_13380 & ~n_13381;
assign n_13384 = n_13383 ^ x115;
assign n_13385 = n_13384 ^ x116;
assign n_13386 = n_13144 ^ n_13384;
assign n_13387 = n_13385 & n_13386;
assign n_13388 = n_13387 ^ x116;
assign n_13389 = n_13388 ^ x117;
assign n_13390 = n_13155 ^ n_13388;
assign n_13391 = n_13389 & n_13390;
assign n_13392 = n_13391 ^ x117;
assign n_13393 = n_13392 ^ x118;
assign n_13394 = n_13392 ^ n_13115;
assign n_13395 = n_13182 & n_13392;
assign n_13396 = n_13393 & n_13394;
assign n_13397 = ~n_13188 & ~n_13395;
assign n_13398 = n_13396 ^ x118;
assign n_13399 = x120 ^ n_13397;
assign n_13400 = n_13145 ^ n_13397;
assign n_13401 = n_13398 ^ x119;
assign n_13402 = ~n_13399 & ~n_13400;
assign n_13403 = n_13402 ^ x120;
assign n_13404 = n_13403 ^ x121;
assign n_13405 = n_13146 ^ n_13403;
assign n_13406 = n_13404 & n_13405;
assign n_13407 = n_13406 ^ x121;
assign n_13408 = n_13407 ^ x122;
assign n_13409 = n_13147 ^ n_13407;
assign n_13410 = n_13408 & n_13409;
assign n_13411 = n_13410 ^ x122;
assign n_13412 = n_13411 ^ x123;
assign n_13413 = n_13148 ^ n_13411;
assign n_13414 = n_13412 & n_13413;
assign n_13415 = n_13414 ^ x123;
assign n_13416 = n_13415 ^ x124;
assign n_13417 = n_13149 ^ n_13415;
assign n_13418 = n_13416 & n_13417;
assign n_13419 = n_13418 ^ x124;
assign n_13420 = n_13419 ^ x125;
assign n_13421 = n_13150 ^ n_13419;
assign n_13422 = n_13420 & n_13421;
assign n_13423 = n_13422 ^ x125;
assign n_13424 = n_13423 ^ x126;
assign n_13425 = n_13029 ^ n_13423;
assign n_13426 = ~x127 & ~n_13424;
assign n_13427 = n_13424 & n_13425;
assign n_13428 = n_13029 & n_13426;
assign n_13429 = n_13426 ^ x127;
assign n_13430 = n_13427 ^ x126;
assign n_13431 = ~x127 & ~n_13430;
assign n_13432 = n_13266 & n_13431;
assign n_13433 = n_13262 & n_13431;
assign n_13434 = n_13226 & n_13431;
assign n_13435 = n_13222 & n_13431;
assign n_13436 = n_13206 & n_13431;
assign n_13437 = ~n_13201 & n_13431;
assign n_13438 = x64 & n_13431;
assign n_13439 = ~n_340 & ~n_13431;
assign n_13440 = x65 & n_13431;
assign n_13441 = ~n_13178 & n_13431;
assign n_13442 = n_13191 & n_13431;
assign n_13443 = n_13195 & n_13431;
assign n_13444 = n_13210 & n_13431;
assign n_13445 = n_13214 & n_13431;
assign n_13446 = n_13218 & n_13431;
assign n_13447 = n_13230 & n_13431;
assign n_13448 = n_13234 & n_13431;
assign n_13449 = n_13238 & n_13431;
assign n_13450 = n_13242 & n_13431;
assign n_13451 = n_13246 & n_13431;
assign n_13452 = n_13250 & n_13431;
assign n_13453 = n_13254 & n_13431;
assign n_13454 = n_13258 & n_13431;
assign n_13455 = n_13270 & n_13431;
assign n_13456 = n_13274 & n_13431;
assign n_13457 = n_13278 & n_13431;
assign n_13458 = n_13282 & n_13431;
assign n_13459 = n_13286 & n_13431;
assign n_13460 = n_13290 & n_13431;
assign n_13461 = n_13294 & n_13431;
assign n_13462 = n_13298 & n_13431;
assign n_13463 = n_13302 & n_13431;
assign n_13464 = n_13306 & n_13431;
assign n_13465 = n_13310 & n_13431;
assign n_13466 = n_13314 & n_13431;
assign n_13467 = n_13318 & n_13431;
assign n_13468 = n_13322 & n_13431;
assign n_13469 = n_13326 & n_13431;
assign n_13470 = n_13330 & n_13431;
assign n_13471 = n_13335 & n_13431;
assign n_13472 = n_13339 & n_13431;
assign n_13473 = n_13342 & n_13431;
assign n_13474 = n_13346 & n_13431;
assign n_13475 = n_13350 & n_13431;
assign n_13476 = n_13354 & n_13431;
assign n_13477 = n_13358 & n_13431;
assign n_13478 = n_13362 & n_13431;
assign n_13479 = n_13366 & n_13431;
assign n_13480 = n_13370 & n_13431;
assign n_13481 = n_13374 & n_13431;
assign n_13482 = ~n_13380 & n_13431;
assign n_13483 = n_13385 & n_13431;
assign n_13484 = n_13389 & n_13431;
assign n_13485 = n_13393 & n_13431;
assign n_13486 = ~n_13399 & n_13431;
assign n_13487 = n_13404 & n_13431;
assign n_13488 = n_13408 & n_13431;
assign n_13489 = n_13412 & n_13431;
assign n_13490 = n_13416 & n_13431;
assign n_13491 = n_13420 & n_13431;
assign y1 = n_13431;
assign n_13492 = n_13203 & n_13431;
assign n_13493 = n_13382 & n_13431;
assign n_13494 = n_13401 & n_13431;
assign n_13495 = n_13432 ^ n_13119;
assign n_13496 = n_13433 ^ n_13113;
assign n_13497 = n_13434 ^ n_13104;
assign n_13498 = n_13435 ^ n_13103;
assign n_13499 = n_13436 ^ n_13099;
assign n_13500 = n_13437 ^ n_13098;
assign n_13501 = ~x1 & n_13438;
assign n_13502 = n_13438 & n_242;
assign n_13503 = n_13439 ^ x65;
assign n_13504 = n_13441 ^ n_13160;
assign n_13505 = n_13442 ^ n_13152;
assign n_13506 = n_13443 ^ n_13095;
assign n_13507 = n_13444 ^ n_13100;
assign n_13508 = n_13445 ^ n_13101;
assign n_13509 = n_13446 ^ n_13102;
assign n_13510 = n_13447 ^ n_13105;
assign n_13511 = n_13448 ^ n_13106;
assign n_13512 = n_13449 ^ n_13107;
assign n_13513 = n_13450 ^ n_13108;
assign n_13514 = n_13451 ^ n_13109;
assign n_13515 = n_13452 ^ n_13110;
assign n_13516 = n_13453 ^ n_13111;
assign n_13517 = n_13454 ^ n_13112;
assign n_13518 = n_13455 ^ n_13120;
assign n_13519 = n_13456 ^ n_13121;
assign n_13520 = n_13457 ^ n_13122;
assign n_13521 = n_13458 ^ n_13123;
assign n_13522 = n_13459 ^ n_13124;
assign n_13523 = n_13460 ^ n_13125;
assign n_13524 = n_13461 ^ n_13126;
assign n_13525 = n_13462 ^ n_13127;
assign n_13526 = n_13463 ^ n_13128;
assign n_13527 = n_13464 ^ n_13129;
assign n_13528 = n_13465 ^ n_13130;
assign n_13529 = n_13466 ^ n_13131;
assign n_13530 = n_13467 ^ n_13132;
assign n_13531 = n_13468 ^ n_13133;
assign n_13532 = n_13469 ^ n_13154;
assign n_13533 = n_13470 ^ n_13134;
assign n_13534 = n_13471 ^ n_13118;
assign n_13535 = n_13472 ^ n_13153;
assign n_13536 = n_13473 ^ n_13135;
assign n_13537 = n_13474 ^ n_13136;
assign n_13538 = n_13475 ^ n_13137;
assign n_13539 = n_13476 ^ n_13138;
assign n_13540 = n_13477 ^ n_13139;
assign n_13541 = n_13478 ^ n_13140;
assign n_13542 = n_13479 ^ n_13141;
assign n_13543 = n_13480 ^ n_13142;
assign n_13544 = n_13481 ^ n_13117;
assign n_13545 = n_13482 ^ n_13143;
assign n_13546 = n_13483 ^ n_13144;
assign n_13547 = n_13484 ^ n_13155;
assign n_13548 = n_13485 ^ n_13115;
assign n_13549 = n_13486 ^ n_13145;
assign n_13550 = n_13487 ^ n_13146;
assign n_13551 = n_13488 ^ n_13147;
assign n_13552 = n_13489 ^ n_13148;
assign n_13553 = n_13490 ^ n_13149;
assign n_13554 = n_13491 ^ n_13150;
assign n_13555 = n_13094 ^ n_13492;
assign n_13556 = n_13116 ^ n_13493;
assign n_13557 = n_13114 ^ n_13494;
assign n_13558 = ~x87 ^ n_13495;
assign n_13559 = n_13495 ^ x87;
assign n_13560 = n_13496 ^ x86;
assign n_13561 = x86 & ~n_13496;
assign n_13562 = ~x77 ^ n_13497;
assign n_13563 = n_13497 ^ x77;
assign n_13564 = n_13498 ^ x76;
assign n_13565 = x76 & ~n_13498;
assign n_13566 = n_13499 ^ x72;
assign n_13567 = n_13500 ^ x71;
assign n_13568 = n_13501 ^ n_13034;
assign n_13569 = ~n_347 & n_13503;
assign n_13570 = n_13560 ^ n_13561;
assign n_13571 = n_13561 ^ n_13495;
assign n_13572 = n_13564 ^ n_13565;
assign n_13573 = n_13565 ^ n_13497;
assign n_13574 = n_13440 ^ n_13568;
assign n_13575 = x65 ^ n_13569;
assign n_13576 = n_13558 & ~n_13570;
assign n_13577 = ~n_13559 & n_13571;
assign n_13578 = n_13562 & ~n_13572;
assign n_13579 = ~n_13563 & n_13573;
assign n_13580 = n_13574 ^ x2;
assign n_13581 = n_13575 ^ x65;
assign n_13582 = n_13577 ^ x87;
assign n_13583 = n_13579 ^ x77;
assign n_13584 = n_13581 ^ x65;
assign n_13585 = ~n_13584 & ~n_13502;
assign n_13586 = x66 ^ n_13585;
assign n_13587 = n_13580 ^ n_13585;
assign n_13588 = ~n_13586 & ~n_13587;
assign n_13589 = n_13588 ^ x66;
assign n_13590 = n_13589 ^ x67;
assign n_13591 = n_13504 ^ n_13589;
assign n_13592 = n_13590 & n_13591;
assign n_13593 = n_13592 ^ x67;
assign n_13594 = n_13593 ^ x68;
assign n_13595 = n_13505 ^ n_13593;
assign n_13596 = n_13594 & ~n_13595;
assign n_13597 = n_13596 ^ x68;
assign n_13598 = n_13597 ^ x69;
assign n_13599 = n_13506 ^ n_13597;
assign n_13600 = n_13598 & ~n_13599;
assign n_13601 = n_13600 ^ x69;
assign n_13602 = n_13601 ^ x70;
assign n_13603 = n_13555 ^ n_13601;
assign n_13604 = n_13602 & n_13603;
assign n_13605 = n_13604 ^ x70;
assign n_13606 = n_13605 ^ n_13500;
assign n_13607 = n_13605 ^ x71;
assign n_13608 = ~n_13567 & n_13606;
assign n_13609 = n_13608 ^ x71;
assign n_13610 = n_13609 ^ n_13499;
assign n_13611 = n_13609 ^ x72;
assign n_13612 = ~n_13566 & n_13610;
assign n_13613 = n_13612 ^ x72;
assign n_13614 = n_13613 ^ x73;
assign n_13615 = n_13507 ^ n_13613;
assign n_13616 = n_13614 & n_13615;
assign n_13617 = n_13616 ^ x73;
assign n_13618 = n_13617 ^ x74;
assign n_13619 = n_13508 ^ n_13617;
assign n_13620 = n_13618 & n_13619;
assign n_13621 = n_13620 ^ x74;
assign n_13622 = n_13621 ^ x75;
assign n_13623 = n_13509 ^ n_13621;
assign n_13624 = n_13622 & n_13623;
assign n_13625 = n_13624 ^ x75;
assign n_13626 = n_13625 ^ x76;
assign n_13627 = n_13625 ^ n_13498;
assign n_13628 = n_13578 & n_13625;
assign n_13629 = n_13626 & n_13627;
assign n_13630 = ~n_13583 & ~n_13628;
assign n_13631 = n_13629 ^ x76;
assign n_13632 = x78 ^ n_13630;
assign n_13633 = n_13510 ^ n_13630;
assign n_13634 = n_13631 ^ x77;
assign n_13635 = ~n_13632 & ~n_13633;
assign n_13636 = n_13635 ^ x78;
assign n_13637 = n_13636 ^ x79;
assign n_13638 = n_13511 ^ n_13636;
assign n_13639 = n_13637 & n_13638;
assign n_13640 = n_13639 ^ x79;
assign n_13641 = n_13640 ^ x80;
assign n_13642 = n_13512 ^ n_13640;
assign n_13643 = n_13641 & n_13642;
assign n_13644 = n_13643 ^ x80;
assign n_13645 = n_13644 ^ x81;
assign n_13646 = n_13513 ^ n_13644;
assign n_13647 = n_13645 & n_13646;
assign n_13648 = n_13647 ^ x81;
assign n_13649 = n_13648 ^ x82;
assign n_13650 = n_13514 ^ n_13648;
assign n_13651 = n_13649 & n_13650;
assign n_13652 = n_13651 ^ x82;
assign n_13653 = n_13652 ^ x83;
assign n_13654 = n_13515 ^ n_13652;
assign n_13655 = n_13653 & n_13654;
assign n_13656 = n_13655 ^ x83;
assign n_13657 = n_13656 ^ x84;
assign n_13658 = n_13516 ^ n_13656;
assign n_13659 = n_13657 & n_13658;
assign n_13660 = n_13659 ^ x84;
assign n_13661 = n_13660 ^ x85;
assign n_13662 = n_13517 ^ n_13660;
assign n_13663 = n_13661 & n_13662;
assign n_13664 = n_13663 ^ x85;
assign n_13665 = n_13664 ^ x86;
assign n_13666 = n_13664 ^ n_13496;
assign n_13667 = n_13576 & n_13664;
assign n_13668 = n_13665 & n_13666;
assign n_13669 = ~n_13582 & ~n_13667;
assign n_13670 = n_13668 ^ x86;
assign n_13671 = x88 ^ n_13669;
assign n_13672 = n_13518 ^ n_13669;
assign n_13673 = n_13670 ^ x87;
assign n_13674 = ~n_13671 & ~n_13672;
assign n_13675 = n_13674 ^ x88;
assign n_13676 = n_13675 ^ x89;
assign n_13677 = n_13519 ^ n_13675;
assign n_13678 = n_13676 & n_13677;
assign n_13679 = n_13678 ^ x89;
assign n_13680 = n_13679 ^ x90;
assign n_13681 = n_13520 ^ n_13679;
assign n_13682 = n_13680 & n_13681;
assign n_13683 = n_13682 ^ x90;
assign n_13684 = n_13683 ^ x91;
assign n_13685 = n_13521 ^ n_13683;
assign n_13686 = n_13684 & n_13685;
assign n_13687 = n_13686 ^ x91;
assign n_13688 = n_13687 ^ x92;
assign n_13689 = n_13522 ^ n_13687;
assign n_13690 = n_13688 & n_13689;
assign n_13691 = n_13690 ^ x92;
assign n_13692 = n_13691 ^ x93;
assign n_13693 = n_13523 ^ n_13691;
assign n_13694 = n_13692 & n_13693;
assign n_13695 = n_13694 ^ x93;
assign n_13696 = n_13695 ^ x94;
assign n_13697 = n_13524 ^ n_13695;
assign n_13698 = n_13696 & n_13697;
assign n_13699 = n_13698 ^ x94;
assign n_13700 = n_13699 ^ x95;
assign n_13701 = n_13525 ^ n_13699;
assign n_13702 = n_13700 & n_13701;
assign n_13703 = n_13702 ^ x95;
assign n_13704 = n_13703 ^ x96;
assign n_13705 = n_13526 ^ n_13703;
assign n_13706 = n_13704 & ~n_13705;
assign n_13707 = n_13706 ^ x96;
assign n_13708 = n_13707 ^ x97;
assign n_13709 = n_13527 ^ n_13707;
assign n_13710 = n_13708 & n_13709;
assign n_13711 = n_13710 ^ x97;
assign n_13712 = n_13711 ^ x98;
assign n_13713 = n_13528 ^ n_13711;
assign n_13714 = n_13712 & n_13713;
assign n_13715 = n_13714 ^ x98;
assign n_13716 = n_13715 ^ x99;
assign n_13717 = n_13529 ^ n_13715;
assign n_13718 = n_13716 & n_13717;
assign n_13719 = n_13718 ^ x99;
assign n_13720 = n_13719 ^ x100;
assign n_13721 = n_13530 ^ n_13719;
assign n_13722 = n_13720 & n_13721;
assign n_13723 = n_13722 ^ x100;
assign n_13724 = n_13723 ^ x101;
assign n_13725 = n_13531 ^ n_13723;
assign n_13726 = n_13724 & n_13725;
assign n_13727 = n_13726 ^ x101;
assign n_13728 = n_13727 ^ x102;
assign n_13729 = n_13532 ^ n_13727;
assign n_13730 = n_13728 & n_13729;
assign n_13731 = n_13730 ^ x102;
assign n_13732 = n_13731 ^ x103;
assign n_13733 = n_13533 ^ n_13731;
assign n_13734 = n_13732 & n_13733;
assign n_13735 = n_13734 ^ x103;
assign n_13736 = n_13735 ^ x104;
assign n_13737 = n_13534 ^ n_13735;
assign n_13738 = n_13736 & n_13737;
assign n_13739 = n_13738 ^ x104;
assign n_13740 = n_13739 ^ x105;
assign n_13741 = n_13535 ^ n_13739;
assign n_13742 = n_13740 & n_13741;
assign n_13743 = n_13742 ^ x105;
assign n_13744 = n_13743 ^ x106;
assign n_13745 = n_13536 ^ n_13743;
assign n_13746 = n_13744 & n_13745;
assign n_13747 = n_13746 ^ x106;
assign n_13748 = n_13747 ^ x107;
assign n_13749 = n_13537 ^ n_13747;
assign n_13750 = n_13748 & n_13749;
assign n_13751 = n_13750 ^ x107;
assign n_13752 = n_13751 ^ x108;
assign n_13753 = n_13538 ^ n_13751;
assign n_13754 = n_13752 & n_13753;
assign n_13755 = n_13754 ^ x108;
assign n_13756 = n_13755 ^ x109;
assign n_13757 = n_13539 ^ n_13755;
assign n_13758 = n_13756 & n_13757;
assign n_13759 = n_13758 ^ x109;
assign n_13760 = n_13759 ^ x110;
assign n_13761 = n_13540 ^ n_13759;
assign n_13762 = n_13760 & n_13761;
assign n_13763 = n_13762 ^ x110;
assign n_13764 = n_13763 ^ x111;
assign n_13765 = n_13541 ^ n_13763;
assign n_13766 = n_13764 & n_13765;
assign n_13767 = n_13766 ^ x111;
assign n_13768 = n_13767 ^ x112;
assign n_13769 = n_13542 ^ n_13767;
assign n_13770 = n_13768 & n_13769;
assign n_13771 = n_13770 ^ x112;
assign n_13772 = n_13771 ^ x113;
assign n_13773 = n_13543 ^ n_13771;
assign n_13774 = n_13772 & n_13773;
assign n_13775 = n_13774 ^ x113;
assign n_13776 = n_13775 ^ x114;
assign n_13777 = n_13544 ^ n_13775;
assign n_13778 = n_13776 & n_13777;
assign n_13779 = n_13778 ^ x114;
assign n_13780 = n_13779 ^ x115;
assign n_13781 = n_13556 ^ n_13779;
assign n_13782 = n_13780 & n_13781;
assign n_13783 = n_13782 ^ x115;
assign n_13784 = n_13783 ^ x116;
assign n_13785 = n_13545 ^ n_13783;
assign n_13786 = n_13784 & n_13785;
assign n_13787 = n_13786 ^ x116;
assign n_13788 = n_13787 ^ x117;
assign n_13789 = n_13546 ^ n_13787;
assign n_13790 = n_13788 & n_13789;
assign n_13791 = n_13790 ^ x117;
assign n_13792 = n_13791 ^ x118;
assign n_13793 = n_13547 ^ n_13791;
assign n_13794 = n_13792 & n_13793;
assign n_13795 = n_13794 ^ x118;
assign n_13796 = n_13795 ^ x119;
assign n_13797 = n_13548 ^ n_13795;
assign n_13798 = n_13796 & n_13797;
assign n_13799 = n_13798 ^ x119;
assign n_13800 = n_13799 ^ x120;
assign n_13801 = n_13557 ^ n_13799;
assign n_13802 = n_13800 & n_13801;
assign n_13803 = n_13802 ^ x120;
assign n_13804 = n_13803 ^ x121;
assign n_13805 = n_13549 ^ n_13803;
assign n_13806 = n_13804 & n_13805;
assign n_13807 = n_13806 ^ x121;
assign n_13808 = n_13807 ^ x122;
assign n_13809 = n_13550 ^ n_13807;
assign n_13810 = n_13808 & n_13809;
assign n_13811 = n_13810 ^ x122;
assign n_13812 = n_13811 ^ x123;
assign n_13813 = n_13551 ^ n_13811;
assign n_13814 = n_13812 & n_13813;
assign n_13815 = n_13814 ^ x123;
assign n_13816 = n_13815 ^ x124;
assign n_13817 = n_13552 ^ n_13815;
assign n_13818 = n_13816 & n_13817;
assign n_13819 = n_13818 ^ x124;
assign n_13820 = n_13819 ^ x125;
assign n_13821 = n_13553 ^ n_13819;
assign n_13822 = n_13820 & n_13821;
assign n_13823 = n_13822 ^ x125;
assign n_13824 = n_13823 ^ x126;
assign n_13825 = n_13554 ^ n_13823;
assign n_13826 = n_13824 & n_13825;
assign n_13827 = n_13826 ^ x126;
assign n_13828 = ~n_13827 & n_13429;
assign n_13829 = ~n_11802 & ~n_13827;
assign n_13830 = n_13828 ^ x127;
assign n_13831 = ~n_13428 & ~n_13829;
assign n_13832 = n_13029 & n_13830;
assign n_13833 = x64 & ~n_13831;
assign n_13834 = x65 & ~n_13831;
assign n_13835 = ~n_13586 & ~n_13831;
assign n_13836 = n_13590 & ~n_13831;
assign n_13837 = n_13594 & ~n_13831;
assign n_13838 = n_13598 & ~n_13831;
assign n_13839 = n_13602 & ~n_13831;
assign n_13840 = n_13607 & ~n_13831;
assign n_13841 = n_13611 & ~n_13831;
assign n_13842 = n_13614 & ~n_13831;
assign n_13843 = n_13618 & ~n_13831;
assign n_13844 = n_13622 & ~n_13831;
assign n_13845 = n_13626 & ~n_13831;
assign n_13846 = ~n_13632 & ~n_13831;
assign n_13847 = n_13637 & ~n_13831;
assign n_13848 = n_13641 & ~n_13831;
assign n_13849 = n_13645 & ~n_13831;
assign n_13850 = n_13649 & ~n_13831;
assign n_13851 = n_13653 & ~n_13831;
assign n_13852 = n_13657 & ~n_13831;
assign n_13853 = n_13661 & ~n_13831;
assign n_13854 = n_13665 & ~n_13831;
assign n_13855 = ~n_13671 & ~n_13831;
assign n_13856 = n_13676 & ~n_13831;
assign n_13857 = n_13680 & ~n_13831;
assign n_13858 = n_13684 & ~n_13831;
assign n_13859 = n_13688 & ~n_13831;
assign n_13860 = n_13692 & ~n_13831;
assign n_13861 = n_13696 & ~n_13831;
assign n_13862 = n_13700 & ~n_13831;
assign n_13863 = n_13704 & ~n_13831;
assign n_13864 = n_13708 & ~n_13831;
assign n_13865 = n_13712 & ~n_13831;
assign n_13866 = n_13716 & ~n_13831;
assign n_13867 = n_13720 & ~n_13831;
assign n_13868 = n_13724 & ~n_13831;
assign n_13869 = n_13728 & ~n_13831;
assign n_13870 = n_13732 & ~n_13831;
assign n_13871 = n_13736 & ~n_13831;
assign n_13872 = n_13740 & ~n_13831;
assign n_13873 = n_13744 & ~n_13831;
assign n_13874 = n_13748 & ~n_13831;
assign n_13875 = n_13752 & ~n_13831;
assign n_13876 = n_13756 & ~n_13831;
assign n_13877 = n_13760 & ~n_13831;
assign n_13878 = n_13764 & ~n_13831;
assign n_13879 = n_13768 & ~n_13831;
assign n_13880 = n_13772 & ~n_13831;
assign n_13881 = n_13776 & ~n_13831;
assign n_13882 = n_13780 & ~n_13831;
assign n_13883 = n_13784 & ~n_13831;
assign n_13884 = n_13788 & ~n_13831;
assign n_13885 = n_13792 & ~n_13831;
assign n_13886 = n_13796 & ~n_13831;
assign n_13887 = n_13800 & ~n_13831;
assign n_13888 = n_13804 & ~n_13831;
assign n_13889 = n_13808 & ~n_13831;
assign n_13890 = n_13812 & ~n_13831;
assign n_13891 = n_13816 & ~n_13831;
assign n_13892 = n_13820 & ~n_13831;
assign n_13893 = n_13824 & ~n_13831;
assign y0 = ~n_13831;
assign n_13894 = n_13634 & ~n_13831;
assign n_13895 = n_13673 & ~n_13831;
assign y127 = n_13832;
assign n_13896 = n_13833 ^ x0;
assign n_13897 = n_13835 ^ n_13580;
assign n_13898 = n_13836 ^ n_13504;
assign n_13899 = n_13837 ^ n_13505;
assign n_13900 = n_13838 ^ n_13506;
assign n_13901 = n_13839 ^ n_13555;
assign n_13902 = n_13840 ^ n_13500;
assign n_13903 = n_13841 ^ n_13499;
assign n_13904 = n_13842 ^ n_13507;
assign n_13905 = n_13843 ^ n_13508;
assign n_13906 = n_13844 ^ n_13509;
assign n_13907 = n_13845 ^ n_13498;
assign n_13908 = n_13846 ^ n_13510;
assign n_13909 = n_13847 ^ n_13511;
assign n_13910 = n_13848 ^ n_13512;
assign n_13911 = n_13849 ^ n_13513;
assign n_13912 = n_13850 ^ n_13514;
assign n_13913 = n_13851 ^ n_13515;
assign n_13914 = n_13852 ^ n_13516;
assign n_13915 = n_13853 ^ n_13517;
assign n_13916 = n_13854 ^ n_13496;
assign n_13917 = n_13855 ^ n_13518;
assign n_13918 = n_13856 ^ n_13519;
assign n_13919 = n_13857 ^ n_13520;
assign n_13920 = n_13858 ^ n_13521;
assign n_13921 = n_13859 ^ n_13522;
assign n_13922 = n_13860 ^ n_13523;
assign n_13923 = n_13861 ^ n_13524;
assign n_13924 = n_13862 ^ n_13525;
assign n_13925 = n_13863 ^ n_13526;
assign n_13926 = n_13864 ^ n_13527;
assign n_13927 = n_13865 ^ n_13528;
assign n_13928 = n_13866 ^ n_13529;
assign n_13929 = n_13867 ^ n_13530;
assign n_13930 = n_13868 ^ n_13531;
assign n_13931 = n_13869 ^ n_13532;
assign n_13932 = n_13870 ^ n_13533;
assign n_13933 = n_13871 ^ n_13534;
assign n_13934 = n_13872 ^ n_13535;
assign n_13935 = n_13873 ^ n_13536;
assign n_13936 = n_13874 ^ n_13537;
assign n_13937 = n_13875 ^ n_13538;
assign n_13938 = n_13876 ^ n_13539;
assign n_13939 = n_13877 ^ n_13540;
assign n_13940 = n_13878 ^ n_13541;
assign n_13941 = n_13879 ^ n_13542;
assign n_13942 = n_13880 ^ n_13543;
assign n_13943 = n_13881 ^ n_13544;
assign n_13944 = n_13882 ^ n_13556;
assign n_13945 = n_13883 ^ n_13545;
assign n_13946 = n_13884 ^ n_13546;
assign n_13947 = n_13885 ^ n_13547;
assign n_13948 = n_13886 ^ n_13548;
assign n_13949 = n_13887 ^ n_13557;
assign n_13950 = n_13888 ^ n_13549;
assign n_13951 = n_13889 ^ n_13550;
assign n_13952 = n_13890 ^ n_13551;
assign n_13953 = n_13891 ^ n_13552;
assign n_13954 = n_13892 ^ n_13553;
assign n_13955 = n_13893 ^ n_13554;
assign n_13956 = n_13497 ^ n_13894;
assign n_13957 = n_13495 ^ n_13895;
assign n_13958 = n_13833 & n_13896;
assign y64 = n_13896;
assign y66 = n_13897;
assign y67 = n_13898;
assign y68 = ~n_13899;
assign y69 = ~n_13900;
assign y70 = n_13901;
assign y71 = n_13902;
assign y72 = n_13903;
assign y73 = n_13904;
assign y74 = n_13905;
assign y75 = n_13906;
assign y76 = n_13907;
assign y78 = n_13908;
assign y79 = n_13909;
assign y80 = n_13910;
assign y81 = n_13911;
assign y82 = n_13912;
assign y83 = n_13913;
assign y84 = n_13914;
assign y85 = n_13915;
assign y86 = n_13916;
assign y88 = n_13917;
assign y89 = n_13918;
assign y90 = n_13919;
assign y91 = n_13920;
assign y92 = n_13921;
assign y93 = n_13922;
assign y94 = n_13923;
assign y95 = n_13924;
assign y96 = ~n_13925;
assign y97 = n_13926;
assign y98 = n_13927;
assign y99 = n_13928;
assign y100 = n_13929;
assign y101 = n_13930;
assign y102 = n_13931;
assign y103 = n_13932;
assign y104 = n_13933;
assign y105 = n_13934;
assign y106 = n_13935;
assign y107 = n_13936;
assign y108 = n_13937;
assign y109 = n_13938;
assign y110 = n_13939;
assign y111 = n_13940;
assign y112 = n_13941;
assign y113 = n_13942;
assign y114 = n_13943;
assign y115 = n_13944;
assign y116 = n_13945;
assign y117 = n_13946;
assign y118 = n_13947;
assign y119 = n_13948;
assign y120 = n_13949;
assign y121 = n_13950;
assign y122 = n_13951;
assign y123 = n_13952;
assign y124 = n_13953;
assign y125 = n_13954;
assign y126 = n_13955;
assign y77 = n_13956;
assign y87 = n_13957;
assign n_13959 = n_13834 ^ n_13958;
assign n_13960 = n_13959 ^ n_13438;
assign n_13961 = n_13960 ^ x1;
assign y65 = n_13961;
endmodule