module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 ;
  assign n17 = x0 & x8 ;
  assign n18 = x1 & x9 ;
  assign n19 = n17 & ~n18 ;
  assign n20 = ~x8 & n18 ;
  assign n21 = ~n19 & ~n20 ;
  assign n23 = x14 ^ x6 ;
  assign n22 = x7 & x15 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = x13 ^ x5 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = ~n25 & n26 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n24 & ~n28 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n30 ^ n22 ;
  assign n32 = x12 ^ x4 ;
  assign n33 = x11 ^ x3 ;
  assign n34 = n32 & n33 ;
  assign n35 = n31 & n34 ;
  assign n36 = n21 & n35 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = x9 ^ x1 ;
  assign n39 = x2 & x10 ;
  assign n40 = ~n38 & ~n39 ;
  assign n41 = n37 & n40 ;
  assign n42 = n41 ^ n37 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = x10 ^ x2 ;
  assign n52 = x4 & x12 ;
  assign n65 = x3 & x11 ;
  assign n66 = n52 & n65 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = n67 ^ n52 ;
  assign n45 = x5 & x13 ;
  assign n46 = x6 & x14 ;
  assign n47 = n45 & n46 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = n45 ^ x5 ;
  assign n51 = n50 ^ x13 ;
  assign n53 = n52 ^ x4 ;
  assign n54 = n53 ^ x12 ;
  assign n55 = n51 & n54 ;
  assign n56 = n55 ^ n51 ;
  assign n57 = n56 ^ n54 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = n58 ^ n54 ;
  assign n60 = n49 & n59 ;
  assign n61 = n60 ^ n49 ;
  assign n62 = n61 ^ n49 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n63 ^ n59 ;
  assign n69 = n68 ^ n64 ;
  assign n70 = ~x3 & ~x11 ;
  assign n71 = n52 & n70 ;
  assign n72 = n71 ^ n70 ;
  assign n73 = n72 ^ n64 ;
  assign n74 = n69 & n73 ;
  assign n75 = n74 ^ n69 ;
  assign n76 = n75 ^ n71 ;
  assign n77 = n76 ^ n64 ;
  assign n78 = n44 & n77 ;
  assign n79 = n78 ^ n44 ;
  assign n80 = n79 ^ n77 ;
  assign n81 = n20 & n35 ;
  assign n82 = n81 ^ n20 ;
  assign n83 = n82 ^ n35 ;
  assign n84 = n80 & ~n83 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = n85 ^ n80 ;
  assign n87 = n86 ^ n83 ;
  assign n88 = ~n43 & n87 ;
  assign n89 = ~x0 & ~x8 ;
  assign n90 = ~n18 & ~n39 ;
  assign n91 = ~n89 & n90 ;
  assign n92 = ~x2 & ~x10 ;
  assign n93 = n92 ^ n91 ;
  assign n94 = ~n91 & n93 ;
  assign n95 = n94 ^ n91 ;
  assign n96 = n95 ^ n77 ;
  assign n97 = n92 ^ n77 ;
  assign n98 = ~n96 & ~n97 ;
  assign n99 = n98 ^ n94 ;
  assign n100 = n99 ^ n77 ;
  assign n109 = x2 & ~n70 ;
  assign n110 = n109 ^ n68 ;
  assign n111 = ~n109 & n110 ;
  assign n112 = n111 ^ n109 ;
  assign n113 = n112 ^ n64 ;
  assign n114 = n69 & n113 ;
  assign n115 = n114 ^ n111 ;
  assign n116 = n115 ^ n64 ;
  assign n101 = ~x1 & ~x9 ;
  assign n102 = ~n17 & ~n101 ;
  assign n103 = ~n89 & ~n102 ;
  assign n104 = ~x0 & x10 ;
  assign n105 = n20 & n104 ;
  assign n106 = n105 ^ n103 ;
  assign n107 = n103 & n106 ;
  assign n108 = n107 ^ n103 ;
  assign n117 = n116 ^ n108 ;
  assign n118 = n116 ^ n105 ;
  assign n119 = n117 & n118 ;
  assign n120 = n119 ^ n107 ;
  assign n121 = n120 ^ n116 ;
  assign n122 = ~n100 & ~n121 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = n88 & n123 ;
  assign n125 = n124 ^ n88 ;
  assign n126 = n125 ^ n88 ;
  assign n127 = n126 ^ n123 ;
  assign n128 = n116 ^ n38 ;
  assign n129 = n70 ^ n68 ;
  assign n130 = n70 & n129 ;
  assign n131 = n130 ^ n68 ;
  assign n132 = n131 ^ n64 ;
  assign n133 = n64 & n132 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = n134 ^ n68 ;
  assign n136 = n135 ^ n44 ;
  assign n137 = n136 ^ n70 ;
  assign n138 = n128 & ~n137 ;
  assign n139 = n138 ^ n128 ;
  assign n142 = x8 ^ x0 ;
  assign n144 = n142 ^ n18 ;
  assign n145 = n144 ^ n35 ;
  assign n140 = n38 & n92 ;
  assign n141 = ~n101 & ~n140 ;
  assign n143 = n142 ^ n141 ;
  assign n146 = n145 ^ n143 ;
  assign n147 = n139 & n146 ;
  assign n148 = n147 ^ n143 ;
  assign n150 = n92 ^ n38 ;
  assign n149 = n128 ^ n35 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = ~n137 & n151 ;
  assign n153 = n152 ^ n151 ;
  assign n154 = n153 ^ n137 ;
  assign n155 = n154 ^ n150 ;
  assign n156 = n137 ^ n35 ;
  assign n157 = n22 & n23 ;
  assign n158 = ~n49 & ~n157 ;
  assign n159 = n51 & ~n158 ;
  assign n160 = ~n52 & ~n159 ;
  assign n161 = n54 & ~n160 ;
  assign n162 = n161 ^ n33 ;
  assign n163 = ~n31 & ~n46 ;
  assign n164 = n25 & ~n163 ;
  assign n165 = ~n45 & ~n164 ;
  assign n166 = n165 ^ n32 ;
  assign n167 = ~n46 & ~n157 ;
  assign n168 = n167 ^ n25 ;
  assign y0 = n127 ;
  assign y1 = n148 ;
  assign y2 = ~n155 ;
  assign y3 = n156 ;
  assign y4 = n162 ;
  assign y5 = ~n166 ;
  assign y6 = ~n168 ;
  assign y7 = n24 ;
endmodule
