module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 ;
  assign n151 = ~x5 & ~x22 ;
  assign n184 = ~x56 & n151 ;
  assign n148 = ~x4 & ~x19 ;
  assign n149 = ~x16 & ~x18 ;
  assign n150 = n148 & n149 ;
  assign n152 = ~x6 & ~x12 ;
  assign n153 = ~x17 & n152 ;
  assign n154 = n151 & n153 ;
  assign n155 = n150 & n154 ;
  assign n156 = ~x8 & ~x21 ;
  assign n157 = ~x7 & ~x13 ;
  assign n172 = x10 & n157 ;
  assign n173 = n156 & n172 ;
  assign n164 = ~x7 & ~x8 ;
  assign n166 = x21 & n164 ;
  assign n165 = x13 & n164 ;
  assign n167 = n166 ^ n165 ;
  assign n162 = ~x21 & n157 ;
  assign n160 = ~x8 & ~x13 ;
  assign n161 = ~x21 & n160 ;
  assign n163 = n162 ^ n161 ;
  assign n168 = n167 ^ n163 ;
  assign n169 = ~x10 & ~x14 ;
  assign n170 = n168 & n169 ;
  assign n158 = x14 & n157 ;
  assign n159 = n156 & n158 ;
  assign n171 = n170 ^ n159 ;
  assign n174 = n173 ^ n171 ;
  assign n175 = ~x9 & ~x11 ;
  assign n178 = ~x56 & n175 ;
  assign n179 = ~n151 & n178 ;
  assign n180 = n174 & n179 ;
  assign n181 = n155 & n180 ;
  assign n176 = n174 & n175 ;
  assign n177 = n155 & n176 ;
  assign n182 = n181 ^ n177 ;
  assign n183 = n182 ^ n178 ;
  assign n185 = n184 ^ n183 ;
  assign n200 = x54 & ~n185 ;
  assign n198 = x0 & ~x54 ;
  assign n186 = ~x14 & ~x22 ;
  assign n187 = n157 & n186 ;
  assign n188 = n175 & n187 ;
  assign n189 = ~x17 & ~x21 ;
  assign n190 = ~x8 & n189 ;
  assign n191 = ~x5 & n152 ;
  assign n192 = n190 & n191 ;
  assign n193 = n188 & n192 ;
  assign n194 = ~x0 & x54 ;
  assign n195 = n150 & n194 ;
  assign n196 = n193 & n195 ;
  assign n197 = ~n185 & n196 ;
  assign n199 = n198 ^ n197 ;
  assign n201 = n200 ^ n199 ;
  assign n202 = ~x3 & ~x129 ;
  assign n203 = ~n201 & n202 ;
  assign n204 = ~x5 & ~x6 ;
  assign n205 = ~x7 & ~x12 ;
  assign n206 = ~n204 & ~n205 ;
  assign n207 = ~x13 & ~n206 ;
  assign n208 = ~x5 & ~x7 ;
  assign n209 = n208 ^ n152 ;
  assign n210 = n207 & n209 ;
  assign n211 = x13 & n152 ;
  assign n212 = n208 & n211 ;
  assign n213 = ~x9 & ~n212 ;
  assign n214 = ~n210 & n213 ;
  assign n215 = n157 & n191 ;
  assign n216 = x9 & ~n215 ;
  assign n217 = ~x10 & x54 ;
  assign n218 = n186 & n217 ;
  assign n219 = ~x8 & ~x11 ;
  assign n220 = n189 & n219 ;
  assign n221 = n218 & n220 ;
  assign n222 = n150 & n221 ;
  assign n223 = ~n216 & n222 ;
  assign n224 = ~n214 & n223 ;
  assign n225 = n157 & n204 ;
  assign n226 = n150 & n225 ;
  assign n227 = ~x14 & n156 ;
  assign n228 = ~x11 & ~x12 ;
  assign n229 = ~x10 & ~x22 ;
  assign n230 = n228 & n229 ;
  assign n231 = n227 & n230 ;
  assign n232 = n226 & n231 ;
  assign n233 = ~x17 & x54 ;
  assign n234 = ~x1 & n233 ;
  assign n235 = ~n232 & n234 ;
  assign n236 = n235 ^ x1 ;
  assign n237 = n202 & n236 ;
  assign n238 = ~n224 & n237 ;
  assign n239 = n238 ^ n202 ;
  assign n240 = ~x38 & ~x50 ;
  assign n241 = ~x40 & ~x46 ;
  assign n242 = n240 & n241 ;
  assign n243 = x41 & x43 ;
  assign n244 = n243 ^ x41 ;
  assign n245 = n244 ^ x43 ;
  assign n246 = ~x42 & ~x44 ;
  assign n247 = ~n245 & n246 ;
  assign n248 = n242 & n247 ;
  assign n249 = ~x47 & ~x48 ;
  assign n250 = n248 & n249 ;
  assign n251 = x15 & x20 ;
  assign n252 = n251 ^ x15 ;
  assign n253 = n252 ^ x20 ;
  assign n254 = x45 & n253 ;
  assign n255 = n254 ^ x45 ;
  assign n256 = n255 ^ n253 ;
  assign n257 = x24 & x49 ;
  assign n258 = n257 ^ x24 ;
  assign n259 = n258 ^ x49 ;
  assign n260 = x82 & ~n259 ;
  assign n261 = ~n256 & n260 ;
  assign n262 = x122 & x127 ;
  assign n263 = ~x82 & ~n262 ;
  assign n264 = x2 & ~n263 ;
  assign n265 = n261 & n264 ;
  assign n266 = n250 & n265 ;
  assign n267 = n266 ^ n264 ;
  assign n272 = ~n256 & n259 ;
  assign n273 = n272 ^ n256 ;
  assign n274 = ~x41 & ~x46 ;
  assign n275 = n240 & n274 ;
  assign n276 = ~x43 & ~x47 ;
  assign n277 = ~x2 & ~x48 ;
  assign n278 = n276 & n277 ;
  assign n279 = n275 & n278 ;
  assign n280 = ~n273 & n279 ;
  assign n281 = ~x40 & n246 ;
  assign n268 = ~x65 & ~n262 ;
  assign n282 = x82 & n268 ;
  assign n283 = n281 & n282 ;
  assign n284 = n280 & n283 ;
  assign n285 = ~n267 & n284 ;
  assign n269 = ~x82 & n268 ;
  assign n270 = ~n267 & n269 ;
  assign n271 = n270 ^ n267 ;
  assign n286 = n285 ^ n271 ;
  assign n287 = ~x129 & n286 ;
  assign n294 = ~x9 & ~x14 ;
  assign n295 = n229 & n294 ;
  assign n296 = ~x12 & n220 ;
  assign n297 = n295 & n296 ;
  assign n288 = x0 & ~x113 ;
  assign n289 = ~x123 & n288 ;
  assign n290 = ~x61 & ~x118 ;
  assign n298 = ~x129 & n290 ;
  assign n299 = ~n289 & n298 ;
  assign n300 = n226 & n299 ;
  assign n301 = n297 & n300 ;
  assign n291 = ~x129 & ~n290 ;
  assign n292 = ~n289 & n291 ;
  assign n293 = n292 ^ x129 ;
  assign n302 = n301 ^ n293 ;
  assign n312 = x4 & ~x54 ;
  assign n316 = n202 & n312 ;
  assign n303 = ~x18 & n148 ;
  assign n304 = ~x16 & x54 ;
  assign n305 = n189 & n304 ;
  assign n306 = n303 & n305 ;
  assign n307 = x10 & ~x22 ;
  assign n308 = n219 & n307 ;
  assign n309 = n306 & n308 ;
  assign n310 = n157 & n294 ;
  assign n311 = n191 & n310 ;
  assign n313 = n202 & ~n312 ;
  assign n314 = n311 & n313 ;
  assign n315 = n309 & n314 ;
  assign n317 = n316 ^ n315 ;
  assign n318 = x5 & ~x54 ;
  assign n319 = ~x13 & n295 ;
  assign n320 = ~x59 & n220 ;
  assign n321 = n319 & n320 ;
  assign n322 = n152 & n208 ;
  assign n323 = n304 & n322 ;
  assign n324 = ~x25 & x28 ;
  assign n325 = ~x29 & n324 ;
  assign n326 = n303 & n325 ;
  assign n327 = n323 & n326 ;
  assign n328 = n321 & n327 ;
  assign n329 = ~n318 & ~n328 ;
  assign n330 = n202 & ~n329 ;
  assign n331 = x6 & ~x54 ;
  assign n332 = ~x28 & ~x29 ;
  assign n333 = x25 & n332 ;
  assign n334 = n303 & n333 ;
  assign n335 = n323 & n334 ;
  assign n336 = n321 & n335 ;
  assign n337 = ~n331 & ~n336 ;
  assign n338 = n202 & ~n337 ;
  assign n339 = x7 & ~x54 ;
  assign n340 = x8 & n306 ;
  assign n341 = ~x11 & n322 ;
  assign n342 = n319 & n341 ;
  assign n343 = n340 & n342 ;
  assign n344 = ~n339 & ~n343 ;
  assign n345 = n202 & ~n344 ;
  assign n346 = x8 & ~x54 ;
  assign n347 = ~x12 & n295 ;
  assign n348 = n225 & n347 ;
  assign n349 = n148 & n304 ;
  assign n350 = ~x17 & ~x18 ;
  assign n351 = n219 & n350 ;
  assign n352 = x21 & n351 ;
  assign n353 = n349 & n352 ;
  assign n354 = n348 & n353 ;
  assign n355 = ~n346 & ~n354 ;
  assign n356 = n202 & ~n355 ;
  assign n357 = x9 & ~x54 ;
  assign n358 = ~x8 & n306 ;
  assign n359 = x11 & n322 ;
  assign n360 = n319 & n359 ;
  assign n361 = n358 & n360 ;
  assign n362 = ~n357 & ~n361 ;
  assign n363 = n202 & ~n362 ;
  assign n364 = x10 & ~x54 ;
  assign n365 = ~x9 & ~x18 ;
  assign n366 = n190 & n365 ;
  assign n367 = n229 & n366 ;
  assign n368 = ~x13 & x14 ;
  assign n369 = n349 & n368 ;
  assign n370 = n341 & n369 ;
  assign n371 = n367 & n370 ;
  assign n372 = ~n364 & ~n371 ;
  assign n373 = n202 & ~n372 ;
  assign n376 = x11 & ~x54 ;
  assign n381 = n202 & n376 ;
  assign n374 = ~x10 & ~x11 ;
  assign n375 = x22 & n374 ;
  assign n377 = n202 & ~n376 ;
  assign n378 = n375 & n377 ;
  assign n379 = n311 & n378 ;
  assign n380 = n358 & n379 ;
  assign n382 = n381 ^ n380 ;
  assign n383 = x12 & ~x54 ;
  assign n384 = x18 & n225 ;
  assign n385 = n295 & n349 ;
  assign n386 = n384 & n385 ;
  assign n387 = n296 & n386 ;
  assign n388 = ~n383 & ~n387 ;
  assign n389 = n202 & ~n388 ;
  assign n390 = ~x25 & ~x28 ;
  assign n391 = x29 & n390 ;
  assign n392 = ~x59 & n229 ;
  assign n393 = n391 & n392 ;
  assign n394 = n306 & n393 ;
  assign n395 = x13 & ~x54 ;
  assign n396 = n219 & ~n395 ;
  assign n397 = n311 & n396 ;
  assign n398 = n394 & n397 ;
  assign n399 = n398 ^ n395 ;
  assign n400 = n202 & n399 ;
  assign n401 = x14 & ~x54 ;
  assign n402 = x13 & ~x16 ;
  assign n403 = n148 & n402 ;
  assign n404 = n218 & n403 ;
  assign n405 = n341 & n404 ;
  assign n406 = n366 & n405 ;
  assign n407 = ~n401 & ~n406 ;
  assign n408 = n202 & ~n407 ;
  assign n413 = ~x70 & ~n262 ;
  assign n416 = n413 ^ x82 ;
  assign n411 = ~x82 & n262 ;
  assign n412 = x15 & n411 ;
  assign n433 = n416 ^ n412 ;
  assign n420 = x45 & n259 ;
  assign n421 = n420 ^ x45 ;
  assign n422 = n421 ^ n259 ;
  assign n423 = x15 & ~n245 ;
  assign n424 = n423 ^ n245 ;
  assign n425 = n249 & ~n424 ;
  assign n426 = n422 & n425 ;
  assign n427 = n426 ^ n425 ;
  assign n409 = n242 & n246 ;
  assign n417 = n413 ^ n409 ;
  assign n418 = n416 & n417 ;
  assign n419 = n418 ^ n409 ;
  assign n428 = n427 ^ n419 ;
  assign n434 = n433 ^ n428 ;
  assign n435 = n427 ^ x82 ;
  assign n436 = n435 ^ n419 ;
  assign n437 = ~n434 & n436 ;
  assign n429 = n419 ^ x82 ;
  assign n414 = n413 ^ n412 ;
  assign n430 = n429 ^ n414 ;
  assign n431 = n428 & ~n430 ;
  assign n438 = n437 ^ n431 ;
  assign n439 = n438 ^ n419 ;
  assign n440 = n439 ^ n433 ;
  assign n441 = n431 ^ n427 ;
  assign n442 = n441 ^ n412 ;
  assign n443 = ~n440 & ~n442 ;
  assign n444 = n443 ^ n437 ;
  assign n432 = n431 ^ n418 ;
  assign n445 = n444 ^ n432 ;
  assign n410 = n409 ^ x82 ;
  assign n415 = n414 ^ n410 ;
  assign n446 = n445 ^ n415 ;
  assign n447 = n446 ^ n412 ;
  assign n468 = n447 ^ x129 ;
  assign n469 = x129 & n468 ;
  assign n448 = ~x48 & n276 ;
  assign n449 = ~n422 & n448 ;
  assign n450 = x15 & ~x40 ;
  assign n451 = n246 & n450 ;
  assign n452 = n275 & n451 ;
  assign n453 = n449 & n452 ;
  assign n454 = n453 ^ x15 ;
  assign n455 = ~x2 & ~x20 ;
  assign n456 = ~n259 & ~n455 ;
  assign n457 = ~x15 & ~x45 ;
  assign n458 = n249 & n457 ;
  assign n459 = n456 & n458 ;
  assign n460 = n248 & n459 ;
  assign n461 = ~n454 & ~n460 ;
  assign n465 = x82 & ~n461 ;
  assign n462 = x82 & ~x129 ;
  assign n463 = ~n461 & n462 ;
  assign n464 = n447 & n463 ;
  assign n466 = n465 ^ n464 ;
  assign n467 = n466 ^ n447 ;
  assign n470 = n469 ^ n467 ;
  assign n471 = n470 ^ n465 ;
  assign n472 = x16 & ~x54 ;
  assign n473 = n219 & n306 ;
  assign n474 = x6 & ~x13 ;
  assign n475 = n208 & n474 ;
  assign n476 = n347 & n475 ;
  assign n477 = n473 & n476 ;
  assign n478 = ~n472 & ~n477 ;
  assign n479 = n202 & ~n478 ;
  assign n480 = x17 & ~x54 ;
  assign n481 = ~x25 & x59 ;
  assign n482 = n156 & n481 ;
  assign n483 = n233 & n332 ;
  assign n484 = n482 & n483 ;
  assign n485 = n150 & n484 ;
  assign n486 = n342 & n485 ;
  assign n487 = ~n480 & ~n486 ;
  assign n488 = n202 & ~n487 ;
  assign n493 = x18 & ~x54 ;
  assign n497 = n202 & n493 ;
  assign n489 = n225 & n303 ;
  assign n490 = n347 & n489 ;
  assign n491 = x16 & x54 ;
  assign n492 = n220 & n491 ;
  assign n494 = n202 & ~n493 ;
  assign n495 = n492 & n494 ;
  assign n496 = n490 & n495 ;
  assign n498 = n497 ^ n496 ;
  assign n502 = x19 & ~x54 ;
  assign n506 = n202 & n502 ;
  assign n499 = x17 & ~x21 ;
  assign n500 = n219 & n499 ;
  assign n501 = n304 & n500 ;
  assign n503 = n202 & ~n502 ;
  assign n504 = n501 & n503 ;
  assign n505 = n490 & n504 ;
  assign n507 = n506 ^ n505 ;
  assign n523 = x20 & x82 ;
  assign n508 = ~x46 & ~x50 ;
  assign n509 = ~x38 & ~x40 ;
  assign n510 = n246 & n509 ;
  assign n511 = n508 & n510 ;
  assign n512 = ~x45 & n249 ;
  assign n513 = ~n245 & ~n259 ;
  assign n514 = n512 & n513 ;
  assign n515 = n511 & n514 ;
  assign n520 = ~x15 & x82 ;
  assign n521 = n515 & n520 ;
  assign n516 = ~x2 & ~x15 ;
  assign n517 = ~x20 & x82 ;
  assign n518 = n516 & n517 ;
  assign n519 = n515 & n518 ;
  assign n522 = n521 ^ n519 ;
  assign n524 = n523 ^ n522 ;
  assign n525 = x20 & n411 ;
  assign n526 = ~x71 & ~n262 ;
  assign n530 = x82 & ~n253 ;
  assign n531 = n526 & n530 ;
  assign n532 = ~n525 & n531 ;
  assign n533 = n515 & n532 ;
  assign n527 = ~x82 & n526 ;
  assign n528 = ~n525 & n527 ;
  assign n529 = n528 ^ n525 ;
  assign n534 = n533 ^ n529 ;
  assign n535 = ~n524 & ~n534 ;
  assign n536 = ~x129 & ~n535 ;
  assign n537 = x21 & ~x54 ;
  assign n538 = ~x4 & x19 ;
  assign n539 = ~x21 & n538 ;
  assign n540 = n304 & n539 ;
  assign n541 = n351 & n540 ;
  assign n542 = n348 & n541 ;
  assign n543 = ~n537 & ~n542 ;
  assign n544 = n202 & ~n543 ;
  assign n545 = x22 & ~x54 ;
  assign n546 = x5 & ~x6 ;
  assign n547 = ~x14 & n546 ;
  assign n548 = n157 & n228 ;
  assign n549 = n547 & n548 ;
  assign n550 = n349 & n549 ;
  assign n551 = n367 & n550 ;
  assign n552 = ~n545 & ~n551 ;
  assign n553 = n202 & ~n552 ;
  assign n554 = ~x23 & x55 ;
  assign n555 = x61 & ~x129 ;
  assign n556 = ~n554 & n555 ;
  assign n563 = ~n245 & n512 ;
  assign n567 = x24 & x82 ;
  assign n568 = n508 & n567 ;
  assign n569 = n510 & n568 ;
  assign n570 = n563 & n569 ;
  assign n571 = ~x129 & ~n570 ;
  assign n557 = x2 & n253 ;
  assign n558 = n557 ^ x2 ;
  assign n559 = n558 ^ n253 ;
  assign n572 = ~x45 & ~x49 ;
  assign n573 = n249 & n572 ;
  assign n574 = ~n559 & n573 ;
  assign n575 = n248 & n574 ;
  assign n576 = x63 & ~n262 ;
  assign n577 = x82 & n576 ;
  assign n584 = ~n575 & n577 ;
  assign n585 = n584 ^ n576 ;
  assign n586 = n571 & ~n585 ;
  assign n560 = ~x49 & ~n559 ;
  assign n561 = x82 & ~n560 ;
  assign n562 = n262 & ~n561 ;
  assign n564 = n409 & n563 ;
  assign n565 = x82 & ~n564 ;
  assign n566 = ~n562 & ~n565 ;
  assign n580 = ~x24 & ~n576 ;
  assign n578 = ~x24 & n577 ;
  assign n579 = ~n575 & n578 ;
  assign n581 = n580 ^ n579 ;
  assign n582 = n571 & n581 ;
  assign n583 = ~n566 & n582 ;
  assign n587 = n586 ^ n583 ;
  assign n638 = x58 ^ x53 ;
  assign n641 = n638 ^ x53 ;
  assign n631 = ~x53 & ~x58 ;
  assign n632 = ~x27 & ~x85 ;
  assign n633 = x25 & ~x116 ;
  assign n634 = ~x26 & n633 ;
  assign n635 = n632 & n634 ;
  assign n636 = ~n631 & ~n635 ;
  assign n637 = n202 & ~n636 ;
  assign n667 = n641 ^ n637 ;
  assign n645 = ~x95 & ~x100 ;
  assign n646 = ~x97 & ~x110 ;
  assign n647 = n645 & n646 ;
  assign n648 = n647 ^ x110 ;
  assign n649 = x25 & n648 ;
  assign n658 = ~x27 & ~n649 ;
  assign n609 = x39 & x52 ;
  assign n610 = n609 ^ x39 ;
  assign n611 = n610 ^ x52 ;
  assign n612 = ~x51 & x116 ;
  assign n613 = ~n611 & n612 ;
  assign n650 = n633 ^ n613 ;
  assign n656 = x27 & ~n650 ;
  assign n651 = ~x51 & ~x52 ;
  assign n652 = x27 & ~x39 ;
  assign n653 = n651 & n652 ;
  assign n654 = ~n650 & n653 ;
  assign n655 = n649 & n654 ;
  assign n657 = n656 ^ n655 ;
  assign n659 = n658 ^ n657 ;
  assign n660 = ~x26 & ~x85 ;
  assign n661 = ~n659 & n660 ;
  assign n598 = x100 & ~x116 ;
  assign n591 = x116 ^ x110 ;
  assign n590 = x116 ^ x96 ;
  assign n592 = n591 ^ n590 ;
  assign n593 = n590 ^ x116 ;
  assign n594 = n592 & ~n593 ;
  assign n595 = n594 ^ n590 ;
  assign n596 = ~x85 & x100 ;
  assign n597 = ~n595 & n596 ;
  assign n599 = n598 ^ n597 ;
  assign n600 = n599 ^ x100 ;
  assign n588 = x85 & ~x116 ;
  assign n589 = x25 & n588 ;
  assign n601 = n600 ^ n589 ;
  assign n602 = x25 & x26 ;
  assign n603 = n588 & n602 ;
  assign n604 = n603 ^ x26 ;
  assign n605 = n604 ^ n600 ;
  assign n606 = n601 & ~n605 ;
  assign n607 = n606 ^ n603 ;
  assign n608 = n607 ^ n600 ;
  assign n614 = x26 & ~x85 ;
  assign n624 = ~n613 & n614 ;
  assign n618 = ~x25 & ~x116 ;
  assign n619 = n614 & n618 ;
  assign n625 = n624 ^ n619 ;
  assign n626 = n608 & n625 ;
  assign n627 = n626 ^ n608 ;
  assign n628 = n627 ^ n625 ;
  assign n620 = x27 & ~n619 ;
  assign n621 = ~n608 & n620 ;
  assign n615 = x27 & n614 ;
  assign n616 = ~n613 & n615 ;
  assign n617 = ~n608 & n616 ;
  assign n622 = n621 ^ n617 ;
  assign n623 = n622 ^ x27 ;
  assign n629 = n628 ^ n623 ;
  assign n642 = n638 ^ n629 ;
  assign n643 = n641 & n642 ;
  assign n644 = n643 ^ n629 ;
  assign n662 = n661 ^ n644 ;
  assign n668 = n667 ^ n662 ;
  assign n669 = n661 ^ x53 ;
  assign n670 = n669 ^ n644 ;
  assign n671 = n668 & ~n670 ;
  assign n663 = n644 ^ x53 ;
  assign n639 = n638 ^ n637 ;
  assign n664 = n663 ^ n639 ;
  assign n665 = n662 & ~n664 ;
  assign n672 = n671 ^ n665 ;
  assign n673 = n672 ^ n644 ;
  assign n674 = n673 ^ n667 ;
  assign n675 = n665 ^ n661 ;
  assign n676 = n675 ^ n637 ;
  assign n677 = ~n674 & ~n676 ;
  assign n678 = n677 ^ n671 ;
  assign n666 = n665 ^ n643 ;
  assign n679 = n678 ^ n666 ;
  assign n630 = n629 ^ x53 ;
  assign n640 = n639 ^ n630 ;
  assign n680 = n679 ^ n640 ;
  assign n681 = n680 ^ n637 ;
  assign n682 = x26 & x116 ;
  assign n683 = n600 & ~n682 ;
  assign n684 = ~n624 & ~n683 ;
  assign n685 = ~x27 & ~x53 ;
  assign n686 = ~x58 & n685 ;
  assign n687 = n202 & n686 ;
  assign n688 = ~n684 & n687 ;
  assign n689 = x85 & n613 ;
  assign n690 = n689 ^ x85 ;
  assign n691 = n690 ^ n613 ;
  assign n692 = x27 & ~n691 ;
  assign n693 = x85 & x116 ;
  assign n694 = x85 & x110 ;
  assign n695 = n694 ^ x85 ;
  assign n696 = n695 ^ x110 ;
  assign n697 = x95 & ~x96 ;
  assign n698 = ~n696 & n697 ;
  assign n699 = ~n693 & ~n698 ;
  assign n700 = ~x27 & ~x100 ;
  assign n701 = ~n699 & n700 ;
  assign n702 = ~n692 & ~n701 ;
  assign n703 = ~x26 & n202 ;
  assign n704 = n631 & n703 ;
  assign n705 = ~n702 & n704 ;
  assign n715 = x51 & ~n611 ;
  assign n716 = n715 ^ n611 ;
  assign n717 = n682 & ~n716 ;
  assign n720 = ~x26 & ~x100 ;
  assign n721 = ~x110 & n720 ;
  assign n722 = n632 & n697 ;
  assign n723 = n721 & n722 ;
  assign n724 = ~n717 & n723 ;
  assign n718 = n632 & n717 ;
  assign n719 = n718 ^ x85 ;
  assign n725 = n724 ^ n719 ;
  assign n726 = n653 ^ x27 ;
  assign n727 = ~x26 & x116 ;
  assign n728 = n726 & n727 ;
  assign n729 = ~n725 & n728 ;
  assign n730 = n729 ^ n725 ;
  assign n734 = ~x26 & ~x39 ;
  assign n735 = n651 & n734 ;
  assign n731 = ~x27 & ~x39 ;
  assign n732 = n651 & n731 ;
  assign n733 = n732 ^ x26 ;
  assign n736 = n735 ^ n733 ;
  assign n737 = n648 & ~n736 ;
  assign n738 = x27 ^ x26 ;
  assign n739 = ~x116 & n738 ;
  assign n740 = x28 & ~n739 ;
  assign n741 = ~n737 & n740 ;
  assign n742 = n741 ^ x28 ;
  assign n743 = x100 & x116 ;
  assign n744 = ~x26 & ~x27 ;
  assign n745 = ~x28 & ~x116 ;
  assign n746 = n744 & ~n745 ;
  assign n747 = ~n743 & n746 ;
  assign n752 = ~x53 & ~x85 ;
  assign n753 = ~n747 & n752 ;
  assign n754 = ~n742 & n753 ;
  assign n755 = ~n730 & n754 ;
  assign n756 = n755 ^ n753 ;
  assign n748 = ~x53 & n747 ;
  assign n749 = ~n742 & n748 ;
  assign n750 = ~n730 & n749 ;
  assign n751 = n750 ^ n748 ;
  assign n757 = n756 ^ n751 ;
  assign n706 = ~x26 & ~x53 ;
  assign n707 = ~x85 & n706 ;
  assign n708 = ~x27 & x28 ;
  assign n709 = ~x116 & n708 ;
  assign n710 = x58 & n709 ;
  assign n711 = n707 & n710 ;
  assign n758 = x53 & n660 ;
  assign n759 = n709 & n758 ;
  assign n760 = ~x58 & n202 ;
  assign n761 = ~n759 & n760 ;
  assign n762 = ~n711 & n761 ;
  assign n763 = ~n757 & n762 ;
  assign n712 = x58 & n202 ;
  assign n713 = ~n711 & n712 ;
  assign n714 = n713 ^ n202 ;
  assign n764 = n763 ^ n714 ;
  assign n765 = x29 & ~x116 ;
  assign n786 = x53 & ~x58 ;
  assign n787 = n765 & n786 ;
  assign n791 = ~x27 & n787 ;
  assign n772 = ~x96 & ~x110 ;
  assign n773 = x97 & ~n772 ;
  assign n774 = x29 & ~x110 ;
  assign n775 = n645 & n774 ;
  assign n776 = ~n773 & n775 ;
  assign n771 = x29 & x110 ;
  assign n777 = n776 ^ n771 ;
  assign n778 = ~x58 & x97 ;
  assign n779 = n645 & n778 ;
  assign n780 = ~n773 & n779 ;
  assign n781 = n780 ^ x58 ;
  assign n782 = ~n777 & ~n781 ;
  assign n783 = x97 & x116 ;
  assign n784 = x58 & ~n765 ;
  assign n785 = ~n783 & n784 ;
  assign n788 = n685 & ~n787 ;
  assign n789 = ~n785 & n788 ;
  assign n790 = ~n782 & n789 ;
  assign n792 = n791 ^ n790 ;
  assign n766 = x85 & n765 ;
  assign n767 = n686 & n766 ;
  assign n793 = x27 & n631 ;
  assign n794 = n765 & n793 ;
  assign n795 = n660 & ~n794 ;
  assign n796 = ~n767 & n795 ;
  assign n797 = ~n792 & n796 ;
  assign n768 = ~x26 & x85 ;
  assign n769 = ~n767 & n768 ;
  assign n770 = n769 ^ x26 ;
  assign n798 = n797 ^ n770 ;
  assign n799 = x26 & ~x27 ;
  assign n800 = ~x85 & n631 ;
  assign n801 = n799 & n800 ;
  assign n802 = n765 & n801 ;
  assign n803 = n202 & ~n802 ;
  assign n804 = n798 & n803 ;
  assign n805 = n804 ^ n202 ;
  assign n806 = ~x30 & ~x109 ;
  assign n807 = ~x60 & x109 ;
  assign n808 = ~n806 & ~n807 ;
  assign n809 = ~x106 & ~n808 ;
  assign n810 = ~x88 & x106 ;
  assign n811 = ~x129 & ~n810 ;
  assign n812 = ~n809 & n811 ;
  assign n813 = ~x31 & ~x109 ;
  assign n814 = ~x30 & x109 ;
  assign n815 = ~n813 & ~n814 ;
  assign n816 = ~x106 & ~n815 ;
  assign n817 = ~x89 & x106 ;
  assign n818 = ~x129 & ~n817 ;
  assign n819 = ~n816 & n818 ;
  assign n820 = ~x32 & ~x109 ;
  assign n821 = ~x31 & x109 ;
  assign n822 = ~n820 & ~n821 ;
  assign n823 = ~x106 & ~n822 ;
  assign n824 = ~x99 & x106 ;
  assign n825 = ~x129 & ~n824 ;
  assign n826 = ~n823 & n825 ;
  assign n827 = ~x33 & ~x109 ;
  assign n828 = ~x32 & x109 ;
  assign n829 = ~n827 & ~n828 ;
  assign n830 = ~x106 & ~n829 ;
  assign n831 = ~x90 & x106 ;
  assign n832 = ~x129 & ~n831 ;
  assign n833 = ~n830 & n832 ;
  assign n834 = ~x34 & ~x109 ;
  assign n835 = ~x33 & x109 ;
  assign n836 = ~n834 & ~n835 ;
  assign n837 = ~x106 & ~n836 ;
  assign n838 = ~x91 & x106 ;
  assign n839 = ~x129 & ~n838 ;
  assign n840 = ~n837 & n839 ;
  assign n841 = ~x35 & ~x109 ;
  assign n842 = ~x34 & x109 ;
  assign n843 = ~n841 & ~n842 ;
  assign n844 = ~x106 & ~n843 ;
  assign n845 = ~x92 & x106 ;
  assign n846 = ~x129 & ~n845 ;
  assign n847 = ~n844 & n846 ;
  assign n848 = ~x36 & ~x109 ;
  assign n849 = ~x35 & x109 ;
  assign n850 = ~n848 & ~n849 ;
  assign n851 = ~x106 & ~n850 ;
  assign n852 = ~x98 & x106 ;
  assign n853 = ~x129 & ~n852 ;
  assign n854 = ~n851 & n853 ;
  assign n855 = ~x37 & ~x109 ;
  assign n856 = ~x36 & x109 ;
  assign n857 = ~n855 & ~n856 ;
  assign n858 = ~x106 & ~n857 ;
  assign n859 = ~x93 & x106 ;
  assign n860 = ~x129 & ~n859 ;
  assign n861 = ~n858 & n860 ;
  assign n862 = ~x24 & ~x45 ;
  assign n863 = ~x49 & ~x50 ;
  assign n864 = n862 & n863 ;
  assign n865 = ~n559 & n864 ;
  assign n866 = n274 & n276 ;
  assign n867 = ~x48 & x82 ;
  assign n868 = n866 & n867 ;
  assign n869 = n865 & n868 ;
  assign n870 = n869 ^ x82 ;
  assign n871 = x82 & ~n281 ;
  assign n872 = n262 & ~n871 ;
  assign n873 = ~n870 & n872 ;
  assign n874 = n873 ^ n871 ;
  assign n875 = x38 & ~n874 ;
  assign n876 = n875 ^ x38 ;
  assign n877 = n876 ^ n874 ;
  assign n888 = ~x44 & x82 ;
  assign n889 = ~x40 & ~x42 ;
  assign n890 = x38 & n889 ;
  assign n891 = n888 & n890 ;
  assign n892 = ~x129 & ~n891 ;
  assign n886 = x74 & ~n262 ;
  assign n893 = n892 ^ n886 ;
  assign n894 = ~n892 & ~n893 ;
  assign n895 = n894 ^ n892 ;
  assign n878 = ~x48 & ~x49 ;
  assign n879 = n862 & n878 ;
  assign n880 = ~n559 & n879 ;
  assign n881 = ~x50 & n866 ;
  assign n882 = n880 & n881 ;
  assign n883 = x82 & n281 ;
  assign n884 = n882 & n883 ;
  assign n885 = n884 ^ x82 ;
  assign n896 = n895 ^ n885 ;
  assign n887 = n886 ^ n885 ;
  assign n897 = n896 ^ n887 ;
  assign n898 = n897 ^ n894 ;
  assign n899 = n898 ^ n885 ;
  assign n900 = n877 & ~n899 ;
  assign n901 = n900 ^ n899 ;
  assign n902 = x109 & n651 ;
  assign n903 = x39 & ~n902 ;
  assign n904 = ~x51 & x109 ;
  assign n905 = ~n611 & n904 ;
  assign n906 = ~x106 & ~n905 ;
  assign n907 = ~n903 & n906 ;
  assign n908 = ~x129 & ~n907 ;
  assign n911 = n261 & n279 ;
  assign n912 = n911 ^ x82 ;
  assign n909 = x82 & ~n246 ;
  assign n913 = ~x40 & n262 ;
  assign n914 = ~n909 & n913 ;
  assign n915 = ~n912 & n914 ;
  assign n910 = ~x40 & n909 ;
  assign n916 = n915 ^ n910 ;
  assign n917 = ~x42 & n888 ;
  assign n918 = x40 & n917 ;
  assign n919 = ~x129 & ~n918 ;
  assign n920 = ~n916 & n919 ;
  assign n923 = n422 & n559 ;
  assign n924 = n923 ^ n422 ;
  assign n925 = n924 ^ n559 ;
  assign n926 = ~x46 & ~n245 ;
  assign n927 = n240 & n249 ;
  assign n928 = n926 & n927 ;
  assign n929 = ~n925 & n928 ;
  assign n930 = n246 & n929 ;
  assign n921 = x73 & ~n262 ;
  assign n931 = x82 & n921 ;
  assign n932 = ~n930 & n931 ;
  assign n933 = n920 & n932 ;
  assign n922 = n920 & ~n921 ;
  assign n934 = n933 ^ n922 ;
  assign n936 = x76 & ~n262 ;
  assign n940 = ~x82 & n936 ;
  assign n935 = ~n273 & n278 ;
  assign n937 = x82 & n936 ;
  assign n938 = n511 & n937 ;
  assign n939 = n935 & n938 ;
  assign n941 = n940 ^ n939 ;
  assign n942 = x82 & n262 ;
  assign n943 = n278 & n942 ;
  assign n944 = ~n273 & n943 ;
  assign n945 = n944 ^ n942 ;
  assign n946 = n945 ^ n262 ;
  assign n950 = ~x41 & ~x82 ;
  assign n947 = ~x41 & x82 ;
  assign n948 = n246 & n947 ;
  assign n949 = n242 & n948 ;
  assign n951 = n950 ^ n949 ;
  assign n952 = ~n946 & n951 ;
  assign n953 = n952 ^ x41 ;
  assign n954 = x41 & n917 ;
  assign n955 = n242 & n954 ;
  assign n956 = ~x129 & ~n955 ;
  assign n957 = ~n953 & n956 ;
  assign n958 = n957 ^ n956 ;
  assign n959 = n941 & n958 ;
  assign n960 = n959 ^ n958 ;
  assign n978 = x42 & n888 ;
  assign n979 = ~x129 & ~n978 ;
  assign n982 = n979 ^ x72 ;
  assign n962 = x44 & x82 ;
  assign n963 = n262 & ~n962 ;
  assign n968 = ~x40 & x82 ;
  assign n969 = n963 & n968 ;
  assign n974 = n929 & n969 ;
  assign n964 = ~x82 & n963 ;
  assign n975 = n974 ^ n964 ;
  assign n976 = n975 ^ n962 ;
  assign n970 = x42 & n969 ;
  assign n971 = n929 & n970 ;
  assign n966 = x42 & ~n962 ;
  assign n965 = x42 & n964 ;
  assign n967 = n966 ^ n965 ;
  assign n972 = n971 ^ n967 ;
  assign n973 = n972 ^ x42 ;
  assign n977 = n976 ^ n973 ;
  assign n992 = n982 ^ n977 ;
  assign n986 = n889 & n929 ;
  assign n983 = n979 ^ n263 ;
  assign n984 = n982 & ~n983 ;
  assign n985 = n984 ^ n263 ;
  assign n987 = n986 ^ n985 ;
  assign n993 = n992 ^ n987 ;
  assign n994 = n986 ^ x72 ;
  assign n995 = n994 ^ n985 ;
  assign n996 = ~n993 & n995 ;
  assign n988 = n985 ^ x72 ;
  assign n980 = n979 ^ n977 ;
  assign n989 = n988 ^ n980 ;
  assign n990 = n987 & n989 ;
  assign n997 = n996 ^ n990 ;
  assign n998 = n997 ^ n985 ;
  assign n999 = n998 ^ n992 ;
  assign n1000 = n990 ^ n986 ;
  assign n1001 = n1000 ^ n977 ;
  assign n1002 = n999 & n1001 ;
  assign n1003 = n1002 ^ n996 ;
  assign n991 = n990 ^ n984 ;
  assign n1004 = n1003 ^ n991 ;
  assign n961 = n263 ^ x72 ;
  assign n981 = n980 ^ n961 ;
  assign n1005 = n1004 ^ n981 ;
  assign n1006 = ~n259 & n455 ;
  assign n1007 = n458 & n1006 ;
  assign n1009 = n411 & ~n1007 ;
  assign n1008 = n262 & n1007 ;
  assign n1010 = n1009 ^ n1008 ;
  assign n1012 = n275 & n281 ;
  assign n1013 = ~x43 & x82 ;
  assign n1014 = ~n1012 & n1013 ;
  assign n1015 = ~n1010 & n1014 ;
  assign n1011 = ~x43 & n1010 ;
  assign n1016 = n1015 ^ n1011 ;
  assign n1025 = n888 & n889 ;
  assign n1026 = n275 & n1025 ;
  assign n1033 = ~x43 & ~x129 ;
  assign n1037 = n1026 & n1033 ;
  assign n1017 = n246 & n968 ;
  assign n1018 = n275 & n1017 ;
  assign n1019 = ~n253 & ~n259 ;
  assign n1020 = ~x2 & ~x45 ;
  assign n1021 = n249 & n1020 ;
  assign n1022 = n1019 & n1021 ;
  assign n1023 = n1018 & n1022 ;
  assign n1024 = n1023 ^ x82 ;
  assign n1027 = x77 & ~n262 ;
  assign n1034 = n1027 & n1033 ;
  assign n1035 = n1026 & n1034 ;
  assign n1036 = ~n1024 & n1035 ;
  assign n1038 = n1037 ^ n1036 ;
  assign n1031 = ~x129 & ~n1026 ;
  assign n1028 = ~x129 & n1027 ;
  assign n1029 = ~n1026 & n1028 ;
  assign n1030 = ~n1024 & n1029 ;
  assign n1032 = n1031 ^ n1030 ;
  assign n1039 = n1038 ^ n1032 ;
  assign n1040 = ~n1016 & n1039 ;
  assign n1041 = ~x67 & ~n262 ;
  assign n1042 = x44 & n262 ;
  assign n1043 = ~n1041 & ~n1042 ;
  assign n1044 = ~x129 & ~n962 ;
  assign n1048 = x82 & n889 ;
  assign n1049 = n1044 & n1048 ;
  assign n1050 = n1043 & n1049 ;
  assign n1051 = n929 & n1050 ;
  assign n1045 = ~x82 & n1044 ;
  assign n1046 = n1043 & n1045 ;
  assign n1047 = n1046 ^ n1044 ;
  assign n1052 = n1051 ^ n1047 ;
  assign n1053 = ~x50 & n510 ;
  assign n1054 = x82 & n274 ;
  assign n1055 = n448 & n1054 ;
  assign n1056 = n1053 & n1055 ;
  assign n1057 = n1056 ^ x82 ;
  assign n1058 = n262 & n455 ;
  assign n1059 = ~n259 & n520 ;
  assign n1060 = n1058 & n1059 ;
  assign n1061 = n1060 ^ n411 ;
  assign n1062 = ~x45 & ~n1061 ;
  assign n1063 = ~n1057 & n1062 ;
  assign n1064 = n1063 ^ x45 ;
  assign n1065 = ~x15 & ~n259 ;
  assign n1066 = n249 & n455 ;
  assign n1067 = n1065 & n1066 ;
  assign n1068 = n248 & n1067 ;
  assign n1069 = x68 & ~n262 ;
  assign n1070 = x82 & n1069 ;
  assign n1071 = ~n1068 & n1070 ;
  assign n1072 = n1071 ^ n1069 ;
  assign n1073 = n274 & n448 ;
  assign n1074 = x45 & x82 ;
  assign n1075 = ~x50 & ~x129 ;
  assign n1076 = n1074 & n1075 ;
  assign n1077 = n510 & n1076 ;
  assign n1078 = n1073 & n1077 ;
  assign n1079 = n1078 ^ x129 ;
  assign n1080 = ~n1072 & ~n1079 ;
  assign n1081 = n1064 & n1080 ;
  assign n1082 = ~n245 & n249 ;
  assign n1090 = x82 & n1082 ;
  assign n1091 = ~n925 & n1090 ;
  assign n1092 = n1091 ^ x82 ;
  assign n1087 = ~x75 & ~x82 ;
  assign n1088 = ~n262 & n1087 ;
  assign n1083 = ~x75 & x82 ;
  assign n1084 = ~n262 & n1083 ;
  assign n1085 = n1082 & n1084 ;
  assign n1086 = ~n925 & n1085 ;
  assign n1089 = n1088 ^ n1086 ;
  assign n1093 = n1092 ^ n1089 ;
  assign n1094 = n511 & n1093 ;
  assign n1096 = ~x75 & n263 ;
  assign n1101 = ~n1094 & ~n1096 ;
  assign n1095 = x82 & n1053 ;
  assign n1097 = x46 & ~n263 ;
  assign n1098 = ~n1096 & n1097 ;
  assign n1099 = ~n1095 & n1098 ;
  assign n1100 = ~n1094 & n1099 ;
  assign n1102 = n1101 ^ n1100 ;
  assign n1103 = ~x129 & ~n1102 ;
  assign n1104 = n248 & n880 ;
  assign n1105 = x82 & ~n1104 ;
  assign n1106 = x64 & ~n262 ;
  assign n1107 = ~n1105 & n1106 ;
  assign n1108 = ~n880 & n942 ;
  assign n1109 = n1108 ^ n262 ;
  assign n1116 = x82 & ~n248 ;
  assign n1117 = n1109 & n1116 ;
  assign n1118 = n1117 ^ n1116 ;
  assign n1119 = n1118 ^ n1109 ;
  assign n1113 = x47 & ~n1109 ;
  assign n1110 = x47 & x82 ;
  assign n1111 = ~n248 & n1110 ;
  assign n1112 = ~n1109 & n1111 ;
  assign n1114 = n1113 ^ n1112 ;
  assign n1115 = n1114 ^ x47 ;
  assign n1120 = n1119 ^ n1115 ;
  assign n1121 = ~x43 & x47 ;
  assign n1122 = n1026 & n1121 ;
  assign n1123 = ~x129 & ~n1122 ;
  assign n1124 = n1120 & n1123 ;
  assign n1125 = n1124 ^ n1123 ;
  assign n1126 = n1107 & n1125 ;
  assign n1127 = n1126 ^ n1125 ;
  assign n1128 = x82 & n866 ;
  assign n1129 = n1053 & n1128 ;
  assign n1130 = n1129 ^ x82 ;
  assign n1132 = ~x45 & x82 ;
  assign n1133 = ~n259 & n1132 ;
  assign n1134 = ~n559 & n1133 ;
  assign n1135 = n1134 ^ x82 ;
  assign n1136 = ~x48 & n262 ;
  assign n1137 = ~n1135 & n1136 ;
  assign n1138 = ~n1130 & n1137 ;
  assign n1131 = ~x48 & n1130 ;
  assign n1139 = n1138 ^ n1131 ;
  assign n1140 = x48 & n276 ;
  assign n1141 = n1026 & n1140 ;
  assign n1142 = ~x129 & ~n1141 ;
  assign n1143 = ~n1139 & n1142 ;
  assign n1146 = ~x47 & n248 ;
  assign n1147 = ~n925 & n1146 ;
  assign n1144 = x62 & ~n262 ;
  assign n1148 = x82 & n1144 ;
  assign n1149 = ~n1147 & n1148 ;
  assign n1150 = n1143 & n1149 ;
  assign n1145 = n1143 & ~n1144 ;
  assign n1151 = n1150 ^ n1145 ;
  assign n1152 = n515 & n559 ;
  assign n1153 = ~x46 & n240 ;
  assign n1154 = ~x24 & ~x40 ;
  assign n1155 = n246 & n1154 ;
  assign n1156 = n1153 & n1155 ;
  assign n1157 = x49 & ~n245 ;
  assign n1158 = n512 & n1157 ;
  assign n1159 = n1156 & n1158 ;
  assign n1160 = n1159 ^ x49 ;
  assign n1161 = x82 & ~n1160 ;
  assign n1162 = ~n1152 & n1161 ;
  assign n1163 = n1162 ^ x82 ;
  assign n1164 = x82 & n508 ;
  assign n1165 = n510 & n1164 ;
  assign n1166 = n514 & n1165 ;
  assign n1167 = n1166 ^ x82 ;
  assign n1168 = x49 & n411 ;
  assign n1169 = ~x69 & ~n262 ;
  assign n1170 = ~n1168 & n1169 ;
  assign n1171 = ~n1167 & n1170 ;
  assign n1172 = n1171 ^ n1168 ;
  assign n1173 = ~x129 & ~n1172 ;
  assign n1174 = ~n1163 & n1173 ;
  assign n1175 = n1174 ^ x129 ;
  assign n1186 = x82 & ~n510 ;
  assign n1190 = ~x50 & ~n262 ;
  assign n1191 = ~n1186 & n1190 ;
  assign n1179 = n278 ^ n274 ;
  assign n1180 = ~n278 & n1179 ;
  assign n1181 = n1180 ^ n274 ;
  assign n1182 = n1181 ^ n273 ;
  assign n1183 = n273 & ~n1182 ;
  assign n1184 = n1183 ^ n1180 ;
  assign n1185 = n1184 ^ n274 ;
  assign n1187 = ~x50 & n942 ;
  assign n1188 = ~n1186 & n1187 ;
  assign n1189 = ~n1185 & n1188 ;
  assign n1192 = n1191 ^ n1189 ;
  assign n1193 = n1192 ^ x50 ;
  assign n1176 = x82 & ~n882 ;
  assign n1177 = x66 & ~n262 ;
  assign n1178 = ~n1176 & n1177 ;
  assign n1194 = n1193 ^ n1178 ;
  assign n1195 = x50 & x82 ;
  assign n1196 = n510 & n1195 ;
  assign n1197 = ~x129 & ~n1196 ;
  assign n1198 = n1197 ^ n1193 ;
  assign n1199 = ~n1197 & n1198 ;
  assign n1200 = n1199 ^ n1193 ;
  assign n1201 = ~n1194 & ~n1200 ;
  assign n1202 = n1201 ^ n1199 ;
  assign n1203 = n1202 ^ n1178 ;
  assign n1204 = x51 & ~x109 ;
  assign n1205 = ~x106 & ~n904 ;
  assign n1206 = ~n1204 & n1205 ;
  assign n1207 = ~x129 & ~n1206 ;
  assign n1208 = x52 & ~n904 ;
  assign n1209 = ~x106 & ~n902 ;
  assign n1210 = ~n1208 & n1209 ;
  assign n1211 = ~x129 & ~n1210 ;
  assign n1212 = ~x116 & n786 ;
  assign n1213 = ~x53 & x97 ;
  assign n1214 = x58 & x116 ;
  assign n1215 = ~x58 & n645 ;
  assign n1216 = n772 & n1215 ;
  assign n1217 = ~n1214 & ~n1216 ;
  assign n1218 = n1213 & ~n1217 ;
  assign n1219 = ~n1212 & ~n1218 ;
  assign n1220 = n632 & n703 ;
  assign n1221 = ~n1219 & n1220 ;
  assign n1222 = ~x129 & ~n263 ;
  assign n1223 = n455 & n1065 ;
  assign n1224 = ~n262 & n1223 ;
  assign n1225 = n564 & n1224 ;
  assign n1226 = n1222 & ~n1225 ;
  assign n1227 = ~x123 & ~x129 ;
  assign n1228 = x114 & ~x122 ;
  assign n1229 = n1227 & n1228 ;
  assign n1230 = ~x26 & x37 ;
  assign n1233 = n800 & n1230 ;
  assign n1231 = n631 & n1230 ;
  assign n1236 = n1233 ^ n1231 ;
  assign n1272 = n1236 ^ x27 ;
  assign n1244 = x116 ^ x58 ;
  assign n1242 = x116 ^ x26 ;
  assign n1243 = n1242 ^ x37 ;
  assign n1245 = n1244 ^ n1243 ;
  assign n1246 = n1245 ^ x37 ;
  assign n1248 = n1246 ^ n1244 ;
  assign n1240 = x116 ^ x94 ;
  assign n1241 = n1240 ^ x116 ;
  assign n1249 = n1248 ^ n1241 ;
  assign n1247 = n1246 ^ n1241 ;
  assign n1250 = n1249 ^ n1247 ;
  assign n1253 = ~n1241 & ~n1249 ;
  assign n1251 = n1246 ^ x37 ;
  assign n1252 = ~x116 & n1251 ;
  assign n1254 = n1253 ^ n1252 ;
  assign n1255 = ~n1250 & n1254 ;
  assign n1256 = n1255 ^ n1253 ;
  assign n1257 = n1256 ^ n1246 ;
  assign n1258 = n1257 ^ x116 ;
  assign n1259 = n1258 ^ x116 ;
  assign n1260 = x53 & ~n1259 ;
  assign n1261 = n1260 ^ x53 ;
  assign n1262 = n1261 ^ n1259 ;
  assign n1263 = ~x58 & n1230 ;
  assign n1264 = n1262 & n1263 ;
  assign n1265 = n1264 ^ n1262 ;
  assign n1266 = n1265 ^ n1263 ;
  assign n1237 = n1233 ^ x85 ;
  assign n1238 = n1236 & n1237 ;
  assign n1239 = n1238 ^ x85 ;
  assign n1267 = n1266 ^ n1239 ;
  assign n1273 = n1272 ^ n1267 ;
  assign n1274 = n1266 ^ n1231 ;
  assign n1275 = n1274 ^ n1239 ;
  assign n1276 = n1273 & n1275 ;
  assign n1268 = n1239 ^ n1231 ;
  assign n1234 = n1233 ^ x27 ;
  assign n1269 = n1268 ^ n1234 ;
  assign n1270 = ~n1267 & n1269 ;
  assign n1277 = n1276 ^ n1270 ;
  assign n1278 = n1277 ^ n1239 ;
  assign n1279 = n1278 ^ n1272 ;
  assign n1280 = n1270 ^ n1266 ;
  assign n1281 = n1280 ^ x27 ;
  assign n1282 = n1279 & ~n1281 ;
  assign n1283 = n1282 ^ n1276 ;
  assign n1271 = n1270 ^ n1238 ;
  assign n1284 = n1283 ^ n1271 ;
  assign n1232 = n1231 ^ x85 ;
  assign n1235 = n1234 ^ n1232 ;
  assign n1285 = n1284 ^ n1235 ;
  assign n1286 = n1285 ^ n1233 ;
  assign n1287 = n202 & ~n1286 ;
  assign n1288 = n1287 ^ n202 ;
  assign n1297 = x85 & n631 ;
  assign n1294 = x26 & ~x53 ;
  assign n1295 = ~x58 & n1294 ;
  assign n1292 = ~x26 & ~x58 ;
  assign n1293 = ~x85 & n1292 ;
  assign n1296 = n1295 ^ n1293 ;
  assign n1298 = n1297 ^ n1296 ;
  assign n1307 = x57 & ~n707 ;
  assign n1308 = n1298 & n1307 ;
  assign n1309 = n1308 ^ n707 ;
  assign n1301 = x60 & n1214 ;
  assign n1304 = ~x57 & n707 ;
  assign n1305 = ~n1301 & n1304 ;
  assign n1299 = x57 & x116 ;
  assign n1300 = ~n1298 & n1299 ;
  assign n1302 = n707 & ~n1301 ;
  assign n1303 = n1300 & n1302 ;
  assign n1306 = n1305 ^ n1303 ;
  assign n1310 = n1309 ^ n1306 ;
  assign n1289 = x57 & ~x58 ;
  assign n1290 = n707 & n1289 ;
  assign n1311 = ~x27 & n202 ;
  assign n1312 = ~n1290 & n1311 ;
  assign n1313 = n1310 & n1312 ;
  assign n1291 = n202 & n1290 ;
  assign n1314 = n1313 ^ n1291 ;
  assign n1315 = x58 & ~x116 ;
  assign n1316 = n744 & n1315 ;
  assign n1317 = ~x58 & n738 ;
  assign n1318 = n613 & n1317 ;
  assign n1319 = ~n1316 & ~n1318 ;
  assign n1320 = n202 & n752 ;
  assign n1321 = ~n1319 & n1320 ;
  assign n1322 = x59 & ~x116 ;
  assign n1338 = x27 & n1322 ;
  assign n1339 = n800 & n1338 ;
  assign n1329 = x96 & n631 ;
  assign n1330 = ~n648 & n1329 ;
  assign n1327 = x59 & n631 ;
  assign n1328 = n648 & n1327 ;
  assign n1331 = n1330 ^ n1328 ;
  assign n1332 = n638 & n1322 ;
  assign n1333 = ~x85 & ~n1332 ;
  assign n1334 = ~n1331 & n1333 ;
  assign n1325 = n1297 & n1322 ;
  assign n1326 = n1325 ^ x85 ;
  assign n1335 = n1334 ^ n1326 ;
  assign n1336 = n744 & ~n1335 ;
  assign n1323 = x26 & n1322 ;
  assign n1324 = n800 & n1323 ;
  assign n1337 = n1336 ^ n1324 ;
  assign n1340 = n1339 ^ n1337 ;
  assign n1341 = n202 & n1340 ;
  assign n1342 = ~x117 & ~x122 ;
  assign n1343 = x60 & ~n1342 ;
  assign n1344 = x123 & n1342 ;
  assign n1345 = ~n1343 & ~n1344 ;
  assign n1346 = ~x114 & ~x122 ;
  assign n1347 = x123 & ~x129 ;
  assign n1348 = n1346 & n1347 ;
  assign n1349 = x136 & ~x137 ;
  assign n1350 = x131 & x132 ;
  assign n1351 = x133 & n1350 ;
  assign n1352 = ~x138 & n1351 ;
  assign n1353 = n1349 & n1352 ;
  assign n1354 = x140 & n1353 ;
  assign n1355 = ~x62 & ~n1353 ;
  assign n1356 = ~x129 & ~n1355 ;
  assign n1357 = ~n1354 & n1356 ;
  assign n1358 = x142 & n1353 ;
  assign n1359 = ~x63 & ~n1353 ;
  assign n1360 = ~x129 & ~n1359 ;
  assign n1361 = ~n1358 & n1360 ;
  assign n1362 = x139 & n1353 ;
  assign n1363 = ~x64 & ~n1353 ;
  assign n1364 = ~x129 & ~n1363 ;
  assign n1365 = ~n1362 & n1364 ;
  assign n1366 = x146 & n1353 ;
  assign n1367 = ~x65 & ~n1353 ;
  assign n1368 = ~x129 & ~n1367 ;
  assign n1369 = ~n1366 & n1368 ;
  assign n1370 = ~x136 & ~x137 ;
  assign n1371 = n1352 & n1370 ;
  assign n1372 = x143 & n1371 ;
  assign n1373 = ~x66 & ~n1371 ;
  assign n1374 = ~x129 & ~n1373 ;
  assign n1375 = ~n1372 & n1374 ;
  assign n1376 = x139 & n1371 ;
  assign n1377 = ~x67 & ~n1371 ;
  assign n1378 = ~x129 & ~n1377 ;
  assign n1379 = ~n1376 & n1378 ;
  assign n1380 = x141 & n1353 ;
  assign n1381 = ~x68 & ~n1353 ;
  assign n1382 = ~x129 & ~n1381 ;
  assign n1383 = ~n1380 & n1382 ;
  assign n1384 = x143 & n1353 ;
  assign n1385 = ~x69 & ~n1353 ;
  assign n1386 = ~x129 & ~n1385 ;
  assign n1387 = ~n1384 & n1386 ;
  assign n1388 = x144 & n1353 ;
  assign n1389 = ~x70 & ~n1353 ;
  assign n1390 = ~x129 & ~n1389 ;
  assign n1391 = ~n1388 & n1390 ;
  assign n1392 = x145 & n1353 ;
  assign n1393 = ~x71 & ~n1353 ;
  assign n1394 = ~x129 & ~n1393 ;
  assign n1395 = ~n1392 & n1394 ;
  assign n1396 = x140 & n1371 ;
  assign n1397 = ~x72 & ~n1371 ;
  assign n1398 = ~x129 & ~n1397 ;
  assign n1399 = ~n1396 & n1398 ;
  assign n1400 = x141 & n1371 ;
  assign n1401 = ~x73 & ~n1371 ;
  assign n1402 = ~x129 & ~n1401 ;
  assign n1403 = ~n1400 & n1402 ;
  assign n1404 = x142 & n1371 ;
  assign n1405 = ~x74 & ~n1371 ;
  assign n1406 = ~x129 & ~n1405 ;
  assign n1407 = ~n1404 & n1406 ;
  assign n1408 = x144 & n1371 ;
  assign n1409 = ~x75 & ~n1371 ;
  assign n1410 = ~x129 & ~n1409 ;
  assign n1411 = ~n1408 & n1410 ;
  assign n1412 = x145 & n1371 ;
  assign n1413 = ~x76 & ~n1371 ;
  assign n1414 = ~x129 & ~n1413 ;
  assign n1415 = ~n1412 & n1414 ;
  assign n1416 = x146 & n1371 ;
  assign n1417 = ~x77 & ~n1371 ;
  assign n1418 = ~x129 & ~n1417 ;
  assign n1419 = ~n1416 & n1418 ;
  assign n1420 = ~x136 & x137 ;
  assign n1421 = n1352 & n1420 ;
  assign n1422 = ~x142 & n1421 ;
  assign n1423 = ~x78 & ~n1421 ;
  assign n1424 = ~x129 & ~n1423 ;
  assign n1425 = ~n1422 & n1424 ;
  assign n1426 = ~x143 & n1421 ;
  assign n1427 = ~x79 & ~n1421 ;
  assign n1428 = ~x129 & ~n1427 ;
  assign n1429 = ~n1426 & n1428 ;
  assign n1430 = ~x144 & n1421 ;
  assign n1431 = ~x80 & ~n1421 ;
  assign n1432 = ~x129 & ~n1431 ;
  assign n1433 = ~n1430 & n1432 ;
  assign n1434 = ~x145 & n1421 ;
  assign n1435 = ~x81 & ~n1421 ;
  assign n1436 = ~x129 & ~n1435 ;
  assign n1437 = ~n1434 & n1436 ;
  assign n1438 = ~x146 & n1421 ;
  assign n1439 = ~x82 & ~n1421 ;
  assign n1440 = ~x129 & ~n1439 ;
  assign n1441 = ~n1438 & n1440 ;
  assign n1442 = x136 & ~x138 ;
  assign n1443 = x31 & n1442 ;
  assign n1444 = x115 & x138 ;
  assign n1445 = ~x87 & ~x138 ;
  assign n1446 = ~x136 & ~n1445 ;
  assign n1447 = ~n1444 & n1446 ;
  assign n1448 = ~n1443 & ~n1447 ;
  assign n1449 = x137 & ~n1448 ;
  assign n1450 = x62 & ~x138 ;
  assign n1451 = ~x89 & x138 ;
  assign n1452 = x136 & ~n1451 ;
  assign n1453 = ~n1450 & n1452 ;
  assign n1454 = x72 & ~x138 ;
  assign n1455 = ~x119 & x138 ;
  assign n1456 = ~x136 & ~n1455 ;
  assign n1457 = ~n1454 & n1456 ;
  assign n1458 = ~n1453 & ~n1457 ;
  assign n1459 = ~x137 & ~n1458 ;
  assign n1460 = ~n1449 & ~n1459 ;
  assign n1461 = ~x141 & n1421 ;
  assign n1462 = ~x84 & ~n1421 ;
  assign n1463 = ~x129 & ~n1462 ;
  assign n1464 = ~n1461 & n1463 ;
  assign n1465 = ~x97 & n645 ;
  assign n1466 = ~n696 & ~n1465 ;
  assign n1467 = x96 & n1466 ;
  assign n1468 = ~n588 & ~n1467 ;
  assign n1469 = n686 & n703 ;
  assign n1470 = ~n1468 & n1469 ;
  assign n1471 = ~x139 & n1421 ;
  assign n1472 = ~x86 & ~n1421 ;
  assign n1473 = ~x129 & ~n1472 ;
  assign n1474 = ~n1471 & n1473 ;
  assign n1475 = ~x140 & n1421 ;
  assign n1476 = ~x87 & ~n1421 ;
  assign n1477 = ~x129 & ~n1476 ;
  assign n1478 = ~n1475 & n1477 ;
  assign n1479 = x137 & n1442 ;
  assign n1480 = n1351 & n1479 ;
  assign n1481 = ~x139 & n1480 ;
  assign n1482 = ~x88 & ~n1480 ;
  assign n1483 = ~x129 & ~n1482 ;
  assign n1484 = ~n1481 & n1483 ;
  assign n1485 = ~x140 & n1480 ;
  assign n1486 = ~x89 & ~n1480 ;
  assign n1487 = ~x129 & ~n1486 ;
  assign n1488 = ~n1485 & n1487 ;
  assign n1489 = ~x142 & n1480 ;
  assign n1490 = ~x90 & ~n1480 ;
  assign n1491 = ~x129 & ~n1490 ;
  assign n1492 = ~n1489 & n1491 ;
  assign n1493 = ~x143 & n1480 ;
  assign n1494 = ~x91 & ~n1480 ;
  assign n1495 = ~x129 & ~n1494 ;
  assign n1496 = ~n1493 & n1495 ;
  assign n1497 = ~x144 & n1480 ;
  assign n1498 = ~x92 & ~n1480 ;
  assign n1499 = ~x129 & ~n1498 ;
  assign n1500 = ~n1497 & n1499 ;
  assign n1501 = ~x146 & n1480 ;
  assign n1502 = ~x93 & ~n1480 ;
  assign n1503 = ~x129 & ~n1502 ;
  assign n1504 = ~n1501 & n1503 ;
  assign n1505 = x82 & x138 ;
  assign n1506 = n1370 & n1505 ;
  assign n1507 = n1351 & n1506 ;
  assign n1508 = ~x142 & n1507 ;
  assign n1509 = ~x94 & ~n1507 ;
  assign n1510 = ~x129 & ~n1509 ;
  assign n1511 = ~n1508 & n1510 ;
  assign n1512 = ~x3 & ~x110 ;
  assign n1513 = ~n1351 & ~n1512 ;
  assign n1514 = ~n1507 & ~n1513 ;
  assign n1515 = x95 & n1514 ;
  assign n1516 = x143 & n1507 ;
  assign n1517 = ~n1515 & ~n1516 ;
  assign n1518 = ~x129 & ~n1517 ;
  assign n1519 = x96 & n1514 ;
  assign n1520 = x146 & n1507 ;
  assign n1521 = ~n1519 & ~n1520 ;
  assign n1522 = ~x129 & ~n1521 ;
  assign n1523 = x97 & n1514 ;
  assign n1524 = x145 & n1507 ;
  assign n1525 = ~n1523 & ~n1524 ;
  assign n1526 = ~x129 & ~n1525 ;
  assign n1527 = ~x145 & n1480 ;
  assign n1528 = ~x98 & ~n1480 ;
  assign n1529 = ~x129 & ~n1528 ;
  assign n1530 = ~n1527 & n1529 ;
  assign n1531 = ~x141 & n1480 ;
  assign n1532 = ~x99 & ~n1480 ;
  assign n1533 = ~x129 & ~n1532 ;
  assign n1534 = ~n1531 & n1533 ;
  assign n1535 = x100 & n1514 ;
  assign n1536 = x144 & n1507 ;
  assign n1537 = ~n1535 & ~n1536 ;
  assign n1538 = ~x129 & ~n1537 ;
  assign n1539 = x37 & n1442 ;
  assign n1540 = ~x96 & x138 ;
  assign n1541 = ~x82 & ~x138 ;
  assign n1542 = ~x136 & ~n1541 ;
  assign n1543 = ~n1540 & n1542 ;
  assign n1544 = ~n1539 & ~n1543 ;
  assign n1545 = x137 & ~n1544 ;
  assign n1546 = x65 & ~x138 ;
  assign n1547 = ~x93 & x138 ;
  assign n1548 = x136 & ~n1547 ;
  assign n1549 = ~n1546 & n1548 ;
  assign n1550 = x77 & ~x138 ;
  assign n1551 = ~x124 & x138 ;
  assign n1552 = ~x136 & ~n1551 ;
  assign n1553 = ~n1550 & n1552 ;
  assign n1554 = ~n1549 & ~n1553 ;
  assign n1555 = ~x137 & ~n1554 ;
  assign n1556 = ~n1545 & ~n1555 ;
  assign n1557 = x91 & n1349 ;
  assign n1558 = x95 & n1420 ;
  assign n1559 = ~n1557 & ~n1558 ;
  assign n1560 = x138 & ~n1559 ;
  assign n1561 = ~x34 & x136 ;
  assign n1562 = ~x79 & ~x136 ;
  assign n1563 = x137 & ~n1562 ;
  assign n1564 = ~n1561 & n1563 ;
  assign n1565 = x69 & x136 ;
  assign n1566 = x66 & ~x136 ;
  assign n1567 = ~x137 & ~n1566 ;
  assign n1568 = ~n1565 & n1567 ;
  assign n1569 = ~n1564 & ~n1568 ;
  assign n1570 = ~x138 & ~n1569 ;
  assign n1571 = ~n1560 & ~n1570 ;
  assign n1572 = x90 & n1349 ;
  assign n1573 = x94 & n1420 ;
  assign n1574 = ~n1572 & ~n1573 ;
  assign n1575 = x138 & ~n1574 ;
  assign n1576 = ~x33 & x136 ;
  assign n1577 = ~x78 & ~x136 ;
  assign n1578 = x137 & ~n1577 ;
  assign n1579 = ~n1576 & n1578 ;
  assign n1580 = x63 & x136 ;
  assign n1581 = x74 & ~x136 ;
  assign n1582 = ~x137 & ~n1581 ;
  assign n1583 = ~n1580 & n1582 ;
  assign n1584 = ~n1579 & ~n1583 ;
  assign n1585 = ~x138 & ~n1584 ;
  assign n1586 = ~n1575 & ~n1585 ;
  assign n1587 = x99 & n1349 ;
  assign n1588 = ~x112 & n1420 ;
  assign n1589 = ~n1587 & ~n1588 ;
  assign n1590 = x138 & ~n1589 ;
  assign n1591 = ~x32 & x136 ;
  assign n1592 = ~x84 & ~x136 ;
  assign n1593 = x137 & ~n1592 ;
  assign n1594 = ~n1591 & n1593 ;
  assign n1595 = x68 & x136 ;
  assign n1596 = x73 & ~x136 ;
  assign n1597 = ~x137 & ~n1596 ;
  assign n1598 = ~n1595 & n1597 ;
  assign n1599 = ~n1594 & ~n1598 ;
  assign n1600 = ~x138 & ~n1599 ;
  assign n1601 = ~n1590 & ~n1600 ;
  assign n1602 = x35 & n1442 ;
  assign n1603 = ~x100 & x138 ;
  assign n1604 = ~x80 & ~x138 ;
  assign n1605 = ~x136 & ~n1604 ;
  assign n1606 = ~n1603 & n1605 ;
  assign n1607 = ~n1602 & ~n1606 ;
  assign n1608 = x137 & ~n1607 ;
  assign n1609 = x70 & ~x138 ;
  assign n1610 = ~x92 & x138 ;
  assign n1611 = x136 & ~n1610 ;
  assign n1612 = ~n1609 & n1611 ;
  assign n1613 = x75 & ~x138 ;
  assign n1614 = ~x125 & x138 ;
  assign n1615 = ~x136 & ~n1614 ;
  assign n1616 = ~n1613 & n1615 ;
  assign n1617 = ~n1612 & ~n1616 ;
  assign n1618 = ~x137 & ~n1617 ;
  assign n1619 = ~n1608 & ~n1618 ;
  assign n1620 = ~x26 & n686 ;
  assign n1621 = n1466 & n1620 ;
  assign n1622 = ~n693 & ~n1621 ;
  assign n1623 = n202 & ~n1622 ;
  assign n1624 = x36 & n1442 ;
  assign n1625 = ~x97 & x138 ;
  assign n1626 = ~x81 & ~x138 ;
  assign n1627 = ~x136 & ~n1626 ;
  assign n1628 = ~n1625 & n1627 ;
  assign n1629 = ~n1624 & ~n1628 ;
  assign n1630 = x137 & ~n1629 ;
  assign n1631 = x71 & ~x138 ;
  assign n1632 = ~x98 & x138 ;
  assign n1633 = x136 & ~n1632 ;
  assign n1634 = ~n1631 & n1633 ;
  assign n1635 = x76 & ~x138 ;
  assign n1636 = ~x23 & x138 ;
  assign n1637 = ~x136 & ~n1636 ;
  assign n1638 = ~n1635 & n1637 ;
  assign n1639 = ~n1634 & ~n1638 ;
  assign n1640 = ~x137 & ~n1639 ;
  assign n1641 = ~n1630 & ~n1640 ;
  assign n1642 = x30 & n1442 ;
  assign n1643 = ~x111 & x138 ;
  assign n1644 = ~x86 & ~x138 ;
  assign n1645 = ~x136 & ~n1644 ;
  assign n1646 = ~n1643 & n1645 ;
  assign n1647 = ~n1642 & ~n1646 ;
  assign n1648 = x137 & ~n1647 ;
  assign n1649 = x64 & ~x138 ;
  assign n1650 = ~x88 & x138 ;
  assign n1651 = x136 & ~n1650 ;
  assign n1652 = ~n1649 & n1651 ;
  assign n1653 = x67 & ~x138 ;
  assign n1654 = ~x120 & x138 ;
  assign n1655 = ~x136 & ~n1654 ;
  assign n1656 = ~n1653 & n1655 ;
  assign n1657 = ~n1652 & ~n1656 ;
  assign n1658 = ~x137 & ~n1657 ;
  assign n1659 = ~n1648 & ~n1658 ;
  assign n1660 = ~x26 & n726 ;
  assign n1661 = ~n799 & ~n1660 ;
  assign n1662 = x116 & n202 ;
  assign n1663 = ~n1661 & n1662 ;
  assign n1664 = ~x53 & x58 ;
  assign n1665 = ~x97 & n1664 ;
  assign n1666 = ~n786 & ~n1665 ;
  assign n1667 = n1662 & ~n1666 ;
  assign n1668 = ~x139 & n1506 ;
  assign n1669 = ~x129 & n1351 ;
  assign n1670 = ~x111 & ~n1506 ;
  assign n1671 = n1669 & ~n1670 ;
  assign n1672 = ~n1668 & n1671 ;
  assign n1673 = x112 & ~n1506 ;
  assign n1674 = ~x141 & n1506 ;
  assign n1675 = n1669 & ~n1674 ;
  assign n1676 = ~n1673 & n1675 ;
  assign n1677 = ~x11 & ~x22 ;
  assign n1678 = x54 & n1677 ;
  assign n1679 = ~x54 & x113 ;
  assign n1680 = n202 & ~n1679 ;
  assign n1681 = ~n1678 & n1680 ;
  assign n1682 = x115 & ~n1506 ;
  assign n1683 = ~x140 & n1506 ;
  assign n1684 = n1669 & ~n1683 ;
  assign n1685 = ~n1682 & n1684 ;
  assign n1686 = x54 & n202 ;
  assign n1687 = ~x4 & ~x9 ;
  assign n1688 = n205 & n1687 ;
  assign n1689 = n1686 & ~n1688 ;
  assign n1690 = x122 & ~x129 ;
  assign n1691 = ~x54 & x118 ;
  assign n1692 = x54 & ~x59 ;
  assign n1693 = n391 & n1692 ;
  assign n1694 = ~n1691 & ~n1693 ;
  assign n1695 = ~x129 & ~n1694 ;
  assign n1696 = ~x129 & ~n645 ;
  assign n1697 = ~x120 & n1512 ;
  assign n1698 = ~x111 & ~x129 ;
  assign n1699 = ~n1697 & n1698 ;
  assign n1700 = x81 & x120 ;
  assign n1701 = ~x129 & n1700 ;
  assign n1702 = ~x129 & ~x134 ;
  assign n1703 = ~x129 & ~x135 ;
  assign n1704 = x57 & ~x129 ;
  assign n1705 = ~x96 & x125 ;
  assign n1706 = ~x3 & ~n1705 ;
  assign n1707 = ~x129 & ~n1706 ;
  assign n1708 = ~x126 & x132 ;
  assign n1709 = x133 & n1708 ;
  assign y0 = x108 ;
  assign y1 = x83 ;
  assign y2 = x104 ;
  assign y3 = x103 ;
  assign y4 = x102 ;
  assign y5 = x105 ;
  assign y6 = x107 ;
  assign y7 = x101 ;
  assign y8 = x126 ;
  assign y9 = x121 ;
  assign y10 = x1 ;
  assign y11 = x0 ;
  assign y12 = ~1'b0 ;
  assign y13 = x130 ;
  assign y14 = x128 ;
  assign y15 = ~n203 ;
  assign y16 = ~n239 ;
  assign y17 = n287 ;
  assign y18 = ~n302 ;
  assign y19 = n317 ;
  assign y20 = n330 ;
  assign y21 = n338 ;
  assign y22 = n345 ;
  assign y23 = n356 ;
  assign y24 = n363 ;
  assign y25 = n373 ;
  assign y26 = n382 ;
  assign y27 = n389 ;
  assign y28 = n400 ;
  assign y29 = n408 ;
  assign y30 = ~n471 ;
  assign y31 = n479 ;
  assign y32 = n488 ;
  assign y33 = n498 ;
  assign y34 = n507 ;
  assign y35 = n536 ;
  assign y36 = n544 ;
  assign y37 = n553 ;
  assign y38 = n556 ;
  assign y39 = n587 ;
  assign y40 = ~n681 ;
  assign y41 = n688 ;
  assign y42 = n705 ;
  assign y43 = n764 ;
  assign y44 = n805 ;
  assign y45 = n812 ;
  assign y46 = n819 ;
  assign y47 = n826 ;
  assign y48 = n833 ;
  assign y49 = n840 ;
  assign y50 = n847 ;
  assign y51 = n854 ;
  assign y52 = n861 ;
  assign y53 = ~n901 ;
  assign y54 = n908 ;
  assign y55 = n934 ;
  assign y56 = n960 ;
  assign y57 = n1005 ;
  assign y58 = n1040 ;
  assign y59 = n1052 ;
  assign y60 = n1081 ;
  assign y61 = n1103 ;
  assign y62 = n1127 ;
  assign y63 = n1151 ;
  assign y64 = ~n1175 ;
  assign y65 = ~n1203 ;
  assign y66 = n1207 ;
  assign y67 = n1211 ;
  assign y68 = n1221 ;
  assign y69 = ~n1226 ;
  assign y70 = n1229 ;
  assign y71 = n1288 ;
  assign y72 = n1314 ;
  assign y73 = n1321 ;
  assign y74 = n1341 ;
  assign y75 = ~n1345 ;
  assign y76 = n1348 ;
  assign y77 = ~n1357 ;
  assign y78 = ~n1361 ;
  assign y79 = ~n1365 ;
  assign y80 = ~n1369 ;
  assign y81 = ~n1375 ;
  assign y82 = ~n1379 ;
  assign y83 = ~n1383 ;
  assign y84 = ~n1387 ;
  assign y85 = ~n1391 ;
  assign y86 = ~n1395 ;
  assign y87 = ~n1399 ;
  assign y88 = ~n1403 ;
  assign y89 = ~n1407 ;
  assign y90 = ~n1411 ;
  assign y91 = ~n1415 ;
  assign y92 = ~n1419 ;
  assign y93 = n1425 ;
  assign y94 = n1429 ;
  assign y95 = n1433 ;
  assign y96 = n1437 ;
  assign y97 = n1441 ;
  assign y98 = ~n1460 ;
  assign y99 = n1464 ;
  assign y100 = n1470 ;
  assign y101 = n1474 ;
  assign y102 = n1478 ;
  assign y103 = n1484 ;
  assign y104 = n1488 ;
  assign y105 = n1492 ;
  assign y106 = n1496 ;
  assign y107 = n1500 ;
  assign y108 = n1504 ;
  assign y109 = n1511 ;
  assign y110 = n1518 ;
  assign y111 = n1522 ;
  assign y112 = n1526 ;
  assign y113 = n1530 ;
  assign y114 = n1534 ;
  assign y115 = n1538 ;
  assign y116 = ~n1556 ;
  assign y117 = ~n1571 ;
  assign y118 = ~n1586 ;
  assign y119 = ~n1601 ;
  assign y120 = ~n1619 ;
  assign y121 = n1623 ;
  assign y122 = ~n1641 ;
  assign y123 = ~n1659 ;
  assign y124 = n1663 ;
  assign y125 = n1667 ;
  assign y126 = n1672 ;
  assign y127 = n1676 ;
  assign y128 = n1681 ;
  assign y129 = ~n1227 ;
  assign y130 = n1685 ;
  assign y131 = n1689 ;
  assign y132 = ~n1690 ;
  assign y133 = n1695 ;
  assign y134 = n1696 ;
  assign y135 = n1699 ;
  assign y136 = n1701 ;
  assign y137 = ~n1702 ;
  assign y138 = ~n1703 ;
  assign y139 = n1704 ;
  assign y140 = n1707 ;
  assign y141 = n1709 ;
endmodule
