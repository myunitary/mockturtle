module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 ;
  assign n210 = ~x31 & x63 ;
  assign n138 = x63 ^ x31 ;
  assign n208 = ~x30 & x62 ;
  assign n209 = ~n138 & n208 ;
  assign n211 = n210 ^ n209 ;
  assign n137 = x62 ^ x30 ;
  assign n139 = ~n137 & ~n138 ;
  assign n205 = ~x29 & x61 ;
  assign n141 = x61 ^ x29 ;
  assign n203 = ~x28 & x60 ;
  assign n204 = ~n141 & n203 ;
  assign n206 = n205 ^ n204 ;
  assign n207 = n139 & n206 ;
  assign n212 = n211 ^ n207 ;
  assign n140 = x60 ^ x28 ;
  assign n142 = ~n140 & ~n141 ;
  assign n143 = n139 & n142 ;
  assign n199 = ~x27 & x59 ;
  assign n145 = x59 ^ x27 ;
  assign n197 = ~x26 & x58 ;
  assign n198 = ~n145 & n197 ;
  assign n200 = n199 ^ n198 ;
  assign n144 = x58 ^ x26 ;
  assign n146 = ~n144 & ~n145 ;
  assign n194 = ~x25 & x57 ;
  assign n148 = x57 ^ x25 ;
  assign n192 = ~x24 & x56 ;
  assign n193 = ~n148 & n192 ;
  assign n195 = n194 ^ n193 ;
  assign n196 = n146 & n195 ;
  assign n201 = n200 ^ n196 ;
  assign n202 = n143 & n201 ;
  assign n213 = n212 ^ n202 ;
  assign n147 = x56 ^ x24 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = n146 & n149 ;
  assign n151 = n143 & n150 ;
  assign n187 = ~x23 & x55 ;
  assign n153 = x55 ^ x23 ;
  assign n185 = ~x22 & x54 ;
  assign n186 = ~n153 & n185 ;
  assign n188 = n187 ^ n186 ;
  assign n152 = x54 ^ x22 ;
  assign n154 = ~n152 & ~n153 ;
  assign n182 = ~x21 & x53 ;
  assign n156 = x53 ^ x21 ;
  assign n180 = ~x20 & x52 ;
  assign n181 = ~n156 & n180 ;
  assign n183 = n182 ^ n181 ;
  assign n184 = n154 & n183 ;
  assign n189 = n188 ^ n184 ;
  assign n155 = x52 ^ x20 ;
  assign n157 = ~n155 & ~n156 ;
  assign n158 = n154 & n157 ;
  assign n176 = ~x19 & x51 ;
  assign n160 = x51 ^ x19 ;
  assign n174 = ~x18 & x50 ;
  assign n175 = ~n160 & n174 ;
  assign n177 = n176 ^ n175 ;
  assign n159 = x50 ^ x18 ;
  assign n161 = ~n159 & ~n160 ;
  assign n171 = ~x17 & x49 ;
  assign n163 = x49 ^ x17 ;
  assign n169 = ~x16 & x48 ;
  assign n170 = ~n163 & n169 ;
  assign n172 = n171 ^ n170 ;
  assign n173 = n161 & n172 ;
  assign n178 = n177 ^ n173 ;
  assign n179 = n158 & n178 ;
  assign n190 = n189 ^ n179 ;
  assign n191 = n151 & n190 ;
  assign n214 = n213 ^ n191 ;
  assign n132 = ~x15 & x47 ;
  assign n99 = x47 ^ x15 ;
  assign n130 = ~x14 & x46 ;
  assign n131 = ~n99 & n130 ;
  assign n133 = n132 ^ n131 ;
  assign n98 = x46 ^ x14 ;
  assign n100 = ~n98 & ~n99 ;
  assign n127 = ~x13 & x45 ;
  assign n102 = x45 ^ x13 ;
  assign n125 = ~x12 & x44 ;
  assign n126 = ~n102 & n125 ;
  assign n128 = n127 ^ n126 ;
  assign n129 = n100 & n128 ;
  assign n134 = n133 ^ n129 ;
  assign n101 = x44 ^ x12 ;
  assign n103 = ~n101 & ~n102 ;
  assign n104 = n100 & n103 ;
  assign n121 = ~x11 & x43 ;
  assign n106 = x43 ^ x11 ;
  assign n119 = ~x10 & x42 ;
  assign n120 = ~n106 & n119 ;
  assign n122 = n121 ^ n120 ;
  assign n105 = x42 ^ x10 ;
  assign n107 = ~n105 & ~n106 ;
  assign n116 = ~x9 & x41 ;
  assign n109 = x41 ^ x9 ;
  assign n114 = ~x8 & x40 ;
  assign n115 = ~n109 & n114 ;
  assign n117 = n116 ^ n115 ;
  assign n118 = n107 & n117 ;
  assign n123 = n122 ^ n118 ;
  assign n124 = n104 & n123 ;
  assign n135 = n134 ^ n124 ;
  assign n94 = ~x7 & x39 ;
  assign n80 = x39 ^ x7 ;
  assign n92 = ~x6 & x38 ;
  assign n93 = ~n80 & n92 ;
  assign n95 = n94 ^ n93 ;
  assign n79 = x38 ^ x6 ;
  assign n81 = ~n79 & ~n80 ;
  assign n89 = ~x5 & x37 ;
  assign n83 = x37 ^ x5 ;
  assign n87 = ~x4 & x36 ;
  assign n88 = ~n83 & n87 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = n81 & n90 ;
  assign n96 = n95 ^ n91 ;
  assign n76 = ~x3 & x35 ;
  assign n71 = x35 ^ x3 ;
  assign n74 = ~x2 & x34 ;
  assign n75 = ~n71 & n74 ;
  assign n77 = n76 ^ n75 ;
  assign n68 = ~x1 & x33 ;
  assign n65 = x33 ^ x1 ;
  assign n66 = ~x0 & x32 ;
  assign n67 = ~n65 & n66 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = x34 ^ x2 ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = n69 & n72 ;
  assign n78 = n77 ^ n73 ;
  assign n82 = x36 ^ x4 ;
  assign n84 = ~n82 & ~n83 ;
  assign n85 = n81 & n84 ;
  assign n86 = n78 & n85 ;
  assign n97 = n96 ^ n86 ;
  assign n108 = x40 ^ x8 ;
  assign n110 = ~n108 & ~n109 ;
  assign n111 = n107 & n110 ;
  assign n112 = n104 & n111 ;
  assign n113 = n97 & n112 ;
  assign n136 = n135 ^ n113 ;
  assign n162 = x48 ^ x16 ;
  assign n164 = ~n162 & ~n163 ;
  assign n165 = n161 & n164 ;
  assign n166 = n158 & n165 ;
  assign n167 = n151 & n166 ;
  assign n168 = n136 & n167 ;
  assign n215 = n214 ^ n168 ;
  assign n216 = x32 ^ x0 ;
  assign n217 = n215 & n216 ;
  assign n218 = n217 ^ x32 ;
  assign n219 = n65 & n215 ;
  assign n220 = n219 ^ x33 ;
  assign n221 = n70 & n215 ;
  assign n222 = n221 ^ x34 ;
  assign n223 = n71 & n215 ;
  assign n224 = n223 ^ x35 ;
  assign n225 = n82 & n215 ;
  assign n226 = n225 ^ x36 ;
  assign n227 = n83 & n215 ;
  assign n228 = n227 ^ x37 ;
  assign n229 = n79 & n215 ;
  assign n230 = n229 ^ x38 ;
  assign n231 = n80 & n215 ;
  assign n232 = n231 ^ x39 ;
  assign n233 = n108 & n215 ;
  assign n234 = n233 ^ x40 ;
  assign n235 = n109 & n215 ;
  assign n236 = n235 ^ x41 ;
  assign n237 = n105 & n215 ;
  assign n238 = n237 ^ x42 ;
  assign n239 = n106 & n215 ;
  assign n240 = n239 ^ x43 ;
  assign n241 = n101 & n215 ;
  assign n242 = n241 ^ x44 ;
  assign n243 = n102 & n215 ;
  assign n244 = n243 ^ x45 ;
  assign n245 = n98 & n215 ;
  assign n246 = n245 ^ x46 ;
  assign n247 = n99 & n215 ;
  assign n248 = n247 ^ x47 ;
  assign n249 = n162 & n215 ;
  assign n250 = n249 ^ x48 ;
  assign n251 = n163 & n215 ;
  assign n252 = n251 ^ x49 ;
  assign n253 = n159 & n215 ;
  assign n254 = n253 ^ x50 ;
  assign n255 = n160 & n215 ;
  assign n256 = n255 ^ x51 ;
  assign n257 = n155 & n215 ;
  assign n258 = n257 ^ x52 ;
  assign n259 = n156 & n215 ;
  assign n260 = n259 ^ x53 ;
  assign n261 = n152 & n215 ;
  assign n262 = n261 ^ x54 ;
  assign n263 = n153 & n215 ;
  assign n264 = n263 ^ x55 ;
  assign n265 = n147 & n215 ;
  assign n266 = n265 ^ x56 ;
  assign n267 = n148 & n215 ;
  assign n268 = n267 ^ x57 ;
  assign n269 = n144 & n215 ;
  assign n270 = n269 ^ x58 ;
  assign n271 = n145 & n215 ;
  assign n272 = n271 ^ x59 ;
  assign n273 = n140 & n215 ;
  assign n274 = n273 ^ x60 ;
  assign n275 = n141 & n215 ;
  assign n276 = n275 ^ x61 ;
  assign n277 = n137 & n215 ;
  assign n278 = n277 ^ x62 ;
  assign n279 = n138 & n215 ;
  assign n280 = n279 ^ x63 ;
  assign y0 = n218 ;
  assign y1 = n220 ;
  assign y2 = n222 ;
  assign y3 = n224 ;
  assign y4 = n226 ;
  assign y5 = n228 ;
  assign y6 = n230 ;
  assign y7 = n232 ;
  assign y8 = n234 ;
  assign y9 = n236 ;
  assign y10 = n238 ;
  assign y11 = n240 ;
  assign y12 = n242 ;
  assign y13 = n244 ;
  assign y14 = n246 ;
  assign y15 = n248 ;
  assign y16 = n250 ;
  assign y17 = n252 ;
  assign y18 = n254 ;
  assign y19 = n256 ;
  assign y20 = n258 ;
  assign y21 = n260 ;
  assign y22 = n262 ;
  assign y23 = n264 ;
  assign y24 = n266 ;
  assign y25 = n268 ;
  assign y26 = n270 ;
  assign y27 = n272 ;
  assign y28 = n274 ;
  assign y29 = n276 ;
  assign y30 = n278 ;
  assign y31 = n280 ;
endmodule
