module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 ;
  assign n33 = x12 & x13 ;
  assign n34 = n33 ^ x12 ;
  assign n35 = n34 ^ x13 ;
  assign n36 = x14 & x15 ;
  assign n37 = n36 ^ x14 ;
  assign n38 = n37 ^ x15 ;
  assign n39 = n35 & n38 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = x8 & x9 ;
  assign n43 = n42 ^ x8 ;
  assign n44 = n43 ^ x9 ;
  assign n45 = x10 & x11 ;
  assign n46 = n45 ^ x10 ;
  assign n47 = n46 ^ x11 ;
  assign n48 = n44 & n47 ;
  assign n49 = n48 ^ n44 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = ~n41 & ~n50 ;
  assign n52 = x4 & x5 ;
  assign n53 = n52 ^ x4 ;
  assign n54 = n53 ^ x5 ;
  assign n55 = x6 & x7 ;
  assign n56 = n55 ^ x6 ;
  assign n57 = n56 ^ x7 ;
  assign n58 = n54 & n57 ;
  assign n59 = n58 ^ n54 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = x0 & x1 ;
  assign n62 = n61 ^ x0 ;
  assign n63 = n62 ^ x1 ;
  assign n64 = x2 & x3 ;
  assign n65 = n64 ^ x2 ;
  assign n66 = n65 ^ x3 ;
  assign n67 = n63 & n66 ;
  assign n68 = n67 ^ n63 ;
  assign n69 = n68 ^ n66 ;
  assign n70 = ~n60 & ~n69 ;
  assign n71 = n51 & n70 ;
  assign n72 = n71 ^ n51 ;
  assign n73 = n72 ^ n70 ;
  assign n74 = x28 & x29 ;
  assign n75 = n74 ^ x28 ;
  assign n76 = n75 ^ x29 ;
  assign n77 = x30 & x31 ;
  assign n78 = n77 ^ x30 ;
  assign n79 = n78 ^ x31 ;
  assign n80 = n76 & n79 ;
  assign n81 = n80 ^ n76 ;
  assign n82 = n81 ^ n79 ;
  assign n83 = x24 & x25 ;
  assign n84 = n83 ^ x24 ;
  assign n85 = n84 ^ x25 ;
  assign n86 = x26 & x27 ;
  assign n87 = n86 ^ x26 ;
  assign n88 = n87 ^ x27 ;
  assign n89 = n85 & n88 ;
  assign n90 = n89 ^ n85 ;
  assign n91 = n90 ^ n88 ;
  assign n92 = ~n82 & ~n91 ;
  assign n93 = x20 & x21 ;
  assign n94 = n93 ^ x20 ;
  assign n95 = n94 ^ x21 ;
  assign n96 = x22 & x23 ;
  assign n97 = n96 ^ x22 ;
  assign n98 = n97 ^ x23 ;
  assign n99 = n95 & n98 ;
  assign n100 = n99 ^ n95 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = x16 & x17 ;
  assign n103 = n102 ^ x16 ;
  assign n104 = n103 ^ x17 ;
  assign n105 = x18 & x19 ;
  assign n106 = n105 ^ x18 ;
  assign n107 = n106 ^ x19 ;
  assign n108 = n104 & n107 ;
  assign n109 = n108 ^ n104 ;
  assign n110 = n109 ^ n107 ;
  assign n111 = ~n101 & ~n110 ;
  assign n112 = n92 & n111 ;
  assign n113 = n112 ^ n92 ;
  assign n114 = n113 ^ n111 ;
  assign n115 = n73 & n114 ;
  assign n116 = n115 ^ n73 ;
  assign n117 = n116 ^ n114 ;
  assign n118 = n115 ^ n114 ;
  assign n119 = n73 & n113 ;
  assign n120 = n119 ^ n113 ;
  assign n121 = n120 ^ n73 ;
  assign n122 = n121 ^ n70 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = 1'b0 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = ~n117 ;
  assign y30 = n118 ;
  assign y31 = n122 ;
endmodule
