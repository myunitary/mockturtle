module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23;
output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24;
wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985, n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, n_4012, n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, n_4021, n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4029, n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4048, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, n_4057, n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077, n_4078, n_4079, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085, n_4086, n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, n_4093, n_4094, n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, n_4102, n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157, n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165, n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220, n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, n_4227, n_4228, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, n_4236, n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, n_4255, n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, n_4264, n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281, n_4282, n_4283, n_4284, n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, n_4291, n_4292, n_4293, n_4294, n_4295, n_4296, n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, n_4303, n_4304, n_4305, n_4306, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312, n_4313, n_4314, n_4315, n_4316, n_4317, n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330, n_4331, n_4332, n_4333, n_4334, n_4335, n_4336, n_4337, n_4338, n_4339, n_4340, n_4341, n_4342, n_4343, n_4344, n_4345, n_4346, n_4347, n_4348, n_4349, n_4350, n_4351, n_4352, n_4353, n_4354, n_4355, n_4356, n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, n_4363, n_4364, n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372, n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380, n_4381, n_4382, n_4383, n_4384, n_4385, n_4386, n_4387, n_4388, n_4389, n_4390, n_4391, n_4392, n_4393, n_4394, n_4395, n_4396, n_4397, n_4398, n_4399, n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4407, n_4408, n_4409, n_4410, n_4411, n_4412, n_4413, n_4414, n_4415, n_4416, n_4417, n_4418, n_4419, n_4420, n_4421, n_4422, n_4423, n_4424, n_4425, n_4426, n_4427, n_4428, n_4429, n_4430, n_4431, n_4432, n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439, n_4440, n_4441, n_4442, n_4443, n_4444, n_4445, n_4446, n_4447, n_4448, n_4449, n_4450, n_4451, n_4452, n_4453, n_4454, n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461, n_4462, n_4463, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469, n_4470, n_4471, n_4472, n_4473, n_4474, n_4475, n_4476, n_4477, n_4478, n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485, n_4486, n_4487, n_4488, n_4489, n_4490, n_4491, n_4492, n_4493, n_4494, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500, n_4501, n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509, n_4510, n_4511, n_4512, n_4513, n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525, n_4526, n_4527, n_4528, n_4529, n_4530, n_4531, n_4532, n_4533, n_4534, n_4535, n_4536, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4543, n_4544, n_4545, n_4546, n_4547, n_4548, n_4549, n_4550, n_4551, n_4552, n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559, n_4560, n_4561, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568, n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575, n_4576, n_4577, n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584, n_4585, n_4586, n_4587, n_4588, n_4589, n_4590, n_4591, n_4592, n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600, n_4601, n_4602, n_4603, n_4604, n_4605, n_4606, n_4607, n_4608, n_4609, n_4610, n_4611, n_4612, n_4613, n_4614, n_4615, n_4616, n_4617, n_4618, n_4619, n_4620, n_4621, n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4629, n_4630, n_4631, n_4632, n_4633, n_4634, n_4635, n_4636, n_4637, n_4638, n_4639, n_4640, n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648, n_4649, n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656, n_4657, n_4658, n_4659, n_4660, n_4661, n_4662, n_4663, n_4664, n_4665, n_4666, n_4667, n_4668, n_4669, n_4670, n_4671, n_4672, n_4673, n_4674, n_4675, n_4676, n_4677, n_4678, n_4679, n_4680, n_4681, n_4682, n_4683, n_4684, n_4685, n_4686, n_4687, n_4688, n_4689, n_4690, n_4691, n_4692, n_4693, n_4694, n_4695, n_4696, n_4697, n_4698, n_4699, n_4700, n_4701, n_4702, n_4703, n_4704, n_4705, n_4706, n_4707, n_4708, n_4709, n_4710, n_4711, n_4712, n_4713, n_4714, n_4715, n_4716, n_4717, n_4718, n_4719, n_4720, n_4721, n_4722, n_4723, n_4724, n_4725, n_4726, n_4727, n_4728, n_4729, n_4730, n_4731, n_4732, n_4733, n_4734, n_4735, n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750, n_4751, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4758, n_4759, n_4760, n_4761, n_4762, n_4763, n_4764, n_4765, n_4766, n_4767, n_4768, n_4769, n_4770, n_4771, n_4772, n_4773, n_4774, n_4775, n_4776, n_4777, n_4778, n_4779, n_4780, n_4781, n_4782, n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790, n_4791, n_4792, n_4793, n_4794, n_4795, n_4796, n_4797, n_4798, n_4799, n_4800, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806, n_4807, n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814, n_4815, n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823, n_4824, n_4825, n_4826, n_4827, n_4828, n_4829, n_4830, n_4831, n_4832, n_4833, n_4834, n_4835, n_4836, n_4837, n_4838, n_4839, n_4840, n_4841, n_4842, n_4843, n_4844, n_4845, n_4846, n_4847, n_4848, n_4849, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855, n_4856, n_4857, n_4858, n_4859, n_4860, n_4861, n_4862, n_4863, n_4864, n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872, n_4873, n_4874, n_4875, n_4876, n_4877, n_4878, n_4879, n_4880, n_4881, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887, n_4888, n_4889, n_4890, n_4891, n_4892, n_4893, n_4894, n_4895, n_4896, n_4897, n_4898, n_4899, n_4900, n_4901, n_4902, n_4903, n_4904, n_4905, n_4906, n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913, n_4914, n_4915, n_4916, n_4917, n_4918, n_4919, n_4920, n_4921, n_4922, n_4923, n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930, n_4931, n_4932, n_4933, n_4934, n_4935, n_4936, n_4937, n_4938, n_4939, n_4940, n_4941, n_4942, n_4943, n_4944, n_4945, n_4946, n_4947, n_4948, n_4949, n_4950, y0, n_4951, n_4952, n_4953, n_4954, n_4955, n_4956, n_4957, n_4958, n_4959, n_4960, n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, n_4969, n_4970, n_4971, n_4972, n_4973, n_4974, n_4975, n_4976, n_4977, n_4978, n_4979, n_4980, n_4981, n_4982, n_4983, n_4984, n_4985, n_4986, n_4987, n_4988, n_4989, n_4990, n_4991, n_4992, n_4993, n_4994, n_4995, n_4996, n_4997, n_4998, y1, n_4999, n_5000, n_5001, n_5002, n_5003, n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010, n_5011, n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018, n_5019, n_5020, n_5021, n_5022, n_5023, y2, n_5024, n_5025, n_5026, n_5027, n_5028, n_5029, n_5030, n_5031, n_5032, n_5033, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040, n_5041, n_5042, n_5043, n_5044, n_5045, n_5046, n_5047, n_5048, n_5049, n_5050, n_5051, n_5052, n_5053, n_5054, n_5055, n_5056, n_5057, n_5058, n_5059, n_5060, n_5061, n_5062, n_5063, n_5064, n_5065, n_5066, n_5067, n_5068, n_5069, n_5070, n_5071, n_5072, n_5073, n_5074, n_5075, n_5076, n_5077, n_5078, n_5079, n_5080, n_5081, n_5082, n_5083, n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091, n_5092, n_5093, n_5094, n_5095, n_5096, n_5097, n_5098, n_5099, n_5100, n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107, n_5108, n_5109, y3, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115, n_5116, n_5117, n_5118, n_5119, n_5120, n_5121, n_5122, n_5123, n_5124, n_5125, y4, n_5126, n_5127, n_5128, n_5129, n_5130, n_5131, n_5132, n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139, n_5140, n_5141, n_5142, n_5143, n_5144, y6, n_5145, n_5146, n_5147, n_5148, n_5149, n_5150, n_5151, n_5152, y5, y7, n_5153, n_5154, n_5155, n_5156, n_5157, n_5158, n_5159, n_5160, n_5161, n_5162, n_5163, n_5164, n_5165, n_5166, n_5167, n_5168, n_5169, n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5176, n_5177, n_5178, n_5179, n_5180, y8, n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192, n_5193, n_5194, y9, n_5195, n_5196, n_5197, n_5198, n_5199, n_5200, n_5201, n_5202, n_5203, n_5204, n_5205, y10, n_5206, n_5207, n_5208, n_5209, y11, n_5210, n_5211, n_5212, n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, y12, n_5219, n_5220, n_5221, n_5222, n_5223, n_5224, n_5225, n_5226, n_5227, y13, n_5228, n_5229, n_5230, n_5231, n_5232, n_5233, n_5234, n_5235, n_5236, y14, n_5237, n_5238, n_5239, n_5240, n_5241, n_5242, n_5243, n_5244, n_5245, y15, n_5246, n_5247, n_5248, n_5249, n_5250, n_5251, n_5252, n_5253, n_5254, y16, n_5255, n_5256, n_5257, n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, y17, n_5264, n_5265, n_5266, n_5267, n_5268, n_5269, n_5270, n_5271, n_5272, n_5273, n_5274, n_5275, n_5276, n_5277, n_5278, n_5279, n_5280, n_5281, n_5282, n_5283, n_5284, n_5285, n_5286, n_5287, n_5288, n_5289, n_5290, y18, n_5291, n_5292, n_5293, y19, n_5294, n_5295, n_5296, n_5297, n_5298, n_5299, n_5300, n_5301, n_5302, n_5303, n_5304, n_5305, n_5306, y22, y24, n_5307, y21, n_5308, y20, y23;
assign n_0 = ~x0 & x1;
assign n_1 = x2 ^ x1;
assign n_2 = x1 & ~x2;
assign n_3 = ~x6 & ~x7;
assign n_4 = ~x12 & ~x13;
assign n_5 = ~x16 & x17;
assign n_6 = x17 ^ x16;
assign n_7 = x18 & ~x19;
assign n_8 = x21 ^ x20;
assign n_9 = x22 ^ x21;
assign n_10 = x19 & ~x22;
assign n_11 = x12 & ~x22;
assign n_12 = x13 & ~x22;
assign n_13 = x6 & ~x22;
assign n_14 = x22 ^ x2;
assign n_15 = x0 & ~x22;
assign n_16 = x22 ^ x1;
assign n_17 = ~x21 & ~x22;
assign n_18 = x23 ^ x22;
assign n_19 = n_0 ^ x0;
assign n_20 = x22 & n_0;
assign n_21 = n_1 & n_0;
assign n_22 = n_2 ^ n_1;
assign n_23 = ~x14 & n_4;
assign n_24 = n_5 ^ x16;
assign n_25 = n_7 ^ x18;
assign n_26 = x22 & n_7;
assign n_27 = n_9 & ~n_8;
assign n_28 = ~x18 & n_10;
assign n_29 = n_10 ^ x19;
assign n_30 = n_10 ^ x22;
assign n_31 = n_15 ^ x0;
assign n_32 = ~x2 & ~n_15;
assign n_33 = n_15 ^ x2;
assign n_34 = ~n_1 & ~n_19;
assign n_35 = n_20 ^ n_1;
assign n_36 = n_21 ^ n_1;
assign n_37 = n_14 & ~n_22;
assign n_38 = n_24 ^ x17;
assign n_39 = n_25 ^ x19;
assign n_40 = ~n_24 & n_25;
assign n_41 = ~n_24 & n_26;
assign n_42 = n_26 ^ n_7;
assign n_43 = n_5 & n_26;
assign n_44 = x2 & ~n_31;
assign n_45 = n_31 ^ x1;
assign n_46 = n_32 ^ n_33;
assign n_47 = ~x3 & n_34;
assign n_48 = n_34 ^ n_19;
assign n_49 = n_19 & n_37;
assign n_50 = n_37 ^ x22;
assign n_51 = n_38 ^ x16;
assign n_52 = n_38 & n_26;
assign n_53 = n_39 ^ x18;
assign n_54 = n_28 ^ n_39;
assign n_55 = n_42 ^ n_30;
assign n_56 = n_44 ^ n_32;
assign n_57 = n_45 ^ n_0;
assign n_58 = ~x4 & n_47;
assign n_59 = ~x22 & ~n_47;
assign n_60 = n_48 ^ n_36;
assign n_61 = n_49 ^ n_34;
assign n_62 = n_26 & n_51;
assign n_63 = ~n_24 & ~n_53;
assign n_64 = n_54 ^ n_29;
assign n_65 = n_5 & n_54;
assign n_66 = n_54 & n_51;
assign n_67 = n_38 & n_54;
assign n_68 = n_55 ^ n_53;
assign n_69 = n_56 ^ n_49;
assign n_70 = n_56 ^ n_48;
assign n_71 = n_46 ^ n_57;
assign n_72 = ~x5 & n_58;
assign n_73 = ~x22 & ~n_58;
assign n_74 = n_59 ^ x4;
assign n_75 = n_60 ^ x0;
assign n_76 = n_61 ^ n_50;
assign n_77 = n_64 ^ n_25;
assign n_78 = n_64 & n_51;
assign n_79 = n_38 & n_64;
assign n_80 = n_5 & n_64;
assign n_81 = n_68 & n_51;
assign n_82 = n_5 & n_68;
assign n_83 = n_38 & n_68;
assign n_84 = ~n_61 & ~n_71;
assign n_85 = ~x22 & ~n_72;
assign n_86 = n_72 & n_3;
assign n_87 = n_73 ^ x5;
assign n_88 = n_76 ^ x3;
assign n_89 = n_84 ^ n_60;
assign n_90 = n_85 ^ x6;
assign n_91 = ~n_85 & ~n_13;
assign n_92 = ~x8 & n_86;
assign n_93 = ~x22 & ~n_86;
assign n_94 = n_74 ^ n_87;
assign n_95 = n_87 & ~n_74;
assign n_96 = n_88 ^ n_74;
assign n_97 = n_89 ^ n_61;
assign n_98 = n_87 ^ n_90;
assign n_99 = n_90 & n_87;
assign n_100 = x7 ^ n_91;
assign n_101 = ~x9 & n_92;
assign n_102 = ~x22 & ~n_92;
assign n_103 = n_93 ^ x8;
assign n_104 = n_94 ^ n_95;
assign n_105 = n_97 ^ n_35;
assign n_106 = n_99 ^ n_98;
assign n_107 = n_100 & n_98;
assign n_108 = n_99 ^ n_100;
assign n_109 = ~x10 & n_101;
assign n_110 = ~x22 & ~n_101;
assign n_111 = n_102 ^ x9;
assign n_112 = n_103 ^ n_100;
assign n_113 = n_100 & ~n_103;
assign n_114 = ~n_103 & n_99;
assign n_115 = n_104 ^ n_95;
assign n_116 = n_69 ^ n_105;
assign n_117 = ~n_103 & ~n_106;
assign n_118 = n_107 ^ n_100;
assign n_119 = ~x11 & n_109;
assign n_120 = ~x22 & ~n_109;
assign n_121 = n_110 ^ x10;
assign n_122 = n_103 ^ n_111;
assign n_123 = n_111 & n_103;
assign n_124 = n_106 & ~n_113;
assign n_125 = n_113 ^ n_112;
assign n_126 = n_114 ^ n_100;
assign n_127 = ~n_88 & n_115;
assign n_128 = n_116 ^ n_84;
assign n_129 = n_117 ^ n_106;
assign n_130 = n_118 ^ n_106;
assign n_131 = n_118 ^ n_99;
assign n_132 = ~x22 & ~n_119;
assign n_133 = n_119 & n_23;
assign n_134 = n_120 ^ x11;
assign n_135 = n_121 ^ n_111;
assign n_136 = n_121 & n_122;
assign n_137 = n_122 ^ n_123;
assign n_138 = n_124 ^ n_113;
assign n_139 = n_124 ^ n_103;
assign n_140 = n_127 ^ n_95;
assign n_141 = n_128 ^ n_34;
assign n_142 = ~n_100 & n_130;
assign n_143 = n_103 & ~n_130;
assign n_144 = n_130 ^ n_103;
assign n_145 = n_132 ^ x12;
assign n_146 = ~n_132 & ~n_11;
assign n_147 = ~x22 & ~n_133;
assign n_148 = ~x15 & n_133;
assign n_149 = n_134 & ~n_122;
assign n_150 = n_121 ^ n_134;
assign n_151 = n_122 ^ n_134;
assign n_152 = n_136 ^ n_122;
assign n_153 = ~n_134 & n_136;
assign n_154 = n_137 ^ n_134;
assign n_155 = n_137 ^ n_121;
assign n_156 = n_138 ^ n_129;
assign n_157 = n_141 ^ n_88;
assign n_158 = ~n_88 & ~n_141;
assign n_159 = ~n_74 & ~n_141;
assign n_160 = n_141 ^ n_87;
assign n_161 = n_142 ^ n_138;
assign n_162 = n_143 ^ n_130;
assign n_163 = n_134 ^ n_145;
assign n_164 = n_145 & n_134;
assign n_165 = x13 ^ n_146;
assign n_166 = ~n_12 & n_146;
assign n_167 = n_147 ^ x15;
assign n_168 = ~x22 & ~n_148;
assign n_169 = ~n_148 & n_51;
assign n_170 = n_148 ^ x16;
assign n_171 = n_148 ^ x18;
assign n_172 = ~n_148 & ~n_6;
assign n_173 = n_149 ^ n_134;
assign n_174 = n_152 ^ n_121;
assign n_175 = n_154 & ~n_155;
assign n_176 = ~n_74 & ~n_157;
assign n_177 = n_87 & n_157;
assign n_178 = n_157 ^ n_87;
assign n_179 = n_158 ^ n_141;
assign n_180 = n_158 ^ n_88;
assign n_181 = n_159 ^ n_88;
assign n_182 = n_159 ^ n_141;
assign n_183 = n_162 ^ n_156;
assign n_184 = n_163 ^ n_164;
assign n_185 = n_164 & n_165;
assign n_186 = n_165 ^ n_164;
assign n_187 = x14 ^ n_166;
assign n_188 = ~n_9 & n_167;
assign n_189 = ~n_167 & n_27;
assign n_190 = ~n_168 & n_39;
assign n_191 = ~n_168 & n_63;
assign n_192 = n_77 & n_169;
assign n_193 = n_42 & n_169;
assign n_194 = ~x17 & ~n_170;
assign n_195 = n_171 ^ x22;
assign n_196 = n_24 ^ n_172;
assign n_197 = n_174 ^ n_137;
assign n_198 = n_175 ^ n_153;
assign n_199 = n_176 ^ n_157;
assign n_200 = n_176 ^ n_74;
assign n_201 = n_177 ^ n_87;
assign n_202 = ~n_74 & ~n_179;
assign n_203 = n_179 ^ n_74;
assign n_204 = n_179 ^ n_87;
assign n_205 = n_183 ^ n_126;
assign n_206 = ~n_184 & ~n_165;
assign n_207 = n_165 ^ n_187;
assign n_208 = ~n_187 & n_165;
assign n_209 = ~n_184 & n_187;
assign n_210 = n_164 & ~n_187;
assign n_211 = n_187 ^ n_184;
assign n_212 = n_87 ^ n_187;
assign n_213 = n_189 ^ n_27;
assign n_214 = ~n_24 & n_190;
assign n_215 = ~x22 & ~n_191;
assign n_216 = n_192 ^ n_191;
assign n_217 = n_194 ^ n_170;
assign n_218 = ~n_55 & n_194;
assign n_219 = n_77 & n_194;
assign n_220 = n_42 & n_194;
assign n_221 = n_28 & n_194;
assign n_222 = n_196 ^ n_171;
assign n_223 = n_170 ^ n_196;
assign n_224 = n_201 ^ n_157;
assign n_225 = n_200 ^ n_202;
assign n_226 = n_202 ^ n_179;
assign n_227 = n_202 ^ n_87;
assign n_228 = ~n_87 & n_202;
assign n_229 = n_181 ^ n_203;
assign n_230 = ~n_203 & n_204;
assign n_231 = n_161 ^ n_205;
assign n_232 = n_206 ^ n_184;
assign n_233 = n_206 ^ n_165;
assign n_234 = n_185 ^ n_206;
assign n_235 = n_207 ^ n_184;
assign n_236 = n_208 ^ n_207;
assign n_237 = n_209 ^ n_184;
assign n_238 = n_185 ^ n_209;
assign n_239 = ~n_165 & n_209;
assign n_240 = n_210 ^ n_164;
assign n_241 = n_193 ^ n_214;
assign n_242 = n_215 ^ x20;
assign n_243 = n_215 ^ x21;
assign n_244 = n_216 & n_213;
assign n_245 = n_189 & n_216;
assign n_246 = n_28 & ~n_217;
assign n_247 = ~n_55 & ~n_217;
assign n_248 = n_77 & ~n_217;
assign n_249 = n_42 & ~n_217;
assign n_250 = n_218 ^ n_78;
assign n_251 = n_219 ^ n_81;
assign n_252 = n_220 ^ n_66;
assign n_253 = n_221 ^ n_62;
assign n_254 = n_195 & n_222;
assign n_255 = ~n_55 & ~n_223;
assign n_256 = n_77 & ~n_223;
assign n_257 = n_42 & ~n_223;
assign n_258 = n_28 & ~n_223;
assign n_259 = n_224 ^ n_87;
assign n_260 = n_225 ^ n_226;
assign n_261 = n_228 ^ n_179;
assign n_262 = n_229 ^ n_182;
assign n_263 = ~n_187 & n_232;
assign n_264 = n_233 ^ n_187;
assign n_265 = n_234 ^ n_187;
assign n_266 = n_240 ^ n_237;
assign n_267 = n_240 ^ n_165;
assign n_268 = n_189 & n_241;
assign n_269 = n_213 & n_241;
assign n_270 = n_241 ^ n_213;
assign n_271 = ~n_9 & n_242;
assign n_272 = ~n_242 & n_167;
assign n_273 = n_8 & n_243;
assign n_274 = n_246 ^ n_52;
assign n_275 = n_247 ^ n_79;
assign n_276 = n_248 ^ n_83;
assign n_277 = n_249 ^ n_67;
assign n_278 = n_27 & n_250;
assign n_279 = n_213 & n_250;
assign n_280 = n_27 & n_251;
assign n_281 = n_189 & n_251;
assign n_282 = ~n_167 & ~n_251;
assign n_283 = n_251 ^ n_241;
assign n_284 = ~n_167 & n_252;
assign n_285 = n_252 & n_189;
assign n_286 = n_252 & n_213;
assign n_287 = ~n_189 & ~n_253;
assign n_288 = n_253 ^ n_189;
assign n_289 = n_253 ^ n_252;
assign n_290 = n_27 & n_253;
assign n_291 = n_188 & n_253;
assign n_292 = n_253 ^ n_216;
assign n_293 = n_254 ^ n_172;
assign n_294 = n_255 ^ n_80;
assign n_295 = n_256 ^ n_82;
assign n_296 = n_257 ^ n_65;
assign n_297 = n_258 ^ n_43;
assign n_298 = n_260 ^ n_87;
assign n_299 = n_87 & ~n_260;
assign n_300 = n_260 ^ n_157;
assign n_301 = n_207 & ~n_266;
assign n_302 = n_211 ^ n_266;
assign n_303 = n_266 ^ n_185;
assign n_304 = n_244 ^ n_269;
assign n_305 = n_269 ^ n_270;
assign n_306 = ~n_271 & ~n_167;
assign n_307 = n_271 ^ n_242;
assign n_308 = n_271 & n_251;
assign n_309 = n_271 & n_252;
assign n_310 = n_271 & n_250;
assign n_311 = n_272 ^ n_167;
assign n_312 = n_273 & n_251;
assign n_313 = n_273 & n_241;
assign n_314 = ~n_273 ^ ~n_252;
assign n_315 = n_274 ^ n_213;
assign n_316 = ~n_213 & ~n_274;
assign n_317 = n_189 & n_274;
assign n_318 = n_271 & n_274;
assign n_319 = n_188 & n_274;
assign n_320 = n_250 ^ n_275;
assign n_321 = n_273 & n_275;
assign n_322 = n_275 ^ n_252;
assign n_323 = n_271 & n_275;
assign n_324 = n_189 & n_275;
assign n_325 = n_275 & n_213;
assign n_326 = n_276 & n_27;
assign n_327 = n_216 ^ n_276;
assign n_328 = n_276 & n_189;
assign n_329 = n_167 ^ ~n_276;
assign n_330 = ~n_167 & n_277;
assign n_331 = n_271 & n_277;
assign n_332 = n_277 ^ n_241;
assign n_333 = n_213 & n_277;
assign n_334 = n_277 ^ n_252;
assign n_335 = n_277 ^ n_271;
assign n_336 = n_189 & n_277;
assign n_337 = n_251 ^ n_277;
assign n_338 = n_278 ^ n_279;
assign n_339 = n_279 ^ n_250;
assign n_340 = n_280 ^ n_281;
assign n_341 = n_283 ^ n_274;
assign n_342 = n_287 ^ n_27;
assign n_343 = n_288 ^ n_287;
assign n_344 = n_271 & n_292;
assign n_345 = ~n_167 & n_292;
assign n_346 = n_293 ^ n_24;
assign n_347 = ~n_271 ^ ~n_294;
assign n_348 = n_294 ^ n_213;
assign n_349 = n_213 & n_294;
assign n_350 = n_294 ^ n_253;
assign n_351 = n_294 ^ n_251;
assign n_352 = n_251 ^ n_295;
assign n_353 = n_213 & n_295;
assign n_354 = n_189 & n_295;
assign n_355 = n_271 & n_295;
assign n_356 = n_167 & n_295;
assign n_357 = n_241 ^ n_295;
assign n_358 = n_213 & n_296;
assign n_359 = n_189 & n_296;
assign n_360 = n_289 ^ n_296;
assign n_361 = ~n_167 & ~n_296;
assign n_362 = n_296 ^ n_274;
assign n_363 = n_296 ^ n_294;
assign n_364 = n_296 ^ n_250;
assign n_365 = ~n_167 & n_297;
assign n_366 = n_213 & n_297;
assign n_367 = n_273 & n_297;
assign n_368 = n_189 & n_297;
assign n_369 = ~n_271 & ~n_297;
assign n_370 = n_297 ^ n_277;
assign n_371 = n_297 ^ n_253;
assign n_372 = n_177 ^ n_299;
assign n_373 = n_299 ^ n_87;
assign n_374 = n_300 ^ n_227;
assign n_375 = n_303 ^ n_301;
assign n_376 = ~n_216 ^ ~n_305;
assign n_377 = n_306 ^ n_167;
assign n_378 = n_306 & n_252;
assign n_379 = ~n_307 & n_282;
assign n_380 = n_189 ^ n_307;
assign n_381 = ~n_307 & ~n_189;
assign n_382 = n_311 ^ n_242;
assign n_383 = n_189 ^ n_311;
assign n_384 = n_311 & n_275;
assign n_385 = n_311 & n_276;
assign n_386 = n_311 & n_241;
assign n_387 = n_315 ^ n_316;
assign n_388 = n_320 ^ n_294;
assign n_389 = n_313 ^ n_321;
assign n_390 = n_312 ^ n_321;
assign n_391 = n_324 ^ n_281;
assign n_392 = n_326 ^ n_216;
assign n_393 = n_328 ^ n_326;
assign n_394 = n_245 ^ n_328;
assign n_395 = n_271 & n_330;
assign n_396 = n_273 & n_330;
assign n_397 = n_307 & n_330;
assign n_398 = n_273 & n_332;
assign n_399 = n_334 ^ n_296;
assign n_400 = n_335 ^ n_331;
assign n_401 = n_338 ^ n_286;
assign n_402 = n_324 ^ n_338;
assign n_403 = n_338 ^ n_281;
assign n_404 = n_339 ^ n_316;
assign n_405 = n_325 ^ n_340;
assign n_406 = n_271 & n_341;
assign n_407 = n_290 ^ n_342;
assign n_408 = n_343 ^ n_290;
assign n_409 = n_345 ^ n_241;
assign n_410 = n_346 ^ x22;
assign n_411 = n_348 ^ n_349;
assign n_412 = n_349 ^ n_285;
assign n_413 = n_319 ^ n_349;
assign n_414 = n_351 ^ n_332;
assign n_415 = n_352 ^ n_327;
assign n_416 = n_188 & n_352;
assign n_417 = n_343 ^ n_353;
assign n_418 = n_280 ^ n_353;
assign n_419 = n_273 & n_356;
assign n_420 = n_279 ^ n_358;
assign n_421 = n_273 & n_360;
assign n_422 = ~n_361 & n_362;
assign n_423 = n_272 & n_362;
assign n_424 = n_307 & n_365;
assign n_425 = n_271 & n_365;
assign n_426 = n_365 ^ n_275;
assign n_427 = n_361 ^ n_365;
assign n_428 = n_366 ^ n_297;
assign n_429 = n_368 ^ n_318;
assign n_430 = n_371 ^ n_274;
assign n_431 = n_372 ^ n_374;
assign n_432 = n_375 ^ n_264;
assign n_433 = n_377 ^ n_271;
assign n_434 = ~n_377 & n_216;
assign n_435 = ~n_377 & n_296;
assign n_436 = n_273 ^ n_377;
assign n_437 = ~n_377 & n_294;
assign n_438 = ~n_377 & n_276;
assign n_439 = ~n_377 & n_253;
assign n_440 = n_189 ^ n_377;
assign n_441 = n_274 ^ n_377;
assign n_442 = n_216 ^ n_377;
assign n_443 = n_213 ^ n_377;
assign n_444 = ~n_377 & n_283;
assign n_445 = n_378 ^ n_284;
assign n_446 = n_378 ^ n_285;
assign n_447 = n_379 ^ n_282;
assign n_448 = n_380 ^ n_381;
assign n_449 = n_216 & n_381;
assign n_450 = n_216 & n_382;
assign n_451 = n_253 & n_382;
assign n_452 = n_241 & n_382;
assign n_453 = n_252 & n_383;
assign n_454 = n_383 & n_283;
assign n_455 = n_387 ^ n_317;
assign n_456 = n_189 & ~n_388;
assign n_457 = n_389 ^ n_343;
assign n_458 = n_244 ^ n_393;
assign n_459 = n_395 ^ n_331;
assign n_460 = n_387 ^ n_395;
assign n_461 = n_359 ^ n_395;
assign n_462 = n_396 ^ n_333;
assign n_463 = n_396 ^ n_286;
assign n_464 = n_325 ^ n_397;
assign n_465 = n_27 & n_399;
assign n_466 = n_400 ^ n_370;
assign n_467 = n_408 ^ n_286;
assign n_468 = ~n_171 & n_410;
assign n_469 = n_412 ^ n_268;
assign n_470 = n_273 & n_415;
assign n_471 = n_418 ^ n_358;
assign n_472 = n_419 ^ n_397;
assign n_473 = n_419 ^ n_387;
assign n_474 = n_420 ^ n_340;
assign n_475 = n_422 ^ n_332;
assign n_476 = n_397 ^ n_424;
assign n_477 = n_425 ^ n_395;
assign n_478 = n_333 ^ n_425;
assign n_479 = n_273 & n_426;
assign n_480 = n_428 ^ n_316;
assign n_481 = n_429 ^ n_353;
assign n_482 = n_431 ^ n_202;
assign n_483 = n_432 ^ n_301;
assign n_484 = n_188 ^ n_433;
assign n_485 = n_433 ^ n_311;
assign n_486 = ~n_433 & n_216;
assign n_487 = ~n_433 & n_296;
assign n_488 = ~n_433 & n_274;
assign n_489 = ~n_433 & n_297;
assign n_490 = ~n_433 & n_275;
assign n_491 = ~n_433 & n_294;
assign n_492 = ~n_433 & n_276;
assign n_493 = ~n_433 & n_295;
assign n_494 = ~n_433 & n_250;
assign n_495 = n_253 ^ n_433;
assign n_496 = ~n_433 & n_251;
assign n_497 = n_433 ^ ~n_363;
assign n_498 = n_368 ^ n_433;
assign n_499 = n_325 ^ n_435;
assign n_500 = n_244 ^ n_435;
assign n_501 = n_435 ^ n_437;
assign n_502 = n_244 ^ n_438;
assign n_503 = n_438 ^ n_216;
assign n_504 = n_439 ^ n_434;
assign n_505 = n_241 & ~n_440;
assign n_506 = ~n_440 & n_334;
assign n_507 = n_442 ^ n_434;
assign n_508 = n_327 & ~n_443;
assign n_509 = n_435 ^ n_445;
assign n_510 = n_445 ^ n_309;
assign n_511 = n_408 ^ n_445;
assign n_512 = n_439 ^ n_445;
assign n_513 = n_451 ^ n_439;
assign n_514 = n_452 ^ n_438;
assign n_515 = n_456 ^ n_189;
assign n_516 = n_394 ^ n_457;
assign n_517 = n_407 ^ n_459;
assign n_518 = n_464 ^ n_424;
assign n_519 = n_466 ^ n_369;
assign n_520 = n_467 ^ n_424;
assign n_521 = n_171 ^ n_468;
assign n_522 = n_470 ^ n_273;
assign n_523 = n_473 ^ n_359;
assign n_524 = n_474 ^ n_324;
assign n_525 = n_475 ^ n_371;
assign n_526 = n_476 ^ n_349;
assign n_527 = n_477 ^ n_397;
assign n_528 = n_478 ^ n_356;
assign n_529 = n_479 ^ n_354;
assign n_530 = ~n_481 ^ ~n_401;
assign n_531 = n_482 ^ n_228;
assign n_532 = n_484 & ~n_216;
assign n_533 = ~n_484 & n_275;
assign n_534 = n_484 ^ n_273;
assign n_535 = ~n_484 & n_253;
assign n_536 = n_216 ^ n_484;
assign n_537 = ~n_484 & n_250;
assign n_538 = n_276 & ~n_484;
assign n_539 = ~n_484 & n_251;
assign n_540 = ~n_484 & n_241;
assign n_541 = ~n_484 & n_294;
assign n_542 = ~n_484 & n_297;
assign n_543 = ~n_484 & n_252;
assign n_544 = ~n_484 & n_277;
assign n_545 = n_354 ^ n_484;
assign n_546 = ~n_484 & n_414;
assign n_547 = ~n_484 & n_364;
assign n_548 = n_279 ^ n_484;
assign n_549 = ~n_484 & n_357;
assign n_550 = n_484 ^ n_307;
assign n_551 = ~n_485 & n_274;
assign n_552 = ~n_485 & n_250;
assign n_553 = n_485 ^ n_307;
assign n_554 = n_297 ^ n_485;
assign n_555 = n_485 & ~n_297;
assign n_556 = n_287 ^ n_485;
assign n_557 = n_485 & n_287;
assign n_558 = ~n_485 & n_251;
assign n_559 = ~n_485 & n_277;
assign n_560 = ~n_485 & n_294;
assign n_561 = ~n_485 & n_296;
assign n_562 = ~n_485 & n_216;
assign n_563 = ~n_485 & n_241;
assign n_564 = ~n_485 & n_371;
assign n_565 = ~n_485 & n_295;
assign n_566 = ~n_485 & n_334;
assign n_567 = n_414 ^ n_485;
assign n_568 = ~n_485 & n_350;
assign n_569 = n_486 ^ n_434;
assign n_570 = n_486 ^ n_216;
assign n_571 = n_313 ^ n_487;
assign n_572 = n_359 ^ n_487;
assign n_573 = n_424 ^ n_487;
assign n_574 = n_488 ^ n_487;
assign n_575 = n_488 ^ n_318;
assign n_576 = n_488 ^ n_310;
assign n_577 = ~n_489 ^ ~n_406;
assign n_578 = n_413 ^ n_489;
assign n_579 = n_384 ^ n_490;
assign n_580 = n_490 ^ n_323;
assign n_581 = n_472 ^ n_490;
assign n_582 = n_279 ^ n_490;
assign n_583 = n_492 ^ n_486;
assign n_584 = n_385 ^ n_492;
assign n_585 = n_492 ^ n_340;
assign n_586 = n_355 ^ n_493;
assign n_587 = n_493 ^ n_437;
assign n_588 = n_343 ^ n_494;
assign n_589 = n_494 ^ n_310;
assign n_590 = n_349 ^ n_494;
assign n_591 = n_494 ^ n_489;
assign n_592 = n_496 ^ n_308;
assign n_593 = n_496 ^ n_330;
assign n_594 = n_496 ^ n_459;
assign n_595 = n_500 ^ n_492;
assign n_596 = n_505 ^ n_268;
assign n_597 = n_503 ^ n_507;
assign n_598 = n_510 ^ n_285;
assign n_599 = n_459 ^ n_510;
assign n_600 = n_494 ^ n_510;
assign n_601 = n_493 ^ n_510;
assign n_602 = n_393 ^ n_510;
assign n_603 = n_489 ^ n_510;
assign n_604 = n_513 ^ n_424;
assign n_605 = n_402 ^ n_515;
assign n_606 = ~n_369 & ~n_517;
assign n_607 = x19 & ~n_521;
assign n_608 = n_521 ^ ~n_40;
assign n_609 = n_522 ^ n_456;
assign n_610 = n_307 & n_525;
assign n_611 = n_27 & n_525;
assign n_612 = ~n_505 ^ ~n_526;
assign n_613 = n_259 ^ n_531;
assign n_614 = n_531 ^ n_202;
assign n_615 = ~n_532 & n_497;
assign n_616 = n_533 ^ n_321;
assign n_617 = n_310 ^ n_533;
assign n_618 = n_396 ^ n_533;
assign n_619 = n_534 ^ n_485;
assign n_620 = ~n_534 & n_253;
assign n_621 = n_276 & ~n_534;
assign n_622 = ~n_534 & n_252;
assign n_623 = ~n_534 & n_216;
assign n_624 = ~n_534 & n_296;
assign n_625 = n_189 ^ n_534;
assign n_626 = ~n_534 & n_295;
assign n_627 = ~n_534 & n_415;
assign n_628 = ~n_534 & n_294;
assign n_629 = n_534 ^ ~n_350;
assign n_630 = ~n_534 & n_370;
assign n_631 = ~n_534 & n_430;
assign n_632 = n_216 ^ n_534;
assign n_633 = n_488 ^ n_535;
assign n_634 = n_535 ^ n_291;
assign n_635 = n_532 ^ n_536;
assign n_636 = n_489 ^ n_537;
assign n_637 = n_537 ^ n_271;
assign n_638 = n_514 ^ n_537;
assign n_639 = n_538 ^ n_281;
assign n_640 = n_333 ^ n_538;
assign n_641 = n_354 ^ n_538;
assign n_642 = n_419 ^ n_538;
assign n_643 = n_539 ^ n_312;
assign n_644 = n_539 ^ n_532;
assign n_645 = n_539 ^ n_537;
assign n_646 = n_319 ^ n_539;
assign n_647 = n_313 ^ n_540;
assign n_648 = n_540 ^ n_368;
assign n_649 = n_454 ^ n_540;
assign n_650 = n_444 ^ n_540;
assign n_651 = n_491 ^ n_541;
assign n_652 = n_541 ^ n_294;
assign n_653 = n_541 ^ n_509;
assign n_654 = n_333 ^ n_541;
assign n_655 = n_359 ^ n_541;
assign n_656 = n_535 ^ n_541;
assign n_657 = n_367 ^ n_542;
assign n_658 = ~n_542 ^ ~n_421;
assign n_659 = n_542 ^ n_509;
assign n_660 = n_542 ^ n_340;
assign n_661 = n_542 ^ n_353;
assign n_662 = n_544 ^ n_543;
assign n_663 = n_245 ^ n_544;
assign n_664 = n_544 ^ n_419;
assign n_665 = n_544 ^ n_453;
assign n_666 = n_547 ^ n_544;
assign n_667 = ~n_550 & n_409;
assign n_668 = n_551 ^ n_274;
assign n_669 = n_539 ^ n_551;
assign n_670 = n_490 ^ n_551;
assign n_671 = n_425 ^ n_551;
assign n_672 = n_387 ^ n_552;
assign n_673 = ~n_553 & n_250;
assign n_674 = ~n_553 & n_275;
assign n_675 = ~n_553 & n_274;
assign n_676 = n_447 ^ n_553;
assign n_677 = ~n_553 & n_276;
assign n_678 = n_484 ^ n_553;
assign n_679 = ~n_553 & n_296;
assign n_680 = ~n_553 & n_295;
assign n_681 = ~n_553 & n_283;
assign n_682 = n_470 ^ n_553;
assign n_683 = n_554 ^ n_555;
assign n_684 = ~n_555 & n_305;
assign n_685 = n_556 ^ n_557;
assign n_686 = n_558 ^ n_279;
assign n_687 = n_558 ^ n_537;
assign n_688 = n_559 ^ n_358;
assign n_689 = n_559 ^ n_490;
assign n_690 = n_344 ^ n_559;
assign n_691 = n_423 ^ n_560;
assign n_692 = n_560 ^ n_439;
assign n_693 = n_561 ^ n_552;
assign n_694 = n_477 ^ n_561;
assign n_695 = n_561 ^ n_533;
assign n_696 = n_367 ^ n_561;
assign n_697 = n_563 ^ n_386;
assign n_698 = n_563 ^ n_424;
assign n_699 = n_563 ^ n_559;
assign n_700 = n_565 ^ n_393;
assign n_701 = n_565 ^ n_533;
assign n_702 = n_565 ^ n_563;
assign n_703 = ~n_377 & n_567;
assign n_704 = n_568 ^ n_538;
assign n_705 = ~n_569 & ~n_450;
assign n_706 = n_572 ^ n_338;
assign n_707 = n_575 ^ n_441;
assign n_708 = n_504 ^ n_575;
assign n_709 = n_575 ^ n_459;
assign n_710 = n_565 ^ n_575;
assign n_711 = n_368 ^ n_579;
assign n_712 = n_286 ^ n_579;
assign n_713 = n_580 ^ n_538;
assign n_714 = n_540 ^ n_580;
assign n_715 = n_420 ^ n_580;
assign n_716 = n_518 ^ n_582;
assign n_717 = n_584 ^ n_353;
assign n_718 = n_336 ^ n_584;
assign n_719 = n_585 ^ n_397;
assign n_720 = n_585 ^ n_387;
assign n_721 = n_585 ^ n_540;
assign n_722 = n_586 ^ n_496;
assign n_723 = n_587 ^ n_538;
assign n_724 = n_589 ^ n_397;
assign n_725 = n_564 ^ n_589;
assign n_726 = n_590 ^ n_586;
assign n_727 = n_592 ^ n_509;
assign n_728 = n_594 ^ n_269;
assign n_729 = n_596 ^ n_452;
assign n_730 = n_543 ^ n_596;
assign n_731 = n_598 ^ n_453;
assign n_732 = n_600 ^ n_487;
assign n_733 = n_604 ^ n_551;
assign n_734 = n_605 ^ n_365;
assign n_735 = n_393 ^ n_605;
assign n_736 = n_605 ^ n_487;
assign n_737 = n_605 ^ n_317;
assign n_738 = n_605 ^ n_435;
assign n_739 = n_607 ^ n_41;
assign n_740 = ~n_10 & n_608;
assign n_741 = n_355 ^ n_609;
assign n_742 = ~n_584 ^ ~n_612;
assign n_743 = n_613 ^ n_373;
assign n_744 = n_572 ^ n_615;
assign n_745 = n_338 ^ n_616;
assign n_746 = n_494 ^ n_616;
assign n_747 = n_535 ^ n_616;
assign n_748 = n_400 ^ n_616;
assign n_749 = n_250 & n_619;
assign n_750 = n_620 ^ n_338;
assign n_751 = n_620 ^ n_580;
assign n_752 = n_537 ^ n_621;
assign n_753 = n_533 ^ n_621;
assign n_754 = n_586 ^ n_621;
assign n_755 = n_596 ^ n_621;
assign n_756 = n_560 ^ n_621;
assign n_757 = n_446 ^ n_622;
assign n_758 = n_552 ^ n_622;
assign n_759 = n_623 ^ n_324;
assign n_760 = n_623 ^ n_317;
assign n_761 = n_458 ^ n_623;
assign n_762 = n_624 ^ n_336;
assign n_763 = n_274 & ~n_625;
assign n_764 = ~n_625 & n_283;
assign n_765 = n_626 ^ n_586;
assign n_766 = n_336 ^ n_626;
assign n_767 = n_268 ^ n_628;
assign n_768 = n_333 ^ n_628;
assign n_769 = n_618 ^ n_628;
assign n_770 = n_573 ^ n_628;
assign n_771 = n_629 & ~n_480;
assign n_772 = n_630 ^ n_393;
assign n_773 = ~n_537 ^ ~n_631;
assign n_774 = n_633 ^ n_620;
assign n_775 = n_633 ^ n_310;
assign n_776 = n_512 ^ n_633;
assign n_777 = n_633 ^ n_340;
assign n_778 = n_634 ^ n_495;
assign n_779 = n_491 ^ n_634;
assign n_780 = n_387 ^ n_635;
assign n_781 = n_620 ^ n_635;
assign n_782 = n_537 ^ n_635;
assign n_783 = n_597 ^ n_635;
assign n_784 = n_638 ^ n_317;
assign n_785 = n_639 ^ n_437;
assign n_786 = ~n_639 ^ n_523;
assign n_787 = n_541 ^ n_639;
assign n_788 = n_498 ^ n_642;
assign n_789 = n_643 ^ n_387;
assign n_790 = n_628 ^ n_643;
assign n_791 = n_449 ^ n_644;
assign n_792 = n_645 ^ n_494;
assign n_793 = n_646 ^ n_488;
assign n_794 = n_647 ^ n_353;
assign n_795 = n_328 ^ n_647;
assign n_796 = n_648 ^ n_424;
assign n_797 = n_651 ^ n_583;
assign n_798 = ~n_655 ^ n_516;
assign n_799 = n_656 ^ n_395;
assign n_800 = ~n_657 ^ ~n_577;
assign n_801 = n_663 ^ n_328;
assign n_802 = n_663 ^ n_490;
assign n_803 = n_663 ^ n_586;
assign n_804 = n_641 ^ n_664;
assign n_805 = n_665 ^ n_451;
assign n_806 = n_666 ^ n_561;
assign n_807 = n_670 ^ n_499;
assign n_808 = n_343 ^ n_673;
assign n_809 = n_624 ^ n_673;
assign n_810 = n_425 ^ n_673;
assign n_811 = n_674 ^ n_635;
assign n_812 = n_628 ^ n_674;
assign n_813 = n_469 ^ n_674;
assign n_814 = n_675 ^ n_353;
assign n_815 = n_560 ^ n_675;
assign n_816 = n_336 ^ n_675;
assign n_817 = n_490 ^ n_675;
assign n_818 = n_462 ^ n_675;
assign n_819 = n_676 ^ n_624;
assign n_820 = n_676 ^ n_448;
assign n_821 = n_676 ^ n_647;
assign n_822 = n_676 ^ n_559;
assign n_823 = n_677 ^ n_584;
assign n_824 = n_294 & ~n_678;
assign n_825 = n_678 & n_422;
assign n_826 = ~n_678 & ~n_337;
assign n_827 = n_679 ^ n_494;
assign n_828 = n_662 ^ n_679;
assign n_829 = n_679 ^ n_634;
assign n_830 = n_679 ^ n_558;
assign n_831 = n_680 ^ n_393;
assign n_832 = n_680 ^ n_676;
assign n_833 = n_681 ^ n_542;
assign n_834 = n_295 & ~n_682;
assign n_835 = ~n_682 & n_357;
assign n_836 = n_340 ^ n_683;
assign n_837 = n_460 ^ n_683;
assign n_838 = n_563 ^ n_683;
assign n_839 = n_336 ^ n_683;
assign n_840 = n_435 ^ n_683;
assign n_841 = n_684 ^ n_324;
assign n_842 = n_684 ^ n_408;
assign n_843 = n_552 ^ n_685;
assign n_844 = n_268 ^ n_685;
assign n_845 = n_685 ^ n_486;
assign n_846 = n_679 ^ n_685;
assign n_847 = n_686 ^ n_340;
assign n_848 = n_688 ^ n_435;
assign n_849 = n_688 ^ n_669;
assign n_850 = ~n_692 ^ ~n_667;
assign n_851 = ~n_694 & ~n_610;
assign n_852 = n_697 ^ n_439;
assign n_853 = n_586 ^ n_697;
assign n_854 = n_691 ^ n_697;
assign n_855 = n_697 ^ n_510;
assign n_856 = n_700 ^ n_552;
assign n_857 = n_703 ^ n_485;
assign n_858 = n_704 ^ n_535;
assign n_859 = n_569 ^ n_705;
assign n_860 = n_706 ^ n_626;
assign n_861 = n_690 ^ n_708;
assign n_862 = n_709 ^ n_349;
assign n_863 = n_710 ^ n_542;
assign n_864 = n_712 ^ n_368;
assign n_865 = n_416 ^ n_712;
assign n_866 = n_713 ^ n_496;
assign n_867 = n_714 ^ n_544;
assign n_868 = n_720 ^ n_331;
assign n_869 = n_721 ^ n_439;
assign n_870 = n_722 ^ n_492;
assign n_871 = n_358 ^ n_724;
assign n_872 = n_725 ^ n_511;
assign n_873 = n_728 ^ n_714;
assign n_874 = n_701 ^ n_728;
assign n_875 = n_729 ^ n_317;
assign n_876 = n_393 ^ n_729;
assign n_877 = n_616 ^ n_731;
assign n_878 = n_279 ^ n_731;
assign n_879 = n_543 ^ n_731;
assign n_880 = n_343 ^ n_731;
assign n_881 = n_477 ^ n_731;
assign n_882 = n_732 ^ n_437;
assign n_883 = n_732 ^ n_489;
assign n_884 = ~n_734 & n_519;
assign n_885 = n_736 ^ n_437;
assign n_886 = n_737 ^ n_579;
assign n_887 = n_737 ^ n_731;
assign n_888 = n_485 & ~n_739;
assign n_889 = n_739 ^ n_274;
assign n_890 = n_352 ^ n_739;
assign n_891 = ~n_433 & n_739;
assign n_892 = n_739 ^ n_253;
assign n_893 = n_189 & n_739;
assign n_894 = n_213 & n_739;
assign n_895 = n_739 ^ n_273;
assign n_896 = ~n_273 & ~n_739;
assign n_897 = ~n_484 & n_739;
assign n_898 = n_739 ^ n_485;
assign n_899 = ~n_553 & n_739;
assign n_900 = n_294 ^ n_739;
assign n_901 = ~n_377 & n_739;
assign n_902 = n_739 ^ n_252;
assign n_903 = n_296 ^ n_739;
assign n_904 = n_739 ^ n_276;
assign n_905 = n_707 ^ n_739;
assign n_906 = n_27 & n_739;
assign n_907 = n_294 ^ n_740;
assign n_908 = ~n_484 & n_740;
assign n_909 = ~n_273 & ~n_740;
assign n_910 = ~n_534 & n_740;
assign n_911 = ~n_553 & n_740;
assign n_912 = ~n_485 & n_740;
assign n_913 = n_275 ^ n_740;
assign n_914 = n_213 ^ n_740;
assign n_915 = ~n_213 & ~n_740;
assign n_916 = n_189 & n_740;
assign n_917 = ~n_377 & n_740;
assign n_918 = n_433 & ~n_740;
assign n_919 = n_377 ^ n_740;
assign n_920 = n_253 ^ n_740;
assign n_921 = n_291 ^ n_740;
assign n_922 = n_274 ^ n_740;
assign n_923 = n_241 ^ n_740;
assign n_924 = n_272 & n_740;
assign n_925 = ~n_381 & n_740;
assign n_926 = n_250 ^ n_740;
assign n_927 = ~n_411 ^ ~n_740;
assign n_928 = n_741 ^ n_438;
assign n_929 = n_745 ^ n_558;
assign n_930 = n_749 ^ n_552;
assign n_931 = n_587 ^ n_749;
assign n_932 = n_751 ^ n_343;
assign n_933 = n_751 ^ n_317;
assign n_934 = n_752 ^ n_279;
assign n_935 = n_753 ^ n_419;
assign n_936 = n_754 ^ n_562;
assign n_937 = n_754 ^ n_596;
assign n_938 = ~n_712 ^ ~n_755;
assign n_939 = n_392 ^ n_757;
assign n_940 = n_368 ^ n_757;
assign n_941 = n_590 ^ n_757;
assign n_942 = n_589 ^ n_757;
assign n_943 = n_683 ^ n_757;
assign n_944 = n_758 ^ n_359;
assign n_945 = n_758 ^ n_488;
assign n_946 = ~n_596 ^ ~n_759;
assign n_947 = ~n_733 ^ ~n_761;
assign n_948 = n_763 ^ n_455;
assign n_949 = n_680 ^ n_763;
assign n_950 = n_699 ^ n_764;
assign n_951 = n_765 ^ n_366;
assign n_952 = n_766 ^ n_269;
assign n_953 = n_768 ^ n_636;
assign n_954 = n_770 ^ n_393;
assign n_955 = n_583 ^ n_772;
assign n_956 = ~n_773 ^ ~n_500;
assign n_957 = n_775 ^ n_437;
assign n_958 = ~n_778 & n_411;
assign n_959 = n_570 ^ n_778;
assign n_960 = n_514 ^ n_780;
assign n_961 = n_780 ^ n_533;
assign n_962 = n_781 ^ n_655;
assign n_963 = n_790 ^ n_354;
assign n_964 = n_791 ^ n_484;
assign n_965 = n_793 ^ n_420;
assign n_966 = n_794 ^ n_596;
assign n_967 = n_795 ^ n_317;
assign n_968 = ~n_795 ^ ~n_461;
assign n_969 = ~n_647 ^ ~n_797;
assign n_970 = ~n_738 ^ ~n_799;
assign n_971 = n_808 ^ n_281;
assign n_972 = n_809 ^ n_765;
assign n_973 = n_810 ^ n_513;
assign n_974 = n_648 ^ n_810;
assign n_975 = n_810 ^ n_572;
assign n_976 = ~n_811 ^ n_417;
assign n_977 = n_462 ^ n_811;
assign n_978 = n_405 ^ n_812;
assign n_979 = ~n_684 ^ ~n_813;
assign n_980 = ~n_811 ^ ~n_814;
assign n_981 = ~n_814 ^ ~n_769;
assign n_982 = n_815 ^ n_477;
assign n_983 = n_328 ^ n_815;
assign n_984 = n_816 ^ n_592;
assign n_985 = n_817 ^ n_593;
assign n_986 = n_819 ^ n_489;
assign n_987 = n_820 ^ n_285;
assign n_988 = n_715 ^ n_821;
assign n_989 = n_760 ^ n_822;
assign n_990 = n_823 ^ n_657;
assign n_991 = n_824 ^ n_652;
assign n_992 = ~n_825 ^ ~n_767;
assign n_993 = n_492 ^ n_825;
assign n_994 = ~n_828 ^ ~n_735;
assign n_995 = n_829 ^ n_571;
assign n_996 = n_830 ^ n_562;
assign n_997 = n_830 ^ n_533;
assign n_998 = n_832 ^ n_313;
assign n_999 = ~n_633 ^ ~n_833;
assign n_1000 = n_636 ^ n_836;
assign n_1001 = n_839 ^ n_535;
assign n_1002 = n_840 ^ n_626;
assign n_1003 = n_733 ^ n_843;
assign n_1004 = n_827 ^ n_844;
assign n_1005 = n_844 ^ n_622;
assign n_1006 = n_573 ^ n_844;
assign n_1007 = n_304 ^ n_845;
assign n_1008 = n_846 ^ n_354;
assign n_1009 = n_848 ^ n_562;
assign n_1010 = ~n_800 ^ n_851;
assign n_1011 = n_852 ^ n_343;
assign n_1012 = n_853 ^ n_685;
assign n_1013 = n_855 ^ n_695;
assign n_1014 = n_661 ^ n_855;
assign n_1015 = n_698 ^ n_858;
assign n_1016 = n_386 ^ n_859;
assign n_1017 = n_338 ^ n_859;
assign n_1018 = n_513 ^ n_859;
assign n_1019 = n_660 ^ n_859;
assign n_1020 = ~n_863 ^ ~n_782;
assign n_1021 = ~n_795 ^ ~n_863;
assign n_1022 = n_463 ^ n_867;
assign n_1023 = n_872 ^ n_286;
assign n_1024 = ~n_873 ^ ~n_659;
assign n_1025 = n_687 ^ n_874;
assign n_1026 = n_875 ^ n_688;
assign n_1027 = n_875 ^ n_717;
assign n_1028 = ~n_876 ^ n_520;
assign n_1029 = n_878 ^ n_291;
assign n_1030 = n_879 ^ n_757;
assign n_1031 = n_880 ^ n_484;
assign n_1032 = n_712 ^ n_880;
assign n_1033 = n_881 ^ n_673;
assign n_1034 = n_529 ^ n_882;
assign n_1035 = ~n_752 ^ ~n_885;
assign n_1036 = n_886 ^ n_336;
assign n_1037 = n_887 ^ n_628;
assign n_1038 = ~n_794 ^ ~n_887;
assign n_1039 = ~n_887 ^ ~n_716;
assign n_1040 = n_668 ^ n_888;
assign n_1041 = ~n_888 & n_376;
assign n_1042 = n_273 & n_889;
assign n_1043 = n_889 ^ n_297;
assign n_1044 = n_890 ^ n_276;
assign n_1045 = n_213 & n_890;
assign n_1046 = n_890 ^ n_274;
assign n_1047 = n_891 ^ n_459;
assign n_1048 = n_891 ^ n_601;
assign n_1049 = n_891 ^ n_675;
assign n_1050 = n_491 ^ n_891;
assign n_1051 = n_592 ^ n_891;
assign n_1052 = n_271 & n_892;
assign n_1053 = ~n_553 & n_892;
assign n_1054 = n_337 ^ n_892;
assign n_1055 = n_893 ^ n_354;
assign n_1056 = n_546 ^ n_893;
assign n_1057 = n_640 ^ n_893;
assign n_1058 = n_893 ^ n_307;
assign n_1059 = n_894 ^ n_286;
assign n_1060 = n_894 ^ n_605;
assign n_1061 = n_548 ^ n_894;
assign n_1062 = n_895 ^ n_896;
assign n_1063 = ~n_896 & ~n_379;
assign n_1064 = n_897 ^ n_730;
assign n_1065 = n_897 ^ n_622;
assign n_1066 = n_897 ^ n_683;
assign n_1067 = ~n_897 ^ ~n_773;
assign n_1068 = n_898 ^ n_888;
assign n_1069 = n_496 ^ n_899;
assign n_1070 = n_680 ^ n_899;
assign n_1071 = n_324 ^ n_899;
assign n_1072 = ~n_900 ^ ~n_609;
assign n_1073 = n_901 ^ n_438;
assign n_1074 = n_901 ^ n_439;
assign n_1075 = n_501 ^ n_901;
assign n_1076 = n_902 ^ n_295;
assign n_1077 = n_902 ^ n_292;
assign n_1078 = n_316 & ~n_902;
assign n_1079 = ~n_382 & n_903;
assign n_1080 = ~n_484 & n_903;
assign n_1081 = ~n_167 & n_904;
assign n_1082 = n_905 ^ n_901;
assign n_1083 = n_390 ^ n_906;
assign n_1084 = n_167 & n_907;
assign n_1085 = ~n_553 & n_907;
assign n_1086 = n_908 ^ n_533;
assign n_1087 = n_559 ^ n_908;
assign n_1088 = n_603 ^ n_908;
assign n_1089 = n_592 ^ n_908;
assign n_1090 = n_542 ^ n_908;
assign n_1091 = n_909 ^ n_510;
assign n_1092 = ~n_909 & ~n_507;
assign n_1093 = ~n_909 & n_748;
assign n_1094 = n_910 ^ n_616;
assign n_1095 = n_910 ^ n_438;
assign n_1096 = n_657 ^ n_910;
assign n_1097 = n_391 ^ n_910;
assign n_1098 = ~n_910 ^ ~n_528;
assign n_1099 = n_621 ^ n_911;
assign n_1100 = n_620 ^ n_911;
assign n_1101 = n_908 ^ n_911;
assign n_1102 = n_325 ^ n_911;
assign n_1103 = n_575 ^ n_912;
assign n_1104 = n_890 ^ n_913;
assign n_1105 = n_913 ^ n_843;
assign n_1106 = n_914 ^ n_915;
assign n_1107 = n_894 ^ n_915;
assign n_1108 = n_269 ^ n_916;
assign n_1109 = n_916 ^ n_552;
assign n_1110 = n_359 ^ n_916;
assign n_1111 = n_916 ^ n_622;
assign n_1112 = n_624 ^ n_916;
assign n_1113 = n_916 ^ n_358;
assign n_1114 = n_917 ^ n_689;
assign n_1115 = n_917 ^ n_589;
assign n_1116 = n_918 ^ n_271;
assign n_1117 = n_676 ^ n_918;
assign n_1118 = ~n_557 & ~n_918;
assign n_1119 = ~n_919 & n_857;
assign n_1120 = n_920 ^ n_295;
assign n_1121 = n_213 & n_920;
assign n_1122 = n_920 ^ n_370;
assign n_1123 = n_242 & n_921;
assign n_1124 = ~n_167 & n_922;
assign n_1125 = ~n_306 & n_922;
assign n_1126 = n_377 ^ ~n_923;
assign n_1127 = n_924 ^ n_628;
assign n_1128 = n_926 ^ n_297;
assign n_1129 = n_926 ^ n_216;
assign n_1130 = ~n_888 & n_927;
assign n_1131 = ~n_611 & ~n_928;
assign n_1132 = ~n_347 ^ n_930;
assign n_1133 = n_930 ^ n_434;
assign n_1134 = n_349 ^ n_930;
assign n_1135 = n_626 ^ n_930;
assign n_1136 = n_846 ^ n_930;
assign n_1137 = n_549 ^ n_933;
assign n_1138 = n_574 ^ n_934;
assign n_1139 = n_935 ^ n_294;
assign n_1140 = n_936 ^ n_674;
assign n_1141 = n_939 ^ n_323;
assign n_1142 = n_588 ^ n_940;
assign n_1143 = ~n_801 ^ ~n_941;
assign n_1144 = ~n_941 ^ n_868;
assign n_1145 = n_943 ^ n_676;
assign n_1146 = n_599 ^ n_944;
assign n_1147 = n_804 ^ n_945;
assign n_1148 = n_789 ^ n_948;
assign n_1149 = ~n_673 ^ ~n_952;
assign n_1150 = n_493 ^ n_958;
assign n_1151 = n_809 ^ n_958;
assign n_1152 = n_711 ^ n_958;
assign n_1153 = n_958 ^ n_683;
assign n_1154 = n_961 ^ n_543;
assign n_1155 = n_963 ^ n_552;
assign n_1156 = n_965 ^ n_859;
assign n_1157 = n_966 ^ n_486;
assign n_1158 = n_967 ^ n_285;
assign n_1159 = n_818 ^ n_973;
assign n_1160 = n_974 ^ n_309;
assign n_1161 = n_975 ^ n_958;
assign n_1162 = ~n_978 ^ ~n_806;
assign n_1163 = n_978 ^ n_563;
assign n_1164 = n_982 ^ n_653;
assign n_1165 = ~n_786 ^ ~n_983;
assign n_1166 = ~n_983 ^ ~n_864;
assign n_1167 = ~n_841 ^ ~n_984;
assign n_1168 = ~n_620 ^ ~n_985;
assign n_1169 = ~n_946 ^ n_986;
assign n_1170 = n_986 ^ n_340;
assign n_1171 = ~n_962 ^ n_988;
assign n_1172 = ~n_957 ^ n_989;
assign n_1173 = ~n_815 ^ ~n_990;
assign n_1174 = n_991 ^ n_627;
assign n_1175 = n_580 ^ n_991;
assign n_1176 = n_991 ^ n_908;
assign n_1177 = n_647 ^ n_991;
assign n_1178 = n_679 ^ n_991;
assign n_1179 = n_366 ^ n_991;
assign n_1180 = n_993 ^ n_534;
assign n_1181 = ~n_995 ^ ~n_403;
assign n_1182 = ~n_805 ^ ~n_996;
assign n_1183 = n_997 ^ n_859;
assign n_1184 = ~n_999 ^ ~n_931;
assign n_1185 = ~n_1001 ^ ~n_977;
assign n_1186 = ~n_1002 ^ ~n_865;
assign n_1187 = ~n_490 ^ n_1007;
assign n_1188 = n_1008 ^ n_244;
assign n_1189 = n_1008 ^ ~n_718;
assign n_1190 = ~n_878 ^ ~n_1009;
assign n_1191 = n_669 ^ n_1011;
assign n_1192 = ~n_768 ^ ~n_1013;
assign n_1193 = ~n_1015 ^ ~n_784;
assign n_1194 = n_1017 ^ n_396;
assign n_1195 = n_1018 ^ n_336;
assign n_1196 = n_1019 ^ ~n_723;
assign n_1197 = n_1019 ^ n_932;
assign n_1198 = ~n_992 ^ ~n_1025;
assign n_1199 = ~n_992 ^ ~n_1028;
assign n_1200 = n_987 ^ n_1029;
assign n_1201 = n_1030 ^ n_628;
assign n_1202 = n_576 ^ n_1030;
assign n_1203 = n_289 & n_1031;
assign n_1204 = ~n_946 ^ ~n_1033;
assign n_1205 = ~n_847 ^ ~n_1034;
assign n_1206 = n_1037 ^ n_623;
assign n_1207 = ~n_1038 ^ ~n_849;
assign n_1208 = ~n_532 & ~n_1040;
assign n_1209 = ~n_1041 ^ n_884;
assign n_1210 = n_1042 ^ n_859;
assign n_1211 = n_1043 & ~n_436;
assign n_1212 = n_307 & n_1044;
assign n_1213 = n_1045 ^ n_496;
assign n_1214 = ~n_433 & n_1046;
assign n_1215 = ~n_534 & n_1046;
assign n_1216 = n_1047 ^ n_675;
assign n_1217 = ~n_1047 ^ n_1006;
assign n_1218 = ~n_771 ^ ~n_1048;
assign n_1219 = n_1050 ^ n_268;
assign n_1220 = n_398 ^ n_1052;
assign n_1221 = n_1053 ^ n_558;
assign n_1222 = n_1053 ^ n_514;
assign n_1223 = ~n_485 & n_1054;
assign n_1224 = n_459 ^ n_1055;
assign n_1225 = n_677 ^ n_1055;
assign n_1226 = n_1055 ^ n_281;
assign n_1227 = n_1051 ^ n_1056;
assign n_1228 = ~n_1057 ^ ~n_744;
assign n_1229 = n_1059 ^ n_445;
assign n_1230 = n_1060 ^ n_333;
assign n_1231 = ~n_1060 ^ ~n_702;
assign n_1232 = ~n_1061 & ~n_404;
assign n_1233 = n_894 ^ n_1062;
assign n_1234 = n_463 ^ n_1062;
assign n_1235 = n_1063 & n_329;
assign n_1236 = n_1062 ^ n_1065;
assign n_1237 = n_1066 ^ n_378;
assign n_1238 = ~n_1067 ^ n_592;
assign n_1239 = n_729 ^ n_1068;
assign n_1240 = n_617 ^ n_1068;
assign n_1241 = n_677 ^ n_1068;
assign n_1242 = n_1068 ^ n_551;
assign n_1243 = n_776 ^ n_1068;
assign n_1244 = n_1068 ^ n_561;
assign n_1245 = n_336 ^ n_1068;
assign n_1246 = n_492 ^ n_1068;
assign n_1247 = n_1018 ^ n_1070;
assign n_1248 = ~n_1070 ^ ~n_524;
assign n_1249 = n_1071 ^ n_493;
assign n_1250 = n_1072 & ~n_707;
assign n_1251 = n_1073 ^ n_486;
assign n_1252 = n_1073 ^ n_697;
assign n_1253 = n_1074 ^ n_875;
assign n_1254 = n_1075 ^ n_697;
assign n_1255 = n_1076 & ~n_545;
assign n_1256 = n_484 & ~n_1077;
assign n_1257 = n_272 & ~n_1078;
assign n_1258 = ~n_377 & ~n_1078;
assign n_1259 = n_1079 ^ n_252;
assign n_1260 = n_1080 ^ n_492;
assign n_1261 = n_1081 ^ n_426;
assign n_1262 = ~n_632 & ~n_1082;
assign n_1263 = ~n_622 ^ ~n_1083;
assign n_1264 = ~n_388 & ~n_1084;
assign n_1265 = n_322 ^ n_1084;
assign n_1266 = n_1085 ^ n_774;
assign n_1267 = n_1086 ^ n_487;
assign n_1268 = ~n_641 ^ ~n_1087;
assign n_1269 = n_1089 ^ n_543;
assign n_1270 = n_1089 ^ n_572;
assign n_1271 = n_1090 ^ n_677;
assign n_1272 = n_1092 ^ n_324;
assign n_1273 = n_325 ^ n_1094;
assign n_1274 = ~n_1095 ^ n_1003;
assign n_1275 = n_830 ^ n_1095;
assign n_1276 = n_624 ^ n_1096;
assign n_1277 = n_506 ^ n_1096;
assign n_1278 = n_1097 ^ n_856;
assign n_1279 = ~n_530 ^ ~n_1098;
assign n_1280 = ~n_1099 ^ ~n_877;
assign n_1281 = n_692 ^ n_1100;
assign n_1282 = n_1023 ^ n_1101;
assign n_1283 = n_1103 ^ n_705;
assign n_1284 = ~n_377 & n_1104;
assign n_1285 = ~n_381 & ~n_1105;
assign n_1286 = n_1106 ^ n_643;
assign n_1287 = n_1106 ^ n_621;
assign n_1288 = n_677 ^ n_1106;
assign n_1289 = ~n_465 ^ ~n_1108;
assign n_1290 = n_1109 ^ n_489;
assign n_1291 = ~n_1109 ^ ~n_736;
assign n_1292 = n_1110 ^ n_674;
assign n_1293 = n_1111 ^ n_584;
assign n_1294 = n_1112 ^ n_502;
assign n_1295 = n_1114 ^ n_616;
assign n_1296 = n_1115 ^ n_437;
assign n_1297 = n_950 ^ n_1115;
assign n_1298 = n_1116 ^ n_919;
assign n_1299 = ~n_826 & n_1117;
assign n_1300 = n_1118 ^ n_1073;
assign n_1301 = n_740 ^ n_1119;
assign n_1302 = ~n_485 & n_1120;
assign n_1303 = n_1121 ^ n_397;
assign n_1304 = ~n_484 & n_1122;
assign n_1305 = ~n_1123 ^ ~n_838;
assign n_1306 = ~n_27 ^ ~n_1124;
assign n_1307 = n_1125 ^ n_739;
assign n_1308 = ~n_888 & n_1126;
assign n_1309 = n_189 & n_1128;
assign n_1310 = n_619 & n_1129;
assign n_1311 = ~n_811 ^ ~n_1130;
assign n_1312 = ~n_1132 & ~n_1091;
assign n_1313 = ~n_1133 ^ ~n_955;
assign n_1314 = n_1133 ^ n_419;
assign n_1315 = n_412 ^ n_1133;
assign n_1316 = ~n_1133 ^ ~n_684;
assign n_1317 = n_1134 ^ n_354;
assign n_1318 = n_1135 ^ n_366;
assign n_1319 = n_1136 ^ n_622;
assign n_1320 = ~n_951 ^ ~n_1138;
assign n_1321 = n_273 & n_1139;
assign n_1322 = ~n_953 ^ ~n_1140;
assign n_1323 = n_1145 ^ n_1047;
assign n_1324 = n_1145 ^ ~n_850;
assign n_1325 = n_971 ^ ~n_1147;
assign n_1326 = n_1148 ^ n_910;
assign n_1327 = ~n_847 ^ ~n_1149;
assign n_1328 = ~n_1149 ^ ~n_947;
assign n_1329 = ~n_1150 ^ ~n_796;
assign n_1330 = ~n_807 ^ ~n_1152;
assign n_1331 = n_1153 ^ n_1085;
assign n_1332 = n_1156 ^ ~n_954;
assign n_1333 = n_1005 ^ ~n_1157;
assign n_1334 = n_1163 ^ n_616;
assign n_1335 = n_294 & n_1164;
assign n_1336 = ~n_1166 ^ ~n_649;
assign n_1337 = n_1170 ^ n_312;
assign n_1338 = n_1170 ^ ~n_1020;
assign n_1339 = ~n_871 ^ ~n_1173;
assign n_1340 = n_1174 ^ n_693;
assign n_1341 = n_958 ^ n_1175;
assign n_1342 = ~n_1175 ^ ~n_976;
assign n_1343 = n_831 ^ n_1175;
assign n_1344 = n_899 ^ n_1176;
assign n_1345 = n_1177 ^ n_541;
assign n_1346 = n_1178 ^ n_677;
assign n_1347 = ~n_1180 & ~n_427;
assign n_1348 = ~n_1168 ^ ~n_1181;
assign n_1349 = n_1183 ^ n_787;
assign n_1350 = ~n_1184 ^ ~n_803;
assign n_1351 = ~n_834 ^ ~n_1187;
assign n_1352 = ~n_981 ^ n_1188;
assign n_1353 = ~n_860 ^ ~n_1189;
assign n_1354 = ~n_1192 ^ ~n_1039;
assign n_1355 = ~n_527 ^ n_1194;
assign n_1356 = n_1195 ^ n_862;
assign n_1357 = ~n_1182 ^ ~n_1197;
assign n_1358 = ~n_1200 ^ ~n_1024;
assign n_1359 = ~n_841 ^ ~n_1202;
assign n_1360 = ~n_1073 ^ ~n_1203;
assign n_1361 = ~n_530 ^ ~n_1205;
assign n_1362 = n_1208 ^ n_353;
assign n_1363 = ~n_1208 ^ ~n_547;
assign n_1364 = ~n_1209 ^ ~n_861;
assign n_1365 = ~n_1211 ^ ~n_1047;
assign n_1366 = ~n_1213 ^ ~n_578;
assign n_1367 = ~n_1214 ^ n_1154;
assign n_1368 = ~n_1215 ^ ~n_869;
assign n_1369 = n_1216 ^ n_596;
assign n_1370 = ~n_1218 ^ ~n_727;
assign n_1371 = ~n_852 ^ ~n_1219;
assign n_1372 = ~n_1220 ^ ~n_1141;
assign n_1373 = ~n_1220 ^ ~n_658;
assign n_1374 = n_1221 ^ n_539;
assign n_1375 = n_1014 ^ n_1222;
assign n_1376 = n_1224 ^ n_912;
assign n_1377 = ~n_1102 ^ ~n_1225;
assign n_1378 = ~n_663 & ~n_1227;
assign n_1379 = ~n_1228 ^ ~n_1204;
assign n_1380 = n_1230 ^ n_622;
assign n_1381 = ~n_1231 ^ n_783;
assign n_1382 = n_1233 ^ n_897;
assign n_1383 = n_473 ^ n_1234;
assign n_1384 = ~n_290 ^ ~n_1235;
assign n_1385 = n_1237 ^ n_901;
assign n_1386 = n_719 ^ n_1238;
assign n_1387 = ~n_871 ^ ~n_1239;
assign n_1388 = n_544 ^ n_1239;
assign n_1389 = ~n_978 ^ ~n_1240;
assign n_1390 = ~n_1219 ^ ~n_1241;
assign n_1391 = n_1241 ^ n_473;
assign n_1392 = ~n_1241 ^ ~n_655;
assign n_1393 = n_1242 ^ n_605;
assign n_1394 = ~n_1181 ^ ~n_1243;
assign n_1395 = n_1244 ^ n_645;
assign n_1396 = n_792 ^ n_1246;
assign n_1397 = n_1247 ^ n_669;
assign n_1398 = ~n_1248 ^ n_1032;
assign n_1399 = ~n_1093 ^ ~n_1249;
assign n_1400 = ~n_785 ^ ~n_1249;
assign n_1401 = n_1049 ^ n_1251;
assign n_1402 = ~n_746 ^ ~n_1252;
assign n_1403 = n_883 ^ n_1253;
assign n_1404 = n_1254 ^ n_244;
assign n_1405 = ~n_636 ^ ~n_1255;
assign n_1406 = ~n_1256 & n_1257;
assign n_1407 = n_1258 ^ n_496;
assign n_1408 = n_942 ^ n_1260;
assign n_1409 = n_1261 & n_1058;
assign n_1410 = n_1262 ^ n_563;
assign n_1411 = ~n_753 & ~n_1263;
assign n_1412 = n_213 & ~n_1264;
assign n_1413 = n_307 & n_1265;
assign n_1414 = n_1267 ^ n_308;
assign n_1415 = ~n_1268 ^ ~n_1159;
assign n_1416 = n_1269 ^ n_674;
assign n_1417 = ~n_777 ^ ~n_1270;
assign n_1418 = n_1191 ^ ~n_1272;
assign n_1419 = ~n_1272 ^ ~n_1226;
assign n_1420 = n_1273 ^ n_1106;
assign n_1421 = n_1276 ^ n_1011;
assign n_1422 = n_566 ^ n_1276;
assign n_1423 = n_1277 ^ n_385;
assign n_1424 = ~n_1201 ^ ~n_1278;
assign n_1425 = ~n_976 ^ ~n_1279;
assign n_1426 = ~n_1280 ^ ~n_980;
assign n_1427 = ~n_1281 ^ ~n_661;
assign n_1428 = ~n_1284 ^ ~n_1146;
assign n_1429 = n_1286 ^ n_824;
assign n_1430 = n_1286 ^ n_893;
assign n_1431 = n_709 ^ n_1286;
assign n_1432 = n_1286 ^ n_910;
assign n_1433 = n_949 ^ n_1287;
assign n_1434 = n_1288 ^ n_434;
assign n_1435 = n_1288 ^ ~n_756;
assign n_1436 = n_1290 ^ n_539;
assign n_1437 = ~n_1291 ^ ~n_972;
assign n_1438 = ~n_508 ^ ~n_1292;
assign n_1439 = ~n_1293 & ~n_1294;
assign n_1440 = ~n_994 ^ ~n_1294;
assign n_1441 = n_1295 ^ n_654;
assign n_1442 = n_1296 ^ n_384;
assign n_1443 = n_990 ^ n_1296;
assign n_1444 = n_1296 ^ n_605;
assign n_1445 = n_1298 ^ n_562;
assign n_1446 = n_1133 ^ n_1298;
assign n_1447 = n_1298 ^ n_505;
assign n_1448 = n_324 ^ n_1298;
assign n_1449 = n_591 ^ n_1298;
assign n_1450 = n_677 ^ n_1298;
assign n_1451 = n_491 ^ n_1298;
assign n_1452 = n_626 ^ n_1298;
assign n_1453 = ~n_278 ^ ~n_1301;
assign n_1454 = n_1302 ^ n_395;
assign n_1455 = ~n_1302 ^ ~n_1165;
assign n_1456 = ~n_679 ^ ~n_1303;
assign n_1457 = ~n_1304 ^ ~n_471;
assign n_1458 = n_1306 & n_1307;
assign n_1459 = ~n_1308 ^ ~n_1036;
assign n_1460 = n_1145 ^ ~n_1309;
assign n_1461 = ~n_1310 ^ n_788;
assign n_1462 = ~n_968 ^ ~n_1311;
assign n_1463 = ~n_1312 ^ ~n_1094;
assign n_1464 = ~n_1111 ^ ~n_1313;
assign n_1465 = n_1314 ^ n_726;
assign n_1466 = n_925 ^ n_1315;
assign n_1467 = ~n_1316 ^ ~n_692;
assign n_1468 = ~n_1317 ^ ~n_747;
assign n_1469 = ~n_670 ^ ~n_1318;
assign n_1470 = ~n_1320 ^ ~n_866;
assign n_1471 = ~n_1021 ^ n_1323;
assign n_1472 = n_1326 ^ n_579;
assign n_1473 = ~n_1230 ^ ~n_1328;
assign n_1474 = ~n_1329 ^ ~n_1001;
assign n_1475 = ~n_1330 ^ ~n_1088;
assign n_1476 = ~n_1297 ^ ~n_1331;
assign n_1477 = n_802 ^ n_1337;
assign n_1478 = ~n_911 ^ ~n_1340;
assign n_1479 = ~n_1340 ^ ~n_1223;
assign n_1480 = ~n_606 ^ ~n_1341;
assign n_1481 = ~n_1184 ^ ~n_1342;
assign n_1482 = ~n_828 ^ ~n_1343;
assign n_1483 = n_1016 ^ ~n_1344;
assign n_1484 = n_618 ^ n_1344;
assign n_1485 = n_1345 ^ n_551;
assign n_1486 = n_1346 ^ n_477;
assign n_1487 = ~n_307 ^ ~n_1347;
assign n_1488 = ~n_1327 & ~n_1348;
assign n_1489 = ~n_1137 ^ n_1349;
assign n_1490 = ~n_1352 ^ ~n_1338;
assign n_1491 = ~n_1218 ^ ~n_1355;
assign n_1492 = ~n_938 ^ n_1356;
assign n_1493 = ~n_1357 ^ ~n_464;
assign n_1494 = ~n_1362 ^ n_1283;
assign n_1495 = ~n_1363 ^ n_1319;
assign n_1496 = ~n_1365 ^ ~n_1266;
assign n_1497 = ~n_1366 ^ ~n_1275;
assign n_1498 = n_1283 ^ ~n_1367;
assign n_1499 = ~n_1368 ^ ~n_1217;
assign n_1500 = ~n_1190 ^ ~n_1369;
assign n_1501 = ~n_1250 & ~n_1370;
assign n_1502 = ~n_499 ^ ~n_1371;
assign n_1503 = ~n_1372 ^ ~n_1000;
assign n_1504 = ~n_1373 & ~n_637;
assign n_1505 = ~n_1373 ^ ~n_1010;
assign n_1506 = ~n_785 ^ ~n_1376;
assign n_1507 = ~n_1377 ^ ~n_1161;
assign n_1508 = ~n_1380 ^ ~n_860;
assign n_1509 = ~n_1249 ^ ~n_1381;
assign n_1510 = n_1100 ^ n_1382;
assign n_1511 = n_1382 ^ n_1177;
assign n_1512 = n_1107 ^ n_1382;
assign n_1513 = n_750 ^ n_1382;
assign n_1514 = ~n_1383 ^ ~n_1305;
assign n_1515 = ~n_1383 ^ ~n_1300;
assign n_1516 = n_1385 ^ n_696;
assign n_1517 = n_1386 ^ ~n_864;
assign n_1518 = ~n_1388 ^ ~n_602;
assign n_1519 = ~n_1388 ^ ~n_1035;
assign n_1520 = ~n_595 ^ n_1391;
assign n_1521 = n_1395 ^ n_338;
assign n_1522 = ~n_1396 ^ ~n_1354;
assign n_1523 = ~n_1398 ^ ~n_1377;
assign n_1524 = ~n_854 ^ ~n_1399;
assign n_1525 = n_1401 ^ n_836;
assign n_1526 = ~n_1401 ^ ~n_659;
assign n_1527 = ~n_1402 ^ ~n_1322;
assign n_1528 = ~n_1402 ^ ~n_1339;
assign n_1529 = ~n_1402 ^ ~n_618;
assign n_1530 = ~n_1185 ^ ~n_1403;
assign n_1531 = ~n_1179 ^ ~n_1404;
assign n_1532 = ~n_1405 ^ ~n_1390;
assign n_1533 = ~n_798 ^ ~n_1406;
assign n_1534 = ~n_873 ^ ~n_1408;
assign n_1535 = ~n_622 ^ ~n_1409;
assign n_1536 = n_515 ^ n_1412;
assign n_1537 = ~n_1272 ^ ~n_1412;
assign n_1538 = n_1413 ^ n_673;
assign n_1539 = ~n_1413 ^ n_998;
assign n_1540 = ~n_509 ^ ~n_1414;
assign n_1541 = ~n_1415 ^ ~n_1358;
assign n_1542 = ~n_1408 ^ ~n_1416;
assign n_1543 = n_1142 ^ n_1420;
assign n_1544 = n_1421 ^ ~n_1369;
assign n_1545 = n_1422 ^ n_491;
assign n_1546 = ~n_1400 ^ ~n_1423;
assign n_1547 = ~n_1351 & ~n_1425;
assign n_1548 = ~n_1426 ^ ~n_861;
assign n_1549 = ~n_717 ^ n_1429;
assign n_1550 = n_1430 ^ n_897;
assign n_1551 = ~n_956 ^ n_1431;
assign n_1552 = n_1005 ^ n_1432;
assign n_1553 = n_1432 ^ ~n_1332;
assign n_1554 = ~n_1424 ^ n_1433;
assign n_1555 = n_1434 ^ ~n_1206;
assign n_1556 = ~n_781 ^ ~n_1435;
assign n_1557 = n_1436 ^ n_1064;
assign n_1558 = ~n_1438 ^ ~n_1069;
assign n_1559 = n_1439 ^ n_1282;
assign n_1560 = ~n_1441 ^ ~n_1299;
assign n_1561 = n_1442 ^ n_343;
assign n_1562 = ~n_1442 ^ ~n_1394;
assign n_1563 = n_842 ^ ~n_1443;
assign n_1564 = n_1127 ^ n_1444;
assign n_1565 = n_1445 ^ n_285;
assign n_1566 = n_831 ^ n_1445;
assign n_1567 = n_1446 ^ n_581;
assign n_1568 = ~n_1149 ^ ~n_1447;
assign n_1569 = ~n_781 ^ ~n_1448;
assign n_1570 = n_1448 ^ n_472;
assign n_1571 = n_664 ^ n_1449;
assign n_1572 = n_650 ^ n_1450;
assign n_1573 = n_1451 ^ n_897;
assign n_1574 = n_1452 ^ n_493;
assign n_1575 = ~n_1362 ^ ~n_1454;
assign n_1576 = ~n_1456 ^ ~n_964;
assign n_1577 = ~n_1457 ^ ~n_762;
assign n_1578 = ~n_1393 ^ ~n_1458;
assign n_1579 = ~n_1459 ^ ~n_870;
assign n_1580 = ~n_1270 & ~n_1461;
assign n_1581 = ~n_1464 ^ ~n_1375;
assign n_1582 = ~n_1196 ^ ~n_1466;
assign n_1583 = ~n_694 ^ ~n_1468;
assign n_1584 = ~n_1469 ^ ~n_1384;
assign n_1585 = n_904 & n_1471;
assign n_1586 = ~n_1472 ^ ~n_929;
assign n_1587 = ~n_1472 ^ ~n_992;
assign n_1588 = ~n_1020 ^ ~n_1475;
assign n_1589 = ~n_1360 ^ n_1477;
assign n_1590 = ~n_1479 ^ ~n_979;
assign n_1591 = ~n_1164 ^ ~n_1480;
assign n_1592 = ~n_1209 ^ ~n_1482;
assign n_1593 = ~n_1483 ^ n_971;
assign n_1594 = ~n_970 ^ ~n_1484;
assign n_1595 = ~n_711 ^ ~n_1485;
assign n_1596 = n_1485 ^ n_488;
assign n_1597 = ~n_1407 ^ ~n_1486;
assign n_1598 = n_1487 & n_1259;
assign n_1599 = ~n_615 ^ n_1488;
assign n_1600 = ~n_1491 ^ ~n_1237;
assign n_1601 = ~n_1492 ^ ~n_1162;
assign n_1602 = ~n_434 ^ ~n_1493;
assign n_1603 = ~n_1471 ^ ~n_1495;
assign n_1604 = ~n_1192 ^ ~n_1497;
assign n_1605 = ~n_1402 ^ ~n_1499;
assign n_1606 = ~n_1502 ^ ~n_1172;
assign n_1607 = ~n_1503 ^ ~n_1506;
assign n_1608 = ~n_1324 ^ ~n_1507;
assign n_1609 = n_1397 ^ ~n_1508;
assign n_1610 = ~n_1428 & ~n_1509;
assign n_1611 = ~n_1026 ^ n_1510;
assign n_1612 = n_1511 ^ n_672;
assign n_1613 = n_1012 ^ n_1513;
assign n_1614 = ~n_1514 ^ n_1378;
assign n_1615 = ~n_1514 ^ ~n_1350;
assign n_1616 = ~n_1515 ^ ~n_1396;
assign n_1617 = ~n_1207 ^ ~n_1516;
assign n_1618 = ~n_1342 ^ ~n_1517;
assign n_1619 = ~n_871 ^ ~n_1518;
assign n_1620 = ~n_1021 ^ ~n_1519;
assign n_1621 = ~n_1520 ^ ~n_1419;
assign n_1622 = ~n_1521 ^ ~n_1410;
assign n_1623 = ~n_1523 ^ ~n_1473;
assign n_1624 = ~n_1524 ^ ~n_1417;
assign n_1625 = ~n_1321 ^ ~n_1525;
assign n_1626 = ~n_1153 ^ ~n_1526;
assign n_1627 = ~n_1333 ^ ~n_1529;
assign n_1628 = ~n_1193 ^ ~n_1531;
assign n_1629 = ~n_1531 ^ ~n_1144;
assign n_1630 = ~n_1532 ^ ~n_1143;
assign n_1631 = ~n_1464 ^ ~n_1533;
assign n_1632 = ~n_1535 ^ ~n_1453;
assign n_1633 = n_1210 ^ ~n_1536;
assign n_1634 = ~n_1474 ^ ~n_1537;
assign n_1635 = ~n_1538 ^ ~n_1496;
assign n_1636 = ~n_1538 ^ ~n_1478;
assign n_1637 = ~n_1539 ^ ~n_1392;
assign n_1638 = ~n_1540 ^ ~n_1463;
assign n_1639 = ~n_1540 ^ ~n_1274;
assign n_1640 = ~n_462 ^ ~n_1543;
assign n_1641 = ~n_1489 ^ ~n_1544;
assign n_1642 = n_1374 ^ n_1545;
assign n_1643 = ~n_1347 ^ ~n_1549;
assign n_1644 = n_960 ^ n_1550;
assign n_1645 = ~n_1351 ^ ~n_1553;
assign n_1646 = n_534 & ~n_1554;
assign n_1647 = ~n_1555 ^ ~n_835;
assign n_1648 = ~n_1556 ^ ~n_1300;
assign n_1649 = ~n_1200 ^ ~n_1558;
assign n_1650 = ~n_1558 & ~n_1199;
assign n_1651 = ~n_1559 ^ ~n_1481;
assign n_1652 = ~n_1560 ^ ~n_1437;
assign n_1653 = n_1433 ^ n_1561;
assign n_1654 = ~n_1494 ^ ~n_1563;
assign n_1655 = n_1565 ^ n_1236;
assign n_1656 = ~n_1566 ^ ~n_1022;
assign n_1657 = n_872 ^ ~n_1567;
assign n_1658 = ~n_1568 ^ n_1561;
assign n_1659 = ~n_1569 ^ ~n_1155;
assign n_1660 = ~n_1570 ^ n_1411;
assign n_1661 = ~n_1057 ^ ~n_1571;
assign n_1662 = ~n_1572 ^ ~n_1158;
assign n_1663 = ~n_1572 ^ ~n_779;
assign n_1664 = n_1245 ^ n_1573;
assign n_1665 = ~n_941 ^ ~n_1574;
assign n_1666 = ~n_742 ^ ~n_1575;
assign n_1667 = ~n_1325 ^ ~n_1576;
assign n_1668 = ~n_1576 ^ ~n_1460;
assign n_1669 = ~n_1293 ^ ~n_1577;
assign n_1670 = ~n_1577 & n_1131;
assign n_1671 = ~n_1540 ^ ~n_1578;
assign n_1672 = ~n_1182 ^ ~n_1579;
assign n_1673 = ~n_1212 ^ n_1580;
assign n_1674 = ~n_1583 ^ ~n_1359;
assign n_1675 = ~n_1583 ^ ~n_1186;
assign n_1676 = ~n_1584 ^ ~n_1160;
assign n_1677 = ~n_1585 ^ ~n_671;
assign n_1678 = ~n_1169 ^ ~n_1586;
assign n_1679 = ~n_1587 ^ ~n_1387;
assign n_1680 = ~n_1455 & ~n_1590;
assign n_1681 = ~n_1591 ^ ~n_1350;
assign n_1682 = ~n_911 ^ ~n_1591;
assign n_1683 = ~n_1582 ^ ~n_1592;
assign n_1684 = ~n_1591 & ~n_1593;
assign n_1685 = ~n_1594 ^ ~n_1028;
assign n_1686 = n_1596 ^ n_948;
assign n_1687 = n_1397 ^ ~n_1597;
assign n_1688 = ~n_349 ^ ~n_1598;
assign n_1689 = ~n_1470 & ~n_1603;
assign n_1690 = n_672 ^ ~n_1604;
assign n_1691 = ~n_1325 ^ ~n_1605;
assign n_1692 = ~n_1426 & ~n_1607;
assign n_1693 = ~n_1608 ^ ~n_1500;
assign n_1694 = ~n_1608 ^ ~n_1546;
assign n_1695 = ~n_1335 ^ ~n_1609;
assign n_1696 = n_1488 & n_1610;
assign n_1697 = ~n_1611 ^ n_837;
assign n_1698 = ~n_1612 ^ ~n_1167;
assign n_1699 = ~n_1554 ^ ~n_1613;
assign n_1700 = ~n_1616 ^ ~n_1476;
assign n_1701 = ~n_1619 ^ ~n_1548;
assign n_1702 = ~n_1171 & ~n_1621;
assign n_1703 = ~n_1622 ^ ~n_1564;
assign n_1704 = ~n_1590 ^ ~n_1624;
assign n_1705 = ~n_1626 ^ ~n_1462;
assign n_1706 = ~n_1622 ^ ~n_1627;
assign n_1707 = ~n_1631 & ~n_1285;
assign n_1708 = ~n_1415 ^ ~n_1632;
assign n_1709 = ~n_1208 & ~n_1633;
assign n_1710 = ~n_1557 ^ ~n_1634;
assign n_1711 = ~n_1638 ^ ~n_1635;
assign n_1712 = ~n_1638 & n_1504;
assign n_1713 = ~n_1173 ^ ~n_1640;
assign n_1714 = ~n_1171 ^ ~n_1642;
assign n_1715 = ~n_490 ^ ~n_1642;
assign n_1716 = n_553 ^ ~n_1643;
assign n_1717 = ~n_1643 & ~n_1527;
assign n_1718 = ~n_1644 ^ ~n_1364;
assign n_1719 = ~n_1618 ^ ~n_1645;
assign n_1720 = ~n_1646 & n_1512;
assign n_1721 = ~n_1647 ^ ~n_1534;
assign n_1722 = ~n_1160 ^ ~n_1648;
assign n_1723 = n_253 & n_1648;
assign n_1724 = ~n_1649 & ~n_1625;
assign n_1725 = ~n_1651 ^ ~n_1630;
assign n_1726 = ~n_1652 ^ ~n_1628;
assign n_1727 = ~n_1653 ^ ~n_1581;
assign n_1728 = ~n_1654 ^ ~n_1595;
assign n_1729 = ~n_1114 ^ n_1655;
assign n_1730 = ~n_1656 ^ ~n_1389;
assign n_1731 = ~n_1633 ^ ~n_1657;
assign n_1732 = ~n_1657 & ~n_1490;
assign n_1733 = ~n_1527 ^ ~n_1658;
assign n_1734 = ~n_1528 ^ ~n_1659;
assign n_1735 = ~n_1660 ^ ~n_1440;
assign n_1736 = ~n_1606 & ~n_1661;
assign n_1737 = ~n_1661 ^ ~n_1232;
assign n_1738 = ~n_1551 ^ ~n_1662;
assign n_1739 = ~n_1165 ^ ~n_1663;
assign n_1740 = ~n_863 ^ ~n_1664;
assign n_1741 = ~n_1427 ^ ~n_1665;
assign n_1742 = ~n_1666 ^ ~n_994;
assign n_1743 = ~n_1668 ^ ~n_1027;
assign n_1744 = ~n_1669 ^ ~n_1637;
assign n_1745 = ~n_1631 & n_1670;
assign n_1746 = ~n_1667 & ~n_1671;
assign n_1747 = ~n_1672 ^ ~n_854;
assign n_1748 = ~n_1618 ^ ~n_1674;
assign n_1749 = ~n_1675 ^ ~n_1552;
assign n_1750 = ~n_1676 ^ ~n_1601;
assign n_1751 = ~n_1678 ^ ~n_969;
assign n_1752 = ~n_1679 ^ ~n_1557;
assign n_1753 = ~n_1682 ^ ~n_1498;
assign n_1754 = ~n_1198 ^ n_1686;
assign n_1755 = ~n_1688 ^ n_1547;
assign n_1756 = ~n_1469 ^ ~n_1693;
assign n_1757 = ~n_992 ^ ~n_1695;
assign n_1758 = ~n_1697 ^ ~n_1428;
assign n_1759 = ~n_1697 ^ ~n_1328;
assign n_1760 = ~n_1698 ^ n_1421;
assign n_1761 = ~n_1554 & ~n_1700;
assign n_1762 = ~n_1701 ^ ~n_1629;
assign n_1763 = ~n_1676 ^ n_1702;
assign n_1764 = ~n_1336 & ~n_1703;
assign n_1765 = ~n_1677 ^ ~n_1704;
assign n_1766 = ~n_1706 ^ ~n_1681;
assign n_1767 = ~n_1687 & n_1707;
assign n_1768 = ~n_1589 ^ ~n_1708;
assign n_1769 = n_1709 ^ ~n_1212;
assign n_1770 = n_1709 ^ ~n_1639;
assign n_1771 = n_1709 ^ ~n_1289;
assign n_1772 = ~n_1710 & ~n_1701;
assign n_1773 = n_165 & ~n_1712;
assign n_1774 = n_273 & n_1712;
assign n_1775 = n_163 & ~n_1712;
assign n_1776 = ~n_145 & ~n_1712;
assign n_1777 = ~n_111 & ~n_1712;
assign n_1778 = ~n_112 & ~n_1712;
assign n_1779 = ~n_100 & ~n_1712;
assign n_1780 = n_90 & ~n_1712;
assign n_1781 = ~n_103 & ~n_1712;
assign n_1782 = n_100 ^ n_1712;
assign n_1783 = n_87 ^ n_1712;
assign n_1784 = ~n_87 & n_1712;
assign n_1785 = ~n_74 & ~n_1712;
assign n_1786 = ~n_88 & ~n_1712;
assign n_1787 = n_88 ^ n_1712;
assign n_1788 = n_135 & ~n_1712;
assign n_1789 = ~n_235 & ~n_1712;
assign n_1790 = n_263 & ~n_1712;
assign n_1791 = ~n_233 & ~n_1712;
assign n_1792 = ~n_1113 ^ n_1712;
assign n_1793 = ~n_1320 ^ ~n_1713;
assign n_1794 = ~n_1600 & ~n_1714;
assign n_1795 = n_1716 & ~n_959;
assign n_1796 = ~n_1599 ^ ~n_1720;
assign n_1797 = ~n_1379 ^ ~n_1720;
assign n_1798 = ~n_742 ^ ~n_1721;
assign n_1799 = ~n_1722 ^ ~n_1685;
assign n_1800 = ~n_1723 ^ ~n_1694;
assign n_1801 = ~n_1602 ^ ~n_1726;
assign n_1802 = ~n_1591 ^ ~n_1727;
assign n_1803 = ~n_1728 ^ ~n_1699;
assign n_1804 = ~n_1728 & ~n_1715;
assign n_1805 = ~n_1361 ^ ~n_1729;
assign n_1806 = ~n_1729 ^ ~n_1542;
assign n_1807 = ~n_1455 ^ ~n_1730;
assign n_1808 = ~n_1418 & ~n_1731;
assign n_1809 = ~n_1733 & ~n_1673;
assign n_1810 = ~n_1734 ^ ~n_1683;
assign n_1811 = ~n_1734 ^ ~n_1685;
assign n_1812 = ~n_1734 & ~n_1614;
assign n_1813 = ~n_1530 ^ ~n_1735;
assign n_1814 = ~n_1688 ^ n_1736;
assign n_1815 = ~n_1737 ^ ~n_1353;
assign n_1816 = ~n_1615 & ~n_1738;
assign n_1817 = ~n_1739 ^ ~n_1522;
assign n_1818 = ~n_1740 ^ ~n_1137;
assign n_1819 = ~n_1415 ^ ~n_1741;
assign n_1820 = ~n_1743 ^ n_1680;
assign n_1821 = x1 & ~n_1745;
assign n_1822 = n_22 & n_1745;
assign n_1823 = ~n_199 & ~n_1745;
assign n_1824 = ~n_226 & ~n_1745;
assign n_1825 = n_87 ^ n_1745;
assign n_1826 = n_157 ^ n_1745;
assign n_1827 = n_531 & ~n_1745;
assign n_1828 = n_159 & ~n_1745;
assign n_1829 = n_98 & ~n_1745;
assign n_1830 = n_144 ^ n_1745;
assign n_1831 = ~n_231 & ~n_1745;
assign n_1832 = n_121 ^ n_1745;
assign n_1833 = n_197 & ~n_1745;
assign n_1834 = n_198 & ~n_1745;
assign n_1835 = n_165 ^ n_1745;
assign n_1836 = ~n_375 & ~n_1745;
assign n_1837 = ~n_165 & n_1745;
assign n_1838 = n_164 & ~n_1745;
assign n_1839 = n_236 & ~n_1745;
assign n_1840 = ~n_187 & n_1745;
assign n_1841 = ~n_1651 ^ ~n_1747;
assign n_1842 = ~n_1749 & ~n_1739;
assign n_1843 = ~n_1697 ^ ~n_1750;
assign n_1844 = ~n_328 ^ ~n_1751;
assign n_1845 = ~n_1752 ^ n_1684;
assign n_1846 = ~n_1753 ^ ~n_1617;
assign n_1847 = ~n_1754 ^ ~n_1465;
assign n_1848 = n_678 & n_1755;
assign n_1849 = ~n_1757 ^ ~n_1151;
assign n_1850 = ~n_1759 ^ ~n_1562;
assign n_1851 = ~n_1760 ^ ~n_1588;
assign n_1852 = ~n_1760 & n_1724;
assign n_1853 = ~n_1493 & n_1761;
assign n_1854 = ~n_1757 & ~n_1762;
assign n_1855 = ~n_1742 ^ ~n_1763;
assign n_1856 = ~n_1530 ^ n_1764;
assign n_1857 = ~n_1721 & ~n_1765;
assign n_1858 = ~n_1766 & ~n_1623;
assign n_1859 = ~n_675 ^ ~n_1769;
assign n_1860 = ~n_1769 & ~n_1711;
assign n_1861 = n_1692 & ~n_1770;
assign n_1862 = n_484 & n_1772;
assign n_1863 = n_1773 ^ n_165;
assign n_1864 = ~n_1774 & ~n_1636;
assign n_1865 = n_1777 ^ n_1712;
assign n_1866 = n_1777 ^ n_111;
assign n_1867 = n_1783 ^ n_1784;
assign n_1868 = n_74 ^ n_1784;
assign n_1869 = n_1785 ^ n_1712;
assign n_1870 = ~n_1758 & ~n_1793;
assign n_1871 = ~n_1733 ^ n_1794;
assign n_1872 = ~n_1795 ^ n_1501;
assign n_1873 = ~n_888 & n_1796;
assign n_1874 = ~n_1796 & ~n_1725;
assign n_1875 = ~n_1797 ^ n_1732;
assign n_1876 = n_216 & n_1797;
assign n_1877 = ~n_1688 ^ ~n_1802;
assign n_1878 = ~n_1803 & ~n_1541;
assign n_1879 = ~n_1691 ^ n_1804;
assign n_1880 = ~n_1805 ^ ~n_1705;
assign n_1881 = ~n_1806 ^ ~n_1620;
assign n_1882 = ~n_1806 ^ ~n_1641;
assign n_1883 = ~n_1652 ^ ~n_1807;
assign n_1884 = n_1808 & ~n_1470;
assign n_1885 = ~n_1753 & n_1809;
assign n_1886 = ~n_1810 ^ ~n_1715;
assign n_1887 = n_1689 & ~n_1811;
assign n_1888 = ~n_1755 & n_1812;
assign n_1889 = ~n_1728 ^ ~n_1813;
assign n_1890 = ~n_1814 ^ n_1767;
assign n_1891 = ~n_1814 ^ ~n_937;
assign n_1892 = ~n_1815 ^ ~n_1334;
assign n_1893 = ~n_1651 ^ ~n_1817;
assign n_1894 = ~n_1632 ^ ~n_1818;
assign n_1895 = ~n_1819 ^ n_1650;
assign n_1896 = ~n_1623 & ~n_1820;
assign n_1897 = n_122 & ~n_1832;
assign n_1898 = n_163 & n_1835;
assign n_1899 = ~n_184 & n_1837;
assign n_1900 = ~n_186 & ~n_1838;
assign n_1901 = n_164 & ~n_1839;
assign n_1902 = n_1840 ^ n_187;
assign n_1903 = ~n_1797 & ~n_1841;
assign n_1904 = ~n_1602 ^ n_1842;
assign n_1905 = ~n_1844 ^ n_1746;
assign n_1906 = ~n_1845 & ~n_1805;
assign n_1907 = ~n_1847 & n_1772;
assign n_1908 = ~n_1847 ^ ~n_1229;
assign n_1909 = ~n_1849 & ~n_1748;
assign n_1910 = ~n_1849 & n_1816;
assign n_1911 = ~n_1850 & n_1717;
assign n_1912 = ~n_1851 & ~n_1798;
assign n_1913 = ~n_1742 & n_1852;
assign n_1914 = ~n_1677 & n_1853;
assign n_1915 = ~n_1742 & ~n_1856;
assign n_1916 = ~n_1859 ^ ~n_1505;
assign n_1917 = ~n_1859 ^ ~n_1792;
assign n_1918 = ~n_1082 & ~n_1862;
assign n_1919 = n_1863 ^ n_145;
assign n_1920 = n_207 & n_1864;
assign n_1921 = n_1712 ^ n_1864;
assign n_1922 = n_1712 ^ n_1864;
assign n_1923 = n_135 & n_1864;
assign n_1924 = ~n_103 ^ n_1864;
assign n_1925 = n_74 ^ n_1864;
assign n_1926 = ~n_187 & n_1864;
assign n_1927 = ~n_1771 & n_1864;
assign n_1928 = n_1866 ^ n_103;
assign n_1929 = ~n_1868 & n_1864;
assign n_1930 = ~n_1751 & n_1870;
assign n_1931 = ~n_1871 ^ n_187;
assign n_1932 = ~n_1872 ^ n_1004;
assign n_1933 = ~n_1873 ^ ~n_1271;
assign n_1934 = n_1871 & ~n_1874;
assign n_1935 = ~n_1871 ^ n_1874;
assign n_1936 = n_145 ^ n_1874;
assign n_1937 = n_165 ^ n_1874;
assign n_1938 = n_134 ^ n_1874;
assign n_1939 = n_121 ^ n_1874;
assign n_1940 = n_103 ^ n_1874;
assign n_1941 = n_111 ^ n_1874;
assign n_1942 = n_100 ^ n_1874;
assign n_1943 = n_87 ^ n_1874;
assign n_1944 = n_90 ^ n_1874;
assign n_1945 = n_74 ^ n_1874;
assign n_1946 = ~n_1872 & ~n_1875;
assign n_1947 = ~n_1876 ^ ~n_1690;
assign n_1948 = ~n_1815 & ~n_1877;
assign n_1949 = ~n_1721 ^ ~n_1880;
assign n_1950 = ~n_1682 ^ ~n_1881;
assign n_1951 = ~n_1623 & ~n_1882;
assign n_1952 = n_1874 & n_1888;
assign n_1953 = n_1874 ^ n_1888;
assign n_1954 = n_1869 ^ n_1888;
assign n_1955 = n_165 & ~n_1888;
assign n_1956 = n_187 ^ n_1888;
assign n_1957 = ~n_134 & ~n_1888;
assign n_1958 = n_145 ^ n_1888;
assign n_1959 = ~n_145 & ~n_1888;
assign n_1960 = n_165 ^ n_1888;
assign n_1961 = ~n_121 & ~n_1888;
assign n_1962 = n_134 ^ n_1888;
assign n_1963 = ~n_111 & ~n_1888;
assign n_1964 = n_121 ^ n_1888;
assign n_1965 = n_100 & ~n_1888;
assign n_1966 = n_103 ^ n_1888;
assign n_1967 = ~n_103 & ~n_1888;
assign n_1968 = n_111 ^ n_1888;
assign n_1969 = ~n_90 & ~n_1888;
assign n_1970 = n_100 ^ n_1888;
assign n_1971 = n_87 & ~n_1888;
assign n_1972 = n_90 ^ n_1888;
assign n_1973 = ~n_1848 & ~n_1889;
assign n_1974 = ~n_1890 ^ n_1888;
assign n_1975 = n_1890 & ~n_1888;
assign n_1976 = ~n_1890 & ~n_1874;
assign n_1977 = n_88 ^ ~n_1890;
assign n_1978 = n_1890 & ~n_88;
assign n_1979 = ~n_1891 & ~n_1719;
assign n_1980 = ~n_1891 & n_1696;
assign n_1981 = ~n_1892 ^ ~n_1799;
assign n_1982 = ~n_1892 & ~n_1846;
assign n_1983 = ~n_1894 ^ ~n_1467;
assign n_1984 = ~n_1844 ^ ~n_1895;
assign n_1985 = n_14 ^ n_1896;
assign n_1986 = n_1 & ~n_1896;
assign n_1987 = ~n_157 & n_1896;
assign n_1988 = n_260 & ~n_1896;
assign n_1989 = ~n_74 & ~n_1896;
assign n_1990 = n_98 & ~n_1896;
assign n_1991 = ~n_130 & ~n_1896;
assign n_1992 = n_100 & ~n_1896;
assign n_1993 = n_139 & ~n_1896;
assign n_1994 = n_121 ^ n_1896;
assign n_1995 = n_197 & ~n_1896;
assign n_1996 = ~n_121 & ~n_1896;
assign n_1997 = n_175 & ~n_1896;
assign n_1998 = n_165 ^ n_1896;
assign n_1999 = n_165 & ~n_1896;
assign n_2000 = ~n_432 & ~n_1896;
assign n_2001 = n_230 & ~n_1896;
assign n_2002 = n_1902 ^ n_1896;
assign n_2003 = ~n_187 & ~n_1905;
assign n_2004 = n_87 & n_1905;
assign n_2005 = ~n_1905 ^ n_88;
assign n_2006 = ~n_1905 ^ n_1888;
assign n_2007 = n_165 ^ n_1906;
assign n_2008 = n_187 ^ n_1906;
assign n_2009 = n_145 ^ n_1906;
assign n_2010 = n_134 ^ n_1906;
assign n_2011 = n_121 ^ n_1906;
assign n_2012 = n_111 ^ n_1906;
assign n_2013 = n_103 ^ n_1906;
assign n_2014 = n_100 ^ n_1906;
assign n_2015 = n_90 ^ n_1906;
assign n_2016 = n_74 ^ n_1906;
assign n_2017 = n_87 ^ n_1906;
assign n_2018 = n_314 & ~n_1906;
assign n_2019 = ~n_1908 ^ ~n_1768;
assign n_2020 = ~n_1908 & ~n_1800;
assign n_2021 = ~n_1871 ^ n_1913;
assign n_2022 = n_187 ^ n_1913;
assign n_2023 = n_165 ^ n_1913;
assign n_2024 = n_1913 ^ n_1874;
assign n_2025 = n_145 ^ n_1913;
assign n_2026 = n_134 ^ n_1913;
assign n_2027 = n_121 ^ n_1913;
assign n_2028 = n_111 ^ n_1913;
assign n_2029 = n_103 ^ n_1913;
assign n_2030 = n_90 ^ n_1913;
assign n_2031 = n_100 ^ n_1913;
assign n_2032 = n_87 ^ n_1913;
assign n_2033 = n_74 ^ n_1913;
assign n_2034 = ~n_1893 & ~n_1918;
assign n_2035 = ~n_1919 & n_1864;
assign n_2036 = n_1920 ^ n_165;
assign n_2037 = n_134 & n_1921;
assign n_2038 = n_1921 & n_90;
assign n_2039 = n_1921 & n_87;
assign n_2040 = ~n_134 & ~n_1922;
assign n_2041 = ~n_1922 & ~n_610;
assign n_2042 = ~n_1922 & n_17;
assign n_2043 = n_1923 ^ n_111;
assign n_2044 = ~n_1924 ^ n_100;
assign n_2045 = ~n_1925 ^ n_1787;
assign n_2046 = n_1926 ^ n_187;
assign n_2047 = n_1926 & n_1791;
assign n_2048 = ~n_307 & n_1927;
assign n_2049 = n_165 ^ n_1927;
assign n_2050 = n_1927 ^ n_1906;
assign n_2051 = n_187 ^ n_1927;
assign n_2052 = n_145 ^ n_1927;
assign n_2053 = n_134 ^ n_1927;
assign n_2054 = n_121 ^ n_1927;
assign n_2055 = n_111 ^ n_1927;
assign n_2056 = n_103 ^ n_1927;
assign n_2057 = n_100 ^ n_1927;
assign n_2058 = n_90 ^ n_1927;
assign n_2059 = n_87 ^ n_1927;
assign n_2060 = n_74 ^ n_1927;
assign n_2061 = n_88 ^ n_1927;
assign n_2062 = n_1928 & n_1864;
assign n_2063 = n_1929 ^ n_74;
assign n_2064 = n_1912 ^ n_1930;
assign n_2065 = ~n_1932 & ~n_1718;
assign n_2066 = ~n_1932 & ~n_1883;
assign n_2067 = ~n_1933 & n_1854;
assign n_2068 = ~n_1934 & ~n_1913;
assign n_2069 = n_88 ^ n_1934;
assign n_2070 = n_1935 & ~n_88;
assign n_2071 = ~n_1947 & ~n_1756;
assign n_2072 = ~n_1947 & ~n_1950;
assign n_2073 = ~n_1952 & ~n_1780;
assign n_2074 = n_1953 ^ n_187;
assign n_2075 = n_1890 & n_1954;
assign n_2076 = n_1955 ^ n_1956;
assign n_2077 = n_1957 ^ n_1958;
assign n_2078 = n_1959 ^ n_1960;
assign n_2079 = n_1961 ^ n_1962;
assign n_2080 = n_1963 ^ n_1964;
assign n_2081 = n_1965 ^ n_1966;
assign n_2082 = n_1967 ^ n_1968;
assign n_2083 = n_1969 ^ n_1970;
assign n_2084 = n_1971 ^ n_90;
assign n_2085 = n_1974 & n_1937;
assign n_2086 = n_1974 & ~n_1936;
assign n_2087 = n_1974 & ~n_1938;
assign n_2088 = n_1974 & ~n_1941;
assign n_2089 = n_1974 & ~n_1940;
assign n_2090 = n_1974 & ~n_1944;
assign n_2091 = n_1974 & n_1942;
assign n_2092 = n_1974 & ~n_1943;
assign n_2093 = n_1974 & ~n_1945;
assign n_2094 = n_1974 & ~n_1939;
assign n_2095 = n_1974 ^ n_1975;
assign n_2096 = n_1953 ^ n_1975;
assign n_2097 = n_1976 ^ n_1874;
assign n_2098 = n_165 & n_1976;
assign n_2099 = n_1974 & n_1977;
assign n_2100 = ~n_1933 & n_1979;
assign n_2101 = n_1980 & n_1885;
assign n_2102 = n_1980 ^ n_1885;
assign n_2103 = ~n_1604 ^ ~n_1983;
assign n_2104 = x1 & n_1985;
assign n_2105 = n_1988 ^ n_1827;
assign n_2106 = n_87 ^ ~n_1988;
assign n_2107 = n_1989 ^ n_87;
assign n_2108 = n_1991 ^ n_1831;
assign n_2109 = n_1992 ^ n_103;
assign n_2110 = n_1993 ^ n_103;
assign n_2111 = n_122 & n_1994;
assign n_2112 = n_1995 ^ n_1834;
assign n_2113 = n_1996 ^ n_134;
assign n_2114 = n_1997 ^ n_134;
assign n_2115 = ~n_1999 & n_1901;
assign n_2116 = n_87 ^ n_2001;
assign n_2117 = n_165 & n_2002;
assign n_2118 = ~n_2003 & ~n_1888;
assign n_2119 = n_1978 ^ n_2004;
assign n_2120 = n_1905 & n_2006;
assign n_2121 = ~n_2018 & ~n_1917;
assign n_2122 = n_2021 & n_1931;
assign n_2123 = n_1935 & n_2023;
assign n_2124 = n_2023 & n_2024;
assign n_2125 = ~n_1935 & n_2024;
assign n_2126 = n_1935 & ~n_2025;
assign n_2127 = n_1935 & ~n_2026;
assign n_2128 = n_1935 & ~n_2027;
assign n_2129 = n_1935 & ~n_2028;
assign n_2130 = n_1935 & ~n_2029;
assign n_2131 = n_1935 & ~n_2030;
assign n_2132 = n_1935 & n_2031;
assign n_2133 = n_1935 & ~n_2032;
assign n_2134 = n_1935 & ~n_2033;
assign n_2135 = n_2035 ^ n_145;
assign n_2136 = n_2037 ^ n_1712;
assign n_2137 = n_2038 ^ n_1712;
assign n_2138 = n_2039 ^ n_1712;
assign n_2139 = ~n_1921 & n_2044;
assign n_2140 = ~n_1921 & n_2045;
assign n_2141 = ~n_1789 ^ n_2046;
assign n_2142 = n_2046 ^ ~n_1790;
assign n_2143 = n_2048 ^ ~n_1776;
assign n_2144 = n_2048 ^ n_1864;
assign n_2145 = n_2048 ^ n_1712;
assign n_2146 = n_2048 ^ ~n_1781;
assign n_2147 = n_2048 ^ ~n_1785;
assign n_2148 = ~n_2048 & ~n_2036;
assign n_2149 = ~n_2048 & n_2043;
assign n_2150 = n_2062 ^ n_103;
assign n_2151 = n_2065 & ~n_1744;
assign n_2152 = n_2065 & n_1884;
assign n_2153 = n_2066 & n_1913;
assign n_2154 = n_2066 ^ n_1913;
assign n_2155 = n_2066 ^ n_1906;
assign n_2156 = n_2066 ^ n_187;
assign n_2157 = n_2068 ^ n_100;
assign n_2158 = n_2068 ^ n_1778;
assign n_2159 = n_2068 & ~n_2070;
assign n_2160 = n_2075 ^ n_1888;
assign n_2161 = ~n_1905 & n_2076;
assign n_2162 = ~n_1905 & ~n_2077;
assign n_2163 = ~n_1905 & n_2078;
assign n_2164 = ~n_1905 & ~n_2079;
assign n_2165 = ~n_1905 & ~n_2080;
assign n_2166 = ~n_1905 & ~n_2081;
assign n_2167 = ~n_1905 & ~n_2082;
assign n_2168 = ~n_1905 & n_2083;
assign n_2169 = ~n_1905 & n_2084;
assign n_2170 = ~n_2095 & ~n_1874;
assign n_2171 = n_2097 ^ n_187;
assign n_2172 = ~n_2098 & n_1888;
assign n_2173 = n_2099 ^ ~n_1890;
assign n_2174 = n_2101 ^ n_2102;
assign n_2175 = ~n_2103 ^ ~n_1677;
assign n_2176 = ~n_87 & n_2105;
assign n_2177 = ~n_2106 ^ n_176;
assign n_2178 = ~n_2106 & ~n_1828;
assign n_2179 = n_2108 ^ n_103;
assign n_2180 = n_2110 & ~n_125;
assign n_2181 = n_2117 ^ n_1896;
assign n_2182 = n_1786 ^ n_2118;
assign n_2183 = n_2120 ^ ~n_1905;
assign n_2184 = n_2101 & n_2121;
assign n_2185 = n_2122 ^ ~n_1871;
assign n_2186 = n_2022 ^ n_2124;
assign n_2187 = n_2125 & ~n_2025;
assign n_2188 = n_2125 & ~n_2026;
assign n_2189 = n_2125 & ~n_2027;
assign n_2190 = n_2125 & ~n_2028;
assign n_2191 = n_2125 & ~n_2029;
assign n_2192 = n_2125 & ~n_2030;
assign n_2193 = n_2125 & ~n_2032;
assign n_2194 = n_2125 & n_2069;
assign n_2195 = n_2125 & ~n_2033;
assign n_2196 = n_2125 & n_2031;
assign n_2197 = n_2139 ^ n_1782;
assign n_2198 = n_2140 ^ n_1787;
assign n_2199 = ~n_2142 & ~n_1791;
assign n_2200 = n_2143 & n_2135;
assign n_2201 = n_145 & n_2144;
assign n_2202 = n_121 & ~n_2144;
assign n_2203 = n_2144 & ~n_100;
assign n_2204 = n_2144 & n_90;
assign n_2205 = n_2144 & ~n_88;
assign n_2206 = n_2145 & ~n_2040;
assign n_2207 = n_2147 & n_2063;
assign n_2208 = ~n_1773 ^ ~n_2148;
assign n_2209 = ~n_1777 ^ ~n_2149;
assign n_2210 = n_2146 & n_2150;
assign n_2211 = ~n_1906 & ~n_2152;
assign n_2212 = n_1906 ^ n_2152;
assign n_2213 = n_1927 ^ n_2152;
assign n_2214 = n_187 ^ n_2152;
assign n_2215 = n_2153 & ~n_1906;
assign n_2216 = n_2153 ^ n_2154;
assign n_2217 = n_2154 & n_2008;
assign n_2218 = n_2154 & n_2007;
assign n_2219 = n_2154 & ~n_2009;
assign n_2220 = n_2154 & ~n_2010;
assign n_2221 = n_2154 & ~n_2011;
assign n_2222 = n_2154 & ~n_2012;
assign n_2223 = n_2154 & ~n_2013;
assign n_2224 = n_2154 & n_2014;
assign n_2225 = n_2154 & ~n_2017;
assign n_2226 = n_2154 & ~n_2016;
assign n_2227 = n_2154 & ~n_88;
assign n_2228 = n_2154 & ~n_2015;
assign n_2229 = n_2155 & n_2156;
assign n_2230 = ~n_112 & n_2157;
assign n_2231 = n_1956 ^ n_2161;
assign n_2232 = n_1958 ^ n_2162;
assign n_2233 = n_1960 ^ n_2163;
assign n_2234 = n_1962 ^ n_2164;
assign n_2235 = n_1964 ^ n_2165;
assign n_2236 = n_1966 ^ n_2166;
assign n_2237 = n_1968 ^ n_2167;
assign n_2238 = n_1970 ^ n_2168;
assign n_2239 = n_1972 ^ n_2169;
assign n_2240 = n_2170 ^ n_1976;
assign n_2241 = ~n_1974 & n_2171;
assign n_2242 = n_2173 & ~n_1874;
assign n_2243 = ~n_2174 & ~n_2121;
assign n_2244 = n_157 & ~n_2178;
assign n_2245 = n_2179 ^ n_100;
assign n_2246 = n_125 ^ n_2180;
assign n_2247 = ~n_184 & n_2181;
assign n_2248 = n_2005 & ~n_2183;
assign n_2249 = ~n_1935 & ~n_2185;
assign n_2250 = ~n_1935 & n_2186;
assign n_2251 = n_2187 ^ n_2123;
assign n_2252 = n_2188 ^ n_2126;
assign n_2253 = n_2189 ^ n_2127;
assign n_2254 = n_2190 ^ n_2128;
assign n_2255 = n_2191 ^ n_2129;
assign n_2256 = n_2192 ^ n_2132;
assign n_2257 = n_2193 ^ n_2131;
assign n_2258 = n_2134 ^ n_2194;
assign n_2259 = n_2195 ^ n_2133;
assign n_2260 = n_2196 ^ n_2130;
assign n_2261 = n_2145 & n_2197;
assign n_2262 = n_2145 & n_2198;
assign n_2263 = ~n_2201 ^ n_2136;
assign n_2264 = n_2202 ^ n_1864;
assign n_2265 = ~n_2203 ^ n_2137;
assign n_2266 = ~n_2204 ^ n_2138;
assign n_2267 = ~n_2208 & ~n_2200;
assign n_2268 = ~n_2211 & ~n_1927;
assign n_2269 = n_2212 & n_2051;
assign n_2270 = n_2212 & n_2049;
assign n_2271 = n_2212 & ~n_2052;
assign n_2272 = n_2212 & ~n_2053;
assign n_2273 = n_2212 & ~n_2054;
assign n_2274 = n_2212 & ~n_2055;
assign n_2275 = n_2212 & ~n_2056;
assign n_2276 = n_2212 & n_2057;
assign n_2277 = n_2212 & ~n_2058;
assign n_2278 = n_2212 & ~n_88;
assign n_2279 = n_2212 & ~n_2059;
assign n_2280 = n_2212 & ~n_2060;
assign n_2281 = n_2213 & n_2050;
assign n_2282 = n_2213 & n_2214;
assign n_2283 = n_2216 ^ n_1906;
assign n_2284 = ~n_2216 & n_1906;
assign n_2285 = n_2229 ^ n_2066;
assign n_2286 = n_2230 ^ n_100;
assign n_2287 = n_2231 & ~n_1712;
assign n_2288 = n_2231 ^ n_1712;
assign n_2289 = ~n_2073 & ~n_2240;
assign n_2290 = n_2240 ^ n_1952;
assign n_2291 = n_2241 ^ n_2074;
assign n_2292 = ~n_2070 & ~n_2242;
assign n_2293 = ~n_2239 & n_2242;
assign n_2294 = n_2243 ^ n_2184;
assign n_2295 = ~n_2115 ^ ~n_2247;
assign n_2296 = n_2248 ^ n_2120;
assign n_2297 = n_1913 ^ n_2249;
assign n_2298 = n_2022 ^ n_2250;
assign n_2299 = n_2234 ^ n_2256;
assign n_2300 = ~n_2258 & ~n_2159;
assign n_2301 = n_2159 ^ n_2258;
assign n_2302 = n_2237 ^ n_2259;
assign n_2303 = n_2264 & n_2206;
assign n_2304 = ~n_1775 & ~n_2268;
assign n_2305 = ~n_2278 & n_2268;
assign n_2306 = n_2049 & n_2281;
assign n_2307 = n_2281 & ~n_2052;
assign n_2308 = n_2281 & ~n_2053;
assign n_2309 = n_2281 & ~n_2054;
assign n_2310 = n_2281 & ~n_2055;
assign n_2311 = n_2281 & ~n_2056;
assign n_2312 = n_2281 & n_2057;
assign n_2313 = n_2281 & ~n_2058;
assign n_2314 = n_2281 & ~n_2059;
assign n_2315 = n_2281 & ~n_2060;
assign n_2316 = n_2281 & n_2061;
assign n_2317 = n_2282 ^ n_2152;
assign n_2318 = n_2283 ^ n_2284;
assign n_2319 = n_2215 ^ n_2284;
assign n_2320 = ~n_2154 & ~n_2285;
assign n_2321 = ~n_2286 & ~n_1712;
assign n_2322 = n_2287 ^ n_2207;
assign n_2323 = n_2288 ^ n_2262;
assign n_2324 = n_2289 ^ n_2210;
assign n_2325 = n_2289 ^ n_2073;
assign n_2326 = n_2096 ^ n_2290;
assign n_2327 = n_2293 ^ n_2238;
assign n_2328 = n_2296 ^ ~n_1905;
assign n_2329 = n_2297 ^ n_1779;
assign n_2330 = n_2298 ^ n_2261;
assign n_2331 = n_2300 ^ n_2236;
assign n_2332 = n_2301 ^ n_2300;
assign n_2333 = ~n_2208 ^ n_2304;
assign n_2334 = ~n_2208 & ~n_2304;
assign n_2335 = n_165 & ~n_2304;
assign n_2336 = n_2305 & ~n_2232;
assign n_2337 = n_2232 ^ n_2305;
assign n_2338 = ~n_2306 ^ ~n_2269;
assign n_2339 = n_2307 ^ n_2270;
assign n_2340 = n_2308 ^ n_2271;
assign n_2341 = n_2309 ^ n_2272;
assign n_2342 = n_2310 ^ n_2273;
assign n_2343 = n_2311 ^ n_2274;
assign n_2344 = n_2312 ^ n_2275;
assign n_2345 = n_2313 ^ n_2276;
assign n_2346 = n_2314 ^ n_2277;
assign n_2347 = n_2315 ^ n_2279;
assign n_2348 = n_2280 ^ n_2316;
assign n_2349 = ~n_2212 & ~n_2317;
assign n_2350 = n_2318 ^ n_121;
assign n_2351 = n_2318 & n_88;
assign n_2352 = n_1788 ^ n_2318;
assign n_2353 = n_2007 & n_2319;
assign n_2354 = n_2319 & ~n_2009;
assign n_2355 = n_2319 & ~n_2010;
assign n_2356 = n_2319 & ~n_2011;
assign n_2357 = n_2319 & ~n_2012;
assign n_2358 = n_2319 & ~n_2013;
assign n_2359 = n_2319 & n_2014;
assign n_2360 = n_2319 & ~n_2015;
assign n_2361 = n_2319 & ~n_2016;
assign n_2362 = n_2319 & ~n_88;
assign n_2363 = n_2319 & ~n_2017;
assign n_2364 = n_1906 ^ n_2320;
assign n_2365 = n_2303 ^ n_2321;
assign n_2366 = n_2326 ^ n_2095;
assign n_2367 = ~n_165 & ~n_2326;
assign n_2368 = n_2326 ^ n_2170;
assign n_2369 = n_2328 ^ n_1888;
assign n_2370 = n_2333 & n_1712;
assign n_2371 = n_2333 ^ n_2334;
assign n_2372 = n_2267 ^ n_2335;
assign n_2373 = n_2336 ^ n_2255;
assign n_2374 = ~n_2338 ^ ~n_2263;
assign n_2375 = n_1865 ^ n_2339;
assign n_2376 = n_2341 ^ n_2289;
assign n_2377 = n_2341 ^ n_2324;
assign n_2378 = n_2342 ^ n_2298;
assign n_2379 = n_2342 ^ n_2330;
assign n_2380 = n_2337 ^ n_2348;
assign n_2381 = n_1927 ^ n_2349;
assign n_2382 = n_135 & n_2350;
assign n_2383 = ~n_2215 & ~n_2351;
assign n_2384 = ~n_2353 ^ ~n_2217;
assign n_2385 = n_2354 ^ n_2218;
assign n_2386 = n_2355 ^ n_2219;
assign n_2387 = n_2356 ^ n_2220;
assign n_2388 = n_2357 ^ n_2221;
assign n_2389 = n_2358 ^ n_2222;
assign n_2390 = n_2359 ^ n_2223;
assign n_2391 = n_2360 ^ n_2224;
assign n_2392 = n_2361 ^ n_2225;
assign n_2393 = n_2226 ^ n_2362;
assign n_2394 = n_2363 ^ n_2228;
assign n_2395 = n_2364 ^ n_1865;
assign n_2396 = ~n_187 & n_2366;
assign n_2397 = ~n_165 & n_2366;
assign n_2398 = n_1869 & ~n_2367;
assign n_2399 = ~n_2368 & ~n_1936;
assign n_2400 = ~n_2368 & ~n_1938;
assign n_2401 = ~n_2368 & ~n_1939;
assign n_2402 = ~n_2368 & ~n_1940;
assign n_2403 = ~n_2368 & n_1942;
assign n_2404 = ~n_2368 & ~n_1943;
assign n_2405 = ~n_2368 & ~n_1944;
assign n_2406 = ~n_2368 & ~n_1945;
assign n_2407 = ~n_88 & ~n_2368;
assign n_2408 = ~n_2368 & ~n_1941;
assign n_2409 = n_74 & n_2369;
assign n_2410 = ~n_2334 & ~n_2370;
assign n_2411 = ~n_134 & n_2371;
assign n_2412 = n_2364 ^ n_2375;
assign n_2413 = ~n_2324 & n_2376;
assign n_2414 = ~n_2330 & n_2378;
assign n_2415 = n_2381 & ~n_2200;
assign n_2416 = n_2381 ^ n_2200;
assign n_2417 = n_2381 & n_2372;
assign n_2418 = n_2382 ^ n_111;
assign n_2419 = ~n_2235 & ~n_2383;
assign n_2420 = n_2235 ^ n_2383;
assign n_2421 = ~n_2384 ^ ~n_2209;
assign n_2422 = n_2340 ^ ~n_2384;
assign n_2423 = n_1779 ^ n_2385;
assign n_2424 = n_2297 ^ n_2385;
assign n_2425 = n_2329 ^ n_2385;
assign n_2426 = ~n_1952 & n_2386;
assign n_2427 = n_2386 ^ n_1780;
assign n_2428 = n_2387 ^ n_2251;
assign n_2429 = n_2343 ^ n_2387;
assign n_2430 = n_2388 ^ n_2252;
assign n_2431 = n_2344 ^ n_2388;
assign n_2432 = n_2389 ^ n_2253;
assign n_2433 = n_2345 ^ n_2389;
assign n_2434 = n_2390 ^ n_2254;
assign n_2435 = n_2346 ^ n_2390;
assign n_2436 = n_2391 ^ n_2255;
assign n_2437 = n_2392 ^ n_2278;
assign n_2438 = n_2278 & n_2392;
assign n_2439 = n_2393 ^ n_2215;
assign n_2440 = n_2260 ^ n_2394;
assign n_2441 = n_2375 & n_2395;
assign n_2442 = n_2396 & ~n_1888;
assign n_2443 = ~n_2290 & ~n_2396;
assign n_2444 = ~n_2397 & ~n_2291;
assign n_2445 = ~n_2398 & ~n_2172;
assign n_2446 = ~n_2399 ^ ~n_2085;
assign n_2447 = n_2400 ^ n_2086;
assign n_2448 = n_2401 ^ n_2087;
assign n_2449 = n_2402 ^ n_2088;
assign n_2450 = n_2403 ^ n_2089;
assign n_2451 = n_2404 ^ n_2090;
assign n_2452 = n_2405 ^ n_2091;
assign n_2453 = n_2406 ^ n_2092;
assign n_2454 = n_2407 ^ n_2170;
assign n_2455 = n_2408 ^ n_2094;
assign n_2456 = n_2004 & ~n_2409;
assign n_2457 = n_1888 ^ n_2409;
assign n_2458 = ~n_2381 & ~n_2410;
assign n_2459 = ~n_2370 & ~n_2411;
assign n_2460 = n_2413 ^ n_2341;
assign n_2461 = n_2414 ^ n_2342;
assign n_2462 = ~n_2333 & n_2415;
assign n_2463 = n_2267 ^ n_2417;
assign n_2464 = n_2418 & ~n_2416;
assign n_2465 = n_2418 ^ n_134;
assign n_2466 = n_2340 ^ n_2421;
assign n_2467 = ~n_2421 & ~n_2422;
assign n_2468 = ~n_2423 & n_2424;
assign n_2469 = n_2377 ^ n_2425;
assign n_2470 = n_2343 ^ n_2428;
assign n_2471 = ~n_2428 & n_2429;
assign n_2472 = n_2344 ^ n_2430;
assign n_2473 = ~n_2430 & n_2431;
assign n_2474 = n_2345 ^ n_2432;
assign n_2475 = ~n_2432 & n_2433;
assign n_2476 = n_2346 ^ n_2434;
assign n_2477 = ~n_2434 & n_2435;
assign n_2478 = n_2436 & ~n_2373;
assign n_2479 = n_2336 ^ n_2436;
assign n_2480 = n_2419 & n_2438;
assign n_2481 = n_2438 ^ n_2437;
assign n_2482 = n_2441 ^ n_2339;
assign n_2483 = n_2442 ^ n_2240;
assign n_2484 = n_1867 & n_2443;
assign n_2485 = n_2443 ^ n_1867;
assign n_2486 = n_1869 ^ n_2444;
assign n_2487 = ~n_2446 ^ n_1786;
assign n_2488 = ~n_2446 ^ n_2118;
assign n_2489 = n_2182 ^ ~n_2446;
assign n_2490 = n_2447 ^ n_2288;
assign n_2491 = n_2447 ^ n_2323;
assign n_2492 = n_2233 ^ n_2448;
assign n_2493 = n_2347 ^ n_2448;
assign n_2494 = n_2234 ^ n_2449;
assign n_2495 = n_2450 ^ n_2257;
assign n_2496 = n_2439 ^ n_2450;
assign n_2497 = n_2236 ^ n_2451;
assign n_2498 = n_2451 & ~n_2236;
assign n_2499 = n_2259 ^ n_2452;
assign n_2500 = n_2238 ^ n_2453;
assign n_2501 = n_2093 ^ n_2454;
assign n_2502 = n_2260 ^ n_2455;
assign n_2503 = n_2456 ^ n_2457;
assign n_2504 = n_2200 & ~n_2459;
assign n_2505 = n_2425 ^ n_2461;
assign n_2506 = n_2334 ^ n_2462;
assign n_2507 = n_2463 & ~n_1712;
assign n_2508 = n_2464 & n_1712;
assign n_2509 = n_2465 & ~n_1712;
assign n_2510 = n_2467 ^ n_2340;
assign n_2511 = n_2468 ^ n_1779;
assign n_2512 = n_2469 ^ n_2461;
assign n_2513 = n_2471 ^ n_2343;
assign n_2514 = n_2473 ^ n_2344;
assign n_2515 = n_2475 ^ n_2345;
assign n_2516 = n_2477 ^ n_2346;
assign n_2517 = n_2478 ^ n_2391;
assign n_2518 = n_2479 ^ n_2205;
assign n_2519 = n_2480 ^ n_2437;
assign n_2520 = ~n_2419 & ~n_2481;
assign n_2521 = n_2482 ^ ~n_2338;
assign n_2522 = n_2482 ^ n_2374;
assign n_2523 = n_2483 ^ n_2484;
assign n_2524 = n_2470 ^ n_2485;
assign n_2525 = n_2472 ^ n_2486;
assign n_2526 = n_2486 & ~n_2160;
assign n_2527 = ~n_2487 & n_2488;
assign n_2528 = n_2489 ^ n_2474;
assign n_2529 = n_2323 & ~n_2490;
assign n_2530 = n_2347 ^ n_2492;
assign n_2531 = ~n_2492 & n_2493;
assign n_2532 = n_2494 ^ n_2256;
assign n_2533 = ~n_2494 & n_2299;
assign n_2534 = n_2439 ^ n_2495;
assign n_2535 = n_2495 & ~n_2496;
assign n_2536 = ~n_2497 & ~n_2331;
assign n_2537 = n_2301 ^ n_2497;
assign n_2538 = n_2499 & n_2302;
assign n_2539 = n_2237 ^ n_2499;
assign n_2540 = n_2500 ^ ~n_2292;
assign n_2541 = n_2500 & ~n_2327;
assign n_2542 = n_2501 ^ n_2500;
assign n_2543 = n_2500 & n_2501;
assign n_2544 = n_2502 ^ n_2394;
assign n_2545 = ~n_2502 & n_2440;
assign n_2546 = ~n_2119 & ~n_2503;
assign n_2547 = ~n_2462 ^ ~n_2504;
assign n_2548 = n_2469 & ~n_2505;
assign n_2549 = ~n_2506 & ~n_2507;
assign n_2550 = ~n_2507 & ~n_2458;
assign n_2551 = n_2418 ^ n_2508;
assign n_2552 = n_2416 ^ n_2509;
assign n_2553 = n_2365 ^ n_2510;
assign n_2554 = n_2510 ^ n_2321;
assign n_2555 = n_2158 ^ n_2511;
assign n_2556 = n_2460 ^ n_2511;
assign n_2557 = n_2379 ^ n_2513;
assign n_2558 = ~n_2265 ^ n_2514;
assign n_2559 = n_2515 ^ ~n_2266;
assign n_2560 = n_2516 ^ n_2287;
assign n_2561 = n_2516 ^ n_2322;
assign n_2562 = n_2476 ^ n_2517;
assign n_2563 = n_2519 ^ n_2520;
assign n_2564 = ~n_2374 & ~n_2521;
assign n_2565 = n_2523 ^ n_2240;
assign n_2566 = ~n_2526 & ~n_2445;
assign n_2567 = n_2527 ^ n_1786;
assign n_2568 = n_2529 ^ n_2447;
assign n_2569 = n_2531 ^ n_2347;
assign n_2570 = n_2532 ^ n_2419;
assign n_2571 = n_2533 ^ n_2449;
assign n_2572 = n_2534 ^ n_2420;
assign n_2573 = n_2420 & n_2534;
assign n_2574 = n_2535 ^ n_2257;
assign n_2575 = n_2536 ^ n_2451;
assign n_2576 = n_2537 ^ n_2292;
assign n_2577 = n_2537 ^ n_2238;
assign n_2578 = n_2537 ^ n_2500;
assign n_2579 = n_2538 ^ n_2452;
assign n_2580 = n_2540 & n_2239;
assign n_2581 = n_2453 ^ n_2541;
assign n_2582 = n_2542 ^ n_2543;
assign n_2583 = ~n_2070 & ~n_2543;
assign n_2584 = n_2545 ^ n_2394;
assign n_2585 = n_2548 ^ n_2377;
assign n_2586 = n_2549 ^ ~n_2141;
assign n_2587 = n_2549 & n_2142;
assign n_2588 = ~n_2547 & n_2550;
assign n_2589 = n_2553 ^ n_2412;
assign n_2590 = ~n_2365 & n_2554;
assign n_2591 = n_2460 ^ n_2555;
assign n_2592 = ~n_2555 & ~n_2556;
assign n_2593 = ~n_2322 & n_2560;
assign n_2594 = n_2563 ^ n_2419;
assign n_2595 = n_2564 ^ n_2482;
assign n_2596 = n_2565 ^ n_2386;
assign n_2597 = n_2565 ^ n_1952;
assign n_2598 = ~n_2265 ^ n_2566;
assign n_2599 = n_2558 ^ n_2566;
assign n_2600 = ~n_2266 ^ n_2567;
assign n_2601 = n_2489 ^ n_2568;
assign n_2602 = n_2569 ^ n_2476;
assign n_2603 = n_2569 ^ n_2562;
assign n_2604 = n_2570 ^ n_2437;
assign n_2605 = n_2571 ^ n_2380;
assign n_2606 = n_2571 ^ n_2348;
assign n_2607 = n_2572 ^ n_2573;
assign n_2608 = n_2574 & ~n_2532;
assign n_2609 = n_2532 ^ n_2574;
assign n_2610 = n_2227 ^ n_2575;
assign n_2611 = n_2537 & ~n_2578;
assign n_2612 = ~n_2537 & n_2581;
assign n_2613 = ~n_2582 & ~n_2242;
assign n_2614 = n_2582 & ~n_2583;
assign n_2615 = n_2518 ^ n_2584;
assign n_2616 = n_2205 ^ n_2584;
assign n_2617 = n_2585 ^ n_2466;
assign n_2618 = ~n_2466 & ~n_2585;
assign n_2619 = ~n_2587 & ~n_2047;
assign n_2620 = n_2590 ^ n_2510;
assign n_2621 = n_2592 ^ n_2460;
assign n_2622 = n_2593 ^ n_2516;
assign n_2623 = n_2595 ^ n_2552;
assign n_2624 = ~n_2427 & n_2596;
assign n_2625 = n_2597 ^ n_2427;
assign n_2626 = ~n_2558 & ~n_2598;
assign n_2627 = ~n_2600 & n_2559;
assign n_2628 = n_2515 ^ n_2600;
assign n_2629 = n_2601 ^ n_2474;
assign n_2630 = ~n_2601 & n_2528;
assign n_2631 = n_2562 & ~n_2602;
assign n_2632 = n_2604 ^ n_2574;
assign n_2633 = n_2380 & n_2606;
assign n_2634 = ~n_2594 & n_2608;
assign n_2635 = n_2520 & ~n_2608;
assign n_2636 = n_2608 ^ n_2609;
assign n_2637 = n_2498 ^ n_2610;
assign n_2638 = n_2611 ^ n_2537;
assign n_2639 = n_2539 ^ n_2612;
assign n_2640 = ~n_2580 ^ ~n_2613;
assign n_2641 = n_2239 & ~n_2614;
assign n_2642 = n_2530 ^ n_2615;
assign n_2643 = n_2518 & ~n_2616;
assign n_2644 = n_2617 ^ n_2618;
assign n_2645 = n_2620 ^ n_2522;
assign n_2646 = n_2352 ^ n_2620;
assign n_2647 = n_2589 ^ n_2621;
assign n_2648 = n_2553 ^ n_2621;
assign n_2649 = n_2622 ^ n_2472;
assign n_2650 = n_2622 ^ n_2525;
assign n_2651 = n_2623 ^ n_134;
assign n_2652 = n_2325 ^ n_2624;
assign n_2653 = n_2626 ^ n_2514;
assign n_2654 = n_2627 ^ n_2567;
assign n_2655 = n_2561 ^ n_2629;
assign n_2656 = n_2630 ^ n_2568;
assign n_2657 = n_2631 ^ n_2517;
assign n_2658 = n_2573 ^ n_2632;
assign n_2659 = n_2633 ^ n_2571;
assign n_2660 = n_2480 & ~n_2636;
assign n_2661 = n_2594 & n_2636;
assign n_2662 = n_2332 & ~n_2637;
assign n_2663 = ~n_2577 & n_2638;
assign n_2664 = n_2639 ^ n_2539;
assign n_2665 = ~n_2640 ^ ~n_2583;
assign n_2666 = n_2643 ^ n_2479;
assign n_2667 = n_2352 ^ n_2645;
assign n_2668 = n_2645 & n_2646;
assign n_2669 = n_2618 ^ n_2647;
assign n_2670 = n_2589 & n_2648;
assign n_2671 = n_2525 & n_2649;
assign n_2672 = n_2628 ^ n_2650;
assign n_2673 = n_2651 ^ n_2465;
assign n_2674 = n_2426 ^ n_2652;
assign n_2675 = n_2653 ^ n_2513;
assign n_2676 = n_2653 ^ n_2557;
assign n_2677 = n_2654 ^ n_2470;
assign n_2678 = n_2654 ^ n_2524;
assign n_2679 = n_2657 ^ n_2561;
assign n_2680 = n_2657 ^ n_2655;
assign n_2681 = n_2530 ^ n_2659;
assign n_2682 = ~n_2634 & ~n_2660;
assign n_2683 = ~n_2661 & ~n_2635;
assign n_2684 = n_2662 ^ n_2498;
assign n_2685 = n_2663 ^ n_2611;
assign n_2686 = n_2665 & ~n_2546;
assign n_2687 = n_2666 ^ n_2603;
assign n_2688 = n_2603 & n_2666;
assign n_2689 = n_2668 ^ n_2646;
assign n_2690 = n_2668 ^ n_2522;
assign n_2691 = n_2670 ^ n_2621;
assign n_2692 = n_2671 ^ n_2622;
assign n_2693 = n_2552 & ~n_2673;
assign n_2694 = n_2512 ^ n_2674;
assign n_2695 = ~n_2557 & n_2675;
assign n_2696 = ~n_2524 & n_2677;
assign n_2697 = n_2678 ^ n_2599;
assign n_2698 = n_2655 & n_2679;
assign n_2699 = n_2681 ^ n_2615;
assign n_2700 = n_2681 & ~n_2642;
assign n_2701 = n_2682 ^ n_2683;
assign n_2702 = ~n_2605 & n_2683;
assign n_2703 = ~n_2227 & ~n_2684;
assign n_2704 = n_2539 ^ n_2684;
assign n_2705 = n_2685 ^ n_2537;
assign n_2706 = n_2687 ^ n_2688;
assign n_2707 = n_2688 ^ n_2680;
assign n_2708 = n_2522 & n_2689;
assign n_2709 = n_2667 ^ n_2691;
assign n_2710 = n_2692 ^ n_2678;
assign n_2711 = n_2551 ^ n_2693;
assign n_2712 = n_2695 ^ n_2653;
assign n_2713 = n_2696 ^ n_2654;
assign n_2714 = n_2692 ^ n_2697;
assign n_2715 = n_2698 ^ n_2657;
assign n_2716 = n_2605 ^ n_2699;
assign n_2717 = n_2700 ^ n_2659;
assign n_2718 = ~n_2699 & n_2701;
assign n_2719 = ~n_2702 & n_2682;
assign n_2720 = n_2575 & ~n_2703;
assign n_2721 = n_2705 ^ n_2500;
assign n_2722 = n_2708 ^ n_2691;
assign n_2723 = ~n_2691 & ~n_2708;
assign n_2724 = n_2708 ^ n_2689;
assign n_2725 = ~n_2697 & n_2710;
assign n_2726 = n_2711 ^ n_2588;
assign n_2727 = n_2712 ^ n_2674;
assign n_2728 = n_2712 ^ n_2694;
assign n_2729 = n_2625 ^ n_2713;
assign n_2730 = n_2714 ^ n_2650;
assign n_2731 = n_2715 ^ n_2650;
assign n_2732 = n_2715 ^ n_2672;
assign n_2733 = n_2717 ^ n_2491;
assign n_2734 = ~n_2491 & n_2717;
assign n_2735 = n_2718 ^ n_2683;
assign n_2736 = n_2699 ^ n_2719;
assign n_2737 = n_2579 ^ n_2720;
assign n_2738 = n_2579 & n_2720;
assign n_2739 = n_2576 & ~n_2721;
assign n_2740 = n_2722 ^ n_2723;
assign n_2741 = ~n_2723 & n_2690;
assign n_2742 = ~n_2691 & n_2724;
assign n_2743 = n_2725 ^ n_2692;
assign n_2744 = n_2694 & ~n_2727;
assign n_2745 = n_2728 ^ n_2713;
assign n_2746 = ~n_2672 & n_2731;
assign n_2747 = n_2733 ^ n_2734;
assign n_2748 = n_2680 ^ ~n_2734;
assign n_2749 = ~n_2716 & n_2735;
assign n_2750 = n_2737 ^ n_2738;
assign n_2751 = n_2632 ^ ~n_2738;
assign n_2752 = n_2537 ^ n_2739;
assign n_2753 = ~n_2623 & n_2740;
assign n_2754 = n_2709 ^ n_2741;
assign n_2755 = n_2742 ^ n_2740;
assign n_2756 = n_2623 & ~n_2742;
assign n_2757 = n_2743 ^ n_2713;
assign n_2758 = n_2743 ^ n_2729;
assign n_2759 = n_2744 ^ n_2712;
assign n_2760 = ~n_2730 & n_2746;
assign n_2761 = n_2746 ^ n_2672;
assign n_2762 = ~n_2680 ^ ~n_2747;
assign n_2763 = n_2748 & n_2706;
assign n_2764 = n_2605 ^ n_2749;
assign n_2765 = ~n_2632 ^ n_2750;
assign n_2766 = n_2751 & n_2607;
assign n_2767 = ~n_2752 & ~n_2641;
assign n_2768 = n_2754 ^ n_2755;
assign n_2769 = ~n_2741 & ~n_2756;
assign n_2770 = n_2729 & n_2757;
assign n_2771 = n_2759 ^ n_2591;
assign n_2772 = n_2760 ^ n_2714;
assign n_2773 = n_2761 ^ n_2715;
assign n_2774 = ~n_2686 & n_2767;
assign n_2775 = ~n_2753 ^ ~n_2768;
assign n_2776 = n_2768 ^ n_2741;
assign n_2777 = n_2770 ^ n_2729;
assign n_2778 = n_2770 ^ n_2743;
assign n_2779 = ~n_2591 & ~n_2771;
assign n_2780 = n_2617 ^ n_2771;
assign n_2781 = n_2773 ^ n_2714;
assign n_2782 = n_2773 ^ n_2656;
assign n_2783 = n_2539 ^ n_2774;
assign n_2784 = ~n_2745 & n_2777;
assign n_2785 = n_2778 ^ n_2728;
assign n_2786 = n_2778 ^ n_2676;
assign n_2787 = n_2779 ^ n_2771;
assign n_2788 = ~n_2647 ^ ~n_2779;
assign n_2789 = n_2644 ^ n_2779;
assign n_2790 = n_2782 ^ n_2746;
assign n_2791 = n_2783 ^ n_2539;
assign n_2792 = n_2784 ^ n_2728;
assign n_2793 = n_2786 ^ n_2777;
assign n_2794 = n_2647 ^ n_2787;
assign n_2795 = n_2788 & n_2644;
assign n_2796 = ~n_2791 & ~n_2664;
assign n_2797 = n_2539 ^ n_2796;
assign n_2798 = n_2704 & ~n_2797;
assign n_2799 = n_2684 ^ n_2798;
assign n_2800 = n_2765 ^ n_2799;
assign n_2801 = n_2799 ^ n_2579;
assign n_2802 = n_2800 & n_2766;
assign n_2803 = n_2737 & n_2801;
assign n_2804 = n_2803 ^ n_2720;
assign n_2805 = n_2804 ^ n_2573;
assign n_2806 = ~n_2658 & ~n_2805;
assign n_2807 = n_2632 ^ n_2806;
assign n_2808 = n_2807 & ~n_2802;
assign n_2809 = ~n_2544 & n_2808;
assign n_2810 = n_2544 ^ n_2808;
assign n_2811 = ~n_2809 & ~n_2764;
assign n_2812 = n_2810 ^ n_2809;
assign n_2813 = n_2812 ^ n_2719;
assign n_2814 = ~n_2736 & n_2813;
assign n_2815 = n_2814 ^ n_2699;
assign n_2816 = ~n_2815 & ~n_2811;
assign n_2817 = n_2762 ^ n_2816;
assign n_2818 = n_2717 ^ n_2816;
assign n_2819 = n_2817 & n_2763;
assign n_2820 = n_2733 & n_2818;
assign n_2821 = n_2820 ^ n_2733;
assign n_2822 = n_2821 ^ n_2816;
assign n_2823 = n_2822 ^ n_2680;
assign n_2824 = n_2822 ^ n_2666;
assign n_2825 = ~n_2707 & n_2823;
assign n_2826 = n_2824 ^ n_2820;
assign n_2827 = n_2825 ^ n_2680;
assign n_2828 = ~n_2687 & n_2826;
assign n_2829 = n_2827 & ~n_2819;
assign n_2830 = n_2828 ^ n_2820;
assign n_2831 = n_2656 ^ n_2829;
assign n_2832 = ~n_2656 & n_2829;
assign n_2833 = n_2830 ^ n_2680;
assign n_2834 = n_2831 & n_2790;
assign n_2835 = n_2732 ^ n_2831;
assign n_2836 = n_2831 ^ n_2832;
assign n_2837 = n_2773 ^ n_2832;
assign n_2838 = n_2833 & n_1973;
assign n_2839 = n_2833 ^ n_1973;
assign n_2840 = n_2834 ^ n_2746;
assign n_2841 = n_2835 ^ ~n_1843;
assign n_2842 = ~n_2772 & ~n_2836;
assign n_2843 = n_2837 & ~n_2781;
assign n_2844 = n_2838 ^ ~n_1843;
assign n_2845 = ~n_165 & ~n_2839;
assign n_2846 = ~n_2839 & n_185;
assign n_2847 = ~n_2839 & n_301;
assign n_2848 = ~n_187 & ~n_2839;
assign n_2849 = n_145 & ~n_2839;
assign n_2850 = n_163 & ~n_2839;
assign n_2851 = n_121 & ~n_2839;
assign n_2852 = n_123 ^ n_2839;
assign n_2853 = ~n_2839 & n_198;
assign n_2854 = ~n_2839 & n_122;
assign n_2855 = ~n_2839 & ~n_231;
assign n_2856 = n_111 & ~n_2839;
assign n_2857 = ~n_2839 & ~n_108;
assign n_2858 = ~n_2839 & n_98;
assign n_2859 = ~n_2839 & n_140;
assign n_2860 = ~n_2839 & n_158;
assign n_2861 = ~n_2839 & ~n_262;
assign n_2862 = n_2840 ^ n_2714;
assign n_2863 = ~n_2841 & n_2839;
assign n_2864 = n_2838 ^ n_2841;
assign n_2865 = n_2841 ^ n_121;
assign n_2866 = n_2843 ^ n_2773;
assign n_2867 = ~n_2841 & ~n_2844;
assign n_2868 = ~n_2845 & ~n_237;
assign n_2869 = n_2846 ^ n_164;
assign n_2870 = ~n_137 & ~n_2851;
assign n_2871 = n_87 & n_2858;
assign n_2872 = n_1858 ^ n_2862;
assign n_2873 = n_2863 ^ n_2839;
assign n_2874 = ~n_2863 & ~n_300;
assign n_2875 = n_2864 & n_208;
assign n_2876 = n_2864 & n_236;
assign n_2877 = n_2864 & n_234;
assign n_2878 = n_2849 ^ n_2864;
assign n_2879 = n_2864 & n_197;
assign n_2880 = n_2864 & n_198;
assign n_2881 = n_2864 & ~n_130;
assign n_2882 = n_2864 & n_98;
assign n_2883 = n_2856 ^ n_2864;
assign n_2884 = n_2864 & n_431;
assign n_2885 = n_2864 & ~n_96;
assign n_2886 = n_2864 & ~n_157;
assign n_2887 = n_2864 & ~n_48;
assign n_2888 = n_123 & n_2865;
assign n_2889 = ~n_2866 & ~n_2842;
assign n_2890 = n_2867 ^ n_2835;
assign n_2891 = ~n_2863 & ~n_2868;
assign n_2892 = n_2873 ^ n_2864;
assign n_2893 = n_207 & n_2873;
assign n_2894 = n_2873 & n_150;
assign n_2895 = ~n_112 & n_2873;
assign n_2896 = n_2873 & n_115;
assign n_2897 = n_87 & ~n_2874;
assign n_2898 = ~n_184 & ~n_2875;
assign n_2899 = n_164 & ~n_2876;
assign n_2900 = ~n_2877 ^ ~n_2847;
assign n_2901 = ~n_163 & n_2878;
assign n_2902 = n_2879 ^ n_2853;
assign n_2903 = n_2881 ^ n_2855;
assign n_2904 = n_2839 & ~n_2882;
assign n_2905 = n_2857 ^ n_2882;
assign n_2906 = ~n_122 & n_2883;
assign n_2907 = n_2859 ^ n_2885;
assign n_2908 = n_2839 & ~n_2886;
assign n_2909 = n_2886 ^ n_2861;
assign n_2910 = n_2888 ^ n_2841;
assign n_2911 = n_2676 ^ n_2889;
assign n_2912 = ~n_2676 & ~n_2889;
assign n_2913 = n_2862 ^ n_2890;
assign n_2914 = n_1858 ^ n_2890;
assign n_2915 = n_2872 ^ n_2890;
assign n_2916 = ~n_2869 & n_2891;
assign n_2917 = n_2898 ^ n_2899;
assign n_2918 = n_165 ^ n_2899;
assign n_2919 = n_2864 ^ n_2901;
assign n_2920 = ~n_131 & ~n_2904;
assign n_2921 = n_2864 ^ n_2906;
assign n_2922 = n_372 & ~n_2908;
assign n_2923 = n_2852 & n_2910;
assign n_2924 = ~n_2911 & ~n_2793;
assign n_2925 = n_2758 ^ n_2911;
assign n_2926 = n_2911 ^ n_2912;
assign n_2927 = n_2778 ^ n_2912;
assign n_2928 = n_2913 & n_2914;
assign n_2929 = n_2915 & ~n_2892;
assign n_2930 = ~n_2915 & n_2864;
assign n_2931 = n_2893 ^ n_2915;
assign n_2932 = ~n_2915 & n_301;
assign n_2933 = ~n_2915 & n_198;
assign n_2934 = n_2894 ^ n_2915;
assign n_2935 = ~n_2915 & n_197;
assign n_2936 = ~n_2915 & ~n_130;
assign n_2937 = n_2895 ^ n_2915;
assign n_2938 = ~n_2915 & ~n_231;
assign n_2939 = ~n_2915 & n_260;
assign n_2940 = n_2896 ^ n_2915;
assign n_2941 = ~n_2915 & n_140;
assign n_2942 = n_0 & ~n_2915;
assign n_2943 = ~n_2841 & n_2915;
assign n_2944 = n_2915 & ~n_48;
assign n_2945 = ~n_187 & n_2916;
assign n_2946 = n_2915 & ~n_2918;
assign n_2947 = n_2845 ^ n_2919;
assign n_2948 = n_103 & n_2920;
assign n_2949 = n_2921 ^ n_2851;
assign n_2950 = n_2839 ^ n_2923;
assign n_2951 = n_2924 ^ n_2777;
assign n_2952 = n_2925 ^ n_1915;
assign n_2953 = n_2792 & n_2926;
assign n_2954 = ~n_2927 & ~n_2785;
assign n_2955 = n_2928 ^ n_2862;
assign n_2956 = n_2929 ^ n_2930;
assign n_2957 = n_163 & ~n_2931;
assign n_2958 = n_122 & ~n_2934;
assign n_2959 = ~n_2935 ^ ~n_2880;
assign n_2960 = n_98 & ~n_2937;
assign n_2961 = n_2939 ^ n_2884;
assign n_2962 = n_2940 ^ n_2907;
assign n_2963 = n_2942 ^ n_2887;
assign n_2964 = n_2943 ^ n_88;
assign n_2965 = n_2946 ^ n_165;
assign n_2966 = n_103 ^ n_2948;
assign n_2967 = ~n_2870 & ~n_2950;
assign n_2968 = n_2951 ^ n_2728;
assign n_2969 = n_2954 ^ n_2778;
assign n_2970 = n_2955 ^ n_2925;
assign n_2971 = n_2955 ^ n_2952;
assign n_2972 = n_207 & ~n_2956;
assign n_2973 = n_150 & ~n_2956;
assign n_2974 = ~n_2956 & n_130;
assign n_2975 = n_2956 ^ n_103;
assign n_2976 = n_2956 ^ n_2864;
assign n_2977 = ~n_2956 & n_115;
assign n_2978 = n_1 & ~n_2956;
assign n_2979 = ~n_2900 ^ ~n_2957;
assign n_2980 = n_2902 ^ n_2958;
assign n_2981 = ~n_2903 ^ ~n_2960;
assign n_2982 = n_157 & ~n_2962;
assign n_2983 = n_2839 & n_2964;
assign n_2984 = n_2917 & ~n_2965;
assign n_2985 = n_134 & n_2967;
assign n_2986 = n_2968 ^ n_1909;
assign n_2987 = n_2969 & ~n_2953;
assign n_2988 = n_2952 & n_2970;
assign n_2989 = ~n_2971 & ~n_2929;
assign n_2990 = n_2971 & ~n_2930;
assign n_2991 = ~n_2971 & n_234;
assign n_2992 = ~n_2971 & n_301;
assign n_2993 = ~n_2971 & n_198;
assign n_2994 = ~n_2971 & n_197;
assign n_2995 = ~n_2971 & n_98;
assign n_2996 = ~n_2971 & ~n_130;
assign n_2997 = ~n_2971 & n_431;
assign n_2998 = ~n_2971 & ~n_96;
assign n_2999 = n_0 & n_2971;
assign n_3000 = ~n_2971 & ~n_48;
assign n_3001 = n_2972 ^ n_2971;
assign n_3002 = n_2973 ^ n_2971;
assign n_3003 = n_100 & n_2974;
assign n_3004 = ~n_2974 & ~n_2975;
assign n_3005 = n_231 & ~n_2976;
assign n_3006 = n_2977 ^ n_2971;
assign n_3007 = n_2978 ^ n_2971;
assign n_3008 = ~n_2979 & ~n_2916;
assign n_3009 = ~n_2979 ^ n_2945;
assign n_3010 = ~n_2981 & n_2966;
assign n_3011 = ~n_2981 ^ n_2948;
assign n_3012 = n_2940 ^ n_2982;
assign n_3013 = n_88 ^ n_2983;
assign n_3014 = n_2898 ^ n_2984;
assign n_3015 = n_134 ^ n_2985;
assign n_3016 = n_2980 ^ n_2985;
assign n_3017 = n_2794 ^ n_2987;
assign n_3018 = n_2759 ^ n_2987;
assign n_3019 = n_2617 ^ n_2987;
assign n_3020 = n_2780 ^ n_2987;
assign n_3021 = n_2988 ^ n_2955;
assign n_3022 = n_2989 ^ n_2990;
assign n_3023 = ~n_2991 ^ ~n_2932;
assign n_3024 = ~n_2994 ^ ~n_2933;
assign n_3025 = n_2996 ^ n_2938;
assign n_3026 = n_2998 ^ n_2941;
assign n_3027 = n_2999 ^ n_2944;
assign n_3028 = n_163 & n_3001;
assign n_3029 = n_122 & ~n_3002;
assign n_3030 = n_2995 ^ n_3004;
assign n_3031 = n_3005 ^ n_2864;
assign n_3032 = ~n_157 & ~n_3006;
assign n_3033 = x0 & ~n_3007;
assign n_3034 = n_3008 ^ n_2839;
assign n_3035 = ~n_3008 & ~n_2848;
assign n_3036 = n_2854 ^ n_3010;
assign n_3037 = n_3010 & n_2854;
assign n_3038 = n_3012 ^ n_2922;
assign n_3039 = n_3012 & n_2897;
assign n_3040 = n_141 & n_3013;
assign n_3041 = n_3015 & ~n_2980;
assign n_3042 = n_3017 & n_2795;
assign n_3043 = n_2771 & ~n_3018;
assign n_3044 = n_2780 & ~n_3019;
assign n_3045 = n_3020 ^ n_1911;
assign n_3046 = n_3021 ^ n_1909;
assign n_3047 = n_3021 ^ n_2986;
assign n_3048 = n_207 & ~n_3022;
assign n_3049 = n_122 & ~n_3022;
assign n_3050 = ~n_103 & ~n_3022;
assign n_3051 = ~n_3022 & n_107;
assign n_3052 = ~n_3022 & n_115;
assign n_3053 = n_134 ^ ~n_3024;
assign n_3054 = n_3026 ^ n_87;
assign n_3055 = ~n_3014 ^ ~n_3028;
assign n_3056 = ~n_2959 ^ ~n_3029;
assign n_3057 = n_3003 ^ n_3031;
assign n_3058 = ~n_2961 ^ ~n_3032;
assign n_3059 = ~n_2963 ^ ~n_3033;
assign n_3060 = n_3036 ^ n_3037;
assign n_3061 = n_87 ^ n_3039;
assign n_3062 = n_2860 ^ n_3040;
assign n_3063 = ~n_2850 & ~n_3041;
assign n_3064 = n_3043 ^ n_2591;
assign n_3065 = n_2789 ^ n_3044;
assign n_3066 = n_2986 & n_3046;
assign n_3067 = ~n_3047 & ~n_2989;
assign n_3068 = n_3047 & ~n_2990;
assign n_3069 = n_3047 & n_234;
assign n_3070 = n_3047 & n_198;
assign n_3071 = n_3047 & n_197;
assign n_3072 = n_3047 & n_122;
assign n_3073 = n_3047 ^ n_121;
assign n_3074 = n_3047 & n_431;
assign n_3075 = n_3047 & n_260;
assign n_3076 = n_3047 & ~n_48;
assign n_3077 = n_3022 ^ n_3047;
assign n_3078 = n_3047 & ~n_75;
assign n_3079 = n_0 & n_3047;
assign n_3080 = n_3047 & n_208;
assign n_3081 = n_187 & n_3047;
assign n_3082 = n_3048 ^ n_3047;
assign n_3083 = n_3050 ^ n_3047;
assign n_3084 = n_3052 ^ n_87;
assign n_3085 = ~n_3055 ^ n_187;
assign n_3086 = n_3055 & ~n_3035;
assign n_3087 = ~n_3056 ^ n_134;
assign n_3088 = n_2936 ^ n_3057;
assign n_3089 = ~n_3058 & ~n_3039;
assign n_3090 = n_2858 ^ ~n_3058;
assign n_3091 = n_3061 ^ ~n_3058;
assign n_3092 = n_3059 & n_3062;
assign n_3093 = n_3064 ^ n_2647;
assign n_3094 = n_3065 ^ n_2647;
assign n_3095 = n_3066 ^ n_2968;
assign n_3096 = n_3067 ^ n_3068;
assign n_3097 = ~n_3069 ^ ~n_2992;
assign n_3098 = ~n_3071 ^ ~n_2993;
assign n_3099 = n_3022 & n_3072;
assign n_3100 = ~n_3053 ^ n_3073;
assign n_3101 = n_3075 ^ n_2997;
assign n_3102 = ~n_60 & ~n_3077;
assign n_3103 = n_3078 ^ x0;
assign n_3104 = n_163 & n_3082;
assign n_3105 = n_98 & n_3083;
assign n_3106 = n_3084 ^ n_3047;
assign n_3107 = n_3008 & n_3085;
assign n_3108 = n_2864 ^ n_3086;
assign n_3109 = n_3087 ^ n_2850;
assign n_3110 = n_3041 & n_3087;
assign n_3111 = ~n_3063 & ~n_3087;
assign n_3112 = n_3030 ^ n_3088;
assign n_3113 = n_3089 ^ n_90;
assign n_3114 = ~n_3089 & n_3090;
assign n_3115 = n_3040 ^ n_3092;
assign n_3116 = n_2669 & n_3093;
assign n_3117 = n_3094 ^ n_1903;
assign n_3118 = n_3095 ^ n_3020;
assign n_3119 = n_3095 ^ n_3045;
assign n_3120 = n_207 & ~n_3096;
assign n_3121 = ~n_121 & ~n_3096;
assign n_3122 = n_130 & ~n_3096;
assign n_3123 = ~n_100 & ~n_3096;
assign n_3124 = n_3096 ^ n_2971;
assign n_3125 = ~n_157 & ~n_3096;
assign n_3126 = ~n_3096 & ~n_3098;
assign n_3127 = ~n_3098 ^ n_134;
assign n_3128 = ~n_3099 ^ ~n_3024;
assign n_3129 = n_3100 ^ n_3073;
assign n_3130 = n_3101 ^ n_87;
assign n_3131 = n_87 & ~n_3101;
assign n_3132 = n_3027 ^ n_3103;
assign n_3133 = ~n_3023 ^ ~n_3104;
assign n_3134 = n_103 ^ n_3105;
assign n_3135 = n_3106 ^ n_3054;
assign n_3136 = n_3107 ^ n_187;
assign n_3137 = ~n_3108 & ~n_3086;
assign n_3138 = n_3109 ^ n_3041;
assign n_3139 = n_2947 ^ n_3111;
assign n_3140 = n_3112 & n_3060;
assign n_3141 = n_3060 ^ n_3112;
assign n_3142 = n_3113 ^ n_3091;
assign n_3143 = n_2871 ^ n_3114;
assign n_3144 = n_3115 ^ n_2909;
assign n_3145 = n_2618 ^ n_3116;
assign n_3146 = ~n_3045 & n_3118;
assign n_3147 = ~n_3119 & ~n_3067;
assign n_3148 = n_3119 & ~n_3068;
assign n_3149 = ~n_3119 & n_198;
assign n_3150 = ~n_3119 & n_197;
assign n_3151 = n_3119 & n_152;
assign n_3152 = ~n_3119 & ~n_231;
assign n_3153 = ~n_3119 & n_98;
assign n_3154 = ~n_3119 & n_431;
assign n_3155 = ~n_3119 & n_260;
assign n_3156 = n_3119 ^ n_74;
assign n_3157 = ~n_3119 & ~n_48;
assign n_3158 = n_0 & ~n_3119;
assign n_3159 = n_3096 ^ n_3119;
assign n_3160 = ~n_3119 & ~n_75;
assign n_3161 = n_165 & ~n_3119;
assign n_3162 = n_3081 ^ n_3119;
assign n_3163 = ~n_3119 & n_301;
assign n_3164 = n_3120 ^ n_3119;
assign n_3165 = ~n_3119 ^ ~n_3121;
assign n_3166 = n_231 & n_3124;
assign n_3167 = n_3126 ^ n_122;
assign n_3168 = ~n_134 & n_3128;
assign n_3169 = ~n_3072 ^ n_3129;
assign n_3170 = n_3130 ^ n_3131;
assign n_3171 = n_3132 ^ n_128;
assign n_3172 = ~n_3133 ^ n_3086;
assign n_3173 = n_3134 ^ n_3051;
assign n_3174 = n_157 & n_3135;
assign n_3175 = n_3034 & ~n_3136;
assign n_3176 = n_187 & n_3137;
assign n_3177 = n_3138 & ~n_3110;
assign n_3178 = n_3140 ^ n_2949;
assign n_3179 = ~n_3037 ^ ~n_3141;
assign n_3180 = n_2839 & n_3142;
assign n_3181 = n_2905 ^ n_3143;
assign n_3182 = ~n_3145 & ~n_3042;
assign n_3183 = n_3146 ^ n_3095;
assign n_3184 = n_3147 ^ n_3148;
assign n_3185 = ~n_3150 ^ ~n_3070;
assign n_3186 = ~n_3096 & n_3151;
assign n_3187 = n_3155 ^ n_3074;
assign n_3188 = ~n_3156 & n_3125;
assign n_3189 = ~n_60 & n_3159;
assign n_3190 = n_3160 ^ n_3000;
assign n_3191 = n_3080 ^ n_3161;
assign n_3192 = n_134 & ~n_3162;
assign n_3193 = n_163 & ~n_3164;
assign n_3194 = n_3166 ^ n_2971;
assign n_3195 = ~n_134 & n_3167;
assign n_3196 = ~n_3169 ^ n_3073;
assign n_3197 = n_3102 ^ n_3171;
assign n_3198 = n_3108 & ~n_3172;
assign n_3199 = n_3173 ^ n_3025;
assign n_3200 = n_3106 ^ n_3174;
assign n_3201 = ~n_3055 ^ n_3175;
assign n_3202 = n_3108 ^ n_3176;
assign n_3203 = n_3180 ^ n_3113;
assign n_3204 = n_2776 & ~n_3182;
assign n_3205 = n_2709 ^ n_3182;
assign n_3206 = n_2775 & ~n_3182;
assign n_3207 = n_3183 ^ n_3094;
assign n_3208 = n_3183 ^ n_3117;
assign n_3209 = n_122 & ~n_3184;
assign n_3210 = n_3184 ^ n_3067;
assign n_3211 = n_130 & ~n_3184;
assign n_3212 = n_100 & ~n_3184;
assign n_3213 = n_3184 ^ n_3047;
assign n_3214 = n_3184 ^ n_3068;
assign n_3215 = n_74 & ~n_3184;
assign n_3216 = n_207 & ~n_3184;
assign n_3217 = ~n_3185 ^ n_134;
assign n_3218 = n_134 ^ n_3186;
assign n_3219 = ~n_3184 & ~n_3187;
assign n_3220 = n_3187 ^ n_87;
assign n_3221 = n_3079 ^ n_3190;
assign n_3222 = ~n_134 & n_3191;
assign n_3223 = n_3119 ^ n_3192;
assign n_3224 = ~n_3097 ^ ~n_3193;
assign n_3225 = n_3194 ^ n_3047;
assign n_3226 = n_122 ^ n_3195;
assign n_3227 = ~n_3049 & n_3196;
assign n_3228 = n_3197 ^ n_2909;
assign n_3229 = n_3198 ^ n_2864;
assign n_3230 = n_3199 ^ n_2949;
assign n_3231 = n_3199 ^ n_3178;
assign n_3232 = n_3200 ^ n_2905;
assign n_3233 = n_3200 ^ n_3181;
assign n_3234 = ~n_3133 ^ n_3202;
assign n_3235 = n_3204 ^ n_2741;
assign n_3236 = n_3205 ^ ~n_2019;
assign n_3237 = ~n_3206 & ~n_2769;
assign n_3238 = n_3117 & ~n_3207;
assign n_3239 = ~n_3208 & ~n_3147;
assign n_3240 = n_3208 & ~n_3148;
assign n_3241 = n_3208 & n_198;
assign n_3242 = n_3208 & n_197;
assign n_3243 = n_3208 ^ n_121;
assign n_3244 = n_3184 ^ n_3208;
assign n_3245 = n_3208 & ~n_130;
assign n_3246 = n_3208 & n_98;
assign n_3247 = n_3208 & n_431;
assign n_3248 = n_3208 & n_260;
assign n_3249 = n_22 & n_3208;
assign n_3250 = n_0 & n_3208;
assign n_3251 = n_3208 & ~n_75;
assign n_3252 = n_3208 & n_234;
assign n_3253 = n_3208 & n_301;
assign n_3254 = ~n_187 & n_3208;
assign n_3255 = n_122 & n_3210;
assign n_3256 = n_3210 ^ n_103;
assign n_3257 = ~n_157 & n_3210;
assign n_3258 = n_231 & ~n_3213;
assign n_3259 = ~n_3214 & ~n_224;
assign n_3260 = n_3208 ^ ~n_3215;
assign n_3261 = n_3216 ^ n_3208;
assign n_3262 = ~n_134 ^ n_3218;
assign n_3263 = n_3219 ^ n_157;
assign n_3264 = n_3221 ^ n_141;
assign n_3265 = n_3161 ^ n_3222;
assign n_3266 = ~n_165 & ~n_3223;
assign n_3267 = ~n_3224 ^ n_2915;
assign n_3268 = n_3123 ^ n_3225;
assign n_3269 = ~n_3165 & n_3226;
assign n_3270 = n_3073 ^ n_3227;
assign n_3271 = n_3144 & n_3228;
assign n_3272 = n_3229 ^ n_2915;
assign n_3273 = n_3178 & ~n_3230;
assign n_3274 = n_3181 & ~n_3232;
assign n_3275 = n_2755 & ~n_3235;
assign n_3276 = n_2711 ^ n_3237;
assign n_3277 = n_2726 ^ n_3237;
assign n_3278 = n_3238 ^ n_3183;
assign n_3279 = n_3239 ^ n_3240;
assign n_3280 = ~n_3242 ^ ~n_3149;
assign n_3281 = n_3209 & ~n_3243;
assign n_3282 = ~n_60 & ~n_3244;
assign n_3283 = n_3245 ^ n_3152;
assign n_3284 = n_3248 ^ n_3154;
assign n_3285 = n_3250 ^ n_3157;
assign n_3286 = n_3251 ^ n_3076;
assign n_3287 = ~n_3252 ^ ~n_3163;
assign n_3288 = n_3255 ^ n_134;
assign n_3289 = n_3256 ^ n_130;
assign n_3290 = n_3131 & ~n_3257;
assign n_3291 = n_3258 ^ n_3047;
assign n_3292 = ~n_3259 ^ ~n_3170;
assign n_3293 = ~n_3262 ^ n_134;
assign n_3294 = n_87 & ~n_3263;
assign n_3295 = n_3189 ^ n_3264;
assign n_3296 = n_3261 ^ n_3265;
assign n_3297 = n_3261 ^ n_3266;
assign n_3298 = n_3268 ^ n_3194;
assign n_3299 = ~n_3270 & ~n_3168;
assign n_3300 = n_3115 ^ n_3271;
assign n_3301 = ~n_187 & n_3272;
assign n_3302 = ~n_3272 & ~n_3267;
assign n_3303 = n_3273 ^ n_3140;
assign n_3304 = n_3274 ^ n_3143;
assign n_3305 = n_2623 ^ n_3275;
assign n_3306 = n_2726 & n_3276;
assign n_3307 = ~n_1886 ^ n_3277;
assign n_3308 = n_3278 ^ n_3205;
assign n_3309 = n_3278 ^ n_3236;
assign n_3310 = n_122 & ~n_3279;
assign n_3311 = n_3279 ^ n_3147;
assign n_3312 = n_98 & ~n_3279;
assign n_3313 = ~n_157 & ~n_3279;
assign n_3314 = n_1 & ~n_3279;
assign n_3315 = n_207 & ~n_3279;
assign n_3316 = n_134 ^ ~n_3280;
assign n_3317 = n_103 ^ ~n_3283;
assign n_3318 = n_3284 ^ n_87;
assign n_3319 = n_3158 ^ n_3286;
assign n_3320 = n_3289 ^ n_3214;
assign n_3321 = n_3291 ^ n_3119;
assign n_3322 = ~n_3292 ^ ~n_3188;
assign n_3323 = ~n_3288 & ~n_3293;
assign n_3324 = n_157 ^ n_3294;
assign n_3325 = n_3295 ^ n_3038;
assign n_3326 = n_3296 ^ n_3261;
assign n_3327 = n_3297 ^ n_3261;
assign n_3328 = n_130 & ~n_3298;
assign n_3329 = n_2947 ^ n_3299;
assign n_3330 = n_3038 ^ n_3300;
assign n_3331 = n_3301 ^ ~n_3224;
assign n_3332 = n_3302 ^ n_2915;
assign n_3333 = n_3016 ^ n_3303;
assign n_3334 = n_3304 ^ n_3011;
assign n_3335 = n_3305 ^ n_1907;
assign n_3336 = n_3306 ^ n_3237;
assign n_3337 = n_3236 & ~n_3308;
assign n_3338 = n_3309 & ~n_3239;
assign n_3339 = ~n_3309 & ~n_3240;
assign n_3340 = n_3309 & n_197;
assign n_3341 = n_3309 ^ n_121;
assign n_3342 = n_3309 & ~n_130;
assign n_3343 = n_3309 ^ n_100;
assign n_3344 = n_3309 & n_431;
assign n_3345 = n_3309 & n_260;
assign n_3346 = n_3309 ^ n_74;
assign n_3347 = x1 & n_3309;
assign n_3348 = n_3309 & ~n_48;
assign n_3349 = n_3309 & n_198;
assign n_3350 = n_3309 & n_234;
assign n_3351 = n_3309 & n_301;
assign n_3352 = ~n_187 & n_3309;
assign n_3353 = n_3309 & n_3208;
assign n_3354 = ~n_3311 & n_173;
assign n_3355 = n_3244 ^ n_3311;
assign n_3356 = n_3311 ^ n_103;
assign n_3357 = n_3312 ^ n_3283;
assign n_3358 = n_3314 ^ n_3309;
assign n_3359 = n_3315 ^ n_3309;
assign n_3360 = n_3319 ^ n_141;
assign n_3361 = ~n_3320 & n_3122;
assign n_3362 = n_3212 ^ n_3321;
assign n_3363 = ~n_3322 ^ ~n_3290;
assign n_3364 = ~n_3262 ^ n_3323;
assign n_3365 = ~n_3260 & ~n_3324;
assign n_3366 = ~n_3326 ^ ~n_3327;
assign n_3367 = n_3225 ^ n_3328;
assign n_3368 = ~n_3329 & ~n_3139;
assign n_3369 = n_3329 ^ n_3111;
assign n_3370 = ~n_3330 & n_3325;
assign n_3371 = ~n_187 & ~n_3332;
assign n_3372 = n_3336 ^ n_2586;
assign n_3373 = n_3336 ^ n_2199;
assign n_3374 = n_3336 & ~n_2619;
assign n_3375 = n_3337 ^ n_3278;
assign n_3376 = n_3338 ^ n_3339;
assign n_3377 = ~n_3340 ^ ~n_3241;
assign n_3378 = n_3310 & n_3341;
assign n_3379 = n_3312 & ~n_3343;
assign n_3380 = n_3345 ^ n_3247;
assign n_3381 = n_3313 & ~n_3346;
assign n_3382 = n_3249 ^ n_3347;
assign n_3383 = ~n_3350 ^ ~n_3253;
assign n_3384 = ~n_3254 & ~n_3352;
assign n_3385 = n_3355 ^ n_3208;
assign n_3386 = n_3355 & ~n_199;
assign n_3387 = x0 & n_3358;
assign n_3388 = n_163 & n_3359;
assign n_3389 = n_3360 ^ n_3282;
assign n_3390 = n_3320 ^ n_3361;
assign n_3391 = n_3362 ^ n_3291;
assign n_3392 = ~n_3363 ^ n_3011;
assign n_3393 = n_3364 ^ n_134;
assign n_3394 = ~n_3366 ^ n_3261;
assign n_3395 = n_3368 ^ n_3299;
assign n_3396 = n_3300 ^ n_3370;
assign n_3397 = n_2971 ^ n_3371;
assign n_3398 = n_3372 ^ n_1878;
assign n_3399 = n_2586 & n_3373;
assign n_3400 = n_1910 ^ n_3374;
assign n_3401 = n_3375 ^ n_3305;
assign n_3402 = n_3375 ^ n_3335;
assign n_3403 = n_122 & ~n_3376;
assign n_3404 = n_3376 ^ n_3239;
assign n_3405 = ~n_3376 & n_130;
assign n_3406 = n_3376 ^ n_3208;
assign n_3407 = ~n_157 & ~n_3376;
assign n_3408 = n_3376 ^ n_3240;
assign n_3409 = n_1 & ~n_3376;
assign n_3410 = n_207 & ~n_3376;
assign n_3411 = n_134 ^ ~n_3377;
assign n_3412 = n_3380 ^ n_87;
assign n_3413 = ~n_87 & n_3380;
assign n_3414 = n_122 & n_3385;
assign n_3415 = n_3385 ^ n_3356;
assign n_3416 = n_201 & n_3385;
assign n_3417 = ~n_3285 ^ ~n_3387;
assign n_3418 = ~n_3287 ^ ~n_3388;
assign n_3419 = n_3203 ^ n_3389;
assign n_3420 = n_3153 ^ n_3390;
assign n_3421 = n_130 & n_3391;
assign n_3422 = n_3392 & n_3334;
assign n_3423 = n_3304 ^ n_3392;
assign n_3424 = n_3393 ^ n_3186;
assign n_3425 = ~n_163 & ~n_3394;
assign n_3426 = n_3009 ^ n_3395;
assign n_3427 = n_3396 ^ n_3203;
assign n_3428 = ~n_187 & n_3397;
assign n_3429 = ~n_3335 & n_3401;
assign n_3430 = n_3402 & ~n_3338;
assign n_3431 = ~n_3402 & ~n_3339;
assign n_3432 = n_3402 ^ n_121;
assign n_3433 = ~n_3402 & n_98;
assign n_3434 = n_87 & ~n_3402;
assign n_3435 = ~n_3402 & n_531;
assign n_3436 = ~n_3402 & n_260;
assign n_3437 = n_3402 ^ n_74;
assign n_3438 = ~n_3402 & ~n_48;
assign n_3439 = n_0 & ~n_3402;
assign n_3440 = ~n_3402 & n_197;
assign n_3441 = ~n_3402 & n_198;
assign n_3442 = ~n_3402 & n_234;
assign n_3443 = ~n_187 & ~n_3402;
assign n_3444 = ~n_3402 & ~n_237;
assign n_3445 = ~n_3402 & ~n_141;
assign n_3446 = n_122 & n_3404;
assign n_3447 = n_3404 & n_98;
assign n_3448 = ~n_157 & n_3404;
assign n_3449 = ~n_3405 & n_144;
assign n_3450 = n_100 & n_3405;
assign n_3451 = ~n_231 & ~n_3406;
assign n_3452 = n_201 & ~n_3408;
assign n_3453 = n_3409 ^ n_3402;
assign n_3454 = n_3410 ^ n_3402;
assign n_3455 = n_3412 ^ n_3413;
assign n_3456 = ~n_134 & n_3414;
assign n_3457 = n_3415 ^ n_130;
assign n_3458 = ~n_3386 ^ ~n_3416;
assign n_3459 = ~n_3417 ^ n_141;
assign n_3460 = ~n_3418 ^ n_3047;
assign n_3461 = n_3420 ^ n_3367;
assign n_3462 = n_3321 ^ n_3421;
assign n_3463 = n_3422 ^ ~n_3363;
assign n_3464 = n_3127 ^ n_3424;
assign n_3465 = n_3261 ^ n_3425;
assign n_3466 = ~n_3419 & n_3427;
assign n_3467 = n_3429 ^ n_3375;
assign n_3468 = n_3430 ^ n_3431;
assign n_3469 = n_3403 & ~n_3432;
assign n_3470 = n_3436 ^ n_3344;
assign n_3471 = n_3407 & ~n_3437;
assign n_3472 = n_3439 ^ n_3348;
assign n_3473 = ~n_3440 ^ ~n_3349;
assign n_3474 = ~n_3442 ^ ~n_3351;
assign n_3475 = n_3443 ^ n_3402;
assign n_3476 = ~n_3443 & n_3384;
assign n_3477 = ~n_206 & ~n_3444;
assign n_3478 = n_3310 ^ n_3446;
assign n_3479 = ~n_3446 & ~n_3316;
assign n_3480 = n_3357 ^ n_3447;
assign n_3481 = ~n_3447 & ~n_3317;
assign n_3482 = n_3448 ^ n_3284;
assign n_3483 = n_3449 ^ n_3433;
assign n_3484 = n_3450 ^ n_130;
assign n_3485 = n_3452 ^ n_3448;
assign n_3486 = n_3453 ^ n_3382;
assign n_3487 = n_163 & ~n_3454;
assign n_3488 = n_3354 ^ n_3456;
assign n_3489 = n_3457 & n_3211;
assign n_3490 = n_3220 ^ ~n_3458;
assign n_3491 = n_3459 ^ n_3233;
assign n_3492 = n_3461 ^ n_3016;
assign n_3493 = n_3461 ^ n_3333;
assign n_3494 = n_3463 ^ ~n_3179;
assign n_3495 = ~n_3464 ^ n_3186;
assign n_3496 = n_3428 ^ n_3465;
assign n_3497 = n_3465 ^ n_3371;
assign n_3498 = n_3389 ^ n_3466;
assign n_3499 = n_3277 ^ n_3467;
assign n_3500 = n_3468 ^ n_3339;
assign n_3501 = n_130 & ~n_3468;
assign n_3502 = n_3468 ^ n_3309;
assign n_3503 = n_3468 ^ n_231;
assign n_3504 = n_100 & ~n_3468;
assign n_3505 = ~n_157 & ~n_3468;
assign n_3506 = n_3468 ^ n_3338;
assign n_3507 = n_1 & ~n_3468;
assign n_3508 = n_122 & ~n_3468;
assign n_3509 = n_163 & ~n_3468;
assign n_3510 = n_3470 ^ n_87;
assign n_3511 = ~n_87 & ~n_3470;
assign n_3512 = ~n_3473 ^ n_134;
assign n_3513 = n_187 ^ ~n_3474;
assign n_3514 = ~n_3280 ^ ~n_3478;
assign n_3515 = ~n_3479 ^ ~n_3378;
assign n_3516 = ~n_103 & n_3480;
assign n_3517 = ~n_3481 ^ ~n_3379;
assign n_3518 = n_3484 ^ n_3451;
assign n_3519 = ~n_3482 & n_3485;
assign n_3520 = ~x0 & ~n_3486;
assign n_3521 = ~n_3383 ^ ~n_3487;
assign n_3522 = n_3217 & ~n_3488;
assign n_3523 = n_3457 ^ n_3489;
assign n_3524 = ~n_3490 ^ n_3386;
assign n_3525 = ~n_3333 & n_3492;
assign n_3526 = ~n_3495 & ~n_3269;
assign n_3527 = ~n_3397 & n_3497;
assign n_3528 = n_3498 ^ n_3233;
assign n_3529 = ~n_3499 & n_3307;
assign n_3530 = ~n_1886 ^ n_3499;
assign n_3531 = n_122 & n_3500;
assign n_3532 = ~n_157 & n_3500;
assign n_3533 = ~n_103 & n_3501;
assign n_3534 = n_3501 ^ n_3503;
assign n_3535 = n_3504 ^ n_3431;
assign n_3536 = ~n_224 & ~n_3506;
assign n_3537 = n_3510 ^ n_3511;
assign n_3538 = ~n_134 & n_3514;
assign n_3539 = ~n_3516 & ~n_3517;
assign n_3540 = n_3342 ^ n_3518;
assign n_3541 = n_3519 ^ n_3452;
assign n_3542 = n_3453 ^ n_3520;
assign n_3543 = n_3354 ^ n_3522;
assign n_3544 = n_3246 ^ n_3523;
assign n_3545 = ~n_3524 & ~n_3365;
assign n_3546 = n_3525 ^ n_3461;
assign n_3547 = n_3009 ^ n_3526;
assign n_3548 = n_3527 ^ n_2971;
assign n_3549 = ~n_3491 & ~n_3528;
assign n_3550 = n_3529 ^ n_3467;
assign n_3551 = n_3530 & ~n_3430;
assign n_3552 = ~n_3530 & ~n_3431;
assign n_3553 = n_3530 & ~n_130;
assign n_3554 = n_3530 & n_98;
assign n_3555 = ~n_3530 & n_614;
assign n_3556 = n_3434 ^ n_3530;
assign n_3557 = n_3530 & ~n_225;
assign n_3558 = n_3530 ^ n_74;
assign n_3559 = n_22 & n_3530;
assign n_3560 = n_0 & n_3530;
assign n_3561 = n_3507 ^ n_3530;
assign n_3562 = n_3530 ^ n_121;
assign n_3563 = n_3530 & n_197;
assign n_3564 = n_3530 & n_198;
assign n_3565 = n_3530 ^ n_165;
assign n_3566 = n_3475 ^ n_3530;
assign n_3567 = ~n_165 & ~n_3530;
assign n_3568 = ~n_187 & ~n_3530;
assign n_3569 = n_3403 ^ n_3531;
assign n_3570 = ~n_3531 & ~n_3411;
assign n_3571 = ~n_3532 & n_3455;
assign n_3572 = n_3533 ^ n_103;
assign n_3573 = ~n_3502 & n_3534;
assign n_3574 = n_130 & n_3535;
assign n_3575 = ~n_3413 ^ ~n_3536;
assign n_3576 = ~n_3538 & ~n_3515;
assign n_3577 = n_3369 ^ n_3539;
assign n_3578 = n_3483 ^ n_3540;
assign n_3579 = n_3541 ^ n_3448;
assign n_3580 = n_3542 ^ n_141;
assign n_3581 = ~n_3543 ^ ~n_3281;
assign n_3582 = n_3544 ^ n_3462;
assign n_3583 = ~n_3179 ^ n_3545;
assign n_3584 = ~n_3547 & ~n_3426;
assign n_3585 = n_3547 ^ n_3395;
assign n_3586 = n_3548 ^ n_3047;
assign n_3587 = n_3459 ^ n_3549;
assign n_3588 = n_3550 ^ n_3372;
assign n_3589 = n_3550 ^ n_3398;
assign n_3590 = n_3552 ^ n_3431;
assign n_3591 = n_3555 ^ n_202;
assign n_3592 = ~n_74 & n_3556;
assign n_3593 = n_3557 ^ n_3435;
assign n_3594 = ~n_3558 & n_3505;
assign n_3595 = n_3560 ^ n_3438;
assign n_3596 = x0 & n_3561;
assign n_3597 = ~n_3562 & n_3508;
assign n_3598 = ~n_3563 ^ ~n_3441;
assign n_3599 = n_3509 & n_3565;
assign n_3600 = ~n_165 & ~n_3566;
assign n_3601 = n_240 & n_3567;
assign n_3602 = ~n_3567 & ~n_3477;
assign n_3603 = ~n_232 & ~n_3568;
assign n_3604 = n_3568 ^ n_187;
assign n_3605 = ~n_3377 ^ ~n_3569;
assign n_3606 = ~n_3570 ^ ~n_3469;
assign n_3607 = ~n_3571 ^ ~n_3471;
assign n_3608 = n_3572 ^ n_3573;
assign n_3609 = n_3431 ^ n_3574;
assign n_3610 = n_3234 ^ n_3576;
assign n_3611 = n_3579 ^ n_3452;
assign n_3612 = ~n_3581 ^ n_3201;
assign n_3613 = n_3582 ^ n_3177;
assign n_3614 = n_3546 ^ n_3582;
assign n_3615 = n_3583 & ~n_3494;
assign n_3616 = n_3463 ^ n_3583;
assign n_3617 = n_3584 ^ n_3526;
assign n_3618 = n_3585 ^ n_3578;
assign n_3619 = ~n_187 & n_3586;
assign n_3620 = ~n_3586 & n_3460;
assign n_3621 = n_3587 ^ n_3423;
assign n_3622 = ~n_3423 & n_3587;
assign n_3623 = ~n_3398 & n_3588;
assign n_3624 = n_3589 & ~n_3551;
assign n_3625 = ~n_3589 & ~n_3552;
assign n_3626 = ~n_3589 & n_98;
assign n_3627 = ~n_3589 & ~n_130;
assign n_3628 = ~n_3589 & n_743;
assign n_3629 = n_3589 ^ n_74;
assign n_3630 = n_3589 & n_202;
assign n_3631 = ~n_3589 & n_531;
assign n_3632 = n_22 & n_3589;
assign n_3633 = x1 & ~n_3589;
assign n_3634 = x0 & ~n_3589;
assign n_3635 = ~n_3589 & ~n_231;
assign n_3636 = n_3589 ^ n_121;
assign n_3637 = ~n_3589 & n_197;
assign n_3638 = ~n_3589 & n_198;
assign n_3639 = n_3589 ^ n_165;
assign n_3640 = n_3589 ^ n_187;
assign n_3641 = ~n_187 & ~n_3589;
assign n_3642 = ~n_3589 & n_301;
assign n_3643 = n_3589 ^ n_103;
assign n_3644 = n_3590 ^ n_3551;
assign n_3645 = ~n_228 & n_3591;
assign n_3646 = n_3530 ^ n_3592;
assign n_3647 = ~n_3472 ^ ~n_3596;
assign n_3648 = ~n_3598 ^ n_134;
assign n_3649 = n_3600 ^ n_3530;
assign n_3650 = n_3601 ^ n_3603;
assign n_3651 = n_3604 ^ n_141;
assign n_3652 = ~n_134 & n_3605;
assign n_3653 = ~n_3607 ^ ~n_3575;
assign n_3654 = n_3554 ^ n_3608;
assign n_3655 = ~n_3318 & ~n_3611;
assign n_3656 = n_3546 ^ n_3613;
assign n_3657 = n_3613 & n_3614;
assign n_3658 = n_3615 ^ n_3545;
assign n_3659 = n_3201 ^ n_3617;
assign n_3660 = n_3612 ^ n_3617;
assign n_3661 = n_3619 ^ ~n_3418;
assign n_3662 = n_3620 ^ n_3047;
assign n_3663 = n_3621 ^ n_3622;
assign n_3664 = n_3623 ^ n_3550;
assign n_3665 = n_3624 ^ n_3625;
assign n_3666 = n_3628 ^ n_613;
assign n_3667 = n_3630 ^ n_179;
assign n_3668 = n_3633 ^ n_3559;
assign n_3669 = ~n_3637 ^ ~n_3564;
assign n_3670 = ~n_3640 & n_238;
assign n_3671 = n_206 & n_3641;
assign n_3672 = n_3468 ^ n_3644;
assign n_3673 = n_201 & ~n_3644;
assign n_3674 = ~n_3644 & n_173;
assign n_3675 = n_228 ^ n_3645;
assign n_3676 = ~n_179 & n_3646;
assign n_3677 = ~n_3647 ^ n_3542;
assign n_3678 = ~n_3647 ^ n_141;
assign n_3679 = n_164 & n_3649;
assign n_3680 = n_160 & ~n_3651;
assign n_3681 = ~n_3652 & ~n_3606;
assign n_3682 = ~n_3653 ^ n_3493;
assign n_3683 = n_3654 ^ n_3609;
assign n_3684 = n_3452 ^ n_3655;
assign n_3685 = n_3657 ^ n_3546;
assign n_3686 = n_3658 ^ n_3231;
assign n_3687 = n_3612 & ~n_3659;
assign n_3688 = n_3662 ^ n_3119;
assign n_3689 = ~n_187 & n_3662;
assign n_3690 = n_3664 ^ n_1910;
assign n_3691 = n_3664 & n_1910;
assign n_3692 = n_3665 ^ n_3551;
assign n_3693 = n_130 & n_3665;
assign n_3694 = n_3665 ^ n_3530;
assign n_3695 = ~n_3665 & n_115;
assign n_3696 = n_1 & ~n_3665;
assign n_3697 = n_207 & n_3665;
assign n_3698 = n_134 ^ ~n_3669;
assign n_3699 = n_3671 ^ n_3650;
assign n_3700 = n_3672 ^ n_3430;
assign n_3701 = ~n_157 & n_3672;
assign n_3702 = n_122 & n_3672;
assign n_3703 = n_163 & n_3672;
assign n_3704 = ~n_3673 ^ n_3537;
assign n_3705 = ~n_3666 & n_3675;
assign n_3706 = ~n_3593 ^ ~n_3676;
assign n_3707 = ~n_3616 ^ n_3677;
assign n_3708 = n_3678 ^ n_3616;
assign n_3709 = n_3678 ^ n_3622;
assign n_3710 = ~n_3679 ^ ~n_3602;
assign n_3711 = n_3680 ^ n_87;
assign n_3712 = n_3331 ^ n_3681;
assign n_3713 = n_3660 ^ n_3683;
assign n_3714 = ~n_3684 ^ ~n_3381;
assign n_3715 = n_3685 ^ n_3539;
assign n_3716 = n_3685 ^ n_3577;
assign n_3717 = n_3687 ^ ~n_3581;
assign n_3718 = ~n_187 & n_3688;
assign n_3719 = n_3689 ^ n_3119;
assign n_3720 = n_3689 ^ ~n_3521;
assign n_3721 = n_3690 & ~n_3400;
assign n_3722 = n_3691 & n_3399;
assign n_3723 = n_3690 ^ n_3691;
assign n_3724 = n_3692 ^ n_3402;
assign n_3725 = ~n_224 & ~n_3692;
assign n_3726 = ~n_3692 & n_173;
assign n_3727 = ~n_3692 & n_302;
assign n_3728 = ~n_103 & n_3693;
assign n_3729 = ~n_142 & ~n_3693;
assign n_3730 = ~n_231 & ~n_3694;
assign n_3731 = n_3695 ^ n_87;
assign n_3732 = n_3697 ^ n_165;
assign n_3733 = ~n_3670 & ~n_3699;
assign n_3734 = n_3700 ^ n_3692;
assign n_3735 = n_130 & ~n_3700;
assign n_3736 = ~n_157 & ~n_3700;
assign n_3737 = ~n_60 & ~n_3700;
assign n_3738 = n_122 & ~n_3700;
assign n_3739 = n_163 & ~n_3700;
assign n_3740 = n_3511 & ~n_3701;
assign n_3741 = n_3702 ^ ~n_3473;
assign n_3742 = n_3674 ^ n_3702;
assign n_3743 = n_3509 ^ n_3703;
assign n_3744 = ~n_3703 & ~n_3513;
assign n_3745 = ~n_3704 ^ ~n_3594;
assign n_3746 = n_3666 ^ n_3705;
assign n_3747 = ~n_3706 ^ n_87;
assign n_3748 = n_3580 & ~n_3707;
assign n_3749 = n_3708 & ~n_3709;
assign n_3750 = ~n_3710 ^ n_187;
assign n_3751 = n_3711 ^ n_3641;
assign n_3752 = ~n_3714 ^ n_3231;
assign n_3753 = ~n_3577 & ~n_3715;
assign n_3754 = n_3234 ^ n_3717;
assign n_3755 = n_3610 ^ n_3717;
assign n_3756 = ~n_3521 ^ n_3718;
assign n_3757 = ~n_3719 & ~n_3720;
assign n_3758 = n_3664 ^ n_3721;
assign n_3759 = ~n_3723 & ~n_3399;
assign n_3760 = n_3728 ^ n_143;
assign n_3761 = n_3729 ^ n_3730;
assign n_3762 = n_3724 ^ n_3734;
assign n_3763 = n_201 & n_3734;
assign n_3764 = n_122 & n_3734;
assign n_3765 = n_163 & n_3734;
assign n_3766 = n_100 & n_3735;
assign n_3767 = n_144 & ~n_3735;
assign n_3768 = ~n_3629 & n_3736;
assign n_3769 = n_3634 ^ n_3737;
assign n_3770 = n_3636 & n_3738;
assign n_3771 = n_3639 & n_3739;
assign n_3772 = n_3741 & n_3742;
assign n_3773 = ~n_3474 ^ ~n_3743;
assign n_3774 = ~n_3744 ^ ~n_3599;
assign n_3775 = ~n_3745 ^ ~n_3740;
assign n_3776 = n_3748 ^ n_3580;
assign n_3777 = n_3749 ^ n_3616;
assign n_3778 = n_3752 & n_3686;
assign n_3779 = n_3658 ^ n_3752;
assign n_3780 = n_3753 ^ n_3685;
assign n_3781 = ~n_3610 & ~n_3754;
assign n_3782 = n_3757 ^ n_3119;
assign n_3783 = n_3758 ^ n_1930;
assign n_3784 = ~n_3758 & ~n_1930;
assign n_3785 = n_3758 & n_3624;
assign n_3786 = n_3759 & ~n_3624;
assign n_3787 = n_3722 ^ n_3759;
assign n_3788 = n_3627 ^ n_3761;
assign n_3789 = ~n_231 & n_3762;
assign n_3790 = ~n_134 & n_3764;
assign n_3791 = n_3765 ^ n_187;
assign n_3792 = n_3766 ^ n_130;
assign n_3793 = n_3767 ^ n_3626;
assign n_3794 = ~n_3725 ^ ~n_3768;
assign n_3795 = n_3769 ^ n_3595;
assign n_3796 = ~n_3727 ^ ~n_3771;
assign n_3797 = n_3772 ^ n_3674;
assign n_3798 = ~n_187 & n_3773;
assign n_3799 = ~n_3775 ^ n_3656;
assign n_3800 = n_3776 & ~n_3663;
assign n_3801 = n_3778 ^ ~n_3714;
assign n_3802 = n_3585 ^ n_3780;
assign n_3803 = n_3618 ^ n_3780;
assign n_3804 = n_3781 ^ n_3576;
assign n_3805 = n_3782 ^ n_3208;
assign n_3806 = n_3783 & n_260;
assign n_3807 = n_3783 ^ n_74;
assign n_3808 = n_3783 & n_228;
assign n_3809 = n_22 & ~n_3783;
assign n_3810 = n_0 & ~n_3783;
assign n_3811 = n_141 ^ n_3783;
assign n_3812 = n_3783 ^ n_100;
assign n_3813 = ~n_3783 & ~n_183;
assign n_3814 = n_3783 & ~n_106;
assign n_3815 = n_3783 ^ n_112;
assign n_3816 = n_103 & n_3783;
assign n_3817 = n_3783 & n_114;
assign n_3818 = n_3783 ^ n_121;
assign n_3819 = ~n_3783 & n_197;
assign n_3820 = ~n_3783 & n_198;
assign n_3821 = n_163 & ~n_3783;
assign n_3822 = ~n_3783 & n_234;
assign n_3823 = ~n_3783 & n_208;
assign n_3824 = n_3641 ^ n_3783;
assign n_3825 = n_3783 ^ n_3589;
assign n_3826 = n_3783 ^ n_3784;
assign n_3827 = ~n_3722 & ~n_3785;
assign n_3828 = n_3786 ^ n_3758;
assign n_3829 = n_3758 ^ n_3787;
assign n_3830 = n_3787 ^ n_1930;
assign n_3831 = n_3726 ^ n_3790;
assign n_3832 = n_3553 ^ n_3792;
assign n_3833 = ~n_3794 & ~n_3763;
assign n_3834 = n_3795 ^ n_141;
assign n_3835 = ~n_3796 ^ n_187;
assign n_3836 = n_3797 ^ n_3702;
assign n_3837 = ~n_3798 & ~n_3774;
assign n_3838 = ~n_3777 & ~n_3800;
assign n_3839 = n_3801 ^ n_3493;
assign n_3840 = n_3801 ^ n_3682;
assign n_3841 = n_3618 & ~n_3802;
assign n_3842 = n_3712 ^ n_3804;
assign n_3843 = n_3331 ^ n_3804;
assign n_3844 = ~n_187 & ~n_3805;
assign n_3845 = ~n_157 & n_3807;
assign n_3846 = n_3808 ^ n_3783;
assign n_3847 = n_98 & n_3812;
assign n_3848 = n_3814 ^ n_117;
assign n_3849 = n_99 & ~n_3816;
assign n_3850 = n_122 & n_3818;
assign n_3851 = n_3642 ^ n_3821;
assign n_3852 = ~n_184 & ~n_3823;
assign n_3853 = ~n_187 & n_3825;
assign n_3854 = ~n_3825 & n_3643;
assign n_3855 = n_3826 ^ n_1912;
assign n_3856 = ~n_1912 & n_3826;
assign n_3857 = n_3828 ^ n_3827;
assign n_3858 = ~n_3829 & ~n_3625;
assign n_3859 = n_3829 & n_98;
assign n_3860 = n_3829 & ~n_202;
assign n_3861 = n_3829 & ~n_260;
assign n_3862 = n_298 ^ n_3829;
assign n_3863 = n_3731 ^ n_3829;
assign n_3864 = n_74 & n_3829;
assign n_3865 = n_3829 & ~n_225;
assign n_3866 = ~n_19 & n_3829;
assign n_3867 = n_3829 ^ n_14;
assign n_3868 = n_3696 ^ n_3829;
assign n_3869 = n_3829 & ~n_130;
assign n_3870 = ~n_3829 & ~n_231;
assign n_3871 = ~n_3829 & n_122;
assign n_3872 = n_3829 & n_197;
assign n_3873 = n_3829 & n_198;
assign n_3874 = n_3732 ^ n_3829;
assign n_3875 = n_3829 & n_234;
assign n_3876 = n_3829 & n_301;
assign n_3877 = n_3589 ^ n_3829;
assign n_3878 = n_3648 & ~n_3831;
assign n_3879 = n_3789 ^ n_3832;
assign n_3880 = ~n_3747 & n_3833;
assign n_3881 = n_3834 ^ n_3779;
assign n_3882 = ~n_187 ^ ~n_3835;
assign n_3883 = n_3836 ^ n_3674;
assign n_3884 = n_141 ^ n_3837;
assign n_3885 = ~n_141 & n_3837;
assign n_3886 = n_3353 & n_3837;
assign n_3887 = n_3779 ^ n_3838;
assign n_3888 = ~n_3682 & ~n_3839;
assign n_3889 = n_3841 ^ n_3578;
assign n_3890 = n_3712 & ~n_3843;
assign n_3891 = n_614 & n_3846;
assign n_3892 = n_3848 & ~n_3815;
assign n_3893 = ~n_108 & ~n_3849;
assign n_3894 = n_3824 ^ n_3853;
assign n_3895 = n_3853 ^ n_103;
assign n_3896 = n_3854 ^ n_103;
assign n_3897 = ~n_3855 & ~n_115;
assign n_3898 = n_3855 & n_743;
assign n_3899 = n_22 & ~n_3855;
assign n_3900 = x1 & n_3855;
assign n_3901 = ~x0 & n_3855;
assign n_3902 = ~n_3855 & n_117;
assign n_3903 = n_3855 & ~n_129;
assign n_3904 = n_3855 ^ n_103;
assign n_3905 = n_122 ^ n_3855;
assign n_3906 = n_3855 & n_197;
assign n_3907 = n_3855 & n_198;
assign n_3908 = n_163 & n_3855;
assign n_3909 = n_3855 ^ n_165;
assign n_3910 = n_3855 & n_185;
assign n_3911 = ~n_187 & n_3855;
assign n_3912 = ~n_3855 & n_240;
assign n_3913 = n_3855 ^ n_3856;
assign n_3914 = n_3857 & n_1930;
assign n_3915 = n_3857 ^ n_3625;
assign n_3916 = n_3858 ^ n_3758;
assign n_3917 = n_1912 ^ n_3858;
assign n_3918 = n_3760 ^ n_3859;
assign n_3919 = ~n_3861 & n_3862;
assign n_3920 = ~n_157 & ~n_3863;
assign n_3921 = n_95 ^ n_3864;
assign n_3922 = n_3865 ^ n_3631;
assign n_3923 = ~n_34 & ~n_3866;
assign n_3924 = x1 & ~n_3867;
assign n_3925 = n_3868 ^ n_3668;
assign n_3926 = n_3869 ^ n_3635;
assign n_3927 = n_3870 ^ n_100;
assign n_3928 = n_3871 ^ n_152;
assign n_3929 = n_3872 ^ n_3638;
assign n_3930 = n_3873 ^ n_3819;
assign n_3931 = n_163 & n_3874;
assign n_3932 = n_3876 ^ n_3822;
assign n_3933 = ~n_187 & n_3877;
assign n_3934 = n_3726 ^ n_3878;
assign n_3935 = n_3879 ^ n_3793;
assign n_3936 = ~n_3794 ^ n_3880;
assign n_3937 = ~n_3882 ^ n_187;
assign n_3938 = n_3512 & ~n_3883;
assign n_3939 = n_3884 ^ n_3208;
assign n_3940 = n_3208 ^ ~n_3884;
assign n_3941 = n_3884 & n_3476;
assign n_3942 = n_3208 & n_3885;
assign n_3943 = n_3885 ^ n_3884;
assign n_3944 = n_3443 & n_3886;
assign n_3945 = n_3445 & n_3886;
assign n_3946 = ~n_3881 & n_3887;
assign n_3947 = n_3888 ^ ~n_3653;
assign n_3948 = n_3660 ^ n_3889;
assign n_3949 = n_3713 ^ n_3889;
assign n_3950 = n_3890 ^ n_3681;
assign n_3951 = n_202 ^ n_3891;
assign n_3952 = n_3813 ^ n_3892;
assign n_3953 = n_3894 ^ n_3855;
assign n_3954 = n_3855 & ~n_3896;
assign n_3955 = n_3896 ^ n_3855;
assign n_3956 = n_3897 ^ n_87;
assign n_3957 = n_3898 ^ n_613;
assign n_3958 = n_3900 ^ n_3809;
assign n_3959 = n_3903 ^ n_3817;
assign n_3960 = n_3904 ^ n_3816;
assign n_3961 = ~n_3855 & ~n_3905;
assign n_3962 = ~n_3906 ^ ~n_3820;
assign n_3963 = n_163 & n_3909;
assign n_3964 = n_3910 ^ n_164;
assign n_3965 = n_3911 ^ n_187;
assign n_3966 = n_3912 ^ n_164;
assign n_3967 = n_3913 & n_1861;
assign n_3968 = n_3913 ^ n_1861;
assign n_3969 = n_3914 ^ n_3827;
assign n_3970 = n_3915 ^ n_3858;
assign n_3971 = n_3917 & n_2064;
assign n_3972 = n_3918 ^ n_3788;
assign n_3973 = ~n_3746 ^ ~n_3920;
assign n_3974 = ~n_3667 & n_3921;
assign n_3975 = n_116 ^ n_3923;
assign n_3976 = ~x0 & n_3925;
assign n_3977 = n_103 ^ ~n_3926;
assign n_3978 = n_3927 ^ n_3893;
assign n_3979 = ~n_3665 & n_3928;
assign n_3980 = ~n_134 & ~n_3929;
assign n_3981 = n_3930 ^ n_134;
assign n_3982 = n_3733 ^ ~n_3931;
assign n_3983 = n_187 ^ ~n_3932;
assign n_3984 = ~n_3934 ^ ~n_3770;
assign n_3985 = n_3755 ^ n_3935;
assign n_3986 = n_3716 ^ n_3936;
assign n_3987 = ~n_3791 & ~n_3937;
assign n_3988 = n_3674 ^ n_3938;
assign n_3989 = ~n_3782 ^ n_3939;
assign n_3990 = n_3782 & n_3940;
assign n_3991 = n_141 & ~n_3941;
assign n_3992 = n_3254 & n_3942;
assign n_3993 = n_3443 ^ n_3942;
assign n_3994 = ~n_3254 & n_3943;
assign n_3995 = n_187 & ~n_3943;
assign n_3996 = ~n_3530 & n_3945;
assign n_3997 = n_3834 ^ n_3946;
assign n_3998 = n_3947 ^ n_3656;
assign n_3999 = n_3947 ^ n_3799;
assign n_4000 = n_3713 & ~n_3948;
assign n_4001 = n_3496 ^ n_3950;
assign n_4002 = n_134 & ~n_3953;
assign n_4003 = n_3955 ^ n_3954;
assign n_4004 = ~n_157 & n_3956;
assign n_4005 = ~n_3951 & ~n_3957;
assign n_4006 = n_90 & n_3960;
assign n_4007 = n_3961 ^ n_3855;
assign n_4008 = n_134 ^ ~n_3962;
assign n_4009 = ~n_3964 ^ ~n_3852;
assign n_4010 = ~n_184 & ~n_3965;
assign n_4011 = ~n_3967 & n_1860;
assign n_4012 = n_3967 ^ n_1860;
assign n_4013 = n_3968 & ~n_48;
assign n_4014 = n_3968 ^ n_14;
assign n_4015 = n_3968 ^ n_87;
assign n_4016 = n_87 & ~n_3968;
assign n_4017 = ~n_3968 & n_531;
assign n_4018 = n_3968 & ~n_130;
assign n_4019 = ~n_3968 & n_122;
assign n_4020 = n_3968 ^ n_121;
assign n_4021 = ~n_3968 & n_197;
assign n_4022 = ~n_3968 & n_198;
assign n_4023 = n_3968 & n_210;
assign n_4024 = ~n_3968 & n_240;
assign n_4025 = ~n_184 & n_3968;
assign n_4026 = ~n_187 & ~n_3968;
assign n_4027 = n_3968 & n_1860;
assign n_4028 = n_3856 & n_3969;
assign n_4029 = n_3970 ^ n_3625;
assign n_4030 = n_3970 & n_122;
assign n_4031 = ~n_3916 & n_3971;
assign n_4032 = ~n_3973 ^ n_3803;
assign n_4033 = ~n_3922 ^ ~n_3974;
assign n_4034 = n_3868 ^ n_3976;
assign n_4035 = n_3952 ^ n_3978;
assign n_4036 = n_3980 ^ n_134;
assign n_4037 = n_3981 ^ n_3855;
assign n_4038 = ~n_3984 ^ n_3661;
assign n_4039 = ~n_3882 ^ n_3987;
assign n_4040 = ~n_3988 ^ ~n_3597;
assign n_4041 = ~n_187 & ~n_3990;
assign n_4042 = n_141 ^ n_3991;
assign n_4043 = ~n_3944 & ~n_3991;
assign n_4044 = n_3992 ^ n_3994;
assign n_4045 = n_3942 ^ n_3994;
assign n_4046 = ~n_3995 & ~n_3996;
assign n_4047 = n_3997 ^ n_3840;
assign n_4048 = ~n_3799 & ~n_3998;
assign n_4049 = n_4000 ^ n_3683;
assign n_4050 = n_4002 ^ n_3855;
assign n_4051 = ~n_187 & ~n_4003;
assign n_4052 = n_4006 ^ n_3816;
assign n_4053 = n_4011 ^ n_1860;
assign n_4054 = n_22 & ~n_4012;
assign n_4055 = n_0 & ~n_4012;
assign n_4056 = n_4012 ^ x22;
assign n_4057 = n_4012 ^ n_74;
assign n_4058 = ~n_4012 & ~n_225;
assign n_4059 = ~n_4012 & n_531;
assign n_4060 = ~n_4012 & n_98;
assign n_4061 = n_144 ^ n_4012;
assign n_4062 = ~n_4012 & n_122;
assign n_4063 = ~n_4012 & n_197;
assign n_4064 = ~n_4012 & n_198;
assign n_4065 = n_4012 & n_234;
assign n_4066 = ~n_4012 & n_301;
assign n_4067 = x1 & n_4014;
assign n_4068 = n_4016 ^ n_4012;
assign n_4069 = ~n_4019 ^ ~n_4008;
assign n_4070 = n_4024 ^ n_4010;
assign n_4071 = n_4025 ^ n_209;
assign n_4072 = ~n_187 & ~n_4027;
assign n_4073 = n_4027 ^ n_3968;
assign n_4074 = ~n_134 & ~n_4027;
assign n_4075 = ~n_4028 & n_1861;
assign n_4076 = ~n_4029 & ~n_3830;
assign n_4077 = n_1 & n_4029;
assign n_4078 = n_4029 ^ n_3624;
assign n_4079 = n_4029 & ~n_483;
assign n_4080 = n_4029 & n_3845;
assign n_4081 = n_4029 & n_3847;
assign n_4082 = n_4029 & n_3850;
assign n_4083 = ~n_4030 ^ ~n_3669;
assign n_4084 = n_1912 ^ n_4031;
assign n_4085 = ~n_4033 ^ n_87;
assign n_4086 = ~n_87 & ~n_4033;
assign n_4087 = n_4034 ^ n_141;
assign n_4088 = n_4036 ^ n_3929;
assign n_4089 = n_4037 & ~n_4007;
assign n_4090 = n_4039 ^ n_187;
assign n_4091 = ~n_4040 ^ n_3496;
assign n_4092 = ~n_3568 ^ ~n_4042;
assign n_4093 = n_3530 & ~n_4042;
assign n_4094 = n_141 ^ n_4043;
assign n_4095 = n_3352 ^ n_4044;
assign n_4096 = ~n_3352 & n_4045;
assign n_4097 = n_4048 ^ ~n_3775;
assign n_4098 = n_3935 ^ n_4049;
assign n_4099 = n_3985 ^ n_4049;
assign n_4100 = ~n_165 & n_4050;
assign n_4101 = ~n_3954 & n_4051;
assign n_4102 = ~n_98 & ~n_4052;
assign n_4103 = n_1916 & ~n_4053;
assign n_4104 = n_4055 ^ n_70;
assign n_4105 = n_4058 ^ n_4017;
assign n_4106 = n_4062 ^ n_3907;
assign n_4107 = n_4063 ^ n_4022;
assign n_4108 = ~n_74 & ~n_4068;
assign n_4109 = ~n_4069 ^ n_4020;
assign n_4110 = n_3966 ^ n_4071;
assign n_4111 = n_4073 ^ n_4012;
assign n_4112 = n_3967 ^ n_4075;
assign n_4113 = n_4076 ^ n_3855;
assign n_4114 = n_4076 & ~n_199;
assign n_4115 = n_4076 ^ n_3858;
assign n_4116 = ~n_112 & n_4076;
assign n_4117 = n_121 & n_4076;
assign n_4118 = ~n_4076 & n_3908;
assign n_4119 = n_4076 & n_3963;
assign n_4120 = n_4077 ^ n_3811;
assign n_4121 = n_122 & ~n_4078;
assign n_4122 = n_3875 ^ n_4079;
assign n_4123 = ~n_134 & n_4083;
assign n_4124 = ~n_4084 & ~n_1861;
assign n_4125 = n_4028 ^ n_4084;
assign n_4126 = n_4085 ^ n_4086;
assign n_4127 = n_4087 ^ n_3840;
assign n_4128 = n_4088 ^ ~n_4082;
assign n_4129 = n_4089 ^ n_3961;
assign n_4130 = n_4090 ^ ~n_3796;
assign n_4131 = n_4091 ^ n_3950;
assign n_4132 = n_4091 & n_4001;
assign n_4133 = ~n_4092 ^ n_4093;
assign n_4134 = n_3993 ^ n_4096;
assign n_4135 = n_4097 ^ n_3936;
assign n_4136 = n_4097 ^ n_3986;
assign n_4137 = n_3985 & n_4098;
assign n_4138 = n_4009 & ~n_4100;
assign n_4139 = n_3959 ^ n_4102;
assign n_4140 = x1 & n_4103;
assign n_4141 = ~n_75 & n_4103;
assign n_4142 = n_22 & n_4103;
assign n_4143 = n_4103 ^ n_4012;
assign n_4144 = ~n_225 & n_4103;
assign n_4145 = n_531 & n_4103;
assign n_4146 = n_87 & n_4103;
assign n_4147 = n_98 & n_4103;
assign n_4148 = n_4103 ^ n_103;
assign n_4149 = ~n_121 & n_4103;
assign n_4150 = n_197 & n_4103;
assign n_4151 = n_198 & n_4103;
assign n_4152 = n_163 & n_4103;
assign n_4153 = n_234 & n_4103;
assign n_4154 = ~n_187 & ~n_4103;
assign n_4155 = ~n_237 & ~n_4103;
assign n_4156 = n_240 & n_4103;
assign n_4157 = ~n_4103 & n_1745;
assign n_4158 = n_4103 & ~n_1902;
assign n_4159 = n_4103 & ~n_1840;
assign n_4160 = n_134 ^ ~n_4107;
assign n_4161 = n_4012 ^ n_4108;
assign n_4162 = n_4070 ^ n_4110;
assign n_4163 = n_4072 & n_4111;
assign n_4164 = n_4111 & ~n_4074;
assign n_4165 = ~n_4112 & n_1860;
assign n_4166 = n_4113 ^ n_84;
assign n_4167 = n_4113 ^ n_89;
assign n_4168 = n_134 & ~n_4113;
assign n_4169 = n_4114 ^ n_4004;
assign n_4170 = n_4115 ^ n_4029;
assign n_4171 = ~n_157 & ~n_4115;
assign n_4172 = ~n_4115 & n_98;
assign n_4173 = ~n_4115 & n_122;
assign n_4174 = n_4116 ^ n_103;
assign n_4175 = ~n_3932 ^ ~n_4118;
assign n_4176 = n_3924 ^ n_4120;
assign n_4177 = ~n_4121 & ~n_3698;
assign n_4178 = n_3851 ^ n_4122;
assign n_4179 = ~n_4124 & n_4011;
assign n_4180 = n_4075 ^ n_4124;
assign n_4181 = n_3967 ^ n_4124;
assign n_4182 = n_4125 ^ n_3969;
assign n_4183 = n_115 & ~n_4125;
assign n_4184 = n_1 & ~n_4125;
assign n_4185 = ~n_112 & ~n_4125;
assign n_4186 = n_4125 & n_4019;
assign n_4187 = n_122 & ~n_4125;
assign n_4188 = n_207 & ~n_4125;
assign n_4189 = ~n_4126 & ~n_4080;
assign n_4190 = ~n_4127 & n_4047;
assign n_4191 = n_4129 ^ n_3855;
assign n_4192 = n_3750 & ~n_4130;
assign n_4193 = n_4132 ^ ~n_4040;
assign n_4194 = ~n_3982 ^ n_4134;
assign n_4195 = n_3986 & ~n_4135;
assign n_4196 = n_4137 ^ n_4049;
assign n_4197 = ~n_100 & n_4139;
assign n_4198 = n_4140 ^ n_4054;
assign n_4199 = n_4141 ^ n_105;
assign n_4200 = n_4142 ^ n_1821;
assign n_4201 = n_74 & ~n_4143;
assign n_4202 = n_4144 ^ n_4059;
assign n_4203 = n_1824 ^ n_4145;
assign n_4204 = n_4146 ^ n_1745;
assign n_4205 = n_4064 ^ n_4150;
assign n_4206 = n_1833 ^ n_4151;
assign n_4207 = n_4153 ^ n_4066;
assign n_4208 = ~n_263 & ~n_4154;
assign n_4209 = n_1902 ^ n_4154;
assign n_4210 = n_165 & n_4155;
assign n_4211 = n_267 & ~n_4156;
assign n_4212 = ~n_4159 & n_1896;
assign n_4213 = ~n_179 & ~n_4161;
assign n_4214 = n_165 & n_4162;
assign n_4215 = n_134 ^ n_4163;
assign n_4216 = n_4103 ^ n_4164;
assign n_4217 = n_4165 ^ n_4075;
assign n_4218 = ~n_4076 & n_4166;
assign n_4219 = n_4076 & n_4167;
assign n_4220 = n_4168 ^ n_4117;
assign n_4221 = ~n_4113 & n_4169;
assign n_4222 = n_201 & ~n_4170;
assign n_4223 = ~n_4170 & n_98;
assign n_4224 = ~n_4170 & n_173;
assign n_4225 = n_4086 & ~n_4171;
assign n_4226 = ~n_4172 & ~n_3977;
assign n_4227 = n_3980 & ~n_4173;
assign n_4228 = n_4174 ^ n_3855;
assign n_4229 = ~n_187 & n_4175;
assign n_4230 = n_4176 ^ n_4120;
assign n_4231 = ~n_4177 ^ ~n_3979;
assign n_4232 = n_4178 & ~n_4133;
assign n_4233 = n_4178 ^ n_187;
assign n_4234 = n_4178 ^ n_4043;
assign n_4235 = n_4178 ^ n_87;
assign n_4236 = ~n_4178 & ~n_4046;
assign n_4237 = ~n_4179 & n_4103;
assign n_4238 = n_1 & n_4180;
assign n_4239 = n_87 & n_4180;
assign n_4240 = n_4180 & ~n_260;
assign n_4241 = n_3855 ^ n_4180;
assign n_4242 = ~n_4180 & n_130;
assign n_4243 = ~n_4180 & n_122;
assign n_4244 = ~n_4180 & n_152;
assign n_4245 = n_207 & n_4180;
assign n_4246 = n_4182 ^ n_3829;
assign n_4247 = n_163 & ~n_4182;
assign n_4248 = n_4183 ^ n_87;
assign n_4249 = n_4184 ^ n_3968;
assign n_4250 = n_4185 ^ n_103;
assign n_4251 = ~n_4186 ^ ~n_3962;
assign n_4252 = n_4187 & ~n_4109;
assign n_4253 = n_4188 ^ n_3968;
assign n_4254 = n_4087 ^ n_4190;
assign n_4255 = n_4191 ^ n_122;
assign n_4256 = ~n_3796 ^ n_4192;
assign n_4257 = n_4038 ^ n_4193;
assign n_4258 = n_3661 ^ n_4193;
assign n_4259 = n_4195 ^ n_4097;
assign n_4260 = n_3842 ^ n_4196;
assign n_4261 = n_4196 ^ n_3972;
assign n_4262 = n_4102 ^ n_4197;
assign n_4263 = n_4013 ^ n_4199;
assign n_4264 = n_4201 ^ n_4012;
assign n_4265 = n_202 & ~n_4204;
assign n_4266 = n_134 ^ ~n_4205;
assign n_4267 = n_4206 ^ n_134;
assign n_4268 = n_134 & n_4206;
assign n_4269 = n_4207 ^ n_187;
assign n_4270 = n_187 & n_4207;
assign n_4271 = n_4208 ^ n_1836;
assign n_4272 = n_239 ^ n_4210;
assign n_4273 = n_1745 & n_4210;
assign n_4274 = n_1900 ^ n_4211;
assign n_4275 = ~n_4105 ^ ~n_4213;
assign n_4276 = n_4110 ^ n_4214;
assign n_4277 = ~n_187 & n_4216;
assign n_4278 = n_4217 & ~n_1916;
assign n_4279 = n_4217 ^ n_4179;
assign n_4280 = n_4218 ^ n_3810;
assign n_4281 = n_4219 ^ n_3901;
assign n_4282 = n_122 & n_4220;
assign n_4283 = n_4004 ^ n_4221;
assign n_4284 = ~n_4222 & n_4189;
assign n_4285 = ~n_4223 ^ ~n_3926;
assign n_4286 = ~n_4128 ^ ~n_4224;
assign n_4287 = ~n_4226 ^ ~n_4081;
assign n_4288 = n_98 & n_4228;
assign n_4289 = ~n_4229 ^ ~n_4119;
assign n_4290 = ~n_4230 ^ ~n_3632;
assign n_4291 = ~n_4231 & ~n_4123;
assign n_4292 = n_4232 ^ n_4093;
assign n_4293 = n_4233 ^ n_4043;
assign n_4294 = n_3530 & n_4234;
assign n_4295 = n_4235 ^ n_4043;
assign n_4296 = ~n_4237 & n_1745;
assign n_4297 = n_4238 ^ x1;
assign n_4298 = n_4240 ^ n_157;
assign n_4299 = n_431 & n_4241;
assign n_4300 = n_231 & ~n_4241;
assign n_4301 = n_144 & ~n_4242;
assign n_4302 = n_100 & n_4242;
assign n_4303 = ~n_4243 & ~n_151;
assign n_4304 = n_4243 ^ n_122;
assign n_4305 = n_4021 ^ n_4244;
assign n_4306 = n_4245 ^ n_165;
assign n_4307 = ~n_224 & ~n_4246;
assign n_4308 = ~n_4247 & ~n_3983;
assign n_4309 = n_4248 ^ n_3968;
assign n_4310 = n_4249 ^ n_3958;
assign n_4311 = n_4250 ^ n_3968;
assign n_4312 = ~n_134 & n_4251;
assign n_4313 = ~n_4069 ^ n_4252;
assign n_4314 = n_163 & n_4253;
assign n_4315 = n_4254 ^ n_3999;
assign n_4316 = ~n_3930 & ~n_4255;
assign n_4317 = n_4256 ^ n_4095;
assign n_4318 = ~n_4038 & n_4258;
assign n_4319 = n_4259 ^ n_3803;
assign n_4320 = n_4259 ^ n_4032;
assign n_4321 = n_4260 ^ n_3972;
assign n_4322 = n_4260 & ~n_4261;
assign n_4323 = ~n_3902 & ~n_4262;
assign n_4324 = ~n_4264 & ~n_261;
assign n_4325 = n_1825 ^ n_4265;
assign n_4326 = n_4267 ^ n_4268;
assign n_4327 = n_4269 ^ n_4270;
assign n_4328 = n_4272 ^ n_1899;
assign n_4329 = ~n_4273 & ~n_4212;
assign n_4330 = ~n_4023 & ~n_4276;
assign n_4331 = n_4278 ^ n_4237;
assign n_4332 = ~n_4278 & ~n_1745;
assign n_4333 = n_4103 ^ n_4279;
assign n_4334 = n_4181 ^ n_4279;
assign n_4335 = n_74 & n_4279;
assign n_4336 = n_4279 & ~n_4275;
assign n_4337 = ~n_144 & ~n_4279;
assign n_4338 = ~n_142 & n_4279;
assign n_4339 = n_4279 ^ n_3968;
assign n_4340 = ~n_121 & n_4279;
assign n_4341 = ~n_234 & n_4279;
assign n_4342 = n_4280 ^ n_4281;
assign n_4343 = n_4284 ^ ~n_4225;
assign n_4344 = ~n_103 & n_4285;
assign n_4345 = ~n_4286 ^ ~n_4227;
assign n_4346 = n_4035 ^ ~n_4288;
assign n_4347 = ~n_4290 ^ n_4120;
assign n_4348 = n_4292 & ~n_3945;
assign n_4349 = n_4294 ^ n_4178;
assign n_4350 = ~n_212 & n_4295;
assign n_4351 = n_4296 & ~n_1896;
assign n_4352 = n_163 & n_4296;
assign n_4353 = ~n_4296 & n_1986;
assign n_4354 = ~n_4296 & ~n_2107;
assign n_4355 = ~n_4296 & ~n_2109;
assign n_4356 = ~n_4296 & ~n_2113;
assign n_4357 = n_4056 ^ n_4297;
assign n_4358 = ~n_4057 & ~n_4298;
assign n_4359 = n_4300 ^ n_3855;
assign n_4360 = n_4301 ^ n_4018;
assign n_4361 = n_4302 ^ n_4180;
assign n_4362 = n_4106 ^ n_4304;
assign n_4363 = n_4306 ^ n_4012;
assign n_4364 = n_4307 ^ n_3919;
assign n_4365 = ~n_4289 & ~n_4308;
assign n_4366 = ~n_157 & n_4309;
assign n_4367 = ~x0 & ~n_4310;
assign n_4368 = n_98 & n_4311;
assign n_4369 = ~n_4313 & ~n_4312;
assign n_4370 = ~n_4138 ^ ~n_4314;
assign n_4371 = n_3981 ^ n_4316;
assign n_4372 = n_4318 ^ ~n_3984;
assign n_4373 = n_4032 & ~n_4319;
assign n_4374 = n_4322 ^ n_3972;
assign n_4375 = ~n_4202 ^ ~n_4324;
assign n_4376 = n_4203 ^ n_4325;
assign n_4377 = n_4328 ^ n_4274;
assign n_4378 = n_1 & ~n_4331;
assign n_4379 = n_4331 ^ n_4217;
assign n_4380 = n_74 & ~n_4331;
assign n_4381 = ~n_157 & ~n_4331;
assign n_4382 = n_103 & n_4331;
assign n_4383 = ~n_142 & ~n_4331;
assign n_4384 = n_4331 ^ n_4012;
assign n_4385 = ~n_4331 & n_1823;
assign n_4386 = ~n_4331 & n_1897;
assign n_4387 = ~n_4331 & n_1898;
assign n_4388 = n_4332 ^ n_4296;
assign n_4389 = ~n_60 & ~n_4333;
assign n_4390 = n_4334 ^ n_4239;
assign n_4391 = n_4103 ^ ~n_4335;
assign n_4392 = n_4336 ^ n_157;
assign n_4393 = n_4061 ^ n_4337;
assign n_4394 = n_231 & ~n_4339;
assign n_4395 = ~n_301 & ~n_4339;
assign n_4396 = n_4340 ^ n_4103;
assign n_4397 = ~n_4341 & ~n_265;
assign n_4398 = ~n_165 & n_4341;
assign n_4399 = n_3975 ^ n_4342;
assign n_4400 = ~n_4287 & ~n_4344;
assign n_4401 = ~n_4345 ^ n_3884;
assign n_4402 = n_3884 & ~n_4345;
assign n_4403 = n_4345 & n_3989;
assign n_4404 = ~n_4346 ^ n_4257;
assign n_4405 = ~x0 & n_4347;
assign n_4406 = ~n_4236 & ~n_4348;
assign n_4407 = n_4094 & ~n_4349;
assign n_4408 = n_4350 ^ n_4043;
assign n_4409 = ~n_48 & n_4351;
assign n_4410 = ~n_4352 & n_2000;
assign n_4411 = ~n_21 & ~n_4353;
assign n_4412 = n_87 ^ n_4354;
assign n_4413 = n_103 ^ n_4355;
assign n_4414 = n_134 ^ n_4356;
assign n_4415 = n_4067 ^ n_4357;
assign n_4416 = n_4299 ^ n_4358;
assign n_4417 = n_4360 ^ n_4060;
assign n_4418 = n_4361 ^ n_4359;
assign n_4419 = n_4303 ^ n_4362;
assign n_4420 = n_163 & n_4363;
assign n_4421 = n_3860 ^ n_4364;
assign n_4422 = n_3751 ^ n_4365;
assign n_4423 = n_3641 ^ n_4365;
assign n_4424 = n_3711 ^ n_4365;
assign n_4425 = ~n_4366 ^ n_4005;
assign n_4426 = n_4249 ^ n_4367;
assign n_4427 = ~n_4368 ^ n_4323;
assign n_4428 = n_4194 ^ n_4369;
assign n_4429 = n_4134 ^ n_4369;
assign n_4430 = ~n_4370 ^ n_3933;
assign n_4431 = ~n_4370 ^ n_187;
assign n_4432 = ~n_4370 ^ n_3589;
assign n_4433 = n_4371 ^ n_4282;
assign n_4434 = n_3756 ^ n_4372;
assign n_4435 = n_4372 ^ n_4291;
assign n_4436 = n_4373 ^ ~n_3973;
assign n_4437 = n_4131 ^ n_4374;
assign n_4438 = n_87 & n_4375;
assign n_4439 = n_4378 ^ n_1745;
assign n_4440 = n_4379 ^ n_4333;
assign n_4441 = ~n_4379 & ~n_4149;
assign n_4442 = ~n_4380 ^ n_1745;
assign n_4443 = n_4381 ^ ~n_4375;
assign n_4444 = n_4382 ^ n_4148;
assign n_4445 = ~n_231 & n_4384;
assign n_4446 = ~n_4270 ^ ~n_4387;
assign n_4447 = n_1 & ~n_4388;
assign n_4448 = n_4388 & n_1896;
assign n_4449 = n_4388 ^ n_4237;
assign n_4450 = n_1826 ^ n_4388;
assign n_4451 = ~n_224 & ~n_4388;
assign n_4452 = n_144 & n_4388;
assign n_4453 = n_130 & ~n_4388;
assign n_4454 = n_4388 ^ n_4103;
assign n_4455 = n_4388 ^ n_4278;
assign n_4456 = ~n_4388 & n_1998;
assign n_4457 = ~n_4388 & n_2111;
assign n_4458 = n_4389 ^ n_97;
assign n_4459 = n_4390 ^ n_3968;
assign n_4460 = n_87 & ~n_4392;
assign n_4461 = n_130 & ~n_4393;
assign n_4462 = n_4394 ^ n_3968;
assign n_4463 = n_4395 ^ n_3968;
assign n_4464 = n_122 & n_4396;
assign n_4465 = n_4397 ^ n_4065;
assign n_4466 = n_4398 ^ n_4279;
assign n_4467 = n_4136 ^ n_4399;
assign n_4468 = n_4131 ^ n_4400;
assign n_4469 = n_4401 ^ n_3844;
assign n_4470 = ~n_3254 & n_4402;
assign n_4471 = ~n_4403 & n_4041;
assign n_4472 = n_4120 ^ n_4405;
assign n_4473 = n_87 ^ n_4406;
assign n_4474 = n_141 ^ n_4407;
assign n_4475 = n_48 ^ n_4409;
assign n_4476 = n_187 & ~n_4410;
assign n_4477 = n_4157 ^ n_4410;
assign n_4478 = n_4158 & ~n_4410;
assign n_4479 = ~n_4103 & ~n_4410;
assign n_4480 = ~n_4209 & ~n_4410;
assign n_4481 = ~n_4157 & n_4410;
assign n_4482 = n_20 ^ n_4411;
assign n_4483 = ~n_4412 & n_180;
assign n_4484 = ~n_99 & ~n_4413;
assign n_4485 = ~n_123 & ~n_4414;
assign n_4486 = n_4415 ^ n_4357;
assign n_4487 = n_4417 ^ n_4418;
assign n_4488 = n_4419 ^ n_4305;
assign n_4489 = ~n_4420 ^ n_4330;
assign n_4490 = n_3806 ^ n_4421;
assign n_4491 = ~n_4423 & n_4424;
assign n_4492 = n_4321 ^ ~n_4425;
assign n_4493 = n_4426 ^ n_141;
assign n_4494 = ~n_4194 & ~n_4429;
assign n_4495 = n_4431 ^ n_3829;
assign n_4496 = ~n_3877 & ~n_4432;
assign n_4497 = n_4317 ^ n_4433;
assign n_4498 = n_4095 ^ n_4433;
assign n_4499 = n_4434 ^ n_4291;
assign n_4500 = n_4434 & ~n_4435;
assign n_4501 = n_3949 ^ n_4436;
assign n_4502 = n_4436 ^ ~n_4343;
assign n_4503 = ~n_4438 ^ ~n_4385;
assign n_4504 = n_4439 ^ n_4198;
assign n_4505 = ~n_199 & n_4440;
assign n_4506 = n_4440 ^ n_4103;
assign n_4507 = n_153 & n_4440;
assign n_4508 = n_122 & ~n_4441;
assign n_4509 = n_87 & n_4443;
assign n_4510 = n_130 & n_4444;
assign n_4511 = n_4445 ^ n_4331;
assign n_4512 = n_4447 ^ n_1896;
assign n_4513 = n_4448 ^ n_4388;
assign n_4514 = n_122 & ~n_4448;
assign n_4515 = n_4449 ^ ~n_4375;
assign n_4516 = n_122 & ~n_4449;
assign n_4517 = ~n_4449 & n_302;
assign n_4518 = ~n_157 & ~n_4450;
assign n_4519 = n_1830 ^ n_4452;
assign n_4520 = n_100 & n_4453;
assign n_4521 = n_231 & ~n_4454;
assign n_4522 = n_122 & n_4455;
assign n_4523 = n_163 & n_4455;
assign n_4524 = n_4456 ^ n_4448;
assign n_4525 = ~n_4268 ^ ~n_4457;
assign n_4526 = n_4458 ^ n_4104;
assign n_4527 = ~n_260 & ~n_4459;
assign n_4528 = n_157 ^ n_4460;
assign n_4529 = n_4061 ^ n_4461;
assign n_4530 = n_4338 ^ n_4462;
assign n_4531 = ~n_4160 & ~n_4464;
assign n_4532 = n_4152 ^ n_4465;
assign n_4533 = n_4466 ^ n_4463;
assign n_4534 = n_4468 ^ n_4374;
assign n_4535 = n_4468 & ~n_4437;
assign n_4536 = ~n_4470 & ~n_4471;
assign n_4537 = n_3999 ^ n_4472;
assign n_4538 = n_4293 & n_4474;
assign n_4539 = n_4475 ^ n_56;
assign n_4540 = n_4476 ^ n_187;
assign n_4541 = ~n_4476 & n_4329;
assign n_4542 = n_4480 ^ n_4410;
assign n_4543 = n_2116 & ~n_4483;
assign n_4544 = n_2246 & ~n_4484;
assign n_4545 = n_2114 & ~n_4485;
assign n_4546 = ~n_4486 ^ ~n_3899;
assign n_4547 = n_4469 ^ n_4487;
assign n_4548 = n_4473 ^ n_4488;
assign n_4549 = n_3895 ^ ~n_4489;
assign n_4550 = ~n_4283 & n_4490;
assign n_4551 = n_4491 ^ n_3641;
assign n_4552 = ~n_4493 & n_4320;
assign n_4553 = n_4320 ^ n_4493;
assign n_4554 = n_4494 ^ n_4369;
assign n_4555 = ~n_4495 & n_4496;
assign n_4556 = n_4317 & n_4498;
assign n_4557 = ~n_4427 ^ n_4499;
assign n_4558 = n_4500 ^ n_4291;
assign n_4559 = n_4501 ^ ~n_4343;
assign n_4560 = ~n_4501 & n_4502;
assign n_4561 = ~x0 & ~n_4504;
assign n_4562 = n_87 & ~n_4506;
assign n_4563 = ~n_4107 ^ ~n_4508;
assign n_4564 = ~n_4375 ^ n_4509;
assign n_4565 = n_4148 ^ n_4510;
assign n_4566 = n_4383 ^ n_4511;
assign n_4567 = n_4512 ^ n_4200;
assign n_4568 = n_4513 ^ n_4332;
assign n_4569 = n_173 & n_4513;
assign n_4570 = n_4456 ^ n_4513;
assign n_4571 = ~n_4514 & ~n_4326;
assign n_4572 = n_157 & ~n_4515;
assign n_4573 = ~n_4516 ^ ~n_4205;
assign n_4574 = ~n_4517 ^ ~n_4446;
assign n_4575 = n_4518 ^ n_1826;
assign n_4576 = n_130 & n_4519;
assign n_4577 = n_4388 ^ n_4520;
assign n_4578 = n_4521 ^ n_4103;
assign n_4579 = ~n_4522 & ~n_4266;
assign n_4580 = ~n_4523 & ~n_4327;
assign n_4581 = n_4524 & ~n_4271;
assign n_4582 = n_4263 ^ n_4526;
assign n_4583 = n_4015 ^ n_4527;
assign n_4584 = ~n_4391 & ~n_4528;
assign n_4585 = n_4147 ^ n_4529;
assign n_4586 = ~n_4507 ^ ~n_4531;
assign n_4587 = n_4532 ^ n_4533;
assign n_4588 = n_4535 ^ n_4400;
assign n_4589 = n_4497 ^ n_4536;
assign n_4590 = ~n_4537 & ~n_4315;
assign n_4591 = n_4408 ^ n_4538;
assign n_4592 = n_4482 ^ n_4539;
assign n_4593 = n_4484 ^ n_4544;
assign n_4594 = ~n_4546 ^ n_4357;
assign n_4595 = n_4099 ^ n_4550;
assign n_4596 = n_4551 ^ n_4430;
assign n_4597 = ~n_4552 & ~n_1981;
assign n_4598 = n_4552 ^ n_4553;
assign n_4599 = ~n_4553 & n_1904;
assign n_4600 = n_4473 ^ n_4554;
assign n_4601 = n_4431 ^ n_4555;
assign n_4602 = n_4556 ^ n_4433;
assign n_4603 = n_4469 ^ n_4558;
assign n_4604 = n_4560 ^ ~n_4343;
assign n_4605 = n_4439 ^ n_4561;
assign n_4606 = ~n_177 & ~n_4562;
assign n_4607 = ~n_134 & n_4563;
assign n_4608 = ~n_4442 & n_4564;
assign n_4609 = n_4565 ^ n_1829;
assign n_4610 = ~x0 & ~n_4567;
assign n_4611 = n_1 & ~n_4568;
assign n_4612 = ~n_4568 & ~n_2177;
assign n_4613 = n_98 & n_4568;
assign n_4614 = n_134 & ~n_4568;
assign n_4615 = n_136 & n_4568;
assign n_4616 = n_207 & n_4568;
assign n_4617 = ~n_4569 ^ ~n_4525;
assign n_4618 = n_302 & n_4570;
assign n_4619 = n_4572 ^ n_4449;
assign n_4620 = ~n_134 & n_4573;
assign n_4621 = ~n_74 & n_4575;
assign n_4622 = n_1830 ^ n_4576;
assign n_4623 = n_4577 ^ n_4578;
assign n_4624 = ~n_4579 ^ ~n_4386;
assign n_4625 = ~n_4574 ^ ~n_4580;
assign n_4626 = n_4377 & ~n_4581;
assign n_4627 = n_4583 ^ n_201;
assign n_4628 = n_4585 ^ n_4530;
assign n_4629 = n_4101 ^ n_4587;
assign n_4630 = ~n_4587 & n_3954;
assign n_4631 = n_4587 & ~n_4051;
assign n_4632 = n_4404 ^ n_4588;
assign n_4633 = ~n_4346 ^ n_4588;
assign n_4634 = n_4472 ^ n_4590;
assign n_4635 = n_4422 ^ n_4591;
assign n_4636 = n_4593 ^ n_4484;
assign n_4637 = ~x0 & ~n_4594;
assign n_4638 = n_4600 ^ n_4488;
assign n_4639 = ~n_4600 & n_4548;
assign n_4640 = n_3895 ^ n_4601;
assign n_4641 = n_4428 ^ n_4602;
assign n_4642 = n_4603 ^ n_4487;
assign n_4643 = n_4603 & n_4547;
assign n_4644 = n_4604 ^ n_4550;
assign n_4645 = n_4595 ^ n_4604;
assign n_4646 = n_4605 ^ n_141;
assign n_4647 = ~n_4275 ^ n_4606;
assign n_4648 = ~n_4586 & ~n_4607;
assign n_4649 = ~n_4503 & ~n_4608;
assign n_4650 = n_4609 ^ n_4566;
assign n_4651 = n_4512 ^ n_4610;
assign n_4652 = n_4611 ^ n_16;
assign n_4653 = n_4612 ^ n_176;
assign n_4654 = ~n_2245 & n_4613;
assign n_4655 = ~n_149 & ~n_4614;
assign n_4656 = n_163 & ~n_4616;
assign n_4657 = ~n_4617 ^ ~n_4571;
assign n_4658 = n_178 & ~n_4619;
assign n_4659 = n_1826 ^ n_4621;
assign n_4660 = n_1990 ^ n_4622;
assign n_4661 = ~n_4624 & ~n_4620;
assign n_4662 = ~n_4625 ^ n_4545;
assign n_4663 = ~n_4625 & ~n_4545;
assign n_4664 = ~n_4618 ^ n_4626;
assign n_4665 = n_4627 ^ n_4416;
assign n_4666 = n_4589 ^ n_4628;
assign n_4667 = n_4628 ^ n_4536;
assign n_4668 = ~n_187 & n_4630;
assign n_4669 = n_4026 & ~n_4630;
assign n_4670 = n_4631 ^ n_4026;
assign n_4671 = ~n_4404 & n_4633;
assign n_4672 = n_4399 ^ n_4634;
assign n_4673 = n_4357 ^ n_4637;
assign n_4674 = n_4639 ^ n_4554;
assign n_4675 = n_4640 ^ ~n_4489;
assign n_4676 = n_4640 & ~n_4549;
assign n_4677 = n_4643 ^ n_4487;
assign n_4678 = n_4595 & n_4644;
assign n_4679 = n_4582 ^ n_4645;
assign n_4680 = n_4505 ^ n_4647;
assign n_4681 = n_4635 ^ n_4648;
assign n_4682 = n_4591 ^ n_4648;
assign n_4683 = n_4641 ^ n_4650;
assign n_4684 = n_4428 ^ n_4650;
assign n_4685 = n_4651 ^ n_141;
assign n_4686 = n_1822 ^ n_4652;
assign n_4687 = ~n_4653 & ~n_2244;
assign n_4688 = n_2179 ^ n_4654;
assign n_4689 = n_2112 ^ n_4655;
assign n_4690 = ~n_2295 ^ ~n_4656;
assign n_4691 = n_4649 & ~n_4658;
assign n_4692 = n_1987 ^ n_4659;
assign n_4693 = n_4660 ^ n_4623;
assign n_4694 = n_4551 ^ n_4661;
assign n_4695 = n_4663 ^ n_4662;
assign n_4696 = ~n_4664 ^ n_4215;
assign n_4697 = n_4534 ^ n_4665;
assign n_4698 = ~n_4589 & ~n_4667;
assign n_4699 = ~n_4631 & ~n_4669;
assign n_4700 = n_4668 ^ n_4670;
assign n_4701 = n_4671 ^ n_4588;
assign n_4702 = n_4672 & ~n_4467;
assign n_4703 = n_4559 ^ n_4673;
assign n_4704 = n_4676 ^ n_4601;
assign n_4705 = n_4666 ^ n_4677;
assign n_4706 = n_4678 ^ n_4604;
assign n_4707 = ~n_4680 & ~n_4584;
assign n_4708 = n_4635 & n_4682;
assign n_4709 = n_4641 & n_4684;
assign n_4710 = n_4686 ^ n_4652;
assign n_4711 = ~n_2176 & ~n_4687;
assign n_4712 = n_4688 ^ n_4674;
assign n_4713 = ~n_4674 & n_4688;
assign n_4714 = n_4689 ^ n_4615;
assign n_4715 = ~n_4690 ^ n_4277;
assign n_4716 = n_187 & n_4690;
assign n_4717 = ~n_4690 ^ n_4103;
assign n_4718 = ~n_4690 ^ n_187;
assign n_4719 = ~n_4690 & n_4164;
assign n_4720 = n_4592 ^ n_4691;
assign n_4721 = n_4692 ^ n_4451;
assign n_4722 = n_4638 ^ n_4693;
assign n_4723 = n_4694 ^ n_4430;
assign n_4724 = n_4694 & ~n_4596;
assign n_4725 = n_4698 ^ n_4628;
assign n_4726 = n_4696 ^ n_4699;
assign n_4727 = ~n_4664 ^ n_4699;
assign n_4728 = n_4557 ^ n_4701;
assign n_4729 = n_4499 ^ n_4701;
assign n_4730 = n_4702 ^ n_4634;
assign n_4731 = ~n_4703 & ~n_4597;
assign n_4732 = n_4629 ^ n_4704;
assign n_4733 = n_4321 ^ n_4706;
assign n_4734 = n_4708 ^ n_4648;
assign n_4735 = n_4709 ^ n_4650;
assign n_4736 = ~n_2104 ^ ~n_4710;
assign n_4737 = n_4705 ^ n_4711;
assign n_4738 = n_4666 ^ n_4711;
assign n_4739 = n_4713 ^ n_4712;
assign n_4740 = n_4629 ^ n_4714;
assign n_4741 = n_4716 ^ n_187;
assign n_4742 = n_4216 & n_4717;
assign n_4743 = n_4716 ^ n_4718;
assign n_4744 = n_1840 ^ ~n_4719;
assign n_4745 = n_4376 ^ n_4721;
assign n_4746 = n_4724 ^ n_4661;
assign n_4747 = n_4683 ^ n_4725;
assign n_4748 = ~n_4725 & ~n_4683;
assign n_4749 = n_4726 ^ n_4695;
assign n_4750 = ~n_4696 & ~n_4727;
assign n_4751 = n_4728 ^ n_4691;
assign n_4752 = n_4557 & n_4729;
assign n_4753 = ~n_4552 & n_4730;
assign n_4754 = ~n_4730 & n_1904;
assign n_4755 = n_4732 ^ n_4714;
assign n_4756 = n_4733 ^ ~n_4425;
assign n_4757 = n_4733 & ~n_4492;
assign n_4758 = n_4734 ^ n_4636;
assign n_4759 = n_4723 ^ n_4734;
assign n_4760 = n_4638 ^ n_4735;
assign n_4761 = ~n_4736 ^ n_4652;
assign n_4762 = ~n_4705 & ~n_4738;
assign n_4763 = ~n_4732 & n_4740;
assign n_4764 = n_4741 ^ n_4540;
assign n_4765 = n_4742 ^ n_4103;
assign n_4766 = n_4479 & ~n_4744;
assign n_4767 = n_4675 ^ n_4746;
assign n_4768 = ~n_4746 & ~n_4675;
assign n_4769 = n_4748 ^ n_4747;
assign n_4770 = n_4750 ^ n_4699;
assign n_4771 = n_4751 ^ n_4592;
assign n_4772 = n_4751 & ~n_4720;
assign n_4773 = n_4752 ^ ~n_4427;
assign n_4774 = ~n_4598 & ~n_4753;
assign n_4775 = ~n_1904 & n_4753;
assign n_4776 = ~n_1981 ^ n_4754;
assign n_4777 = ~n_4754 & ~n_1981;
assign n_4778 = n_4598 & ~n_4754;
assign n_4779 = n_4646 ^ n_4756;
assign n_4780 = n_4757 ^ n_4706;
assign n_4781 = n_4723 ^ n_4758;
assign n_4782 = n_4758 & n_4759;
assign n_4783 = n_4760 ^ n_4693;
assign n_4784 = ~n_4760 & ~n_4722;
assign n_4785 = ~x0 & n_4761;
assign n_4786 = n_4762 ^ n_4711;
assign n_4787 = n_4763 ^ n_4704;
assign n_4788 = ~n_187 & ~n_4765;
assign n_4789 = n_4768 ^ n_4767;
assign n_4790 = ~n_4768 & ~n_4755;
assign n_4791 = n_4715 ^ n_4770;
assign n_4792 = n_4772 ^ n_4592;
assign n_4793 = n_4642 & ~n_4773;
assign n_4794 = n_4773 ^ n_4642;
assign n_4795 = n_4774 ^ n_4559;
assign n_4796 = n_4776 ^ n_4777;
assign n_4797 = n_4777 & ~n_4599;
assign n_4798 = ~n_4778 ^ n_4731;
assign n_4799 = n_4697 ^ n_4780;
assign n_4800 = n_4665 ^ n_4780;
assign n_4801 = ~n_4781 & ~n_4713;
assign n_4802 = n_4782 ^ n_4723;
assign n_4803 = n_4783 ^ n_4769;
assign n_4804 = n_4784 ^ n_4735;
assign n_4805 = n_4652 ^ n_4785;
assign n_4806 = n_4786 ^ n_4543;
assign n_4807 = ~n_4786 & n_4543;
assign n_4808 = n_4700 ^ n_4787;
assign n_4809 = ~n_4787 & n_4700;
assign n_4810 = n_4743 ^ n_4788;
assign n_4811 = ~n_4792 & ~n_4745;
assign n_4812 = n_4745 ^ n_4792;
assign n_4813 = n_4793 ^ n_4794;
assign n_4814 = n_4703 & ~n_4795;
assign n_4815 = n_4796 ^ n_4730;
assign n_4816 = ~n_4798 & ~n_4775;
assign n_4817 = n_4685 ^ n_4799;
assign n_4818 = ~n_4697 & ~n_4800;
assign n_4819 = ~n_4657 ^ n_4802;
assign n_4820 = ~n_4802 & ~n_4657;
assign n_4821 = n_4681 ^ n_4804;
assign n_4822 = n_4804 & ~n_4681;
assign n_4823 = n_4805 ^ n_4707;
assign n_4824 = ~n_4805 & ~n_4707;
assign n_4825 = n_4806 ^ n_4747;
assign n_4826 = n_4807 ^ n_4806;
assign n_4827 = ~n_4807 & n_4783;
assign n_4828 = ~n_4808 & n_4726;
assign n_4829 = ~n_4809 & ~n_4726;
assign n_4830 = n_4726 ^ n_4809;
assign n_4831 = n_4809 ^ n_4808;
assign n_4832 = n_4810 ^ ~n_4690;
assign n_4833 = n_4793 ^ n_4811;
assign n_4834 = ~n_4811 ^ n_4737;
assign n_4835 = n_4811 ^ n_4812;
assign n_4836 = ~n_4813 & n_4737;
assign n_4837 = n_4673 ^ n_4814;
assign n_4838 = ~n_4553 & ~n_4815;
assign n_4839 = n_4818 ^ n_4780;
assign n_4840 = n_4819 ^ n_4767;
assign n_4841 = n_4820 ^ n_4819;
assign n_4842 = ~n_4820 ^ ~n_4755;
assign n_4843 = n_4821 ^ n_4712;
assign n_4844 = n_4713 ^ n_4822;
assign n_4845 = n_4822 & ~n_4713;
assign n_4846 = n_4822 ^ n_4821;
assign n_4847 = n_4824 ^ n_4823;
assign n_4848 = n_4826 & n_4769;
assign n_4849 = ~n_4748 & ~n_4827;
assign n_4850 = n_4828 ^ n_4663;
assign n_4851 = n_4695 & n_4829;
assign n_4852 = n_4829 ^ n_4809;
assign n_4853 = n_4830 ^ n_4829;
assign n_4854 = n_4830 & ~n_4749;
assign n_4855 = ~n_4158 & n_4832;
assign n_4856 = ~n_4832 & n_4542;
assign n_4857 = n_4832 & ~n_4481;
assign n_4858 = ~n_4793 & n_4834;
assign n_4859 = n_4813 ^ n_4835;
assign n_4860 = n_4582 ^ n_4837;
assign n_4861 = n_4679 ^ n_4837;
assign n_4862 = n_4838 ^ n_4796;
assign n_4863 = n_4632 ^ n_4839;
assign n_4864 = ~n_4839 & n_4632;
assign n_4865 = ~n_4768 & n_4841;
assign n_4866 = n_4789 & n_4842;
assign n_4867 = n_4844 ^ n_4845;
assign n_4868 = ~n_4845 ^ ~n_4801;
assign n_4869 = ~n_4712 & n_4846;
assign n_4870 = ~n_4846 & n_4739;
assign n_4871 = ~n_4781 & ~n_4846;
assign n_4872 = ~n_4783 ^ ~n_4848;
assign n_4873 = n_4850 ^ n_4662;
assign n_4874 = n_4851 ^ n_4829;
assign n_4875 = ~n_4695 & ~n_4852;
assign n_4876 = n_4828 ^ n_4853;
assign n_4877 = n_4854 ^ n_4809;
assign n_4878 = ~n_4855 & ~n_4157;
assign n_4879 = n_4855 ^ n_4832;
assign n_4880 = n_4856 ^ n_4857;
assign n_4881 = n_4857 ^ n_4480;
assign n_4882 = n_4833 ^ n_4859;
assign n_4883 = ~n_4835 & ~n_4859;
assign n_4884 = n_4679 & n_4860;
assign n_4885 = n_4861 ^ n_2072;
assign n_4886 = ~n_4598 & n_4862;
assign n_4887 = n_4823 ^ n_4863;
assign n_4888 = n_4864 ^ n_4863;
assign n_4889 = n_4755 ^ ~n_4865;
assign n_4890 = n_4821 & n_4867;
assign n_4891 = n_4739 & n_4868;
assign n_4892 = n_4870 ^ n_4781;
assign n_4893 = ~n_4870 ^ ~n_4871;
assign n_4894 = ~n_4867 & n_4871;
assign n_4895 = ~n_4828 & n_4873;
assign n_4896 = n_4875 ^ n_4809;
assign n_4897 = n_4874 ^ n_4876;
assign n_4898 = n_4876 ^ n_4663;
assign n_4899 = ~n_4663 & ~n_4876;
assign n_4900 = ~n_4477 & ~n_4878;
assign n_4901 = n_4879 ^ n_4766;
assign n_4902 = ~n_4737 ^ ~n_4883;
assign n_4903 = n_4884 ^ n_4837;
assign n_4904 = n_4552 ^ n_4886;
assign n_4905 = ~n_4888 & ~n_4847;
assign n_4906 = ~n_4771 & ~n_4888;
assign n_4907 = n_4869 ^ n_4892;
assign n_4908 = ~n_4868 ^ ~n_4893;
assign n_4909 = ~n_4891 & ~n_4894;
assign n_4910 = n_4895 ^ n_4850;
assign n_4911 = n_4898 ^ n_4899;
assign n_4912 = ~n_4899 & ~n_4877;
assign n_4913 = ~n_4764 & ~n_4900;
assign n_4914 = ~n_4901 & n_4880;
assign n_4915 = n_4779 ^ n_4903;
assign n_4916 = n_4646 ^ n_4903;
assign n_4917 = n_4703 & ~n_4904;
assign n_4918 = ~n_4829 & n_4911;
assign n_4919 = n_4478 ^ n_4913;
assign n_4920 = n_4915 ^ n_1946;
assign n_4921 = n_4915 & n_1946;
assign n_4922 = n_4779 & ~n_4916;
assign n_4923 = ~n_4917 & ~n_4816;
assign n_4924 = n_4919 ^ n_4879;
assign n_4925 = n_4921 ^ n_4920;
assign n_4926 = n_4922 ^ n_4903;
assign n_4927 = ~n_4923 & ~n_4797;
assign n_4928 = n_4924 ^ n_4914;
assign n_4929 = n_4817 ^ n_4926;
assign n_4930 = n_4685 ^ n_4926;
assign n_4931 = n_2072 ^ n_4927;
assign n_4932 = n_4929 ^ ~n_2175;
assign n_4933 = n_4817 & ~n_4930;
assign n_4934 = ~n_4931 & ~n_4885;
assign n_4935 = ~n_4920 & ~n_4932;
assign n_4936 = n_4933 ^ n_4926;
assign n_4937 = n_4934 ^ n_4885;
assign n_4938 = n_4934 ^ n_4927;
assign n_4939 = n_4935 ^ n_4925;
assign n_4940 = n_4887 ^ n_4936;
assign n_4941 = n_4805 ^ n_4936;
assign n_4942 = n_4936 & n_4824;
assign n_4943 = ~n_4936 & n_4905;
assign n_4944 = n_4920 ^ n_4937;
assign n_4945 = ~n_4861 & ~n_4937;
assign n_4946 = ~n_4921 & n_4938;
assign n_4947 = n_4940 ^ ~n_1801;
assign n_4948 = ~n_4823 & ~n_4941;
assign n_4949 = ~n_4771 ^ ~n_4942;
assign n_4950 = ~n_4864 & ~n_4943;
assign y0 = n_4944;
assign n_4951 = n_4945 ^ n_4937;
assign n_4952 = n_4945 ^ n_18;
assign n_4953 = n_4945 ^ n_4920;
assign n_4954 = ~n_4945 & n_4946;
assign n_4955 = n_4946 ^ n_4935;
assign n_4956 = n_4948 ^ n_4936;
assign n_4957 = n_4949 & n_4950;
assign n_4958 = n_4920 & n_4951;
assign n_4959 = n_18 & ~n_4951;
assign n_4960 = ~n_4951 & ~n_4939;
assign n_4961 = ~n_4952 & ~n_4953;
assign n_4962 = n_4932 & n_4954;
assign n_4963 = n_4945 & ~n_4955;
assign n_4964 = n_4956 & n_4888;
assign n_4965 = n_4942 ^ n_4956;
assign n_4966 = n_4956 & ~n_4906;
assign n_4967 = n_4958 ^ n_4920;
assign n_4968 = n_4958 & ~n_4938;
assign n_4969 = n_4925 ^ n_4961;
assign n_4970 = n_4925 & n_4962;
assign n_4971 = n_4864 & ~n_4965;
assign n_4972 = ~n_4957 & ~n_4966;
assign n_4973 = n_4967 ^ n_4959;
assign n_4974 = n_4932 & n_4968;
assign n_4975 = n_4968 ^ n_4921;
assign n_4976 = n_4960 ^ n_4970;
assign n_4977 = n_4971 ^ n_4942;
assign n_4978 = n_4882 ^ n_4972;
assign n_4979 = n_4745 ^ n_4972;
assign n_4980 = n_4792 ^ n_4972;
assign n_4981 = n_4902 & n_4972;
assign n_4982 = n_4932 ^ n_4973;
assign n_4983 = n_4974 ^ n_4963;
assign n_4984 = n_4975 ^ n_4967;
assign n_4985 = n_18 & n_4976;
assign n_4986 = ~n_4977 & ~n_4943;
assign n_4987 = n_4978 ^ ~n_1855;
assign n_4988 = ~n_1855 & ~n_4978;
assign n_4989 = n_4979 ^ n_4792;
assign n_4990 = n_4979 & n_4980;
assign n_4991 = n_4858 & ~n_4981;
assign n_4992 = n_4982 ^ n_4969;
assign n_4993 = ~n_18 & ~n_4983;
assign n_4994 = n_4984 ^ ~n_2175;
assign n_4995 = ~n_4964 & n_4986;
assign n_4996 = n_4987 ^ n_4988;
assign n_4997 = ~n_4882 & n_4989;
assign n_4998 = n_4990 ^ n_4972;
assign y1 = n_4992;
assign n_4999 = n_4985 ^ n_4993;
assign n_5000 = n_4932 & ~n_4994;
assign n_5001 = n_4771 ^ n_4995;
assign n_5002 = n_4997 ^ n_4833;
assign n_5003 = ~n_4836 & ~n_4998;
assign n_5004 = n_5000 ^ n_4929;
assign n_5005 = n_5001 ^ ~n_1984;
assign n_5006 = n_1984 & n_5001;
assign n_5007 = n_4737 ^ n_5002;
assign n_5008 = ~n_4991 & ~n_5003;
assign n_5009 = n_5004 ^ n_4947;
assign n_5010 = n_5004 ^ n_4940;
assign n_5011 = n_5006 ^ n_5005;
assign n_5012 = n_4976 & ~n_5006;
assign n_5013 = n_5007 ^ n_1857;
assign n_5014 = n_4825 ^ n_5008;
assign n_5015 = n_4748 ^ n_5008;
assign n_5016 = n_4786 ^ n_5008;
assign n_5017 = n_4999 ^ n_5009;
assign n_5018 = ~n_5009 & ~n_5005;
assign n_5019 = ~n_4947 & n_5010;
assign n_5020 = n_5014 ^ n_2071;
assign n_5021 = n_5015 ^ n_4747;
assign n_5022 = n_5015 & n_4872;
assign n_5023 = n_4806 & n_5016;
assign y2 = n_5017;
assign n_5024 = n_5019 ^ n_5004;
assign n_5025 = n_5021 ^ n_4748;
assign n_5026 = ~n_5022 & n_4849;
assign n_5027 = n_5023 ^ n_5008;
assign n_5028 = n_5009 & n_5024;
assign n_5029 = n_5024 ^ n_18;
assign n_5030 = ~n_18 & n_5024;
assign n_5031 = ~n_5024 & ~n_5011;
assign n_5032 = n_4825 & n_5025;
assign n_5033 = n_4803 & ~n_5027;
assign n_5034 = n_5028 ^ n_5024;
assign n_5035 = n_4983 & ~n_5028;
assign n_5036 = n_4976 & n_5028;
assign n_5037 = n_5029 ^ n_5030;
assign n_5038 = ~n_5006 & ~n_5031;
assign n_5039 = n_5032 ^ n_5015;
assign n_5040 = ~n_5033 & ~n_5026;
assign n_5041 = n_5034 ^ n_5009;
assign n_5042 = n_5030 & ~n_5035;
assign n_5043 = n_5005 & n_5036;
assign n_5044 = n_5037 ^ n_5028;
assign n_5045 = n_5038 ^ n_4988;
assign n_5046 = n_4988 & n_5038;
assign n_5047 = n_5013 ^ n_5038;
assign n_5048 = n_4826 ^ n_5039;
assign n_5049 = n_4843 ^ n_5040;
assign n_5050 = n_4712 ^ n_5040;
assign n_5051 = n_4908 & n_5040;
assign n_5052 = ~n_4993 & ~n_5041;
assign n_5053 = n_5018 ^ n_5041;
assign n_5054 = n_5041 & n_5031;
assign n_5055 = ~n_4976 & n_5044;
assign n_5056 = n_5045 ^ n_5046;
assign n_5057 = ~n_4996 ^ n_5047;
assign n_5058 = n_4783 ^ n_5048;
assign n_5059 = n_5049 ^ n_1982;
assign n_5060 = n_1982 & n_5049;
assign n_5061 = n_4843 & n_5050;
assign n_5062 = ~n_5051 & n_4909;
assign n_5063 = n_4983 & ~n_5053;
assign n_5064 = n_5054 & n_5012;
assign n_5065 = n_5055 ^ n_5028;
assign n_5066 = n_4996 ^ n_5056;
assign n_5067 = n_5056 & ~n_4996;
assign n_5068 = ~n_5056 ^ ~n_5013;
assign n_5069 = ~n_5057 ^ n_5038;
assign n_5070 = n_5058 ^ n_2020;
assign n_5071 = n_5060 ^ n_5059;
assign n_5072 = n_5061 ^ n_4890;
assign n_5073 = n_4840 ^ n_5062;
assign n_5074 = n_4819 ^ n_5062;
assign n_5075 = n_4802 ^ n_5062;
assign n_5076 = ~n_4657 ^ n_5062;
assign n_5077 = n_4889 & ~n_5062;
assign n_5078 = ~n_18 & ~n_5063;
assign n_5079 = ~n_5046 & n_5063;
assign n_5080 = n_5043 ^ n_5064;
assign n_5081 = ~n_5052 & ~n_5065;
assign n_5082 = n_5066 ^ n_5046;
assign n_5083 = n_5067 ^ n_5066;
assign n_5084 = n_5007 ^ n_5067;
assign n_5085 = n_5072 ^ n_4907;
assign n_5086 = n_5073 ^ n_1887;
assign n_5087 = ~n_4840 & ~n_5074;
assign n_5088 = ~n_5075 & n_5076;
assign n_5089 = n_4866 & ~n_5077;
assign n_5090 = n_5068 & n_5079;
assign n_5091 = n_18 & ~n_5080;
assign n_5092 = n_5081 & ~n_5042;
assign n_5093 = ~n_5082 & n_5013;
assign n_5094 = n_5013 & ~n_5084;
assign n_5095 = n_1951 ^ n_5085;
assign n_5096 = n_4768 ^ n_5087;
assign n_5097 = n_5088 ^ n_5062;
assign n_5098 = ~n_5069 & n_5090;
assign n_5099 = n_5091 ^ n_18;
assign n_5100 = n_5067 ^ n_5091;
assign n_5101 = n_5005 ^ n_5092;
assign n_5102 = n_5093 ^ n_5066;
assign n_5103 = n_5094 ^ n_5067;
assign n_5104 = n_5095 ^ n_5060;
assign n_5105 = ~n_5071 & n_5095;
assign n_5106 = n_4841 ^ n_5096;
assign n_5107 = ~n_4790 & n_5097;
assign n_5108 = n_5078 ^ n_5099;
assign n_5109 = n_5082 & n_5100;
assign y3 = ~n_5101;
assign n_5110 = n_5080 & ~n_5102;
assign n_5111 = n_5020 ^ n_5103;
assign n_5112 = n_5014 ^ n_5103;
assign n_5113 = n_4755 ^ n_5106;
assign n_5114 = ~n_5089 & ~n_5107;
assign n_5115 = n_5108 ^ n_5082;
assign n_5116 = n_5083 ^ n_5109;
assign n_5117 = n_18 & ~n_5110;
assign n_5118 = n_5111 & n_5098;
assign n_5119 = ~n_5111 & n_5110;
assign n_5120 = n_5020 & ~n_5112;
assign n_5121 = n_2151 ^ n_5113;
assign n_5122 = n_4662 ^ n_5114;
assign n_5123 = n_4808 ^ n_5114;
assign n_5124 = ~n_4831 & ~n_5114;
assign n_5125 = n_4918 & ~n_5114;
assign y4 = ~n_5115;
assign n_5126 = ~n_5078 & n_5116;
assign n_5127 = ~n_5117 & ~n_5098;
assign n_5128 = ~n_18 & ~n_5118;
assign n_5129 = n_5120 ^ n_5103;
assign n_5130 = n_4808 ^ n_5122;
assign n_5131 = ~n_5123 & ~n_4910;
assign n_5132 = n_4695 ^ n_5124;
assign n_5133 = n_5124 & n_4695;
assign n_5134 = ~n_5125 & n_4912;
assign n_5135 = n_5100 ^ n_5126;
assign n_5136 = n_5111 ^ n_5127;
assign n_5137 = ~n_5128 & ~n_5119;
assign n_5138 = n_5070 ^ n_5129;
assign n_5139 = n_5058 ^ n_5129;
assign n_5140 = n_5130 ^ n_2067;
assign n_5141 = n_4850 ^ n_5131;
assign n_5142 = ~n_5132 & ~n_4896;
assign n_5143 = ~n_5133 & n_5134;
assign n_5144 = n_5013 ^ n_5135;
assign y6 = ~n_5136;
assign n_5145 = n_5138 ^ n_5137;
assign n_5146 = ~n_5138 & n_5118;
assign n_5147 = n_5138 & n_5119;
assign n_5148 = ~n_5070 & n_5139;
assign n_5149 = n_5141 ^ n_4897;
assign n_5150 = n_4829 ^ n_5142;
assign n_5151 = n_4791 ^ n_5143;
assign n_5152 = n_4770 ^ n_5143;
assign y5 = n_5144;
assign y7 = ~n_5145;
assign n_5153 = ~n_18 & ~n_5146;
assign n_5154 = n_18 & ~n_5147;
assign n_5155 = n_5148 ^ n_5129;
assign n_5156 = n_5149 ^ n_5150;
assign n_5157 = n_5151 ^ ~n_1879;
assign n_5158 = n_4791 & ~n_5152;
assign n_5159 = n_5153 ^ n_18;
assign n_5160 = n_5154 ^ n_5059;
assign n_5161 = n_5155 ^ n_5059;
assign n_5162 = ~n_5059 & n_5155;
assign n_5163 = n_5095 ^ n_5155;
assign n_5164 = n_5060 ^ n_5155;
assign n_5165 = n_5156 ^ n_1914;
assign n_5166 = n_5158 ^ n_5143;
assign n_5167 = n_5159 ^ n_5154;
assign n_5168 = n_5160 ^ n_5153;
assign n_5169 = n_5146 & ~n_5162;
assign n_5170 = n_5104 & n_5163;
assign n_5171 = n_5162 ^ n_5164;
assign n_5172 = n_5166 & ~n_4881;
assign n_5173 = ~n_5166 & n_4928;
assign n_5174 = n_5167 ^ n_5161;
assign n_5175 = n_5161 & ~n_5168;
assign n_5176 = n_5170 ^ n_5071;
assign n_5177 = n_5105 ^ n_5170;
assign n_5178 = n_5171 ^ n_1951;
assign n_5179 = ~n_4856 & ~n_5172;
assign n_5180 = n_4924 ^ n_5173;
assign y8 = n_5174;
assign n_5181 = n_5175 ^ n_5153;
assign n_5182 = n_5095 & n_5176;
assign n_5183 = n_5147 & n_5177;
assign n_5184 = n_5095 & ~n_5178;
assign n_5185 = n_5179 ^ n_4541;
assign n_5186 = n_5180 ^ n_2100;
assign n_5187 = n_5071 ^ n_5181;
assign n_5188 = n_5182 ^ n_5071;
assign n_5189 = n_5184 ^ n_5085;
assign n_5190 = n_5185 ^ n_2034;
assign n_5191 = n_5095 ^ n_5187;
assign n_5192 = n_5169 & ~n_5188;
assign n_5193 = n_5086 ^ n_5189;
assign n_5194 = n_5073 ^ n_5189;
assign y9 = n_5191;
assign n_5195 = ~n_18 & ~n_5192;
assign n_5196 = ~n_5193 & n_5192;
assign n_5197 = n_5193 & n_5183;
assign n_5198 = ~n_5086 & n_5194;
assign n_5199 = ~n_5195 & ~n_5183;
assign n_5200 = ~n_18 & ~n_5196;
assign n_5201 = n_5198 ^ n_5189;
assign n_5202 = n_5193 ^ n_5199;
assign n_5203 = ~n_5200 & ~n_5197;
assign n_5204 = n_5121 ^ n_5201;
assign n_5205 = n_5113 ^ n_5201;
assign y10 = ~n_5202;
assign n_5206 = n_5204 ^ n_5203;
assign n_5207 = ~n_5204 & n_5196;
assign n_5208 = n_5204 & n_5197;
assign n_5209 = ~n_5121 & n_5205;
assign y11 = ~n_5206;
assign n_5210 = ~n_18 & ~n_5207;
assign n_5211 = n_5209 ^ n_5201;
assign n_5212 = ~n_5210 & ~n_5208;
assign n_5213 = n_5140 ^ n_5211;
assign n_5214 = n_5130 ^ n_5211;
assign n_5215 = n_5213 ^ n_5212;
assign n_5216 = ~n_5213 & n_5207;
assign n_5217 = n_5213 & n_5208;
assign n_5218 = ~n_5140 & n_5214;
assign y12 = ~n_5215;
assign n_5219 = ~n_18 & ~n_5216;
assign n_5220 = n_5218 ^ n_5211;
assign n_5221 = ~n_5219 & ~n_5217;
assign n_5222 = n_5165 ^ n_5220;
assign n_5223 = n_5156 ^ n_5220;
assign n_5224 = n_5222 ^ n_5221;
assign n_5225 = ~n_5222 & n_5216;
assign n_5226 = n_5222 & n_5217;
assign n_5227 = ~n_5165 & n_5223;
assign y13 = ~n_5224;
assign n_5228 = ~n_18 & ~n_5225;
assign n_5229 = n_5227 ^ n_5220;
assign n_5230 = ~n_5228 & ~n_5226;
assign n_5231 = n_5157 ^ n_5229;
assign n_5232 = n_5151 ^ n_5229;
assign n_5233 = n_5231 ^ n_5230;
assign n_5234 = ~n_5231 & n_5226;
assign n_5235 = n_5231 & n_5225;
assign n_5236 = n_5157 & ~n_5232;
assign y14 = n_5233;
assign n_5237 = n_18 & ~n_5234;
assign n_5238 = n_5236 ^ n_5229;
assign n_5239 = ~n_5237 & ~n_5235;
assign n_5240 = n_5186 ^ n_5238;
assign n_5241 = n_5180 ^ n_5238;
assign n_5242 = n_5240 ^ n_5239;
assign n_5243 = n_5240 & n_5235;
assign n_5244 = ~n_5240 & n_5234;
assign n_5245 = n_5186 & ~n_5241;
assign y15 = ~n_5242;
assign n_5246 = ~n_18 & ~n_5243;
assign n_5247 = n_5245 ^ n_5238;
assign n_5248 = ~n_5246 & ~n_5244;
assign n_5249 = n_5190 ^ n_5247;
assign n_5250 = n_5185 ^ n_5247;
assign n_5251 = n_5249 ^ n_5248;
assign n_5252 = n_5249 & n_5244;
assign n_5253 = ~n_5249 & n_5243;
assign n_5254 = ~n_5190 & n_5250;
assign y16 = ~n_5251;
assign n_5255 = n_18 & ~n_5252;
assign n_5256 = n_5254 ^ n_5247;
assign n_5257 = ~n_5255 & ~n_5253;
assign n_5258 = ~n_1949 ^ n_5256;
assign n_5259 = n_5256 & ~n_1949;
assign n_5260 = n_5257 ^ n_5258;
assign n_5261 = n_5258 & n_5253;
assign n_5262 = n_5259 ^ n_5258;
assign n_5263 = n_5252 & n_5259;
assign y17 = ~n_5260;
assign n_5264 = n_5262 ^ n_5253;
assign n_5265 = n_5255 & ~n_5262;
assign n_5266 = ~n_1948 ^ n_5262;
assign n_5267 = n_1948 ^ ~n_5263;
assign n_5268 = n_5264 ^ n_5261;
assign n_5269 = n_5263 ^ n_5265;
assign n_5270 = n_5252 & n_5266;
assign n_5271 = n_5268 ^ n_5253;
assign n_5272 = ~n_5261 ^ ~n_5270;
assign n_5273 = ~n_18 & n_5271;
assign n_5274 = ~n_1948 & ~n_5271;
assign n_5275 = n_5272 & n_5267;
assign n_5276 = ~n_5273 & ~n_5269;
assign n_5277 = n_5274 ^ n_1980;
assign n_5278 = ~n_5274 & ~n_2102;
assign n_5279 = n_5274 ^ n_18;
assign n_5280 = n_5274 & n_2243;
assign n_5281 = ~n_5274 & n_2294;
assign n_5282 = n_18 & ~n_5275;
assign n_5283 = n_1948 ^ n_5276;
assign n_5284 = n_2174 ^ n_5278;
assign n_5285 = n_2041 ^ n_5280;
assign n_5286 = ~n_5280 & n_2041;
assign n_5287 = n_2243 ^ n_5281;
assign n_5288 = n_5282 ^ n_5277;
assign n_5289 = n_5282 ^ n_18;
assign n_5290 = n_5279 ^ n_5282;
assign y18 = ~n_5283;
assign n_5291 = n_5286 ^ n_5285;
assign n_5292 = ~n_17 & n_5286;
assign n_5293 = n_5287 & n_5275;
assign y19 = ~n_5288;
assign n_5294 = n_5289 ^ n_1980;
assign n_5295 = ~n_5284 & n_5290;
assign n_5296 = ~n_5289 & n_5291;
assign n_5297 = n_18 & ~n_5293;
assign n_5298 = n_5292 & n_5293;
assign n_5299 = n_5277 & ~n_5294;
assign n_5300 = n_18 ^ n_5295;
assign n_5301 = n_5296 ^ n_18;
assign n_5302 = n_5285 ^ n_5297;
assign n_5303 = n_18 & ~n_5298;
assign n_5304 = n_5299 ^ n_18;
assign n_5305 = n_5300 ^ n_2121;
assign n_5306 = ~n_2042 & ~n_5301;
assign y22 = ~n_5302;
assign y24 = n_5303;
assign n_5307 = n_5304 ^ n_1885;
assign y21 = ~n_5305;
assign n_5308 = ~n_5306 & ~n_5298;
assign y20 = ~n_5307;
assign y23 = n_5308;
endmodule