module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 ;
  assign n18 = x9 ^ x1 ;
  assign n17 = x0 & x8 ;
  assign n19 = n18 ^ n17 ;
  assign n22 = x10 ^ x2 ;
  assign n21 = x1 & x9 ;
  assign n23 = n22 ^ n21 ;
  assign n20 = n17 & n18 ;
  assign n24 = n23 ^ n20 ;
  assign n31 = x11 ^ x3 ;
  assign n30 = x2 & x10 ;
  assign n32 = n31 ^ n30 ;
  assign n28 = n21 & n22 ;
  assign n25 = x0 & n18 ;
  assign n26 = x8 & n22 ;
  assign n27 = n25 & n26 ;
  assign n29 = n28 ^ n27 ;
  assign n33 = n32 ^ n29 ;
  assign n38 = x12 ^ x4 ;
  assign n37 = x3 & x11 ;
  assign n39 = n38 ^ n37 ;
  assign n35 = n29 & n32 ;
  assign n34 = n30 & n31 ;
  assign n36 = n35 ^ n34 ;
  assign n40 = n39 ^ n36 ;
  assign n48 = x13 ^ x5 ;
  assign n47 = x4 & x12 ;
  assign n49 = n48 ^ n47 ;
  assign n44 = n34 & n39 ;
  assign n43 = n37 & n38 ;
  assign n45 = n44 ^ n43 ;
  assign n41 = n32 & n39 ;
  assign n42 = n29 & n41 ;
  assign n46 = n45 ^ n42 ;
  assign n50 = n49 ^ n46 ;
  assign n55 = x14 ^ x6 ;
  assign n54 = x5 & x13 ;
  assign n56 = n55 ^ n54 ;
  assign n52 = n46 & n49 ;
  assign n51 = n47 & n48 ;
  assign n53 = n52 ^ n51 ;
  assign n57 = n56 ^ n53 ;
  assign n65 = x15 ^ x7 ;
  assign n64 = x6 & x14 ;
  assign n66 = n65 ^ n64 ;
  assign n61 = n51 & n56 ;
  assign n60 = n54 & n55 ;
  assign n62 = n61 ^ n60 ;
  assign n58 = n49 & n56 ;
  assign n59 = n46 & n58 ;
  assign n63 = n62 ^ n59 ;
  assign n67 = n66 ^ n63 ;
  assign n74 = x7 & x15 ;
  assign n75 = n74 ^ n65 ;
  assign n71 = n62 & n66 ;
  assign n70 = n64 & n65 ;
  assign n72 = n71 ^ n70 ;
  assign n68 = n58 & n66 ;
  assign n69 = n46 & n68 ;
  assign n73 = n72 ^ n69 ;
  assign n76 = n75 ^ n73 ;
  assign y0 = n19 ;
  assign y1 = n24 ;
  assign y2 = n33 ;
  assign y3 = n40 ;
  assign y4 = n50 ;
  assign y5 = n57 ;
  assign y6 = n67 ;
  assign y7 = n76 ;
endmodule
