module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 ;
  assign n15 = x1 & x9 ;
  assign n16 = n15 ^ x9 ;
  assign n202 = x0 & x2 ;
  assign n203 = n202 ^ x0 ;
  assign n204 = n203 ^ x2 ;
  assign n214 = n16 & ~n204 ;
  assign n215 = ~x5 & x6 ;
  assign n216 = ~n214 & n215 ;
  assign n217 = n216 ^ x6 ;
  assign n218 = x9 ^ x0 ;
  assign n219 = x1 & x5 ;
  assign n220 = x2 & n219 ;
  assign n221 = ~n218 & n220 ;
  assign n222 = n217 & n221 ;
  assign n223 = n222 ^ n217 ;
  assign n224 = n223 ^ n221 ;
  assign n225 = x8 & ~n224 ;
  assign n226 = n225 ^ x8 ;
  assign n11 = x0 & x9 ;
  assign n12 = n11 ^ x9 ;
  assign n227 = ~x1 & ~n12 ;
  assign n228 = ~x8 & ~n227 ;
  assign n24 = n11 ^ x0 ;
  assign n229 = ~x1 & x2 ;
  assign n230 = n24 & n229 ;
  assign n231 = ~n228 & ~n230 ;
  assign n232 = ~x5 & ~n231 ;
  assign n233 = n226 & n232 ;
  assign n234 = n233 ^ n226 ;
  assign n235 = n234 ^ n232 ;
  assign n236 = x3 & ~n235 ;
  assign n237 = n236 ^ x3 ;
  assign n238 = x2 & n24 ;
  assign n239 = n238 ^ x2 ;
  assign n240 = n239 ^ n24 ;
  assign n241 = x1 & ~x3 ;
  assign n242 = ~n12 & n241 ;
  assign n243 = ~n240 & n242 ;
  assign n244 = n243 ^ n240 ;
  assign n245 = ~x2 & ~x6 ;
  assign n246 = ~n24 & n245 ;
  assign n247 = n246 ^ x6 ;
  assign n248 = x5 & ~n247 ;
  assign n249 = n248 ^ x5 ;
  assign n250 = ~n244 & n249 ;
  assign n251 = n250 ^ n249 ;
  assign n125 = x2 & x9 ;
  assign n28 = n15 ^ x1 ;
  assign n252 = ~x2 & n28 ;
  assign n253 = ~n125 & ~n252 ;
  assign n254 = x0 & x3 ;
  assign n255 = n254 ^ x0 ;
  assign n256 = n255 ^ x3 ;
  assign n257 = x6 & ~n256 ;
  assign n258 = ~n253 & n257 ;
  assign n259 = n251 & n258 ;
  assign n260 = n259 ^ n251 ;
  assign n261 = n260 ^ n258 ;
  assign n262 = x8 & ~n261 ;
  assign n263 = n262 ^ x8 ;
  assign n264 = x1 & ~x8 ;
  assign n265 = x2 & ~x3 ;
  assign n266 = n16 & n265 ;
  assign n267 = ~n264 & ~n266 ;
  assign n268 = ~x0 & ~n267 ;
  assign n269 = x2 & x6 ;
  assign n270 = n269 ^ x6 ;
  assign n271 = x3 & n270 ;
  assign n272 = n271 ^ x3 ;
  assign n273 = n28 ^ x9 ;
  assign n274 = ~n125 & ~n273 ;
  assign n275 = ~n272 & n274 ;
  assign n276 = n275 ^ n125 ;
  assign n277 = x8 & ~n276 ;
  assign n278 = n277 ^ x8 ;
  assign n279 = n278 ^ n276 ;
  assign n280 = n268 & n279 ;
  assign n281 = n280 ^ n268 ;
  assign n282 = n281 ^ n279 ;
  assign n283 = x8 & ~n273 ;
  assign n284 = n283 ^ n273 ;
  assign n285 = x2 & x3 ;
  assign n286 = n285 ^ x2 ;
  assign n287 = n286 ^ x3 ;
  assign n288 = ~x0 & ~n287 ;
  assign n289 = ~n284 & n288 ;
  assign n290 = ~x5 & ~n289 ;
  assign n291 = n282 & n290 ;
  assign n292 = n291 ^ n289 ;
  assign n293 = n263 & n292 ;
  assign n294 = n293 ^ n263 ;
  assign n295 = n294 ^ n292 ;
  assign n296 = n237 & n295 ;
  assign n297 = n296 ^ n237 ;
  assign n298 = n297 ^ n295 ;
  assign n318 = x7 & n298 ;
  assign n319 = n318 ^ x7 ;
  assign n320 = n319 ^ x7 ;
  assign n321 = n320 ^ n298 ;
  assign n13 = x1 & n12 ;
  assign n14 = n13 ^ x1 ;
  assign n17 = x3 & x5 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = n18 ^ x5 ;
  assign n20 = n16 & ~n19 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n14 & ~n21 ;
  assign n23 = n22 ^ n21 ;
  assign n25 = x1 & n24 ;
  assign n26 = n25 ^ x1 ;
  assign n27 = n26 ^ n24 ;
  assign n29 = x7 & n28 ;
  assign n30 = n29 ^ x7 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = ~n27 & ~n31 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = ~n23 & ~n33 ;
  assign n35 = n34 ^ n23 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = x2 & ~n36 ;
  assign n38 = n37 ^ x2 ;
  assign n39 = n38 ^ n36 ;
  assign n41 = x2 ^ x0 ;
  assign n60 = x5 ^ x2 ;
  assign n58 = x5 ^ x1 ;
  assign n59 = n58 ^ x5 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = n59 ^ x5 ;
  assign n63 = ~n61 & ~n62 ;
  assign n64 = n63 ^ n59 ;
  assign n65 = ~n41 & ~n64 ;
  assign n66 = n65 ^ x2 ;
  assign n67 = n66 ^ x5 ;
  assign n68 = n67 ^ x5 ;
  assign n73 = n68 ^ x9 ;
  assign n43 = x9 ^ x2 ;
  assign n42 = n41 ^ x2 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n43 ^ x2 ;
  assign n46 = n44 & n45 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = n47 ^ n43 ;
  assign n49 = x9 ^ x3 ;
  assign n50 = x1 & n49 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n48 & n51 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n53 ^ x1 ;
  assign n55 = n54 ^ n49 ;
  assign n56 = n55 ^ x9 ;
  assign n57 = n56 ^ x9 ;
  assign n99 = n56 & n57 ;
  assign n100 = n99 ^ n56 ;
  assign n101 = n100 ^ n56 ;
  assign n102 = n101 ^ n68 ;
  assign n103 = ~n73 & ~n102 ;
  assign n104 = n103 ^ n73 ;
  assign n105 = n104 ^ n100 ;
  assign n106 = n105 ^ n68 ;
  assign n74 = n73 ^ n56 ;
  assign n89 = n74 ^ x7 ;
  assign n75 = n74 ^ n56 ;
  assign n82 = n75 ^ x7 ;
  assign n83 = ~n75 & ~n82 ;
  assign n69 = n68 ^ n57 ;
  assign n91 = n83 ^ n69 ;
  assign n70 = n69 ^ n68 ;
  assign n90 = n70 ^ x7 ;
  assign n92 = n91 ^ n90 ;
  assign n93 = n89 & ~n92 ;
  assign n77 = n74 ^ n70 ;
  assign n78 = n77 ^ n75 ;
  assign n79 = n75 ^ n70 ;
  assign n80 = n79 ^ x7 ;
  assign n81 = ~n78 & ~n80 ;
  assign n84 = n83 ^ n81 ;
  assign n85 = n84 ^ n69 ;
  assign n76 = n75 ^ n74 ;
  assign n86 = n85 ^ n76 ;
  assign n87 = n81 ^ n69 ;
  assign n88 = n86 & ~n87 ;
  assign n94 = n93 ^ n88 ;
  assign n95 = n94 ^ n83 ;
  assign n71 = n70 ^ n69 ;
  assign n72 = n71 ^ x7 ;
  assign n96 = n95 ^ n72 ;
  assign n97 = n96 ^ x7 ;
  assign n98 = n97 ^ x7 ;
  assign n107 = n106 ^ n98 ;
  assign n115 = n39 & ~n107 ;
  assign n116 = n115 ^ n39 ;
  assign n117 = n116 ^ n39 ;
  assign n118 = n117 ^ n107 ;
  assign n40 = n39 ^ x8 ;
  assign n108 = n107 ^ x8 ;
  assign n109 = n107 & ~n108 ;
  assign n110 = n109 ^ x8 ;
  assign n111 = ~n40 & ~n110 ;
  assign n112 = n111 ^ n109 ;
  assign n113 = n112 ^ n39 ;
  assign n114 = n113 ^ x8 ;
  assign n119 = n118 ^ n114 ;
  assign n120 = n119 ^ x6 ;
  assign n182 = x6 & n120 ;
  assign n129 = x0 & ~x2 ;
  assign n131 = x9 ^ x5 ;
  assign n132 = n131 ^ x9 ;
  assign n130 = x9 ^ x7 ;
  assign n133 = n132 ^ n130 ;
  assign n135 = n133 ^ x9 ;
  assign n137 = n135 ^ n133 ;
  assign n134 = n133 ^ n132 ;
  assign n138 = n134 ^ n133 ;
  assign n139 = ~n137 & n138 ;
  assign n140 = n139 ^ n133 ;
  assign n143 = n139 ^ n134 ;
  assign n141 = n131 ^ x1 ;
  assign n142 = n141 ^ n135 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = ~n140 & n144 ;
  assign n146 = n145 ^ n139 ;
  assign n136 = n135 ^ n134 ;
  assign n147 = n146 ^ n136 ;
  assign n150 = n143 ^ n135 ;
  assign n151 = n141 ^ n134 ;
  assign n148 = n133 ^ x8 ;
  assign n152 = n151 ^ n148 ;
  assign n153 = ~n150 & n152 ;
  assign n154 = n153 ^ n145 ;
  assign n155 = n154 ^ n139 ;
  assign n149 = n148 ^ n134 ;
  assign n156 = n155 ^ n149 ;
  assign n157 = ~n147 & ~n156 ;
  assign n158 = n157 ^ n145 ;
  assign n159 = n158 ^ n133 ;
  assign n160 = n159 ^ n131 ;
  assign n161 = n160 ^ x9 ;
  assign n162 = n161 ^ n141 ;
  assign n163 = n162 ^ n135 ;
  assign n164 = n163 ^ n134 ;
  assign n165 = n164 ^ n133 ;
  assign n166 = n129 & ~n165 ;
  assign n167 = n166 ^ n129 ;
  assign n121 = x5 & x7 ;
  assign n122 = n121 ^ x7 ;
  assign n123 = x8 & n122 ;
  assign n124 = ~x0 & ~x1 ;
  assign n126 = n125 ^ x2 ;
  assign n127 = n124 & n126 ;
  assign n128 = n123 & n127 ;
  assign n168 = n167 ^ n128 ;
  assign n169 = n128 ^ x3 ;
  assign n170 = x3 & ~n169 ;
  assign n171 = n170 ^ x3 ;
  assign n172 = n171 ^ n167 ;
  assign n173 = n168 & ~n172 ;
  assign n174 = n173 ^ n170 ;
  assign n175 = n174 ^ n167 ;
  assign n176 = n175 ^ x6 ;
  assign n177 = ~x6 & ~n176 ;
  assign n178 = n177 ^ n119 ;
  assign n179 = ~n120 & n178 ;
  assign n180 = n179 ^ n177 ;
  assign n181 = n180 ^ n175 ;
  assign n183 = n182 ^ n181 ;
  assign n184 = n183 ^ n175 ;
  assign n322 = x4 & ~n184 ;
  assign n323 = n322 ^ x4 ;
  assign n324 = n323 ^ n184 ;
  assign n325 = n321 & n324 ;
  assign n326 = n325 ^ n324 ;
  assign n327 = n326 ^ x4 ;
  assign n186 = ~x6 & x8 ;
  assign n187 = x5 & ~n186 ;
  assign n188 = x4 & x8 ;
  assign n189 = x6 & x9 ;
  assign n190 = n189 ^ x6 ;
  assign n191 = n190 ^ x9 ;
  assign n192 = ~n188 & n191 ;
  assign n193 = n187 & ~n192 ;
  assign n194 = x6 & ~x9 ;
  assign n195 = x4 & x9 ;
  assign n196 = ~n194 & ~n195 ;
  assign n197 = x5 & x6 ;
  assign n198 = ~x8 & ~n197 ;
  assign n199 = ~n196 & n198 ;
  assign n200 = ~n193 & ~n199 ;
  assign n201 = ~x1 & ~x3 ;
  assign n205 = ~x7 & ~n204 ;
  assign n206 = n201 & n205 ;
  assign n207 = ~n200 & n206 ;
  assign n210 = n207 ^ n184 ;
  assign n304 = n210 ^ x4 ;
  assign n211 = n207 ^ x7 ;
  assign n212 = n210 & ~n211 ;
  assign n213 = n212 ^ x7 ;
  assign n299 = n298 ^ n213 ;
  assign n305 = n304 ^ n299 ;
  assign n306 = n298 ^ n184 ;
  assign n307 = n306 ^ n213 ;
  assign n308 = n305 & ~n307 ;
  assign n300 = n213 ^ n184 ;
  assign n208 = n207 ^ x4 ;
  assign n301 = n300 ^ n208 ;
  assign n302 = ~n299 & n301 ;
  assign n309 = n308 ^ n302 ;
  assign n310 = n309 ^ n213 ;
  assign n311 = n310 ^ n304 ;
  assign n312 = n302 ^ n298 ;
  assign n313 = n312 ^ x4 ;
  assign n314 = n311 & ~n313 ;
  assign n315 = n314 ^ n308 ;
  assign n303 = n302 ^ n212 ;
  assign n316 = n315 ^ n303 ;
  assign n185 = n184 ^ x7 ;
  assign n209 = n208 ^ n185 ;
  assign n317 = n316 ^ n209 ;
  assign n328 = n327 ^ n317 ;
  assign n329 = n328 ^ n207 ;
  assign n343 = n218 ^ x9 ;
  assign n347 = x9 ^ x6 ;
  assign n342 = x6 ^ x5 ;
  assign n348 = n347 ^ n342 ;
  assign n349 = n348 ^ x8 ;
  assign n350 = n349 ^ x8 ;
  assign n351 = n350 ^ n218 ;
  assign n352 = n351 ^ n343 ;
  assign n353 = n349 & n352 ;
  assign n354 = n353 ^ n349 ;
  assign n355 = n354 ^ n343 ;
  assign n356 = n355 ^ n349 ;
  assign n357 = n343 & n356 ;
  assign n358 = n357 ^ n343 ;
  assign n359 = n358 ^ n356 ;
  assign n345 = n342 ^ x9 ;
  assign n346 = ~n342 & ~n345 ;
  assign n360 = n359 ^ n346 ;
  assign n361 = n360 ^ n354 ;
  assign n344 = n343 ^ n342 ;
  assign n362 = n361 ^ n344 ;
  assign n364 = n359 ^ n343 ;
  assign n363 = n351 ^ n349 ;
  assign n365 = n364 ^ n363 ;
  assign n366 = ~n362 & ~n365 ;
  assign n367 = n366 ^ n362 ;
  assign n368 = n367 ^ n359 ;
  assign n369 = n368 ^ n355 ;
  assign n370 = n369 ^ x5 ;
  assign n371 = n370 ^ x9 ;
  assign n372 = n371 ^ x9 ;
  assign n373 = n43 & n218 ;
  assign n374 = n373 ^ n218 ;
  assign n375 = n374 ^ n43 ;
  assign n376 = x9 ^ x8 ;
  assign n377 = x5 & n376 ;
  assign n378 = n377 ^ x5 ;
  assign n379 = ~n375 & n378 ;
  assign n380 = x2 & n379 ;
  assign n381 = n380 ^ x2 ;
  assign n382 = n372 & n381 ;
  assign n383 = n382 ^ n379 ;
  assign n384 = n126 & n186 ;
  assign n385 = ~x1 & ~n384 ;
  assign n386 = n383 & n385 ;
  assign n387 = n386 ^ n384 ;
  assign n460 = n387 ^ x1 ;
  assign n330 = ~x2 & n124 ;
  assign n331 = x5 ^ x4 ;
  assign n332 = x8 & n331 ;
  assign n333 = n332 ^ x5 ;
  assign n334 = ~n191 & ~n333 ;
  assign n335 = n334 ^ n191 ;
  assign n336 = x4 & n189 ;
  assign n337 = ~n335 & n336 ;
  assign n338 = n337 ^ n335 ;
  assign n339 = n338 ^ n336 ;
  assign n340 = n330 & n339 ;
  assign n341 = n340 ^ n330 ;
  assign n440 = n341 ^ x4 ;
  assign n461 = n460 ^ n440 ;
  assign n388 = n387 ^ n341 ;
  assign n446 = n388 ^ x4 ;
  assign n399 = x8 ^ x0 ;
  assign n397 = n376 ^ n347 ;
  assign n393 = n347 ^ n131 ;
  assign n394 = n393 ^ x8 ;
  assign n395 = n394 ^ x9 ;
  assign n396 = n395 ^ n376 ;
  assign n398 = n397 ^ n396 ;
  assign n400 = n399 ^ n398 ;
  assign n401 = n400 ^ n398 ;
  assign n402 = n400 ^ n397 ;
  assign n403 = n401 & n402 ;
  assign n404 = n403 ^ n400 ;
  assign n412 = n402 ^ n401 ;
  assign n413 = n412 ^ n400 ;
  assign n405 = n400 ^ n376 ;
  assign n406 = n405 ^ n402 ;
  assign n407 = n406 ^ n401 ;
  assign n408 = n400 ^ x9 ;
  assign n409 = n408 ^ n402 ;
  assign n410 = n409 ^ n401 ;
  assign n411 = n407 & n410 ;
  assign n414 = n413 ^ n411 ;
  assign n415 = n404 & n414 ;
  assign n416 = n415 ^ n400 ;
  assign n417 = n416 ^ n400 ;
  assign n418 = x2 & ~n417 ;
  assign n419 = n418 ^ x2 ;
  assign n420 = n419 ^ n417 ;
  assign n421 = x0 & x6 ;
  assign n422 = n421 ^ x6 ;
  assign n423 = x2 & n422 ;
  assign n424 = n423 ^ x2 ;
  assign n425 = n424 ^ n422 ;
  assign n426 = x5 & x8 ;
  assign n427 = n426 ^ x8 ;
  assign n428 = ~x6 & ~x8 ;
  assign n429 = n427 & ~n428 ;
  assign n430 = n425 & n429 ;
  assign n431 = n430 ^ n428 ;
  assign n432 = x9 & ~n431 ;
  assign n433 = n432 ^ x9 ;
  assign n434 = n433 ^ n431 ;
  assign n435 = n420 & n434 ;
  assign n436 = n435 ^ n420 ;
  assign n437 = n436 ^ n434 ;
  assign n389 = n341 ^ x1 ;
  assign n390 = n388 & n389 ;
  assign n391 = n390 ^ n388 ;
  assign n392 = n391 ^ x1 ;
  assign n438 = n437 ^ n392 ;
  assign n447 = n446 ^ n438 ;
  assign n448 = n437 ^ n387 ;
  assign n449 = n448 ^ n392 ;
  assign n450 = ~n447 & ~n449 ;
  assign n439 = n392 ^ n387 ;
  assign n441 = n440 ^ n439 ;
  assign n442 = ~n438 & n441 ;
  assign n443 = n442 ^ n438 ;
  assign n444 = n443 ^ n441 ;
  assign n451 = n450 ^ n444 ;
  assign n452 = n451 ^ n392 ;
  assign n453 = n452 ^ n446 ;
  assign n454 = n444 ^ n437 ;
  assign n455 = n454 ^ x4 ;
  assign n456 = n453 & ~n455 ;
  assign n457 = n456 ^ n455 ;
  assign n458 = n457 ^ n450 ;
  assign n445 = n444 ^ n391 ;
  assign n459 = n458 ^ n445 ;
  assign n462 = n461 ^ n459 ;
  assign n463 = n462 ^ n341 ;
  assign n574 = x3 & ~n463 ;
  assign n575 = n574 ^ x3 ;
  assign n576 = n575 ^ n463 ;
  assign n464 = n463 ^ x3 ;
  assign n465 = x2 & x8 ;
  assign n475 = n465 ^ x8 ;
  assign n476 = n475 ^ x0 ;
  assign n477 = x5 ^ x0 ;
  assign n478 = n477 ^ x0 ;
  assign n479 = n477 & n478 ;
  assign n480 = n479 ^ n477 ;
  assign n481 = n480 ^ n475 ;
  assign n482 = n476 & n481 ;
  assign n483 = n482 ^ n479 ;
  assign n484 = n483 ^ n475 ;
  assign n487 = n484 ^ x1 ;
  assign n466 = n465 ^ x2 ;
  assign n467 = n466 ^ x8 ;
  assign n468 = x5 & ~n467 ;
  assign n469 = x5 ^ x3 ;
  assign n470 = x8 & n469 ;
  assign n471 = n470 ^ n469 ;
  assign n472 = n471 ^ x5 ;
  assign n473 = x0 & n472 ;
  assign n474 = ~n468 & ~n473 ;
  assign n485 = n484 ^ n474 ;
  assign n486 = n485 ^ n484 ;
  assign n488 = n487 ^ n486 ;
  assign n489 = n486 ^ n484 ;
  assign n490 = n488 & ~n489 ;
  assign n491 = n490 ^ n486 ;
  assign n492 = x3 & x8 ;
  assign n493 = ~x2 & ~n492 ;
  assign n494 = ~x0 & ~n493 ;
  assign n495 = ~x6 & ~n494 ;
  assign n496 = n491 & n495 ;
  assign n497 = n496 ^ x6 ;
  assign n498 = ~x5 & ~x9 ;
  assign n499 = x8 ^ x2 ;
  assign n500 = n499 ^ x8 ;
  assign n501 = n500 ^ x1 ;
  assign n504 = n501 ^ n500 ;
  assign n502 = n501 ^ x8 ;
  assign n505 = n504 ^ n502 ;
  assign n506 = n504 ^ x6 ;
  assign n507 = n505 ^ x3 ;
  assign n508 = n506 & n507 ;
  assign n509 = n508 ^ x6 ;
  assign n510 = n509 ^ n505 ;
  assign n511 = n505 & ~n510 ;
  assign n512 = n511 ^ n508 ;
  assign n513 = n512 ^ x6 ;
  assign n503 = n502 ^ n501 ;
  assign n514 = n513 ^ n503 ;
  assign n515 = n504 ^ n501 ;
  assign n517 = n502 ^ x6 ;
  assign n516 = n504 ^ x3 ;
  assign n518 = n517 ^ n516 ;
  assign n519 = ~n515 & ~n518 ;
  assign n520 = n519 ^ n511 ;
  assign n521 = n520 ^ n508 ;
  assign n522 = n514 & n521 ;
  assign n523 = x0 & x8 ;
  assign n524 = n523 ^ x8 ;
  assign n525 = ~x2 & ~n524 ;
  assign n526 = x0 & x1 ;
  assign n527 = ~x1 & ~x6 ;
  assign n528 = ~n526 & ~n527 ;
  assign n529 = n525 & n528 ;
  assign n530 = n522 & n529 ;
  assign n531 = n530 ^ n522 ;
  assign n532 = n531 ^ n529 ;
  assign n533 = n498 & n532 ;
  assign n534 = n533 ^ x9 ;
  assign n535 = ~n497 & ~n534 ;
  assign n536 = n535 ^ n534 ;
  assign n542 = x1 & x3 ;
  assign n543 = n542 ^ x3 ;
  assign n544 = ~n467 & n543 ;
  assign n545 = x0 & ~n219 ;
  assign n546 = ~n544 & n545 ;
  assign n547 = n546 ^ x0 ;
  assign n538 = x1 & x2 ;
  assign n548 = x3 & ~x5 ;
  assign n549 = n538 & n548 ;
  assign n550 = n549 ^ x5 ;
  assign n551 = n287 & ~n550 ;
  assign n552 = n551 ^ n287 ;
  assign n553 = n547 & n552 ;
  assign n554 = n553 ^ n547 ;
  assign n555 = n554 ^ n552 ;
  assign n556 = x6 & ~n555 ;
  assign n557 = n556 ^ x6 ;
  assign n537 = n426 ^ x5 ;
  assign n539 = x3 & n538 ;
  assign n540 = n537 & n539 ;
  assign n541 = x9 & ~n540 ;
  assign n558 = n557 ^ n541 ;
  assign n559 = n541 ^ x4 ;
  assign n560 = x4 & n559 ;
  assign n561 = n560 ^ x4 ;
  assign n562 = n561 ^ n557 ;
  assign n563 = ~n558 & ~n562 ;
  assign n564 = n563 ^ n560 ;
  assign n565 = n564 ^ n557 ;
  assign n566 = ~n536 & n565 ;
  assign n567 = n566 ^ n565 ;
  assign n568 = n567 ^ x3 ;
  assign n569 = ~n567 & ~n568 ;
  assign n570 = n569 ^ x3 ;
  assign n571 = ~n464 & n570 ;
  assign n572 = n571 ^ n569 ;
  assign n573 = n572 ^ n463 ;
  assign n577 = n576 ^ n573 ;
  assign n578 = n577 ^ n567 ;
  assign n597 = x7 & ~n578 ;
  assign n598 = n597 ^ x7 ;
  assign n599 = n598 ^ n578 ;
  assign n579 = n578 ^ x7 ;
  assign n580 = n28 & n475 ;
  assign n581 = ~n240 & ~n526 ;
  assign n582 = x2 & ~n124 ;
  assign n583 = ~x8 & ~n582 ;
  assign n584 = ~n581 & n583 ;
  assign n585 = ~n580 & ~n584 ;
  assign n586 = x7 & ~n585 ;
  assign n587 = ~n127 & ~n586 ;
  assign n588 = ~x6 & ~n19 ;
  assign n589 = ~x4 & n588 ;
  assign n590 = ~n587 & n589 ;
  assign n591 = n590 ^ x7 ;
  assign n592 = ~n590 & ~n591 ;
  assign n593 = n592 ^ x7 ;
  assign n594 = ~n579 & n593 ;
  assign n595 = n594 ^ n592 ;
  assign n596 = n595 ^ n578 ;
  assign n600 = n599 ^ n596 ;
  assign n601 = n600 ^ n590 ;
  assign n602 = x2 & ~n186 ;
  assign n603 = x1 & ~n602 ;
  assign n604 = x5 & ~n493 ;
  assign n605 = ~n603 & n604 ;
  assign n606 = x3 & ~x8 ;
  assign n607 = ~n28 & ~n606 ;
  assign n608 = x3 & ~x9 ;
  assign n609 = ~x6 & ~n608 ;
  assign n610 = ~n607 & n609 ;
  assign n611 = x3 & x9 ;
  assign n612 = n611 ^ x9 ;
  assign n613 = x1 & n612 ;
  assign n614 = x6 & ~x8 ;
  assign n615 = ~x4 & n614 ;
  assign n616 = n613 & n615 ;
  assign n617 = n616 ^ x4 ;
  assign n618 = n610 & ~n617 ;
  assign n619 = n618 ^ n617 ;
  assign n620 = n605 & ~n619 ;
  assign n621 = n620 ^ n619 ;
  assign n622 = x1 & x8 ;
  assign n623 = n622 ^ x1 ;
  assign n624 = n623 ^ x8 ;
  assign n625 = ~x3 & n215 ;
  assign n626 = ~n624 & n625 ;
  assign n632 = x8 ^ x3 ;
  assign n633 = n632 ^ x8 ;
  assign n648 = n633 ^ x1 ;
  assign n634 = n633 ^ x8 ;
  assign n641 = n634 ^ x1 ;
  assign n642 = n634 & n641 ;
  assign n627 = x8 ^ x5 ;
  assign n628 = n627 ^ x2 ;
  assign n650 = n642 ^ n628 ;
  assign n629 = n628 ^ n627 ;
  assign n649 = n629 ^ x1 ;
  assign n651 = n650 ^ n649 ;
  assign n652 = ~n648 & ~n651 ;
  assign n636 = n633 ^ n629 ;
  assign n637 = n636 ^ n634 ;
  assign n638 = n634 ^ n629 ;
  assign n639 = n638 ^ x1 ;
  assign n640 = ~n637 & n639 ;
  assign n643 = n642 ^ n640 ;
  assign n644 = n643 ^ n628 ;
  assign n635 = n634 ^ n633 ;
  assign n645 = n644 ^ n635 ;
  assign n646 = n640 ^ n628 ;
  assign n647 = n645 & ~n646 ;
  assign n653 = n652 ^ n647 ;
  assign n654 = n653 ^ n642 ;
  assign n630 = n629 ^ n628 ;
  assign n631 = n630 ^ x1 ;
  assign n655 = n654 ^ n631 ;
  assign n656 = ~x9 & n655 ;
  assign n657 = ~n626 & n656 ;
  assign n658 = n657 ^ x9 ;
  assign n661 = ~x6 & ~x9 ;
  assign n659 = x9 ^ x1 ;
  assign n660 = n376 & n659 ;
  assign n663 = n661 ^ n660 ;
  assign n662 = n660 & n661 ;
  assign n664 = n663 ^ n662 ;
  assign n665 = ~n43 & n664 ;
  assign n666 = n665 ^ n43 ;
  assign n667 = n666 ^ x9 ;
  assign n668 = x3 & n667 ;
  assign n669 = n668 ^ x3 ;
  assign n670 = n658 & ~n669 ;
  assign n671 = ~n621 & n670 ;
  assign n672 = x8 & x9 ;
  assign n673 = ~n614 & ~n672 ;
  assign n674 = ~x5 & ~n673 ;
  assign n675 = ~x2 & n201 ;
  assign n676 = ~n674 & n675 ;
  assign n677 = x4 & ~n676 ;
  assign n678 = ~x0 & ~n677 ;
  assign n679 = n671 & n678 ;
  assign n680 = n679 ^ n678 ;
  assign n683 = n672 ^ x8 ;
  assign n684 = n683 ^ x9 ;
  assign n685 = x5 & n684 ;
  assign n686 = n685 ^ x5 ;
  assign n687 = n686 ^ x5 ;
  assign n681 = x0 & x5 ;
  assign n682 = n672 & n681 ;
  assign n688 = n687 ^ n682 ;
  assign n689 = x1 & ~x5 ;
  assign n690 = ~n125 & n689 ;
  assign n691 = n690 ^ x1 ;
  assign n692 = n688 & n691 ;
  assign n693 = n692 ^ n691 ;
  assign n694 = n376 ^ n273 ;
  assign n695 = n376 ^ x2 ;
  assign n696 = ~x2 & n695 ;
  assign n697 = n696 ^ x2 ;
  assign n698 = n697 ^ n273 ;
  assign n699 = ~n694 & ~n698 ;
  assign n700 = n699 ^ n696 ;
  assign n701 = n700 ^ n273 ;
  assign n702 = x3 & ~n701 ;
  assign n703 = n702 ^ x3 ;
  assign n704 = n703 ^ n701 ;
  assign n705 = n693 & n704 ;
  assign n706 = n705 ^ n704 ;
  assign n707 = n706 ^ x3 ;
  assign n708 = n622 ^ x8 ;
  assign n709 = x9 & n287 ;
  assign n710 = n709 ^ x9 ;
  assign n711 = n710 ^ x9 ;
  assign n712 = n708 & n711 ;
  assign n713 = x5 & n543 ;
  assign n714 = n713 ^ x5 ;
  assign n715 = x2 & n684 ;
  assign n716 = n715 ^ x2 ;
  assign n717 = n716 ^ n684 ;
  assign n718 = n714 & ~n717 ;
  assign n719 = n718 ^ n717 ;
  assign n720 = n712 & ~n719 ;
  assign n721 = n720 ^ n712 ;
  assign n722 = n721 ^ n719 ;
  assign n723 = x0 & n722 ;
  assign n724 = n723 ^ x0 ;
  assign n725 = n707 & n724 ;
  assign n726 = n725 ^ n724 ;
  assign n727 = n726 ^ n707 ;
  assign n728 = n727 ^ n724 ;
  assign n729 = n728 ^ x6 ;
  assign n732 = n376 ^ x9 ;
  assign n730 = n659 ^ x9 ;
  assign n733 = n732 ^ n730 ;
  assign n731 = n730 ^ n347 ;
  assign n734 = n733 ^ n731 ;
  assign n738 = n733 & n734 ;
  assign n739 = n738 ^ n733 ;
  assign n736 = n730 ^ x9 ;
  assign n737 = n736 ^ x2 ;
  assign n740 = n739 ^ n737 ;
  assign n741 = x2 & n740 ;
  assign n742 = n741 ^ x2 ;
  assign n744 = n742 ^ n731 ;
  assign n750 = n742 ^ n730 ;
  assign n751 = n750 ^ x2 ;
  assign n752 = n744 & n751 ;
  assign n753 = n752 ^ n744 ;
  assign n745 = n744 ^ x2 ;
  assign n746 = n738 ^ n730 ;
  assign n747 = n746 ^ n734 ;
  assign n748 = n745 & n747 ;
  assign n749 = n748 ^ n745 ;
  assign n754 = n753 ^ n749 ;
  assign n743 = n742 ^ n738 ;
  assign n755 = n754 ^ n743 ;
  assign n735 = n734 ^ x2 ;
  assign n756 = n755 ^ n735 ;
  assign n757 = n756 ^ x2 ;
  assign n758 = n757 ^ n376 ;
  assign n759 = n758 ^ x9 ;
  assign n760 = x3 & n759 ;
  assign n761 = n760 ^ x3 ;
  assign n762 = n761 ^ x3 ;
  assign n768 = n659 ^ x8 ;
  assign n769 = n347 ^ x9 ;
  assign n763 = x6 ^ x3 ;
  assign n764 = n763 ^ x9 ;
  assign n765 = n764 ^ x9 ;
  assign n766 = n765 ^ n347 ;
  assign n770 = n769 ^ n766 ;
  assign n771 = x8 & n770 ;
  assign n772 = n771 ^ n770 ;
  assign n773 = n772 ^ n347 ;
  assign n774 = n768 & n773 ;
  assign n775 = n774 ^ n773 ;
  assign n776 = n775 ^ n772 ;
  assign n767 = ~x8 & n766 ;
  assign n777 = n776 ^ n767 ;
  assign n778 = n777 ^ n659 ;
  assign n779 = n778 ^ x8 ;
  assign n780 = n779 ^ x9 ;
  assign n781 = n780 ^ n347 ;
  assign n782 = x0 & ~x5 ;
  assign n783 = ~x2 & n782 ;
  assign n784 = ~n781 & n783 ;
  assign n785 = n784 ^ n782 ;
  assign n786 = n762 & n785 ;
  assign n787 = n786 ^ n785 ;
  assign n788 = n787 ^ n782 ;
  assign n789 = n788 ^ x6 ;
  assign n790 = n788 & n789 ;
  assign n791 = n790 ^ n788 ;
  assign n792 = n791 ^ n788 ;
  assign n793 = n792 ^ n728 ;
  assign n794 = n729 & n793 ;
  assign n795 = n794 ^ n729 ;
  assign n796 = n795 ^ n791 ;
  assign n797 = n796 ^ n728 ;
  assign n798 = ~x4 & ~x7 ;
  assign n799 = ~n797 & n798 ;
  assign n800 = n799 ^ x7 ;
  assign n801 = n680 & ~n800 ;
  assign n802 = n801 ^ n800 ;
  assign n803 = n802 ^ x7 ;
  assign n804 = x7 & n672 ;
  assign n805 = x0 & ~n804 ;
  assign n806 = n14 & ~n805 ;
  assign n807 = n24 & ~n624 ;
  assign n808 = ~n806 & ~n807 ;
  assign n809 = ~x5 & ~x6 ;
  assign n810 = ~x4 & ~n287 ;
  assign n811 = n809 & n810 ;
  assign n812 = ~n808 & n811 ;
  assign n813 = ~n803 & n812 ;
  assign n814 = n813 ^ n812 ;
  assign n815 = n814 ^ n803 ;
  assign n816 = n815 ^ n812 ;
  assign n817 = n672 ^ x9 ;
  assign n818 = ~x3 & x5 ;
  assign n819 = n817 & n818 ;
  assign n820 = n819 ^ x3 ;
  assign n821 = x2 & ~n820 ;
  assign n822 = n821 ^ x2 ;
  assign n823 = n822 ^ n820 ;
  assign n824 = ~x6 & ~n606 ;
  assign n825 = ~n18 & ~n824 ;
  assign n826 = n823 & n825 ;
  assign n827 = n826 ^ n823 ;
  assign n828 = n827 ^ n825 ;
  assign n829 = n469 ^ n60 ;
  assign n830 = n60 ^ x5 ;
  assign n831 = n829 & n830 ;
  assign n832 = n831 ^ n60 ;
  assign n833 = ~x8 & n832 ;
  assign n834 = n833 ^ x2 ;
  assign n835 = n834 ^ x5 ;
  assign n836 = x9 & ~n835 ;
  assign n837 = n836 ^ x9 ;
  assign n838 = n837 ^ n835 ;
  assign n839 = x1 & ~n838 ;
  assign n840 = ~n828 & n839 ;
  assign n841 = n840 ^ x1 ;
  assign n842 = n468 & n527 ;
  assign n843 = ~n625 & ~n842 ;
  assign n844 = ~x9 & ~n843 ;
  assign n845 = n841 & n844 ;
  assign n846 = n845 ^ n841 ;
  assign n847 = n846 ^ n844 ;
  assign n848 = x0 & ~n847 ;
  assign n849 = n848 ^ x0 ;
  assign n850 = x3 & x6 ;
  assign n851 = n850 ^ x3 ;
  assign n852 = x2 & n851 ;
  assign n853 = n215 & n287 ;
  assign n854 = ~n852 & ~n853 ;
  assign n855 = x9 & ~n854 ;
  assign n856 = ~x9 & n215 ;
  assign n857 = ~n851 & ~n856 ;
  assign n858 = ~x8 & ~n857 ;
  assign n859 = ~n855 & ~n858 ;
  assign n860 = ~x1 & ~n859 ;
  assign n861 = n622 & n856 ;
  assign n862 = x5 & x9 ;
  assign n863 = n862 ^ x5 ;
  assign n864 = n863 ^ x9 ;
  assign n865 = ~n428 & n864 ;
  assign n866 = ~x2 & ~n865 ;
  assign n867 = ~x6 & ~n862 ;
  assign n868 = ~n15 & ~n426 ;
  assign n869 = n867 & ~n868 ;
  assign n870 = ~n866 & ~n869 ;
  assign n871 = x3 & ~n870 ;
  assign n872 = ~n861 & ~n871 ;
  assign n873 = ~n860 & n872 ;
  assign n874 = n849 & n873 ;
  assign n875 = n874 ^ n873 ;
  assign n876 = x4 & n875 ;
  assign n877 = n876 ^ x4 ;
  assign n878 = n877 ^ n875 ;
  assign n902 = x6 & n287 ;
  assign n903 = ~n608 & ~n902 ;
  assign n906 = n903 ^ x1 ;
  assign n884 = n376 ^ n131 ;
  assign n885 = n884 ^ x2 ;
  assign n886 = n884 & n885 ;
  assign n879 = n347 ^ x2 ;
  assign n880 = n132 ^ x2 ;
  assign n881 = n879 & ~n880 ;
  assign n882 = ~n376 & n881 ;
  assign n887 = n886 ^ n882 ;
  assign n888 = n887 ^ n881 ;
  assign n889 = n888 ^ n885 ;
  assign n891 = n886 ^ n881 ;
  assign n890 = n131 ^ x2 ;
  assign n892 = n891 ^ n890 ;
  assign n893 = n889 & ~n892 ;
  assign n894 = n893 ^ n886 ;
  assign n883 = n882 ^ n881 ;
  assign n895 = n894 ^ n883 ;
  assign n896 = n895 ^ n885 ;
  assign n897 = ~x3 & ~n614 ;
  assign n898 = ~n187 & ~n897 ;
  assign n899 = n896 & n898 ;
  assign n900 = n899 ^ n896 ;
  assign n901 = n900 ^ n898 ;
  assign n904 = n903 ^ n901 ;
  assign n905 = n904 ^ n903 ;
  assign n907 = n906 ^ n905 ;
  assign n908 = n905 ^ n903 ;
  assign n909 = ~n907 & ~n908 ;
  assign n910 = n909 ^ n905 ;
  assign n911 = x2 & n215 ;
  assign n912 = ~x4 & ~n911 ;
  assign n913 = ~n910 & n912 ;
  assign n914 = n913 ^ x4 ;
  assign n915 = ~x5 & ~n672 ;
  assign n916 = ~x1 & ~x2 ;
  assign n917 = ~x3 & x4 ;
  assign n918 = n916 & n917 ;
  assign n919 = ~n915 & n918 ;
  assign n920 = ~n342 & n919 ;
  assign n921 = ~n914 & n920 ;
  assign n922 = n921 ^ n914 ;
  assign n923 = n922 ^ n920 ;
  assign n924 = x0 & n923 ;
  assign n925 = n924 ^ x0 ;
  assign n926 = n925 ^ n923 ;
  assign n927 = ~x7 & n926 ;
  assign n928 = n878 & n927 ;
  assign n929 = n928 ^ x7 ;
  assign n930 = ~x4 & n582 ;
  assign n931 = x4 ^ x3 ;
  assign n932 = n330 & n931 ;
  assign n933 = ~n930 & ~n932 ;
  assign n934 = ~x7 & n197 ;
  assign n935 = ~n933 & n934 ;
  assign n936 = x3 & ~x4 ;
  assign n937 = ~n330 & n936 ;
  assign n938 = n330 & n917 ;
  assign n939 = ~n937 & ~n938 ;
  assign n940 = n934 & ~n939 ;
  assign n941 = x4 & n124 ;
  assign n942 = ~n287 & n941 ;
  assign n943 = ~n197 & ~n942 ;
  assign n944 = ~x7 & ~n943 ;
  assign n990 = n421 ^ x0 ;
  assign n991 = n990 ^ x6 ;
  assign n992 = ~n624 & ~n991 ;
  assign n993 = n992 ^ n991 ;
  assign n994 = ~n538 & n659 ;
  assign n995 = n993 & n994 ;
  assign n996 = n995 ^ n659 ;
  assign n997 = x0 & ~x1 ;
  assign n998 = n684 & n997 ;
  assign n999 = n998 ^ x0 ;
  assign n1000 = n28 & n999 ;
  assign n1001 = n1000 ^ n999 ;
  assign n1002 = n996 & n1001 ;
  assign n1003 = n1002 ^ n996 ;
  assign n1004 = n1003 ^ n1001 ;
  assign n1005 = x5 & ~n1004 ;
  assign n1006 = n1005 ^ x5 ;
  assign n1007 = n1006 ^ n1004 ;
  assign n1008 = n202 ^ x2 ;
  assign n1009 = n264 & ~n1008 ;
  assign n1010 = x6 & x8 ;
  assign n1011 = n129 & n1010 ;
  assign n1012 = n1009 & n1011 ;
  assign n1013 = n1012 ^ n1009 ;
  assign n1014 = n1013 ^ n1011 ;
  assign n1015 = x9 & ~n1014 ;
  assign n1016 = n1015 ^ x9 ;
  assign n1017 = ~x0 & ~x8 ;
  assign n1018 = n28 & ~n782 ;
  assign n1019 = ~n1017 & n1018 ;
  assign n1020 = n1016 & n1019 ;
  assign n1021 = n1020 ^ n1016 ;
  assign n1022 = n1021 ^ n1019 ;
  assign n1023 = n1007 & ~n1022 ;
  assign n1024 = n1023 ^ n1022 ;
  assign n1025 = x3 & ~n1024 ;
  assign n1026 = n1025 ^ x3 ;
  assign n980 = n12 & n465 ;
  assign n981 = ~x0 & ~n614 ;
  assign n982 = ~x2 & ~x9 ;
  assign n983 = ~n426 & n982 ;
  assign n984 = ~n981 & n983 ;
  assign n985 = ~n980 & ~n984 ;
  assign n946 = n218 ^ x2 ;
  assign n947 = n946 ^ x5 ;
  assign n948 = n947 ^ x2 ;
  assign n951 = n948 ^ x5 ;
  assign n952 = n951 ^ x9 ;
  assign n953 = n952 ^ x6 ;
  assign n954 = x9 & n953 ;
  assign n955 = n954 ^ x6 ;
  assign n956 = n955 ^ x9 ;
  assign n957 = ~x6 & ~n956 ;
  assign n949 = n948 ^ n60 ;
  assign n950 = n60 & n949 ;
  assign n958 = n957 ^ n950 ;
  assign n959 = n958 ^ n954 ;
  assign n945 = n60 ^ x6 ;
  assign n960 = n959 ^ n945 ;
  assign n962 = n957 ^ x6 ;
  assign n961 = n952 ^ x9 ;
  assign n963 = n962 ^ n961 ;
  assign n964 = ~n960 & n963 ;
  assign n965 = n964 ^ n957 ;
  assign n966 = n965 ^ n955 ;
  assign n967 = n966 ^ n218 ;
  assign n968 = n967 ^ x2 ;
  assign n969 = n968 ^ x5 ;
  assign n970 = n969 ^ n947 ;
  assign n971 = x8 & n970 ;
  assign n972 = n971 ^ x8 ;
  assign n973 = n972 ^ n970 ;
  assign n974 = x9 & n523 ;
  assign n975 = ~n715 & ~n974 ;
  assign n976 = x6 & ~n975 ;
  assign n977 = ~n973 & n976 ;
  assign n978 = n977 ^ n973 ;
  assign n979 = n978 ^ n976 ;
  assign n986 = n985 ^ n979 ;
  assign n987 = x1 & n986 ;
  assign n988 = n987 ^ n986 ;
  assign n989 = n988 ^ n979 ;
  assign n1027 = n1026 ^ n989 ;
  assign n1028 = n989 ^ x7 ;
  assign n1029 = x7 & n1028 ;
  assign n1030 = n1029 ^ x7 ;
  assign n1031 = n1030 ^ n1026 ;
  assign n1032 = ~n1027 & ~n1031 ;
  assign n1033 = n1032 ^ n1029 ;
  assign n1034 = n1033 ^ n1026 ;
  assign n1039 = x6 & n879 ;
  assign n1040 = n1039 ^ x6 ;
  assign n1041 = n1040 ^ n879 ;
  assign n1042 = n1041 ^ x2 ;
  assign n1043 = n1042 ^ x6 ;
  assign n1044 = x2 & ~n1043 ;
  assign n1045 = n1044 ^ x2 ;
  assign n1035 = n58 ^ x9 ;
  assign n1036 = n1035 ^ x5 ;
  assign n1037 = n1036 ^ n131 ;
  assign n1038 = ~n131 & n1037 ;
  assign n1046 = n1045 ^ n1038 ;
  assign n1047 = n1046 ^ n1041 ;
  assign n1048 = n1047 ^ n890 ;
  assign n1050 = n1045 ^ x2 ;
  assign n1049 = n347 ^ x6 ;
  assign n1051 = n1050 ^ n1049 ;
  assign n1052 = ~n1048 & n1051 ;
  assign n1053 = n1052 ^ n1051 ;
  assign n1054 = n1053 ^ n1045 ;
  assign n1055 = n1054 ^ n1042 ;
  assign n1056 = n1055 ^ x1 ;
  assign n1057 = n1056 ^ x5 ;
  assign n1058 = n1057 ^ x9 ;
  assign n1059 = n1058 ^ n1035 ;
  assign n1060 = n1059 ^ x0 ;
  assign n1063 = n864 & n1008 ;
  assign n1061 = ~x0 & x2 ;
  assign n1062 = n864 & n1061 ;
  assign n1064 = n1063 ^ n1062 ;
  assign n1065 = n1064 ^ n1059 ;
  assign n1066 = ~n1060 & ~n1065 ;
  assign n1067 = n1066 ^ n1062 ;
  assign n1068 = n1067 ^ n1059 ;
  assign n1069 = x8 & ~n1068 ;
  assign n1070 = n1069 ^ x8 ;
  assign n1071 = n1070 ^ x8 ;
  assign n1073 = x6 & ~n376 ;
  assign n1074 = ~n499 & n1073 ;
  assign n1075 = n946 ^ n41 ;
  assign n1077 = ~x1 & ~x8 ;
  assign n1076 = x2 & ~n946 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1079 = ~n1075 & n1078 ;
  assign n1080 = n1079 ^ n1076 ;
  assign n1081 = x5 & ~n1080 ;
  assign n1082 = n1081 ^ x5 ;
  assign n1083 = n1074 & n1082 ;
  assign n1084 = n1083 ^ n1074 ;
  assign n1085 = n1084 ^ n1082 ;
  assign n1093 = n1071 & ~n1085 ;
  assign n1094 = n1093 ^ n1085 ;
  assign n1072 = n1071 ^ x7 ;
  assign n1086 = n1085 ^ x7 ;
  assign n1087 = n1085 & ~n1086 ;
  assign n1088 = n1087 ^ x7 ;
  assign n1089 = ~n1072 & ~n1088 ;
  assign n1090 = n1089 ^ n1087 ;
  assign n1091 = n1090 ^ n1071 ;
  assign n1092 = n1091 ^ x7 ;
  assign n1095 = n1094 ^ n1092 ;
  assign n1108 = n43 ^ x9 ;
  assign n1106 = n732 ^ n43 ;
  assign n1109 = n1108 ^ n1106 ;
  assign n1110 = n1108 ^ x7 ;
  assign n1111 = x2 ^ x1 ;
  assign n1112 = n1111 ^ x9 ;
  assign n1113 = n1112 ^ x9 ;
  assign n1114 = n1113 ^ n1109 ;
  assign n1115 = n1110 & ~n1114 ;
  assign n1116 = n1115 ^ x7 ;
  assign n1117 = n1116 ^ n1109 ;
  assign n1118 = ~n1109 & ~n1117 ;
  assign n1119 = n1118 ^ n1115 ;
  assign n1120 = n1119 ^ x7 ;
  assign n1107 = n1106 ^ n43 ;
  assign n1121 = n1120 ^ n1107 ;
  assign n1122 = n1108 ^ n43 ;
  assign n1124 = n1106 ^ x7 ;
  assign n1123 = n1113 ^ n1108 ;
  assign n1125 = n1124 ^ n1123 ;
  assign n1126 = n1122 & ~n1125 ;
  assign n1127 = n1126 ^ n1118 ;
  assign n1128 = n1127 ^ n1115 ;
  assign n1129 = ~n1121 & n1128 ;
  assign n1130 = n1129 ^ x9 ;
  assign n1131 = n1130 ^ n1112 ;
  assign n1132 = x0 & ~n1131 ;
  assign n1133 = n1132 ^ x0 ;
  assign n1134 = n1133 ^ n1131 ;
  assign n1096 = n15 & n523 ;
  assign n1097 = n1096 ^ n684 ;
  assign n1098 = ~x2 & x7 ;
  assign n1099 = n1098 ^ n684 ;
  assign n1100 = ~n1098 & ~n1099 ;
  assign n1101 = n1100 ^ n1098 ;
  assign n1102 = n1101 ^ n1096 ;
  assign n1103 = ~n1097 & n1102 ;
  assign n1104 = n1103 ^ n1100 ;
  assign n1105 = n1104 ^ n1096 ;
  assign n1135 = n1134 ^ n1105 ;
  assign n1136 = n1105 ^ n809 ;
  assign n1137 = ~n809 & n1136 ;
  assign n1138 = n1137 ^ n809 ;
  assign n1139 = n1138 ^ n1134 ;
  assign n1140 = n1135 & n1139 ;
  assign n1141 = n1140 ^ n1137 ;
  assign n1142 = n1141 ^ n1134 ;
  assign n1146 = n1095 & n1142 ;
  assign n1147 = n1146 ^ n1142 ;
  assign n1148 = n1147 ^ n1142 ;
  assign n1149 = n1148 ^ n1095 ;
  assign n1143 = x3 & ~n1142 ;
  assign n1144 = n1095 & n1143 ;
  assign n1145 = n1144 ^ x3 ;
  assign n1150 = n1149 ^ n1145 ;
  assign n1151 = x4 & n1150 ;
  assign n1152 = n1151 ^ n1150 ;
  assign n1153 = n1034 & n1152 ;
  assign n1154 = n1153 ^ n1152 ;
  assign n1155 = n1154 ^ x4 ;
  assign n1156 = n944 & n1155 ;
  assign n1157 = n1156 ^ n944 ;
  assign n1158 = n1157 ^ n944 ;
  assign n1159 = n1158 ^ n1155 ;
  assign n1160 = n376 & n1008 ;
  assign n1161 = x8 & n129 ;
  assign n1162 = x7 & x9 ;
  assign n1163 = n1162 ^ x7 ;
  assign n1164 = n1161 & n1163 ;
  assign n1165 = ~n1160 & ~n1164 ;
  assign n1166 = n201 & n809 ;
  assign n1167 = ~n1165 & n1166 ;
  assign n1362 = n1167 ^ x7 ;
  assign n1168 = ~x5 & ~x7 ;
  assign n1169 = n938 & n1168 ;
  assign n1170 = ~x6 & n1169 ;
  assign n1342 = n1170 ^ x4 ;
  assign n1363 = n1362 ^ n1342 ;
  assign n1171 = n1170 ^ n1167 ;
  assign n1348 = n1171 ^ x4 ;
  assign n1227 = ~n376 & n422 ;
  assign n1228 = n399 ^ n376 ;
  assign n1229 = n1228 ^ n732 ;
  assign n1230 = n732 ^ n376 ;
  assign n1231 = n1229 & ~n1230 ;
  assign n1232 = n1231 ^ n732 ;
  assign n1233 = n245 & ~n1232 ;
  assign n1234 = n1227 & n1233 ;
  assign n1235 = n1234 ^ n1227 ;
  assign n1236 = n1235 ^ n1233 ;
  assign n1237 = x3 & ~n1236 ;
  assign n1238 = n1237 ^ x3 ;
  assign n1239 = ~x9 & ~n399 ;
  assign n1240 = x6 ^ x2 ;
  assign n1241 = n1240 ^ x6 ;
  assign n1198 = x8 ^ x6 ;
  assign n1242 = n1241 ^ n1198 ;
  assign n1243 = n1241 ^ x6 ;
  assign n1244 = n1242 & ~n1243 ;
  assign n1245 = n1244 ^ n1241 ;
  assign n1246 = n1239 & ~n1245 ;
  assign n1189 = n492 ^ x3 ;
  assign n1190 = n1189 ^ x8 ;
  assign n1247 = ~x6 & n1190 ;
  assign n1248 = n715 & ~n1247 ;
  assign n1249 = n1246 & n1248 ;
  assign n1250 = n1249 ^ n1246 ;
  assign n1251 = n1250 ^ n1248 ;
  assign n1252 = n1238 & ~n1251 ;
  assign n1253 = n1252 ^ n1251 ;
  assign n1254 = n1253 ^ x1 ;
  assign n1199 = n1198 ^ n376 ;
  assign n1200 = n1198 ^ x9 ;
  assign n1201 = n376 ^ x0 ;
  assign n1202 = n1201 ^ n49 ;
  assign n1203 = n1202 ^ n49 ;
  assign n1204 = n1200 & n1203 ;
  assign n1205 = n1204 ^ n1198 ;
  assign n1206 = n1199 & n1205 ;
  assign n1207 = n1206 ^ n1205 ;
  assign n1208 = n1207 ^ n1200 ;
  assign n1209 = n1198 & n1202 ;
  assign n1210 = n1209 ^ n1199 ;
  assign n1211 = n1208 & n1210 ;
  assign n1212 = n1211 ^ n1208 ;
  assign n1213 = n1212 ^ n1209 ;
  assign n1214 = n1213 ^ n1198 ;
  assign n1215 = n1214 ^ x8 ;
  assign n1216 = n1215 ^ n1198 ;
  assign n1191 = ~n191 & n1190 ;
  assign n1192 = n1191 ^ n191 ;
  assign n1217 = n1216 ^ n1192 ;
  assign n1218 = n1192 ^ x2 ;
  assign n1219 = x2 & n1218 ;
  assign n1220 = n1219 ^ x2 ;
  assign n1221 = n1220 ^ n1216 ;
  assign n1222 = ~n1217 & ~n1221 ;
  assign n1223 = n1222 ^ n1219 ;
  assign n1224 = n1223 ^ n1216 ;
  assign n1175 = n672 ^ x3 ;
  assign n1176 = n1175 ^ x6 ;
  assign n1179 = n672 ^ x6 ;
  assign n1177 = n672 ^ n523 ;
  assign n1178 = n1177 ^ n672 ;
  assign n1180 = n1179 ^ n1178 ;
  assign n1181 = n1179 ^ n672 ;
  assign n1182 = n1180 & ~n1181 ;
  assign n1183 = n1182 ^ n1179 ;
  assign n1184 = ~n1176 & ~n1183 ;
  assign n1185 = n1184 ^ x6 ;
  assign n1186 = n1185 ^ n672 ;
  assign n1187 = n1186 ^ n672 ;
  assign n1188 = n1187 ^ x2 ;
  assign n1193 = x2 & ~n1192 ;
  assign n1194 = n1193 ^ n1187 ;
  assign n1195 = n1188 & n1194 ;
  assign n1196 = n1195 ^ n1188 ;
  assign n1197 = n1196 ^ n1194 ;
  assign n1225 = n1224 ^ n1197 ;
  assign n1226 = n1225 ^ n1187 ;
  assign n1255 = n1254 ^ n1226 ;
  assign n1256 = x1 & n1255 ;
  assign n1257 = n1256 ^ n1254 ;
  assign n1258 = x3 & ~n467 ;
  assign n1259 = n194 & n1258 ;
  assign n1260 = ~x5 & ~n1259 ;
  assign n1261 = ~n1257 & n1260 ;
  assign n1262 = n1261 ^ x5 ;
  assign n1316 = x2 & ~n684 ;
  assign n1317 = n254 & n1316 ;
  assign n1318 = ~n285 & n376 ;
  assign n1319 = ~x2 & ~n254 ;
  assign n1320 = x5 & ~n1319 ;
  assign n1321 = ~n1318 & n1320 ;
  assign n1322 = ~n1317 & ~n1321 ;
  assign n1325 = n1322 ^ x1 ;
  assign n1265 = n17 & n126 ;
  assign n1266 = n1265 ^ n17 ;
  assign n1267 = n1266 ^ n126 ;
  assign n1268 = x0 & ~n1267 ;
  assign n1269 = n1268 ^ x0 ;
  assign n1270 = n1269 ^ n1267 ;
  assign n1313 = n1270 ^ x8 ;
  assign n1278 = n60 ^ x9 ;
  assign n1279 = n1278 ^ x5 ;
  assign n1280 = n1279 ^ x8 ;
  assign n1281 = n1280 ^ n377 ;
  assign n1282 = n1278 ^ x0 ;
  assign n1283 = n1282 ^ x5 ;
  assign n1284 = n732 & ~n1283 ;
  assign n1285 = n1284 ^ n1280 ;
  assign n1286 = ~n1281 & ~n1285 ;
  assign n1287 = n1286 ^ n1280 ;
  assign n1288 = x3 & n1287 ;
  assign n1289 = n1288 ^ x3 ;
  assign n1290 = n1289 ^ n1287 ;
  assign n1263 = n17 & n982 ;
  assign n1291 = n1290 ^ n1263 ;
  assign n1314 = n1313 ^ n1291 ;
  assign n1264 = n1263 ^ x8 ;
  assign n1297 = n1290 ^ n1264 ;
  assign n1274 = x2 & x5 ;
  assign n1275 = n1274 ^ x5 ;
  assign n1276 = x3 & n1275 ;
  assign n1271 = n1270 ^ n1263 ;
  assign n1272 = n1264 & n1271 ;
  assign n1273 = n1272 ^ n1270 ;
  assign n1277 = n1276 ^ n1273 ;
  assign n1298 = n1297 ^ n1277 ;
  assign n1299 = n1276 ^ x8 ;
  assign n1300 = n1299 ^ n1273 ;
  assign n1301 = n1298 & n1300 ;
  assign n1302 = n1301 ^ n1298 ;
  assign n1292 = n1273 ^ x8 ;
  assign n1293 = n1292 ^ n1291 ;
  assign n1294 = n1277 & n1293 ;
  assign n1295 = n1294 ^ n1277 ;
  assign n1303 = n1302 ^ n1295 ;
  assign n1304 = n1303 ^ n1273 ;
  assign n1305 = n1304 ^ n1297 ;
  assign n1306 = n1295 ^ n1276 ;
  assign n1307 = n1306 ^ n1290 ;
  assign n1308 = n1305 & n1307 ;
  assign n1309 = n1308 ^ n1305 ;
  assign n1310 = n1309 ^ n1307 ;
  assign n1311 = n1310 ^ n1302 ;
  assign n1296 = n1295 ^ n1272 ;
  assign n1312 = n1311 ^ n1296 ;
  assign n1315 = n1314 ^ n1312 ;
  assign n1323 = n1322 ^ n1315 ;
  assign n1324 = n1323 ^ n1322 ;
  assign n1326 = n1325 ^ n1324 ;
  assign n1327 = n1325 ^ n1322 ;
  assign n1328 = ~n1326 & n1327 ;
  assign n1329 = n1328 ^ n1327 ;
  assign n1330 = n1329 ^ n1325 ;
  assign n1331 = x8 & n862 ;
  assign n1332 = n285 & n1331 ;
  assign n1333 = ~x6 & ~n1332 ;
  assign n1334 = n1330 & n1333 ;
  assign n1335 = n1334 ^ x6 ;
  assign n1336 = n1262 & n1335 ;
  assign n1337 = n1336 ^ n1262 ;
  assign n1338 = n1337 ^ n1335 ;
  assign n1339 = n1338 ^ n1262 ;
  assign n1340 = n1339 ^ n1335 ;
  assign n1172 = n1170 ^ x7 ;
  assign n1173 = n1171 & n1172 ;
  assign n1174 = n1173 ^ x7 ;
  assign n1341 = n1340 ^ n1174 ;
  assign n1349 = n1348 ^ n1341 ;
  assign n1350 = n1340 ^ n1167 ;
  assign n1351 = n1350 ^ n1174 ;
  assign n1352 = ~n1349 & ~n1351 ;
  assign n1343 = n1174 ^ n1167 ;
  assign n1344 = n1343 ^ n1342 ;
  assign n1345 = ~n1341 & n1344 ;
  assign n1346 = n1345 ^ n1344 ;
  assign n1353 = n1352 ^ n1346 ;
  assign n1354 = n1353 ^ n1174 ;
  assign n1355 = n1354 ^ n1348 ;
  assign n1356 = n1346 ^ n1340 ;
  assign n1357 = n1356 ^ x4 ;
  assign n1358 = n1355 & ~n1357 ;
  assign n1359 = n1358 ^ n1355 ;
  assign n1360 = n1359 ^ n1352 ;
  assign n1347 = n1346 ^ n1173 ;
  assign n1361 = n1360 ^ n1347 ;
  assign n1364 = n1363 ^ n1361 ;
  assign n1365 = n1364 ^ n1170 ;
  assign n1382 = x3 ^ x1 ;
  assign n1383 = x5 & n1382 ;
  assign n1384 = n1383 ^ x3 ;
  assign n1445 = n1384 ^ x8 ;
  assign n1413 = n830 ^ n58 ;
  assign n1409 = n477 ^ x5 ;
  assign n1411 = n1409 ^ x5 ;
  assign n1410 = n1409 ^ x3 ;
  assign n1412 = n1411 ^ n1410 ;
  assign n1414 = n1413 ^ n1412 ;
  assign n1415 = n1412 ^ n830 ;
  assign n1416 = ~n1414 & n1415 ;
  assign n1417 = n1416 ^ n1412 ;
  assign n1425 = n1415 ^ n1414 ;
  assign n1426 = n1425 ^ n1412 ;
  assign n1418 = n1412 ^ n1410 ;
  assign n1419 = n1418 ^ n1415 ;
  assign n1420 = n1419 ^ n1414 ;
  assign n1421 = n1412 ^ n1409 ;
  assign n1422 = n1421 ^ n1415 ;
  assign n1423 = n1422 ^ n1414 ;
  assign n1424 = n1420 & n1423 ;
  assign n1427 = n1426 ^ n1424 ;
  assign n1428 = ~n1417 & n1427 ;
  assign n1429 = n1428 ^ n1412 ;
  assign n1430 = n1429 ^ n1412 ;
  assign n1431 = x8 & ~n1430 ;
  assign n1432 = n1431 ^ x8 ;
  assign n1433 = ~x5 & ~n524 ;
  assign n1434 = ~n17 & n538 ;
  assign n1435 = ~n1433 & n1434 ;
  assign n1436 = n1432 & n1435 ;
  assign n1437 = n1436 ^ n1432 ;
  assign n1438 = n1437 ^ n1435 ;
  assign n1397 = n1274 ^ x2 ;
  assign n1398 = ~n17 & ~n1397 ;
  assign n1399 = ~n475 & n542 ;
  assign n1400 = n1399 ^ x1 ;
  assign n1401 = n1398 & n1400 ;
  assign n1402 = n1401 ^ n1400 ;
  assign n1403 = ~x0 & x5 ;
  assign n1404 = n475 & ~n1403 ;
  assign n1405 = n543 & n1404 ;
  assign n1406 = n1402 & n1405 ;
  assign n1407 = n1406 ^ n1402 ;
  assign n1408 = n1407 ^ n1405 ;
  assign n1439 = n1438 ^ n1408 ;
  assign n1440 = x9 & ~n1439 ;
  assign n1441 = n1440 ^ x9 ;
  assign n1442 = n1441 ^ n1439 ;
  assign n1443 = n1442 ^ n1408 ;
  assign n1368 = n1275 ^ x9 ;
  assign n1366 = n1275 ^ x3 ;
  assign n1367 = n1366 ^ n1275 ;
  assign n1369 = n1368 ^ n1367 ;
  assign n1370 = n1367 ^ n1275 ;
  assign n1371 = ~n1369 & ~n1370 ;
  assign n1372 = n1371 ^ n1367 ;
  assign n1373 = ~x0 & ~n659 ;
  assign n1374 = ~n1372 & n1373 ;
  assign n1375 = n219 ^ x1 ;
  assign n1376 = n1375 ^ x5 ;
  assign n1377 = n659 & n1376 ;
  assign n1378 = n265 & ~n1377 ;
  assign n1379 = n1374 & n1378 ;
  assign n1380 = n1379 ^ n1374 ;
  assign n1381 = n1380 ^ n1378 ;
  assign n1385 = n1384 ^ n1381 ;
  assign n1387 = ~x2 & n273 ;
  assign n1388 = ~n612 & n1387 ;
  assign n1386 = x8 & n1384 ;
  assign n1389 = n1388 ^ n1386 ;
  assign n1390 = n1386 ^ x8 ;
  assign n1391 = n1390 ^ n1384 ;
  assign n1392 = ~n1389 & n1391 ;
  assign n1393 = n1392 ^ n1388 ;
  assign n1394 = n1393 ^ n1384 ;
  assign n1395 = ~n1385 & ~n1394 ;
  assign n1396 = n1395 ^ n1386 ;
  assign n1444 = n1443 ^ n1396 ;
  assign n1446 = n1445 ^ n1444 ;
  assign n1451 = ~n1384 & n1388 ;
  assign n1452 = ~n1381 & n1451 ;
  assign n1453 = n1452 ^ n1381 ;
  assign n1454 = x8 & ~n1453 ;
  assign n1455 = n1454 ^ x8 ;
  assign n1456 = n1455 ^ n1453 ;
  assign n1447 = n1443 ^ x6 ;
  assign n1448 = x6 & n1447 ;
  assign n1449 = n1448 ^ x6 ;
  assign n1450 = n1449 ^ x6 ;
  assign n1457 = n1456 ^ n1450 ;
  assign n1458 = ~n1446 & n1457 ;
  assign n1459 = n1458 ^ n1446 ;
  assign n1460 = n1459 ^ n1449 ;
  assign n1461 = n1460 ^ n1456 ;
  assign n1462 = ~x6 & ~n264 ;
  assign n1463 = ~n999 & n1462 ;
  assign n1464 = x6 & n16 ;
  assign n1465 = n1464 ^ x6 ;
  assign n1466 = ~n28 & n524 ;
  assign n1467 = n1465 & ~n1466 ;
  assign n1468 = ~x2 & ~n1467 ;
  assign n1469 = n18 & ~n1468 ;
  assign n1470 = ~n1463 & n1469 ;
  assign n1471 = ~n1461 & n1470 ;
  assign n1472 = n1471 ^ n1461 ;
  assign n1473 = n1472 ^ n1470 ;
  assign n1474 = n1473 ^ x7 ;
  assign n1475 = n1111 ^ n376 ;
  assign n1476 = n1475 ^ n695 ;
  assign n1478 = n1476 ^ x9 ;
  assign n1477 = n1476 ^ n1475 ;
  assign n1479 = n1478 ^ n1477 ;
  assign n1486 = n1479 ^ n1478 ;
  assign n1483 = n1111 ^ x0 ;
  assign n1484 = n1483 ^ n376 ;
  assign n1481 = n1476 ^ n376 ;
  assign n1482 = n1481 ^ n1478 ;
  assign n1485 = n1484 ^ n1482 ;
  assign n1487 = n1486 ^ n1485 ;
  assign n1488 = n1482 ^ n1479 ;
  assign n1489 = n1482 ^ n1476 ;
  assign n1490 = ~n1488 & ~n1489 ;
  assign n1491 = n1490 ^ n1478 ;
  assign n1492 = n1491 ^ n1489 ;
  assign n1493 = n1487 & ~n1492 ;
  assign n1494 = n1493 ^ n1490 ;
  assign n1480 = n1479 ^ n1476 ;
  assign n1495 = n1494 ^ n1480 ;
  assign n1496 = n1478 ^ n1476 ;
  assign n1497 = n1496 ^ n1479 ;
  assign n1498 = n1497 ^ n1485 ;
  assign n1499 = ~n1484 & n1498 ;
  assign n1500 = n1499 ^ n1493 ;
  assign n1501 = n1500 ^ n1478 ;
  assign n1502 = n1501 ^ n1488 ;
  assign n1503 = n1495 & ~n1502 ;
  assign n1504 = n1503 ^ n1493 ;
  assign n1505 = n1504 ^ n1478 ;
  assign n1506 = n1505 ^ n1488 ;
  assign n1507 = n1506 ^ n1111 ;
  assign n1508 = n1507 ^ n1111 ;
  assign n1509 = n1508 ^ n1484 ;
  assign n1512 = n588 & ~n1509 ;
  assign n1513 = n1512 ^ n588 ;
  assign n1510 = x7 & n588 ;
  assign n1511 = n1509 & n1510 ;
  assign n1514 = n1513 ^ n1511 ;
  assign n1515 = n1514 ^ n1473 ;
  assign n1516 = ~n1474 & ~n1515 ;
  assign n1517 = n1516 ^ n1515 ;
  assign n1518 = n1517 ^ n1511 ;
  assign n1519 = n1518 ^ n1473 ;
  assign n1520 = ~x4 & ~n1169 ;
  assign n1521 = n1519 & n1520 ;
  assign n1522 = n1521 ^ n1169 ;
  assign n1523 = x3 & ~n189 ;
  assign n1524 = n524 & ~n867 ;
  assign n1525 = n1523 & ~n1524 ;
  assign n1526 = ~n809 & n917 ;
  assign n1527 = ~x2 & ~n1526 ;
  assign n1528 = ~n1525 & n1527 ;
  assign n1529 = n265 & n684 ;
  assign n1530 = ~n915 & n1529 ;
  assign n1531 = ~n1528 & ~n1530 ;
  assign n1532 = ~x1 & ~n1531 ;
  assign n1533 = ~x3 & n864 ;
  assign n1534 = n524 & ~n1523 ;
  assign n1535 = ~n1533 & ~n1534 ;
  assign n1536 = ~x2 & ~n1535 ;
  assign n1537 = n852 & n915 ;
  assign n1538 = ~x6 & ~n1331 ;
  assign n1539 = ~x3 & ~n1538 ;
  assign n1540 = ~n1537 & ~n1539 ;
  assign n1541 = ~n1536 & n1540 ;
  assign n1542 = x1 & ~n1541 ;
  assign n1543 = x1 & n684 ;
  assign n1544 = n1543 ^ n684 ;
  assign n1545 = n782 & n852 ;
  assign n1546 = ~x7 & ~n1545 ;
  assign n1547 = ~n1544 & ~n1546 ;
  assign n1548 = ~x7 & ~n675 ;
  assign n1549 = x0 & ~n1548 ;
  assign n1550 = ~x5 & ~n265 ;
  assign n1551 = x6 & ~n1550 ;
  assign n1552 = x4 & ~n675 ;
  assign n1553 = x7 & ~n265 ;
  assign n1554 = ~n1552 & ~n1553 ;
  assign n1555 = ~n1551 & n1554 ;
  assign n1556 = ~n1549 & n1555 ;
  assign n1557 = ~n1547 & n1556 ;
  assign n1558 = ~n1542 & n1557 ;
  assign n1559 = ~n1532 & n1558 ;
  assign n1560 = ~x7 & n809 ;
  assign n1561 = x8 & ~n14 ;
  assign n1562 = x2 & n936 ;
  assign n1563 = n27 & n1562 ;
  assign n1564 = ~n1561 & n1563 ;
  assign n1565 = ~n938 & ~n1564 ;
  assign n1566 = n1560 & ~n1565 ;
  assign y0 = ~n329 ;
  assign y1 = n601 ;
  assign y2 = n816 ;
  assign y3 = ~n929 ;
  assign y4 = n935 ;
  assign y5 = n940 ;
  assign y6 = n1159 ;
  assign y7 = ~n1365 ;
  assign y8 = ~n1522 ;
  assign y9 = n1559 ;
  assign y10 = n1566 ;
endmodule
