module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 ;
  assign n545 = ~x30 & ~x542 ;
  assign n546 = x30 & x542 ;
  assign n547 = ~n545 & ~n546 ;
  assign n548 = ~x29 & ~x541 ;
  assign n549 = x29 & x541 ;
  assign n550 = ~n548 & ~n549 ;
  assign n551 = n547 & n550 ;
  assign n552 = ~n547 & ~n550 ;
  assign n553 = ~n551 & ~n552 ;
  assign n554 = ~x31 & ~x543 ;
  assign n555 = x31 & x543 ;
  assign n556 = ~n554 & ~n555 ;
  assign n557 = ~n553 & ~n556 ;
  assign n558 = n553 & n556 ;
  assign n559 = ~n557 & ~n558 ;
  assign n560 = ~x25 & ~x537 ;
  assign n561 = x25 & x537 ;
  assign n562 = ~n560 & ~n561 ;
  assign n563 = ~n559 & ~n562 ;
  assign n564 = n559 & n562 ;
  assign n565 = ~n563 & ~n564 ;
  assign n566 = ~x27 & ~x539 ;
  assign n567 = x27 & x539 ;
  assign n568 = ~n566 & ~n567 ;
  assign n569 = ~x26 & ~x538 ;
  assign n570 = x26 & x538 ;
  assign n571 = ~n569 & ~n570 ;
  assign n572 = ~n568 & ~n571 ;
  assign n573 = n568 & n571 ;
  assign n574 = ~n572 & ~n573 ;
  assign n575 = ~x28 & ~x540 ;
  assign n576 = x28 & x540 ;
  assign n577 = ~n575 & ~n576 ;
  assign n578 = ~n574 & ~n577 ;
  assign n579 = n574 & n577 ;
  assign n580 = ~n578 & ~n579 ;
  assign n581 = n565 & ~n580 ;
  assign n582 = ~n563 & ~n581 ;
  assign n583 = ~n551 & ~n558 ;
  assign n584 = ~n582 & n583 ;
  assign n585 = n582 & ~n583 ;
  assign n586 = ~n584 & ~n585 ;
  assign n587 = ~n573 & ~n579 ;
  assign n588 = n586 & n587 ;
  assign n589 = ~n584 & ~n588 ;
  assign n590 = ~n586 & ~n587 ;
  assign n591 = ~n588 & ~n590 ;
  assign n592 = ~n565 & n580 ;
  assign n593 = ~n581 & ~n592 ;
  assign n594 = ~x17 & ~x529 ;
  assign n595 = x17 & x529 ;
  assign n596 = ~n594 & ~n595 ;
  assign n597 = n593 & ~n596 ;
  assign n598 = ~x23 & ~x535 ;
  assign n599 = x23 & x535 ;
  assign n600 = ~n598 & ~n599 ;
  assign n601 = ~x22 & ~x534 ;
  assign n602 = x22 & x534 ;
  assign n603 = ~n601 & ~n602 ;
  assign n604 = ~n600 & ~n603 ;
  assign n605 = n600 & n603 ;
  assign n606 = ~n604 & ~n605 ;
  assign n607 = ~x24 & ~x536 ;
  assign n608 = x24 & x536 ;
  assign n609 = ~n607 & ~n608 ;
  assign n610 = ~n606 & ~n609 ;
  assign n611 = n606 & n609 ;
  assign n612 = ~n610 & ~n611 ;
  assign n613 = ~x18 & ~x530 ;
  assign n614 = x18 & x530 ;
  assign n615 = ~n613 & ~n614 ;
  assign n616 = ~n612 & ~n615 ;
  assign n617 = n612 & n615 ;
  assign n618 = ~n616 & ~n617 ;
  assign n619 = ~x20 & ~x532 ;
  assign n620 = x20 & x532 ;
  assign n621 = ~n619 & ~n620 ;
  assign n622 = ~x19 & ~x531 ;
  assign n623 = x19 & x531 ;
  assign n624 = ~n622 & ~n623 ;
  assign n625 = ~n621 & ~n624 ;
  assign n626 = n621 & n624 ;
  assign n627 = ~n625 & ~n626 ;
  assign n628 = ~x21 & ~x533 ;
  assign n629 = x21 & x533 ;
  assign n630 = ~n628 & ~n629 ;
  assign n631 = ~n627 & ~n630 ;
  assign n632 = n627 & n630 ;
  assign n633 = ~n631 & ~n632 ;
  assign n634 = n618 & ~n633 ;
  assign n635 = ~n618 & n633 ;
  assign n636 = ~n634 & ~n635 ;
  assign n637 = ~n593 & n596 ;
  assign n638 = ~n597 & ~n637 ;
  assign n639 = n636 & n638 ;
  assign n640 = ~n597 & ~n639 ;
  assign n641 = n591 & ~n640 ;
  assign n642 = ~n616 & ~n634 ;
  assign n643 = ~n605 & ~n611 ;
  assign n644 = ~n642 & n643 ;
  assign n645 = n642 & ~n643 ;
  assign n646 = ~n644 & ~n645 ;
  assign n647 = ~n626 & ~n632 ;
  assign n648 = n646 & n647 ;
  assign n649 = ~n646 & ~n647 ;
  assign n650 = ~n648 & ~n649 ;
  assign n651 = ~n591 & n640 ;
  assign n652 = ~n641 & ~n651 ;
  assign n653 = n650 & n652 ;
  assign n654 = ~n641 & ~n653 ;
  assign n655 = ~n589 & ~n654 ;
  assign n656 = n589 & n654 ;
  assign n657 = ~n655 & ~n656 ;
  assign n658 = ~n644 & ~n648 ;
  assign n659 = n657 & ~n658 ;
  assign n660 = ~n655 & ~n659 ;
  assign n661 = ~n657 & n658 ;
  assign n662 = ~n659 & ~n661 ;
  assign n663 = ~n650 & ~n652 ;
  assign n664 = ~n653 & ~n663 ;
  assign n665 = ~n636 & ~n638 ;
  assign n666 = ~n639 & ~n665 ;
  assign n667 = ~x1 & ~x513 ;
  assign n668 = x1 & x513 ;
  assign n669 = ~n667 & ~n668 ;
  assign n670 = n666 & ~n669 ;
  assign n671 = ~x8 & ~x520 ;
  assign n672 = x8 & x520 ;
  assign n673 = ~n671 & ~n672 ;
  assign n674 = ~x7 & ~x519 ;
  assign n675 = x7 & x519 ;
  assign n676 = ~n674 & ~n675 ;
  assign n677 = ~n673 & ~n676 ;
  assign n678 = n673 & n676 ;
  assign n679 = ~n677 & ~n678 ;
  assign n680 = ~x9 & ~x521 ;
  assign n681 = x9 & x521 ;
  assign n682 = ~n680 & ~n681 ;
  assign n683 = ~n679 & ~n682 ;
  assign n684 = n679 & n682 ;
  assign n685 = ~n683 & ~n684 ;
  assign n686 = ~x3 & ~x515 ;
  assign n687 = x3 & x515 ;
  assign n688 = ~n686 & ~n687 ;
  assign n689 = ~n685 & ~n688 ;
  assign n690 = n685 & n688 ;
  assign n691 = ~n689 & ~n690 ;
  assign n692 = ~x5 & ~x517 ;
  assign n693 = x5 & x517 ;
  assign n694 = ~n692 & ~n693 ;
  assign n695 = ~x4 & ~x516 ;
  assign n696 = x4 & x516 ;
  assign n697 = ~n695 & ~n696 ;
  assign n698 = ~n694 & ~n697 ;
  assign n699 = n694 & n697 ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = ~x6 & ~x518 ;
  assign n702 = x6 & x518 ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = ~n700 & ~n703 ;
  assign n705 = n700 & n703 ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = n691 & ~n706 ;
  assign n708 = ~n691 & n706 ;
  assign n709 = ~n707 & ~n708 ;
  assign n710 = ~x15 & ~x527 ;
  assign n711 = x15 & x527 ;
  assign n712 = ~n710 & ~n711 ;
  assign n713 = ~x14 & ~x526 ;
  assign n714 = x14 & x526 ;
  assign n715 = ~n713 & ~n714 ;
  assign n716 = ~n712 & ~n715 ;
  assign n717 = n712 & n715 ;
  assign n718 = ~n716 & ~n717 ;
  assign n719 = ~x16 & ~x528 ;
  assign n720 = x16 & x528 ;
  assign n721 = ~n719 & ~n720 ;
  assign n722 = ~n718 & ~n721 ;
  assign n723 = n718 & n721 ;
  assign n724 = ~n722 & ~n723 ;
  assign n725 = ~x10 & ~x522 ;
  assign n726 = x10 & x522 ;
  assign n727 = ~n725 & ~n726 ;
  assign n728 = ~n724 & ~n727 ;
  assign n729 = n724 & n727 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = ~x12 & ~x524 ;
  assign n732 = x12 & x524 ;
  assign n733 = ~n731 & ~n732 ;
  assign n734 = ~x11 & ~x523 ;
  assign n735 = x11 & x523 ;
  assign n736 = ~n734 & ~n735 ;
  assign n737 = ~n733 & ~n736 ;
  assign n738 = n733 & n736 ;
  assign n739 = ~n737 & ~n738 ;
  assign n740 = ~x13 & ~x525 ;
  assign n741 = x13 & x525 ;
  assign n742 = ~n740 & ~n741 ;
  assign n743 = ~n739 & ~n742 ;
  assign n744 = n739 & n742 ;
  assign n745 = ~n743 & ~n744 ;
  assign n746 = n730 & ~n745 ;
  assign n747 = ~n730 & n745 ;
  assign n748 = ~n746 & ~n747 ;
  assign n749 = ~x2 & ~x514 ;
  assign n750 = x2 & x514 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = n748 & ~n751 ;
  assign n753 = ~n748 & n751 ;
  assign n754 = ~n752 & ~n753 ;
  assign n755 = n709 & n754 ;
  assign n756 = ~n709 & ~n754 ;
  assign n757 = ~n755 & ~n756 ;
  assign n758 = ~n666 & n669 ;
  assign n759 = ~n670 & ~n758 ;
  assign n760 = n757 & n759 ;
  assign n761 = ~n670 & ~n760 ;
  assign n762 = n664 & ~n761 ;
  assign n763 = ~n689 & ~n707 ;
  assign n764 = ~n678 & ~n684 ;
  assign n765 = ~n763 & n764 ;
  assign n766 = n763 & ~n764 ;
  assign n767 = ~n765 & ~n766 ;
  assign n768 = ~n699 & ~n705 ;
  assign n769 = n767 & n768 ;
  assign n770 = ~n767 & ~n768 ;
  assign n771 = ~n769 & ~n770 ;
  assign n772 = ~n728 & ~n746 ;
  assign n773 = ~n717 & ~n723 ;
  assign n774 = ~n772 & n773 ;
  assign n775 = n772 & ~n773 ;
  assign n776 = ~n774 & ~n775 ;
  assign n777 = ~n738 & ~n744 ;
  assign n778 = n776 & n777 ;
  assign n779 = ~n776 & ~n777 ;
  assign n780 = ~n778 & ~n779 ;
  assign n781 = ~n752 & ~n755 ;
  assign n782 = n780 & ~n781 ;
  assign n783 = ~n780 & n781 ;
  assign n784 = ~n782 & ~n783 ;
  assign n785 = n771 & n784 ;
  assign n786 = ~n771 & ~n784 ;
  assign n787 = ~n785 & ~n786 ;
  assign n788 = ~n664 & n761 ;
  assign n789 = ~n762 & ~n788 ;
  assign n790 = n787 & n789 ;
  assign n791 = ~n762 & ~n790 ;
  assign n792 = n662 & ~n791 ;
  assign n793 = ~n774 & ~n778 ;
  assign n794 = ~n782 & ~n785 ;
  assign n795 = ~n793 & ~n794 ;
  assign n796 = n793 & n794 ;
  assign n797 = ~n795 & ~n796 ;
  assign n798 = ~n765 & ~n769 ;
  assign n799 = n797 & ~n798 ;
  assign n800 = ~n797 & n798 ;
  assign n801 = ~n799 & ~n800 ;
  assign n802 = ~n662 & n791 ;
  assign n803 = ~n792 & ~n802 ;
  assign n804 = n801 & n803 ;
  assign n805 = ~n792 & ~n804 ;
  assign n806 = ~n660 & ~n805 ;
  assign n807 = n660 & n805 ;
  assign n808 = ~n806 & ~n807 ;
  assign n809 = ~n795 & ~n799 ;
  assign n810 = n808 & ~n809 ;
  assign n811 = ~n808 & n809 ;
  assign n812 = ~n810 & ~n811 ;
  assign n813 = ~n801 & ~n803 ;
  assign n814 = ~n804 & ~n813 ;
  assign n815 = ~n787 & ~n789 ;
  assign n816 = ~n790 & ~n815 ;
  assign n817 = ~n757 & ~n759 ;
  assign n818 = ~n760 & ~n817 ;
  assign n819 = ~x0 & ~x512 ;
  assign n820 = x0 & x512 ;
  assign n821 = ~n819 & ~n820 ;
  assign n822 = ~n818 & n821 ;
  assign n823 = ~n816 & n822 ;
  assign n824 = ~n814 & n823 ;
  assign n825 = ~n812 & n824 ;
  assign n826 = ~n806 & ~n810 ;
  assign n827 = n825 & n826 ;
  assign n828 = ~x510 & ~x542 ;
  assign n829 = x510 & x542 ;
  assign n830 = ~n828 & ~n829 ;
  assign n831 = ~x509 & ~x541 ;
  assign n832 = x509 & x541 ;
  assign n833 = ~n831 & ~n832 ;
  assign n834 = n830 & n833 ;
  assign n835 = ~n830 & ~n833 ;
  assign n836 = ~n834 & ~n835 ;
  assign n837 = ~x511 & ~x543 ;
  assign n838 = x511 & x543 ;
  assign n839 = ~n837 & ~n838 ;
  assign n840 = n836 & n839 ;
  assign n841 = ~n834 & ~n840 ;
  assign n842 = ~n836 & ~n839 ;
  assign n843 = ~n840 & ~n842 ;
  assign n844 = ~x505 & ~x537 ;
  assign n845 = x505 & x537 ;
  assign n846 = ~n844 & ~n845 ;
  assign n847 = n843 & n846 ;
  assign n848 = ~x507 & ~x539 ;
  assign n849 = x507 & x539 ;
  assign n850 = ~n848 & ~n849 ;
  assign n851 = ~x506 & ~x538 ;
  assign n852 = x506 & x538 ;
  assign n853 = ~n851 & ~n852 ;
  assign n854 = ~n850 & ~n853 ;
  assign n855 = n850 & n853 ;
  assign n856 = ~n854 & ~n855 ;
  assign n857 = ~x508 & ~x540 ;
  assign n858 = x508 & x540 ;
  assign n859 = ~n857 & ~n858 ;
  assign n860 = ~n856 & ~n859 ;
  assign n861 = n856 & n859 ;
  assign n862 = ~n860 & ~n861 ;
  assign n863 = ~n843 & ~n846 ;
  assign n864 = ~n847 & ~n863 ;
  assign n865 = n862 & n864 ;
  assign n866 = ~n847 & ~n865 ;
  assign n867 = n841 & n866 ;
  assign n868 = ~n841 & ~n866 ;
  assign n869 = ~n867 & ~n868 ;
  assign n870 = ~n855 & ~n861 ;
  assign n871 = n869 & n870 ;
  assign n872 = ~n867 & ~n871 ;
  assign n873 = ~n869 & ~n870 ;
  assign n874 = ~n871 & ~n873 ;
  assign n875 = ~n862 & ~n864 ;
  assign n876 = ~n865 & ~n875 ;
  assign n877 = ~x497 & ~x529 ;
  assign n878 = x497 & x529 ;
  assign n879 = ~n877 & ~n878 ;
  assign n880 = n876 & n879 ;
  assign n881 = ~x503 & ~x535 ;
  assign n882 = x503 & x535 ;
  assign n883 = ~n881 & ~n882 ;
  assign n884 = ~x502 & ~x534 ;
  assign n885 = x502 & x534 ;
  assign n886 = ~n884 & ~n885 ;
  assign n887 = ~n883 & ~n886 ;
  assign n888 = n883 & n886 ;
  assign n889 = ~n887 & ~n888 ;
  assign n890 = ~x504 & ~x536 ;
  assign n891 = x504 & x536 ;
  assign n892 = ~n890 & ~n891 ;
  assign n893 = ~n889 & ~n892 ;
  assign n894 = n889 & n892 ;
  assign n895 = ~n893 & ~n894 ;
  assign n896 = ~x498 & ~x530 ;
  assign n897 = x498 & x530 ;
  assign n898 = ~n896 & ~n897 ;
  assign n899 = ~n895 & ~n898 ;
  assign n900 = n895 & n898 ;
  assign n901 = ~n899 & ~n900 ;
  assign n902 = ~x500 & ~x532 ;
  assign n903 = x500 & x532 ;
  assign n904 = ~n902 & ~n903 ;
  assign n905 = ~x499 & ~x531 ;
  assign n906 = x499 & x531 ;
  assign n907 = ~n905 & ~n906 ;
  assign n908 = ~n904 & ~n907 ;
  assign n909 = n904 & n907 ;
  assign n910 = ~n908 & ~n909 ;
  assign n911 = ~x501 & ~x533 ;
  assign n912 = x501 & x533 ;
  assign n913 = ~n911 & ~n912 ;
  assign n914 = ~n910 & ~n913 ;
  assign n915 = n910 & n913 ;
  assign n916 = ~n914 & ~n915 ;
  assign n917 = n901 & ~n916 ;
  assign n918 = ~n901 & n916 ;
  assign n919 = ~n917 & ~n918 ;
  assign n920 = ~n876 & ~n879 ;
  assign n921 = ~n880 & ~n920 ;
  assign n922 = ~n919 & n921 ;
  assign n923 = ~n880 & ~n922 ;
  assign n924 = n874 & n923 ;
  assign n925 = ~n874 & ~n923 ;
  assign n926 = ~n899 & ~n917 ;
  assign n927 = ~n888 & ~n894 ;
  assign n928 = ~n926 & n927 ;
  assign n929 = n926 & ~n927 ;
  assign n930 = ~n928 & ~n929 ;
  assign n931 = ~n909 & ~n915 ;
  assign n932 = n930 & n931 ;
  assign n933 = ~n930 & ~n931 ;
  assign n934 = ~n932 & ~n933 ;
  assign n935 = ~n925 & n934 ;
  assign n936 = ~n924 & ~n935 ;
  assign n937 = ~n872 & ~n936 ;
  assign n938 = n872 & n936 ;
  assign n939 = ~n937 & ~n938 ;
  assign n940 = ~n928 & ~n932 ;
  assign n941 = n939 & ~n940 ;
  assign n942 = ~n937 & ~n941 ;
  assign n943 = ~n939 & n940 ;
  assign n944 = ~n941 & ~n943 ;
  assign n945 = n919 & ~n921 ;
  assign n946 = ~n922 & ~n945 ;
  assign n947 = ~x481 & ~x513 ;
  assign n948 = x481 & x513 ;
  assign n949 = ~n947 & ~n948 ;
  assign n950 = n946 & n949 ;
  assign n951 = ~x488 & ~x520 ;
  assign n952 = x488 & x520 ;
  assign n953 = ~n951 & ~n952 ;
  assign n954 = ~x487 & ~x519 ;
  assign n955 = x487 & x519 ;
  assign n956 = ~n954 & ~n955 ;
  assign n957 = ~n953 & ~n956 ;
  assign n958 = n953 & n956 ;
  assign n959 = ~n957 & ~n958 ;
  assign n960 = ~x489 & ~x521 ;
  assign n961 = x489 & x521 ;
  assign n962 = ~n960 & ~n961 ;
  assign n963 = ~n959 & ~n962 ;
  assign n964 = n959 & n962 ;
  assign n965 = ~n963 & ~n964 ;
  assign n966 = ~x483 & ~x515 ;
  assign n967 = x483 & x515 ;
  assign n968 = ~n966 & ~n967 ;
  assign n969 = ~n965 & ~n968 ;
  assign n970 = n965 & n968 ;
  assign n971 = ~n969 & ~n970 ;
  assign n972 = ~x485 & ~x517 ;
  assign n973 = x485 & x517 ;
  assign n974 = ~n972 & ~n973 ;
  assign n975 = ~x484 & ~x516 ;
  assign n976 = x484 & x516 ;
  assign n977 = ~n975 & ~n976 ;
  assign n978 = ~n974 & ~n977 ;
  assign n979 = n974 & n977 ;
  assign n980 = ~n978 & ~n979 ;
  assign n981 = ~x486 & ~x518 ;
  assign n982 = x486 & x518 ;
  assign n983 = ~n981 & ~n982 ;
  assign n984 = ~n980 & ~n983 ;
  assign n985 = n980 & n983 ;
  assign n986 = ~n984 & ~n985 ;
  assign n987 = n971 & ~n986 ;
  assign n988 = ~n971 & n986 ;
  assign n989 = ~n987 & ~n988 ;
  assign n990 = ~x495 & ~x527 ;
  assign n991 = x495 & x527 ;
  assign n992 = ~n990 & ~n991 ;
  assign n993 = ~x494 & ~x526 ;
  assign n994 = x494 & x526 ;
  assign n995 = ~n993 & ~n994 ;
  assign n996 = ~n992 & ~n995 ;
  assign n997 = n992 & n995 ;
  assign n998 = ~n996 & ~n997 ;
  assign n999 = ~x496 & ~x528 ;
  assign n1000 = x496 & x528 ;
  assign n1001 = ~n999 & ~n1000 ;
  assign n1002 = ~n998 & ~n1001 ;
  assign n1003 = n998 & n1001 ;
  assign n1004 = ~n1002 & ~n1003 ;
  assign n1005 = ~x490 & ~x522 ;
  assign n1006 = x490 & x522 ;
  assign n1007 = ~n1005 & ~n1006 ;
  assign n1008 = ~n1004 & ~n1007 ;
  assign n1009 = n1004 & n1007 ;
  assign n1010 = ~n1008 & ~n1009 ;
  assign n1011 = ~x492 & ~x524 ;
  assign n1012 = x492 & x524 ;
  assign n1013 = ~n1011 & ~n1012 ;
  assign n1014 = ~x491 & ~x523 ;
  assign n1015 = x491 & x523 ;
  assign n1016 = ~n1014 & ~n1015 ;
  assign n1017 = ~n1013 & ~n1016 ;
  assign n1018 = n1013 & n1016 ;
  assign n1019 = ~n1017 & ~n1018 ;
  assign n1020 = ~x493 & ~x525 ;
  assign n1021 = x493 & x525 ;
  assign n1022 = ~n1020 & ~n1021 ;
  assign n1023 = ~n1019 & ~n1022 ;
  assign n1024 = n1019 & n1022 ;
  assign n1025 = ~n1023 & ~n1024 ;
  assign n1026 = n1010 & ~n1025 ;
  assign n1027 = ~n1010 & n1025 ;
  assign n1028 = ~n1026 & ~n1027 ;
  assign n1029 = ~x482 & ~x514 ;
  assign n1030 = x482 & x514 ;
  assign n1031 = ~n1029 & ~n1030 ;
  assign n1032 = n1028 & ~n1031 ;
  assign n1033 = ~n1028 & n1031 ;
  assign n1034 = ~n1032 & ~n1033 ;
  assign n1035 = n989 & n1034 ;
  assign n1036 = ~n989 & ~n1034 ;
  assign n1037 = ~n1035 & ~n1036 ;
  assign n1038 = ~n946 & ~n949 ;
  assign n1039 = ~n950 & ~n1038 ;
  assign n1040 = ~n1037 & n1039 ;
  assign n1041 = ~n950 & ~n1040 ;
  assign n1042 = ~n924 & ~n925 ;
  assign n1043 = n934 & n1042 ;
  assign n1044 = ~n934 & ~n1042 ;
  assign n1045 = ~n1043 & ~n1044 ;
  assign n1046 = ~n1041 & ~n1045 ;
  assign n1047 = n1041 & n1045 ;
  assign n1048 = ~n969 & ~n987 ;
  assign n1049 = ~n958 & ~n964 ;
  assign n1050 = ~n1048 & n1049 ;
  assign n1051 = n1048 & ~n1049 ;
  assign n1052 = ~n1050 & ~n1051 ;
  assign n1053 = ~n979 & ~n985 ;
  assign n1054 = n1052 & n1053 ;
  assign n1055 = ~n1052 & ~n1053 ;
  assign n1056 = ~n1054 & ~n1055 ;
  assign n1057 = ~n1008 & ~n1026 ;
  assign n1058 = ~n997 & ~n1003 ;
  assign n1059 = ~n1057 & n1058 ;
  assign n1060 = n1057 & ~n1058 ;
  assign n1061 = ~n1059 & ~n1060 ;
  assign n1062 = ~n1018 & ~n1024 ;
  assign n1063 = n1061 & n1062 ;
  assign n1064 = ~n1061 & ~n1062 ;
  assign n1065 = ~n1063 & ~n1064 ;
  assign n1066 = ~n1032 & ~n1035 ;
  assign n1067 = n1065 & ~n1066 ;
  assign n1068 = ~n1065 & n1066 ;
  assign n1069 = ~n1067 & ~n1068 ;
  assign n1070 = n1056 & ~n1069 ;
  assign n1071 = ~n1056 & n1069 ;
  assign n1072 = ~n1070 & ~n1071 ;
  assign n1073 = ~n1047 & n1072 ;
  assign n1074 = ~n1046 & ~n1073 ;
  assign n1075 = ~n944 & ~n1074 ;
  assign n1076 = n944 & n1074 ;
  assign n1077 = ~n1059 & ~n1063 ;
  assign n1078 = ~n1068 & ~n1071 ;
  assign n1079 = ~n1077 & n1078 ;
  assign n1080 = n1077 & ~n1078 ;
  assign n1081 = ~n1079 & ~n1080 ;
  assign n1082 = ~n1050 & ~n1054 ;
  assign n1083 = n1081 & ~n1082 ;
  assign n1084 = ~n1081 & n1082 ;
  assign n1085 = ~n1083 & ~n1084 ;
  assign n1086 = ~n1076 & ~n1085 ;
  assign n1087 = ~n1075 & ~n1086 ;
  assign n1088 = ~n942 & n1087 ;
  assign n1089 = n942 & ~n1087 ;
  assign n1090 = ~n1088 & ~n1089 ;
  assign n1091 = ~n1079 & ~n1083 ;
  assign n1092 = n1090 & ~n1091 ;
  assign n1093 = ~n1088 & ~n1092 ;
  assign n1094 = ~n1090 & n1091 ;
  assign n1095 = ~n1092 & ~n1094 ;
  assign n1096 = n1037 & ~n1039 ;
  assign n1097 = ~n1040 & ~n1096 ;
  assign n1098 = ~x480 & ~x512 ;
  assign n1099 = x480 & x512 ;
  assign n1100 = ~n1098 & ~n1099 ;
  assign n1101 = n1097 & n1100 ;
  assign n1102 = ~n1046 & ~n1047 ;
  assign n1103 = n1072 & n1102 ;
  assign n1104 = ~n1072 & ~n1102 ;
  assign n1105 = ~n1103 & ~n1104 ;
  assign n1106 = n1101 & n1105 ;
  assign n1107 = ~n1075 & ~n1076 ;
  assign n1108 = ~n1085 & n1107 ;
  assign n1109 = n1085 & ~n1107 ;
  assign n1110 = ~n1108 & ~n1109 ;
  assign n1111 = n1106 & n1110 ;
  assign n1112 = ~n1095 & n1111 ;
  assign n1113 = n1093 & n1112 ;
  assign n1114 = ~x478 & ~x542 ;
  assign n1115 = x478 & x542 ;
  assign n1116 = ~n1114 & ~n1115 ;
  assign n1117 = ~x477 & ~x541 ;
  assign n1118 = x477 & x541 ;
  assign n1119 = ~n1117 & ~n1118 ;
  assign n1120 = n1116 & n1119 ;
  assign n1121 = ~n1116 & ~n1119 ;
  assign n1122 = ~n1120 & ~n1121 ;
  assign n1123 = ~x479 & ~x543 ;
  assign n1124 = x479 & x543 ;
  assign n1125 = ~n1123 & ~n1124 ;
  assign n1126 = n1122 & n1125 ;
  assign n1127 = ~n1120 & ~n1126 ;
  assign n1128 = ~n1122 & ~n1125 ;
  assign n1129 = ~n1126 & ~n1128 ;
  assign n1130 = ~x473 & ~x537 ;
  assign n1131 = x473 & x537 ;
  assign n1132 = ~n1130 & ~n1131 ;
  assign n1133 = n1129 & n1132 ;
  assign n1134 = ~n1129 & ~n1132 ;
  assign n1135 = ~x475 & ~x539 ;
  assign n1136 = x475 & x539 ;
  assign n1137 = ~n1135 & ~n1136 ;
  assign n1138 = ~x474 & ~x538 ;
  assign n1139 = x474 & x538 ;
  assign n1140 = ~n1138 & ~n1139 ;
  assign n1141 = ~n1137 & ~n1140 ;
  assign n1142 = n1137 & n1140 ;
  assign n1143 = ~n1141 & ~n1142 ;
  assign n1144 = ~x476 & ~x540 ;
  assign n1145 = x476 & x540 ;
  assign n1146 = ~n1144 & ~n1145 ;
  assign n1147 = ~n1143 & ~n1146 ;
  assign n1148 = n1143 & n1146 ;
  assign n1149 = ~n1147 & ~n1148 ;
  assign n1150 = ~n1134 & n1149 ;
  assign n1151 = ~n1133 & ~n1150 ;
  assign n1152 = n1127 & n1151 ;
  assign n1153 = ~n1127 & ~n1151 ;
  assign n1154 = ~n1152 & ~n1153 ;
  assign n1155 = ~n1142 & ~n1148 ;
  assign n1156 = n1154 & n1155 ;
  assign n1157 = ~n1152 & ~n1156 ;
  assign n1158 = ~n1154 & ~n1155 ;
  assign n1159 = ~n1156 & ~n1158 ;
  assign n1160 = ~n1133 & ~n1134 ;
  assign n1161 = ~n1149 & n1160 ;
  assign n1162 = n1149 & ~n1160 ;
  assign n1163 = ~n1161 & ~n1162 ;
  assign n1164 = ~x465 & ~x529 ;
  assign n1165 = x465 & x529 ;
  assign n1166 = ~n1164 & ~n1165 ;
  assign n1167 = ~n1163 & n1166 ;
  assign n1168 = n1163 & ~n1166 ;
  assign n1169 = ~x471 & ~x535 ;
  assign n1170 = x471 & x535 ;
  assign n1171 = ~n1169 & ~n1170 ;
  assign n1172 = ~x470 & ~x534 ;
  assign n1173 = x470 & x534 ;
  assign n1174 = ~n1172 & ~n1173 ;
  assign n1175 = ~n1171 & ~n1174 ;
  assign n1176 = n1171 & n1174 ;
  assign n1177 = ~n1175 & ~n1176 ;
  assign n1178 = ~x472 & ~x536 ;
  assign n1179 = x472 & x536 ;
  assign n1180 = ~n1178 & ~n1179 ;
  assign n1181 = ~n1177 & ~n1180 ;
  assign n1182 = n1177 & n1180 ;
  assign n1183 = ~n1181 & ~n1182 ;
  assign n1184 = ~x466 & ~x530 ;
  assign n1185 = x466 & x530 ;
  assign n1186 = ~n1184 & ~n1185 ;
  assign n1187 = ~n1183 & ~n1186 ;
  assign n1188 = n1183 & n1186 ;
  assign n1189 = ~n1187 & ~n1188 ;
  assign n1190 = ~x468 & ~x532 ;
  assign n1191 = x468 & x532 ;
  assign n1192 = ~n1190 & ~n1191 ;
  assign n1193 = ~x467 & ~x531 ;
  assign n1194 = x467 & x531 ;
  assign n1195 = ~n1193 & ~n1194 ;
  assign n1196 = ~n1192 & ~n1195 ;
  assign n1197 = n1192 & n1195 ;
  assign n1198 = ~n1196 & ~n1197 ;
  assign n1199 = ~x469 & ~x533 ;
  assign n1200 = x469 & x533 ;
  assign n1201 = ~n1199 & ~n1200 ;
  assign n1202 = ~n1198 & ~n1201 ;
  assign n1203 = n1198 & n1201 ;
  assign n1204 = ~n1202 & ~n1203 ;
  assign n1205 = n1189 & ~n1204 ;
  assign n1206 = ~n1189 & n1204 ;
  assign n1207 = ~n1205 & ~n1206 ;
  assign n1208 = ~n1168 & ~n1207 ;
  assign n1209 = ~n1167 & ~n1208 ;
  assign n1210 = n1159 & n1209 ;
  assign n1211 = ~n1159 & ~n1209 ;
  assign n1212 = ~n1187 & ~n1205 ;
  assign n1213 = ~n1176 & ~n1182 ;
  assign n1214 = ~n1212 & n1213 ;
  assign n1215 = n1212 & ~n1213 ;
  assign n1216 = ~n1214 & ~n1215 ;
  assign n1217 = ~n1197 & ~n1203 ;
  assign n1218 = n1216 & n1217 ;
  assign n1219 = ~n1216 & ~n1217 ;
  assign n1220 = ~n1218 & ~n1219 ;
  assign n1221 = ~n1211 & n1220 ;
  assign n1222 = ~n1210 & ~n1221 ;
  assign n1223 = ~n1157 & ~n1222 ;
  assign n1224 = n1157 & n1222 ;
  assign n1225 = ~n1223 & ~n1224 ;
  assign n1226 = ~n1214 & ~n1218 ;
  assign n1227 = n1225 & ~n1226 ;
  assign n1228 = ~n1223 & ~n1227 ;
  assign n1229 = ~n1225 & n1226 ;
  assign n1230 = ~n1227 & ~n1229 ;
  assign n1231 = ~x449 & ~x513 ;
  assign n1232 = x449 & x513 ;
  assign n1233 = ~n1231 & ~n1232 ;
  assign n1234 = ~n1167 & ~n1168 ;
  assign n1235 = ~n1207 & n1234 ;
  assign n1236 = n1207 & ~n1234 ;
  assign n1237 = ~n1235 & ~n1236 ;
  assign n1238 = ~n1233 & ~n1237 ;
  assign n1239 = n1233 & n1237 ;
  assign n1240 = ~x456 & ~x520 ;
  assign n1241 = x456 & x520 ;
  assign n1242 = ~n1240 & ~n1241 ;
  assign n1243 = ~x455 & ~x519 ;
  assign n1244 = x455 & x519 ;
  assign n1245 = ~n1243 & ~n1244 ;
  assign n1246 = ~n1242 & ~n1245 ;
  assign n1247 = n1242 & n1245 ;
  assign n1248 = ~n1246 & ~n1247 ;
  assign n1249 = ~x457 & ~x521 ;
  assign n1250 = x457 & x521 ;
  assign n1251 = ~n1249 & ~n1250 ;
  assign n1252 = ~n1248 & ~n1251 ;
  assign n1253 = n1248 & n1251 ;
  assign n1254 = ~n1252 & ~n1253 ;
  assign n1255 = ~x451 & ~x515 ;
  assign n1256 = x451 & x515 ;
  assign n1257 = ~n1255 & ~n1256 ;
  assign n1258 = ~n1254 & ~n1257 ;
  assign n1259 = n1254 & n1257 ;
  assign n1260 = ~n1258 & ~n1259 ;
  assign n1261 = ~x453 & ~x517 ;
  assign n1262 = x453 & x517 ;
  assign n1263 = ~n1261 & ~n1262 ;
  assign n1264 = ~x452 & ~x516 ;
  assign n1265 = x452 & x516 ;
  assign n1266 = ~n1264 & ~n1265 ;
  assign n1267 = ~n1263 & ~n1266 ;
  assign n1268 = n1263 & n1266 ;
  assign n1269 = ~n1267 & ~n1268 ;
  assign n1270 = ~x454 & ~x518 ;
  assign n1271 = x454 & x518 ;
  assign n1272 = ~n1270 & ~n1271 ;
  assign n1273 = ~n1269 & ~n1272 ;
  assign n1274 = n1269 & n1272 ;
  assign n1275 = ~n1273 & ~n1274 ;
  assign n1276 = n1260 & ~n1275 ;
  assign n1277 = ~n1260 & n1275 ;
  assign n1278 = ~n1276 & ~n1277 ;
  assign n1279 = ~x463 & ~x527 ;
  assign n1280 = x463 & x527 ;
  assign n1281 = ~n1279 & ~n1280 ;
  assign n1282 = ~x462 & ~x526 ;
  assign n1283 = x462 & x526 ;
  assign n1284 = ~n1282 & ~n1283 ;
  assign n1285 = ~n1281 & ~n1284 ;
  assign n1286 = n1281 & n1284 ;
  assign n1287 = ~n1285 & ~n1286 ;
  assign n1288 = ~x464 & ~x528 ;
  assign n1289 = x464 & x528 ;
  assign n1290 = ~n1288 & ~n1289 ;
  assign n1291 = ~n1287 & ~n1290 ;
  assign n1292 = n1287 & n1290 ;
  assign n1293 = ~n1291 & ~n1292 ;
  assign n1294 = ~x458 & ~x522 ;
  assign n1295 = x458 & x522 ;
  assign n1296 = ~n1294 & ~n1295 ;
  assign n1297 = ~n1293 & ~n1296 ;
  assign n1298 = n1293 & n1296 ;
  assign n1299 = ~n1297 & ~n1298 ;
  assign n1300 = ~x460 & ~x524 ;
  assign n1301 = x460 & x524 ;
  assign n1302 = ~n1300 & ~n1301 ;
  assign n1303 = ~x459 & ~x523 ;
  assign n1304 = x459 & x523 ;
  assign n1305 = ~n1303 & ~n1304 ;
  assign n1306 = ~n1302 & ~n1305 ;
  assign n1307 = n1302 & n1305 ;
  assign n1308 = ~n1306 & ~n1307 ;
  assign n1309 = ~x461 & ~x525 ;
  assign n1310 = x461 & x525 ;
  assign n1311 = ~n1309 & ~n1310 ;
  assign n1312 = ~n1308 & ~n1311 ;
  assign n1313 = n1308 & n1311 ;
  assign n1314 = ~n1312 & ~n1313 ;
  assign n1315 = n1299 & ~n1314 ;
  assign n1316 = ~n1299 & n1314 ;
  assign n1317 = ~n1315 & ~n1316 ;
  assign n1318 = ~x450 & ~x514 ;
  assign n1319 = x450 & x514 ;
  assign n1320 = ~n1318 & ~n1319 ;
  assign n1321 = n1317 & ~n1320 ;
  assign n1322 = ~n1317 & n1320 ;
  assign n1323 = ~n1321 & ~n1322 ;
  assign n1324 = n1278 & n1323 ;
  assign n1325 = ~n1278 & ~n1323 ;
  assign n1326 = ~n1324 & ~n1325 ;
  assign n1327 = ~n1239 & n1326 ;
  assign n1328 = ~n1238 & ~n1327 ;
  assign n1329 = ~n1210 & ~n1211 ;
  assign n1330 = ~n1220 & n1329 ;
  assign n1331 = n1220 & ~n1329 ;
  assign n1332 = ~n1330 & ~n1331 ;
  assign n1333 = n1328 & n1332 ;
  assign n1334 = ~n1328 & ~n1332 ;
  assign n1335 = ~n1258 & ~n1276 ;
  assign n1336 = ~n1247 & ~n1253 ;
  assign n1337 = ~n1335 & n1336 ;
  assign n1338 = n1335 & ~n1336 ;
  assign n1339 = ~n1337 & ~n1338 ;
  assign n1340 = ~n1268 & ~n1274 ;
  assign n1341 = n1339 & n1340 ;
  assign n1342 = ~n1339 & ~n1340 ;
  assign n1343 = ~n1341 & ~n1342 ;
  assign n1344 = ~n1297 & ~n1315 ;
  assign n1345 = ~n1286 & ~n1292 ;
  assign n1346 = ~n1344 & n1345 ;
  assign n1347 = n1344 & ~n1345 ;
  assign n1348 = ~n1346 & ~n1347 ;
  assign n1349 = ~n1307 & ~n1313 ;
  assign n1350 = n1348 & n1349 ;
  assign n1351 = ~n1348 & ~n1349 ;
  assign n1352 = ~n1350 & ~n1351 ;
  assign n1353 = ~n1321 & ~n1324 ;
  assign n1354 = n1352 & ~n1353 ;
  assign n1355 = ~n1352 & n1353 ;
  assign n1356 = ~n1354 & ~n1355 ;
  assign n1357 = n1343 & n1356 ;
  assign n1358 = ~n1343 & ~n1356 ;
  assign n1359 = ~n1357 & ~n1358 ;
  assign n1360 = ~n1334 & ~n1359 ;
  assign n1361 = ~n1333 & ~n1360 ;
  assign n1362 = ~n1230 & ~n1361 ;
  assign n1363 = n1230 & n1361 ;
  assign n1364 = ~n1343 & ~n1354 ;
  assign n1365 = ~n1355 & ~n1364 ;
  assign n1366 = ~n1346 & ~n1350 ;
  assign n1367 = n1365 & ~n1366 ;
  assign n1368 = ~n1365 & n1366 ;
  assign n1369 = ~n1367 & ~n1368 ;
  assign n1370 = ~n1337 & ~n1341 ;
  assign n1371 = n1369 & ~n1370 ;
  assign n1372 = ~n1369 & n1370 ;
  assign n1373 = ~n1371 & ~n1372 ;
  assign n1374 = ~n1363 & ~n1373 ;
  assign n1375 = ~n1362 & ~n1374 ;
  assign n1376 = ~n1228 & n1375 ;
  assign n1377 = n1228 & ~n1375 ;
  assign n1378 = ~n1376 & ~n1377 ;
  assign n1379 = ~n1367 & ~n1371 ;
  assign n1380 = n1378 & ~n1379 ;
  assign n1381 = ~n1376 & ~n1380 ;
  assign n1382 = ~n1378 & n1379 ;
  assign n1383 = ~n1380 & ~n1382 ;
  assign n1384 = ~x448 & ~x512 ;
  assign n1385 = x448 & x512 ;
  assign n1386 = ~n1384 & ~n1385 ;
  assign n1387 = ~n1238 & ~n1239 ;
  assign n1388 = n1326 & n1387 ;
  assign n1389 = ~n1326 & ~n1387 ;
  assign n1390 = ~n1388 & ~n1389 ;
  assign n1391 = n1386 & ~n1390 ;
  assign n1392 = ~n1333 & ~n1334 ;
  assign n1393 = ~n1359 & n1392 ;
  assign n1394 = n1359 & ~n1392 ;
  assign n1395 = ~n1393 & ~n1394 ;
  assign n1396 = n1391 & n1395 ;
  assign n1397 = ~n1362 & ~n1363 ;
  assign n1398 = ~n1373 & n1397 ;
  assign n1399 = n1373 & ~n1397 ;
  assign n1400 = ~n1398 & ~n1399 ;
  assign n1401 = n1396 & n1400 ;
  assign n1402 = ~n1383 & n1401 ;
  assign n1403 = n1381 & n1402 ;
  assign n1404 = n1113 & n1403 ;
  assign n1405 = ~x446 & ~x542 ;
  assign n1406 = x446 & x542 ;
  assign n1407 = ~n1405 & ~n1406 ;
  assign n1408 = ~x445 & ~x541 ;
  assign n1409 = x445 & x541 ;
  assign n1410 = ~n1408 & ~n1409 ;
  assign n1411 = n1407 & n1410 ;
  assign n1412 = ~n1407 & ~n1410 ;
  assign n1413 = ~n1411 & ~n1412 ;
  assign n1414 = ~x447 & ~x543 ;
  assign n1415 = x447 & x543 ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = ~n1413 & ~n1416 ;
  assign n1418 = n1413 & n1416 ;
  assign n1419 = ~n1417 & ~n1418 ;
  assign n1420 = ~x441 & ~x537 ;
  assign n1421 = x441 & x537 ;
  assign n1422 = ~n1420 & ~n1421 ;
  assign n1423 = ~n1419 & ~n1422 ;
  assign n1424 = n1419 & n1422 ;
  assign n1425 = ~n1423 & ~n1424 ;
  assign n1426 = ~x443 & ~x539 ;
  assign n1427 = x443 & x539 ;
  assign n1428 = ~n1426 & ~n1427 ;
  assign n1429 = ~x442 & ~x538 ;
  assign n1430 = x442 & x538 ;
  assign n1431 = ~n1429 & ~n1430 ;
  assign n1432 = ~n1428 & ~n1431 ;
  assign n1433 = n1428 & n1431 ;
  assign n1434 = ~n1432 & ~n1433 ;
  assign n1435 = ~x444 & ~x540 ;
  assign n1436 = x444 & x540 ;
  assign n1437 = ~n1435 & ~n1436 ;
  assign n1438 = ~n1434 & ~n1437 ;
  assign n1439 = n1434 & n1437 ;
  assign n1440 = ~n1438 & ~n1439 ;
  assign n1441 = n1425 & ~n1440 ;
  assign n1442 = ~n1423 & ~n1441 ;
  assign n1443 = ~n1411 & ~n1418 ;
  assign n1444 = ~n1442 & n1443 ;
  assign n1445 = n1442 & ~n1443 ;
  assign n1446 = ~n1444 & ~n1445 ;
  assign n1447 = ~n1433 & ~n1439 ;
  assign n1448 = n1446 & n1447 ;
  assign n1449 = ~n1444 & ~n1448 ;
  assign n1450 = ~n1446 & ~n1447 ;
  assign n1451 = ~n1448 & ~n1450 ;
  assign n1452 = ~n1425 & n1440 ;
  assign n1453 = ~n1441 & ~n1452 ;
  assign n1454 = ~x433 & ~x529 ;
  assign n1455 = x433 & x529 ;
  assign n1456 = ~n1454 & ~n1455 ;
  assign n1457 = n1453 & ~n1456 ;
  assign n1458 = ~x439 & ~x535 ;
  assign n1459 = x439 & x535 ;
  assign n1460 = ~n1458 & ~n1459 ;
  assign n1461 = ~x438 & ~x534 ;
  assign n1462 = x438 & x534 ;
  assign n1463 = ~n1461 & ~n1462 ;
  assign n1464 = ~n1460 & ~n1463 ;
  assign n1465 = n1460 & n1463 ;
  assign n1466 = ~n1464 & ~n1465 ;
  assign n1467 = ~x440 & ~x536 ;
  assign n1468 = x440 & x536 ;
  assign n1469 = ~n1467 & ~n1468 ;
  assign n1470 = ~n1466 & ~n1469 ;
  assign n1471 = n1466 & n1469 ;
  assign n1472 = ~n1470 & ~n1471 ;
  assign n1473 = ~x434 & ~x530 ;
  assign n1474 = x434 & x530 ;
  assign n1475 = ~n1473 & ~n1474 ;
  assign n1476 = ~n1472 & ~n1475 ;
  assign n1477 = n1472 & n1475 ;
  assign n1478 = ~n1476 & ~n1477 ;
  assign n1479 = ~x436 & ~x532 ;
  assign n1480 = x436 & x532 ;
  assign n1481 = ~n1479 & ~n1480 ;
  assign n1482 = ~x435 & ~x531 ;
  assign n1483 = x435 & x531 ;
  assign n1484 = ~n1482 & ~n1483 ;
  assign n1485 = ~n1481 & ~n1484 ;
  assign n1486 = n1481 & n1484 ;
  assign n1487 = ~n1485 & ~n1486 ;
  assign n1488 = ~x437 & ~x533 ;
  assign n1489 = x437 & x533 ;
  assign n1490 = ~n1488 & ~n1489 ;
  assign n1491 = ~n1487 & ~n1490 ;
  assign n1492 = n1487 & n1490 ;
  assign n1493 = ~n1491 & ~n1492 ;
  assign n1494 = n1478 & ~n1493 ;
  assign n1495 = ~n1478 & n1493 ;
  assign n1496 = ~n1494 & ~n1495 ;
  assign n1497 = ~n1453 & n1456 ;
  assign n1498 = ~n1457 & ~n1497 ;
  assign n1499 = n1496 & n1498 ;
  assign n1500 = ~n1457 & ~n1499 ;
  assign n1501 = n1451 & ~n1500 ;
  assign n1502 = ~n1476 & ~n1494 ;
  assign n1503 = ~n1465 & ~n1471 ;
  assign n1504 = ~n1502 & n1503 ;
  assign n1505 = n1502 & ~n1503 ;
  assign n1506 = ~n1504 & ~n1505 ;
  assign n1507 = ~n1486 & ~n1492 ;
  assign n1508 = n1506 & n1507 ;
  assign n1509 = ~n1506 & ~n1507 ;
  assign n1510 = ~n1508 & ~n1509 ;
  assign n1511 = ~n1451 & n1500 ;
  assign n1512 = ~n1501 & ~n1511 ;
  assign n1513 = n1510 & n1512 ;
  assign n1514 = ~n1501 & ~n1513 ;
  assign n1515 = ~n1449 & ~n1514 ;
  assign n1516 = n1449 & n1514 ;
  assign n1517 = ~n1515 & ~n1516 ;
  assign n1518 = ~n1504 & ~n1508 ;
  assign n1519 = n1517 & ~n1518 ;
  assign n1520 = ~n1515 & ~n1519 ;
  assign n1521 = ~n1517 & n1518 ;
  assign n1522 = ~n1519 & ~n1521 ;
  assign n1523 = ~n1510 & ~n1512 ;
  assign n1524 = ~n1513 & ~n1523 ;
  assign n1525 = ~n1496 & ~n1498 ;
  assign n1526 = ~n1499 & ~n1525 ;
  assign n1527 = ~x417 & ~x513 ;
  assign n1528 = x417 & x513 ;
  assign n1529 = ~n1527 & ~n1528 ;
  assign n1530 = n1526 & ~n1529 ;
  assign n1531 = ~x424 & ~x520 ;
  assign n1532 = x424 & x520 ;
  assign n1533 = ~n1531 & ~n1532 ;
  assign n1534 = ~x423 & ~x519 ;
  assign n1535 = x423 & x519 ;
  assign n1536 = ~n1534 & ~n1535 ;
  assign n1537 = ~n1533 & ~n1536 ;
  assign n1538 = n1533 & n1536 ;
  assign n1539 = ~n1537 & ~n1538 ;
  assign n1540 = ~x425 & ~x521 ;
  assign n1541 = x425 & x521 ;
  assign n1542 = ~n1540 & ~n1541 ;
  assign n1543 = ~n1539 & ~n1542 ;
  assign n1544 = n1539 & n1542 ;
  assign n1545 = ~n1543 & ~n1544 ;
  assign n1546 = ~x419 & ~x515 ;
  assign n1547 = x419 & x515 ;
  assign n1548 = ~n1546 & ~n1547 ;
  assign n1549 = ~n1545 & ~n1548 ;
  assign n1550 = n1545 & n1548 ;
  assign n1551 = ~n1549 & ~n1550 ;
  assign n1552 = ~x421 & ~x517 ;
  assign n1553 = x421 & x517 ;
  assign n1554 = ~n1552 & ~n1553 ;
  assign n1555 = ~x420 & ~x516 ;
  assign n1556 = x420 & x516 ;
  assign n1557 = ~n1555 & ~n1556 ;
  assign n1558 = ~n1554 & ~n1557 ;
  assign n1559 = n1554 & n1557 ;
  assign n1560 = ~n1558 & ~n1559 ;
  assign n1561 = ~x422 & ~x518 ;
  assign n1562 = x422 & x518 ;
  assign n1563 = ~n1561 & ~n1562 ;
  assign n1564 = ~n1560 & ~n1563 ;
  assign n1565 = n1560 & n1563 ;
  assign n1566 = ~n1564 & ~n1565 ;
  assign n1567 = n1551 & ~n1566 ;
  assign n1568 = ~n1551 & n1566 ;
  assign n1569 = ~n1567 & ~n1568 ;
  assign n1570 = ~x431 & ~x527 ;
  assign n1571 = x431 & x527 ;
  assign n1572 = ~n1570 & ~n1571 ;
  assign n1573 = ~x430 & ~x526 ;
  assign n1574 = x430 & x526 ;
  assign n1575 = ~n1573 & ~n1574 ;
  assign n1576 = ~n1572 & ~n1575 ;
  assign n1577 = n1572 & n1575 ;
  assign n1578 = ~n1576 & ~n1577 ;
  assign n1579 = ~x432 & ~x528 ;
  assign n1580 = x432 & x528 ;
  assign n1581 = ~n1579 & ~n1580 ;
  assign n1582 = ~n1578 & ~n1581 ;
  assign n1583 = n1578 & n1581 ;
  assign n1584 = ~n1582 & ~n1583 ;
  assign n1585 = ~x426 & ~x522 ;
  assign n1586 = x426 & x522 ;
  assign n1587 = ~n1585 & ~n1586 ;
  assign n1588 = ~n1584 & ~n1587 ;
  assign n1589 = n1584 & n1587 ;
  assign n1590 = ~n1588 & ~n1589 ;
  assign n1591 = ~x428 & ~x524 ;
  assign n1592 = x428 & x524 ;
  assign n1593 = ~n1591 & ~n1592 ;
  assign n1594 = ~x427 & ~x523 ;
  assign n1595 = x427 & x523 ;
  assign n1596 = ~n1594 & ~n1595 ;
  assign n1597 = ~n1593 & ~n1596 ;
  assign n1598 = n1593 & n1596 ;
  assign n1599 = ~n1597 & ~n1598 ;
  assign n1600 = ~x429 & ~x525 ;
  assign n1601 = x429 & x525 ;
  assign n1602 = ~n1600 & ~n1601 ;
  assign n1603 = ~n1599 & ~n1602 ;
  assign n1604 = n1599 & n1602 ;
  assign n1605 = ~n1603 & ~n1604 ;
  assign n1606 = n1590 & ~n1605 ;
  assign n1607 = ~n1590 & n1605 ;
  assign n1608 = ~n1606 & ~n1607 ;
  assign n1609 = ~x418 & ~x514 ;
  assign n1610 = x418 & x514 ;
  assign n1611 = ~n1609 & ~n1610 ;
  assign n1612 = n1608 & ~n1611 ;
  assign n1613 = ~n1608 & n1611 ;
  assign n1614 = ~n1612 & ~n1613 ;
  assign n1615 = n1569 & n1614 ;
  assign n1616 = ~n1569 & ~n1614 ;
  assign n1617 = ~n1615 & ~n1616 ;
  assign n1618 = ~n1526 & n1529 ;
  assign n1619 = ~n1530 & ~n1618 ;
  assign n1620 = n1617 & n1619 ;
  assign n1621 = ~n1530 & ~n1620 ;
  assign n1622 = n1524 & ~n1621 ;
  assign n1623 = ~n1549 & ~n1567 ;
  assign n1624 = ~n1538 & ~n1544 ;
  assign n1625 = ~n1623 & n1624 ;
  assign n1626 = n1623 & ~n1624 ;
  assign n1627 = ~n1625 & ~n1626 ;
  assign n1628 = ~n1559 & ~n1565 ;
  assign n1629 = n1627 & n1628 ;
  assign n1630 = ~n1627 & ~n1628 ;
  assign n1631 = ~n1629 & ~n1630 ;
  assign n1632 = ~n1588 & ~n1606 ;
  assign n1633 = ~n1577 & ~n1583 ;
  assign n1634 = ~n1632 & n1633 ;
  assign n1635 = n1632 & ~n1633 ;
  assign n1636 = ~n1634 & ~n1635 ;
  assign n1637 = ~n1598 & ~n1604 ;
  assign n1638 = n1636 & n1637 ;
  assign n1639 = ~n1636 & ~n1637 ;
  assign n1640 = ~n1638 & ~n1639 ;
  assign n1641 = ~n1612 & ~n1615 ;
  assign n1642 = n1640 & ~n1641 ;
  assign n1643 = ~n1640 & n1641 ;
  assign n1644 = ~n1642 & ~n1643 ;
  assign n1645 = n1631 & n1644 ;
  assign n1646 = ~n1631 & ~n1644 ;
  assign n1647 = ~n1645 & ~n1646 ;
  assign n1648 = ~n1524 & n1621 ;
  assign n1649 = ~n1622 & ~n1648 ;
  assign n1650 = n1647 & n1649 ;
  assign n1651 = ~n1622 & ~n1650 ;
  assign n1652 = n1522 & ~n1651 ;
  assign n1653 = ~n1634 & ~n1638 ;
  assign n1654 = ~n1642 & ~n1645 ;
  assign n1655 = ~n1653 & ~n1654 ;
  assign n1656 = n1653 & n1654 ;
  assign n1657 = ~n1655 & ~n1656 ;
  assign n1658 = ~n1625 & ~n1629 ;
  assign n1659 = n1657 & ~n1658 ;
  assign n1660 = ~n1657 & n1658 ;
  assign n1661 = ~n1659 & ~n1660 ;
  assign n1662 = ~n1522 & n1651 ;
  assign n1663 = ~n1652 & ~n1662 ;
  assign n1664 = n1661 & n1663 ;
  assign n1665 = ~n1652 & ~n1664 ;
  assign n1666 = ~n1520 & ~n1665 ;
  assign n1667 = n1520 & n1665 ;
  assign n1668 = ~n1666 & ~n1667 ;
  assign n1669 = ~n1655 & ~n1659 ;
  assign n1670 = n1668 & ~n1669 ;
  assign n1671 = ~n1666 & ~n1670 ;
  assign n1672 = ~n1668 & n1669 ;
  assign n1673 = ~n1670 & ~n1672 ;
  assign n1674 = ~n1661 & ~n1663 ;
  assign n1675 = ~n1664 & ~n1674 ;
  assign n1676 = ~n1647 & ~n1649 ;
  assign n1677 = ~n1650 & ~n1676 ;
  assign n1678 = ~n1617 & ~n1619 ;
  assign n1679 = ~n1620 & ~n1678 ;
  assign n1680 = ~x416 & ~x512 ;
  assign n1681 = x416 & x512 ;
  assign n1682 = ~n1680 & ~n1681 ;
  assign n1683 = ~n1679 & n1682 ;
  assign n1684 = ~n1677 & n1683 ;
  assign n1685 = ~n1675 & n1684 ;
  assign n1686 = ~n1673 & n1685 ;
  assign n1687 = n1671 & n1686 ;
  assign n1688 = n1404 & n1687 ;
  assign n1689 = ~x414 & ~x542 ;
  assign n1690 = x414 & x542 ;
  assign n1691 = ~n1689 & ~n1690 ;
  assign n1692 = ~x413 & ~x541 ;
  assign n1693 = x413 & x541 ;
  assign n1694 = ~n1692 & ~n1693 ;
  assign n1695 = n1691 & n1694 ;
  assign n1696 = ~n1691 & ~n1694 ;
  assign n1697 = ~n1695 & ~n1696 ;
  assign n1698 = ~x415 & ~x543 ;
  assign n1699 = x415 & x543 ;
  assign n1700 = ~n1698 & ~n1699 ;
  assign n1701 = ~n1697 & ~n1700 ;
  assign n1702 = n1697 & n1700 ;
  assign n1703 = ~n1701 & ~n1702 ;
  assign n1704 = ~x409 & ~x537 ;
  assign n1705 = x409 & x537 ;
  assign n1706 = ~n1704 & ~n1705 ;
  assign n1707 = ~n1703 & ~n1706 ;
  assign n1708 = n1703 & n1706 ;
  assign n1709 = ~n1707 & ~n1708 ;
  assign n1710 = ~x411 & ~x539 ;
  assign n1711 = x411 & x539 ;
  assign n1712 = ~n1710 & ~n1711 ;
  assign n1713 = ~x410 & ~x538 ;
  assign n1714 = x410 & x538 ;
  assign n1715 = ~n1713 & ~n1714 ;
  assign n1716 = ~n1712 & ~n1715 ;
  assign n1717 = n1712 & n1715 ;
  assign n1718 = ~n1716 & ~n1717 ;
  assign n1719 = ~x412 & ~x540 ;
  assign n1720 = x412 & x540 ;
  assign n1721 = ~n1719 & ~n1720 ;
  assign n1722 = ~n1718 & ~n1721 ;
  assign n1723 = n1718 & n1721 ;
  assign n1724 = ~n1722 & ~n1723 ;
  assign n1725 = n1709 & ~n1724 ;
  assign n1726 = ~n1707 & ~n1725 ;
  assign n1727 = ~n1695 & ~n1702 ;
  assign n1728 = ~n1726 & n1727 ;
  assign n1729 = n1726 & ~n1727 ;
  assign n1730 = ~n1728 & ~n1729 ;
  assign n1731 = ~n1717 & ~n1723 ;
  assign n1732 = n1730 & n1731 ;
  assign n1733 = ~n1728 & ~n1732 ;
  assign n1734 = ~n1730 & ~n1731 ;
  assign n1735 = ~n1732 & ~n1734 ;
  assign n1736 = ~n1709 & n1724 ;
  assign n1737 = ~n1725 & ~n1736 ;
  assign n1738 = ~x401 & ~x529 ;
  assign n1739 = x401 & x529 ;
  assign n1740 = ~n1738 & ~n1739 ;
  assign n1741 = n1737 & ~n1740 ;
  assign n1742 = ~x407 & ~x535 ;
  assign n1743 = x407 & x535 ;
  assign n1744 = ~n1742 & ~n1743 ;
  assign n1745 = ~x406 & ~x534 ;
  assign n1746 = x406 & x534 ;
  assign n1747 = ~n1745 & ~n1746 ;
  assign n1748 = ~n1744 & ~n1747 ;
  assign n1749 = n1744 & n1747 ;
  assign n1750 = ~n1748 & ~n1749 ;
  assign n1751 = ~x408 & ~x536 ;
  assign n1752 = x408 & x536 ;
  assign n1753 = ~n1751 & ~n1752 ;
  assign n1754 = ~n1750 & ~n1753 ;
  assign n1755 = n1750 & n1753 ;
  assign n1756 = ~n1754 & ~n1755 ;
  assign n1757 = ~x402 & ~x530 ;
  assign n1758 = x402 & x530 ;
  assign n1759 = ~n1757 & ~n1758 ;
  assign n1760 = ~n1756 & ~n1759 ;
  assign n1761 = n1756 & n1759 ;
  assign n1762 = ~n1760 & ~n1761 ;
  assign n1763 = ~x404 & ~x532 ;
  assign n1764 = x404 & x532 ;
  assign n1765 = ~n1763 & ~n1764 ;
  assign n1766 = ~x403 & ~x531 ;
  assign n1767 = x403 & x531 ;
  assign n1768 = ~n1766 & ~n1767 ;
  assign n1769 = ~n1765 & ~n1768 ;
  assign n1770 = n1765 & n1768 ;
  assign n1771 = ~n1769 & ~n1770 ;
  assign n1772 = ~x405 & ~x533 ;
  assign n1773 = x405 & x533 ;
  assign n1774 = ~n1772 & ~n1773 ;
  assign n1775 = ~n1771 & ~n1774 ;
  assign n1776 = n1771 & n1774 ;
  assign n1777 = ~n1775 & ~n1776 ;
  assign n1778 = n1762 & ~n1777 ;
  assign n1779 = ~n1762 & n1777 ;
  assign n1780 = ~n1778 & ~n1779 ;
  assign n1781 = ~n1737 & n1740 ;
  assign n1782 = ~n1741 & ~n1781 ;
  assign n1783 = n1780 & n1782 ;
  assign n1784 = ~n1741 & ~n1783 ;
  assign n1785 = n1735 & ~n1784 ;
  assign n1786 = ~n1760 & ~n1778 ;
  assign n1787 = ~n1749 & ~n1755 ;
  assign n1788 = ~n1786 & n1787 ;
  assign n1789 = n1786 & ~n1787 ;
  assign n1790 = ~n1788 & ~n1789 ;
  assign n1791 = ~n1770 & ~n1776 ;
  assign n1792 = n1790 & n1791 ;
  assign n1793 = ~n1790 & ~n1791 ;
  assign n1794 = ~n1792 & ~n1793 ;
  assign n1795 = ~n1735 & n1784 ;
  assign n1796 = ~n1785 & ~n1795 ;
  assign n1797 = n1794 & n1796 ;
  assign n1798 = ~n1785 & ~n1797 ;
  assign n1799 = ~n1733 & ~n1798 ;
  assign n1800 = n1733 & n1798 ;
  assign n1801 = ~n1799 & ~n1800 ;
  assign n1802 = ~n1788 & ~n1792 ;
  assign n1803 = n1801 & ~n1802 ;
  assign n1804 = ~n1799 & ~n1803 ;
  assign n1805 = ~n1801 & n1802 ;
  assign n1806 = ~n1803 & ~n1805 ;
  assign n1807 = ~n1794 & ~n1796 ;
  assign n1808 = ~n1797 & ~n1807 ;
  assign n1809 = ~n1780 & ~n1782 ;
  assign n1810 = ~n1783 & ~n1809 ;
  assign n1811 = ~x385 & ~x513 ;
  assign n1812 = x385 & x513 ;
  assign n1813 = ~n1811 & ~n1812 ;
  assign n1814 = n1810 & ~n1813 ;
  assign n1815 = ~x392 & ~x520 ;
  assign n1816 = x392 & x520 ;
  assign n1817 = ~n1815 & ~n1816 ;
  assign n1818 = ~x391 & ~x519 ;
  assign n1819 = x391 & x519 ;
  assign n1820 = ~n1818 & ~n1819 ;
  assign n1821 = ~n1817 & ~n1820 ;
  assign n1822 = n1817 & n1820 ;
  assign n1823 = ~n1821 & ~n1822 ;
  assign n1824 = ~x393 & ~x521 ;
  assign n1825 = x393 & x521 ;
  assign n1826 = ~n1824 & ~n1825 ;
  assign n1827 = ~n1823 & ~n1826 ;
  assign n1828 = n1823 & n1826 ;
  assign n1829 = ~n1827 & ~n1828 ;
  assign n1830 = ~x387 & ~x515 ;
  assign n1831 = x387 & x515 ;
  assign n1832 = ~n1830 & ~n1831 ;
  assign n1833 = ~n1829 & ~n1832 ;
  assign n1834 = n1829 & n1832 ;
  assign n1835 = ~n1833 & ~n1834 ;
  assign n1836 = ~x389 & ~x517 ;
  assign n1837 = x389 & x517 ;
  assign n1838 = ~n1836 & ~n1837 ;
  assign n1839 = ~x388 & ~x516 ;
  assign n1840 = x388 & x516 ;
  assign n1841 = ~n1839 & ~n1840 ;
  assign n1842 = ~n1838 & ~n1841 ;
  assign n1843 = n1838 & n1841 ;
  assign n1844 = ~n1842 & ~n1843 ;
  assign n1845 = ~x390 & ~x518 ;
  assign n1846 = x390 & x518 ;
  assign n1847 = ~n1845 & ~n1846 ;
  assign n1848 = ~n1844 & ~n1847 ;
  assign n1849 = n1844 & n1847 ;
  assign n1850 = ~n1848 & ~n1849 ;
  assign n1851 = n1835 & ~n1850 ;
  assign n1852 = ~n1835 & n1850 ;
  assign n1853 = ~n1851 & ~n1852 ;
  assign n1854 = ~x399 & ~x527 ;
  assign n1855 = x399 & x527 ;
  assign n1856 = ~n1854 & ~n1855 ;
  assign n1857 = ~x398 & ~x526 ;
  assign n1858 = x398 & x526 ;
  assign n1859 = ~n1857 & ~n1858 ;
  assign n1860 = ~n1856 & ~n1859 ;
  assign n1861 = n1856 & n1859 ;
  assign n1862 = ~n1860 & ~n1861 ;
  assign n1863 = ~x400 & ~x528 ;
  assign n1864 = x400 & x528 ;
  assign n1865 = ~n1863 & ~n1864 ;
  assign n1866 = ~n1862 & ~n1865 ;
  assign n1867 = n1862 & n1865 ;
  assign n1868 = ~n1866 & ~n1867 ;
  assign n1869 = ~x394 & ~x522 ;
  assign n1870 = x394 & x522 ;
  assign n1871 = ~n1869 & ~n1870 ;
  assign n1872 = ~n1868 & ~n1871 ;
  assign n1873 = n1868 & n1871 ;
  assign n1874 = ~n1872 & ~n1873 ;
  assign n1875 = ~x396 & ~x524 ;
  assign n1876 = x396 & x524 ;
  assign n1877 = ~n1875 & ~n1876 ;
  assign n1878 = ~x395 & ~x523 ;
  assign n1879 = x395 & x523 ;
  assign n1880 = ~n1878 & ~n1879 ;
  assign n1881 = ~n1877 & ~n1880 ;
  assign n1882 = n1877 & n1880 ;
  assign n1883 = ~n1881 & ~n1882 ;
  assign n1884 = ~x397 & ~x525 ;
  assign n1885 = x397 & x525 ;
  assign n1886 = ~n1884 & ~n1885 ;
  assign n1887 = ~n1883 & ~n1886 ;
  assign n1888 = n1883 & n1886 ;
  assign n1889 = ~n1887 & ~n1888 ;
  assign n1890 = n1874 & ~n1889 ;
  assign n1891 = ~n1874 & n1889 ;
  assign n1892 = ~n1890 & ~n1891 ;
  assign n1893 = ~x386 & ~x514 ;
  assign n1894 = x386 & x514 ;
  assign n1895 = ~n1893 & ~n1894 ;
  assign n1896 = n1892 & ~n1895 ;
  assign n1897 = ~n1892 & n1895 ;
  assign n1898 = ~n1896 & ~n1897 ;
  assign n1899 = n1853 & n1898 ;
  assign n1900 = ~n1853 & ~n1898 ;
  assign n1901 = ~n1899 & ~n1900 ;
  assign n1902 = ~n1810 & n1813 ;
  assign n1903 = ~n1814 & ~n1902 ;
  assign n1904 = n1901 & n1903 ;
  assign n1905 = ~n1814 & ~n1904 ;
  assign n1906 = n1808 & ~n1905 ;
  assign n1907 = ~n1833 & ~n1851 ;
  assign n1908 = ~n1822 & ~n1828 ;
  assign n1909 = ~n1907 & n1908 ;
  assign n1910 = n1907 & ~n1908 ;
  assign n1911 = ~n1909 & ~n1910 ;
  assign n1912 = ~n1843 & ~n1849 ;
  assign n1913 = n1911 & n1912 ;
  assign n1914 = ~n1911 & ~n1912 ;
  assign n1915 = ~n1913 & ~n1914 ;
  assign n1916 = ~n1872 & ~n1890 ;
  assign n1917 = ~n1861 & ~n1867 ;
  assign n1918 = ~n1916 & n1917 ;
  assign n1919 = n1916 & ~n1917 ;
  assign n1920 = ~n1918 & ~n1919 ;
  assign n1921 = ~n1882 & ~n1888 ;
  assign n1922 = n1920 & n1921 ;
  assign n1923 = ~n1920 & ~n1921 ;
  assign n1924 = ~n1922 & ~n1923 ;
  assign n1925 = ~n1896 & ~n1899 ;
  assign n1926 = n1924 & ~n1925 ;
  assign n1927 = ~n1924 & n1925 ;
  assign n1928 = ~n1926 & ~n1927 ;
  assign n1929 = n1915 & n1928 ;
  assign n1930 = ~n1915 & ~n1928 ;
  assign n1931 = ~n1929 & ~n1930 ;
  assign n1932 = ~n1808 & n1905 ;
  assign n1933 = ~n1906 & ~n1932 ;
  assign n1934 = n1931 & n1933 ;
  assign n1935 = ~n1906 & ~n1934 ;
  assign n1936 = n1806 & ~n1935 ;
  assign n1937 = ~n1918 & ~n1922 ;
  assign n1938 = ~n1926 & ~n1929 ;
  assign n1939 = ~n1937 & ~n1938 ;
  assign n1940 = n1937 & n1938 ;
  assign n1941 = ~n1939 & ~n1940 ;
  assign n1942 = ~n1909 & ~n1913 ;
  assign n1943 = n1941 & ~n1942 ;
  assign n1944 = ~n1941 & n1942 ;
  assign n1945 = ~n1943 & ~n1944 ;
  assign n1946 = ~n1806 & n1935 ;
  assign n1947 = ~n1936 & ~n1946 ;
  assign n1948 = n1945 & n1947 ;
  assign n1949 = ~n1936 & ~n1948 ;
  assign n1950 = ~n1804 & ~n1949 ;
  assign n1951 = n1804 & n1949 ;
  assign n1952 = ~n1950 & ~n1951 ;
  assign n1953 = ~n1939 & ~n1943 ;
  assign n1954 = n1952 & ~n1953 ;
  assign n1955 = ~n1950 & ~n1954 ;
  assign n1956 = ~n1952 & n1953 ;
  assign n1957 = ~n1954 & ~n1956 ;
  assign n1958 = ~n1945 & ~n1947 ;
  assign n1959 = ~n1948 & ~n1958 ;
  assign n1960 = ~n1931 & ~n1933 ;
  assign n1961 = ~n1934 & ~n1960 ;
  assign n1962 = ~n1901 & ~n1903 ;
  assign n1963 = ~n1904 & ~n1962 ;
  assign n1964 = ~x384 & ~x512 ;
  assign n1965 = x384 & x512 ;
  assign n1966 = ~n1964 & ~n1965 ;
  assign n1967 = ~n1963 & n1966 ;
  assign n1968 = ~n1961 & n1967 ;
  assign n1969 = ~n1959 & n1968 ;
  assign n1970 = ~n1957 & n1969 ;
  assign n1971 = n1955 & n1970 ;
  assign n1972 = n1688 & n1971 ;
  assign n1973 = ~x382 & ~x542 ;
  assign n1974 = x382 & x542 ;
  assign n1975 = ~n1973 & ~n1974 ;
  assign n1976 = ~x381 & ~x541 ;
  assign n1977 = x381 & x541 ;
  assign n1978 = ~n1976 & ~n1977 ;
  assign n1979 = n1975 & n1978 ;
  assign n1980 = ~n1975 & ~n1978 ;
  assign n1981 = ~n1979 & ~n1980 ;
  assign n1982 = ~x383 & ~x543 ;
  assign n1983 = x383 & x543 ;
  assign n1984 = ~n1982 & ~n1983 ;
  assign n1985 = ~n1981 & ~n1984 ;
  assign n1986 = n1981 & n1984 ;
  assign n1987 = ~n1985 & ~n1986 ;
  assign n1988 = ~x377 & ~x537 ;
  assign n1989 = x377 & x537 ;
  assign n1990 = ~n1988 & ~n1989 ;
  assign n1991 = ~n1987 & ~n1990 ;
  assign n1992 = n1987 & n1990 ;
  assign n1993 = ~n1991 & ~n1992 ;
  assign n1994 = ~x379 & ~x539 ;
  assign n1995 = x379 & x539 ;
  assign n1996 = ~n1994 & ~n1995 ;
  assign n1997 = ~x378 & ~x538 ;
  assign n1998 = x378 & x538 ;
  assign n1999 = ~n1997 & ~n1998 ;
  assign n2000 = ~n1996 & ~n1999 ;
  assign n2001 = n1996 & n1999 ;
  assign n2002 = ~n2000 & ~n2001 ;
  assign n2003 = ~x380 & ~x540 ;
  assign n2004 = x380 & x540 ;
  assign n2005 = ~n2003 & ~n2004 ;
  assign n2006 = ~n2002 & ~n2005 ;
  assign n2007 = n2002 & n2005 ;
  assign n2008 = ~n2006 & ~n2007 ;
  assign n2009 = n1993 & ~n2008 ;
  assign n2010 = ~n1991 & ~n2009 ;
  assign n2011 = ~n1979 & ~n1986 ;
  assign n2012 = ~n2010 & n2011 ;
  assign n2013 = n2010 & ~n2011 ;
  assign n2014 = ~n2012 & ~n2013 ;
  assign n2015 = ~n2001 & ~n2007 ;
  assign n2016 = n2014 & n2015 ;
  assign n2017 = ~n2012 & ~n2016 ;
  assign n2018 = ~n2014 & ~n2015 ;
  assign n2019 = ~n2016 & ~n2018 ;
  assign n2020 = ~n1993 & n2008 ;
  assign n2021 = ~n2009 & ~n2020 ;
  assign n2022 = ~x369 & ~x529 ;
  assign n2023 = x369 & x529 ;
  assign n2024 = ~n2022 & ~n2023 ;
  assign n2025 = n2021 & ~n2024 ;
  assign n2026 = ~x375 & ~x535 ;
  assign n2027 = x375 & x535 ;
  assign n2028 = ~n2026 & ~n2027 ;
  assign n2029 = ~x374 & ~x534 ;
  assign n2030 = x374 & x534 ;
  assign n2031 = ~n2029 & ~n2030 ;
  assign n2032 = ~n2028 & ~n2031 ;
  assign n2033 = n2028 & n2031 ;
  assign n2034 = ~n2032 & ~n2033 ;
  assign n2035 = ~x376 & ~x536 ;
  assign n2036 = x376 & x536 ;
  assign n2037 = ~n2035 & ~n2036 ;
  assign n2038 = ~n2034 & ~n2037 ;
  assign n2039 = n2034 & n2037 ;
  assign n2040 = ~n2038 & ~n2039 ;
  assign n2041 = ~x370 & ~x530 ;
  assign n2042 = x370 & x530 ;
  assign n2043 = ~n2041 & ~n2042 ;
  assign n2044 = ~n2040 & ~n2043 ;
  assign n2045 = n2040 & n2043 ;
  assign n2046 = ~n2044 & ~n2045 ;
  assign n2047 = ~x372 & ~x532 ;
  assign n2048 = x372 & x532 ;
  assign n2049 = ~n2047 & ~n2048 ;
  assign n2050 = ~x371 & ~x531 ;
  assign n2051 = x371 & x531 ;
  assign n2052 = ~n2050 & ~n2051 ;
  assign n2053 = ~n2049 & ~n2052 ;
  assign n2054 = n2049 & n2052 ;
  assign n2055 = ~n2053 & ~n2054 ;
  assign n2056 = ~x373 & ~x533 ;
  assign n2057 = x373 & x533 ;
  assign n2058 = ~n2056 & ~n2057 ;
  assign n2059 = ~n2055 & ~n2058 ;
  assign n2060 = n2055 & n2058 ;
  assign n2061 = ~n2059 & ~n2060 ;
  assign n2062 = n2046 & ~n2061 ;
  assign n2063 = ~n2046 & n2061 ;
  assign n2064 = ~n2062 & ~n2063 ;
  assign n2065 = ~n2021 & n2024 ;
  assign n2066 = ~n2025 & ~n2065 ;
  assign n2067 = n2064 & n2066 ;
  assign n2068 = ~n2025 & ~n2067 ;
  assign n2069 = n2019 & ~n2068 ;
  assign n2070 = ~n2044 & ~n2062 ;
  assign n2071 = ~n2033 & ~n2039 ;
  assign n2072 = ~n2070 & n2071 ;
  assign n2073 = n2070 & ~n2071 ;
  assign n2074 = ~n2072 & ~n2073 ;
  assign n2075 = ~n2054 & ~n2060 ;
  assign n2076 = n2074 & n2075 ;
  assign n2077 = ~n2074 & ~n2075 ;
  assign n2078 = ~n2076 & ~n2077 ;
  assign n2079 = ~n2019 & n2068 ;
  assign n2080 = ~n2069 & ~n2079 ;
  assign n2081 = n2078 & n2080 ;
  assign n2082 = ~n2069 & ~n2081 ;
  assign n2083 = ~n2017 & ~n2082 ;
  assign n2084 = n2017 & n2082 ;
  assign n2085 = ~n2083 & ~n2084 ;
  assign n2086 = ~n2072 & ~n2076 ;
  assign n2087 = n2085 & ~n2086 ;
  assign n2088 = ~n2083 & ~n2087 ;
  assign n2089 = ~n2085 & n2086 ;
  assign n2090 = ~n2087 & ~n2089 ;
  assign n2091 = ~n2078 & ~n2080 ;
  assign n2092 = ~n2081 & ~n2091 ;
  assign n2093 = ~n2064 & ~n2066 ;
  assign n2094 = ~n2067 & ~n2093 ;
  assign n2095 = ~x353 & ~x513 ;
  assign n2096 = x353 & x513 ;
  assign n2097 = ~n2095 & ~n2096 ;
  assign n2098 = n2094 & ~n2097 ;
  assign n2099 = ~x360 & ~x520 ;
  assign n2100 = x360 & x520 ;
  assign n2101 = ~n2099 & ~n2100 ;
  assign n2102 = ~x359 & ~x519 ;
  assign n2103 = x359 & x519 ;
  assign n2104 = ~n2102 & ~n2103 ;
  assign n2105 = ~n2101 & ~n2104 ;
  assign n2106 = n2101 & n2104 ;
  assign n2107 = ~n2105 & ~n2106 ;
  assign n2108 = ~x361 & ~x521 ;
  assign n2109 = x361 & x521 ;
  assign n2110 = ~n2108 & ~n2109 ;
  assign n2111 = ~n2107 & ~n2110 ;
  assign n2112 = n2107 & n2110 ;
  assign n2113 = ~n2111 & ~n2112 ;
  assign n2114 = ~x355 & ~x515 ;
  assign n2115 = x355 & x515 ;
  assign n2116 = ~n2114 & ~n2115 ;
  assign n2117 = ~n2113 & ~n2116 ;
  assign n2118 = n2113 & n2116 ;
  assign n2119 = ~n2117 & ~n2118 ;
  assign n2120 = ~x357 & ~x517 ;
  assign n2121 = x357 & x517 ;
  assign n2122 = ~n2120 & ~n2121 ;
  assign n2123 = ~x356 & ~x516 ;
  assign n2124 = x356 & x516 ;
  assign n2125 = ~n2123 & ~n2124 ;
  assign n2126 = ~n2122 & ~n2125 ;
  assign n2127 = n2122 & n2125 ;
  assign n2128 = ~n2126 & ~n2127 ;
  assign n2129 = ~x358 & ~x518 ;
  assign n2130 = x358 & x518 ;
  assign n2131 = ~n2129 & ~n2130 ;
  assign n2132 = ~n2128 & ~n2131 ;
  assign n2133 = n2128 & n2131 ;
  assign n2134 = ~n2132 & ~n2133 ;
  assign n2135 = n2119 & ~n2134 ;
  assign n2136 = ~n2119 & n2134 ;
  assign n2137 = ~n2135 & ~n2136 ;
  assign n2138 = ~x367 & ~x527 ;
  assign n2139 = x367 & x527 ;
  assign n2140 = ~n2138 & ~n2139 ;
  assign n2141 = ~x366 & ~x526 ;
  assign n2142 = x366 & x526 ;
  assign n2143 = ~n2141 & ~n2142 ;
  assign n2144 = ~n2140 & ~n2143 ;
  assign n2145 = n2140 & n2143 ;
  assign n2146 = ~n2144 & ~n2145 ;
  assign n2147 = ~x368 & ~x528 ;
  assign n2148 = x368 & x528 ;
  assign n2149 = ~n2147 & ~n2148 ;
  assign n2150 = ~n2146 & ~n2149 ;
  assign n2151 = n2146 & n2149 ;
  assign n2152 = ~n2150 & ~n2151 ;
  assign n2153 = ~x362 & ~x522 ;
  assign n2154 = x362 & x522 ;
  assign n2155 = ~n2153 & ~n2154 ;
  assign n2156 = ~n2152 & ~n2155 ;
  assign n2157 = n2152 & n2155 ;
  assign n2158 = ~n2156 & ~n2157 ;
  assign n2159 = ~x364 & ~x524 ;
  assign n2160 = x364 & x524 ;
  assign n2161 = ~n2159 & ~n2160 ;
  assign n2162 = ~x363 & ~x523 ;
  assign n2163 = x363 & x523 ;
  assign n2164 = ~n2162 & ~n2163 ;
  assign n2165 = ~n2161 & ~n2164 ;
  assign n2166 = n2161 & n2164 ;
  assign n2167 = ~n2165 & ~n2166 ;
  assign n2168 = ~x365 & ~x525 ;
  assign n2169 = x365 & x525 ;
  assign n2170 = ~n2168 & ~n2169 ;
  assign n2171 = ~n2167 & ~n2170 ;
  assign n2172 = n2167 & n2170 ;
  assign n2173 = ~n2171 & ~n2172 ;
  assign n2174 = n2158 & ~n2173 ;
  assign n2175 = ~n2158 & n2173 ;
  assign n2176 = ~n2174 & ~n2175 ;
  assign n2177 = ~x354 & ~x514 ;
  assign n2178 = x354 & x514 ;
  assign n2179 = ~n2177 & ~n2178 ;
  assign n2180 = n2176 & ~n2179 ;
  assign n2181 = ~n2176 & n2179 ;
  assign n2182 = ~n2180 & ~n2181 ;
  assign n2183 = n2137 & n2182 ;
  assign n2184 = ~n2137 & ~n2182 ;
  assign n2185 = ~n2183 & ~n2184 ;
  assign n2186 = ~n2094 & n2097 ;
  assign n2187 = ~n2098 & ~n2186 ;
  assign n2188 = n2185 & n2187 ;
  assign n2189 = ~n2098 & ~n2188 ;
  assign n2190 = n2092 & ~n2189 ;
  assign n2191 = ~n2117 & ~n2135 ;
  assign n2192 = ~n2106 & ~n2112 ;
  assign n2193 = ~n2191 & n2192 ;
  assign n2194 = n2191 & ~n2192 ;
  assign n2195 = ~n2193 & ~n2194 ;
  assign n2196 = ~n2127 & ~n2133 ;
  assign n2197 = n2195 & n2196 ;
  assign n2198 = ~n2195 & ~n2196 ;
  assign n2199 = ~n2197 & ~n2198 ;
  assign n2200 = ~n2156 & ~n2174 ;
  assign n2201 = ~n2145 & ~n2151 ;
  assign n2202 = ~n2200 & n2201 ;
  assign n2203 = n2200 & ~n2201 ;
  assign n2204 = ~n2202 & ~n2203 ;
  assign n2205 = ~n2166 & ~n2172 ;
  assign n2206 = n2204 & n2205 ;
  assign n2207 = ~n2204 & ~n2205 ;
  assign n2208 = ~n2206 & ~n2207 ;
  assign n2209 = ~n2180 & ~n2183 ;
  assign n2210 = n2208 & ~n2209 ;
  assign n2211 = ~n2208 & n2209 ;
  assign n2212 = ~n2210 & ~n2211 ;
  assign n2213 = n2199 & n2212 ;
  assign n2214 = ~n2199 & ~n2212 ;
  assign n2215 = ~n2213 & ~n2214 ;
  assign n2216 = ~n2092 & n2189 ;
  assign n2217 = ~n2190 & ~n2216 ;
  assign n2218 = n2215 & n2217 ;
  assign n2219 = ~n2190 & ~n2218 ;
  assign n2220 = n2090 & ~n2219 ;
  assign n2221 = ~n2202 & ~n2206 ;
  assign n2222 = ~n2210 & ~n2213 ;
  assign n2223 = ~n2221 & ~n2222 ;
  assign n2224 = n2221 & n2222 ;
  assign n2225 = ~n2223 & ~n2224 ;
  assign n2226 = ~n2193 & ~n2197 ;
  assign n2227 = n2225 & ~n2226 ;
  assign n2228 = ~n2225 & n2226 ;
  assign n2229 = ~n2227 & ~n2228 ;
  assign n2230 = ~n2090 & n2219 ;
  assign n2231 = ~n2220 & ~n2230 ;
  assign n2232 = n2229 & n2231 ;
  assign n2233 = ~n2220 & ~n2232 ;
  assign n2234 = ~n2088 & ~n2233 ;
  assign n2235 = n2088 & n2233 ;
  assign n2236 = ~n2234 & ~n2235 ;
  assign n2237 = ~n2223 & ~n2227 ;
  assign n2238 = n2236 & ~n2237 ;
  assign n2239 = ~n2234 & ~n2238 ;
  assign n2240 = ~n2236 & n2237 ;
  assign n2241 = ~n2238 & ~n2240 ;
  assign n2242 = ~n2229 & ~n2231 ;
  assign n2243 = ~n2232 & ~n2242 ;
  assign n2244 = ~n2215 & ~n2217 ;
  assign n2245 = ~n2218 & ~n2244 ;
  assign n2246 = ~n2185 & ~n2187 ;
  assign n2247 = ~n2188 & ~n2246 ;
  assign n2248 = ~x352 & ~x512 ;
  assign n2249 = x352 & x512 ;
  assign n2250 = ~n2248 & ~n2249 ;
  assign n2251 = ~n2247 & n2250 ;
  assign n2252 = ~n2245 & n2251 ;
  assign n2253 = ~n2243 & n2252 ;
  assign n2254 = ~n2241 & n2253 ;
  assign n2255 = n2239 & n2254 ;
  assign n2256 = n1972 & n2255 ;
  assign n2257 = ~x350 & ~x542 ;
  assign n2258 = x350 & x542 ;
  assign n2259 = ~n2257 & ~n2258 ;
  assign n2260 = ~x349 & ~x541 ;
  assign n2261 = x349 & x541 ;
  assign n2262 = ~n2260 & ~n2261 ;
  assign n2263 = n2259 & n2262 ;
  assign n2264 = ~n2259 & ~n2262 ;
  assign n2265 = ~n2263 & ~n2264 ;
  assign n2266 = ~x351 & ~x543 ;
  assign n2267 = x351 & x543 ;
  assign n2268 = ~n2266 & ~n2267 ;
  assign n2269 = ~n2265 & ~n2268 ;
  assign n2270 = n2265 & n2268 ;
  assign n2271 = ~n2269 & ~n2270 ;
  assign n2272 = ~x345 & ~x537 ;
  assign n2273 = x345 & x537 ;
  assign n2274 = ~n2272 & ~n2273 ;
  assign n2275 = ~n2271 & ~n2274 ;
  assign n2276 = n2271 & n2274 ;
  assign n2277 = ~n2275 & ~n2276 ;
  assign n2278 = ~x347 & ~x539 ;
  assign n2279 = x347 & x539 ;
  assign n2280 = ~n2278 & ~n2279 ;
  assign n2281 = ~x346 & ~x538 ;
  assign n2282 = x346 & x538 ;
  assign n2283 = ~n2281 & ~n2282 ;
  assign n2284 = ~n2280 & ~n2283 ;
  assign n2285 = n2280 & n2283 ;
  assign n2286 = ~n2284 & ~n2285 ;
  assign n2287 = ~x348 & ~x540 ;
  assign n2288 = x348 & x540 ;
  assign n2289 = ~n2287 & ~n2288 ;
  assign n2290 = ~n2286 & ~n2289 ;
  assign n2291 = n2286 & n2289 ;
  assign n2292 = ~n2290 & ~n2291 ;
  assign n2293 = n2277 & ~n2292 ;
  assign n2294 = ~n2275 & ~n2293 ;
  assign n2295 = ~n2263 & ~n2270 ;
  assign n2296 = ~n2294 & n2295 ;
  assign n2297 = n2294 & ~n2295 ;
  assign n2298 = ~n2296 & ~n2297 ;
  assign n2299 = ~n2285 & ~n2291 ;
  assign n2300 = n2298 & n2299 ;
  assign n2301 = ~n2296 & ~n2300 ;
  assign n2302 = ~n2298 & ~n2299 ;
  assign n2303 = ~n2300 & ~n2302 ;
  assign n2304 = ~n2277 & n2292 ;
  assign n2305 = ~n2293 & ~n2304 ;
  assign n2306 = ~x337 & ~x529 ;
  assign n2307 = x337 & x529 ;
  assign n2308 = ~n2306 & ~n2307 ;
  assign n2309 = n2305 & ~n2308 ;
  assign n2310 = ~x343 & ~x535 ;
  assign n2311 = x343 & x535 ;
  assign n2312 = ~n2310 & ~n2311 ;
  assign n2313 = ~x342 & ~x534 ;
  assign n2314 = x342 & x534 ;
  assign n2315 = ~n2313 & ~n2314 ;
  assign n2316 = ~n2312 & ~n2315 ;
  assign n2317 = n2312 & n2315 ;
  assign n2318 = ~n2316 & ~n2317 ;
  assign n2319 = ~x344 & ~x536 ;
  assign n2320 = x344 & x536 ;
  assign n2321 = ~n2319 & ~n2320 ;
  assign n2322 = ~n2318 & ~n2321 ;
  assign n2323 = n2318 & n2321 ;
  assign n2324 = ~n2322 & ~n2323 ;
  assign n2325 = ~x338 & ~x530 ;
  assign n2326 = x338 & x530 ;
  assign n2327 = ~n2325 & ~n2326 ;
  assign n2328 = ~n2324 & ~n2327 ;
  assign n2329 = n2324 & n2327 ;
  assign n2330 = ~n2328 & ~n2329 ;
  assign n2331 = ~x340 & ~x532 ;
  assign n2332 = x340 & x532 ;
  assign n2333 = ~n2331 & ~n2332 ;
  assign n2334 = ~x339 & ~x531 ;
  assign n2335 = x339 & x531 ;
  assign n2336 = ~n2334 & ~n2335 ;
  assign n2337 = ~n2333 & ~n2336 ;
  assign n2338 = n2333 & n2336 ;
  assign n2339 = ~n2337 & ~n2338 ;
  assign n2340 = ~x341 & ~x533 ;
  assign n2341 = x341 & x533 ;
  assign n2342 = ~n2340 & ~n2341 ;
  assign n2343 = ~n2339 & ~n2342 ;
  assign n2344 = n2339 & n2342 ;
  assign n2345 = ~n2343 & ~n2344 ;
  assign n2346 = n2330 & ~n2345 ;
  assign n2347 = ~n2330 & n2345 ;
  assign n2348 = ~n2346 & ~n2347 ;
  assign n2349 = ~n2305 & n2308 ;
  assign n2350 = ~n2309 & ~n2349 ;
  assign n2351 = n2348 & n2350 ;
  assign n2352 = ~n2309 & ~n2351 ;
  assign n2353 = n2303 & ~n2352 ;
  assign n2354 = ~n2328 & ~n2346 ;
  assign n2355 = ~n2317 & ~n2323 ;
  assign n2356 = ~n2354 & n2355 ;
  assign n2357 = n2354 & ~n2355 ;
  assign n2358 = ~n2356 & ~n2357 ;
  assign n2359 = ~n2338 & ~n2344 ;
  assign n2360 = n2358 & n2359 ;
  assign n2361 = ~n2358 & ~n2359 ;
  assign n2362 = ~n2360 & ~n2361 ;
  assign n2363 = ~n2303 & n2352 ;
  assign n2364 = ~n2353 & ~n2363 ;
  assign n2365 = n2362 & n2364 ;
  assign n2366 = ~n2353 & ~n2365 ;
  assign n2367 = ~n2301 & ~n2366 ;
  assign n2368 = n2301 & n2366 ;
  assign n2369 = ~n2367 & ~n2368 ;
  assign n2370 = ~n2356 & ~n2360 ;
  assign n2371 = n2369 & ~n2370 ;
  assign n2372 = ~n2367 & ~n2371 ;
  assign n2373 = ~n2369 & n2370 ;
  assign n2374 = ~n2371 & ~n2373 ;
  assign n2375 = ~n2362 & ~n2364 ;
  assign n2376 = ~n2365 & ~n2375 ;
  assign n2377 = ~n2348 & ~n2350 ;
  assign n2378 = ~n2351 & ~n2377 ;
  assign n2379 = ~x321 & ~x513 ;
  assign n2380 = x321 & x513 ;
  assign n2381 = ~n2379 & ~n2380 ;
  assign n2382 = n2378 & ~n2381 ;
  assign n2383 = ~x328 & ~x520 ;
  assign n2384 = x328 & x520 ;
  assign n2385 = ~n2383 & ~n2384 ;
  assign n2386 = ~x327 & ~x519 ;
  assign n2387 = x327 & x519 ;
  assign n2388 = ~n2386 & ~n2387 ;
  assign n2389 = ~n2385 & ~n2388 ;
  assign n2390 = n2385 & n2388 ;
  assign n2391 = ~n2389 & ~n2390 ;
  assign n2392 = ~x329 & ~x521 ;
  assign n2393 = x329 & x521 ;
  assign n2394 = ~n2392 & ~n2393 ;
  assign n2395 = ~n2391 & ~n2394 ;
  assign n2396 = n2391 & n2394 ;
  assign n2397 = ~n2395 & ~n2396 ;
  assign n2398 = ~x323 & ~x515 ;
  assign n2399 = x323 & x515 ;
  assign n2400 = ~n2398 & ~n2399 ;
  assign n2401 = ~n2397 & ~n2400 ;
  assign n2402 = n2397 & n2400 ;
  assign n2403 = ~n2401 & ~n2402 ;
  assign n2404 = ~x325 & ~x517 ;
  assign n2405 = x325 & x517 ;
  assign n2406 = ~n2404 & ~n2405 ;
  assign n2407 = ~x324 & ~x516 ;
  assign n2408 = x324 & x516 ;
  assign n2409 = ~n2407 & ~n2408 ;
  assign n2410 = ~n2406 & ~n2409 ;
  assign n2411 = n2406 & n2409 ;
  assign n2412 = ~n2410 & ~n2411 ;
  assign n2413 = ~x326 & ~x518 ;
  assign n2414 = x326 & x518 ;
  assign n2415 = ~n2413 & ~n2414 ;
  assign n2416 = ~n2412 & ~n2415 ;
  assign n2417 = n2412 & n2415 ;
  assign n2418 = ~n2416 & ~n2417 ;
  assign n2419 = n2403 & ~n2418 ;
  assign n2420 = ~n2403 & n2418 ;
  assign n2421 = ~n2419 & ~n2420 ;
  assign n2422 = ~x335 & ~x527 ;
  assign n2423 = x335 & x527 ;
  assign n2424 = ~n2422 & ~n2423 ;
  assign n2425 = ~x334 & ~x526 ;
  assign n2426 = x334 & x526 ;
  assign n2427 = ~n2425 & ~n2426 ;
  assign n2428 = ~n2424 & ~n2427 ;
  assign n2429 = n2424 & n2427 ;
  assign n2430 = ~n2428 & ~n2429 ;
  assign n2431 = ~x336 & ~x528 ;
  assign n2432 = x336 & x528 ;
  assign n2433 = ~n2431 & ~n2432 ;
  assign n2434 = ~n2430 & ~n2433 ;
  assign n2435 = n2430 & n2433 ;
  assign n2436 = ~n2434 & ~n2435 ;
  assign n2437 = ~x330 & ~x522 ;
  assign n2438 = x330 & x522 ;
  assign n2439 = ~n2437 & ~n2438 ;
  assign n2440 = ~n2436 & ~n2439 ;
  assign n2441 = n2436 & n2439 ;
  assign n2442 = ~n2440 & ~n2441 ;
  assign n2443 = ~x332 & ~x524 ;
  assign n2444 = x332 & x524 ;
  assign n2445 = ~n2443 & ~n2444 ;
  assign n2446 = ~x331 & ~x523 ;
  assign n2447 = x331 & x523 ;
  assign n2448 = ~n2446 & ~n2447 ;
  assign n2449 = ~n2445 & ~n2448 ;
  assign n2450 = n2445 & n2448 ;
  assign n2451 = ~n2449 & ~n2450 ;
  assign n2452 = ~x333 & ~x525 ;
  assign n2453 = x333 & x525 ;
  assign n2454 = ~n2452 & ~n2453 ;
  assign n2455 = ~n2451 & ~n2454 ;
  assign n2456 = n2451 & n2454 ;
  assign n2457 = ~n2455 & ~n2456 ;
  assign n2458 = n2442 & ~n2457 ;
  assign n2459 = ~n2442 & n2457 ;
  assign n2460 = ~n2458 & ~n2459 ;
  assign n2461 = ~x322 & ~x514 ;
  assign n2462 = x322 & x514 ;
  assign n2463 = ~n2461 & ~n2462 ;
  assign n2464 = n2460 & ~n2463 ;
  assign n2465 = ~n2460 & n2463 ;
  assign n2466 = ~n2464 & ~n2465 ;
  assign n2467 = n2421 & n2466 ;
  assign n2468 = ~n2421 & ~n2466 ;
  assign n2469 = ~n2467 & ~n2468 ;
  assign n2470 = ~n2378 & n2381 ;
  assign n2471 = ~n2382 & ~n2470 ;
  assign n2472 = n2469 & n2471 ;
  assign n2473 = ~n2382 & ~n2472 ;
  assign n2474 = n2376 & ~n2473 ;
  assign n2475 = ~n2401 & ~n2419 ;
  assign n2476 = ~n2390 & ~n2396 ;
  assign n2477 = ~n2475 & n2476 ;
  assign n2478 = n2475 & ~n2476 ;
  assign n2479 = ~n2477 & ~n2478 ;
  assign n2480 = ~n2411 & ~n2417 ;
  assign n2481 = n2479 & n2480 ;
  assign n2482 = ~n2479 & ~n2480 ;
  assign n2483 = ~n2481 & ~n2482 ;
  assign n2484 = ~n2440 & ~n2458 ;
  assign n2485 = ~n2429 & ~n2435 ;
  assign n2486 = ~n2484 & n2485 ;
  assign n2487 = n2484 & ~n2485 ;
  assign n2488 = ~n2486 & ~n2487 ;
  assign n2489 = ~n2450 & ~n2456 ;
  assign n2490 = n2488 & n2489 ;
  assign n2491 = ~n2488 & ~n2489 ;
  assign n2492 = ~n2490 & ~n2491 ;
  assign n2493 = ~n2464 & ~n2467 ;
  assign n2494 = n2492 & ~n2493 ;
  assign n2495 = ~n2492 & n2493 ;
  assign n2496 = ~n2494 & ~n2495 ;
  assign n2497 = n2483 & n2496 ;
  assign n2498 = ~n2483 & ~n2496 ;
  assign n2499 = ~n2497 & ~n2498 ;
  assign n2500 = ~n2376 & n2473 ;
  assign n2501 = ~n2474 & ~n2500 ;
  assign n2502 = n2499 & n2501 ;
  assign n2503 = ~n2474 & ~n2502 ;
  assign n2504 = n2374 & ~n2503 ;
  assign n2505 = ~n2486 & ~n2490 ;
  assign n2506 = ~n2494 & ~n2497 ;
  assign n2507 = ~n2505 & ~n2506 ;
  assign n2508 = n2505 & n2506 ;
  assign n2509 = ~n2507 & ~n2508 ;
  assign n2510 = ~n2477 & ~n2481 ;
  assign n2511 = n2509 & ~n2510 ;
  assign n2512 = ~n2509 & n2510 ;
  assign n2513 = ~n2511 & ~n2512 ;
  assign n2514 = ~n2374 & n2503 ;
  assign n2515 = ~n2504 & ~n2514 ;
  assign n2516 = n2513 & n2515 ;
  assign n2517 = ~n2504 & ~n2516 ;
  assign n2518 = ~n2372 & ~n2517 ;
  assign n2519 = n2372 & n2517 ;
  assign n2520 = ~n2518 & ~n2519 ;
  assign n2521 = ~n2507 & ~n2511 ;
  assign n2522 = n2520 & ~n2521 ;
  assign n2523 = ~n2518 & ~n2522 ;
  assign n2524 = ~n2520 & n2521 ;
  assign n2525 = ~n2522 & ~n2524 ;
  assign n2526 = ~n2513 & ~n2515 ;
  assign n2527 = ~n2516 & ~n2526 ;
  assign n2528 = ~n2499 & ~n2501 ;
  assign n2529 = ~n2502 & ~n2528 ;
  assign n2530 = ~n2469 & ~n2471 ;
  assign n2531 = ~n2472 & ~n2530 ;
  assign n2532 = ~x320 & ~x512 ;
  assign n2533 = x320 & x512 ;
  assign n2534 = ~n2532 & ~n2533 ;
  assign n2535 = ~n2531 & n2534 ;
  assign n2536 = ~n2529 & n2535 ;
  assign n2537 = ~n2527 & n2536 ;
  assign n2538 = ~n2525 & n2537 ;
  assign n2539 = n2523 & n2538 ;
  assign n2540 = n2256 & n2539 ;
  assign n2541 = ~x318 & ~x542 ;
  assign n2542 = x318 & x542 ;
  assign n2543 = ~n2541 & ~n2542 ;
  assign n2544 = ~x317 & ~x541 ;
  assign n2545 = x317 & x541 ;
  assign n2546 = ~n2544 & ~n2545 ;
  assign n2547 = n2543 & n2546 ;
  assign n2548 = ~n2543 & ~n2546 ;
  assign n2549 = ~n2547 & ~n2548 ;
  assign n2550 = ~x319 & ~x543 ;
  assign n2551 = x319 & x543 ;
  assign n2552 = ~n2550 & ~n2551 ;
  assign n2553 = ~n2549 & ~n2552 ;
  assign n2554 = n2549 & n2552 ;
  assign n2555 = ~n2553 & ~n2554 ;
  assign n2556 = ~x313 & ~x537 ;
  assign n2557 = x313 & x537 ;
  assign n2558 = ~n2556 & ~n2557 ;
  assign n2559 = ~n2555 & ~n2558 ;
  assign n2560 = n2555 & n2558 ;
  assign n2561 = ~n2559 & ~n2560 ;
  assign n2562 = ~x315 & ~x539 ;
  assign n2563 = x315 & x539 ;
  assign n2564 = ~n2562 & ~n2563 ;
  assign n2565 = ~x314 & ~x538 ;
  assign n2566 = x314 & x538 ;
  assign n2567 = ~n2565 & ~n2566 ;
  assign n2568 = ~n2564 & ~n2567 ;
  assign n2569 = n2564 & n2567 ;
  assign n2570 = ~n2568 & ~n2569 ;
  assign n2571 = ~x316 & ~x540 ;
  assign n2572 = x316 & x540 ;
  assign n2573 = ~n2571 & ~n2572 ;
  assign n2574 = ~n2570 & ~n2573 ;
  assign n2575 = n2570 & n2573 ;
  assign n2576 = ~n2574 & ~n2575 ;
  assign n2577 = n2561 & ~n2576 ;
  assign n2578 = ~n2559 & ~n2577 ;
  assign n2579 = ~n2547 & ~n2554 ;
  assign n2580 = ~n2578 & n2579 ;
  assign n2581 = n2578 & ~n2579 ;
  assign n2582 = ~n2580 & ~n2581 ;
  assign n2583 = ~n2569 & ~n2575 ;
  assign n2584 = n2582 & n2583 ;
  assign n2585 = ~n2580 & ~n2584 ;
  assign n2586 = ~n2582 & ~n2583 ;
  assign n2587 = ~n2584 & ~n2586 ;
  assign n2588 = ~n2561 & n2576 ;
  assign n2589 = ~n2577 & ~n2588 ;
  assign n2590 = ~x305 & ~x529 ;
  assign n2591 = x305 & x529 ;
  assign n2592 = ~n2590 & ~n2591 ;
  assign n2593 = n2589 & ~n2592 ;
  assign n2594 = ~x311 & ~x535 ;
  assign n2595 = x311 & x535 ;
  assign n2596 = ~n2594 & ~n2595 ;
  assign n2597 = ~x310 & ~x534 ;
  assign n2598 = x310 & x534 ;
  assign n2599 = ~n2597 & ~n2598 ;
  assign n2600 = ~n2596 & ~n2599 ;
  assign n2601 = n2596 & n2599 ;
  assign n2602 = ~n2600 & ~n2601 ;
  assign n2603 = ~x312 & ~x536 ;
  assign n2604 = x312 & x536 ;
  assign n2605 = ~n2603 & ~n2604 ;
  assign n2606 = ~n2602 & ~n2605 ;
  assign n2607 = n2602 & n2605 ;
  assign n2608 = ~n2606 & ~n2607 ;
  assign n2609 = ~x306 & ~x530 ;
  assign n2610 = x306 & x530 ;
  assign n2611 = ~n2609 & ~n2610 ;
  assign n2612 = ~n2608 & ~n2611 ;
  assign n2613 = n2608 & n2611 ;
  assign n2614 = ~n2612 & ~n2613 ;
  assign n2615 = ~x308 & ~x532 ;
  assign n2616 = x308 & x532 ;
  assign n2617 = ~n2615 & ~n2616 ;
  assign n2618 = ~x307 & ~x531 ;
  assign n2619 = x307 & x531 ;
  assign n2620 = ~n2618 & ~n2619 ;
  assign n2621 = ~n2617 & ~n2620 ;
  assign n2622 = n2617 & n2620 ;
  assign n2623 = ~n2621 & ~n2622 ;
  assign n2624 = ~x309 & ~x533 ;
  assign n2625 = x309 & x533 ;
  assign n2626 = ~n2624 & ~n2625 ;
  assign n2627 = ~n2623 & ~n2626 ;
  assign n2628 = n2623 & n2626 ;
  assign n2629 = ~n2627 & ~n2628 ;
  assign n2630 = n2614 & ~n2629 ;
  assign n2631 = ~n2614 & n2629 ;
  assign n2632 = ~n2630 & ~n2631 ;
  assign n2633 = ~n2589 & n2592 ;
  assign n2634 = ~n2593 & ~n2633 ;
  assign n2635 = n2632 & n2634 ;
  assign n2636 = ~n2593 & ~n2635 ;
  assign n2637 = n2587 & ~n2636 ;
  assign n2638 = ~n2612 & ~n2630 ;
  assign n2639 = ~n2601 & ~n2607 ;
  assign n2640 = ~n2638 & n2639 ;
  assign n2641 = n2638 & ~n2639 ;
  assign n2642 = ~n2640 & ~n2641 ;
  assign n2643 = ~n2622 & ~n2628 ;
  assign n2644 = n2642 & n2643 ;
  assign n2645 = ~n2642 & ~n2643 ;
  assign n2646 = ~n2644 & ~n2645 ;
  assign n2647 = ~n2587 & n2636 ;
  assign n2648 = ~n2637 & ~n2647 ;
  assign n2649 = n2646 & n2648 ;
  assign n2650 = ~n2637 & ~n2649 ;
  assign n2651 = ~n2585 & ~n2650 ;
  assign n2652 = n2585 & n2650 ;
  assign n2653 = ~n2651 & ~n2652 ;
  assign n2654 = ~n2640 & ~n2644 ;
  assign n2655 = n2653 & ~n2654 ;
  assign n2656 = ~n2651 & ~n2655 ;
  assign n2657 = ~n2653 & n2654 ;
  assign n2658 = ~n2655 & ~n2657 ;
  assign n2659 = ~n2646 & ~n2648 ;
  assign n2660 = ~n2649 & ~n2659 ;
  assign n2661 = ~n2632 & ~n2634 ;
  assign n2662 = ~n2635 & ~n2661 ;
  assign n2663 = ~x289 & ~x513 ;
  assign n2664 = x289 & x513 ;
  assign n2665 = ~n2663 & ~n2664 ;
  assign n2666 = n2662 & ~n2665 ;
  assign n2667 = ~x296 & ~x520 ;
  assign n2668 = x296 & x520 ;
  assign n2669 = ~n2667 & ~n2668 ;
  assign n2670 = ~x295 & ~x519 ;
  assign n2671 = x295 & x519 ;
  assign n2672 = ~n2670 & ~n2671 ;
  assign n2673 = ~n2669 & ~n2672 ;
  assign n2674 = n2669 & n2672 ;
  assign n2675 = ~n2673 & ~n2674 ;
  assign n2676 = ~x297 & ~x521 ;
  assign n2677 = x297 & x521 ;
  assign n2678 = ~n2676 & ~n2677 ;
  assign n2679 = ~n2675 & ~n2678 ;
  assign n2680 = n2675 & n2678 ;
  assign n2681 = ~n2679 & ~n2680 ;
  assign n2682 = ~x291 & ~x515 ;
  assign n2683 = x291 & x515 ;
  assign n2684 = ~n2682 & ~n2683 ;
  assign n2685 = ~n2681 & ~n2684 ;
  assign n2686 = n2681 & n2684 ;
  assign n2687 = ~n2685 & ~n2686 ;
  assign n2688 = ~x293 & ~x517 ;
  assign n2689 = x293 & x517 ;
  assign n2690 = ~n2688 & ~n2689 ;
  assign n2691 = ~x292 & ~x516 ;
  assign n2692 = x292 & x516 ;
  assign n2693 = ~n2691 & ~n2692 ;
  assign n2694 = ~n2690 & ~n2693 ;
  assign n2695 = n2690 & n2693 ;
  assign n2696 = ~n2694 & ~n2695 ;
  assign n2697 = ~x294 & ~x518 ;
  assign n2698 = x294 & x518 ;
  assign n2699 = ~n2697 & ~n2698 ;
  assign n2700 = ~n2696 & ~n2699 ;
  assign n2701 = n2696 & n2699 ;
  assign n2702 = ~n2700 & ~n2701 ;
  assign n2703 = n2687 & ~n2702 ;
  assign n2704 = ~n2687 & n2702 ;
  assign n2705 = ~n2703 & ~n2704 ;
  assign n2706 = ~x303 & ~x527 ;
  assign n2707 = x303 & x527 ;
  assign n2708 = ~n2706 & ~n2707 ;
  assign n2709 = ~x302 & ~x526 ;
  assign n2710 = x302 & x526 ;
  assign n2711 = ~n2709 & ~n2710 ;
  assign n2712 = ~n2708 & ~n2711 ;
  assign n2713 = n2708 & n2711 ;
  assign n2714 = ~n2712 & ~n2713 ;
  assign n2715 = ~x304 & ~x528 ;
  assign n2716 = x304 & x528 ;
  assign n2717 = ~n2715 & ~n2716 ;
  assign n2718 = ~n2714 & ~n2717 ;
  assign n2719 = n2714 & n2717 ;
  assign n2720 = ~n2718 & ~n2719 ;
  assign n2721 = ~x298 & ~x522 ;
  assign n2722 = x298 & x522 ;
  assign n2723 = ~n2721 & ~n2722 ;
  assign n2724 = ~n2720 & ~n2723 ;
  assign n2725 = n2720 & n2723 ;
  assign n2726 = ~n2724 & ~n2725 ;
  assign n2727 = ~x300 & ~x524 ;
  assign n2728 = x300 & x524 ;
  assign n2729 = ~n2727 & ~n2728 ;
  assign n2730 = ~x299 & ~x523 ;
  assign n2731 = x299 & x523 ;
  assign n2732 = ~n2730 & ~n2731 ;
  assign n2733 = ~n2729 & ~n2732 ;
  assign n2734 = n2729 & n2732 ;
  assign n2735 = ~n2733 & ~n2734 ;
  assign n2736 = ~x301 & ~x525 ;
  assign n2737 = x301 & x525 ;
  assign n2738 = ~n2736 & ~n2737 ;
  assign n2739 = ~n2735 & ~n2738 ;
  assign n2740 = n2735 & n2738 ;
  assign n2741 = ~n2739 & ~n2740 ;
  assign n2742 = n2726 & ~n2741 ;
  assign n2743 = ~n2726 & n2741 ;
  assign n2744 = ~n2742 & ~n2743 ;
  assign n2745 = ~x290 & ~x514 ;
  assign n2746 = x290 & x514 ;
  assign n2747 = ~n2745 & ~n2746 ;
  assign n2748 = n2744 & ~n2747 ;
  assign n2749 = ~n2744 & n2747 ;
  assign n2750 = ~n2748 & ~n2749 ;
  assign n2751 = n2705 & n2750 ;
  assign n2752 = ~n2705 & ~n2750 ;
  assign n2753 = ~n2751 & ~n2752 ;
  assign n2754 = ~n2662 & n2665 ;
  assign n2755 = ~n2666 & ~n2754 ;
  assign n2756 = n2753 & n2755 ;
  assign n2757 = ~n2666 & ~n2756 ;
  assign n2758 = n2660 & ~n2757 ;
  assign n2759 = ~n2685 & ~n2703 ;
  assign n2760 = ~n2674 & ~n2680 ;
  assign n2761 = ~n2759 & n2760 ;
  assign n2762 = n2759 & ~n2760 ;
  assign n2763 = ~n2761 & ~n2762 ;
  assign n2764 = ~n2695 & ~n2701 ;
  assign n2765 = n2763 & n2764 ;
  assign n2766 = ~n2763 & ~n2764 ;
  assign n2767 = ~n2765 & ~n2766 ;
  assign n2768 = ~n2724 & ~n2742 ;
  assign n2769 = ~n2713 & ~n2719 ;
  assign n2770 = ~n2768 & n2769 ;
  assign n2771 = n2768 & ~n2769 ;
  assign n2772 = ~n2770 & ~n2771 ;
  assign n2773 = ~n2734 & ~n2740 ;
  assign n2774 = n2772 & n2773 ;
  assign n2775 = ~n2772 & ~n2773 ;
  assign n2776 = ~n2774 & ~n2775 ;
  assign n2777 = ~n2748 & ~n2751 ;
  assign n2778 = n2776 & ~n2777 ;
  assign n2779 = ~n2776 & n2777 ;
  assign n2780 = ~n2778 & ~n2779 ;
  assign n2781 = n2767 & n2780 ;
  assign n2782 = ~n2767 & ~n2780 ;
  assign n2783 = ~n2781 & ~n2782 ;
  assign n2784 = ~n2660 & n2757 ;
  assign n2785 = ~n2758 & ~n2784 ;
  assign n2786 = n2783 & n2785 ;
  assign n2787 = ~n2758 & ~n2786 ;
  assign n2788 = n2658 & ~n2787 ;
  assign n2789 = ~n2770 & ~n2774 ;
  assign n2790 = ~n2778 & ~n2781 ;
  assign n2791 = ~n2789 & ~n2790 ;
  assign n2792 = n2789 & n2790 ;
  assign n2793 = ~n2791 & ~n2792 ;
  assign n2794 = ~n2761 & ~n2765 ;
  assign n2795 = n2793 & ~n2794 ;
  assign n2796 = ~n2793 & n2794 ;
  assign n2797 = ~n2795 & ~n2796 ;
  assign n2798 = ~n2658 & n2787 ;
  assign n2799 = ~n2788 & ~n2798 ;
  assign n2800 = n2797 & n2799 ;
  assign n2801 = ~n2788 & ~n2800 ;
  assign n2802 = ~n2656 & ~n2801 ;
  assign n2803 = n2656 & n2801 ;
  assign n2804 = ~n2802 & ~n2803 ;
  assign n2805 = ~n2791 & ~n2795 ;
  assign n2806 = n2804 & ~n2805 ;
  assign n2807 = ~n2802 & ~n2806 ;
  assign n2808 = ~n2804 & n2805 ;
  assign n2809 = ~n2806 & ~n2808 ;
  assign n2810 = ~n2797 & ~n2799 ;
  assign n2811 = ~n2800 & ~n2810 ;
  assign n2812 = ~n2783 & ~n2785 ;
  assign n2813 = ~n2786 & ~n2812 ;
  assign n2814 = ~n2753 & ~n2755 ;
  assign n2815 = ~n2756 & ~n2814 ;
  assign n2816 = ~x288 & ~x512 ;
  assign n2817 = x288 & x512 ;
  assign n2818 = ~n2816 & ~n2817 ;
  assign n2819 = ~n2815 & n2818 ;
  assign n2820 = ~n2813 & n2819 ;
  assign n2821 = ~n2811 & n2820 ;
  assign n2822 = ~n2809 & n2821 ;
  assign n2823 = n2807 & n2822 ;
  assign n2824 = n2540 & n2823 ;
  assign n2825 = ~x286 & ~x542 ;
  assign n2826 = x286 & x542 ;
  assign n2827 = ~n2825 & ~n2826 ;
  assign n2828 = ~x285 & ~x541 ;
  assign n2829 = x285 & x541 ;
  assign n2830 = ~n2828 & ~n2829 ;
  assign n2831 = n2827 & n2830 ;
  assign n2832 = ~n2827 & ~n2830 ;
  assign n2833 = ~n2831 & ~n2832 ;
  assign n2834 = ~x287 & ~x543 ;
  assign n2835 = x287 & x543 ;
  assign n2836 = ~n2834 & ~n2835 ;
  assign n2837 = ~n2833 & ~n2836 ;
  assign n2838 = n2833 & n2836 ;
  assign n2839 = ~n2837 & ~n2838 ;
  assign n2840 = ~x281 & ~x537 ;
  assign n2841 = x281 & x537 ;
  assign n2842 = ~n2840 & ~n2841 ;
  assign n2843 = ~n2839 & ~n2842 ;
  assign n2844 = n2839 & n2842 ;
  assign n2845 = ~n2843 & ~n2844 ;
  assign n2846 = ~x283 & ~x539 ;
  assign n2847 = x283 & x539 ;
  assign n2848 = ~n2846 & ~n2847 ;
  assign n2849 = ~x282 & ~x538 ;
  assign n2850 = x282 & x538 ;
  assign n2851 = ~n2849 & ~n2850 ;
  assign n2852 = ~n2848 & ~n2851 ;
  assign n2853 = n2848 & n2851 ;
  assign n2854 = ~n2852 & ~n2853 ;
  assign n2855 = ~x284 & ~x540 ;
  assign n2856 = x284 & x540 ;
  assign n2857 = ~n2855 & ~n2856 ;
  assign n2858 = ~n2854 & ~n2857 ;
  assign n2859 = n2854 & n2857 ;
  assign n2860 = ~n2858 & ~n2859 ;
  assign n2861 = n2845 & ~n2860 ;
  assign n2862 = ~n2843 & ~n2861 ;
  assign n2863 = ~n2831 & ~n2838 ;
  assign n2864 = ~n2862 & n2863 ;
  assign n2865 = n2862 & ~n2863 ;
  assign n2866 = ~n2864 & ~n2865 ;
  assign n2867 = ~n2853 & ~n2859 ;
  assign n2868 = n2866 & n2867 ;
  assign n2869 = ~n2864 & ~n2868 ;
  assign n2870 = ~n2866 & ~n2867 ;
  assign n2871 = ~n2868 & ~n2870 ;
  assign n2872 = ~n2845 & n2860 ;
  assign n2873 = ~n2861 & ~n2872 ;
  assign n2874 = ~x273 & ~x529 ;
  assign n2875 = x273 & x529 ;
  assign n2876 = ~n2874 & ~n2875 ;
  assign n2877 = n2873 & ~n2876 ;
  assign n2878 = ~x279 & ~x535 ;
  assign n2879 = x279 & x535 ;
  assign n2880 = ~n2878 & ~n2879 ;
  assign n2881 = ~x278 & ~x534 ;
  assign n2882 = x278 & x534 ;
  assign n2883 = ~n2881 & ~n2882 ;
  assign n2884 = ~n2880 & ~n2883 ;
  assign n2885 = n2880 & n2883 ;
  assign n2886 = ~n2884 & ~n2885 ;
  assign n2887 = ~x280 & ~x536 ;
  assign n2888 = x280 & x536 ;
  assign n2889 = ~n2887 & ~n2888 ;
  assign n2890 = ~n2886 & ~n2889 ;
  assign n2891 = n2886 & n2889 ;
  assign n2892 = ~n2890 & ~n2891 ;
  assign n2893 = ~x274 & ~x530 ;
  assign n2894 = x274 & x530 ;
  assign n2895 = ~n2893 & ~n2894 ;
  assign n2896 = ~n2892 & ~n2895 ;
  assign n2897 = n2892 & n2895 ;
  assign n2898 = ~n2896 & ~n2897 ;
  assign n2899 = ~x276 & ~x532 ;
  assign n2900 = x276 & x532 ;
  assign n2901 = ~n2899 & ~n2900 ;
  assign n2902 = ~x275 & ~x531 ;
  assign n2903 = x275 & x531 ;
  assign n2904 = ~n2902 & ~n2903 ;
  assign n2905 = ~n2901 & ~n2904 ;
  assign n2906 = n2901 & n2904 ;
  assign n2907 = ~n2905 & ~n2906 ;
  assign n2908 = ~x277 & ~x533 ;
  assign n2909 = x277 & x533 ;
  assign n2910 = ~n2908 & ~n2909 ;
  assign n2911 = ~n2907 & ~n2910 ;
  assign n2912 = n2907 & n2910 ;
  assign n2913 = ~n2911 & ~n2912 ;
  assign n2914 = n2898 & ~n2913 ;
  assign n2915 = ~n2898 & n2913 ;
  assign n2916 = ~n2914 & ~n2915 ;
  assign n2917 = ~n2873 & n2876 ;
  assign n2918 = ~n2877 & ~n2917 ;
  assign n2919 = n2916 & n2918 ;
  assign n2920 = ~n2877 & ~n2919 ;
  assign n2921 = n2871 & ~n2920 ;
  assign n2922 = ~n2896 & ~n2914 ;
  assign n2923 = ~n2885 & ~n2891 ;
  assign n2924 = ~n2922 & n2923 ;
  assign n2925 = n2922 & ~n2923 ;
  assign n2926 = ~n2924 & ~n2925 ;
  assign n2927 = ~n2906 & ~n2912 ;
  assign n2928 = n2926 & n2927 ;
  assign n2929 = ~n2926 & ~n2927 ;
  assign n2930 = ~n2928 & ~n2929 ;
  assign n2931 = ~n2871 & n2920 ;
  assign n2932 = ~n2921 & ~n2931 ;
  assign n2933 = n2930 & n2932 ;
  assign n2934 = ~n2921 & ~n2933 ;
  assign n2935 = ~n2869 & ~n2934 ;
  assign n2936 = n2869 & n2934 ;
  assign n2937 = ~n2935 & ~n2936 ;
  assign n2938 = ~n2924 & ~n2928 ;
  assign n2939 = n2937 & ~n2938 ;
  assign n2940 = ~n2935 & ~n2939 ;
  assign n2941 = ~n2937 & n2938 ;
  assign n2942 = ~n2939 & ~n2941 ;
  assign n2943 = ~n2930 & ~n2932 ;
  assign n2944 = ~n2933 & ~n2943 ;
  assign n2945 = ~n2916 & ~n2918 ;
  assign n2946 = ~n2919 & ~n2945 ;
  assign n2947 = ~x257 & ~x513 ;
  assign n2948 = x257 & x513 ;
  assign n2949 = ~n2947 & ~n2948 ;
  assign n2950 = n2946 & ~n2949 ;
  assign n2951 = ~x264 & ~x520 ;
  assign n2952 = x264 & x520 ;
  assign n2953 = ~n2951 & ~n2952 ;
  assign n2954 = ~x263 & ~x519 ;
  assign n2955 = x263 & x519 ;
  assign n2956 = ~n2954 & ~n2955 ;
  assign n2957 = ~n2953 & ~n2956 ;
  assign n2958 = n2953 & n2956 ;
  assign n2959 = ~n2957 & ~n2958 ;
  assign n2960 = ~x265 & ~x521 ;
  assign n2961 = x265 & x521 ;
  assign n2962 = ~n2960 & ~n2961 ;
  assign n2963 = ~n2959 & ~n2962 ;
  assign n2964 = n2959 & n2962 ;
  assign n2965 = ~n2963 & ~n2964 ;
  assign n2966 = ~x259 & ~x515 ;
  assign n2967 = x259 & x515 ;
  assign n2968 = ~n2966 & ~n2967 ;
  assign n2969 = ~n2965 & ~n2968 ;
  assign n2970 = n2965 & n2968 ;
  assign n2971 = ~n2969 & ~n2970 ;
  assign n2972 = ~x261 & ~x517 ;
  assign n2973 = x261 & x517 ;
  assign n2974 = ~n2972 & ~n2973 ;
  assign n2975 = ~x260 & ~x516 ;
  assign n2976 = x260 & x516 ;
  assign n2977 = ~n2975 & ~n2976 ;
  assign n2978 = ~n2974 & ~n2977 ;
  assign n2979 = n2974 & n2977 ;
  assign n2980 = ~n2978 & ~n2979 ;
  assign n2981 = ~x262 & ~x518 ;
  assign n2982 = x262 & x518 ;
  assign n2983 = ~n2981 & ~n2982 ;
  assign n2984 = ~n2980 & ~n2983 ;
  assign n2985 = n2980 & n2983 ;
  assign n2986 = ~n2984 & ~n2985 ;
  assign n2987 = n2971 & ~n2986 ;
  assign n2988 = ~n2971 & n2986 ;
  assign n2989 = ~n2987 & ~n2988 ;
  assign n2990 = ~x271 & ~x527 ;
  assign n2991 = x271 & x527 ;
  assign n2992 = ~n2990 & ~n2991 ;
  assign n2993 = ~x270 & ~x526 ;
  assign n2994 = x270 & x526 ;
  assign n2995 = ~n2993 & ~n2994 ;
  assign n2996 = ~n2992 & ~n2995 ;
  assign n2997 = n2992 & n2995 ;
  assign n2998 = ~n2996 & ~n2997 ;
  assign n2999 = ~x272 & ~x528 ;
  assign n3000 = x272 & x528 ;
  assign n3001 = ~n2999 & ~n3000 ;
  assign n3002 = ~n2998 & ~n3001 ;
  assign n3003 = n2998 & n3001 ;
  assign n3004 = ~n3002 & ~n3003 ;
  assign n3005 = ~x266 & ~x522 ;
  assign n3006 = x266 & x522 ;
  assign n3007 = ~n3005 & ~n3006 ;
  assign n3008 = ~n3004 & ~n3007 ;
  assign n3009 = n3004 & n3007 ;
  assign n3010 = ~n3008 & ~n3009 ;
  assign n3011 = ~x268 & ~x524 ;
  assign n3012 = x268 & x524 ;
  assign n3013 = ~n3011 & ~n3012 ;
  assign n3014 = ~x267 & ~x523 ;
  assign n3015 = x267 & x523 ;
  assign n3016 = ~n3014 & ~n3015 ;
  assign n3017 = ~n3013 & ~n3016 ;
  assign n3018 = n3013 & n3016 ;
  assign n3019 = ~n3017 & ~n3018 ;
  assign n3020 = ~x269 & ~x525 ;
  assign n3021 = x269 & x525 ;
  assign n3022 = ~n3020 & ~n3021 ;
  assign n3023 = ~n3019 & ~n3022 ;
  assign n3024 = n3019 & n3022 ;
  assign n3025 = ~n3023 & ~n3024 ;
  assign n3026 = n3010 & ~n3025 ;
  assign n3027 = ~n3010 & n3025 ;
  assign n3028 = ~n3026 & ~n3027 ;
  assign n3029 = ~x258 & ~x514 ;
  assign n3030 = x258 & x514 ;
  assign n3031 = ~n3029 & ~n3030 ;
  assign n3032 = n3028 & ~n3031 ;
  assign n3033 = ~n3028 & n3031 ;
  assign n3034 = ~n3032 & ~n3033 ;
  assign n3035 = n2989 & n3034 ;
  assign n3036 = ~n2989 & ~n3034 ;
  assign n3037 = ~n3035 & ~n3036 ;
  assign n3038 = ~n2946 & n2949 ;
  assign n3039 = ~n2950 & ~n3038 ;
  assign n3040 = n3037 & n3039 ;
  assign n3041 = ~n2950 & ~n3040 ;
  assign n3042 = n2944 & ~n3041 ;
  assign n3043 = ~n2969 & ~n2987 ;
  assign n3044 = ~n2958 & ~n2964 ;
  assign n3045 = ~n3043 & n3044 ;
  assign n3046 = n3043 & ~n3044 ;
  assign n3047 = ~n3045 & ~n3046 ;
  assign n3048 = ~n2979 & ~n2985 ;
  assign n3049 = n3047 & n3048 ;
  assign n3050 = ~n3047 & ~n3048 ;
  assign n3051 = ~n3049 & ~n3050 ;
  assign n3052 = ~n3008 & ~n3026 ;
  assign n3053 = ~n2997 & ~n3003 ;
  assign n3054 = ~n3052 & n3053 ;
  assign n3055 = n3052 & ~n3053 ;
  assign n3056 = ~n3054 & ~n3055 ;
  assign n3057 = ~n3018 & ~n3024 ;
  assign n3058 = n3056 & n3057 ;
  assign n3059 = ~n3056 & ~n3057 ;
  assign n3060 = ~n3058 & ~n3059 ;
  assign n3061 = ~n3032 & ~n3035 ;
  assign n3062 = n3060 & ~n3061 ;
  assign n3063 = ~n3060 & n3061 ;
  assign n3064 = ~n3062 & ~n3063 ;
  assign n3065 = n3051 & n3064 ;
  assign n3066 = ~n3051 & ~n3064 ;
  assign n3067 = ~n3065 & ~n3066 ;
  assign n3068 = ~n2944 & n3041 ;
  assign n3069 = ~n3042 & ~n3068 ;
  assign n3070 = n3067 & n3069 ;
  assign n3071 = ~n3042 & ~n3070 ;
  assign n3072 = n2942 & ~n3071 ;
  assign n3073 = ~n3054 & ~n3058 ;
  assign n3074 = ~n3062 & ~n3065 ;
  assign n3075 = ~n3073 & ~n3074 ;
  assign n3076 = n3073 & n3074 ;
  assign n3077 = ~n3075 & ~n3076 ;
  assign n3078 = ~n3045 & ~n3049 ;
  assign n3079 = n3077 & ~n3078 ;
  assign n3080 = ~n3077 & n3078 ;
  assign n3081 = ~n3079 & ~n3080 ;
  assign n3082 = ~n2942 & n3071 ;
  assign n3083 = ~n3072 & ~n3082 ;
  assign n3084 = n3081 & n3083 ;
  assign n3085 = ~n3072 & ~n3084 ;
  assign n3086 = ~n2940 & ~n3085 ;
  assign n3087 = n2940 & n3085 ;
  assign n3088 = ~n3086 & ~n3087 ;
  assign n3089 = ~n3075 & ~n3079 ;
  assign n3090 = n3088 & ~n3089 ;
  assign n3091 = ~n3086 & ~n3090 ;
  assign n3092 = ~n3088 & n3089 ;
  assign n3093 = ~n3090 & ~n3092 ;
  assign n3094 = ~n3081 & ~n3083 ;
  assign n3095 = ~n3084 & ~n3094 ;
  assign n3096 = ~n3067 & ~n3069 ;
  assign n3097 = ~n3070 & ~n3096 ;
  assign n3098 = ~n3037 & ~n3039 ;
  assign n3099 = ~n3040 & ~n3098 ;
  assign n3100 = ~x256 & ~x512 ;
  assign n3101 = x256 & x512 ;
  assign n3102 = ~n3100 & ~n3101 ;
  assign n3103 = ~n3099 & n3102 ;
  assign n3104 = ~n3097 & n3103 ;
  assign n3105 = ~n3095 & n3104 ;
  assign n3106 = ~n3093 & n3105 ;
  assign n3107 = n3091 & n3106 ;
  assign n3108 = n2824 & n3107 ;
  assign n3109 = ~x254 & ~x542 ;
  assign n3110 = x254 & x542 ;
  assign n3111 = ~n3109 & ~n3110 ;
  assign n3112 = ~x253 & ~x541 ;
  assign n3113 = x253 & x541 ;
  assign n3114 = ~n3112 & ~n3113 ;
  assign n3115 = n3111 & n3114 ;
  assign n3116 = ~n3111 & ~n3114 ;
  assign n3117 = ~n3115 & ~n3116 ;
  assign n3118 = ~x255 & ~x543 ;
  assign n3119 = x255 & x543 ;
  assign n3120 = ~n3118 & ~n3119 ;
  assign n3121 = ~n3117 & ~n3120 ;
  assign n3122 = n3117 & n3120 ;
  assign n3123 = ~n3121 & ~n3122 ;
  assign n3124 = ~x249 & ~x537 ;
  assign n3125 = x249 & x537 ;
  assign n3126 = ~n3124 & ~n3125 ;
  assign n3127 = ~n3123 & ~n3126 ;
  assign n3128 = n3123 & n3126 ;
  assign n3129 = ~n3127 & ~n3128 ;
  assign n3130 = ~x251 & ~x539 ;
  assign n3131 = x251 & x539 ;
  assign n3132 = ~n3130 & ~n3131 ;
  assign n3133 = ~x250 & ~x538 ;
  assign n3134 = x250 & x538 ;
  assign n3135 = ~n3133 & ~n3134 ;
  assign n3136 = ~n3132 & ~n3135 ;
  assign n3137 = n3132 & n3135 ;
  assign n3138 = ~n3136 & ~n3137 ;
  assign n3139 = ~x252 & ~x540 ;
  assign n3140 = x252 & x540 ;
  assign n3141 = ~n3139 & ~n3140 ;
  assign n3142 = ~n3138 & ~n3141 ;
  assign n3143 = n3138 & n3141 ;
  assign n3144 = ~n3142 & ~n3143 ;
  assign n3145 = n3129 & ~n3144 ;
  assign n3146 = ~n3127 & ~n3145 ;
  assign n3147 = ~n3115 & ~n3122 ;
  assign n3148 = ~n3146 & n3147 ;
  assign n3149 = n3146 & ~n3147 ;
  assign n3150 = ~n3148 & ~n3149 ;
  assign n3151 = ~n3137 & ~n3143 ;
  assign n3152 = n3150 & n3151 ;
  assign n3153 = ~n3148 & ~n3152 ;
  assign n3154 = ~n3150 & ~n3151 ;
  assign n3155 = ~n3152 & ~n3154 ;
  assign n3156 = ~n3129 & n3144 ;
  assign n3157 = ~n3145 & ~n3156 ;
  assign n3158 = ~x241 & ~x529 ;
  assign n3159 = x241 & x529 ;
  assign n3160 = ~n3158 & ~n3159 ;
  assign n3161 = n3157 & ~n3160 ;
  assign n3162 = ~x247 & ~x535 ;
  assign n3163 = x247 & x535 ;
  assign n3164 = ~n3162 & ~n3163 ;
  assign n3165 = ~x246 & ~x534 ;
  assign n3166 = x246 & x534 ;
  assign n3167 = ~n3165 & ~n3166 ;
  assign n3168 = ~n3164 & ~n3167 ;
  assign n3169 = n3164 & n3167 ;
  assign n3170 = ~n3168 & ~n3169 ;
  assign n3171 = ~x248 & ~x536 ;
  assign n3172 = x248 & x536 ;
  assign n3173 = ~n3171 & ~n3172 ;
  assign n3174 = ~n3170 & ~n3173 ;
  assign n3175 = n3170 & n3173 ;
  assign n3176 = ~n3174 & ~n3175 ;
  assign n3177 = ~x242 & ~x530 ;
  assign n3178 = x242 & x530 ;
  assign n3179 = ~n3177 & ~n3178 ;
  assign n3180 = ~n3176 & ~n3179 ;
  assign n3181 = n3176 & n3179 ;
  assign n3182 = ~n3180 & ~n3181 ;
  assign n3183 = ~x244 & ~x532 ;
  assign n3184 = x244 & x532 ;
  assign n3185 = ~n3183 & ~n3184 ;
  assign n3186 = ~x243 & ~x531 ;
  assign n3187 = x243 & x531 ;
  assign n3188 = ~n3186 & ~n3187 ;
  assign n3189 = ~n3185 & ~n3188 ;
  assign n3190 = n3185 & n3188 ;
  assign n3191 = ~n3189 & ~n3190 ;
  assign n3192 = ~x245 & ~x533 ;
  assign n3193 = x245 & x533 ;
  assign n3194 = ~n3192 & ~n3193 ;
  assign n3195 = ~n3191 & ~n3194 ;
  assign n3196 = n3191 & n3194 ;
  assign n3197 = ~n3195 & ~n3196 ;
  assign n3198 = n3182 & ~n3197 ;
  assign n3199 = ~n3182 & n3197 ;
  assign n3200 = ~n3198 & ~n3199 ;
  assign n3201 = ~n3157 & n3160 ;
  assign n3202 = ~n3161 & ~n3201 ;
  assign n3203 = n3200 & n3202 ;
  assign n3204 = ~n3161 & ~n3203 ;
  assign n3205 = n3155 & ~n3204 ;
  assign n3206 = ~n3180 & ~n3198 ;
  assign n3207 = ~n3169 & ~n3175 ;
  assign n3208 = ~n3206 & n3207 ;
  assign n3209 = n3206 & ~n3207 ;
  assign n3210 = ~n3208 & ~n3209 ;
  assign n3211 = ~n3190 & ~n3196 ;
  assign n3212 = n3210 & n3211 ;
  assign n3213 = ~n3210 & ~n3211 ;
  assign n3214 = ~n3212 & ~n3213 ;
  assign n3215 = ~n3155 & n3204 ;
  assign n3216 = ~n3205 & ~n3215 ;
  assign n3217 = n3214 & n3216 ;
  assign n3218 = ~n3205 & ~n3217 ;
  assign n3219 = ~n3153 & ~n3218 ;
  assign n3220 = n3153 & n3218 ;
  assign n3221 = ~n3219 & ~n3220 ;
  assign n3222 = ~n3208 & ~n3212 ;
  assign n3223 = n3221 & ~n3222 ;
  assign n3224 = ~n3219 & ~n3223 ;
  assign n3225 = ~n3221 & n3222 ;
  assign n3226 = ~n3223 & ~n3225 ;
  assign n3227 = ~n3214 & ~n3216 ;
  assign n3228 = ~n3217 & ~n3227 ;
  assign n3229 = ~n3200 & ~n3202 ;
  assign n3230 = ~n3203 & ~n3229 ;
  assign n3231 = ~x225 & ~x513 ;
  assign n3232 = x225 & x513 ;
  assign n3233 = ~n3231 & ~n3232 ;
  assign n3234 = n3230 & ~n3233 ;
  assign n3235 = ~x232 & ~x520 ;
  assign n3236 = x232 & x520 ;
  assign n3237 = ~n3235 & ~n3236 ;
  assign n3238 = ~x231 & ~x519 ;
  assign n3239 = x231 & x519 ;
  assign n3240 = ~n3238 & ~n3239 ;
  assign n3241 = ~n3237 & ~n3240 ;
  assign n3242 = n3237 & n3240 ;
  assign n3243 = ~n3241 & ~n3242 ;
  assign n3244 = ~x233 & ~x521 ;
  assign n3245 = x233 & x521 ;
  assign n3246 = ~n3244 & ~n3245 ;
  assign n3247 = ~n3243 & ~n3246 ;
  assign n3248 = n3243 & n3246 ;
  assign n3249 = ~n3247 & ~n3248 ;
  assign n3250 = ~x227 & ~x515 ;
  assign n3251 = x227 & x515 ;
  assign n3252 = ~n3250 & ~n3251 ;
  assign n3253 = ~n3249 & ~n3252 ;
  assign n3254 = n3249 & n3252 ;
  assign n3255 = ~n3253 & ~n3254 ;
  assign n3256 = ~x229 & ~x517 ;
  assign n3257 = x229 & x517 ;
  assign n3258 = ~n3256 & ~n3257 ;
  assign n3259 = ~x228 & ~x516 ;
  assign n3260 = x228 & x516 ;
  assign n3261 = ~n3259 & ~n3260 ;
  assign n3262 = ~n3258 & ~n3261 ;
  assign n3263 = n3258 & n3261 ;
  assign n3264 = ~n3262 & ~n3263 ;
  assign n3265 = ~x230 & ~x518 ;
  assign n3266 = x230 & x518 ;
  assign n3267 = ~n3265 & ~n3266 ;
  assign n3268 = ~n3264 & ~n3267 ;
  assign n3269 = n3264 & n3267 ;
  assign n3270 = ~n3268 & ~n3269 ;
  assign n3271 = n3255 & ~n3270 ;
  assign n3272 = ~n3255 & n3270 ;
  assign n3273 = ~n3271 & ~n3272 ;
  assign n3274 = ~x239 & ~x527 ;
  assign n3275 = x239 & x527 ;
  assign n3276 = ~n3274 & ~n3275 ;
  assign n3277 = ~x238 & ~x526 ;
  assign n3278 = x238 & x526 ;
  assign n3279 = ~n3277 & ~n3278 ;
  assign n3280 = ~n3276 & ~n3279 ;
  assign n3281 = n3276 & n3279 ;
  assign n3282 = ~n3280 & ~n3281 ;
  assign n3283 = ~x240 & ~x528 ;
  assign n3284 = x240 & x528 ;
  assign n3285 = ~n3283 & ~n3284 ;
  assign n3286 = ~n3282 & ~n3285 ;
  assign n3287 = n3282 & n3285 ;
  assign n3288 = ~n3286 & ~n3287 ;
  assign n3289 = ~x234 & ~x522 ;
  assign n3290 = x234 & x522 ;
  assign n3291 = ~n3289 & ~n3290 ;
  assign n3292 = ~n3288 & ~n3291 ;
  assign n3293 = n3288 & n3291 ;
  assign n3294 = ~n3292 & ~n3293 ;
  assign n3295 = ~x236 & ~x524 ;
  assign n3296 = x236 & x524 ;
  assign n3297 = ~n3295 & ~n3296 ;
  assign n3298 = ~x235 & ~x523 ;
  assign n3299 = x235 & x523 ;
  assign n3300 = ~n3298 & ~n3299 ;
  assign n3301 = ~n3297 & ~n3300 ;
  assign n3302 = n3297 & n3300 ;
  assign n3303 = ~n3301 & ~n3302 ;
  assign n3304 = ~x237 & ~x525 ;
  assign n3305 = x237 & x525 ;
  assign n3306 = ~n3304 & ~n3305 ;
  assign n3307 = ~n3303 & ~n3306 ;
  assign n3308 = n3303 & n3306 ;
  assign n3309 = ~n3307 & ~n3308 ;
  assign n3310 = n3294 & ~n3309 ;
  assign n3311 = ~n3294 & n3309 ;
  assign n3312 = ~n3310 & ~n3311 ;
  assign n3313 = ~x226 & ~x514 ;
  assign n3314 = x226 & x514 ;
  assign n3315 = ~n3313 & ~n3314 ;
  assign n3316 = n3312 & ~n3315 ;
  assign n3317 = ~n3312 & n3315 ;
  assign n3318 = ~n3316 & ~n3317 ;
  assign n3319 = n3273 & n3318 ;
  assign n3320 = ~n3273 & ~n3318 ;
  assign n3321 = ~n3319 & ~n3320 ;
  assign n3322 = ~n3230 & n3233 ;
  assign n3323 = ~n3234 & ~n3322 ;
  assign n3324 = n3321 & n3323 ;
  assign n3325 = ~n3234 & ~n3324 ;
  assign n3326 = n3228 & ~n3325 ;
  assign n3327 = ~n3253 & ~n3271 ;
  assign n3328 = ~n3242 & ~n3248 ;
  assign n3329 = ~n3327 & n3328 ;
  assign n3330 = n3327 & ~n3328 ;
  assign n3331 = ~n3329 & ~n3330 ;
  assign n3332 = ~n3263 & ~n3269 ;
  assign n3333 = n3331 & n3332 ;
  assign n3334 = ~n3331 & ~n3332 ;
  assign n3335 = ~n3333 & ~n3334 ;
  assign n3336 = ~n3292 & ~n3310 ;
  assign n3337 = ~n3281 & ~n3287 ;
  assign n3338 = ~n3336 & n3337 ;
  assign n3339 = n3336 & ~n3337 ;
  assign n3340 = ~n3338 & ~n3339 ;
  assign n3341 = ~n3302 & ~n3308 ;
  assign n3342 = n3340 & n3341 ;
  assign n3343 = ~n3340 & ~n3341 ;
  assign n3344 = ~n3342 & ~n3343 ;
  assign n3345 = ~n3316 & ~n3319 ;
  assign n3346 = n3344 & ~n3345 ;
  assign n3347 = ~n3344 & n3345 ;
  assign n3348 = ~n3346 & ~n3347 ;
  assign n3349 = n3335 & n3348 ;
  assign n3350 = ~n3335 & ~n3348 ;
  assign n3351 = ~n3349 & ~n3350 ;
  assign n3352 = ~n3228 & n3325 ;
  assign n3353 = ~n3326 & ~n3352 ;
  assign n3354 = n3351 & n3353 ;
  assign n3355 = ~n3326 & ~n3354 ;
  assign n3356 = n3226 & ~n3355 ;
  assign n3357 = ~n3338 & ~n3342 ;
  assign n3358 = ~n3346 & ~n3349 ;
  assign n3359 = ~n3357 & ~n3358 ;
  assign n3360 = n3357 & n3358 ;
  assign n3361 = ~n3359 & ~n3360 ;
  assign n3362 = ~n3329 & ~n3333 ;
  assign n3363 = n3361 & ~n3362 ;
  assign n3364 = ~n3361 & n3362 ;
  assign n3365 = ~n3363 & ~n3364 ;
  assign n3366 = ~n3226 & n3355 ;
  assign n3367 = ~n3356 & ~n3366 ;
  assign n3368 = n3365 & n3367 ;
  assign n3369 = ~n3356 & ~n3368 ;
  assign n3370 = ~n3224 & ~n3369 ;
  assign n3371 = n3224 & n3369 ;
  assign n3372 = ~n3370 & ~n3371 ;
  assign n3373 = ~n3359 & ~n3363 ;
  assign n3374 = n3372 & ~n3373 ;
  assign n3375 = ~n3370 & ~n3374 ;
  assign n3376 = ~n3372 & n3373 ;
  assign n3377 = ~n3374 & ~n3376 ;
  assign n3378 = ~n3365 & ~n3367 ;
  assign n3379 = ~n3368 & ~n3378 ;
  assign n3380 = ~n3351 & ~n3353 ;
  assign n3381 = ~n3354 & ~n3380 ;
  assign n3382 = ~n3321 & ~n3323 ;
  assign n3383 = ~n3324 & ~n3382 ;
  assign n3384 = ~x224 & ~x512 ;
  assign n3385 = x224 & x512 ;
  assign n3386 = ~n3384 & ~n3385 ;
  assign n3387 = ~n3383 & n3386 ;
  assign n3388 = ~n3381 & n3387 ;
  assign n3389 = ~n3379 & n3388 ;
  assign n3390 = ~n3377 & n3389 ;
  assign n3391 = n3375 & n3390 ;
  assign n3392 = n3108 & n3391 ;
  assign n3393 = ~x222 & ~x542 ;
  assign n3394 = x222 & x542 ;
  assign n3395 = ~n3393 & ~n3394 ;
  assign n3396 = ~x221 & ~x541 ;
  assign n3397 = x221 & x541 ;
  assign n3398 = ~n3396 & ~n3397 ;
  assign n3399 = n3395 & n3398 ;
  assign n3400 = ~n3395 & ~n3398 ;
  assign n3401 = ~n3399 & ~n3400 ;
  assign n3402 = ~x223 & ~x543 ;
  assign n3403 = x223 & x543 ;
  assign n3404 = ~n3402 & ~n3403 ;
  assign n3405 = ~n3401 & ~n3404 ;
  assign n3406 = n3401 & n3404 ;
  assign n3407 = ~n3405 & ~n3406 ;
  assign n3408 = ~x217 & ~x537 ;
  assign n3409 = x217 & x537 ;
  assign n3410 = ~n3408 & ~n3409 ;
  assign n3411 = ~n3407 & ~n3410 ;
  assign n3412 = n3407 & n3410 ;
  assign n3413 = ~n3411 & ~n3412 ;
  assign n3414 = ~x219 & ~x539 ;
  assign n3415 = x219 & x539 ;
  assign n3416 = ~n3414 & ~n3415 ;
  assign n3417 = ~x218 & ~x538 ;
  assign n3418 = x218 & x538 ;
  assign n3419 = ~n3417 & ~n3418 ;
  assign n3420 = ~n3416 & ~n3419 ;
  assign n3421 = n3416 & n3419 ;
  assign n3422 = ~n3420 & ~n3421 ;
  assign n3423 = ~x220 & ~x540 ;
  assign n3424 = x220 & x540 ;
  assign n3425 = ~n3423 & ~n3424 ;
  assign n3426 = ~n3422 & ~n3425 ;
  assign n3427 = n3422 & n3425 ;
  assign n3428 = ~n3426 & ~n3427 ;
  assign n3429 = n3413 & ~n3428 ;
  assign n3430 = ~n3411 & ~n3429 ;
  assign n3431 = ~n3399 & ~n3406 ;
  assign n3432 = ~n3430 & n3431 ;
  assign n3433 = n3430 & ~n3431 ;
  assign n3434 = ~n3432 & ~n3433 ;
  assign n3435 = ~n3421 & ~n3427 ;
  assign n3436 = n3434 & n3435 ;
  assign n3437 = ~n3432 & ~n3436 ;
  assign n3438 = ~n3434 & ~n3435 ;
  assign n3439 = ~n3436 & ~n3438 ;
  assign n3440 = ~n3413 & n3428 ;
  assign n3441 = ~n3429 & ~n3440 ;
  assign n3442 = ~x209 & ~x529 ;
  assign n3443 = x209 & x529 ;
  assign n3444 = ~n3442 & ~n3443 ;
  assign n3445 = n3441 & ~n3444 ;
  assign n3446 = ~x215 & ~x535 ;
  assign n3447 = x215 & x535 ;
  assign n3448 = ~n3446 & ~n3447 ;
  assign n3449 = ~x214 & ~x534 ;
  assign n3450 = x214 & x534 ;
  assign n3451 = ~n3449 & ~n3450 ;
  assign n3452 = ~n3448 & ~n3451 ;
  assign n3453 = n3448 & n3451 ;
  assign n3454 = ~n3452 & ~n3453 ;
  assign n3455 = ~x216 & ~x536 ;
  assign n3456 = x216 & x536 ;
  assign n3457 = ~n3455 & ~n3456 ;
  assign n3458 = ~n3454 & ~n3457 ;
  assign n3459 = n3454 & n3457 ;
  assign n3460 = ~n3458 & ~n3459 ;
  assign n3461 = ~x210 & ~x530 ;
  assign n3462 = x210 & x530 ;
  assign n3463 = ~n3461 & ~n3462 ;
  assign n3464 = ~n3460 & ~n3463 ;
  assign n3465 = n3460 & n3463 ;
  assign n3466 = ~n3464 & ~n3465 ;
  assign n3467 = ~x212 & ~x532 ;
  assign n3468 = x212 & x532 ;
  assign n3469 = ~n3467 & ~n3468 ;
  assign n3470 = ~x211 & ~x531 ;
  assign n3471 = x211 & x531 ;
  assign n3472 = ~n3470 & ~n3471 ;
  assign n3473 = ~n3469 & ~n3472 ;
  assign n3474 = n3469 & n3472 ;
  assign n3475 = ~n3473 & ~n3474 ;
  assign n3476 = ~x213 & ~x533 ;
  assign n3477 = x213 & x533 ;
  assign n3478 = ~n3476 & ~n3477 ;
  assign n3479 = ~n3475 & ~n3478 ;
  assign n3480 = n3475 & n3478 ;
  assign n3481 = ~n3479 & ~n3480 ;
  assign n3482 = n3466 & ~n3481 ;
  assign n3483 = ~n3466 & n3481 ;
  assign n3484 = ~n3482 & ~n3483 ;
  assign n3485 = ~n3441 & n3444 ;
  assign n3486 = ~n3445 & ~n3485 ;
  assign n3487 = n3484 & n3486 ;
  assign n3488 = ~n3445 & ~n3487 ;
  assign n3489 = n3439 & ~n3488 ;
  assign n3490 = ~n3464 & ~n3482 ;
  assign n3491 = ~n3453 & ~n3459 ;
  assign n3492 = ~n3490 & n3491 ;
  assign n3493 = n3490 & ~n3491 ;
  assign n3494 = ~n3492 & ~n3493 ;
  assign n3495 = ~n3474 & ~n3480 ;
  assign n3496 = n3494 & n3495 ;
  assign n3497 = ~n3494 & ~n3495 ;
  assign n3498 = ~n3496 & ~n3497 ;
  assign n3499 = ~n3439 & n3488 ;
  assign n3500 = ~n3489 & ~n3499 ;
  assign n3501 = n3498 & n3500 ;
  assign n3502 = ~n3489 & ~n3501 ;
  assign n3503 = ~n3437 & ~n3502 ;
  assign n3504 = n3437 & n3502 ;
  assign n3505 = ~n3503 & ~n3504 ;
  assign n3506 = ~n3492 & ~n3496 ;
  assign n3507 = n3505 & ~n3506 ;
  assign n3508 = ~n3503 & ~n3507 ;
  assign n3509 = ~n3505 & n3506 ;
  assign n3510 = ~n3507 & ~n3509 ;
  assign n3511 = ~n3498 & ~n3500 ;
  assign n3512 = ~n3501 & ~n3511 ;
  assign n3513 = ~n3484 & ~n3486 ;
  assign n3514 = ~n3487 & ~n3513 ;
  assign n3515 = ~x193 & ~x513 ;
  assign n3516 = x193 & x513 ;
  assign n3517 = ~n3515 & ~n3516 ;
  assign n3518 = n3514 & ~n3517 ;
  assign n3519 = ~x200 & ~x520 ;
  assign n3520 = x200 & x520 ;
  assign n3521 = ~n3519 & ~n3520 ;
  assign n3522 = ~x199 & ~x519 ;
  assign n3523 = x199 & x519 ;
  assign n3524 = ~n3522 & ~n3523 ;
  assign n3525 = ~n3521 & ~n3524 ;
  assign n3526 = n3521 & n3524 ;
  assign n3527 = ~n3525 & ~n3526 ;
  assign n3528 = ~x201 & ~x521 ;
  assign n3529 = x201 & x521 ;
  assign n3530 = ~n3528 & ~n3529 ;
  assign n3531 = ~n3527 & ~n3530 ;
  assign n3532 = n3527 & n3530 ;
  assign n3533 = ~n3531 & ~n3532 ;
  assign n3534 = ~x195 & ~x515 ;
  assign n3535 = x195 & x515 ;
  assign n3536 = ~n3534 & ~n3535 ;
  assign n3537 = ~n3533 & ~n3536 ;
  assign n3538 = n3533 & n3536 ;
  assign n3539 = ~n3537 & ~n3538 ;
  assign n3540 = ~x197 & ~x517 ;
  assign n3541 = x197 & x517 ;
  assign n3542 = ~n3540 & ~n3541 ;
  assign n3543 = ~x196 & ~x516 ;
  assign n3544 = x196 & x516 ;
  assign n3545 = ~n3543 & ~n3544 ;
  assign n3546 = ~n3542 & ~n3545 ;
  assign n3547 = n3542 & n3545 ;
  assign n3548 = ~n3546 & ~n3547 ;
  assign n3549 = ~x198 & ~x518 ;
  assign n3550 = x198 & x518 ;
  assign n3551 = ~n3549 & ~n3550 ;
  assign n3552 = ~n3548 & ~n3551 ;
  assign n3553 = n3548 & n3551 ;
  assign n3554 = ~n3552 & ~n3553 ;
  assign n3555 = n3539 & ~n3554 ;
  assign n3556 = ~n3539 & n3554 ;
  assign n3557 = ~n3555 & ~n3556 ;
  assign n3558 = ~x207 & ~x527 ;
  assign n3559 = x207 & x527 ;
  assign n3560 = ~n3558 & ~n3559 ;
  assign n3561 = ~x206 & ~x526 ;
  assign n3562 = x206 & x526 ;
  assign n3563 = ~n3561 & ~n3562 ;
  assign n3564 = ~n3560 & ~n3563 ;
  assign n3565 = n3560 & n3563 ;
  assign n3566 = ~n3564 & ~n3565 ;
  assign n3567 = ~x208 & ~x528 ;
  assign n3568 = x208 & x528 ;
  assign n3569 = ~n3567 & ~n3568 ;
  assign n3570 = ~n3566 & ~n3569 ;
  assign n3571 = n3566 & n3569 ;
  assign n3572 = ~n3570 & ~n3571 ;
  assign n3573 = ~x202 & ~x522 ;
  assign n3574 = x202 & x522 ;
  assign n3575 = ~n3573 & ~n3574 ;
  assign n3576 = ~n3572 & ~n3575 ;
  assign n3577 = n3572 & n3575 ;
  assign n3578 = ~n3576 & ~n3577 ;
  assign n3579 = ~x204 & ~x524 ;
  assign n3580 = x204 & x524 ;
  assign n3581 = ~n3579 & ~n3580 ;
  assign n3582 = ~x203 & ~x523 ;
  assign n3583 = x203 & x523 ;
  assign n3584 = ~n3582 & ~n3583 ;
  assign n3585 = ~n3581 & ~n3584 ;
  assign n3586 = n3581 & n3584 ;
  assign n3587 = ~n3585 & ~n3586 ;
  assign n3588 = ~x205 & ~x525 ;
  assign n3589 = x205 & x525 ;
  assign n3590 = ~n3588 & ~n3589 ;
  assign n3591 = ~n3587 & ~n3590 ;
  assign n3592 = n3587 & n3590 ;
  assign n3593 = ~n3591 & ~n3592 ;
  assign n3594 = n3578 & ~n3593 ;
  assign n3595 = ~n3578 & n3593 ;
  assign n3596 = ~n3594 & ~n3595 ;
  assign n3597 = ~x194 & ~x514 ;
  assign n3598 = x194 & x514 ;
  assign n3599 = ~n3597 & ~n3598 ;
  assign n3600 = n3596 & ~n3599 ;
  assign n3601 = ~n3596 & n3599 ;
  assign n3602 = ~n3600 & ~n3601 ;
  assign n3603 = n3557 & n3602 ;
  assign n3604 = ~n3557 & ~n3602 ;
  assign n3605 = ~n3603 & ~n3604 ;
  assign n3606 = ~n3514 & n3517 ;
  assign n3607 = ~n3518 & ~n3606 ;
  assign n3608 = n3605 & n3607 ;
  assign n3609 = ~n3518 & ~n3608 ;
  assign n3610 = n3512 & ~n3609 ;
  assign n3611 = ~n3537 & ~n3555 ;
  assign n3612 = ~n3526 & ~n3532 ;
  assign n3613 = ~n3611 & n3612 ;
  assign n3614 = n3611 & ~n3612 ;
  assign n3615 = ~n3613 & ~n3614 ;
  assign n3616 = ~n3547 & ~n3553 ;
  assign n3617 = n3615 & n3616 ;
  assign n3618 = ~n3615 & ~n3616 ;
  assign n3619 = ~n3617 & ~n3618 ;
  assign n3620 = ~n3576 & ~n3594 ;
  assign n3621 = ~n3565 & ~n3571 ;
  assign n3622 = ~n3620 & n3621 ;
  assign n3623 = n3620 & ~n3621 ;
  assign n3624 = ~n3622 & ~n3623 ;
  assign n3625 = ~n3586 & ~n3592 ;
  assign n3626 = n3624 & n3625 ;
  assign n3627 = ~n3624 & ~n3625 ;
  assign n3628 = ~n3626 & ~n3627 ;
  assign n3629 = ~n3600 & ~n3603 ;
  assign n3630 = n3628 & ~n3629 ;
  assign n3631 = ~n3628 & n3629 ;
  assign n3632 = ~n3630 & ~n3631 ;
  assign n3633 = n3619 & n3632 ;
  assign n3634 = ~n3619 & ~n3632 ;
  assign n3635 = ~n3633 & ~n3634 ;
  assign n3636 = ~n3512 & n3609 ;
  assign n3637 = ~n3610 & ~n3636 ;
  assign n3638 = n3635 & n3637 ;
  assign n3639 = ~n3610 & ~n3638 ;
  assign n3640 = n3510 & ~n3639 ;
  assign n3641 = ~n3622 & ~n3626 ;
  assign n3642 = ~n3630 & ~n3633 ;
  assign n3643 = ~n3641 & ~n3642 ;
  assign n3644 = n3641 & n3642 ;
  assign n3645 = ~n3643 & ~n3644 ;
  assign n3646 = ~n3613 & ~n3617 ;
  assign n3647 = n3645 & ~n3646 ;
  assign n3648 = ~n3645 & n3646 ;
  assign n3649 = ~n3647 & ~n3648 ;
  assign n3650 = ~n3510 & n3639 ;
  assign n3651 = ~n3640 & ~n3650 ;
  assign n3652 = n3649 & n3651 ;
  assign n3653 = ~n3640 & ~n3652 ;
  assign n3654 = ~n3508 & ~n3653 ;
  assign n3655 = n3508 & n3653 ;
  assign n3656 = ~n3654 & ~n3655 ;
  assign n3657 = ~n3643 & ~n3647 ;
  assign n3658 = n3656 & ~n3657 ;
  assign n3659 = ~n3654 & ~n3658 ;
  assign n3660 = ~n3656 & n3657 ;
  assign n3661 = ~n3658 & ~n3660 ;
  assign n3662 = ~n3649 & ~n3651 ;
  assign n3663 = ~n3652 & ~n3662 ;
  assign n3664 = ~n3635 & ~n3637 ;
  assign n3665 = ~n3638 & ~n3664 ;
  assign n3666 = ~n3605 & ~n3607 ;
  assign n3667 = ~n3608 & ~n3666 ;
  assign n3668 = ~x192 & ~x512 ;
  assign n3669 = x192 & x512 ;
  assign n3670 = ~n3668 & ~n3669 ;
  assign n3671 = ~n3667 & n3670 ;
  assign n3672 = ~n3665 & n3671 ;
  assign n3673 = ~n3663 & n3672 ;
  assign n3674 = ~n3661 & n3673 ;
  assign n3675 = n3659 & n3674 ;
  assign n3676 = n3392 & n3675 ;
  assign n3677 = ~x190 & ~x542 ;
  assign n3678 = x190 & x542 ;
  assign n3679 = ~n3677 & ~n3678 ;
  assign n3680 = ~x189 & ~x541 ;
  assign n3681 = x189 & x541 ;
  assign n3682 = ~n3680 & ~n3681 ;
  assign n3683 = n3679 & n3682 ;
  assign n3684 = ~n3679 & ~n3682 ;
  assign n3685 = ~n3683 & ~n3684 ;
  assign n3686 = ~x191 & ~x543 ;
  assign n3687 = x191 & x543 ;
  assign n3688 = ~n3686 & ~n3687 ;
  assign n3689 = ~n3685 & ~n3688 ;
  assign n3690 = n3685 & n3688 ;
  assign n3691 = ~n3689 & ~n3690 ;
  assign n3692 = ~x185 & ~x537 ;
  assign n3693 = x185 & x537 ;
  assign n3694 = ~n3692 & ~n3693 ;
  assign n3695 = ~n3691 & ~n3694 ;
  assign n3696 = n3691 & n3694 ;
  assign n3697 = ~n3695 & ~n3696 ;
  assign n3698 = ~x187 & ~x539 ;
  assign n3699 = x187 & x539 ;
  assign n3700 = ~n3698 & ~n3699 ;
  assign n3701 = ~x186 & ~x538 ;
  assign n3702 = x186 & x538 ;
  assign n3703 = ~n3701 & ~n3702 ;
  assign n3704 = ~n3700 & ~n3703 ;
  assign n3705 = n3700 & n3703 ;
  assign n3706 = ~n3704 & ~n3705 ;
  assign n3707 = ~x188 & ~x540 ;
  assign n3708 = x188 & x540 ;
  assign n3709 = ~n3707 & ~n3708 ;
  assign n3710 = ~n3706 & ~n3709 ;
  assign n3711 = n3706 & n3709 ;
  assign n3712 = ~n3710 & ~n3711 ;
  assign n3713 = n3697 & ~n3712 ;
  assign n3714 = ~n3695 & ~n3713 ;
  assign n3715 = ~n3683 & ~n3690 ;
  assign n3716 = ~n3714 & n3715 ;
  assign n3717 = n3714 & ~n3715 ;
  assign n3718 = ~n3716 & ~n3717 ;
  assign n3719 = ~n3705 & ~n3711 ;
  assign n3720 = n3718 & n3719 ;
  assign n3721 = ~n3716 & ~n3720 ;
  assign n3722 = ~n3718 & ~n3719 ;
  assign n3723 = ~n3720 & ~n3722 ;
  assign n3724 = ~n3697 & n3712 ;
  assign n3725 = ~n3713 & ~n3724 ;
  assign n3726 = ~x177 & ~x529 ;
  assign n3727 = x177 & x529 ;
  assign n3728 = ~n3726 & ~n3727 ;
  assign n3729 = n3725 & ~n3728 ;
  assign n3730 = ~x183 & ~x535 ;
  assign n3731 = x183 & x535 ;
  assign n3732 = ~n3730 & ~n3731 ;
  assign n3733 = ~x182 & ~x534 ;
  assign n3734 = x182 & x534 ;
  assign n3735 = ~n3733 & ~n3734 ;
  assign n3736 = ~n3732 & ~n3735 ;
  assign n3737 = n3732 & n3735 ;
  assign n3738 = ~n3736 & ~n3737 ;
  assign n3739 = ~x184 & ~x536 ;
  assign n3740 = x184 & x536 ;
  assign n3741 = ~n3739 & ~n3740 ;
  assign n3742 = ~n3738 & ~n3741 ;
  assign n3743 = n3738 & n3741 ;
  assign n3744 = ~n3742 & ~n3743 ;
  assign n3745 = ~x178 & ~x530 ;
  assign n3746 = x178 & x530 ;
  assign n3747 = ~n3745 & ~n3746 ;
  assign n3748 = ~n3744 & ~n3747 ;
  assign n3749 = n3744 & n3747 ;
  assign n3750 = ~n3748 & ~n3749 ;
  assign n3751 = ~x180 & ~x532 ;
  assign n3752 = x180 & x532 ;
  assign n3753 = ~n3751 & ~n3752 ;
  assign n3754 = ~x179 & ~x531 ;
  assign n3755 = x179 & x531 ;
  assign n3756 = ~n3754 & ~n3755 ;
  assign n3757 = ~n3753 & ~n3756 ;
  assign n3758 = n3753 & n3756 ;
  assign n3759 = ~n3757 & ~n3758 ;
  assign n3760 = ~x181 & ~x533 ;
  assign n3761 = x181 & x533 ;
  assign n3762 = ~n3760 & ~n3761 ;
  assign n3763 = ~n3759 & ~n3762 ;
  assign n3764 = n3759 & n3762 ;
  assign n3765 = ~n3763 & ~n3764 ;
  assign n3766 = n3750 & ~n3765 ;
  assign n3767 = ~n3750 & n3765 ;
  assign n3768 = ~n3766 & ~n3767 ;
  assign n3769 = ~n3725 & n3728 ;
  assign n3770 = ~n3729 & ~n3769 ;
  assign n3771 = n3768 & n3770 ;
  assign n3772 = ~n3729 & ~n3771 ;
  assign n3773 = n3723 & ~n3772 ;
  assign n3774 = ~n3748 & ~n3766 ;
  assign n3775 = ~n3737 & ~n3743 ;
  assign n3776 = ~n3774 & n3775 ;
  assign n3777 = n3774 & ~n3775 ;
  assign n3778 = ~n3776 & ~n3777 ;
  assign n3779 = ~n3758 & ~n3764 ;
  assign n3780 = n3778 & n3779 ;
  assign n3781 = ~n3778 & ~n3779 ;
  assign n3782 = ~n3780 & ~n3781 ;
  assign n3783 = ~n3723 & n3772 ;
  assign n3784 = ~n3773 & ~n3783 ;
  assign n3785 = n3782 & n3784 ;
  assign n3786 = ~n3773 & ~n3785 ;
  assign n3787 = ~n3721 & ~n3786 ;
  assign n3788 = n3721 & n3786 ;
  assign n3789 = ~n3787 & ~n3788 ;
  assign n3790 = ~n3776 & ~n3780 ;
  assign n3791 = n3789 & ~n3790 ;
  assign n3792 = ~n3787 & ~n3791 ;
  assign n3793 = ~n3789 & n3790 ;
  assign n3794 = ~n3791 & ~n3793 ;
  assign n3795 = ~n3782 & ~n3784 ;
  assign n3796 = ~n3785 & ~n3795 ;
  assign n3797 = ~n3768 & ~n3770 ;
  assign n3798 = ~n3771 & ~n3797 ;
  assign n3799 = ~x161 & ~x513 ;
  assign n3800 = x161 & x513 ;
  assign n3801 = ~n3799 & ~n3800 ;
  assign n3802 = n3798 & ~n3801 ;
  assign n3803 = ~x168 & ~x520 ;
  assign n3804 = x168 & x520 ;
  assign n3805 = ~n3803 & ~n3804 ;
  assign n3806 = ~x167 & ~x519 ;
  assign n3807 = x167 & x519 ;
  assign n3808 = ~n3806 & ~n3807 ;
  assign n3809 = ~n3805 & ~n3808 ;
  assign n3810 = n3805 & n3808 ;
  assign n3811 = ~n3809 & ~n3810 ;
  assign n3812 = ~x169 & ~x521 ;
  assign n3813 = x169 & x521 ;
  assign n3814 = ~n3812 & ~n3813 ;
  assign n3815 = ~n3811 & ~n3814 ;
  assign n3816 = n3811 & n3814 ;
  assign n3817 = ~n3815 & ~n3816 ;
  assign n3818 = ~x163 & ~x515 ;
  assign n3819 = x163 & x515 ;
  assign n3820 = ~n3818 & ~n3819 ;
  assign n3821 = ~n3817 & ~n3820 ;
  assign n3822 = n3817 & n3820 ;
  assign n3823 = ~n3821 & ~n3822 ;
  assign n3824 = ~x165 & ~x517 ;
  assign n3825 = x165 & x517 ;
  assign n3826 = ~n3824 & ~n3825 ;
  assign n3827 = ~x164 & ~x516 ;
  assign n3828 = x164 & x516 ;
  assign n3829 = ~n3827 & ~n3828 ;
  assign n3830 = ~n3826 & ~n3829 ;
  assign n3831 = n3826 & n3829 ;
  assign n3832 = ~n3830 & ~n3831 ;
  assign n3833 = ~x166 & ~x518 ;
  assign n3834 = x166 & x518 ;
  assign n3835 = ~n3833 & ~n3834 ;
  assign n3836 = ~n3832 & ~n3835 ;
  assign n3837 = n3832 & n3835 ;
  assign n3838 = ~n3836 & ~n3837 ;
  assign n3839 = n3823 & ~n3838 ;
  assign n3840 = ~n3823 & n3838 ;
  assign n3841 = ~n3839 & ~n3840 ;
  assign n3842 = ~x175 & ~x527 ;
  assign n3843 = x175 & x527 ;
  assign n3844 = ~n3842 & ~n3843 ;
  assign n3845 = ~x174 & ~x526 ;
  assign n3846 = x174 & x526 ;
  assign n3847 = ~n3845 & ~n3846 ;
  assign n3848 = ~n3844 & ~n3847 ;
  assign n3849 = n3844 & n3847 ;
  assign n3850 = ~n3848 & ~n3849 ;
  assign n3851 = ~x176 & ~x528 ;
  assign n3852 = x176 & x528 ;
  assign n3853 = ~n3851 & ~n3852 ;
  assign n3854 = ~n3850 & ~n3853 ;
  assign n3855 = n3850 & n3853 ;
  assign n3856 = ~n3854 & ~n3855 ;
  assign n3857 = ~x170 & ~x522 ;
  assign n3858 = x170 & x522 ;
  assign n3859 = ~n3857 & ~n3858 ;
  assign n3860 = ~n3856 & ~n3859 ;
  assign n3861 = n3856 & n3859 ;
  assign n3862 = ~n3860 & ~n3861 ;
  assign n3863 = ~x172 & ~x524 ;
  assign n3864 = x172 & x524 ;
  assign n3865 = ~n3863 & ~n3864 ;
  assign n3866 = ~x171 & ~x523 ;
  assign n3867 = x171 & x523 ;
  assign n3868 = ~n3866 & ~n3867 ;
  assign n3869 = ~n3865 & ~n3868 ;
  assign n3870 = n3865 & n3868 ;
  assign n3871 = ~n3869 & ~n3870 ;
  assign n3872 = ~x173 & ~x525 ;
  assign n3873 = x173 & x525 ;
  assign n3874 = ~n3872 & ~n3873 ;
  assign n3875 = ~n3871 & ~n3874 ;
  assign n3876 = n3871 & n3874 ;
  assign n3877 = ~n3875 & ~n3876 ;
  assign n3878 = n3862 & ~n3877 ;
  assign n3879 = ~n3862 & n3877 ;
  assign n3880 = ~n3878 & ~n3879 ;
  assign n3881 = ~x162 & ~x514 ;
  assign n3882 = x162 & x514 ;
  assign n3883 = ~n3881 & ~n3882 ;
  assign n3884 = n3880 & ~n3883 ;
  assign n3885 = ~n3880 & n3883 ;
  assign n3886 = ~n3884 & ~n3885 ;
  assign n3887 = n3841 & n3886 ;
  assign n3888 = ~n3841 & ~n3886 ;
  assign n3889 = ~n3887 & ~n3888 ;
  assign n3890 = ~n3798 & n3801 ;
  assign n3891 = ~n3802 & ~n3890 ;
  assign n3892 = n3889 & n3891 ;
  assign n3893 = ~n3802 & ~n3892 ;
  assign n3894 = n3796 & ~n3893 ;
  assign n3895 = ~n3821 & ~n3839 ;
  assign n3896 = ~n3810 & ~n3816 ;
  assign n3897 = ~n3895 & n3896 ;
  assign n3898 = n3895 & ~n3896 ;
  assign n3899 = ~n3897 & ~n3898 ;
  assign n3900 = ~n3831 & ~n3837 ;
  assign n3901 = n3899 & n3900 ;
  assign n3902 = ~n3899 & ~n3900 ;
  assign n3903 = ~n3901 & ~n3902 ;
  assign n3904 = ~n3860 & ~n3878 ;
  assign n3905 = ~n3849 & ~n3855 ;
  assign n3906 = ~n3904 & n3905 ;
  assign n3907 = n3904 & ~n3905 ;
  assign n3908 = ~n3906 & ~n3907 ;
  assign n3909 = ~n3870 & ~n3876 ;
  assign n3910 = n3908 & n3909 ;
  assign n3911 = ~n3908 & ~n3909 ;
  assign n3912 = ~n3910 & ~n3911 ;
  assign n3913 = ~n3884 & ~n3887 ;
  assign n3914 = n3912 & ~n3913 ;
  assign n3915 = ~n3912 & n3913 ;
  assign n3916 = ~n3914 & ~n3915 ;
  assign n3917 = n3903 & n3916 ;
  assign n3918 = ~n3903 & ~n3916 ;
  assign n3919 = ~n3917 & ~n3918 ;
  assign n3920 = ~n3796 & n3893 ;
  assign n3921 = ~n3894 & ~n3920 ;
  assign n3922 = n3919 & n3921 ;
  assign n3923 = ~n3894 & ~n3922 ;
  assign n3924 = n3794 & ~n3923 ;
  assign n3925 = ~n3906 & ~n3910 ;
  assign n3926 = ~n3914 & ~n3917 ;
  assign n3927 = ~n3925 & ~n3926 ;
  assign n3928 = n3925 & n3926 ;
  assign n3929 = ~n3927 & ~n3928 ;
  assign n3930 = ~n3897 & ~n3901 ;
  assign n3931 = n3929 & ~n3930 ;
  assign n3932 = ~n3929 & n3930 ;
  assign n3933 = ~n3931 & ~n3932 ;
  assign n3934 = ~n3794 & n3923 ;
  assign n3935 = ~n3924 & ~n3934 ;
  assign n3936 = n3933 & n3935 ;
  assign n3937 = ~n3924 & ~n3936 ;
  assign n3938 = ~n3792 & ~n3937 ;
  assign n3939 = n3792 & n3937 ;
  assign n3940 = ~n3938 & ~n3939 ;
  assign n3941 = ~n3927 & ~n3931 ;
  assign n3942 = n3940 & ~n3941 ;
  assign n3943 = ~n3938 & ~n3942 ;
  assign n3944 = ~n3940 & n3941 ;
  assign n3945 = ~n3942 & ~n3944 ;
  assign n3946 = ~n3933 & ~n3935 ;
  assign n3947 = ~n3936 & ~n3946 ;
  assign n3948 = ~n3919 & ~n3921 ;
  assign n3949 = ~n3922 & ~n3948 ;
  assign n3950 = ~n3889 & ~n3891 ;
  assign n3951 = ~n3892 & ~n3950 ;
  assign n3952 = ~x160 & ~x512 ;
  assign n3953 = x160 & x512 ;
  assign n3954 = ~n3952 & ~n3953 ;
  assign n3955 = ~n3951 & n3954 ;
  assign n3956 = ~n3949 & n3955 ;
  assign n3957 = ~n3947 & n3956 ;
  assign n3958 = ~n3945 & n3957 ;
  assign n3959 = n3943 & n3958 ;
  assign n3960 = n3676 & n3959 ;
  assign n3961 = ~x158 & ~x542 ;
  assign n3962 = x158 & x542 ;
  assign n3963 = ~n3961 & ~n3962 ;
  assign n3964 = ~x157 & ~x541 ;
  assign n3965 = x157 & x541 ;
  assign n3966 = ~n3964 & ~n3965 ;
  assign n3967 = n3963 & n3966 ;
  assign n3968 = ~n3963 & ~n3966 ;
  assign n3969 = ~n3967 & ~n3968 ;
  assign n3970 = ~x159 & ~x543 ;
  assign n3971 = x159 & x543 ;
  assign n3972 = ~n3970 & ~n3971 ;
  assign n3973 = ~n3969 & ~n3972 ;
  assign n3974 = n3969 & n3972 ;
  assign n3975 = ~n3973 & ~n3974 ;
  assign n3976 = ~x153 & ~x537 ;
  assign n3977 = x153 & x537 ;
  assign n3978 = ~n3976 & ~n3977 ;
  assign n3979 = ~n3975 & ~n3978 ;
  assign n3980 = n3975 & n3978 ;
  assign n3981 = ~n3979 & ~n3980 ;
  assign n3982 = ~x155 & ~x539 ;
  assign n3983 = x155 & x539 ;
  assign n3984 = ~n3982 & ~n3983 ;
  assign n3985 = ~x154 & ~x538 ;
  assign n3986 = x154 & x538 ;
  assign n3987 = ~n3985 & ~n3986 ;
  assign n3988 = ~n3984 & ~n3987 ;
  assign n3989 = n3984 & n3987 ;
  assign n3990 = ~n3988 & ~n3989 ;
  assign n3991 = ~x156 & ~x540 ;
  assign n3992 = x156 & x540 ;
  assign n3993 = ~n3991 & ~n3992 ;
  assign n3994 = ~n3990 & ~n3993 ;
  assign n3995 = n3990 & n3993 ;
  assign n3996 = ~n3994 & ~n3995 ;
  assign n3997 = n3981 & ~n3996 ;
  assign n3998 = ~n3979 & ~n3997 ;
  assign n3999 = ~n3967 & ~n3974 ;
  assign n4000 = ~n3998 & n3999 ;
  assign n4001 = n3998 & ~n3999 ;
  assign n4002 = ~n4000 & ~n4001 ;
  assign n4003 = ~n3989 & ~n3995 ;
  assign n4004 = n4002 & n4003 ;
  assign n4005 = ~n4000 & ~n4004 ;
  assign n4006 = ~n4002 & ~n4003 ;
  assign n4007 = ~n4004 & ~n4006 ;
  assign n4008 = ~n3981 & n3996 ;
  assign n4009 = ~n3997 & ~n4008 ;
  assign n4010 = ~x145 & ~x529 ;
  assign n4011 = x145 & x529 ;
  assign n4012 = ~n4010 & ~n4011 ;
  assign n4013 = n4009 & ~n4012 ;
  assign n4014 = ~x151 & ~x535 ;
  assign n4015 = x151 & x535 ;
  assign n4016 = ~n4014 & ~n4015 ;
  assign n4017 = ~x150 & ~x534 ;
  assign n4018 = x150 & x534 ;
  assign n4019 = ~n4017 & ~n4018 ;
  assign n4020 = ~n4016 & ~n4019 ;
  assign n4021 = n4016 & n4019 ;
  assign n4022 = ~n4020 & ~n4021 ;
  assign n4023 = ~x152 & ~x536 ;
  assign n4024 = x152 & x536 ;
  assign n4025 = ~n4023 & ~n4024 ;
  assign n4026 = ~n4022 & ~n4025 ;
  assign n4027 = n4022 & n4025 ;
  assign n4028 = ~n4026 & ~n4027 ;
  assign n4029 = ~x146 & ~x530 ;
  assign n4030 = x146 & x530 ;
  assign n4031 = ~n4029 & ~n4030 ;
  assign n4032 = ~n4028 & ~n4031 ;
  assign n4033 = n4028 & n4031 ;
  assign n4034 = ~n4032 & ~n4033 ;
  assign n4035 = ~x148 & ~x532 ;
  assign n4036 = x148 & x532 ;
  assign n4037 = ~n4035 & ~n4036 ;
  assign n4038 = ~x147 & ~x531 ;
  assign n4039 = x147 & x531 ;
  assign n4040 = ~n4038 & ~n4039 ;
  assign n4041 = ~n4037 & ~n4040 ;
  assign n4042 = n4037 & n4040 ;
  assign n4043 = ~n4041 & ~n4042 ;
  assign n4044 = ~x149 & ~x533 ;
  assign n4045 = x149 & x533 ;
  assign n4046 = ~n4044 & ~n4045 ;
  assign n4047 = ~n4043 & ~n4046 ;
  assign n4048 = n4043 & n4046 ;
  assign n4049 = ~n4047 & ~n4048 ;
  assign n4050 = n4034 & ~n4049 ;
  assign n4051 = ~n4034 & n4049 ;
  assign n4052 = ~n4050 & ~n4051 ;
  assign n4053 = ~n4009 & n4012 ;
  assign n4054 = ~n4013 & ~n4053 ;
  assign n4055 = n4052 & n4054 ;
  assign n4056 = ~n4013 & ~n4055 ;
  assign n4057 = n4007 & ~n4056 ;
  assign n4058 = ~n4032 & ~n4050 ;
  assign n4059 = ~n4021 & ~n4027 ;
  assign n4060 = ~n4058 & n4059 ;
  assign n4061 = n4058 & ~n4059 ;
  assign n4062 = ~n4060 & ~n4061 ;
  assign n4063 = ~n4042 & ~n4048 ;
  assign n4064 = n4062 & n4063 ;
  assign n4065 = ~n4062 & ~n4063 ;
  assign n4066 = ~n4064 & ~n4065 ;
  assign n4067 = ~n4007 & n4056 ;
  assign n4068 = ~n4057 & ~n4067 ;
  assign n4069 = n4066 & n4068 ;
  assign n4070 = ~n4057 & ~n4069 ;
  assign n4071 = ~n4005 & ~n4070 ;
  assign n4072 = n4005 & n4070 ;
  assign n4073 = ~n4071 & ~n4072 ;
  assign n4074 = ~n4060 & ~n4064 ;
  assign n4075 = n4073 & ~n4074 ;
  assign n4076 = ~n4071 & ~n4075 ;
  assign n4077 = ~n4073 & n4074 ;
  assign n4078 = ~n4075 & ~n4077 ;
  assign n4079 = ~n4066 & ~n4068 ;
  assign n4080 = ~n4069 & ~n4079 ;
  assign n4081 = ~n4052 & ~n4054 ;
  assign n4082 = ~n4055 & ~n4081 ;
  assign n4083 = ~x129 & ~x513 ;
  assign n4084 = x129 & x513 ;
  assign n4085 = ~n4083 & ~n4084 ;
  assign n4086 = n4082 & ~n4085 ;
  assign n4087 = ~x136 & ~x520 ;
  assign n4088 = x136 & x520 ;
  assign n4089 = ~n4087 & ~n4088 ;
  assign n4090 = ~x135 & ~x519 ;
  assign n4091 = x135 & x519 ;
  assign n4092 = ~n4090 & ~n4091 ;
  assign n4093 = ~n4089 & ~n4092 ;
  assign n4094 = n4089 & n4092 ;
  assign n4095 = ~n4093 & ~n4094 ;
  assign n4096 = ~x137 & ~x521 ;
  assign n4097 = x137 & x521 ;
  assign n4098 = ~n4096 & ~n4097 ;
  assign n4099 = ~n4095 & ~n4098 ;
  assign n4100 = n4095 & n4098 ;
  assign n4101 = ~n4099 & ~n4100 ;
  assign n4102 = ~x131 & ~x515 ;
  assign n4103 = x131 & x515 ;
  assign n4104 = ~n4102 & ~n4103 ;
  assign n4105 = ~n4101 & ~n4104 ;
  assign n4106 = n4101 & n4104 ;
  assign n4107 = ~n4105 & ~n4106 ;
  assign n4108 = ~x133 & ~x517 ;
  assign n4109 = x133 & x517 ;
  assign n4110 = ~n4108 & ~n4109 ;
  assign n4111 = ~x132 & ~x516 ;
  assign n4112 = x132 & x516 ;
  assign n4113 = ~n4111 & ~n4112 ;
  assign n4114 = ~n4110 & ~n4113 ;
  assign n4115 = n4110 & n4113 ;
  assign n4116 = ~n4114 & ~n4115 ;
  assign n4117 = ~x134 & ~x518 ;
  assign n4118 = x134 & x518 ;
  assign n4119 = ~n4117 & ~n4118 ;
  assign n4120 = ~n4116 & ~n4119 ;
  assign n4121 = n4116 & n4119 ;
  assign n4122 = ~n4120 & ~n4121 ;
  assign n4123 = n4107 & ~n4122 ;
  assign n4124 = ~n4107 & n4122 ;
  assign n4125 = ~n4123 & ~n4124 ;
  assign n4126 = ~x143 & ~x527 ;
  assign n4127 = x143 & x527 ;
  assign n4128 = ~n4126 & ~n4127 ;
  assign n4129 = ~x142 & ~x526 ;
  assign n4130 = x142 & x526 ;
  assign n4131 = ~n4129 & ~n4130 ;
  assign n4132 = ~n4128 & ~n4131 ;
  assign n4133 = n4128 & n4131 ;
  assign n4134 = ~n4132 & ~n4133 ;
  assign n4135 = ~x144 & ~x528 ;
  assign n4136 = x144 & x528 ;
  assign n4137 = ~n4135 & ~n4136 ;
  assign n4138 = ~n4134 & ~n4137 ;
  assign n4139 = n4134 & n4137 ;
  assign n4140 = ~n4138 & ~n4139 ;
  assign n4141 = ~x138 & ~x522 ;
  assign n4142 = x138 & x522 ;
  assign n4143 = ~n4141 & ~n4142 ;
  assign n4144 = ~n4140 & ~n4143 ;
  assign n4145 = n4140 & n4143 ;
  assign n4146 = ~n4144 & ~n4145 ;
  assign n4147 = ~x140 & ~x524 ;
  assign n4148 = x140 & x524 ;
  assign n4149 = ~n4147 & ~n4148 ;
  assign n4150 = ~x139 & ~x523 ;
  assign n4151 = x139 & x523 ;
  assign n4152 = ~n4150 & ~n4151 ;
  assign n4153 = ~n4149 & ~n4152 ;
  assign n4154 = n4149 & n4152 ;
  assign n4155 = ~n4153 & ~n4154 ;
  assign n4156 = ~x141 & ~x525 ;
  assign n4157 = x141 & x525 ;
  assign n4158 = ~n4156 & ~n4157 ;
  assign n4159 = ~n4155 & ~n4158 ;
  assign n4160 = n4155 & n4158 ;
  assign n4161 = ~n4159 & ~n4160 ;
  assign n4162 = n4146 & ~n4161 ;
  assign n4163 = ~n4146 & n4161 ;
  assign n4164 = ~n4162 & ~n4163 ;
  assign n4165 = ~x130 & ~x514 ;
  assign n4166 = x130 & x514 ;
  assign n4167 = ~n4165 & ~n4166 ;
  assign n4168 = n4164 & ~n4167 ;
  assign n4169 = ~n4164 & n4167 ;
  assign n4170 = ~n4168 & ~n4169 ;
  assign n4171 = n4125 & n4170 ;
  assign n4172 = ~n4125 & ~n4170 ;
  assign n4173 = ~n4171 & ~n4172 ;
  assign n4174 = ~n4082 & n4085 ;
  assign n4175 = ~n4086 & ~n4174 ;
  assign n4176 = n4173 & n4175 ;
  assign n4177 = ~n4086 & ~n4176 ;
  assign n4178 = n4080 & ~n4177 ;
  assign n4179 = ~n4105 & ~n4123 ;
  assign n4180 = ~n4094 & ~n4100 ;
  assign n4181 = ~n4179 & n4180 ;
  assign n4182 = n4179 & ~n4180 ;
  assign n4183 = ~n4181 & ~n4182 ;
  assign n4184 = ~n4115 & ~n4121 ;
  assign n4185 = n4183 & n4184 ;
  assign n4186 = ~n4183 & ~n4184 ;
  assign n4187 = ~n4185 & ~n4186 ;
  assign n4188 = ~n4144 & ~n4162 ;
  assign n4189 = ~n4133 & ~n4139 ;
  assign n4190 = ~n4188 & n4189 ;
  assign n4191 = n4188 & ~n4189 ;
  assign n4192 = ~n4190 & ~n4191 ;
  assign n4193 = ~n4154 & ~n4160 ;
  assign n4194 = n4192 & n4193 ;
  assign n4195 = ~n4192 & ~n4193 ;
  assign n4196 = ~n4194 & ~n4195 ;
  assign n4197 = ~n4168 & ~n4171 ;
  assign n4198 = n4196 & ~n4197 ;
  assign n4199 = ~n4196 & n4197 ;
  assign n4200 = ~n4198 & ~n4199 ;
  assign n4201 = n4187 & n4200 ;
  assign n4202 = ~n4187 & ~n4200 ;
  assign n4203 = ~n4201 & ~n4202 ;
  assign n4204 = ~n4080 & n4177 ;
  assign n4205 = ~n4178 & ~n4204 ;
  assign n4206 = n4203 & n4205 ;
  assign n4207 = ~n4178 & ~n4206 ;
  assign n4208 = n4078 & ~n4207 ;
  assign n4209 = ~n4190 & ~n4194 ;
  assign n4210 = ~n4198 & ~n4201 ;
  assign n4211 = ~n4209 & ~n4210 ;
  assign n4212 = n4209 & n4210 ;
  assign n4213 = ~n4211 & ~n4212 ;
  assign n4214 = ~n4181 & ~n4185 ;
  assign n4215 = n4213 & ~n4214 ;
  assign n4216 = ~n4213 & n4214 ;
  assign n4217 = ~n4215 & ~n4216 ;
  assign n4218 = ~n4078 & n4207 ;
  assign n4219 = ~n4208 & ~n4218 ;
  assign n4220 = n4217 & n4219 ;
  assign n4221 = ~n4208 & ~n4220 ;
  assign n4222 = ~n4076 & ~n4221 ;
  assign n4223 = n4076 & n4221 ;
  assign n4224 = ~n4222 & ~n4223 ;
  assign n4225 = ~n4211 & ~n4215 ;
  assign n4226 = n4224 & ~n4225 ;
  assign n4227 = ~n4222 & ~n4226 ;
  assign n4228 = ~n4224 & n4225 ;
  assign n4229 = ~n4226 & ~n4228 ;
  assign n4230 = ~n4217 & ~n4219 ;
  assign n4231 = ~n4220 & ~n4230 ;
  assign n4232 = ~n4203 & ~n4205 ;
  assign n4233 = ~n4206 & ~n4232 ;
  assign n4234 = ~n4173 & ~n4175 ;
  assign n4235 = ~n4176 & ~n4234 ;
  assign n4236 = ~x128 & ~x512 ;
  assign n4237 = x128 & x512 ;
  assign n4238 = ~n4236 & ~n4237 ;
  assign n4239 = ~n4235 & n4238 ;
  assign n4240 = ~n4233 & n4239 ;
  assign n4241 = ~n4231 & n4240 ;
  assign n4242 = ~n4229 & n4241 ;
  assign n4243 = n4227 & n4242 ;
  assign n4244 = n3960 & n4243 ;
  assign n4245 = ~x126 & ~x542 ;
  assign n4246 = x126 & x542 ;
  assign n4247 = ~n4245 & ~n4246 ;
  assign n4248 = ~x125 & ~x541 ;
  assign n4249 = x125 & x541 ;
  assign n4250 = ~n4248 & ~n4249 ;
  assign n4251 = n4247 & n4250 ;
  assign n4252 = ~n4247 & ~n4250 ;
  assign n4253 = ~n4251 & ~n4252 ;
  assign n4254 = ~x127 & ~x543 ;
  assign n4255 = x127 & x543 ;
  assign n4256 = ~n4254 & ~n4255 ;
  assign n4257 = ~n4253 & ~n4256 ;
  assign n4258 = n4253 & n4256 ;
  assign n4259 = ~n4257 & ~n4258 ;
  assign n4260 = ~x121 & ~x537 ;
  assign n4261 = x121 & x537 ;
  assign n4262 = ~n4260 & ~n4261 ;
  assign n4263 = ~n4259 & ~n4262 ;
  assign n4264 = n4259 & n4262 ;
  assign n4265 = ~n4263 & ~n4264 ;
  assign n4266 = ~x123 & ~x539 ;
  assign n4267 = x123 & x539 ;
  assign n4268 = ~n4266 & ~n4267 ;
  assign n4269 = ~x122 & ~x538 ;
  assign n4270 = x122 & x538 ;
  assign n4271 = ~n4269 & ~n4270 ;
  assign n4272 = ~n4268 & ~n4271 ;
  assign n4273 = n4268 & n4271 ;
  assign n4274 = ~n4272 & ~n4273 ;
  assign n4275 = ~x124 & ~x540 ;
  assign n4276 = x124 & x540 ;
  assign n4277 = ~n4275 & ~n4276 ;
  assign n4278 = ~n4274 & ~n4277 ;
  assign n4279 = n4274 & n4277 ;
  assign n4280 = ~n4278 & ~n4279 ;
  assign n4281 = n4265 & ~n4280 ;
  assign n4282 = ~n4263 & ~n4281 ;
  assign n4283 = ~n4251 & ~n4258 ;
  assign n4284 = ~n4282 & n4283 ;
  assign n4285 = n4282 & ~n4283 ;
  assign n4286 = ~n4284 & ~n4285 ;
  assign n4287 = ~n4273 & ~n4279 ;
  assign n4288 = n4286 & n4287 ;
  assign n4289 = ~n4284 & ~n4288 ;
  assign n4290 = ~n4286 & ~n4287 ;
  assign n4291 = ~n4288 & ~n4290 ;
  assign n4292 = ~n4265 & n4280 ;
  assign n4293 = ~n4281 & ~n4292 ;
  assign n4294 = ~x113 & ~x529 ;
  assign n4295 = x113 & x529 ;
  assign n4296 = ~n4294 & ~n4295 ;
  assign n4297 = n4293 & ~n4296 ;
  assign n4298 = ~x119 & ~x535 ;
  assign n4299 = x119 & x535 ;
  assign n4300 = ~n4298 & ~n4299 ;
  assign n4301 = ~x118 & ~x534 ;
  assign n4302 = x118 & x534 ;
  assign n4303 = ~n4301 & ~n4302 ;
  assign n4304 = ~n4300 & ~n4303 ;
  assign n4305 = n4300 & n4303 ;
  assign n4306 = ~n4304 & ~n4305 ;
  assign n4307 = ~x120 & ~x536 ;
  assign n4308 = x120 & x536 ;
  assign n4309 = ~n4307 & ~n4308 ;
  assign n4310 = ~n4306 & ~n4309 ;
  assign n4311 = n4306 & n4309 ;
  assign n4312 = ~n4310 & ~n4311 ;
  assign n4313 = ~x114 & ~x530 ;
  assign n4314 = x114 & x530 ;
  assign n4315 = ~n4313 & ~n4314 ;
  assign n4316 = ~n4312 & ~n4315 ;
  assign n4317 = n4312 & n4315 ;
  assign n4318 = ~n4316 & ~n4317 ;
  assign n4319 = ~x116 & ~x532 ;
  assign n4320 = x116 & x532 ;
  assign n4321 = ~n4319 & ~n4320 ;
  assign n4322 = ~x115 & ~x531 ;
  assign n4323 = x115 & x531 ;
  assign n4324 = ~n4322 & ~n4323 ;
  assign n4325 = ~n4321 & ~n4324 ;
  assign n4326 = n4321 & n4324 ;
  assign n4327 = ~n4325 & ~n4326 ;
  assign n4328 = ~x117 & ~x533 ;
  assign n4329 = x117 & x533 ;
  assign n4330 = ~n4328 & ~n4329 ;
  assign n4331 = ~n4327 & ~n4330 ;
  assign n4332 = n4327 & n4330 ;
  assign n4333 = ~n4331 & ~n4332 ;
  assign n4334 = n4318 & ~n4333 ;
  assign n4335 = ~n4318 & n4333 ;
  assign n4336 = ~n4334 & ~n4335 ;
  assign n4337 = ~n4293 & n4296 ;
  assign n4338 = ~n4297 & ~n4337 ;
  assign n4339 = n4336 & n4338 ;
  assign n4340 = ~n4297 & ~n4339 ;
  assign n4341 = n4291 & ~n4340 ;
  assign n4342 = ~n4316 & ~n4334 ;
  assign n4343 = ~n4305 & ~n4311 ;
  assign n4344 = ~n4342 & n4343 ;
  assign n4345 = n4342 & ~n4343 ;
  assign n4346 = ~n4344 & ~n4345 ;
  assign n4347 = ~n4326 & ~n4332 ;
  assign n4348 = n4346 & n4347 ;
  assign n4349 = ~n4346 & ~n4347 ;
  assign n4350 = ~n4348 & ~n4349 ;
  assign n4351 = ~n4291 & n4340 ;
  assign n4352 = ~n4341 & ~n4351 ;
  assign n4353 = n4350 & n4352 ;
  assign n4354 = ~n4341 & ~n4353 ;
  assign n4355 = ~n4289 & ~n4354 ;
  assign n4356 = n4289 & n4354 ;
  assign n4357 = ~n4355 & ~n4356 ;
  assign n4358 = ~n4344 & ~n4348 ;
  assign n4359 = n4357 & ~n4358 ;
  assign n4360 = ~n4355 & ~n4359 ;
  assign n4361 = ~n4357 & n4358 ;
  assign n4362 = ~n4359 & ~n4361 ;
  assign n4363 = ~n4350 & ~n4352 ;
  assign n4364 = ~n4353 & ~n4363 ;
  assign n4365 = ~n4336 & ~n4338 ;
  assign n4366 = ~n4339 & ~n4365 ;
  assign n4367 = ~x97 & ~x513 ;
  assign n4368 = x97 & x513 ;
  assign n4369 = ~n4367 & ~n4368 ;
  assign n4370 = n4366 & ~n4369 ;
  assign n4371 = ~x104 & ~x520 ;
  assign n4372 = x104 & x520 ;
  assign n4373 = ~n4371 & ~n4372 ;
  assign n4374 = ~x103 & ~x519 ;
  assign n4375 = x103 & x519 ;
  assign n4376 = ~n4374 & ~n4375 ;
  assign n4377 = ~n4373 & ~n4376 ;
  assign n4378 = n4373 & n4376 ;
  assign n4379 = ~n4377 & ~n4378 ;
  assign n4380 = ~x105 & ~x521 ;
  assign n4381 = x105 & x521 ;
  assign n4382 = ~n4380 & ~n4381 ;
  assign n4383 = ~n4379 & ~n4382 ;
  assign n4384 = n4379 & n4382 ;
  assign n4385 = ~n4383 & ~n4384 ;
  assign n4386 = ~x99 & ~x515 ;
  assign n4387 = x99 & x515 ;
  assign n4388 = ~n4386 & ~n4387 ;
  assign n4389 = ~n4385 & ~n4388 ;
  assign n4390 = n4385 & n4388 ;
  assign n4391 = ~n4389 & ~n4390 ;
  assign n4392 = ~x101 & ~x517 ;
  assign n4393 = x101 & x517 ;
  assign n4394 = ~n4392 & ~n4393 ;
  assign n4395 = ~x100 & ~x516 ;
  assign n4396 = x100 & x516 ;
  assign n4397 = ~n4395 & ~n4396 ;
  assign n4398 = ~n4394 & ~n4397 ;
  assign n4399 = n4394 & n4397 ;
  assign n4400 = ~n4398 & ~n4399 ;
  assign n4401 = ~x102 & ~x518 ;
  assign n4402 = x102 & x518 ;
  assign n4403 = ~n4401 & ~n4402 ;
  assign n4404 = ~n4400 & ~n4403 ;
  assign n4405 = n4400 & n4403 ;
  assign n4406 = ~n4404 & ~n4405 ;
  assign n4407 = n4391 & ~n4406 ;
  assign n4408 = ~n4391 & n4406 ;
  assign n4409 = ~n4407 & ~n4408 ;
  assign n4410 = ~x111 & ~x527 ;
  assign n4411 = x111 & x527 ;
  assign n4412 = ~n4410 & ~n4411 ;
  assign n4413 = ~x110 & ~x526 ;
  assign n4414 = x110 & x526 ;
  assign n4415 = ~n4413 & ~n4414 ;
  assign n4416 = ~n4412 & ~n4415 ;
  assign n4417 = n4412 & n4415 ;
  assign n4418 = ~n4416 & ~n4417 ;
  assign n4419 = ~x112 & ~x528 ;
  assign n4420 = x112 & x528 ;
  assign n4421 = ~n4419 & ~n4420 ;
  assign n4422 = ~n4418 & ~n4421 ;
  assign n4423 = n4418 & n4421 ;
  assign n4424 = ~n4422 & ~n4423 ;
  assign n4425 = ~x106 & ~x522 ;
  assign n4426 = x106 & x522 ;
  assign n4427 = ~n4425 & ~n4426 ;
  assign n4428 = ~n4424 & ~n4427 ;
  assign n4429 = n4424 & n4427 ;
  assign n4430 = ~n4428 & ~n4429 ;
  assign n4431 = ~x108 & ~x524 ;
  assign n4432 = x108 & x524 ;
  assign n4433 = ~n4431 & ~n4432 ;
  assign n4434 = ~x107 & ~x523 ;
  assign n4435 = x107 & x523 ;
  assign n4436 = ~n4434 & ~n4435 ;
  assign n4437 = ~n4433 & ~n4436 ;
  assign n4438 = n4433 & n4436 ;
  assign n4439 = ~n4437 & ~n4438 ;
  assign n4440 = ~x109 & ~x525 ;
  assign n4441 = x109 & x525 ;
  assign n4442 = ~n4440 & ~n4441 ;
  assign n4443 = ~n4439 & ~n4442 ;
  assign n4444 = n4439 & n4442 ;
  assign n4445 = ~n4443 & ~n4444 ;
  assign n4446 = n4430 & ~n4445 ;
  assign n4447 = ~n4430 & n4445 ;
  assign n4448 = ~n4446 & ~n4447 ;
  assign n4449 = ~x98 & ~x514 ;
  assign n4450 = x98 & x514 ;
  assign n4451 = ~n4449 & ~n4450 ;
  assign n4452 = n4448 & ~n4451 ;
  assign n4453 = ~n4448 & n4451 ;
  assign n4454 = ~n4452 & ~n4453 ;
  assign n4455 = n4409 & n4454 ;
  assign n4456 = ~n4409 & ~n4454 ;
  assign n4457 = ~n4455 & ~n4456 ;
  assign n4458 = ~n4366 & n4369 ;
  assign n4459 = ~n4370 & ~n4458 ;
  assign n4460 = n4457 & n4459 ;
  assign n4461 = ~n4370 & ~n4460 ;
  assign n4462 = n4364 & ~n4461 ;
  assign n4463 = ~n4389 & ~n4407 ;
  assign n4464 = ~n4378 & ~n4384 ;
  assign n4465 = ~n4463 & n4464 ;
  assign n4466 = n4463 & ~n4464 ;
  assign n4467 = ~n4465 & ~n4466 ;
  assign n4468 = ~n4399 & ~n4405 ;
  assign n4469 = n4467 & n4468 ;
  assign n4470 = ~n4467 & ~n4468 ;
  assign n4471 = ~n4469 & ~n4470 ;
  assign n4472 = ~n4428 & ~n4446 ;
  assign n4473 = ~n4417 & ~n4423 ;
  assign n4474 = ~n4472 & n4473 ;
  assign n4475 = n4472 & ~n4473 ;
  assign n4476 = ~n4474 & ~n4475 ;
  assign n4477 = ~n4438 & ~n4444 ;
  assign n4478 = n4476 & n4477 ;
  assign n4479 = ~n4476 & ~n4477 ;
  assign n4480 = ~n4478 & ~n4479 ;
  assign n4481 = ~n4452 & ~n4455 ;
  assign n4482 = n4480 & ~n4481 ;
  assign n4483 = ~n4480 & n4481 ;
  assign n4484 = ~n4482 & ~n4483 ;
  assign n4485 = n4471 & n4484 ;
  assign n4486 = ~n4471 & ~n4484 ;
  assign n4487 = ~n4485 & ~n4486 ;
  assign n4488 = ~n4364 & n4461 ;
  assign n4489 = ~n4462 & ~n4488 ;
  assign n4490 = n4487 & n4489 ;
  assign n4491 = ~n4462 & ~n4490 ;
  assign n4492 = n4362 & ~n4491 ;
  assign n4493 = ~n4474 & ~n4478 ;
  assign n4494 = ~n4482 & ~n4485 ;
  assign n4495 = ~n4493 & ~n4494 ;
  assign n4496 = n4493 & n4494 ;
  assign n4497 = ~n4495 & ~n4496 ;
  assign n4498 = ~n4465 & ~n4469 ;
  assign n4499 = n4497 & ~n4498 ;
  assign n4500 = ~n4497 & n4498 ;
  assign n4501 = ~n4499 & ~n4500 ;
  assign n4502 = ~n4362 & n4491 ;
  assign n4503 = ~n4492 & ~n4502 ;
  assign n4504 = n4501 & n4503 ;
  assign n4505 = ~n4492 & ~n4504 ;
  assign n4506 = ~n4360 & ~n4505 ;
  assign n4507 = n4360 & n4505 ;
  assign n4508 = ~n4506 & ~n4507 ;
  assign n4509 = ~n4495 & ~n4499 ;
  assign n4510 = n4508 & ~n4509 ;
  assign n4511 = ~n4506 & ~n4510 ;
  assign n4512 = ~n4508 & n4509 ;
  assign n4513 = ~n4510 & ~n4512 ;
  assign n4514 = ~n4501 & ~n4503 ;
  assign n4515 = ~n4504 & ~n4514 ;
  assign n4516 = ~n4487 & ~n4489 ;
  assign n4517 = ~n4490 & ~n4516 ;
  assign n4518 = ~n4457 & ~n4459 ;
  assign n4519 = ~n4460 & ~n4518 ;
  assign n4520 = ~x96 & ~x512 ;
  assign n4521 = x96 & x512 ;
  assign n4522 = ~n4520 & ~n4521 ;
  assign n4523 = ~n4519 & n4522 ;
  assign n4524 = ~n4517 & n4523 ;
  assign n4525 = ~n4515 & n4524 ;
  assign n4526 = ~n4513 & n4525 ;
  assign n4527 = n4511 & n4526 ;
  assign n4528 = n4244 & n4527 ;
  assign n4529 = ~x94 & ~x542 ;
  assign n4530 = x94 & x542 ;
  assign n4531 = ~n4529 & ~n4530 ;
  assign n4532 = ~x93 & ~x541 ;
  assign n4533 = x93 & x541 ;
  assign n4534 = ~n4532 & ~n4533 ;
  assign n4535 = n4531 & n4534 ;
  assign n4536 = ~n4531 & ~n4534 ;
  assign n4537 = ~n4535 & ~n4536 ;
  assign n4538 = ~x95 & ~x543 ;
  assign n4539 = x95 & x543 ;
  assign n4540 = ~n4538 & ~n4539 ;
  assign n4541 = ~n4537 & ~n4540 ;
  assign n4542 = n4537 & n4540 ;
  assign n4543 = ~n4541 & ~n4542 ;
  assign n4544 = ~x89 & ~x537 ;
  assign n4545 = x89 & x537 ;
  assign n4546 = ~n4544 & ~n4545 ;
  assign n4547 = ~n4543 & ~n4546 ;
  assign n4548 = n4543 & n4546 ;
  assign n4549 = ~n4547 & ~n4548 ;
  assign n4550 = ~x91 & ~x539 ;
  assign n4551 = x91 & x539 ;
  assign n4552 = ~n4550 & ~n4551 ;
  assign n4553 = ~x90 & ~x538 ;
  assign n4554 = x90 & x538 ;
  assign n4555 = ~n4553 & ~n4554 ;
  assign n4556 = ~n4552 & ~n4555 ;
  assign n4557 = n4552 & n4555 ;
  assign n4558 = ~n4556 & ~n4557 ;
  assign n4559 = ~x92 & ~x540 ;
  assign n4560 = x92 & x540 ;
  assign n4561 = ~n4559 & ~n4560 ;
  assign n4562 = ~n4558 & ~n4561 ;
  assign n4563 = n4558 & n4561 ;
  assign n4564 = ~n4562 & ~n4563 ;
  assign n4565 = n4549 & ~n4564 ;
  assign n4566 = ~n4547 & ~n4565 ;
  assign n4567 = ~n4535 & ~n4542 ;
  assign n4568 = ~n4566 & n4567 ;
  assign n4569 = n4566 & ~n4567 ;
  assign n4570 = ~n4568 & ~n4569 ;
  assign n4571 = ~n4557 & ~n4563 ;
  assign n4572 = n4570 & n4571 ;
  assign n4573 = ~n4568 & ~n4572 ;
  assign n4574 = ~n4570 & ~n4571 ;
  assign n4575 = ~n4572 & ~n4574 ;
  assign n4576 = ~n4549 & n4564 ;
  assign n4577 = ~n4565 & ~n4576 ;
  assign n4578 = ~x81 & ~x529 ;
  assign n4579 = x81 & x529 ;
  assign n4580 = ~n4578 & ~n4579 ;
  assign n4581 = n4577 & ~n4580 ;
  assign n4582 = ~x87 & ~x535 ;
  assign n4583 = x87 & x535 ;
  assign n4584 = ~n4582 & ~n4583 ;
  assign n4585 = ~x86 & ~x534 ;
  assign n4586 = x86 & x534 ;
  assign n4587 = ~n4585 & ~n4586 ;
  assign n4588 = ~n4584 & ~n4587 ;
  assign n4589 = n4584 & n4587 ;
  assign n4590 = ~n4588 & ~n4589 ;
  assign n4591 = ~x88 & ~x536 ;
  assign n4592 = x88 & x536 ;
  assign n4593 = ~n4591 & ~n4592 ;
  assign n4594 = ~n4590 & ~n4593 ;
  assign n4595 = n4590 & n4593 ;
  assign n4596 = ~n4594 & ~n4595 ;
  assign n4597 = ~x82 & ~x530 ;
  assign n4598 = x82 & x530 ;
  assign n4599 = ~n4597 & ~n4598 ;
  assign n4600 = ~n4596 & ~n4599 ;
  assign n4601 = n4596 & n4599 ;
  assign n4602 = ~n4600 & ~n4601 ;
  assign n4603 = ~x84 & ~x532 ;
  assign n4604 = x84 & x532 ;
  assign n4605 = ~n4603 & ~n4604 ;
  assign n4606 = ~x83 & ~x531 ;
  assign n4607 = x83 & x531 ;
  assign n4608 = ~n4606 & ~n4607 ;
  assign n4609 = ~n4605 & ~n4608 ;
  assign n4610 = n4605 & n4608 ;
  assign n4611 = ~n4609 & ~n4610 ;
  assign n4612 = ~x85 & ~x533 ;
  assign n4613 = x85 & x533 ;
  assign n4614 = ~n4612 & ~n4613 ;
  assign n4615 = ~n4611 & ~n4614 ;
  assign n4616 = n4611 & n4614 ;
  assign n4617 = ~n4615 & ~n4616 ;
  assign n4618 = n4602 & ~n4617 ;
  assign n4619 = ~n4602 & n4617 ;
  assign n4620 = ~n4618 & ~n4619 ;
  assign n4621 = ~n4577 & n4580 ;
  assign n4622 = ~n4581 & ~n4621 ;
  assign n4623 = n4620 & n4622 ;
  assign n4624 = ~n4581 & ~n4623 ;
  assign n4625 = n4575 & ~n4624 ;
  assign n4626 = ~n4600 & ~n4618 ;
  assign n4627 = ~n4589 & ~n4595 ;
  assign n4628 = ~n4626 & n4627 ;
  assign n4629 = n4626 & ~n4627 ;
  assign n4630 = ~n4628 & ~n4629 ;
  assign n4631 = ~n4610 & ~n4616 ;
  assign n4632 = n4630 & n4631 ;
  assign n4633 = ~n4630 & ~n4631 ;
  assign n4634 = ~n4632 & ~n4633 ;
  assign n4635 = ~n4575 & n4624 ;
  assign n4636 = ~n4625 & ~n4635 ;
  assign n4637 = n4634 & n4636 ;
  assign n4638 = ~n4625 & ~n4637 ;
  assign n4639 = ~n4573 & ~n4638 ;
  assign n4640 = n4573 & n4638 ;
  assign n4641 = ~n4639 & ~n4640 ;
  assign n4642 = ~n4628 & ~n4632 ;
  assign n4643 = n4641 & ~n4642 ;
  assign n4644 = ~n4639 & ~n4643 ;
  assign n4645 = ~n4641 & n4642 ;
  assign n4646 = ~n4643 & ~n4645 ;
  assign n4647 = ~n4634 & ~n4636 ;
  assign n4648 = ~n4637 & ~n4647 ;
  assign n4649 = ~n4620 & ~n4622 ;
  assign n4650 = ~n4623 & ~n4649 ;
  assign n4651 = ~x65 & ~x513 ;
  assign n4652 = x65 & x513 ;
  assign n4653 = ~n4651 & ~n4652 ;
  assign n4654 = n4650 & ~n4653 ;
  assign n4655 = ~x72 & ~x520 ;
  assign n4656 = x72 & x520 ;
  assign n4657 = ~n4655 & ~n4656 ;
  assign n4658 = ~x71 & ~x519 ;
  assign n4659 = x71 & x519 ;
  assign n4660 = ~n4658 & ~n4659 ;
  assign n4661 = ~n4657 & ~n4660 ;
  assign n4662 = n4657 & n4660 ;
  assign n4663 = ~n4661 & ~n4662 ;
  assign n4664 = ~x73 & ~x521 ;
  assign n4665 = x73 & x521 ;
  assign n4666 = ~n4664 & ~n4665 ;
  assign n4667 = ~n4663 & ~n4666 ;
  assign n4668 = n4663 & n4666 ;
  assign n4669 = ~n4667 & ~n4668 ;
  assign n4670 = ~x67 & ~x515 ;
  assign n4671 = x67 & x515 ;
  assign n4672 = ~n4670 & ~n4671 ;
  assign n4673 = ~n4669 & ~n4672 ;
  assign n4674 = n4669 & n4672 ;
  assign n4675 = ~n4673 & ~n4674 ;
  assign n4676 = ~x69 & ~x517 ;
  assign n4677 = x69 & x517 ;
  assign n4678 = ~n4676 & ~n4677 ;
  assign n4679 = ~x68 & ~x516 ;
  assign n4680 = x68 & x516 ;
  assign n4681 = ~n4679 & ~n4680 ;
  assign n4682 = ~n4678 & ~n4681 ;
  assign n4683 = n4678 & n4681 ;
  assign n4684 = ~n4682 & ~n4683 ;
  assign n4685 = ~x70 & ~x518 ;
  assign n4686 = x70 & x518 ;
  assign n4687 = ~n4685 & ~n4686 ;
  assign n4688 = ~n4684 & ~n4687 ;
  assign n4689 = n4684 & n4687 ;
  assign n4690 = ~n4688 & ~n4689 ;
  assign n4691 = n4675 & ~n4690 ;
  assign n4692 = ~n4675 & n4690 ;
  assign n4693 = ~n4691 & ~n4692 ;
  assign n4694 = ~x79 & ~x527 ;
  assign n4695 = x79 & x527 ;
  assign n4696 = ~n4694 & ~n4695 ;
  assign n4697 = ~x78 & ~x526 ;
  assign n4698 = x78 & x526 ;
  assign n4699 = ~n4697 & ~n4698 ;
  assign n4700 = ~n4696 & ~n4699 ;
  assign n4701 = n4696 & n4699 ;
  assign n4702 = ~n4700 & ~n4701 ;
  assign n4703 = ~x80 & ~x528 ;
  assign n4704 = x80 & x528 ;
  assign n4705 = ~n4703 & ~n4704 ;
  assign n4706 = ~n4702 & ~n4705 ;
  assign n4707 = n4702 & n4705 ;
  assign n4708 = ~n4706 & ~n4707 ;
  assign n4709 = ~x74 & ~x522 ;
  assign n4710 = x74 & x522 ;
  assign n4711 = ~n4709 & ~n4710 ;
  assign n4712 = ~n4708 & ~n4711 ;
  assign n4713 = n4708 & n4711 ;
  assign n4714 = ~n4712 & ~n4713 ;
  assign n4715 = ~x76 & ~x524 ;
  assign n4716 = x76 & x524 ;
  assign n4717 = ~n4715 & ~n4716 ;
  assign n4718 = ~x75 & ~x523 ;
  assign n4719 = x75 & x523 ;
  assign n4720 = ~n4718 & ~n4719 ;
  assign n4721 = ~n4717 & ~n4720 ;
  assign n4722 = n4717 & n4720 ;
  assign n4723 = ~n4721 & ~n4722 ;
  assign n4724 = ~x77 & ~x525 ;
  assign n4725 = x77 & x525 ;
  assign n4726 = ~n4724 & ~n4725 ;
  assign n4727 = ~n4723 & ~n4726 ;
  assign n4728 = n4723 & n4726 ;
  assign n4729 = ~n4727 & ~n4728 ;
  assign n4730 = n4714 & ~n4729 ;
  assign n4731 = ~n4714 & n4729 ;
  assign n4732 = ~n4730 & ~n4731 ;
  assign n4733 = ~x66 & ~x514 ;
  assign n4734 = x66 & x514 ;
  assign n4735 = ~n4733 & ~n4734 ;
  assign n4736 = n4732 & ~n4735 ;
  assign n4737 = ~n4732 & n4735 ;
  assign n4738 = ~n4736 & ~n4737 ;
  assign n4739 = n4693 & n4738 ;
  assign n4740 = ~n4693 & ~n4738 ;
  assign n4741 = ~n4739 & ~n4740 ;
  assign n4742 = ~n4650 & n4653 ;
  assign n4743 = ~n4654 & ~n4742 ;
  assign n4744 = n4741 & n4743 ;
  assign n4745 = ~n4654 & ~n4744 ;
  assign n4746 = n4648 & ~n4745 ;
  assign n4747 = ~n4673 & ~n4691 ;
  assign n4748 = ~n4662 & ~n4668 ;
  assign n4749 = ~n4747 & n4748 ;
  assign n4750 = n4747 & ~n4748 ;
  assign n4751 = ~n4749 & ~n4750 ;
  assign n4752 = ~n4683 & ~n4689 ;
  assign n4753 = n4751 & n4752 ;
  assign n4754 = ~n4751 & ~n4752 ;
  assign n4755 = ~n4753 & ~n4754 ;
  assign n4756 = ~n4712 & ~n4730 ;
  assign n4757 = ~n4701 & ~n4707 ;
  assign n4758 = ~n4756 & n4757 ;
  assign n4759 = n4756 & ~n4757 ;
  assign n4760 = ~n4758 & ~n4759 ;
  assign n4761 = ~n4722 & ~n4728 ;
  assign n4762 = n4760 & n4761 ;
  assign n4763 = ~n4760 & ~n4761 ;
  assign n4764 = ~n4762 & ~n4763 ;
  assign n4765 = ~n4736 & ~n4739 ;
  assign n4766 = n4764 & ~n4765 ;
  assign n4767 = ~n4764 & n4765 ;
  assign n4768 = ~n4766 & ~n4767 ;
  assign n4769 = n4755 & n4768 ;
  assign n4770 = ~n4755 & ~n4768 ;
  assign n4771 = ~n4769 & ~n4770 ;
  assign n4772 = ~n4648 & n4745 ;
  assign n4773 = ~n4746 & ~n4772 ;
  assign n4774 = n4771 & n4773 ;
  assign n4775 = ~n4746 & ~n4774 ;
  assign n4776 = n4646 & ~n4775 ;
  assign n4777 = ~n4758 & ~n4762 ;
  assign n4778 = ~n4766 & ~n4769 ;
  assign n4779 = ~n4777 & ~n4778 ;
  assign n4780 = n4777 & n4778 ;
  assign n4781 = ~n4779 & ~n4780 ;
  assign n4782 = ~n4749 & ~n4753 ;
  assign n4783 = n4781 & ~n4782 ;
  assign n4784 = ~n4781 & n4782 ;
  assign n4785 = ~n4783 & ~n4784 ;
  assign n4786 = ~n4646 & n4775 ;
  assign n4787 = ~n4776 & ~n4786 ;
  assign n4788 = n4785 & n4787 ;
  assign n4789 = ~n4776 & ~n4788 ;
  assign n4790 = ~n4644 & ~n4789 ;
  assign n4791 = n4644 & n4789 ;
  assign n4792 = ~n4790 & ~n4791 ;
  assign n4793 = ~n4779 & ~n4783 ;
  assign n4794 = n4792 & ~n4793 ;
  assign n4795 = ~n4790 & ~n4794 ;
  assign n4796 = ~n4792 & n4793 ;
  assign n4797 = ~n4794 & ~n4796 ;
  assign n4798 = ~n4785 & ~n4787 ;
  assign n4799 = ~n4788 & ~n4798 ;
  assign n4800 = ~n4741 & ~n4743 ;
  assign n4801 = ~n4744 & ~n4800 ;
  assign n4802 = ~x64 & ~x512 ;
  assign n4803 = x64 & x512 ;
  assign n4804 = ~n4802 & ~n4803 ;
  assign n4805 = ~n4801 & n4804 ;
  assign n4806 = ~n4771 & ~n4773 ;
  assign n4807 = ~n4774 & ~n4806 ;
  assign n4808 = n4805 & ~n4807 ;
  assign n4809 = ~n4799 & n4808 ;
  assign n4810 = ~n4797 & n4809 ;
  assign n4811 = n4795 & n4810 ;
  assign n4812 = n4528 & n4811 ;
  assign n4813 = ~x62 & ~x542 ;
  assign n4814 = x62 & x542 ;
  assign n4815 = ~n4813 & ~n4814 ;
  assign n4816 = ~x61 & ~x541 ;
  assign n4817 = x61 & x541 ;
  assign n4818 = ~n4816 & ~n4817 ;
  assign n4819 = ~n4815 & ~n4818 ;
  assign n4820 = n4815 & n4818 ;
  assign n4821 = ~n4819 & ~n4820 ;
  assign n4822 = ~x63 & ~x543 ;
  assign n4823 = x63 & x543 ;
  assign n4824 = ~n4822 & ~n4823 ;
  assign n4825 = ~n4821 & ~n4824 ;
  assign n4826 = n4821 & n4824 ;
  assign n4827 = ~n4825 & ~n4826 ;
  assign n4828 = ~x57 & ~x537 ;
  assign n4829 = x57 & x537 ;
  assign n4830 = ~n4828 & ~n4829 ;
  assign n4831 = ~n4827 & ~n4830 ;
  assign n4832 = n4827 & n4830 ;
  assign n4833 = ~n4831 & ~n4832 ;
  assign n4834 = ~x59 & ~x539 ;
  assign n4835 = x59 & x539 ;
  assign n4836 = ~n4834 & ~n4835 ;
  assign n4837 = ~x58 & ~x538 ;
  assign n4838 = x58 & x538 ;
  assign n4839 = ~n4837 & ~n4838 ;
  assign n4840 = ~n4836 & ~n4839 ;
  assign n4841 = n4836 & n4839 ;
  assign n4842 = ~n4840 & ~n4841 ;
  assign n4843 = ~x60 & ~x540 ;
  assign n4844 = x60 & x540 ;
  assign n4845 = ~n4843 & ~n4844 ;
  assign n4846 = ~n4842 & ~n4845 ;
  assign n4847 = n4842 & n4845 ;
  assign n4848 = ~n4846 & ~n4847 ;
  assign n4849 = n4833 & ~n4848 ;
  assign n4850 = ~n4831 & ~n4849 ;
  assign n4851 = ~n4820 & ~n4826 ;
  assign n4852 = ~n4850 & n4851 ;
  assign n4853 = n4850 & ~n4851 ;
  assign n4854 = ~n4852 & ~n4853 ;
  assign n4855 = ~n4841 & ~n4847 ;
  assign n4856 = n4854 & n4855 ;
  assign n4857 = ~n4852 & ~n4856 ;
  assign n4858 = ~n4854 & ~n4855 ;
  assign n4859 = ~n4856 & ~n4858 ;
  assign n4860 = ~n4833 & n4848 ;
  assign n4861 = ~n4849 & ~n4860 ;
  assign n4862 = ~x49 & ~x529 ;
  assign n4863 = x49 & x529 ;
  assign n4864 = ~n4862 & ~n4863 ;
  assign n4865 = n4861 & ~n4864 ;
  assign n4866 = ~x55 & ~x535 ;
  assign n4867 = x55 & x535 ;
  assign n4868 = ~n4866 & ~n4867 ;
  assign n4869 = ~x54 & ~x534 ;
  assign n4870 = x54 & x534 ;
  assign n4871 = ~n4869 & ~n4870 ;
  assign n4872 = ~n4868 & ~n4871 ;
  assign n4873 = n4868 & n4871 ;
  assign n4874 = ~n4872 & ~n4873 ;
  assign n4875 = ~x56 & ~x536 ;
  assign n4876 = x56 & x536 ;
  assign n4877 = ~n4875 & ~n4876 ;
  assign n4878 = ~n4874 & ~n4877 ;
  assign n4879 = n4874 & n4877 ;
  assign n4880 = ~n4878 & ~n4879 ;
  assign n4881 = ~x50 & ~x530 ;
  assign n4882 = x50 & x530 ;
  assign n4883 = ~n4881 & ~n4882 ;
  assign n4884 = ~n4880 & ~n4883 ;
  assign n4885 = n4880 & n4883 ;
  assign n4886 = ~n4884 & ~n4885 ;
  assign n4887 = ~x52 & ~x532 ;
  assign n4888 = x52 & x532 ;
  assign n4889 = ~n4887 & ~n4888 ;
  assign n4890 = ~x51 & ~x531 ;
  assign n4891 = x51 & x531 ;
  assign n4892 = ~n4890 & ~n4891 ;
  assign n4893 = ~n4889 & ~n4892 ;
  assign n4894 = n4889 & n4892 ;
  assign n4895 = ~n4893 & ~n4894 ;
  assign n4896 = ~x53 & ~x533 ;
  assign n4897 = x53 & x533 ;
  assign n4898 = ~n4896 & ~n4897 ;
  assign n4899 = ~n4895 & ~n4898 ;
  assign n4900 = n4895 & n4898 ;
  assign n4901 = ~n4899 & ~n4900 ;
  assign n4902 = n4886 & ~n4901 ;
  assign n4903 = ~n4886 & n4901 ;
  assign n4904 = ~n4902 & ~n4903 ;
  assign n4905 = ~n4861 & n4864 ;
  assign n4906 = ~n4865 & ~n4905 ;
  assign n4907 = n4904 & n4906 ;
  assign n4908 = ~n4865 & ~n4907 ;
  assign n4909 = n4859 & ~n4908 ;
  assign n4910 = ~n4884 & ~n4902 ;
  assign n4911 = ~n4873 & ~n4879 ;
  assign n4912 = ~n4910 & n4911 ;
  assign n4913 = n4910 & ~n4911 ;
  assign n4914 = ~n4912 & ~n4913 ;
  assign n4915 = ~n4894 & ~n4900 ;
  assign n4916 = n4914 & n4915 ;
  assign n4917 = ~n4914 & ~n4915 ;
  assign n4918 = ~n4916 & ~n4917 ;
  assign n4919 = ~n4859 & n4908 ;
  assign n4920 = ~n4909 & ~n4919 ;
  assign n4921 = n4918 & n4920 ;
  assign n4922 = ~n4909 & ~n4921 ;
  assign n4923 = ~n4857 & ~n4922 ;
  assign n4924 = n4857 & n4922 ;
  assign n4925 = ~n4923 & ~n4924 ;
  assign n4926 = ~n4912 & ~n4916 ;
  assign n4927 = n4925 & ~n4926 ;
  assign n4928 = ~n4923 & ~n4927 ;
  assign n4929 = ~n4925 & n4926 ;
  assign n4930 = ~n4927 & ~n4929 ;
  assign n4931 = ~n4918 & ~n4920 ;
  assign n4932 = ~n4921 & ~n4931 ;
  assign n4933 = ~n4904 & ~n4906 ;
  assign n4934 = ~n4907 & ~n4933 ;
  assign n4935 = ~x33 & ~x513 ;
  assign n4936 = x33 & x513 ;
  assign n4937 = ~n4935 & ~n4936 ;
  assign n4938 = n4934 & ~n4937 ;
  assign n4939 = ~x40 & ~x520 ;
  assign n4940 = x40 & x520 ;
  assign n4941 = ~n4939 & ~n4940 ;
  assign n4942 = ~x39 & ~x519 ;
  assign n4943 = x39 & x519 ;
  assign n4944 = ~n4942 & ~n4943 ;
  assign n4945 = ~n4941 & ~n4944 ;
  assign n4946 = n4941 & n4944 ;
  assign n4947 = ~n4945 & ~n4946 ;
  assign n4948 = ~x41 & ~x521 ;
  assign n4949 = x41 & x521 ;
  assign n4950 = ~n4948 & ~n4949 ;
  assign n4951 = ~n4947 & ~n4950 ;
  assign n4952 = n4947 & n4950 ;
  assign n4953 = ~n4951 & ~n4952 ;
  assign n4954 = ~x35 & ~x515 ;
  assign n4955 = x35 & x515 ;
  assign n4956 = ~n4954 & ~n4955 ;
  assign n4957 = ~n4953 & ~n4956 ;
  assign n4958 = n4953 & n4956 ;
  assign n4959 = ~n4957 & ~n4958 ;
  assign n4960 = ~x37 & ~x517 ;
  assign n4961 = x37 & x517 ;
  assign n4962 = ~n4960 & ~n4961 ;
  assign n4963 = ~x36 & ~x516 ;
  assign n4964 = x36 & x516 ;
  assign n4965 = ~n4963 & ~n4964 ;
  assign n4966 = ~n4962 & ~n4965 ;
  assign n4967 = n4962 & n4965 ;
  assign n4968 = ~n4966 & ~n4967 ;
  assign n4969 = ~x38 & ~x518 ;
  assign n4970 = x38 & x518 ;
  assign n4971 = ~n4969 & ~n4970 ;
  assign n4972 = ~n4968 & ~n4971 ;
  assign n4973 = n4968 & n4971 ;
  assign n4974 = ~n4972 & ~n4973 ;
  assign n4975 = n4959 & ~n4974 ;
  assign n4976 = ~n4959 & n4974 ;
  assign n4977 = ~n4975 & ~n4976 ;
  assign n4978 = ~x47 & ~x527 ;
  assign n4979 = x47 & x527 ;
  assign n4980 = ~n4978 & ~n4979 ;
  assign n4981 = ~x46 & ~x526 ;
  assign n4982 = x46 & x526 ;
  assign n4983 = ~n4981 & ~n4982 ;
  assign n4984 = ~n4980 & ~n4983 ;
  assign n4985 = n4980 & n4983 ;
  assign n4986 = ~n4984 & ~n4985 ;
  assign n4987 = ~x48 & ~x528 ;
  assign n4988 = x48 & x528 ;
  assign n4989 = ~n4987 & ~n4988 ;
  assign n4990 = ~n4986 & ~n4989 ;
  assign n4991 = n4986 & n4989 ;
  assign n4992 = ~n4990 & ~n4991 ;
  assign n4993 = ~x42 & ~x522 ;
  assign n4994 = x42 & x522 ;
  assign n4995 = ~n4993 & ~n4994 ;
  assign n4996 = ~n4992 & ~n4995 ;
  assign n4997 = n4992 & n4995 ;
  assign n4998 = ~n4996 & ~n4997 ;
  assign n4999 = ~x44 & ~x524 ;
  assign n5000 = x44 & x524 ;
  assign n5001 = ~n4999 & ~n5000 ;
  assign n5002 = ~x43 & ~x523 ;
  assign n5003 = x43 & x523 ;
  assign n5004 = ~n5002 & ~n5003 ;
  assign n5005 = ~n5001 & ~n5004 ;
  assign n5006 = n5001 & n5004 ;
  assign n5007 = ~n5005 & ~n5006 ;
  assign n5008 = ~x45 & ~x525 ;
  assign n5009 = x45 & x525 ;
  assign n5010 = ~n5008 & ~n5009 ;
  assign n5011 = ~n5007 & ~n5010 ;
  assign n5012 = n5007 & n5010 ;
  assign n5013 = ~n5011 & ~n5012 ;
  assign n5014 = n4998 & ~n5013 ;
  assign n5015 = ~n4998 & n5013 ;
  assign n5016 = ~n5014 & ~n5015 ;
  assign n5017 = ~x34 & ~x514 ;
  assign n5018 = x34 & x514 ;
  assign n5019 = ~n5017 & ~n5018 ;
  assign n5020 = n5016 & ~n5019 ;
  assign n5021 = ~n5016 & n5019 ;
  assign n5022 = ~n5020 & ~n5021 ;
  assign n5023 = n4977 & n5022 ;
  assign n5024 = ~n4977 & ~n5022 ;
  assign n5025 = ~n5023 & ~n5024 ;
  assign n5026 = ~n4934 & n4937 ;
  assign n5027 = ~n4938 & ~n5026 ;
  assign n5028 = n5025 & n5027 ;
  assign n5029 = ~n4938 & ~n5028 ;
  assign n5030 = n4932 & ~n5029 ;
  assign n5031 = ~n4957 & ~n4975 ;
  assign n5032 = ~n4946 & ~n4952 ;
  assign n5033 = ~n5031 & n5032 ;
  assign n5034 = n5031 & ~n5032 ;
  assign n5035 = ~n5033 & ~n5034 ;
  assign n5036 = ~n4967 & ~n4973 ;
  assign n5037 = n5035 & n5036 ;
  assign n5038 = ~n5035 & ~n5036 ;
  assign n5039 = ~n5037 & ~n5038 ;
  assign n5040 = ~n4996 & ~n5014 ;
  assign n5041 = ~n4985 & ~n4991 ;
  assign n5042 = ~n5040 & n5041 ;
  assign n5043 = n5040 & ~n5041 ;
  assign n5044 = ~n5042 & ~n5043 ;
  assign n5045 = ~n5006 & ~n5012 ;
  assign n5046 = n5044 & n5045 ;
  assign n5047 = ~n5044 & ~n5045 ;
  assign n5048 = ~n5046 & ~n5047 ;
  assign n5049 = ~n5020 & ~n5023 ;
  assign n5050 = n5048 & ~n5049 ;
  assign n5051 = ~n5048 & n5049 ;
  assign n5052 = ~n5050 & ~n5051 ;
  assign n5053 = n5039 & n5052 ;
  assign n5054 = ~n5039 & ~n5052 ;
  assign n5055 = ~n5053 & ~n5054 ;
  assign n5056 = ~n4932 & n5029 ;
  assign n5057 = ~n5030 & ~n5056 ;
  assign n5058 = n5055 & n5057 ;
  assign n5059 = ~n5030 & ~n5058 ;
  assign n5060 = n4930 & ~n5059 ;
  assign n5061 = ~n5042 & ~n5046 ;
  assign n5062 = ~n5050 & ~n5053 ;
  assign n5063 = ~n5061 & ~n5062 ;
  assign n5064 = n5061 & n5062 ;
  assign n5065 = ~n5063 & ~n5064 ;
  assign n5066 = ~n5033 & ~n5037 ;
  assign n5067 = n5065 & ~n5066 ;
  assign n5068 = ~n5065 & n5066 ;
  assign n5069 = ~n5067 & ~n5068 ;
  assign n5070 = ~n4930 & n5059 ;
  assign n5071 = ~n5060 & ~n5070 ;
  assign n5072 = n5069 & n5071 ;
  assign n5073 = ~n5060 & ~n5072 ;
  assign n5074 = ~n4928 & ~n5073 ;
  assign n5075 = n4928 & n5073 ;
  assign n5076 = ~n5074 & ~n5075 ;
  assign n5077 = ~n5063 & ~n5067 ;
  assign n5078 = n5076 & ~n5077 ;
  assign n5079 = ~n5074 & ~n5078 ;
  assign n5080 = ~n5076 & n5077 ;
  assign n5081 = ~n5078 & ~n5080 ;
  assign n5082 = ~n5069 & ~n5071 ;
  assign n5083 = ~n5072 & ~n5082 ;
  assign n5084 = ~n5025 & ~n5027 ;
  assign n5085 = ~n5028 & ~n5084 ;
  assign n5086 = ~x32 & ~x512 ;
  assign n5087 = x32 & x512 ;
  assign n5088 = ~n5086 & ~n5087 ;
  assign n5089 = ~n5085 & n5088 ;
  assign n5090 = ~n5055 & ~n5057 ;
  assign n5091 = ~n5058 & ~n5090 ;
  assign n5092 = n5089 & ~n5091 ;
  assign n5093 = ~n5083 & n5092 ;
  assign n5094 = ~n5081 & n5093 ;
  assign n5095 = n5079 & n5094 ;
  assign n5096 = n4812 & n5095 ;
  assign n5097 = ~n827 & n5096 ;
  assign n5098 = n816 & ~n822 ;
  assign n5099 = ~n823 & ~n5098 ;
  assign n5100 = ~n4805 & n4807 ;
  assign n5101 = ~n4808 & ~n5100 ;
  assign n5102 = ~n4528 & n4811 ;
  assign n5103 = n4517 & ~n4523 ;
  assign n5104 = ~n4524 & ~n5103 ;
  assign n5105 = ~n4244 & n4527 ;
  assign n5106 = ~n1381 & ~n1402 ;
  assign n5107 = ~n1093 & ~n1112 ;
  assign n5108 = ~n5106 & ~n5107 ;
  assign n5109 = ~n1404 & n5108 ;
  assign n5110 = ~n1404 & n1687 ;
  assign n5111 = ~n1671 & ~n1686 ;
  assign n5112 = ~n1687 & ~n5111 ;
  assign n5113 = n5109 & ~n5112 ;
  assign n5114 = n1404 & ~n1687 ;
  assign n5115 = n1677 & ~n1683 ;
  assign n5116 = ~n1684 & ~n5115 ;
  assign n5117 = ~n1391 & ~n1395 ;
  assign n5118 = ~n1396 & ~n5117 ;
  assign n5119 = n1113 & ~n1403 ;
  assign n5120 = ~n1113 & ~n5107 ;
  assign n5121 = ~n1403 & ~n5106 ;
  assign n5122 = n5120 & ~n5121 ;
  assign n5123 = n1383 & ~n1401 ;
  assign n5124 = ~n1402 & ~n5123 ;
  assign n5125 = ~n1396 & ~n1400 ;
  assign n5126 = ~n1401 & ~n5125 ;
  assign n5127 = ~n1097 & ~n1100 ;
  assign n5128 = ~n1101 & ~n5127 ;
  assign n5129 = ~n1386 & n1390 ;
  assign n5130 = ~n1391 & ~n5129 ;
  assign n5131 = ~n5128 & n5130 ;
  assign n5132 = n1395 & n5131 ;
  assign n5133 = ~n1101 & ~n1105 ;
  assign n5134 = ~n1106 & ~n5133 ;
  assign n5135 = ~n5118 & ~n5131 ;
  assign n5136 = ~n5134 & ~n5135 ;
  assign n5137 = ~n5132 & ~n5136 ;
  assign n5138 = n5126 & ~n5137 ;
  assign n5139 = ~n5126 & n5137 ;
  assign n5140 = ~n1106 & ~n1110 ;
  assign n5141 = ~n1111 & ~n5140 ;
  assign n5142 = ~n5139 & ~n5141 ;
  assign n5143 = ~n5138 & ~n5142 ;
  assign n5144 = ~n5124 & n5143 ;
  assign n5145 = n1095 & ~n1111 ;
  assign n5146 = ~n1112 & ~n5145 ;
  assign n5147 = n5124 & ~n5143 ;
  assign n5148 = n5146 & ~n5147 ;
  assign n5149 = ~n5144 & ~n5148 ;
  assign n5150 = ~n5122 & n5149 ;
  assign n5151 = ~n1113 & n1403 ;
  assign n5152 = ~n5120 & n5121 ;
  assign n5153 = ~n5151 & ~n5152 ;
  assign n5154 = ~n5150 & n5153 ;
  assign n5155 = ~n5119 & ~n5154 ;
  assign n5156 = ~n5118 & ~n5155 ;
  assign n5157 = ~n5134 & n5155 ;
  assign n5158 = ~n5156 & ~n5157 ;
  assign n5159 = ~n5116 & n5158 ;
  assign n5160 = n1679 & ~n1682 ;
  assign n5161 = ~n1683 & ~n5160 ;
  assign n5162 = ~n5130 & ~n5155 ;
  assign n5163 = ~n5128 & n5155 ;
  assign n5164 = ~n5162 & ~n5163 ;
  assign n5165 = n5161 & ~n5164 ;
  assign n5166 = ~n5159 & n5165 ;
  assign n5167 = n1675 & ~n1684 ;
  assign n5168 = ~n1685 & ~n5167 ;
  assign n5169 = ~n5126 & ~n5155 ;
  assign n5170 = ~n5141 & n5155 ;
  assign n5171 = ~n5169 & ~n5170 ;
  assign n5172 = n5168 & ~n5171 ;
  assign n5173 = n5116 & ~n5158 ;
  assign n5174 = ~n5172 & ~n5173 ;
  assign n5175 = ~n5166 & n5174 ;
  assign n5176 = n1673 & ~n1685 ;
  assign n5177 = ~n1686 & ~n5176 ;
  assign n5178 = ~n5124 & ~n5155 ;
  assign n5179 = ~n5146 & n5155 ;
  assign n5180 = ~n5178 & ~n5179 ;
  assign n5181 = ~n5177 & n5180 ;
  assign n5182 = ~n5168 & n5171 ;
  assign n5183 = ~n5181 & ~n5182 ;
  assign n5184 = ~n5175 & n5183 ;
  assign n5185 = n5177 & ~n5180 ;
  assign n5186 = ~n5109 & n5112 ;
  assign n5187 = ~n5185 & ~n5186 ;
  assign n5188 = ~n5184 & n5187 ;
  assign n5189 = ~n5114 & ~n5188 ;
  assign n5190 = ~n5113 & n5189 ;
  assign n5191 = ~n5110 & ~n5190 ;
  assign n5192 = n5109 & ~n5191 ;
  assign n5193 = n5112 & ~n5189 ;
  assign n5194 = ~n5192 & ~n5193 ;
  assign n5195 = ~n1688 & n1971 ;
  assign n5196 = n1961 & ~n1967 ;
  assign n5197 = ~n1968 & ~n5196 ;
  assign n5198 = ~n5116 & n5191 ;
  assign n5199 = ~n5158 & ~n5191 ;
  assign n5200 = ~n5198 & ~n5199 ;
  assign n5201 = ~n5197 & n5200 ;
  assign n5202 = n1963 & ~n1966 ;
  assign n5203 = ~n1967 & ~n5202 ;
  assign n5204 = n5164 & ~n5191 ;
  assign n5205 = n5161 & n5191 ;
  assign n5206 = ~n5204 & ~n5205 ;
  assign n5207 = n5203 & n5206 ;
  assign n5208 = ~n5201 & n5207 ;
  assign n5209 = n1959 & ~n1968 ;
  assign n5210 = ~n1969 & ~n5209 ;
  assign n5211 = ~n5168 & n5191 ;
  assign n5212 = ~n5171 & ~n5191 ;
  assign n5213 = ~n5211 & ~n5212 ;
  assign n5214 = n5210 & ~n5213 ;
  assign n5215 = n5197 & ~n5200 ;
  assign n5216 = ~n5214 & ~n5215 ;
  assign n5217 = ~n5208 & n5216 ;
  assign n5218 = n1957 & ~n1969 ;
  assign n5219 = ~n1970 & ~n5218 ;
  assign n5220 = ~n5177 & n5191 ;
  assign n5221 = ~n5180 & ~n5191 ;
  assign n5222 = ~n5220 & ~n5221 ;
  assign n5223 = ~n5219 & n5222 ;
  assign n5224 = ~n5210 & n5213 ;
  assign n5225 = ~n5223 & ~n5224 ;
  assign n5226 = ~n5217 & n5225 ;
  assign n5227 = ~n1955 & ~n1970 ;
  assign n5228 = ~n1971 & ~n5227 ;
  assign n5229 = n5194 & n5228 ;
  assign n5230 = n5219 & ~n5222 ;
  assign n5231 = ~n5229 & ~n5230 ;
  assign n5232 = ~n5226 & n5231 ;
  assign n5233 = n1688 & ~n1971 ;
  assign n5234 = ~n5194 & ~n5228 ;
  assign n5235 = ~n5233 & ~n5234 ;
  assign n5236 = ~n5232 & n5235 ;
  assign n5237 = ~n5195 & ~n5236 ;
  assign n5238 = ~n5194 & ~n5237 ;
  assign n5239 = n5228 & ~n5236 ;
  assign n5240 = ~n5238 & ~n5239 ;
  assign n5241 = ~n1972 & n2255 ;
  assign n5242 = ~n2239 & ~n2254 ;
  assign n5243 = ~n2255 & ~n5242 ;
  assign n5244 = ~n5240 & ~n5243 ;
  assign n5245 = n1972 & ~n2255 ;
  assign n5246 = n2245 & ~n2251 ;
  assign n5247 = ~n2252 & ~n5246 ;
  assign n5248 = ~n5197 & n5237 ;
  assign n5249 = ~n5200 & ~n5237 ;
  assign n5250 = ~n5248 & ~n5249 ;
  assign n5251 = ~n5247 & n5250 ;
  assign n5252 = n2247 & ~n2250 ;
  assign n5253 = ~n2251 & ~n5252 ;
  assign n5254 = n5206 & ~n5237 ;
  assign n5255 = ~n5203 & n5237 ;
  assign n5256 = ~n5254 & ~n5255 ;
  assign n5257 = n5253 & ~n5256 ;
  assign n5258 = ~n5251 & n5257 ;
  assign n5259 = n2243 & ~n2252 ;
  assign n5260 = ~n2253 & ~n5259 ;
  assign n5261 = n5213 & ~n5237 ;
  assign n5262 = n5210 & n5237 ;
  assign n5263 = ~n5261 & ~n5262 ;
  assign n5264 = n5260 & n5263 ;
  assign n5265 = n5247 & ~n5250 ;
  assign n5266 = ~n5264 & ~n5265 ;
  assign n5267 = ~n5258 & n5266 ;
  assign n5268 = n2241 & ~n2253 ;
  assign n5269 = ~n2254 & ~n5268 ;
  assign n5270 = ~n5219 & n5237 ;
  assign n5271 = ~n5222 & ~n5237 ;
  assign n5272 = ~n5270 & ~n5271 ;
  assign n5273 = ~n5269 & n5272 ;
  assign n5274 = ~n5260 & ~n5263 ;
  assign n5275 = ~n5273 & ~n5274 ;
  assign n5276 = ~n5267 & n5275 ;
  assign n5277 = n5269 & ~n5272 ;
  assign n5278 = n5240 & n5243 ;
  assign n5279 = ~n5277 & ~n5278 ;
  assign n5280 = ~n5276 & n5279 ;
  assign n5281 = ~n5245 & ~n5280 ;
  assign n5282 = ~n5244 & n5281 ;
  assign n5283 = ~n5241 & ~n5282 ;
  assign n5284 = ~n5240 & ~n5283 ;
  assign n5285 = n5243 & ~n5281 ;
  assign n5286 = ~n5284 & ~n5285 ;
  assign n5287 = ~n2256 & n2539 ;
  assign n5288 = n2529 & ~n2535 ;
  assign n5289 = ~n2536 & ~n5288 ;
  assign n5290 = ~n5247 & n5283 ;
  assign n5291 = ~n5250 & ~n5283 ;
  assign n5292 = ~n5290 & ~n5291 ;
  assign n5293 = ~n5289 & n5292 ;
  assign n5294 = n2531 & ~n2534 ;
  assign n5295 = ~n2535 & ~n5294 ;
  assign n5296 = n5256 & ~n5283 ;
  assign n5297 = n5253 & n5283 ;
  assign n5298 = ~n5296 & ~n5297 ;
  assign n5299 = n5295 & n5298 ;
  assign n5300 = ~n5293 & n5299 ;
  assign n5301 = n2527 & ~n2536 ;
  assign n5302 = ~n2537 & ~n5301 ;
  assign n5303 = ~n5260 & n5283 ;
  assign n5304 = n5263 & ~n5283 ;
  assign n5305 = ~n5303 & ~n5304 ;
  assign n5306 = n5302 & ~n5305 ;
  assign n5307 = n5289 & ~n5292 ;
  assign n5308 = ~n5306 & ~n5307 ;
  assign n5309 = ~n5300 & n5308 ;
  assign n5310 = n2525 & ~n2537 ;
  assign n5311 = ~n2538 & ~n5310 ;
  assign n5312 = ~n5269 & n5283 ;
  assign n5313 = ~n5272 & ~n5283 ;
  assign n5314 = ~n5312 & ~n5313 ;
  assign n5315 = ~n5311 & n5314 ;
  assign n5316 = ~n5302 & n5305 ;
  assign n5317 = ~n5315 & ~n5316 ;
  assign n5318 = ~n5309 & n5317 ;
  assign n5319 = ~n2523 & ~n2538 ;
  assign n5320 = ~n2539 & ~n5319 ;
  assign n5321 = n5286 & n5320 ;
  assign n5322 = n5311 & ~n5314 ;
  assign n5323 = ~n5321 & ~n5322 ;
  assign n5324 = ~n5318 & n5323 ;
  assign n5325 = n2256 & ~n2539 ;
  assign n5326 = ~n5286 & ~n5320 ;
  assign n5327 = ~n5325 & ~n5326 ;
  assign n5328 = ~n5324 & n5327 ;
  assign n5329 = ~n5287 & ~n5328 ;
  assign n5330 = ~n5286 & ~n5329 ;
  assign n5331 = n5320 & ~n5328 ;
  assign n5332 = ~n5330 & ~n5331 ;
  assign n5333 = ~n2540 & n2823 ;
  assign n5334 = ~n2807 & ~n2822 ;
  assign n5335 = ~n2823 & ~n5334 ;
  assign n5336 = ~n5332 & ~n5335 ;
  assign n5337 = n2540 & ~n2823 ;
  assign n5338 = n2813 & ~n2819 ;
  assign n5339 = ~n2820 & ~n5338 ;
  assign n5340 = ~n5289 & n5329 ;
  assign n5341 = ~n5292 & ~n5329 ;
  assign n5342 = ~n5340 & ~n5341 ;
  assign n5343 = ~n5339 & n5342 ;
  assign n5344 = n2815 & ~n2818 ;
  assign n5345 = ~n2819 & ~n5344 ;
  assign n5346 = n5298 & ~n5329 ;
  assign n5347 = ~n5295 & n5329 ;
  assign n5348 = ~n5346 & ~n5347 ;
  assign n5349 = n5345 & ~n5348 ;
  assign n5350 = ~n5343 & n5349 ;
  assign n5351 = n2811 & ~n2820 ;
  assign n5352 = ~n2821 & ~n5351 ;
  assign n5353 = n5305 & ~n5329 ;
  assign n5354 = n5302 & n5329 ;
  assign n5355 = ~n5353 & ~n5354 ;
  assign n5356 = n5352 & n5355 ;
  assign n5357 = n5339 & ~n5342 ;
  assign n5358 = ~n5356 & ~n5357 ;
  assign n5359 = ~n5350 & n5358 ;
  assign n5360 = n2809 & ~n2821 ;
  assign n5361 = ~n2822 & ~n5360 ;
  assign n5362 = ~n5311 & n5329 ;
  assign n5363 = ~n5314 & ~n5329 ;
  assign n5364 = ~n5362 & ~n5363 ;
  assign n5365 = ~n5361 & n5364 ;
  assign n5366 = ~n5352 & ~n5355 ;
  assign n5367 = ~n5365 & ~n5366 ;
  assign n5368 = ~n5359 & n5367 ;
  assign n5369 = n5361 & ~n5364 ;
  assign n5370 = n5332 & n5335 ;
  assign n5371 = ~n5369 & ~n5370 ;
  assign n5372 = ~n5368 & n5371 ;
  assign n5373 = ~n5337 & ~n5372 ;
  assign n5374 = ~n5336 & n5373 ;
  assign n5375 = ~n5333 & ~n5374 ;
  assign n5376 = ~n5332 & ~n5375 ;
  assign n5377 = n5335 & ~n5373 ;
  assign n5378 = ~n5376 & ~n5377 ;
  assign n5379 = ~n2824 & n3107 ;
  assign n5380 = n3097 & ~n3103 ;
  assign n5381 = ~n3104 & ~n5380 ;
  assign n5382 = ~n5339 & n5375 ;
  assign n5383 = ~n5342 & ~n5375 ;
  assign n5384 = ~n5382 & ~n5383 ;
  assign n5385 = ~n5381 & n5384 ;
  assign n5386 = n3099 & ~n3102 ;
  assign n5387 = ~n3103 & ~n5386 ;
  assign n5388 = n5348 & ~n5375 ;
  assign n5389 = n5345 & n5375 ;
  assign n5390 = ~n5388 & ~n5389 ;
  assign n5391 = n5387 & n5390 ;
  assign n5392 = ~n5385 & n5391 ;
  assign n5393 = n3095 & ~n3104 ;
  assign n5394 = ~n3105 & ~n5393 ;
  assign n5395 = ~n5352 & n5375 ;
  assign n5396 = n5355 & ~n5375 ;
  assign n5397 = ~n5395 & ~n5396 ;
  assign n5398 = n5394 & ~n5397 ;
  assign n5399 = n5381 & ~n5384 ;
  assign n5400 = ~n5398 & ~n5399 ;
  assign n5401 = ~n5392 & n5400 ;
  assign n5402 = n3093 & ~n3105 ;
  assign n5403 = ~n3106 & ~n5402 ;
  assign n5404 = ~n5361 & n5375 ;
  assign n5405 = ~n5364 & ~n5375 ;
  assign n5406 = ~n5404 & ~n5405 ;
  assign n5407 = ~n5403 & n5406 ;
  assign n5408 = ~n5394 & n5397 ;
  assign n5409 = ~n5407 & ~n5408 ;
  assign n5410 = ~n5401 & n5409 ;
  assign n5411 = ~n3091 & ~n3106 ;
  assign n5412 = ~n3107 & ~n5411 ;
  assign n5413 = n5378 & n5412 ;
  assign n5414 = n5403 & ~n5406 ;
  assign n5415 = ~n5413 & ~n5414 ;
  assign n5416 = ~n5410 & n5415 ;
  assign n5417 = n2824 & ~n3107 ;
  assign n5418 = ~n5378 & ~n5412 ;
  assign n5419 = ~n5417 & ~n5418 ;
  assign n5420 = ~n5416 & n5419 ;
  assign n5421 = ~n5379 & ~n5420 ;
  assign n5422 = ~n5378 & ~n5421 ;
  assign n5423 = n5412 & ~n5420 ;
  assign n5424 = ~n5422 & ~n5423 ;
  assign n5425 = ~n3108 & n3391 ;
  assign n5426 = ~n3375 & ~n3390 ;
  assign n5427 = ~n3391 & ~n5426 ;
  assign n5428 = ~n5424 & ~n5427 ;
  assign n5429 = n3108 & ~n3391 ;
  assign n5430 = n3381 & ~n3387 ;
  assign n5431 = ~n3388 & ~n5430 ;
  assign n5432 = ~n5381 & n5421 ;
  assign n5433 = ~n5384 & ~n5421 ;
  assign n5434 = ~n5432 & ~n5433 ;
  assign n5435 = ~n5431 & n5434 ;
  assign n5436 = n3383 & ~n3386 ;
  assign n5437 = ~n3387 & ~n5436 ;
  assign n5438 = n5390 & ~n5421 ;
  assign n5439 = ~n5387 & n5421 ;
  assign n5440 = ~n5438 & ~n5439 ;
  assign n5441 = n5437 & ~n5440 ;
  assign n5442 = ~n5435 & n5441 ;
  assign n5443 = n3379 & ~n3388 ;
  assign n5444 = ~n3389 & ~n5443 ;
  assign n5445 = n5397 & ~n5421 ;
  assign n5446 = n5394 & n5421 ;
  assign n5447 = ~n5445 & ~n5446 ;
  assign n5448 = n5444 & n5447 ;
  assign n5449 = n5431 & ~n5434 ;
  assign n5450 = ~n5448 & ~n5449 ;
  assign n5451 = ~n5442 & n5450 ;
  assign n5452 = n3377 & ~n3389 ;
  assign n5453 = ~n3390 & ~n5452 ;
  assign n5454 = ~n5403 & n5421 ;
  assign n5455 = ~n5406 & ~n5421 ;
  assign n5456 = ~n5454 & ~n5455 ;
  assign n5457 = ~n5453 & n5456 ;
  assign n5458 = ~n5444 & ~n5447 ;
  assign n5459 = ~n5457 & ~n5458 ;
  assign n5460 = ~n5451 & n5459 ;
  assign n5461 = n5453 & ~n5456 ;
  assign n5462 = n5424 & n5427 ;
  assign n5463 = ~n5461 & ~n5462 ;
  assign n5464 = ~n5460 & n5463 ;
  assign n5465 = ~n5429 & ~n5464 ;
  assign n5466 = ~n5428 & n5465 ;
  assign n5467 = ~n5425 & ~n5466 ;
  assign n5468 = ~n5424 & ~n5467 ;
  assign n5469 = n5427 & ~n5465 ;
  assign n5470 = ~n5468 & ~n5469 ;
  assign n5471 = ~n3392 & n3675 ;
  assign n5472 = n3665 & ~n3671 ;
  assign n5473 = ~n3672 & ~n5472 ;
  assign n5474 = ~n5431 & n5467 ;
  assign n5475 = ~n5434 & ~n5467 ;
  assign n5476 = ~n5474 & ~n5475 ;
  assign n5477 = ~n5473 & n5476 ;
  assign n5478 = n3667 & ~n3670 ;
  assign n5479 = ~n3671 & ~n5478 ;
  assign n5480 = n5440 & ~n5467 ;
  assign n5481 = n5437 & n5467 ;
  assign n5482 = ~n5480 & ~n5481 ;
  assign n5483 = n5479 & n5482 ;
  assign n5484 = ~n5477 & n5483 ;
  assign n5485 = n3663 & ~n3672 ;
  assign n5486 = ~n3673 & ~n5485 ;
  assign n5487 = ~n5444 & n5467 ;
  assign n5488 = n5447 & ~n5467 ;
  assign n5489 = ~n5487 & ~n5488 ;
  assign n5490 = n5486 & ~n5489 ;
  assign n5491 = n5473 & ~n5476 ;
  assign n5492 = ~n5490 & ~n5491 ;
  assign n5493 = ~n5484 & n5492 ;
  assign n5494 = n3661 & ~n3673 ;
  assign n5495 = ~n3674 & ~n5494 ;
  assign n5496 = ~n5453 & n5467 ;
  assign n5497 = ~n5456 & ~n5467 ;
  assign n5498 = ~n5496 & ~n5497 ;
  assign n5499 = ~n5495 & n5498 ;
  assign n5500 = ~n5486 & n5489 ;
  assign n5501 = ~n5499 & ~n5500 ;
  assign n5502 = ~n5493 & n5501 ;
  assign n5503 = ~n3659 & ~n3674 ;
  assign n5504 = ~n3675 & ~n5503 ;
  assign n5505 = n5470 & n5504 ;
  assign n5506 = n5495 & ~n5498 ;
  assign n5507 = ~n5505 & ~n5506 ;
  assign n5508 = ~n5502 & n5507 ;
  assign n5509 = n3392 & ~n3675 ;
  assign n5510 = ~n5470 & ~n5504 ;
  assign n5511 = ~n5509 & ~n5510 ;
  assign n5512 = ~n5508 & n5511 ;
  assign n5513 = ~n5471 & ~n5512 ;
  assign n5514 = ~n5470 & ~n5513 ;
  assign n5515 = n5504 & ~n5512 ;
  assign n5516 = ~n5514 & ~n5515 ;
  assign n5517 = ~n3676 & n3959 ;
  assign n5518 = ~n3943 & ~n3958 ;
  assign n5519 = ~n3959 & ~n5518 ;
  assign n5520 = ~n5516 & ~n5519 ;
  assign n5521 = n3676 & ~n3959 ;
  assign n5522 = n3949 & ~n3955 ;
  assign n5523 = ~n3956 & ~n5522 ;
  assign n5524 = ~n5473 & n5513 ;
  assign n5525 = ~n5476 & ~n5513 ;
  assign n5526 = ~n5524 & ~n5525 ;
  assign n5527 = ~n5523 & n5526 ;
  assign n5528 = n3951 & ~n3954 ;
  assign n5529 = ~n3955 & ~n5528 ;
  assign n5530 = n5482 & ~n5513 ;
  assign n5531 = ~n5479 & n5513 ;
  assign n5532 = ~n5530 & ~n5531 ;
  assign n5533 = n5529 & ~n5532 ;
  assign n5534 = ~n5527 & n5533 ;
  assign n5535 = n3947 & ~n3956 ;
  assign n5536 = ~n3957 & ~n5535 ;
  assign n5537 = n5489 & ~n5513 ;
  assign n5538 = n5486 & n5513 ;
  assign n5539 = ~n5537 & ~n5538 ;
  assign n5540 = n5536 & n5539 ;
  assign n5541 = n5523 & ~n5526 ;
  assign n5542 = ~n5540 & ~n5541 ;
  assign n5543 = ~n5534 & n5542 ;
  assign n5544 = n3945 & ~n3957 ;
  assign n5545 = ~n3958 & ~n5544 ;
  assign n5546 = ~n5495 & n5513 ;
  assign n5547 = ~n5498 & ~n5513 ;
  assign n5548 = ~n5546 & ~n5547 ;
  assign n5549 = ~n5545 & n5548 ;
  assign n5550 = ~n5536 & ~n5539 ;
  assign n5551 = ~n5549 & ~n5550 ;
  assign n5552 = ~n5543 & n5551 ;
  assign n5553 = n5545 & ~n5548 ;
  assign n5554 = n5516 & n5519 ;
  assign n5555 = ~n5553 & ~n5554 ;
  assign n5556 = ~n5552 & n5555 ;
  assign n5557 = ~n5521 & ~n5556 ;
  assign n5558 = ~n5520 & n5557 ;
  assign n5559 = ~n5517 & ~n5558 ;
  assign n5560 = ~n5516 & ~n5559 ;
  assign n5561 = n5519 & ~n5557 ;
  assign n5562 = ~n5560 & ~n5561 ;
  assign n5563 = ~n3960 & n4243 ;
  assign n5564 = n4233 & ~n4239 ;
  assign n5565 = ~n4240 & ~n5564 ;
  assign n5566 = ~n5523 & n5559 ;
  assign n5567 = ~n5526 & ~n5559 ;
  assign n5568 = ~n5566 & ~n5567 ;
  assign n5569 = ~n5565 & n5568 ;
  assign n5570 = n4235 & ~n4238 ;
  assign n5571 = ~n4239 & ~n5570 ;
  assign n5572 = n5532 & ~n5559 ;
  assign n5573 = n5529 & n5559 ;
  assign n5574 = ~n5572 & ~n5573 ;
  assign n5575 = n5571 & n5574 ;
  assign n5576 = ~n5569 & n5575 ;
  assign n5577 = n4231 & ~n4240 ;
  assign n5578 = ~n4241 & ~n5577 ;
  assign n5579 = ~n5536 & n5559 ;
  assign n5580 = n5539 & ~n5559 ;
  assign n5581 = ~n5579 & ~n5580 ;
  assign n5582 = n5578 & ~n5581 ;
  assign n5583 = n5565 & ~n5568 ;
  assign n5584 = ~n5582 & ~n5583 ;
  assign n5585 = ~n5576 & n5584 ;
  assign n5586 = n4229 & ~n4241 ;
  assign n5587 = ~n4242 & ~n5586 ;
  assign n5588 = ~n5545 & n5559 ;
  assign n5589 = ~n5548 & ~n5559 ;
  assign n5590 = ~n5588 & ~n5589 ;
  assign n5591 = ~n5587 & n5590 ;
  assign n5592 = ~n5578 & n5581 ;
  assign n5593 = ~n5591 & ~n5592 ;
  assign n5594 = ~n5585 & n5593 ;
  assign n5595 = ~n4227 & ~n4242 ;
  assign n5596 = ~n4243 & ~n5595 ;
  assign n5597 = n5562 & n5596 ;
  assign n5598 = n5587 & ~n5590 ;
  assign n5599 = ~n5597 & ~n5598 ;
  assign n5600 = ~n5594 & n5599 ;
  assign n5601 = n3960 & ~n4243 ;
  assign n5602 = ~n5562 & ~n5596 ;
  assign n5603 = ~n5601 & ~n5602 ;
  assign n5604 = ~n5600 & n5603 ;
  assign n5605 = ~n5563 & ~n5604 ;
  assign n5606 = ~n5562 & ~n5605 ;
  assign n5607 = n5596 & ~n5604 ;
  assign n5608 = ~n5606 & ~n5607 ;
  assign n5609 = ~n4511 & ~n4526 ;
  assign n5610 = ~n4527 & ~n5609 ;
  assign n5611 = ~n5608 & ~n5610 ;
  assign n5612 = n4244 & ~n4527 ;
  assign n5613 = ~n5565 & n5605 ;
  assign n5614 = ~n5568 & ~n5605 ;
  assign n5615 = ~n5613 & ~n5614 ;
  assign n5616 = ~n5104 & n5615 ;
  assign n5617 = n4519 & ~n4522 ;
  assign n5618 = ~n4523 & ~n5617 ;
  assign n5619 = n5574 & ~n5605 ;
  assign n5620 = ~n5571 & n5605 ;
  assign n5621 = ~n5619 & ~n5620 ;
  assign n5622 = n5618 & ~n5621 ;
  assign n5623 = ~n5616 & n5622 ;
  assign n5624 = n4515 & ~n4524 ;
  assign n5625 = ~n4525 & ~n5624 ;
  assign n5626 = n5581 & ~n5605 ;
  assign n5627 = n5578 & n5605 ;
  assign n5628 = ~n5626 & ~n5627 ;
  assign n5629 = n5625 & n5628 ;
  assign n5630 = n5104 & ~n5615 ;
  assign n5631 = ~n5629 & ~n5630 ;
  assign n5632 = ~n5623 & n5631 ;
  assign n5633 = n4513 & ~n4525 ;
  assign n5634 = ~n4526 & ~n5633 ;
  assign n5635 = ~n5587 & n5605 ;
  assign n5636 = ~n5590 & ~n5605 ;
  assign n5637 = ~n5635 & ~n5636 ;
  assign n5638 = ~n5634 & n5637 ;
  assign n5639 = ~n5625 & ~n5628 ;
  assign n5640 = ~n5638 & ~n5639 ;
  assign n5641 = ~n5632 & n5640 ;
  assign n5642 = n5634 & ~n5637 ;
  assign n5643 = n5608 & n5610 ;
  assign n5644 = ~n5642 & ~n5643 ;
  assign n5645 = ~n5641 & n5644 ;
  assign n5646 = ~n5612 & ~n5645 ;
  assign n5647 = ~n5611 & n5646 ;
  assign n5648 = ~n5105 & ~n5647 ;
  assign n5649 = ~n5104 & n5648 ;
  assign n5650 = ~n5615 & ~n5648 ;
  assign n5651 = ~n5649 & ~n5650 ;
  assign n5652 = ~n5101 & n5651 ;
  assign n5653 = n4801 & ~n4804 ;
  assign n5654 = ~n4805 & ~n5653 ;
  assign n5655 = n5621 & ~n5648 ;
  assign n5656 = n5618 & n5648 ;
  assign n5657 = ~n5655 & ~n5656 ;
  assign n5658 = n5654 & n5657 ;
  assign n5659 = ~n5652 & n5658 ;
  assign n5660 = n4799 & ~n4808 ;
  assign n5661 = ~n4809 & ~n5660 ;
  assign n5662 = ~n5625 & n5648 ;
  assign n5663 = n5628 & ~n5648 ;
  assign n5664 = ~n5662 & ~n5663 ;
  assign n5665 = n5661 & ~n5664 ;
  assign n5666 = n5101 & ~n5651 ;
  assign n5667 = ~n5665 & ~n5666 ;
  assign n5668 = ~n5659 & n5667 ;
  assign n5669 = n4797 & ~n4809 ;
  assign n5670 = ~n4810 & ~n5669 ;
  assign n5671 = ~n5634 & n5648 ;
  assign n5672 = ~n5637 & ~n5648 ;
  assign n5673 = ~n5671 & ~n5672 ;
  assign n5674 = ~n5670 & n5673 ;
  assign n5675 = ~n5661 & n5664 ;
  assign n5676 = ~n5674 & ~n5675 ;
  assign n5677 = ~n5668 & n5676 ;
  assign n5678 = ~n5608 & ~n5648 ;
  assign n5679 = n5610 & ~n5646 ;
  assign n5680 = ~n5678 & ~n5679 ;
  assign n5681 = ~n4795 & ~n4810 ;
  assign n5682 = ~n4811 & ~n5681 ;
  assign n5683 = n5680 & n5682 ;
  assign n5684 = n5670 & ~n5673 ;
  assign n5685 = ~n5683 & ~n5684 ;
  assign n5686 = ~n5677 & n5685 ;
  assign n5687 = n4528 & ~n4811 ;
  assign n5688 = ~n5680 & ~n5682 ;
  assign n5689 = ~n5687 & ~n5688 ;
  assign n5690 = ~n5686 & n5689 ;
  assign n5691 = ~n5102 & ~n5690 ;
  assign n5692 = ~n5101 & n5691 ;
  assign n5693 = ~n5651 & ~n5691 ;
  assign n5694 = ~n5692 & ~n5693 ;
  assign n5695 = ~n4812 & n5095 ;
  assign n5696 = ~n5680 & ~n5691 ;
  assign n5697 = n5682 & ~n5690 ;
  assign n5698 = ~n5696 & ~n5697 ;
  assign n5699 = ~n5079 & ~n5094 ;
  assign n5700 = ~n5095 & ~n5699 ;
  assign n5701 = ~n5698 & ~n5700 ;
  assign n5702 = n4812 & ~n5095 ;
  assign n5703 = ~n5089 & n5091 ;
  assign n5704 = ~n5092 & ~n5703 ;
  assign n5705 = n5694 & ~n5704 ;
  assign n5706 = n5085 & ~n5088 ;
  assign n5707 = ~n5089 & ~n5706 ;
  assign n5708 = n5657 & ~n5691 ;
  assign n5709 = ~n5654 & n5691 ;
  assign n5710 = ~n5708 & ~n5709 ;
  assign n5711 = n5707 & ~n5710 ;
  assign n5712 = ~n5705 & n5711 ;
  assign n5713 = n5083 & ~n5092 ;
  assign n5714 = ~n5093 & ~n5713 ;
  assign n5715 = n5664 & ~n5691 ;
  assign n5716 = n5661 & n5691 ;
  assign n5717 = ~n5715 & ~n5716 ;
  assign n5718 = n5714 & n5717 ;
  assign n5719 = ~n5694 & n5704 ;
  assign n5720 = ~n5718 & ~n5719 ;
  assign n5721 = ~n5712 & n5720 ;
  assign n5722 = n5081 & ~n5093 ;
  assign n5723 = ~n5094 & ~n5722 ;
  assign n5724 = ~n5670 & n5691 ;
  assign n5725 = ~n5673 & ~n5691 ;
  assign n5726 = ~n5724 & ~n5725 ;
  assign n5727 = ~n5723 & n5726 ;
  assign n5728 = ~n5714 & ~n5717 ;
  assign n5729 = ~n5727 & ~n5728 ;
  assign n5730 = ~n5721 & n5729 ;
  assign n5731 = n5723 & ~n5726 ;
  assign n5732 = n5698 & n5700 ;
  assign n5733 = ~n5731 & ~n5732 ;
  assign n5734 = ~n5730 & n5733 ;
  assign n5735 = ~n5702 & ~n5734 ;
  assign n5736 = ~n5701 & n5735 ;
  assign n5737 = ~n5695 & ~n5736 ;
  assign n5738 = n5694 & ~n5737 ;
  assign n5739 = n5704 & n5737 ;
  assign n5740 = ~n5738 & ~n5739 ;
  assign n5741 = n5099 & n5740 ;
  assign n5742 = n5710 & ~n5737 ;
  assign n5743 = n5707 & n5737 ;
  assign n5744 = n818 & ~n821 ;
  assign n5745 = ~n822 & ~n5744 ;
  assign n5746 = ~n5743 & n5745 ;
  assign n5747 = ~n5742 & n5746 ;
  assign n5748 = ~n5741 & ~n5747 ;
  assign n5749 = ~n5099 & ~n5740 ;
  assign n5750 = n814 & ~n823 ;
  assign n5751 = ~n824 & ~n5750 ;
  assign n5752 = ~n5717 & ~n5737 ;
  assign n5753 = n5714 & n5737 ;
  assign n5754 = ~n5752 & ~n5753 ;
  assign n5755 = ~n5751 & ~n5754 ;
  assign n5756 = ~n5749 & ~n5755 ;
  assign n5757 = ~n5748 & n5756 ;
  assign n5758 = n812 & ~n824 ;
  assign n5759 = ~n825 & ~n5758 ;
  assign n5760 = ~n5723 & n5737 ;
  assign n5761 = ~n5726 & ~n5737 ;
  assign n5762 = ~n5760 & ~n5761 ;
  assign n5763 = n5759 & ~n5762 ;
  assign n5764 = n5751 & n5754 ;
  assign n5765 = ~n5763 & ~n5764 ;
  assign n5766 = ~n5757 & n5765 ;
  assign n5767 = ~n5759 & n5762 ;
  assign n5768 = ~n825 & ~n826 ;
  assign n5769 = ~n827 & ~n5768 ;
  assign n5770 = ~n5698 & ~n5737 ;
  assign n5771 = n5700 & ~n5735 ;
  assign n5772 = ~n5770 & ~n5771 ;
  assign n5773 = ~n5769 & ~n5772 ;
  assign n5774 = ~n5767 & ~n5773 ;
  assign n5775 = ~n5766 & n5774 ;
  assign n5776 = n827 & ~n5096 ;
  assign n5777 = n5769 & n5772 ;
  assign n5778 = ~n5776 & ~n5777 ;
  assign n5779 = ~n5775 & n5778 ;
  assign n5780 = ~n5097 & ~n5779 ;
  assign n5781 = ~x0 & ~n5780 ;
  assign n5782 = ~x32 & n5737 ;
  assign n5783 = ~x192 & n5513 ;
  assign n5784 = ~x320 & n5329 ;
  assign n5785 = ~x416 & n5191 ;
  assign n5786 = x448 & ~n5155 ;
  assign n5787 = x480 & n5155 ;
  assign n5788 = ~n5786 & ~n5787 ;
  assign n5789 = ~n5191 & n5788 ;
  assign n5790 = ~n5785 & ~n5789 ;
  assign n5791 = ~n5237 & n5790 ;
  assign n5792 = x384 & n5237 ;
  assign n5793 = ~n5791 & ~n5792 ;
  assign n5794 = ~n5283 & ~n5793 ;
  assign n5795 = x352 & n5283 ;
  assign n5796 = ~n5794 & ~n5795 ;
  assign n5797 = ~n5329 & n5796 ;
  assign n5798 = ~n5784 & ~n5797 ;
  assign n5799 = ~n5375 & ~n5798 ;
  assign n5800 = ~x288 & n5375 ;
  assign n5801 = ~n5799 & ~n5800 ;
  assign n5802 = ~n5421 & ~n5801 ;
  assign n5803 = ~x256 & n5421 ;
  assign n5804 = ~n5802 & ~n5803 ;
  assign n5805 = ~n5467 & n5804 ;
  assign n5806 = x224 & n5467 ;
  assign n5807 = ~n5805 & ~n5806 ;
  assign n5808 = ~n5513 & n5807 ;
  assign n5809 = ~n5783 & ~n5808 ;
  assign n5810 = ~n5559 & ~n5809 ;
  assign n5811 = ~x160 & n5559 ;
  assign n5812 = ~n5810 & ~n5811 ;
  assign n5813 = ~n5605 & n5812 ;
  assign n5814 = x128 & n5605 ;
  assign n5815 = ~n5813 & ~n5814 ;
  assign n5816 = ~n5648 & ~n5815 ;
  assign n5817 = x96 & n5648 ;
  assign n5818 = ~n5816 & ~n5817 ;
  assign n5819 = ~n5691 & ~n5818 ;
  assign n5820 = x64 & n5691 ;
  assign n5821 = ~n5819 & ~n5820 ;
  assign n5822 = ~n5737 & n5821 ;
  assign n5823 = ~n5782 & ~n5822 ;
  assign n5824 = n5780 & ~n5823 ;
  assign n5825 = ~n5781 & ~n5824 ;
  assign n5826 = ~x1 & ~n5780 ;
  assign n5827 = ~x33 & n5737 ;
  assign n5828 = ~x193 & n5513 ;
  assign n5829 = ~x321 & n5329 ;
  assign n5830 = ~x417 & n5191 ;
  assign n5831 = x449 & ~n5155 ;
  assign n5832 = x481 & n5155 ;
  assign n5833 = ~n5831 & ~n5832 ;
  assign n5834 = ~n5191 & n5833 ;
  assign n5835 = ~n5830 & ~n5834 ;
  assign n5836 = ~n5237 & n5835 ;
  assign n5837 = x385 & n5237 ;
  assign n5838 = ~n5836 & ~n5837 ;
  assign n5839 = ~n5283 & ~n5838 ;
  assign n5840 = x353 & n5283 ;
  assign n5841 = ~n5839 & ~n5840 ;
  assign n5842 = ~n5329 & n5841 ;
  assign n5843 = ~n5829 & ~n5842 ;
  assign n5844 = ~n5375 & ~n5843 ;
  assign n5845 = ~x289 & n5375 ;
  assign n5846 = ~n5844 & ~n5845 ;
  assign n5847 = ~n5421 & ~n5846 ;
  assign n5848 = ~x257 & n5421 ;
  assign n5849 = ~n5847 & ~n5848 ;
  assign n5850 = ~n5467 & n5849 ;
  assign n5851 = x225 & n5467 ;
  assign n5852 = ~n5850 & ~n5851 ;
  assign n5853 = ~n5513 & n5852 ;
  assign n5854 = ~n5828 & ~n5853 ;
  assign n5855 = ~n5559 & ~n5854 ;
  assign n5856 = ~x161 & n5559 ;
  assign n5857 = ~n5855 & ~n5856 ;
  assign n5858 = ~n5605 & n5857 ;
  assign n5859 = x129 & n5605 ;
  assign n5860 = ~n5858 & ~n5859 ;
  assign n5861 = ~n5648 & ~n5860 ;
  assign n5862 = x97 & n5648 ;
  assign n5863 = ~n5861 & ~n5862 ;
  assign n5864 = ~n5691 & ~n5863 ;
  assign n5865 = x65 & n5691 ;
  assign n5866 = ~n5864 & ~n5865 ;
  assign n5867 = ~n5737 & n5866 ;
  assign n5868 = ~n5827 & ~n5867 ;
  assign n5869 = n5780 & ~n5868 ;
  assign n5870 = ~n5826 & ~n5869 ;
  assign n5871 = ~x2 & ~n5780 ;
  assign n5872 = ~x34 & n5737 ;
  assign n5873 = ~x194 & n5513 ;
  assign n5874 = ~x322 & n5329 ;
  assign n5875 = ~x418 & n5191 ;
  assign n5876 = x450 & ~n5155 ;
  assign n5877 = x482 & n5155 ;
  assign n5878 = ~n5876 & ~n5877 ;
  assign n5879 = ~n5191 & n5878 ;
  assign n5880 = ~n5875 & ~n5879 ;
  assign n5881 = ~n5237 & n5880 ;
  assign n5882 = x386 & n5237 ;
  assign n5883 = ~n5881 & ~n5882 ;
  assign n5884 = ~n5283 & ~n5883 ;
  assign n5885 = x354 & n5283 ;
  assign n5886 = ~n5884 & ~n5885 ;
  assign n5887 = ~n5329 & n5886 ;
  assign n5888 = ~n5874 & ~n5887 ;
  assign n5889 = ~n5375 & ~n5888 ;
  assign n5890 = ~x290 & n5375 ;
  assign n5891 = ~n5889 & ~n5890 ;
  assign n5892 = ~n5421 & ~n5891 ;
  assign n5893 = ~x258 & n5421 ;
  assign n5894 = ~n5892 & ~n5893 ;
  assign n5895 = ~n5467 & n5894 ;
  assign n5896 = x226 & n5467 ;
  assign n5897 = ~n5895 & ~n5896 ;
  assign n5898 = ~n5513 & n5897 ;
  assign n5899 = ~n5873 & ~n5898 ;
  assign n5900 = ~n5559 & ~n5899 ;
  assign n5901 = ~x162 & n5559 ;
  assign n5902 = ~n5900 & ~n5901 ;
  assign n5903 = ~n5605 & n5902 ;
  assign n5904 = x130 & n5605 ;
  assign n5905 = ~n5903 & ~n5904 ;
  assign n5906 = ~n5648 & ~n5905 ;
  assign n5907 = x98 & n5648 ;
  assign n5908 = ~n5906 & ~n5907 ;
  assign n5909 = ~n5691 & ~n5908 ;
  assign n5910 = x66 & n5691 ;
  assign n5911 = ~n5909 & ~n5910 ;
  assign n5912 = ~n5737 & n5911 ;
  assign n5913 = ~n5872 & ~n5912 ;
  assign n5914 = n5780 & ~n5913 ;
  assign n5915 = ~n5871 & ~n5914 ;
  assign n5916 = ~x3 & ~n5780 ;
  assign n5917 = ~x35 & n5737 ;
  assign n5918 = ~x195 & n5513 ;
  assign n5919 = ~x323 & n5329 ;
  assign n5920 = ~x419 & n5191 ;
  assign n5921 = x451 & ~n5155 ;
  assign n5922 = x483 & n5155 ;
  assign n5923 = ~n5921 & ~n5922 ;
  assign n5924 = ~n5191 & n5923 ;
  assign n5925 = ~n5920 & ~n5924 ;
  assign n5926 = ~n5237 & n5925 ;
  assign n5927 = x387 & n5237 ;
  assign n5928 = ~n5926 & ~n5927 ;
  assign n5929 = ~n5283 & ~n5928 ;
  assign n5930 = x355 & n5283 ;
  assign n5931 = ~n5929 & ~n5930 ;
  assign n5932 = ~n5329 & n5931 ;
  assign n5933 = ~n5919 & ~n5932 ;
  assign n5934 = ~n5375 & ~n5933 ;
  assign n5935 = ~x291 & n5375 ;
  assign n5936 = ~n5934 & ~n5935 ;
  assign n5937 = ~n5421 & ~n5936 ;
  assign n5938 = ~x259 & n5421 ;
  assign n5939 = ~n5937 & ~n5938 ;
  assign n5940 = ~n5467 & n5939 ;
  assign n5941 = x227 & n5467 ;
  assign n5942 = ~n5940 & ~n5941 ;
  assign n5943 = ~n5513 & n5942 ;
  assign n5944 = ~n5918 & ~n5943 ;
  assign n5945 = ~n5559 & ~n5944 ;
  assign n5946 = ~x163 & n5559 ;
  assign n5947 = ~n5945 & ~n5946 ;
  assign n5948 = ~n5605 & n5947 ;
  assign n5949 = x131 & n5605 ;
  assign n5950 = ~n5948 & ~n5949 ;
  assign n5951 = ~n5648 & ~n5950 ;
  assign n5952 = x99 & n5648 ;
  assign n5953 = ~n5951 & ~n5952 ;
  assign n5954 = ~n5691 & ~n5953 ;
  assign n5955 = x67 & n5691 ;
  assign n5956 = ~n5954 & ~n5955 ;
  assign n5957 = ~n5737 & n5956 ;
  assign n5958 = ~n5917 & ~n5957 ;
  assign n5959 = n5780 & ~n5958 ;
  assign n5960 = ~n5916 & ~n5959 ;
  assign n5961 = ~x4 & ~n5780 ;
  assign n5962 = ~x36 & n5737 ;
  assign n5963 = ~x196 & n5513 ;
  assign n5964 = ~x324 & n5329 ;
  assign n5965 = ~x420 & n5191 ;
  assign n5966 = x452 & ~n5155 ;
  assign n5967 = x484 & n5155 ;
  assign n5968 = ~n5966 & ~n5967 ;
  assign n5969 = ~n5191 & n5968 ;
  assign n5970 = ~n5965 & ~n5969 ;
  assign n5971 = ~n5237 & n5970 ;
  assign n5972 = x388 & n5237 ;
  assign n5973 = ~n5971 & ~n5972 ;
  assign n5974 = ~n5283 & ~n5973 ;
  assign n5975 = x356 & n5283 ;
  assign n5976 = ~n5974 & ~n5975 ;
  assign n5977 = ~n5329 & n5976 ;
  assign n5978 = ~n5964 & ~n5977 ;
  assign n5979 = ~n5375 & ~n5978 ;
  assign n5980 = ~x292 & n5375 ;
  assign n5981 = ~n5979 & ~n5980 ;
  assign n5982 = ~n5421 & ~n5981 ;
  assign n5983 = ~x260 & n5421 ;
  assign n5984 = ~n5982 & ~n5983 ;
  assign n5985 = ~n5467 & n5984 ;
  assign n5986 = x228 & n5467 ;
  assign n5987 = ~n5985 & ~n5986 ;
  assign n5988 = ~n5513 & n5987 ;
  assign n5989 = ~n5963 & ~n5988 ;
  assign n5990 = ~n5559 & ~n5989 ;
  assign n5991 = ~x164 & n5559 ;
  assign n5992 = ~n5990 & ~n5991 ;
  assign n5993 = ~n5605 & n5992 ;
  assign n5994 = x132 & n5605 ;
  assign n5995 = ~n5993 & ~n5994 ;
  assign n5996 = ~n5648 & ~n5995 ;
  assign n5997 = x100 & n5648 ;
  assign n5998 = ~n5996 & ~n5997 ;
  assign n5999 = ~n5691 & ~n5998 ;
  assign n6000 = x68 & n5691 ;
  assign n6001 = ~n5999 & ~n6000 ;
  assign n6002 = ~n5737 & n6001 ;
  assign n6003 = ~n5962 & ~n6002 ;
  assign n6004 = n5780 & ~n6003 ;
  assign n6005 = ~n5961 & ~n6004 ;
  assign n6006 = ~x5 & ~n5780 ;
  assign n6007 = ~x37 & n5737 ;
  assign n6008 = ~x197 & n5513 ;
  assign n6009 = ~x325 & n5329 ;
  assign n6010 = ~x421 & n5191 ;
  assign n6011 = x453 & ~n5155 ;
  assign n6012 = x485 & n5155 ;
  assign n6013 = ~n6011 & ~n6012 ;
  assign n6014 = ~n5191 & n6013 ;
  assign n6015 = ~n6010 & ~n6014 ;
  assign n6016 = ~n5237 & n6015 ;
  assign n6017 = x389 & n5237 ;
  assign n6018 = ~n6016 & ~n6017 ;
  assign n6019 = ~n5283 & ~n6018 ;
  assign n6020 = x357 & n5283 ;
  assign n6021 = ~n6019 & ~n6020 ;
  assign n6022 = ~n5329 & n6021 ;
  assign n6023 = ~n6009 & ~n6022 ;
  assign n6024 = ~n5375 & ~n6023 ;
  assign n6025 = ~x293 & n5375 ;
  assign n6026 = ~n6024 & ~n6025 ;
  assign n6027 = ~n5421 & ~n6026 ;
  assign n6028 = ~x261 & n5421 ;
  assign n6029 = ~n6027 & ~n6028 ;
  assign n6030 = ~n5467 & n6029 ;
  assign n6031 = x229 & n5467 ;
  assign n6032 = ~n6030 & ~n6031 ;
  assign n6033 = ~n5513 & n6032 ;
  assign n6034 = ~n6008 & ~n6033 ;
  assign n6035 = ~n5559 & ~n6034 ;
  assign n6036 = ~x165 & n5559 ;
  assign n6037 = ~n6035 & ~n6036 ;
  assign n6038 = ~n5605 & n6037 ;
  assign n6039 = x133 & n5605 ;
  assign n6040 = ~n6038 & ~n6039 ;
  assign n6041 = ~n5648 & ~n6040 ;
  assign n6042 = x101 & n5648 ;
  assign n6043 = ~n6041 & ~n6042 ;
  assign n6044 = ~n5691 & ~n6043 ;
  assign n6045 = x69 & n5691 ;
  assign n6046 = ~n6044 & ~n6045 ;
  assign n6047 = ~n5737 & n6046 ;
  assign n6048 = ~n6007 & ~n6047 ;
  assign n6049 = n5780 & ~n6048 ;
  assign n6050 = ~n6006 & ~n6049 ;
  assign n6051 = ~x6 & ~n5780 ;
  assign n6052 = ~x38 & n5737 ;
  assign n6053 = ~x198 & n5513 ;
  assign n6054 = ~x326 & n5329 ;
  assign n6055 = ~x422 & n5191 ;
  assign n6056 = x454 & ~n5155 ;
  assign n6057 = x486 & n5155 ;
  assign n6058 = ~n6056 & ~n6057 ;
  assign n6059 = ~n5191 & n6058 ;
  assign n6060 = ~n6055 & ~n6059 ;
  assign n6061 = ~n5237 & n6060 ;
  assign n6062 = x390 & n5237 ;
  assign n6063 = ~n6061 & ~n6062 ;
  assign n6064 = ~n5283 & ~n6063 ;
  assign n6065 = x358 & n5283 ;
  assign n6066 = ~n6064 & ~n6065 ;
  assign n6067 = ~n5329 & n6066 ;
  assign n6068 = ~n6054 & ~n6067 ;
  assign n6069 = ~n5375 & ~n6068 ;
  assign n6070 = ~x294 & n5375 ;
  assign n6071 = ~n6069 & ~n6070 ;
  assign n6072 = ~n5421 & ~n6071 ;
  assign n6073 = ~x262 & n5421 ;
  assign n6074 = ~n6072 & ~n6073 ;
  assign n6075 = ~n5467 & n6074 ;
  assign n6076 = x230 & n5467 ;
  assign n6077 = ~n6075 & ~n6076 ;
  assign n6078 = ~n5513 & n6077 ;
  assign n6079 = ~n6053 & ~n6078 ;
  assign n6080 = ~n5559 & ~n6079 ;
  assign n6081 = ~x166 & n5559 ;
  assign n6082 = ~n6080 & ~n6081 ;
  assign n6083 = ~n5605 & n6082 ;
  assign n6084 = x134 & n5605 ;
  assign n6085 = ~n6083 & ~n6084 ;
  assign n6086 = ~n5648 & ~n6085 ;
  assign n6087 = x102 & n5648 ;
  assign n6088 = ~n6086 & ~n6087 ;
  assign n6089 = ~n5691 & ~n6088 ;
  assign n6090 = x70 & n5691 ;
  assign n6091 = ~n6089 & ~n6090 ;
  assign n6092 = ~n5737 & n6091 ;
  assign n6093 = ~n6052 & ~n6092 ;
  assign n6094 = n5780 & ~n6093 ;
  assign n6095 = ~n6051 & ~n6094 ;
  assign n6096 = ~x7 & ~n5780 ;
  assign n6097 = ~x39 & n5737 ;
  assign n6098 = ~x199 & n5513 ;
  assign n6099 = ~x327 & n5329 ;
  assign n6100 = ~x423 & n5191 ;
  assign n6101 = x455 & ~n5155 ;
  assign n6102 = x487 & n5155 ;
  assign n6103 = ~n6101 & ~n6102 ;
  assign n6104 = ~n5191 & n6103 ;
  assign n6105 = ~n6100 & ~n6104 ;
  assign n6106 = ~n5237 & n6105 ;
  assign n6107 = x391 & n5237 ;
  assign n6108 = ~n6106 & ~n6107 ;
  assign n6109 = ~n5283 & ~n6108 ;
  assign n6110 = x359 & n5283 ;
  assign n6111 = ~n6109 & ~n6110 ;
  assign n6112 = ~n5329 & n6111 ;
  assign n6113 = ~n6099 & ~n6112 ;
  assign n6114 = ~n5375 & ~n6113 ;
  assign n6115 = ~x295 & n5375 ;
  assign n6116 = ~n6114 & ~n6115 ;
  assign n6117 = ~n5421 & ~n6116 ;
  assign n6118 = ~x263 & n5421 ;
  assign n6119 = ~n6117 & ~n6118 ;
  assign n6120 = ~n5467 & n6119 ;
  assign n6121 = x231 & n5467 ;
  assign n6122 = ~n6120 & ~n6121 ;
  assign n6123 = ~n5513 & n6122 ;
  assign n6124 = ~n6098 & ~n6123 ;
  assign n6125 = ~n5559 & ~n6124 ;
  assign n6126 = ~x167 & n5559 ;
  assign n6127 = ~n6125 & ~n6126 ;
  assign n6128 = ~n5605 & n6127 ;
  assign n6129 = x135 & n5605 ;
  assign n6130 = ~n6128 & ~n6129 ;
  assign n6131 = ~n5648 & ~n6130 ;
  assign n6132 = x103 & n5648 ;
  assign n6133 = ~n6131 & ~n6132 ;
  assign n6134 = ~n5691 & ~n6133 ;
  assign n6135 = x71 & n5691 ;
  assign n6136 = ~n6134 & ~n6135 ;
  assign n6137 = ~n5737 & n6136 ;
  assign n6138 = ~n6097 & ~n6137 ;
  assign n6139 = n5780 & ~n6138 ;
  assign n6140 = ~n6096 & ~n6139 ;
  assign n6141 = ~x8 & ~n5780 ;
  assign n6142 = ~x40 & n5737 ;
  assign n6143 = ~x200 & n5513 ;
  assign n6144 = ~x328 & n5329 ;
  assign n6145 = ~x424 & n5191 ;
  assign n6146 = x456 & ~n5155 ;
  assign n6147 = x488 & n5155 ;
  assign n6148 = ~n6146 & ~n6147 ;
  assign n6149 = ~n5191 & n6148 ;
  assign n6150 = ~n6145 & ~n6149 ;
  assign n6151 = ~n5237 & n6150 ;
  assign n6152 = x392 & n5237 ;
  assign n6153 = ~n6151 & ~n6152 ;
  assign n6154 = ~n5283 & ~n6153 ;
  assign n6155 = x360 & n5283 ;
  assign n6156 = ~n6154 & ~n6155 ;
  assign n6157 = ~n5329 & n6156 ;
  assign n6158 = ~n6144 & ~n6157 ;
  assign n6159 = ~n5375 & ~n6158 ;
  assign n6160 = ~x296 & n5375 ;
  assign n6161 = ~n6159 & ~n6160 ;
  assign n6162 = ~n5421 & ~n6161 ;
  assign n6163 = ~x264 & n5421 ;
  assign n6164 = ~n6162 & ~n6163 ;
  assign n6165 = ~n5467 & n6164 ;
  assign n6166 = x232 & n5467 ;
  assign n6167 = ~n6165 & ~n6166 ;
  assign n6168 = ~n5513 & n6167 ;
  assign n6169 = ~n6143 & ~n6168 ;
  assign n6170 = ~n5559 & ~n6169 ;
  assign n6171 = ~x168 & n5559 ;
  assign n6172 = ~n6170 & ~n6171 ;
  assign n6173 = ~n5605 & n6172 ;
  assign n6174 = x136 & n5605 ;
  assign n6175 = ~n6173 & ~n6174 ;
  assign n6176 = ~n5648 & ~n6175 ;
  assign n6177 = x104 & n5648 ;
  assign n6178 = ~n6176 & ~n6177 ;
  assign n6179 = ~n5691 & ~n6178 ;
  assign n6180 = x72 & n5691 ;
  assign n6181 = ~n6179 & ~n6180 ;
  assign n6182 = ~n5737 & n6181 ;
  assign n6183 = ~n6142 & ~n6182 ;
  assign n6184 = n5780 & ~n6183 ;
  assign n6185 = ~n6141 & ~n6184 ;
  assign n6186 = ~x9 & ~n5780 ;
  assign n6187 = ~x41 & n5737 ;
  assign n6188 = ~x201 & n5513 ;
  assign n6189 = ~x329 & n5329 ;
  assign n6190 = ~x425 & n5191 ;
  assign n6191 = x457 & ~n5155 ;
  assign n6192 = x489 & n5155 ;
  assign n6193 = ~n6191 & ~n6192 ;
  assign n6194 = ~n5191 & n6193 ;
  assign n6195 = ~n6190 & ~n6194 ;
  assign n6196 = ~n5237 & n6195 ;
  assign n6197 = x393 & n5237 ;
  assign n6198 = ~n6196 & ~n6197 ;
  assign n6199 = ~n5283 & ~n6198 ;
  assign n6200 = x361 & n5283 ;
  assign n6201 = ~n6199 & ~n6200 ;
  assign n6202 = ~n5329 & n6201 ;
  assign n6203 = ~n6189 & ~n6202 ;
  assign n6204 = ~n5375 & ~n6203 ;
  assign n6205 = ~x297 & n5375 ;
  assign n6206 = ~n6204 & ~n6205 ;
  assign n6207 = ~n5421 & ~n6206 ;
  assign n6208 = ~x265 & n5421 ;
  assign n6209 = ~n6207 & ~n6208 ;
  assign n6210 = ~n5467 & n6209 ;
  assign n6211 = x233 & n5467 ;
  assign n6212 = ~n6210 & ~n6211 ;
  assign n6213 = ~n5513 & n6212 ;
  assign n6214 = ~n6188 & ~n6213 ;
  assign n6215 = ~n5559 & ~n6214 ;
  assign n6216 = ~x169 & n5559 ;
  assign n6217 = ~n6215 & ~n6216 ;
  assign n6218 = ~n5605 & n6217 ;
  assign n6219 = x137 & n5605 ;
  assign n6220 = ~n6218 & ~n6219 ;
  assign n6221 = ~n5648 & ~n6220 ;
  assign n6222 = x105 & n5648 ;
  assign n6223 = ~n6221 & ~n6222 ;
  assign n6224 = ~n5691 & ~n6223 ;
  assign n6225 = x73 & n5691 ;
  assign n6226 = ~n6224 & ~n6225 ;
  assign n6227 = ~n5737 & n6226 ;
  assign n6228 = ~n6187 & ~n6227 ;
  assign n6229 = n5780 & ~n6228 ;
  assign n6230 = ~n6186 & ~n6229 ;
  assign n6231 = ~x10 & ~n5780 ;
  assign n6232 = ~x42 & n5737 ;
  assign n6233 = ~x202 & n5513 ;
  assign n6234 = ~x330 & n5329 ;
  assign n6235 = ~x426 & n5191 ;
  assign n6236 = x458 & ~n5155 ;
  assign n6237 = x490 & n5155 ;
  assign n6238 = ~n6236 & ~n6237 ;
  assign n6239 = ~n5191 & n6238 ;
  assign n6240 = ~n6235 & ~n6239 ;
  assign n6241 = ~n5237 & n6240 ;
  assign n6242 = x394 & n5237 ;
  assign n6243 = ~n6241 & ~n6242 ;
  assign n6244 = ~n5283 & ~n6243 ;
  assign n6245 = x362 & n5283 ;
  assign n6246 = ~n6244 & ~n6245 ;
  assign n6247 = ~n5329 & n6246 ;
  assign n6248 = ~n6234 & ~n6247 ;
  assign n6249 = ~n5375 & ~n6248 ;
  assign n6250 = ~x298 & n5375 ;
  assign n6251 = ~n6249 & ~n6250 ;
  assign n6252 = ~n5421 & ~n6251 ;
  assign n6253 = ~x266 & n5421 ;
  assign n6254 = ~n6252 & ~n6253 ;
  assign n6255 = ~n5467 & n6254 ;
  assign n6256 = x234 & n5467 ;
  assign n6257 = ~n6255 & ~n6256 ;
  assign n6258 = ~n5513 & n6257 ;
  assign n6259 = ~n6233 & ~n6258 ;
  assign n6260 = ~n5559 & ~n6259 ;
  assign n6261 = ~x170 & n5559 ;
  assign n6262 = ~n6260 & ~n6261 ;
  assign n6263 = ~n5605 & n6262 ;
  assign n6264 = x138 & n5605 ;
  assign n6265 = ~n6263 & ~n6264 ;
  assign n6266 = ~n5648 & ~n6265 ;
  assign n6267 = x106 & n5648 ;
  assign n6268 = ~n6266 & ~n6267 ;
  assign n6269 = ~n5691 & ~n6268 ;
  assign n6270 = x74 & n5691 ;
  assign n6271 = ~n6269 & ~n6270 ;
  assign n6272 = ~n5737 & n6271 ;
  assign n6273 = ~n6232 & ~n6272 ;
  assign n6274 = n5780 & ~n6273 ;
  assign n6275 = ~n6231 & ~n6274 ;
  assign n6276 = ~x11 & ~n5780 ;
  assign n6277 = ~x43 & n5737 ;
  assign n6278 = ~x203 & n5513 ;
  assign n6279 = ~x331 & n5329 ;
  assign n6280 = ~x427 & n5191 ;
  assign n6281 = x459 & ~n5155 ;
  assign n6282 = x491 & n5155 ;
  assign n6283 = ~n6281 & ~n6282 ;
  assign n6284 = ~n5191 & n6283 ;
  assign n6285 = ~n6280 & ~n6284 ;
  assign n6286 = ~n5237 & n6285 ;
  assign n6287 = x395 & n5237 ;
  assign n6288 = ~n6286 & ~n6287 ;
  assign n6289 = ~n5283 & ~n6288 ;
  assign n6290 = x363 & n5283 ;
  assign n6291 = ~n6289 & ~n6290 ;
  assign n6292 = ~n5329 & n6291 ;
  assign n6293 = ~n6279 & ~n6292 ;
  assign n6294 = ~n5375 & ~n6293 ;
  assign n6295 = ~x299 & n5375 ;
  assign n6296 = ~n6294 & ~n6295 ;
  assign n6297 = ~n5421 & ~n6296 ;
  assign n6298 = ~x267 & n5421 ;
  assign n6299 = ~n6297 & ~n6298 ;
  assign n6300 = ~n5467 & n6299 ;
  assign n6301 = x235 & n5467 ;
  assign n6302 = ~n6300 & ~n6301 ;
  assign n6303 = ~n5513 & n6302 ;
  assign n6304 = ~n6278 & ~n6303 ;
  assign n6305 = ~n5559 & ~n6304 ;
  assign n6306 = ~x171 & n5559 ;
  assign n6307 = ~n6305 & ~n6306 ;
  assign n6308 = ~n5605 & n6307 ;
  assign n6309 = x139 & n5605 ;
  assign n6310 = ~n6308 & ~n6309 ;
  assign n6311 = ~n5648 & ~n6310 ;
  assign n6312 = x107 & n5648 ;
  assign n6313 = ~n6311 & ~n6312 ;
  assign n6314 = ~n5691 & ~n6313 ;
  assign n6315 = x75 & n5691 ;
  assign n6316 = ~n6314 & ~n6315 ;
  assign n6317 = ~n5737 & n6316 ;
  assign n6318 = ~n6277 & ~n6317 ;
  assign n6319 = n5780 & ~n6318 ;
  assign n6320 = ~n6276 & ~n6319 ;
  assign n6321 = ~x12 & ~n5780 ;
  assign n6322 = ~x44 & n5737 ;
  assign n6323 = ~x204 & n5513 ;
  assign n6324 = ~x332 & n5329 ;
  assign n6325 = ~x428 & n5191 ;
  assign n6326 = x460 & ~n5155 ;
  assign n6327 = x492 & n5155 ;
  assign n6328 = ~n6326 & ~n6327 ;
  assign n6329 = ~n5191 & n6328 ;
  assign n6330 = ~n6325 & ~n6329 ;
  assign n6331 = ~n5237 & n6330 ;
  assign n6332 = x396 & n5237 ;
  assign n6333 = ~n6331 & ~n6332 ;
  assign n6334 = ~n5283 & ~n6333 ;
  assign n6335 = x364 & n5283 ;
  assign n6336 = ~n6334 & ~n6335 ;
  assign n6337 = ~n5329 & n6336 ;
  assign n6338 = ~n6324 & ~n6337 ;
  assign n6339 = ~n5375 & ~n6338 ;
  assign n6340 = ~x300 & n5375 ;
  assign n6341 = ~n6339 & ~n6340 ;
  assign n6342 = ~n5421 & ~n6341 ;
  assign n6343 = ~x268 & n5421 ;
  assign n6344 = ~n6342 & ~n6343 ;
  assign n6345 = ~n5467 & n6344 ;
  assign n6346 = x236 & n5467 ;
  assign n6347 = ~n6345 & ~n6346 ;
  assign n6348 = ~n5513 & n6347 ;
  assign n6349 = ~n6323 & ~n6348 ;
  assign n6350 = ~n5559 & ~n6349 ;
  assign n6351 = ~x172 & n5559 ;
  assign n6352 = ~n6350 & ~n6351 ;
  assign n6353 = ~n5605 & n6352 ;
  assign n6354 = x140 & n5605 ;
  assign n6355 = ~n6353 & ~n6354 ;
  assign n6356 = ~n5648 & ~n6355 ;
  assign n6357 = x108 & n5648 ;
  assign n6358 = ~n6356 & ~n6357 ;
  assign n6359 = ~n5691 & ~n6358 ;
  assign n6360 = x76 & n5691 ;
  assign n6361 = ~n6359 & ~n6360 ;
  assign n6362 = ~n5737 & n6361 ;
  assign n6363 = ~n6322 & ~n6362 ;
  assign n6364 = n5780 & ~n6363 ;
  assign n6365 = ~n6321 & ~n6364 ;
  assign n6366 = ~x13 & ~n5780 ;
  assign n6367 = ~x45 & n5737 ;
  assign n6368 = ~x205 & n5513 ;
  assign n6369 = ~x333 & n5329 ;
  assign n6370 = ~x429 & n5191 ;
  assign n6371 = x461 & ~n5155 ;
  assign n6372 = x493 & n5155 ;
  assign n6373 = ~n6371 & ~n6372 ;
  assign n6374 = ~n5191 & n6373 ;
  assign n6375 = ~n6370 & ~n6374 ;
  assign n6376 = ~n5237 & n6375 ;
  assign n6377 = x397 & n5237 ;
  assign n6378 = ~n6376 & ~n6377 ;
  assign n6379 = ~n5283 & ~n6378 ;
  assign n6380 = x365 & n5283 ;
  assign n6381 = ~n6379 & ~n6380 ;
  assign n6382 = ~n5329 & n6381 ;
  assign n6383 = ~n6369 & ~n6382 ;
  assign n6384 = ~n5375 & ~n6383 ;
  assign n6385 = ~x301 & n5375 ;
  assign n6386 = ~n6384 & ~n6385 ;
  assign n6387 = ~n5421 & ~n6386 ;
  assign n6388 = ~x269 & n5421 ;
  assign n6389 = ~n6387 & ~n6388 ;
  assign n6390 = ~n5467 & n6389 ;
  assign n6391 = x237 & n5467 ;
  assign n6392 = ~n6390 & ~n6391 ;
  assign n6393 = ~n5513 & n6392 ;
  assign n6394 = ~n6368 & ~n6393 ;
  assign n6395 = ~n5559 & ~n6394 ;
  assign n6396 = ~x173 & n5559 ;
  assign n6397 = ~n6395 & ~n6396 ;
  assign n6398 = ~n5605 & n6397 ;
  assign n6399 = x141 & n5605 ;
  assign n6400 = ~n6398 & ~n6399 ;
  assign n6401 = ~n5648 & ~n6400 ;
  assign n6402 = x109 & n5648 ;
  assign n6403 = ~n6401 & ~n6402 ;
  assign n6404 = ~n5691 & ~n6403 ;
  assign n6405 = x77 & n5691 ;
  assign n6406 = ~n6404 & ~n6405 ;
  assign n6407 = ~n5737 & n6406 ;
  assign n6408 = ~n6367 & ~n6407 ;
  assign n6409 = n5780 & ~n6408 ;
  assign n6410 = ~n6366 & ~n6409 ;
  assign n6411 = ~x14 & ~n5780 ;
  assign n6412 = ~x46 & n5737 ;
  assign n6413 = ~x206 & n5513 ;
  assign n6414 = ~x334 & n5329 ;
  assign n6415 = ~x430 & n5191 ;
  assign n6416 = x462 & ~n5155 ;
  assign n6417 = x494 & n5155 ;
  assign n6418 = ~n6416 & ~n6417 ;
  assign n6419 = ~n5191 & n6418 ;
  assign n6420 = ~n6415 & ~n6419 ;
  assign n6421 = ~n5237 & n6420 ;
  assign n6422 = x398 & n5237 ;
  assign n6423 = ~n6421 & ~n6422 ;
  assign n6424 = ~n5283 & ~n6423 ;
  assign n6425 = x366 & n5283 ;
  assign n6426 = ~n6424 & ~n6425 ;
  assign n6427 = ~n5329 & n6426 ;
  assign n6428 = ~n6414 & ~n6427 ;
  assign n6429 = ~n5375 & ~n6428 ;
  assign n6430 = ~x302 & n5375 ;
  assign n6431 = ~n6429 & ~n6430 ;
  assign n6432 = ~n5421 & ~n6431 ;
  assign n6433 = ~x270 & n5421 ;
  assign n6434 = ~n6432 & ~n6433 ;
  assign n6435 = ~n5467 & n6434 ;
  assign n6436 = x238 & n5467 ;
  assign n6437 = ~n6435 & ~n6436 ;
  assign n6438 = ~n5513 & n6437 ;
  assign n6439 = ~n6413 & ~n6438 ;
  assign n6440 = ~n5559 & ~n6439 ;
  assign n6441 = ~x174 & n5559 ;
  assign n6442 = ~n6440 & ~n6441 ;
  assign n6443 = ~n5605 & n6442 ;
  assign n6444 = x142 & n5605 ;
  assign n6445 = ~n6443 & ~n6444 ;
  assign n6446 = ~n5648 & ~n6445 ;
  assign n6447 = x110 & n5648 ;
  assign n6448 = ~n6446 & ~n6447 ;
  assign n6449 = ~n5691 & ~n6448 ;
  assign n6450 = x78 & n5691 ;
  assign n6451 = ~n6449 & ~n6450 ;
  assign n6452 = ~n5737 & n6451 ;
  assign n6453 = ~n6412 & ~n6452 ;
  assign n6454 = n5780 & ~n6453 ;
  assign n6455 = ~n6411 & ~n6454 ;
  assign n6456 = ~x15 & ~n5780 ;
  assign n6457 = ~x47 & n5737 ;
  assign n6458 = ~x207 & n5513 ;
  assign n6459 = ~x335 & n5329 ;
  assign n6460 = ~x431 & n5191 ;
  assign n6461 = x463 & ~n5155 ;
  assign n6462 = x495 & n5155 ;
  assign n6463 = ~n6461 & ~n6462 ;
  assign n6464 = ~n5191 & n6463 ;
  assign n6465 = ~n6460 & ~n6464 ;
  assign n6466 = ~n5237 & n6465 ;
  assign n6467 = x399 & n5237 ;
  assign n6468 = ~n6466 & ~n6467 ;
  assign n6469 = ~n5283 & ~n6468 ;
  assign n6470 = x367 & n5283 ;
  assign n6471 = ~n6469 & ~n6470 ;
  assign n6472 = ~n5329 & n6471 ;
  assign n6473 = ~n6459 & ~n6472 ;
  assign n6474 = ~n5375 & ~n6473 ;
  assign n6475 = ~x303 & n5375 ;
  assign n6476 = ~n6474 & ~n6475 ;
  assign n6477 = ~n5421 & ~n6476 ;
  assign n6478 = ~x271 & n5421 ;
  assign n6479 = ~n6477 & ~n6478 ;
  assign n6480 = ~n5467 & n6479 ;
  assign n6481 = x239 & n5467 ;
  assign n6482 = ~n6480 & ~n6481 ;
  assign n6483 = ~n5513 & n6482 ;
  assign n6484 = ~n6458 & ~n6483 ;
  assign n6485 = ~n5559 & ~n6484 ;
  assign n6486 = ~x175 & n5559 ;
  assign n6487 = ~n6485 & ~n6486 ;
  assign n6488 = ~n5605 & n6487 ;
  assign n6489 = x143 & n5605 ;
  assign n6490 = ~n6488 & ~n6489 ;
  assign n6491 = ~n5648 & ~n6490 ;
  assign n6492 = x111 & n5648 ;
  assign n6493 = ~n6491 & ~n6492 ;
  assign n6494 = ~n5691 & ~n6493 ;
  assign n6495 = x79 & n5691 ;
  assign n6496 = ~n6494 & ~n6495 ;
  assign n6497 = ~n5737 & n6496 ;
  assign n6498 = ~n6457 & ~n6497 ;
  assign n6499 = n5780 & ~n6498 ;
  assign n6500 = ~n6456 & ~n6499 ;
  assign n6501 = ~x16 & ~n5780 ;
  assign n6502 = ~x48 & n5737 ;
  assign n6503 = ~x208 & n5513 ;
  assign n6504 = ~x336 & n5329 ;
  assign n6505 = ~x432 & n5191 ;
  assign n6506 = x464 & ~n5155 ;
  assign n6507 = x496 & n5155 ;
  assign n6508 = ~n6506 & ~n6507 ;
  assign n6509 = ~n5191 & n6508 ;
  assign n6510 = ~n6505 & ~n6509 ;
  assign n6511 = ~n5237 & n6510 ;
  assign n6512 = x400 & n5237 ;
  assign n6513 = ~n6511 & ~n6512 ;
  assign n6514 = ~n5283 & ~n6513 ;
  assign n6515 = x368 & n5283 ;
  assign n6516 = ~n6514 & ~n6515 ;
  assign n6517 = ~n5329 & n6516 ;
  assign n6518 = ~n6504 & ~n6517 ;
  assign n6519 = ~n5375 & ~n6518 ;
  assign n6520 = ~x304 & n5375 ;
  assign n6521 = ~n6519 & ~n6520 ;
  assign n6522 = ~n5421 & ~n6521 ;
  assign n6523 = ~x272 & n5421 ;
  assign n6524 = ~n6522 & ~n6523 ;
  assign n6525 = ~n5467 & n6524 ;
  assign n6526 = x240 & n5467 ;
  assign n6527 = ~n6525 & ~n6526 ;
  assign n6528 = ~n5513 & n6527 ;
  assign n6529 = ~n6503 & ~n6528 ;
  assign n6530 = ~n5559 & ~n6529 ;
  assign n6531 = ~x176 & n5559 ;
  assign n6532 = ~n6530 & ~n6531 ;
  assign n6533 = ~n5605 & n6532 ;
  assign n6534 = x144 & n5605 ;
  assign n6535 = ~n6533 & ~n6534 ;
  assign n6536 = ~n5648 & ~n6535 ;
  assign n6537 = x112 & n5648 ;
  assign n6538 = ~n6536 & ~n6537 ;
  assign n6539 = ~n5691 & ~n6538 ;
  assign n6540 = x80 & n5691 ;
  assign n6541 = ~n6539 & ~n6540 ;
  assign n6542 = ~n5737 & n6541 ;
  assign n6543 = ~n6502 & ~n6542 ;
  assign n6544 = n5780 & ~n6543 ;
  assign n6545 = ~n6501 & ~n6544 ;
  assign n6546 = ~x17 & ~n5780 ;
  assign n6547 = ~x49 & n5737 ;
  assign n6548 = ~x209 & n5513 ;
  assign n6549 = ~x337 & n5329 ;
  assign n6550 = ~x433 & n5191 ;
  assign n6551 = x465 & ~n5155 ;
  assign n6552 = x497 & n5155 ;
  assign n6553 = ~n6551 & ~n6552 ;
  assign n6554 = ~n5191 & n6553 ;
  assign n6555 = ~n6550 & ~n6554 ;
  assign n6556 = ~n5237 & n6555 ;
  assign n6557 = x401 & n5237 ;
  assign n6558 = ~n6556 & ~n6557 ;
  assign n6559 = ~n5283 & ~n6558 ;
  assign n6560 = x369 & n5283 ;
  assign n6561 = ~n6559 & ~n6560 ;
  assign n6562 = ~n5329 & n6561 ;
  assign n6563 = ~n6549 & ~n6562 ;
  assign n6564 = ~n5375 & ~n6563 ;
  assign n6565 = ~x305 & n5375 ;
  assign n6566 = ~n6564 & ~n6565 ;
  assign n6567 = ~n5421 & ~n6566 ;
  assign n6568 = ~x273 & n5421 ;
  assign n6569 = ~n6567 & ~n6568 ;
  assign n6570 = ~n5467 & n6569 ;
  assign n6571 = x241 & n5467 ;
  assign n6572 = ~n6570 & ~n6571 ;
  assign n6573 = ~n5513 & n6572 ;
  assign n6574 = ~n6548 & ~n6573 ;
  assign n6575 = ~n5559 & ~n6574 ;
  assign n6576 = ~x177 & n5559 ;
  assign n6577 = ~n6575 & ~n6576 ;
  assign n6578 = ~n5605 & n6577 ;
  assign n6579 = x145 & n5605 ;
  assign n6580 = ~n6578 & ~n6579 ;
  assign n6581 = ~n5648 & ~n6580 ;
  assign n6582 = x113 & n5648 ;
  assign n6583 = ~n6581 & ~n6582 ;
  assign n6584 = ~n5691 & ~n6583 ;
  assign n6585 = x81 & n5691 ;
  assign n6586 = ~n6584 & ~n6585 ;
  assign n6587 = ~n5737 & n6586 ;
  assign n6588 = ~n6547 & ~n6587 ;
  assign n6589 = n5780 & ~n6588 ;
  assign n6590 = ~n6546 & ~n6589 ;
  assign n6591 = ~x18 & ~n5780 ;
  assign n6592 = ~x50 & n5737 ;
  assign n6593 = ~x210 & n5513 ;
  assign n6594 = ~x338 & n5329 ;
  assign n6595 = ~x434 & n5191 ;
  assign n6596 = x466 & ~n5155 ;
  assign n6597 = x498 & n5155 ;
  assign n6598 = ~n6596 & ~n6597 ;
  assign n6599 = ~n5191 & n6598 ;
  assign n6600 = ~n6595 & ~n6599 ;
  assign n6601 = ~n5237 & n6600 ;
  assign n6602 = x402 & n5237 ;
  assign n6603 = ~n6601 & ~n6602 ;
  assign n6604 = ~n5283 & ~n6603 ;
  assign n6605 = x370 & n5283 ;
  assign n6606 = ~n6604 & ~n6605 ;
  assign n6607 = ~n5329 & n6606 ;
  assign n6608 = ~n6594 & ~n6607 ;
  assign n6609 = ~n5375 & ~n6608 ;
  assign n6610 = ~x306 & n5375 ;
  assign n6611 = ~n6609 & ~n6610 ;
  assign n6612 = ~n5421 & ~n6611 ;
  assign n6613 = ~x274 & n5421 ;
  assign n6614 = ~n6612 & ~n6613 ;
  assign n6615 = ~n5467 & n6614 ;
  assign n6616 = x242 & n5467 ;
  assign n6617 = ~n6615 & ~n6616 ;
  assign n6618 = ~n5513 & n6617 ;
  assign n6619 = ~n6593 & ~n6618 ;
  assign n6620 = ~n5559 & ~n6619 ;
  assign n6621 = ~x178 & n5559 ;
  assign n6622 = ~n6620 & ~n6621 ;
  assign n6623 = ~n5605 & n6622 ;
  assign n6624 = x146 & n5605 ;
  assign n6625 = ~n6623 & ~n6624 ;
  assign n6626 = ~n5648 & ~n6625 ;
  assign n6627 = x114 & n5648 ;
  assign n6628 = ~n6626 & ~n6627 ;
  assign n6629 = ~n5691 & ~n6628 ;
  assign n6630 = x82 & n5691 ;
  assign n6631 = ~n6629 & ~n6630 ;
  assign n6632 = ~n5737 & n6631 ;
  assign n6633 = ~n6592 & ~n6632 ;
  assign n6634 = n5780 & ~n6633 ;
  assign n6635 = ~n6591 & ~n6634 ;
  assign n6636 = ~x19 & ~n5780 ;
  assign n6637 = ~x51 & n5737 ;
  assign n6638 = ~x211 & n5513 ;
  assign n6639 = ~x339 & n5329 ;
  assign n6640 = ~x435 & n5191 ;
  assign n6641 = x467 & ~n5155 ;
  assign n6642 = x499 & n5155 ;
  assign n6643 = ~n6641 & ~n6642 ;
  assign n6644 = ~n5191 & n6643 ;
  assign n6645 = ~n6640 & ~n6644 ;
  assign n6646 = ~n5237 & n6645 ;
  assign n6647 = x403 & n5237 ;
  assign n6648 = ~n6646 & ~n6647 ;
  assign n6649 = ~n5283 & ~n6648 ;
  assign n6650 = x371 & n5283 ;
  assign n6651 = ~n6649 & ~n6650 ;
  assign n6652 = ~n5329 & n6651 ;
  assign n6653 = ~n6639 & ~n6652 ;
  assign n6654 = ~n5375 & ~n6653 ;
  assign n6655 = ~x307 & n5375 ;
  assign n6656 = ~n6654 & ~n6655 ;
  assign n6657 = ~n5421 & ~n6656 ;
  assign n6658 = ~x275 & n5421 ;
  assign n6659 = ~n6657 & ~n6658 ;
  assign n6660 = ~n5467 & n6659 ;
  assign n6661 = x243 & n5467 ;
  assign n6662 = ~n6660 & ~n6661 ;
  assign n6663 = ~n5513 & n6662 ;
  assign n6664 = ~n6638 & ~n6663 ;
  assign n6665 = ~n5559 & ~n6664 ;
  assign n6666 = ~x179 & n5559 ;
  assign n6667 = ~n6665 & ~n6666 ;
  assign n6668 = ~n5605 & n6667 ;
  assign n6669 = x147 & n5605 ;
  assign n6670 = ~n6668 & ~n6669 ;
  assign n6671 = ~n5648 & ~n6670 ;
  assign n6672 = x115 & n5648 ;
  assign n6673 = ~n6671 & ~n6672 ;
  assign n6674 = ~n5691 & ~n6673 ;
  assign n6675 = x83 & n5691 ;
  assign n6676 = ~n6674 & ~n6675 ;
  assign n6677 = ~n5737 & n6676 ;
  assign n6678 = ~n6637 & ~n6677 ;
  assign n6679 = n5780 & ~n6678 ;
  assign n6680 = ~n6636 & ~n6679 ;
  assign n6681 = ~x20 & ~n5780 ;
  assign n6682 = ~x52 & n5737 ;
  assign n6683 = ~x212 & n5513 ;
  assign n6684 = ~x340 & n5329 ;
  assign n6685 = ~x436 & n5191 ;
  assign n6686 = x468 & ~n5155 ;
  assign n6687 = x500 & n5155 ;
  assign n6688 = ~n6686 & ~n6687 ;
  assign n6689 = ~n5191 & n6688 ;
  assign n6690 = ~n6685 & ~n6689 ;
  assign n6691 = ~n5237 & n6690 ;
  assign n6692 = x404 & n5237 ;
  assign n6693 = ~n6691 & ~n6692 ;
  assign n6694 = ~n5283 & ~n6693 ;
  assign n6695 = x372 & n5283 ;
  assign n6696 = ~n6694 & ~n6695 ;
  assign n6697 = ~n5329 & n6696 ;
  assign n6698 = ~n6684 & ~n6697 ;
  assign n6699 = ~n5375 & ~n6698 ;
  assign n6700 = ~x308 & n5375 ;
  assign n6701 = ~n6699 & ~n6700 ;
  assign n6702 = ~n5421 & ~n6701 ;
  assign n6703 = ~x276 & n5421 ;
  assign n6704 = ~n6702 & ~n6703 ;
  assign n6705 = ~n5467 & n6704 ;
  assign n6706 = x244 & n5467 ;
  assign n6707 = ~n6705 & ~n6706 ;
  assign n6708 = ~n5513 & n6707 ;
  assign n6709 = ~n6683 & ~n6708 ;
  assign n6710 = ~n5559 & ~n6709 ;
  assign n6711 = ~x180 & n5559 ;
  assign n6712 = ~n6710 & ~n6711 ;
  assign n6713 = ~n5605 & n6712 ;
  assign n6714 = x148 & n5605 ;
  assign n6715 = ~n6713 & ~n6714 ;
  assign n6716 = ~n5648 & ~n6715 ;
  assign n6717 = x116 & n5648 ;
  assign n6718 = ~n6716 & ~n6717 ;
  assign n6719 = ~n5691 & ~n6718 ;
  assign n6720 = x84 & n5691 ;
  assign n6721 = ~n6719 & ~n6720 ;
  assign n6722 = ~n5737 & n6721 ;
  assign n6723 = ~n6682 & ~n6722 ;
  assign n6724 = n5780 & ~n6723 ;
  assign n6725 = ~n6681 & ~n6724 ;
  assign n6726 = ~x21 & ~n5780 ;
  assign n6727 = ~x53 & n5737 ;
  assign n6728 = ~x213 & n5513 ;
  assign n6729 = ~x341 & n5329 ;
  assign n6730 = ~x437 & n5191 ;
  assign n6731 = x469 & ~n5155 ;
  assign n6732 = x501 & n5155 ;
  assign n6733 = ~n6731 & ~n6732 ;
  assign n6734 = ~n5191 & n6733 ;
  assign n6735 = ~n6730 & ~n6734 ;
  assign n6736 = ~n5237 & n6735 ;
  assign n6737 = x405 & n5237 ;
  assign n6738 = ~n6736 & ~n6737 ;
  assign n6739 = ~n5283 & ~n6738 ;
  assign n6740 = x373 & n5283 ;
  assign n6741 = ~n6739 & ~n6740 ;
  assign n6742 = ~n5329 & n6741 ;
  assign n6743 = ~n6729 & ~n6742 ;
  assign n6744 = ~n5375 & ~n6743 ;
  assign n6745 = ~x309 & n5375 ;
  assign n6746 = ~n6744 & ~n6745 ;
  assign n6747 = ~n5421 & ~n6746 ;
  assign n6748 = ~x277 & n5421 ;
  assign n6749 = ~n6747 & ~n6748 ;
  assign n6750 = ~n5467 & n6749 ;
  assign n6751 = x245 & n5467 ;
  assign n6752 = ~n6750 & ~n6751 ;
  assign n6753 = ~n5513 & n6752 ;
  assign n6754 = ~n6728 & ~n6753 ;
  assign n6755 = ~n5559 & ~n6754 ;
  assign n6756 = ~x181 & n5559 ;
  assign n6757 = ~n6755 & ~n6756 ;
  assign n6758 = ~n5605 & n6757 ;
  assign n6759 = x149 & n5605 ;
  assign n6760 = ~n6758 & ~n6759 ;
  assign n6761 = ~n5648 & ~n6760 ;
  assign n6762 = x117 & n5648 ;
  assign n6763 = ~n6761 & ~n6762 ;
  assign n6764 = ~n5691 & ~n6763 ;
  assign n6765 = x85 & n5691 ;
  assign n6766 = ~n6764 & ~n6765 ;
  assign n6767 = ~n5737 & n6766 ;
  assign n6768 = ~n6727 & ~n6767 ;
  assign n6769 = n5780 & ~n6768 ;
  assign n6770 = ~n6726 & ~n6769 ;
  assign n6771 = ~x22 & ~n5780 ;
  assign n6772 = ~x54 & n5737 ;
  assign n6773 = ~x214 & n5513 ;
  assign n6774 = ~x342 & n5329 ;
  assign n6775 = ~x438 & n5191 ;
  assign n6776 = x470 & ~n5155 ;
  assign n6777 = x502 & n5155 ;
  assign n6778 = ~n6776 & ~n6777 ;
  assign n6779 = ~n5191 & n6778 ;
  assign n6780 = ~n6775 & ~n6779 ;
  assign n6781 = ~n5237 & n6780 ;
  assign n6782 = x406 & n5237 ;
  assign n6783 = ~n6781 & ~n6782 ;
  assign n6784 = ~n5283 & ~n6783 ;
  assign n6785 = x374 & n5283 ;
  assign n6786 = ~n6784 & ~n6785 ;
  assign n6787 = ~n5329 & n6786 ;
  assign n6788 = ~n6774 & ~n6787 ;
  assign n6789 = ~n5375 & ~n6788 ;
  assign n6790 = ~x310 & n5375 ;
  assign n6791 = ~n6789 & ~n6790 ;
  assign n6792 = ~n5421 & ~n6791 ;
  assign n6793 = ~x278 & n5421 ;
  assign n6794 = ~n6792 & ~n6793 ;
  assign n6795 = ~n5467 & n6794 ;
  assign n6796 = x246 & n5467 ;
  assign n6797 = ~n6795 & ~n6796 ;
  assign n6798 = ~n5513 & n6797 ;
  assign n6799 = ~n6773 & ~n6798 ;
  assign n6800 = ~n5559 & ~n6799 ;
  assign n6801 = ~x182 & n5559 ;
  assign n6802 = ~n6800 & ~n6801 ;
  assign n6803 = ~n5605 & n6802 ;
  assign n6804 = x150 & n5605 ;
  assign n6805 = ~n6803 & ~n6804 ;
  assign n6806 = ~n5648 & ~n6805 ;
  assign n6807 = x118 & n5648 ;
  assign n6808 = ~n6806 & ~n6807 ;
  assign n6809 = ~n5691 & ~n6808 ;
  assign n6810 = x86 & n5691 ;
  assign n6811 = ~n6809 & ~n6810 ;
  assign n6812 = ~n5737 & n6811 ;
  assign n6813 = ~n6772 & ~n6812 ;
  assign n6814 = n5780 & ~n6813 ;
  assign n6815 = ~n6771 & ~n6814 ;
  assign n6816 = ~x23 & ~n5780 ;
  assign n6817 = ~x55 & n5737 ;
  assign n6818 = ~x215 & n5513 ;
  assign n6819 = ~x343 & n5329 ;
  assign n6820 = ~x439 & n5191 ;
  assign n6821 = x471 & ~n5155 ;
  assign n6822 = x503 & n5155 ;
  assign n6823 = ~n6821 & ~n6822 ;
  assign n6824 = ~n5191 & n6823 ;
  assign n6825 = ~n6820 & ~n6824 ;
  assign n6826 = ~n5237 & n6825 ;
  assign n6827 = x407 & n5237 ;
  assign n6828 = ~n6826 & ~n6827 ;
  assign n6829 = ~n5283 & ~n6828 ;
  assign n6830 = x375 & n5283 ;
  assign n6831 = ~n6829 & ~n6830 ;
  assign n6832 = ~n5329 & n6831 ;
  assign n6833 = ~n6819 & ~n6832 ;
  assign n6834 = ~n5375 & ~n6833 ;
  assign n6835 = ~x311 & n5375 ;
  assign n6836 = ~n6834 & ~n6835 ;
  assign n6837 = ~n5421 & ~n6836 ;
  assign n6838 = ~x279 & n5421 ;
  assign n6839 = ~n6837 & ~n6838 ;
  assign n6840 = ~n5467 & n6839 ;
  assign n6841 = x247 & n5467 ;
  assign n6842 = ~n6840 & ~n6841 ;
  assign n6843 = ~n5513 & n6842 ;
  assign n6844 = ~n6818 & ~n6843 ;
  assign n6845 = ~n5559 & ~n6844 ;
  assign n6846 = ~x183 & n5559 ;
  assign n6847 = ~n6845 & ~n6846 ;
  assign n6848 = ~n5605 & n6847 ;
  assign n6849 = x151 & n5605 ;
  assign n6850 = ~n6848 & ~n6849 ;
  assign n6851 = ~n5648 & ~n6850 ;
  assign n6852 = x119 & n5648 ;
  assign n6853 = ~n6851 & ~n6852 ;
  assign n6854 = ~n5691 & ~n6853 ;
  assign n6855 = x87 & n5691 ;
  assign n6856 = ~n6854 & ~n6855 ;
  assign n6857 = ~n5737 & n6856 ;
  assign n6858 = ~n6817 & ~n6857 ;
  assign n6859 = n5780 & ~n6858 ;
  assign n6860 = ~n6816 & ~n6859 ;
  assign n6861 = ~x24 & ~n5780 ;
  assign n6862 = ~x56 & n5737 ;
  assign n6863 = ~x216 & n5513 ;
  assign n6864 = ~x344 & n5329 ;
  assign n6865 = ~x440 & n5191 ;
  assign n6866 = x472 & ~n5155 ;
  assign n6867 = x504 & n5155 ;
  assign n6868 = ~n6866 & ~n6867 ;
  assign n6869 = ~n5191 & n6868 ;
  assign n6870 = ~n6865 & ~n6869 ;
  assign n6871 = ~n5237 & n6870 ;
  assign n6872 = x408 & n5237 ;
  assign n6873 = ~n6871 & ~n6872 ;
  assign n6874 = ~n5283 & ~n6873 ;
  assign n6875 = x376 & n5283 ;
  assign n6876 = ~n6874 & ~n6875 ;
  assign n6877 = ~n5329 & n6876 ;
  assign n6878 = ~n6864 & ~n6877 ;
  assign n6879 = ~n5375 & ~n6878 ;
  assign n6880 = ~x312 & n5375 ;
  assign n6881 = ~n6879 & ~n6880 ;
  assign n6882 = ~n5421 & ~n6881 ;
  assign n6883 = ~x280 & n5421 ;
  assign n6884 = ~n6882 & ~n6883 ;
  assign n6885 = ~n5467 & n6884 ;
  assign n6886 = x248 & n5467 ;
  assign n6887 = ~n6885 & ~n6886 ;
  assign n6888 = ~n5513 & n6887 ;
  assign n6889 = ~n6863 & ~n6888 ;
  assign n6890 = ~n5559 & ~n6889 ;
  assign n6891 = ~x184 & n5559 ;
  assign n6892 = ~n6890 & ~n6891 ;
  assign n6893 = ~n5605 & n6892 ;
  assign n6894 = x152 & n5605 ;
  assign n6895 = ~n6893 & ~n6894 ;
  assign n6896 = ~n5648 & ~n6895 ;
  assign n6897 = x120 & n5648 ;
  assign n6898 = ~n6896 & ~n6897 ;
  assign n6899 = ~n5691 & ~n6898 ;
  assign n6900 = x88 & n5691 ;
  assign n6901 = ~n6899 & ~n6900 ;
  assign n6902 = ~n5737 & n6901 ;
  assign n6903 = ~n6862 & ~n6902 ;
  assign n6904 = n5780 & ~n6903 ;
  assign n6905 = ~n6861 & ~n6904 ;
  assign n6906 = ~x25 & ~n5780 ;
  assign n6907 = ~x57 & n5737 ;
  assign n6908 = ~x217 & n5513 ;
  assign n6909 = ~x345 & n5329 ;
  assign n6910 = ~x441 & n5191 ;
  assign n6911 = x473 & ~n5155 ;
  assign n6912 = x505 & n5155 ;
  assign n6913 = ~n6911 & ~n6912 ;
  assign n6914 = ~n5191 & n6913 ;
  assign n6915 = ~n6910 & ~n6914 ;
  assign n6916 = ~n5237 & n6915 ;
  assign n6917 = x409 & n5237 ;
  assign n6918 = ~n6916 & ~n6917 ;
  assign n6919 = ~n5283 & ~n6918 ;
  assign n6920 = x377 & n5283 ;
  assign n6921 = ~n6919 & ~n6920 ;
  assign n6922 = ~n5329 & n6921 ;
  assign n6923 = ~n6909 & ~n6922 ;
  assign n6924 = ~n5375 & ~n6923 ;
  assign n6925 = ~x313 & n5375 ;
  assign n6926 = ~n6924 & ~n6925 ;
  assign n6927 = ~n5421 & ~n6926 ;
  assign n6928 = ~x281 & n5421 ;
  assign n6929 = ~n6927 & ~n6928 ;
  assign n6930 = ~n5467 & n6929 ;
  assign n6931 = x249 & n5467 ;
  assign n6932 = ~n6930 & ~n6931 ;
  assign n6933 = ~n5513 & n6932 ;
  assign n6934 = ~n6908 & ~n6933 ;
  assign n6935 = ~n5559 & ~n6934 ;
  assign n6936 = ~x185 & n5559 ;
  assign n6937 = ~n6935 & ~n6936 ;
  assign n6938 = ~n5605 & n6937 ;
  assign n6939 = x153 & n5605 ;
  assign n6940 = ~n6938 & ~n6939 ;
  assign n6941 = ~n5648 & ~n6940 ;
  assign n6942 = x121 & n5648 ;
  assign n6943 = ~n6941 & ~n6942 ;
  assign n6944 = ~n5691 & ~n6943 ;
  assign n6945 = x89 & n5691 ;
  assign n6946 = ~n6944 & ~n6945 ;
  assign n6947 = ~n5737 & n6946 ;
  assign n6948 = ~n6907 & ~n6947 ;
  assign n6949 = n5780 & ~n6948 ;
  assign n6950 = ~n6906 & ~n6949 ;
  assign n6951 = ~x26 & ~n5780 ;
  assign n6952 = ~x58 & n5737 ;
  assign n6953 = ~x218 & n5513 ;
  assign n6954 = ~x346 & n5329 ;
  assign n6955 = ~x442 & n5191 ;
  assign n6956 = x474 & ~n5155 ;
  assign n6957 = x506 & n5155 ;
  assign n6958 = ~n6956 & ~n6957 ;
  assign n6959 = ~n5191 & n6958 ;
  assign n6960 = ~n6955 & ~n6959 ;
  assign n6961 = ~n5237 & n6960 ;
  assign n6962 = x410 & n5237 ;
  assign n6963 = ~n6961 & ~n6962 ;
  assign n6964 = ~n5283 & ~n6963 ;
  assign n6965 = x378 & n5283 ;
  assign n6966 = ~n6964 & ~n6965 ;
  assign n6967 = ~n5329 & n6966 ;
  assign n6968 = ~n6954 & ~n6967 ;
  assign n6969 = ~n5375 & ~n6968 ;
  assign n6970 = ~x314 & n5375 ;
  assign n6971 = ~n6969 & ~n6970 ;
  assign n6972 = ~n5421 & ~n6971 ;
  assign n6973 = ~x282 & n5421 ;
  assign n6974 = ~n6972 & ~n6973 ;
  assign n6975 = ~n5467 & n6974 ;
  assign n6976 = x250 & n5467 ;
  assign n6977 = ~n6975 & ~n6976 ;
  assign n6978 = ~n5513 & n6977 ;
  assign n6979 = ~n6953 & ~n6978 ;
  assign n6980 = ~n5559 & ~n6979 ;
  assign n6981 = ~x186 & n5559 ;
  assign n6982 = ~n6980 & ~n6981 ;
  assign n6983 = ~n5605 & n6982 ;
  assign n6984 = x154 & n5605 ;
  assign n6985 = ~n6983 & ~n6984 ;
  assign n6986 = ~n5648 & ~n6985 ;
  assign n6987 = x122 & n5648 ;
  assign n6988 = ~n6986 & ~n6987 ;
  assign n6989 = ~n5691 & ~n6988 ;
  assign n6990 = x90 & n5691 ;
  assign n6991 = ~n6989 & ~n6990 ;
  assign n6992 = ~n5737 & n6991 ;
  assign n6993 = ~n6952 & ~n6992 ;
  assign n6994 = n5780 & ~n6993 ;
  assign n6995 = ~n6951 & ~n6994 ;
  assign n6996 = ~x27 & ~n5780 ;
  assign n6997 = ~x59 & n5737 ;
  assign n6998 = ~x219 & n5513 ;
  assign n6999 = ~x347 & n5329 ;
  assign n7000 = ~x443 & n5191 ;
  assign n7001 = x475 & ~n5155 ;
  assign n7002 = x507 & n5155 ;
  assign n7003 = ~n7001 & ~n7002 ;
  assign n7004 = ~n5191 & n7003 ;
  assign n7005 = ~n7000 & ~n7004 ;
  assign n7006 = ~n5237 & n7005 ;
  assign n7007 = x411 & n5237 ;
  assign n7008 = ~n7006 & ~n7007 ;
  assign n7009 = ~n5283 & ~n7008 ;
  assign n7010 = x379 & n5283 ;
  assign n7011 = ~n7009 & ~n7010 ;
  assign n7012 = ~n5329 & n7011 ;
  assign n7013 = ~n6999 & ~n7012 ;
  assign n7014 = ~n5375 & ~n7013 ;
  assign n7015 = ~x315 & n5375 ;
  assign n7016 = ~n7014 & ~n7015 ;
  assign n7017 = ~n5421 & ~n7016 ;
  assign n7018 = ~x283 & n5421 ;
  assign n7019 = ~n7017 & ~n7018 ;
  assign n7020 = ~n5467 & n7019 ;
  assign n7021 = x251 & n5467 ;
  assign n7022 = ~n7020 & ~n7021 ;
  assign n7023 = ~n5513 & n7022 ;
  assign n7024 = ~n6998 & ~n7023 ;
  assign n7025 = ~n5559 & ~n7024 ;
  assign n7026 = ~x187 & n5559 ;
  assign n7027 = ~n7025 & ~n7026 ;
  assign n7028 = ~n5605 & n7027 ;
  assign n7029 = x155 & n5605 ;
  assign n7030 = ~n7028 & ~n7029 ;
  assign n7031 = ~n5648 & ~n7030 ;
  assign n7032 = x123 & n5648 ;
  assign n7033 = ~n7031 & ~n7032 ;
  assign n7034 = ~n5691 & ~n7033 ;
  assign n7035 = x91 & n5691 ;
  assign n7036 = ~n7034 & ~n7035 ;
  assign n7037 = ~n5737 & n7036 ;
  assign n7038 = ~n6997 & ~n7037 ;
  assign n7039 = n5780 & ~n7038 ;
  assign n7040 = ~n6996 & ~n7039 ;
  assign n7041 = ~x28 & ~n5780 ;
  assign n7042 = ~x60 & n5737 ;
  assign n7043 = ~x220 & n5513 ;
  assign n7044 = ~x348 & n5329 ;
  assign n7045 = ~x444 & n5191 ;
  assign n7046 = x476 & ~n5155 ;
  assign n7047 = x508 & n5155 ;
  assign n7048 = ~n7046 & ~n7047 ;
  assign n7049 = ~n5191 & n7048 ;
  assign n7050 = ~n7045 & ~n7049 ;
  assign n7051 = ~n5237 & n7050 ;
  assign n7052 = x412 & n5237 ;
  assign n7053 = ~n7051 & ~n7052 ;
  assign n7054 = ~n5283 & ~n7053 ;
  assign n7055 = x380 & n5283 ;
  assign n7056 = ~n7054 & ~n7055 ;
  assign n7057 = ~n5329 & n7056 ;
  assign n7058 = ~n7044 & ~n7057 ;
  assign n7059 = ~n5375 & ~n7058 ;
  assign n7060 = ~x316 & n5375 ;
  assign n7061 = ~n7059 & ~n7060 ;
  assign n7062 = ~n5421 & ~n7061 ;
  assign n7063 = ~x284 & n5421 ;
  assign n7064 = ~n7062 & ~n7063 ;
  assign n7065 = ~n5467 & n7064 ;
  assign n7066 = x252 & n5467 ;
  assign n7067 = ~n7065 & ~n7066 ;
  assign n7068 = ~n5513 & n7067 ;
  assign n7069 = ~n7043 & ~n7068 ;
  assign n7070 = ~n5559 & ~n7069 ;
  assign n7071 = ~x188 & n5559 ;
  assign n7072 = ~n7070 & ~n7071 ;
  assign n7073 = ~n5605 & n7072 ;
  assign n7074 = x156 & n5605 ;
  assign n7075 = ~n7073 & ~n7074 ;
  assign n7076 = ~n5648 & ~n7075 ;
  assign n7077 = x124 & n5648 ;
  assign n7078 = ~n7076 & ~n7077 ;
  assign n7079 = ~n5691 & ~n7078 ;
  assign n7080 = x92 & n5691 ;
  assign n7081 = ~n7079 & ~n7080 ;
  assign n7082 = ~n5737 & n7081 ;
  assign n7083 = ~n7042 & ~n7082 ;
  assign n7084 = n5780 & ~n7083 ;
  assign n7085 = ~n7041 & ~n7084 ;
  assign n7086 = ~x29 & ~n5780 ;
  assign n7087 = ~x61 & n5737 ;
  assign n7088 = ~x221 & n5513 ;
  assign n7089 = ~x349 & n5329 ;
  assign n7090 = ~x445 & n5191 ;
  assign n7091 = x477 & ~n5155 ;
  assign n7092 = x509 & n5155 ;
  assign n7093 = ~n7091 & ~n7092 ;
  assign n7094 = ~n5191 & n7093 ;
  assign n7095 = ~n7090 & ~n7094 ;
  assign n7096 = ~n5237 & n7095 ;
  assign n7097 = x413 & n5237 ;
  assign n7098 = ~n7096 & ~n7097 ;
  assign n7099 = ~n5283 & ~n7098 ;
  assign n7100 = x381 & n5283 ;
  assign n7101 = ~n7099 & ~n7100 ;
  assign n7102 = ~n5329 & n7101 ;
  assign n7103 = ~n7089 & ~n7102 ;
  assign n7104 = ~n5375 & ~n7103 ;
  assign n7105 = ~x317 & n5375 ;
  assign n7106 = ~n7104 & ~n7105 ;
  assign n7107 = ~n5421 & ~n7106 ;
  assign n7108 = ~x285 & n5421 ;
  assign n7109 = ~n7107 & ~n7108 ;
  assign n7110 = ~n5467 & n7109 ;
  assign n7111 = x253 & n5467 ;
  assign n7112 = ~n7110 & ~n7111 ;
  assign n7113 = ~n5513 & n7112 ;
  assign n7114 = ~n7088 & ~n7113 ;
  assign n7115 = ~n5559 & ~n7114 ;
  assign n7116 = ~x189 & n5559 ;
  assign n7117 = ~n7115 & ~n7116 ;
  assign n7118 = ~n5605 & n7117 ;
  assign n7119 = x157 & n5605 ;
  assign n7120 = ~n7118 & ~n7119 ;
  assign n7121 = ~n5648 & ~n7120 ;
  assign n7122 = x125 & n5648 ;
  assign n7123 = ~n7121 & ~n7122 ;
  assign n7124 = ~n5691 & ~n7123 ;
  assign n7125 = x93 & n5691 ;
  assign n7126 = ~n7124 & ~n7125 ;
  assign n7127 = ~n5737 & n7126 ;
  assign n7128 = ~n7087 & ~n7127 ;
  assign n7129 = n5780 & ~n7128 ;
  assign n7130 = ~n7086 & ~n7129 ;
  assign n7131 = ~x30 & ~n5780 ;
  assign n7132 = ~x62 & n5737 ;
  assign n7133 = ~x222 & n5513 ;
  assign n7134 = ~x350 & n5329 ;
  assign n7135 = ~x446 & n5191 ;
  assign n7136 = x478 & ~n5155 ;
  assign n7137 = x510 & n5155 ;
  assign n7138 = ~n7136 & ~n7137 ;
  assign n7139 = ~n5191 & n7138 ;
  assign n7140 = ~n7135 & ~n7139 ;
  assign n7141 = ~n5237 & n7140 ;
  assign n7142 = x414 & n5237 ;
  assign n7143 = ~n7141 & ~n7142 ;
  assign n7144 = ~n5283 & ~n7143 ;
  assign n7145 = x382 & n5283 ;
  assign n7146 = ~n7144 & ~n7145 ;
  assign n7147 = ~n5329 & n7146 ;
  assign n7148 = ~n7134 & ~n7147 ;
  assign n7149 = ~n5375 & ~n7148 ;
  assign n7150 = ~x318 & n5375 ;
  assign n7151 = ~n7149 & ~n7150 ;
  assign n7152 = ~n5421 & ~n7151 ;
  assign n7153 = ~x286 & n5421 ;
  assign n7154 = ~n7152 & ~n7153 ;
  assign n7155 = ~n5467 & n7154 ;
  assign n7156 = x254 & n5467 ;
  assign n7157 = ~n7155 & ~n7156 ;
  assign n7158 = ~n5513 & n7157 ;
  assign n7159 = ~n7133 & ~n7158 ;
  assign n7160 = ~n5559 & ~n7159 ;
  assign n7161 = ~x190 & n5559 ;
  assign n7162 = ~n7160 & ~n7161 ;
  assign n7163 = ~n5605 & n7162 ;
  assign n7164 = x158 & n5605 ;
  assign n7165 = ~n7163 & ~n7164 ;
  assign n7166 = ~n5648 & ~n7165 ;
  assign n7167 = x126 & n5648 ;
  assign n7168 = ~n7166 & ~n7167 ;
  assign n7169 = ~n5691 & ~n7168 ;
  assign n7170 = x94 & n5691 ;
  assign n7171 = ~n7169 & ~n7170 ;
  assign n7172 = ~n5737 & n7171 ;
  assign n7173 = ~n7132 & ~n7172 ;
  assign n7174 = n5780 & ~n7173 ;
  assign n7175 = ~n7131 & ~n7174 ;
  assign n7176 = ~x31 & ~n5780 ;
  assign n7177 = ~x63 & n5737 ;
  assign n7178 = ~x223 & n5513 ;
  assign n7179 = ~x351 & n5329 ;
  assign n7180 = ~x447 & n5191 ;
  assign n7181 = x479 & ~n5155 ;
  assign n7182 = x511 & n5155 ;
  assign n7183 = ~n7181 & ~n7182 ;
  assign n7184 = ~n5191 & n7183 ;
  assign n7185 = ~n7180 & ~n7184 ;
  assign n7186 = ~n5237 & n7185 ;
  assign n7187 = x415 & n5237 ;
  assign n7188 = ~n7186 & ~n7187 ;
  assign n7189 = ~n5283 & ~n7188 ;
  assign n7190 = x383 & n5283 ;
  assign n7191 = ~n7189 & ~n7190 ;
  assign n7192 = ~n5329 & n7191 ;
  assign n7193 = ~n7179 & ~n7192 ;
  assign n7194 = ~n5375 & ~n7193 ;
  assign n7195 = ~x319 & n5375 ;
  assign n7196 = ~n7194 & ~n7195 ;
  assign n7197 = ~n5421 & ~n7196 ;
  assign n7198 = ~x287 & n5421 ;
  assign n7199 = ~n7197 & ~n7198 ;
  assign n7200 = ~n5467 & n7199 ;
  assign n7201 = x255 & n5467 ;
  assign n7202 = ~n7200 & ~n7201 ;
  assign n7203 = ~n5513 & n7202 ;
  assign n7204 = ~n7178 & ~n7203 ;
  assign n7205 = ~n5559 & ~n7204 ;
  assign n7206 = ~x191 & n5559 ;
  assign n7207 = ~n7205 & ~n7206 ;
  assign n7208 = ~n5605 & n7207 ;
  assign n7209 = x159 & n5605 ;
  assign n7210 = ~n7208 & ~n7209 ;
  assign n7211 = ~n5648 & ~n7210 ;
  assign n7212 = x127 & n5648 ;
  assign n7213 = ~n7211 & ~n7212 ;
  assign n7214 = ~n5691 & ~n7213 ;
  assign n7215 = x95 & n5691 ;
  assign n7216 = ~n7214 & ~n7215 ;
  assign n7217 = ~n5737 & n7216 ;
  assign n7218 = ~n7177 & ~n7217 ;
  assign n7219 = n5780 & ~n7218 ;
  assign n7220 = ~n7176 & ~n7219 ;
  assign y0 = n5825 ;
  assign y1 = n5870 ;
  assign y2 = n5915 ;
  assign y3 = n5960 ;
  assign y4 = n6005 ;
  assign y5 = n6050 ;
  assign y6 = n6095 ;
  assign y7 = n6140 ;
  assign y8 = n6185 ;
  assign y9 = n6230 ;
  assign y10 = n6275 ;
  assign y11 = n6320 ;
  assign y12 = n6365 ;
  assign y13 = n6410 ;
  assign y14 = n6455 ;
  assign y15 = n6500 ;
  assign y16 = n6545 ;
  assign y17 = n6590 ;
  assign y18 = n6635 ;
  assign y19 = n6680 ;
  assign y20 = n6725 ;
  assign y21 = n6770 ;
  assign y22 = n6815 ;
  assign y23 = n6860 ;
  assign y24 = n6905 ;
  assign y25 = n6950 ;
  assign y26 = n6995 ;
  assign y27 = n7040 ;
  assign y28 = n7085 ;
  assign y29 = n7130 ;
  assign y30 = n7175 ;
  assign y31 = n7220 ;
endmodule
