module and_ary_16( a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, b11, b12, b13, b14, b15, d0 );
  input a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15;
  input b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, b11, b12, b13, b14, b15;
  output d0;
  wire c0, c1, c2, c3, c4, c5, c6, c7, c8, c9, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c20, c21, c22, c23, c24, c25, c26, c27, c28, c29;
  assign c0 = a0 & b0 ;
  assign c1 = a1 & b1 ;
  assign c2 = a2 & b2 ;
  assign c3 = a3 & b3 ;
  assign c4 = a4 & b4 ;
  assign c5 = a5 & b5 ;
  assign c6 = a6 & b6 ;
  assign c7 = a7 & b7 ;
  assign c8 = a8 & b8 ;
  assign c9 = a9 & b9 ;
  assign c10 = a10 & b10 ;
  assign c11 = a11 & b11 ;
  assign c12 = a12 & b12 ;
  assign c13 = a13 & b13 ;
  assign c14 = a14 & b14 ;
  assign c15 = a15 & b15 ;
  assign c16 = c0 & c1 ;
  assign c17 = c2 & c3 ;
  assign c18 = c4 & c5 ;
  assign c19 = c6 & c7 ;
  assign c20 = c8 & c9 ;
  assign c21 = c10 & c11 ;
  assign c22 = c12 & c13 ;
  assign c23 = c14 & c15 ;
  assign c24 = c16 & c17 ;
  assign c25 = c18 & c19 ;
  assign c26 = c20 & c21 ;
  assign c27 = c22 & c23 ;
  assign c28 = c24 & c25 ;
  assign c29 = c26 & c27 ;
  assign d0 = c28 & c29 ;
endmodule
