module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 ;
  assign n159 = x0 & ~x40 ;
  assign n126 = x40 ^ x0 ;
  assign n157 = x1 & ~x41 ;
  assign n158 = ~n126 & n157 ;
  assign n160 = n159 ^ n158 ;
  assign n127 = x41 ^ x1 ;
  assign n128 = ~n126 & ~n127 ;
  assign n154 = x2 & ~x42 ;
  assign n129 = x42 ^ x2 ;
  assign n152 = x3 & ~x43 ;
  assign n153 = ~n129 & n152 ;
  assign n155 = n154 ^ n153 ;
  assign n156 = n128 & n155 ;
  assign n161 = n160 ^ n156 ;
  assign n130 = x43 ^ x3 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = n128 & n131 ;
  assign n148 = x4 & ~x44 ;
  assign n133 = x44 ^ x4 ;
  assign n146 = x5 & ~x45 ;
  assign n147 = ~n133 & n146 ;
  assign n149 = n148 ^ n147 ;
  assign n134 = x45 ^ x5 ;
  assign n135 = ~n133 & ~n134 ;
  assign n143 = x6 & ~x46 ;
  assign n136 = x46 ^ x6 ;
  assign n141 = x7 & ~x47 ;
  assign n142 = ~n136 & n141 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = n135 & n144 ;
  assign n150 = n149 ^ n145 ;
  assign n151 = n132 & n150 ;
  assign n162 = n161 ^ n151 ;
  assign n137 = x47 ^ x7 ;
  assign n138 = ~n136 & ~n137 ;
  assign n139 = n135 & n138 ;
  assign n140 = n132 & n139 ;
  assign n163 = n162 ^ n140 ;
  assign n546 = x0 & ~x24 ;
  assign n513 = x24 ^ x0 ;
  assign n544 = x1 & ~x25 ;
  assign n545 = ~n513 & n544 ;
  assign n547 = n546 ^ n545 ;
  assign n514 = x25 ^ x1 ;
  assign n515 = ~n513 & ~n514 ;
  assign n541 = x2 & ~x26 ;
  assign n516 = x26 ^ x2 ;
  assign n539 = x3 & ~x27 ;
  assign n540 = ~n516 & n539 ;
  assign n542 = n541 ^ n540 ;
  assign n543 = n515 & n542 ;
  assign n548 = n547 ^ n543 ;
  assign n517 = x27 ^ x3 ;
  assign n518 = ~n516 & ~n517 ;
  assign n519 = n515 & n518 ;
  assign n535 = x4 & ~x28 ;
  assign n520 = x28 ^ x4 ;
  assign n533 = x5 & ~x29 ;
  assign n534 = ~n520 & n533 ;
  assign n536 = n535 ^ n534 ;
  assign n521 = x29 ^ x5 ;
  assign n522 = ~n520 & ~n521 ;
  assign n530 = x6 & ~x30 ;
  assign n523 = x30 ^ x6 ;
  assign n528 = x7 & ~x31 ;
  assign n529 = ~n523 & n528 ;
  assign n531 = n530 ^ n529 ;
  assign n532 = n522 & n531 ;
  assign n537 = n536 ^ n532 ;
  assign n538 = n519 & n537 ;
  assign n549 = n548 ^ n538 ;
  assign n524 = x31 ^ x7 ;
  assign n525 = ~n523 & ~n524 ;
  assign n526 = n522 & n525 ;
  assign n527 = n519 & n526 ;
  assign n550 = n549 ^ n527 ;
  assign n742 = ~n163 & n550 ;
  assign n371 = x0 & ~x32 ;
  assign n338 = x32 ^ x0 ;
  assign n369 = x1 & ~x33 ;
  assign n370 = ~n338 & n369 ;
  assign n372 = n371 ^ n370 ;
  assign n339 = x33 ^ x1 ;
  assign n340 = ~n338 & ~n339 ;
  assign n366 = x2 & ~x34 ;
  assign n341 = x34 ^ x2 ;
  assign n364 = x3 & ~x35 ;
  assign n365 = ~n341 & n364 ;
  assign n367 = n366 ^ n365 ;
  assign n368 = n340 & n367 ;
  assign n373 = n372 ^ n368 ;
  assign n342 = x35 ^ x3 ;
  assign n343 = ~n341 & ~n342 ;
  assign n344 = n340 & n343 ;
  assign n360 = x4 & ~x36 ;
  assign n345 = x36 ^ x4 ;
  assign n358 = x5 & ~x37 ;
  assign n359 = ~n345 & n358 ;
  assign n361 = n360 ^ n359 ;
  assign n346 = x37 ^ x5 ;
  assign n347 = ~n345 & ~n346 ;
  assign n355 = x6 & ~x38 ;
  assign n348 = x38 ^ x6 ;
  assign n353 = x7 & ~x39 ;
  assign n354 = ~n348 & n353 ;
  assign n356 = n355 ^ n354 ;
  assign n357 = n347 & n356 ;
  assign n362 = n361 ^ n357 ;
  assign n363 = n344 & n362 ;
  assign n374 = n373 ^ n363 ;
  assign n349 = x39 ^ x7 ;
  assign n350 = ~n348 & ~n349 ;
  assign n351 = n347 & n350 ;
  assign n352 = n344 & n351 ;
  assign n375 = n374 ^ n352 ;
  assign n741 = ~n375 & n550 ;
  assign n743 = n742 ^ n741 ;
  assign n731 = n375 ^ n163 ;
  assign n736 = n550 & n731 ;
  assign n744 = n743 ^ n736 ;
  assign n702 = x0 & ~x8 ;
  assign n669 = x8 ^ x0 ;
  assign n700 = x1 & ~x9 ;
  assign n701 = ~n669 & n700 ;
  assign n703 = n702 ^ n701 ;
  assign n670 = x9 ^ x1 ;
  assign n671 = ~n669 & ~n670 ;
  assign n697 = x2 & ~x10 ;
  assign n672 = x10 ^ x2 ;
  assign n695 = x3 & ~x11 ;
  assign n696 = ~n672 & n695 ;
  assign n698 = n697 ^ n696 ;
  assign n699 = n671 & n698 ;
  assign n704 = n703 ^ n699 ;
  assign n673 = x11 ^ x3 ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = n671 & n674 ;
  assign n691 = x4 & ~x12 ;
  assign n676 = x12 ^ x4 ;
  assign n689 = x5 & ~x13 ;
  assign n690 = ~n676 & n689 ;
  assign n692 = n691 ^ n690 ;
  assign n677 = x13 ^ x5 ;
  assign n678 = ~n676 & ~n677 ;
  assign n686 = x6 & ~x14 ;
  assign n679 = x14 ^ x6 ;
  assign n684 = x7 & ~x15 ;
  assign n685 = ~n679 & n684 ;
  assign n687 = n686 ^ n685 ;
  assign n688 = n678 & n687 ;
  assign n693 = n692 ^ n688 ;
  assign n694 = n675 & n693 ;
  assign n705 = n704 ^ n694 ;
  assign n680 = x15 ^ x7 ;
  assign n681 = ~n679 & ~n680 ;
  assign n682 = n678 & n681 ;
  assign n683 = n675 & n682 ;
  assign n706 = n705 ^ n683 ;
  assign n604 = x0 & ~x16 ;
  assign n571 = x16 ^ x0 ;
  assign n602 = x1 & ~x17 ;
  assign n603 = ~n571 & n602 ;
  assign n605 = n604 ^ n603 ;
  assign n572 = x17 ^ x1 ;
  assign n573 = ~n571 & ~n572 ;
  assign n599 = x2 & ~x18 ;
  assign n574 = x18 ^ x2 ;
  assign n597 = x3 & ~x19 ;
  assign n598 = ~n574 & n597 ;
  assign n600 = n599 ^ n598 ;
  assign n601 = n573 & n600 ;
  assign n606 = n605 ^ n601 ;
  assign n575 = x19 ^ x3 ;
  assign n576 = ~n574 & ~n575 ;
  assign n577 = n573 & n576 ;
  assign n593 = x4 & ~x20 ;
  assign n578 = x20 ^ x4 ;
  assign n591 = x5 & ~x21 ;
  assign n592 = ~n578 & n591 ;
  assign n594 = n593 ^ n592 ;
  assign n579 = x21 ^ x5 ;
  assign n580 = ~n578 & ~n579 ;
  assign n588 = x6 & ~x22 ;
  assign n581 = x22 ^ x6 ;
  assign n586 = x7 & ~x23 ;
  assign n587 = ~n581 & n586 ;
  assign n589 = n588 ^ n587 ;
  assign n590 = n580 & n589 ;
  assign n595 = n594 ^ n590 ;
  assign n596 = n577 & n595 ;
  assign n607 = n606 ^ n596 ;
  assign n582 = x23 ^ x7 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = n580 & n583 ;
  assign n585 = n577 & n584 ;
  assign n608 = n607 ^ n585 ;
  assign n730 = n706 ^ n608 ;
  assign n732 = n731 ^ n550 ;
  assign n733 = n730 & n732 ;
  assign n729 = n608 & n706 ;
  assign n734 = n733 ^ n729 ;
  assign n735 = n163 & n375 ;
  assign n737 = n736 ^ n735 ;
  assign n738 = n737 ^ n733 ;
  assign n739 = n734 & n738 ;
  assign n740 = n739 ^ n733 ;
  assign n745 = n744 ^ n740 ;
  assign n746 = n737 ^ n734 ;
  assign n747 = n732 ^ n730 ;
  assign n748 = x0 & ~n747 ;
  assign n749 = ~n746 & n748 ;
  assign n750 = ~n745 & n749 ;
  assign n120 = x8 & ~x40 ;
  assign n87 = x40 ^ x8 ;
  assign n118 = x9 & ~x41 ;
  assign n119 = ~n87 & n118 ;
  assign n121 = n120 ^ n119 ;
  assign n88 = x41 ^ x9 ;
  assign n89 = ~n87 & ~n88 ;
  assign n115 = x10 & ~x42 ;
  assign n90 = x42 ^ x10 ;
  assign n113 = x11 & ~x43 ;
  assign n114 = ~n90 & n113 ;
  assign n116 = n115 ^ n114 ;
  assign n117 = n89 & n116 ;
  assign n122 = n121 ^ n117 ;
  assign n91 = x43 ^ x11 ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = n89 & n92 ;
  assign n109 = x12 & ~x44 ;
  assign n94 = x44 ^ x12 ;
  assign n107 = x13 & ~x45 ;
  assign n108 = ~n94 & n107 ;
  assign n110 = n109 ^ n108 ;
  assign n95 = x45 ^ x13 ;
  assign n96 = ~n94 & ~n95 ;
  assign n104 = x14 & ~x46 ;
  assign n97 = x46 ^ x14 ;
  assign n102 = x15 & ~x47 ;
  assign n103 = ~n97 & n102 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n96 & n105 ;
  assign n111 = n110 ^ n106 ;
  assign n112 = n93 & n111 ;
  assign n123 = n122 ^ n112 ;
  assign n98 = x47 ^ x15 ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = n96 & n99 ;
  assign n101 = n93 & n100 ;
  assign n124 = n123 ^ n101 ;
  assign n507 = x8 & ~x24 ;
  assign n474 = x24 ^ x8 ;
  assign n505 = x9 & ~x25 ;
  assign n506 = ~n474 & n505 ;
  assign n508 = n507 ^ n506 ;
  assign n475 = x25 ^ x9 ;
  assign n476 = ~n474 & ~n475 ;
  assign n502 = x10 & ~x26 ;
  assign n477 = x26 ^ x10 ;
  assign n500 = x11 & ~x27 ;
  assign n501 = ~n477 & n500 ;
  assign n503 = n502 ^ n501 ;
  assign n504 = n476 & n503 ;
  assign n509 = n508 ^ n504 ;
  assign n478 = x27 ^ x11 ;
  assign n479 = ~n477 & ~n478 ;
  assign n480 = n476 & n479 ;
  assign n496 = x12 & ~x28 ;
  assign n481 = x28 ^ x12 ;
  assign n494 = x13 & ~x29 ;
  assign n495 = ~n481 & n494 ;
  assign n497 = n496 ^ n495 ;
  assign n482 = x29 ^ x13 ;
  assign n483 = ~n481 & ~n482 ;
  assign n491 = x14 & ~x30 ;
  assign n484 = x30 ^ x14 ;
  assign n489 = x15 & ~x31 ;
  assign n490 = ~n484 & n489 ;
  assign n492 = n491 ^ n490 ;
  assign n493 = n483 & n492 ;
  assign n498 = n497 ^ n493 ;
  assign n499 = n480 & n498 ;
  assign n510 = n509 ^ n499 ;
  assign n485 = x31 ^ x15 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = n483 & n486 ;
  assign n488 = n480 & n487 ;
  assign n511 = n510 ^ n488 ;
  assign n720 = ~n124 & n511 ;
  assign n332 = x8 & ~x32 ;
  assign n299 = x32 ^ x8 ;
  assign n330 = x9 & ~x33 ;
  assign n331 = ~n299 & n330 ;
  assign n333 = n332 ^ n331 ;
  assign n300 = x33 ^ x9 ;
  assign n301 = ~n299 & ~n300 ;
  assign n327 = x10 & ~x34 ;
  assign n302 = x34 ^ x10 ;
  assign n325 = x11 & ~x35 ;
  assign n326 = ~n302 & n325 ;
  assign n328 = n327 ^ n326 ;
  assign n329 = n301 & n328 ;
  assign n334 = n333 ^ n329 ;
  assign n303 = x35 ^ x11 ;
  assign n304 = ~n302 & ~n303 ;
  assign n305 = n301 & n304 ;
  assign n321 = x12 & ~x36 ;
  assign n306 = x36 ^ x12 ;
  assign n319 = x13 & ~x37 ;
  assign n320 = ~n306 & n319 ;
  assign n322 = n321 ^ n320 ;
  assign n307 = x37 ^ x13 ;
  assign n308 = ~n306 & ~n307 ;
  assign n316 = x14 & ~x38 ;
  assign n309 = x38 ^ x14 ;
  assign n314 = x15 & ~x39 ;
  assign n315 = ~n309 & n314 ;
  assign n317 = n316 ^ n315 ;
  assign n318 = n308 & n317 ;
  assign n323 = n322 ^ n318 ;
  assign n324 = n305 & n323 ;
  assign n335 = n334 ^ n324 ;
  assign n310 = x39 ^ x15 ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = n308 & n311 ;
  assign n313 = n305 & n312 ;
  assign n336 = n335 ^ n313 ;
  assign n719 = ~n336 & n511 ;
  assign n721 = n720 ^ n719 ;
  assign n709 = n336 ^ n124 ;
  assign n714 = n511 & n709 ;
  assign n722 = n721 ^ n714 ;
  assign n642 = x8 & ~x16 ;
  assign n609 = x16 ^ x8 ;
  assign n640 = x9 & ~x17 ;
  assign n641 = ~n609 & n640 ;
  assign n643 = n642 ^ n641 ;
  assign n610 = x17 ^ x9 ;
  assign n611 = ~n609 & ~n610 ;
  assign n637 = x10 & ~x18 ;
  assign n612 = x18 ^ x10 ;
  assign n635 = x11 & ~x19 ;
  assign n636 = ~n612 & n635 ;
  assign n638 = n637 ^ n636 ;
  assign n639 = n611 & n638 ;
  assign n644 = n643 ^ n639 ;
  assign n613 = x19 ^ x11 ;
  assign n614 = ~n612 & ~n613 ;
  assign n615 = n611 & n614 ;
  assign n631 = x12 & ~x20 ;
  assign n616 = x20 ^ x12 ;
  assign n629 = x13 & ~x21 ;
  assign n630 = ~n616 & n629 ;
  assign n632 = n631 ^ n630 ;
  assign n617 = x21 ^ x13 ;
  assign n618 = ~n616 & ~n617 ;
  assign n626 = x14 & ~x22 ;
  assign n619 = x22 ^ x14 ;
  assign n624 = x15 & ~x23 ;
  assign n625 = ~n619 & n624 ;
  assign n627 = n626 ^ n625 ;
  assign n628 = n618 & n627 ;
  assign n633 = n632 ^ n628 ;
  assign n634 = n615 & n633 ;
  assign n645 = n644 ^ n634 ;
  assign n620 = x23 ^ x15 ;
  assign n621 = ~n619 & ~n620 ;
  assign n622 = n618 & n621 ;
  assign n623 = n615 & n622 ;
  assign n646 = n645 ^ n623 ;
  assign n708 = n706 ^ n646 ;
  assign n710 = n709 ^ n511 ;
  assign n711 = ~n708 & n710 ;
  assign n707 = n646 & ~n706 ;
  assign n712 = n711 ^ n707 ;
  assign n713 = n124 & n336 ;
  assign n715 = n714 ^ n713 ;
  assign n716 = n715 ^ n711 ;
  assign n717 = n712 & n716 ;
  assign n718 = n717 ^ n711 ;
  assign n723 = n722 ^ n718 ;
  assign n724 = n715 ^ n712 ;
  assign n725 = n710 ^ n708 ;
  assign n726 = x8 & n725 ;
  assign n727 = ~n724 & n726 ;
  assign n728 = ~n723 & n727 ;
  assign n751 = n750 ^ n728 ;
  assign n82 = x16 & ~x40 ;
  assign n49 = x40 ^ x16 ;
  assign n80 = x17 & ~x41 ;
  assign n81 = ~n49 & n80 ;
  assign n83 = n82 ^ n81 ;
  assign n50 = x41 ^ x17 ;
  assign n51 = ~n49 & ~n50 ;
  assign n77 = x18 & ~x42 ;
  assign n52 = x42 ^ x18 ;
  assign n75 = x19 & ~x43 ;
  assign n76 = ~n52 & n75 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = n51 & n78 ;
  assign n84 = n83 ^ n79 ;
  assign n53 = x43 ^ x19 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n51 & n54 ;
  assign n71 = x20 & ~x44 ;
  assign n56 = x44 ^ x20 ;
  assign n69 = x21 & ~x45 ;
  assign n70 = ~n56 & n69 ;
  assign n72 = n71 ^ n70 ;
  assign n57 = x45 ^ x21 ;
  assign n58 = ~n56 & ~n57 ;
  assign n66 = x22 & ~x46 ;
  assign n59 = x46 ^ x22 ;
  assign n64 = x23 & ~x47 ;
  assign n65 = ~n59 & n64 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = n58 & n67 ;
  assign n73 = n72 ^ n68 ;
  assign n74 = n55 & n73 ;
  assign n85 = n84 ^ n74 ;
  assign n60 = x47 ^ x23 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = n58 & n61 ;
  assign n63 = n55 & n62 ;
  assign n86 = n85 ^ n63 ;
  assign n469 = x16 & ~x24 ;
  assign n436 = x24 ^ x16 ;
  assign n467 = x17 & ~x25 ;
  assign n468 = ~n436 & n467 ;
  assign n470 = n469 ^ n468 ;
  assign n437 = x25 ^ x17 ;
  assign n438 = ~n436 & ~n437 ;
  assign n464 = x18 & ~x26 ;
  assign n439 = x26 ^ x18 ;
  assign n462 = x19 & ~x27 ;
  assign n463 = ~n439 & n462 ;
  assign n465 = n464 ^ n463 ;
  assign n466 = n438 & n465 ;
  assign n471 = n470 ^ n466 ;
  assign n440 = x27 ^ x19 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = n438 & n441 ;
  assign n458 = x20 & ~x28 ;
  assign n443 = x28 ^ x20 ;
  assign n456 = x21 & ~x29 ;
  assign n457 = ~n443 & n456 ;
  assign n459 = n458 ^ n457 ;
  assign n444 = x29 ^ x21 ;
  assign n445 = ~n443 & ~n444 ;
  assign n453 = x22 & ~x30 ;
  assign n446 = x30 ^ x22 ;
  assign n451 = x23 & ~x31 ;
  assign n452 = ~n446 & n451 ;
  assign n454 = n453 ^ n452 ;
  assign n455 = n445 & n454 ;
  assign n460 = n459 ^ n455 ;
  assign n461 = n442 & n460 ;
  assign n472 = n471 ^ n461 ;
  assign n447 = x31 ^ x23 ;
  assign n448 = ~n446 & ~n447 ;
  assign n449 = n445 & n448 ;
  assign n450 = n442 & n449 ;
  assign n473 = n472 ^ n450 ;
  assign n660 = ~n86 & n473 ;
  assign n294 = x16 & ~x32 ;
  assign n261 = x32 ^ x16 ;
  assign n292 = x17 & ~x33 ;
  assign n293 = ~n261 & n292 ;
  assign n295 = n294 ^ n293 ;
  assign n262 = x33 ^ x17 ;
  assign n263 = ~n261 & ~n262 ;
  assign n289 = x18 & ~x34 ;
  assign n264 = x34 ^ x18 ;
  assign n287 = x19 & ~x35 ;
  assign n288 = ~n264 & n287 ;
  assign n290 = n289 ^ n288 ;
  assign n291 = n263 & n290 ;
  assign n296 = n295 ^ n291 ;
  assign n265 = x35 ^ x19 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = n263 & n266 ;
  assign n283 = x20 & ~x36 ;
  assign n268 = x36 ^ x20 ;
  assign n281 = x21 & ~x37 ;
  assign n282 = ~n268 & n281 ;
  assign n284 = n283 ^ n282 ;
  assign n269 = x37 ^ x21 ;
  assign n270 = ~n268 & ~n269 ;
  assign n278 = x22 & ~x38 ;
  assign n271 = x38 ^ x22 ;
  assign n276 = x23 & ~x39 ;
  assign n277 = ~n271 & n276 ;
  assign n279 = n278 ^ n277 ;
  assign n280 = n270 & n279 ;
  assign n285 = n284 ^ n280 ;
  assign n286 = n267 & n285 ;
  assign n297 = n296 ^ n286 ;
  assign n272 = x39 ^ x23 ;
  assign n273 = ~n271 & ~n272 ;
  assign n274 = n270 & n273 ;
  assign n275 = n267 & n274 ;
  assign n298 = n297 ^ n275 ;
  assign n659 = ~n298 & n473 ;
  assign n661 = n660 ^ n659 ;
  assign n649 = n298 ^ n86 ;
  assign n654 = n473 & n649 ;
  assign n662 = n661 ^ n654 ;
  assign n648 = n646 ^ n608 ;
  assign n650 = n649 ^ n473 ;
  assign n651 = n648 & n650 ;
  assign n647 = ~n608 & ~n646 ;
  assign n652 = n651 ^ n647 ;
  assign n653 = n86 & n298 ;
  assign n655 = n654 ^ n653 ;
  assign n656 = n655 ^ n651 ;
  assign n657 = n652 & n656 ;
  assign n658 = n657 ^ n651 ;
  assign n663 = n662 ^ n658 ;
  assign n664 = n655 ^ n652 ;
  assign n665 = n650 ^ n648 ;
  assign n666 = x16 & ~n665 ;
  assign n667 = ~n664 & n666 ;
  assign n668 = ~n663 & n667 ;
  assign n752 = n751 ^ n668 ;
  assign n562 = ~n473 & ~n550 ;
  assign n561 = ~n511 & ~n550 ;
  assign n563 = n562 ^ n561 ;
  assign n512 = n511 ^ n473 ;
  assign n554 = n512 & ~n550 ;
  assign n564 = n563 ^ n554 ;
  assign n553 = ~n473 & ~n511 ;
  assign n555 = n554 ^ n553 ;
  assign n410 = x24 & ~x32 ;
  assign n377 = x32 ^ x24 ;
  assign n408 = x25 & ~x33 ;
  assign n409 = ~n377 & n408 ;
  assign n411 = n410 ^ n409 ;
  assign n378 = x33 ^ x25 ;
  assign n379 = ~n377 & ~n378 ;
  assign n405 = x26 & ~x34 ;
  assign n380 = x34 ^ x26 ;
  assign n403 = x27 & ~x35 ;
  assign n404 = ~n380 & n403 ;
  assign n406 = n405 ^ n404 ;
  assign n407 = n379 & n406 ;
  assign n412 = n411 ^ n407 ;
  assign n381 = x35 ^ x27 ;
  assign n382 = ~n380 & ~n381 ;
  assign n383 = n379 & n382 ;
  assign n399 = x28 & ~x36 ;
  assign n384 = x36 ^ x28 ;
  assign n397 = x29 & ~x37 ;
  assign n398 = ~n384 & n397 ;
  assign n400 = n399 ^ n398 ;
  assign n385 = x37 ^ x29 ;
  assign n386 = ~n384 & ~n385 ;
  assign n394 = x30 & ~x38 ;
  assign n387 = x38 ^ x30 ;
  assign n392 = x31 & ~x39 ;
  assign n393 = ~n387 & n392 ;
  assign n395 = n394 ^ n393 ;
  assign n396 = n386 & n395 ;
  assign n401 = n400 ^ n396 ;
  assign n402 = n383 & n401 ;
  assign n413 = n412 ^ n402 ;
  assign n388 = x39 ^ x31 ;
  assign n389 = ~n387 & ~n388 ;
  assign n390 = n386 & n389 ;
  assign n391 = n383 & n390 ;
  assign n414 = n413 ^ n391 ;
  assign n236 = x24 & ~x40 ;
  assign n203 = x40 ^ x24 ;
  assign n234 = x25 & ~x41 ;
  assign n235 = ~n203 & n234 ;
  assign n237 = n236 ^ n235 ;
  assign n204 = x41 ^ x25 ;
  assign n205 = ~n203 & ~n204 ;
  assign n231 = x26 & ~x42 ;
  assign n206 = x42 ^ x26 ;
  assign n229 = x27 & ~x43 ;
  assign n230 = ~n206 & n229 ;
  assign n232 = n231 ^ n230 ;
  assign n233 = n205 & n232 ;
  assign n238 = n237 ^ n233 ;
  assign n207 = x43 ^ x27 ;
  assign n208 = ~n206 & ~n207 ;
  assign n209 = n205 & n208 ;
  assign n225 = x28 & ~x44 ;
  assign n210 = x44 ^ x28 ;
  assign n223 = x29 & ~x45 ;
  assign n224 = ~n210 & n223 ;
  assign n226 = n225 ^ n224 ;
  assign n211 = x45 ^ x29 ;
  assign n212 = ~n210 & ~n211 ;
  assign n220 = x30 & ~x46 ;
  assign n213 = x46 ^ x30 ;
  assign n218 = x31 & ~x47 ;
  assign n219 = ~n213 & n218 ;
  assign n221 = n220 ^ n219 ;
  assign n222 = n212 & n221 ;
  assign n227 = n226 ^ n222 ;
  assign n228 = n209 & n227 ;
  assign n239 = n238 ^ n228 ;
  assign n214 = x47 ^ x31 ;
  assign n215 = ~n213 & ~n214 ;
  assign n216 = n212 & n215 ;
  assign n217 = n209 & n216 ;
  assign n240 = n239 ^ n217 ;
  assign n435 = n414 ^ n240 ;
  assign n551 = n550 ^ n512 ;
  assign n552 = n435 & ~n551 ;
  assign n556 = n555 ^ n552 ;
  assign n557 = n240 & n414 ;
  assign n558 = n557 ^ n552 ;
  assign n559 = n556 & n558 ;
  assign n560 = n559 ^ n552 ;
  assign n565 = n564 ^ n560 ;
  assign n566 = n557 ^ n556 ;
  assign n567 = n551 ^ n435 ;
  assign n568 = x24 & n567 ;
  assign n569 = ~n566 & n568 ;
  assign n570 = ~n565 & n569 ;
  assign n753 = n752 ^ n570 ;
  assign n426 = ~n298 & ~n375 ;
  assign n425 = ~n336 & ~n375 ;
  assign n427 = n426 ^ n425 ;
  assign n337 = n336 ^ n298 ;
  assign n418 = n337 & ~n375 ;
  assign n428 = n427 ^ n418 ;
  assign n417 = ~n298 & ~n336 ;
  assign n419 = n418 ^ n417 ;
  assign n376 = n375 ^ n337 ;
  assign n198 = x32 & ~x40 ;
  assign n165 = x40 ^ x32 ;
  assign n196 = x33 & ~x41 ;
  assign n197 = ~n165 & n196 ;
  assign n199 = n198 ^ n197 ;
  assign n166 = x41 ^ x33 ;
  assign n167 = ~n165 & ~n166 ;
  assign n193 = x34 & ~x42 ;
  assign n168 = x42 ^ x34 ;
  assign n191 = x35 & ~x43 ;
  assign n192 = ~n168 & n191 ;
  assign n194 = n193 ^ n192 ;
  assign n195 = n167 & n194 ;
  assign n200 = n199 ^ n195 ;
  assign n169 = x43 ^ x35 ;
  assign n170 = ~n168 & ~n169 ;
  assign n171 = n167 & n170 ;
  assign n187 = x36 & ~x44 ;
  assign n172 = x44 ^ x36 ;
  assign n185 = x37 & ~x45 ;
  assign n186 = ~n172 & n185 ;
  assign n188 = n187 ^ n186 ;
  assign n173 = x45 ^ x37 ;
  assign n174 = ~n172 & ~n173 ;
  assign n182 = x38 & ~x46 ;
  assign n175 = x46 ^ x38 ;
  assign n180 = x39 & ~x47 ;
  assign n181 = ~n175 & n180 ;
  assign n183 = n182 ^ n181 ;
  assign n184 = n174 & n183 ;
  assign n189 = n188 ^ n184 ;
  assign n190 = n171 & n189 ;
  assign n201 = n200 ^ n190 ;
  assign n176 = x47 ^ x39 ;
  assign n177 = ~n175 & ~n176 ;
  assign n178 = n174 & n177 ;
  assign n179 = n171 & n178 ;
  assign n202 = n201 ^ n179 ;
  assign n415 = n414 ^ n202 ;
  assign n416 = ~n376 & ~n415 ;
  assign n420 = n419 ^ n416 ;
  assign n421 = n202 & ~n414 ;
  assign n422 = n421 ^ n416 ;
  assign n423 = n420 & n422 ;
  assign n424 = n423 ^ n416 ;
  assign n429 = n428 ^ n424 ;
  assign n430 = n421 ^ n420 ;
  assign n431 = n415 ^ n376 ;
  assign n432 = x32 & ~n431 ;
  assign n433 = ~n430 & n432 ;
  assign n434 = ~n429 & n433 ;
  assign n754 = n753 ^ n434 ;
  assign n252 = ~n86 & ~n163 ;
  assign n251 = ~n124 & ~n163 ;
  assign n253 = n252 ^ n251 ;
  assign n125 = n124 ^ n86 ;
  assign n244 = n125 & ~n163 ;
  assign n254 = n253 ^ n244 ;
  assign n243 = ~n86 & ~n124 ;
  assign n245 = n244 ^ n243 ;
  assign n164 = n163 ^ n125 ;
  assign n241 = n240 ^ n202 ;
  assign n242 = ~n164 & n241 ;
  assign n246 = n245 ^ n242 ;
  assign n247 = ~n202 & ~n240 ;
  assign n248 = n247 ^ n242 ;
  assign n249 = n246 & n248 ;
  assign n250 = n249 ^ n242 ;
  assign n255 = n254 ^ n250 ;
  assign n256 = n247 ^ n246 ;
  assign n257 = n241 ^ n164 ;
  assign n258 = x40 & n257 ;
  assign n259 = ~n256 & n258 ;
  assign n260 = ~n255 & n259 ;
  assign n755 = n754 ^ n260 ;
  assign n771 = x1 & ~n747 ;
  assign n772 = ~n746 & n771 ;
  assign n773 = ~n745 & n772 ;
  assign n768 = x9 & n725 ;
  assign n769 = ~n724 & n768 ;
  assign n770 = ~n723 & n769 ;
  assign n774 = n773 ^ n770 ;
  assign n765 = x17 & ~n665 ;
  assign n766 = ~n664 & n765 ;
  assign n767 = ~n663 & n766 ;
  assign n775 = n774 ^ n767 ;
  assign n762 = x25 & n567 ;
  assign n763 = ~n566 & n762 ;
  assign n764 = ~n565 & n763 ;
  assign n776 = n775 ^ n764 ;
  assign n759 = x33 & ~n431 ;
  assign n760 = ~n430 & n759 ;
  assign n761 = ~n429 & n760 ;
  assign n777 = n776 ^ n761 ;
  assign n756 = x41 & n257 ;
  assign n757 = ~n256 & n756 ;
  assign n758 = ~n255 & n757 ;
  assign n778 = n777 ^ n758 ;
  assign n794 = x2 & ~n747 ;
  assign n795 = ~n746 & n794 ;
  assign n796 = ~n745 & n795 ;
  assign n791 = x10 & n725 ;
  assign n792 = ~n724 & n791 ;
  assign n793 = ~n723 & n792 ;
  assign n797 = n796 ^ n793 ;
  assign n788 = x18 & ~n665 ;
  assign n789 = ~n664 & n788 ;
  assign n790 = ~n663 & n789 ;
  assign n798 = n797 ^ n790 ;
  assign n785 = x26 & n567 ;
  assign n786 = ~n566 & n785 ;
  assign n787 = ~n565 & n786 ;
  assign n799 = n798 ^ n787 ;
  assign n782 = x34 & ~n431 ;
  assign n783 = ~n430 & n782 ;
  assign n784 = ~n429 & n783 ;
  assign n800 = n799 ^ n784 ;
  assign n779 = x42 & n257 ;
  assign n780 = ~n256 & n779 ;
  assign n781 = ~n255 & n780 ;
  assign n801 = n800 ^ n781 ;
  assign n817 = x3 & ~n747 ;
  assign n818 = ~n746 & n817 ;
  assign n819 = ~n745 & n818 ;
  assign n814 = x11 & n725 ;
  assign n815 = ~n724 & n814 ;
  assign n816 = ~n723 & n815 ;
  assign n820 = n819 ^ n816 ;
  assign n811 = x19 & ~n665 ;
  assign n812 = ~n664 & n811 ;
  assign n813 = ~n663 & n812 ;
  assign n821 = n820 ^ n813 ;
  assign n808 = x27 & n567 ;
  assign n809 = ~n566 & n808 ;
  assign n810 = ~n565 & n809 ;
  assign n822 = n821 ^ n810 ;
  assign n805 = x35 & ~n431 ;
  assign n806 = ~n430 & n805 ;
  assign n807 = ~n429 & n806 ;
  assign n823 = n822 ^ n807 ;
  assign n802 = x43 & n257 ;
  assign n803 = ~n256 & n802 ;
  assign n804 = ~n255 & n803 ;
  assign n824 = n823 ^ n804 ;
  assign n840 = x4 & ~n747 ;
  assign n841 = ~n746 & n840 ;
  assign n842 = ~n745 & n841 ;
  assign n837 = x12 & n725 ;
  assign n838 = ~n724 & n837 ;
  assign n839 = ~n723 & n838 ;
  assign n843 = n842 ^ n839 ;
  assign n834 = x20 & ~n665 ;
  assign n835 = ~n664 & n834 ;
  assign n836 = ~n663 & n835 ;
  assign n844 = n843 ^ n836 ;
  assign n831 = x28 & n567 ;
  assign n832 = ~n566 & n831 ;
  assign n833 = ~n565 & n832 ;
  assign n845 = n844 ^ n833 ;
  assign n828 = x36 & ~n431 ;
  assign n829 = ~n430 & n828 ;
  assign n830 = ~n429 & n829 ;
  assign n846 = n845 ^ n830 ;
  assign n825 = x44 & n257 ;
  assign n826 = ~n256 & n825 ;
  assign n827 = ~n255 & n826 ;
  assign n847 = n846 ^ n827 ;
  assign n863 = x5 & ~n747 ;
  assign n864 = ~n746 & n863 ;
  assign n865 = ~n745 & n864 ;
  assign n860 = x13 & n725 ;
  assign n861 = ~n724 & n860 ;
  assign n862 = ~n723 & n861 ;
  assign n866 = n865 ^ n862 ;
  assign n857 = x21 & ~n665 ;
  assign n858 = ~n664 & n857 ;
  assign n859 = ~n663 & n858 ;
  assign n867 = n866 ^ n859 ;
  assign n854 = x29 & n567 ;
  assign n855 = ~n566 & n854 ;
  assign n856 = ~n565 & n855 ;
  assign n868 = n867 ^ n856 ;
  assign n851 = x37 & ~n431 ;
  assign n852 = ~n430 & n851 ;
  assign n853 = ~n429 & n852 ;
  assign n869 = n868 ^ n853 ;
  assign n848 = x45 & n257 ;
  assign n849 = ~n256 & n848 ;
  assign n850 = ~n255 & n849 ;
  assign n870 = n869 ^ n850 ;
  assign n886 = x6 & ~n747 ;
  assign n887 = ~n746 & n886 ;
  assign n888 = ~n745 & n887 ;
  assign n883 = x14 & n725 ;
  assign n884 = ~n724 & n883 ;
  assign n885 = ~n723 & n884 ;
  assign n889 = n888 ^ n885 ;
  assign n880 = x22 & ~n665 ;
  assign n881 = ~n664 & n880 ;
  assign n882 = ~n663 & n881 ;
  assign n890 = n889 ^ n882 ;
  assign n877 = x30 & n567 ;
  assign n878 = ~n566 & n877 ;
  assign n879 = ~n565 & n878 ;
  assign n891 = n890 ^ n879 ;
  assign n874 = x38 & ~n431 ;
  assign n875 = ~n430 & n874 ;
  assign n876 = ~n429 & n875 ;
  assign n892 = n891 ^ n876 ;
  assign n871 = x46 & n257 ;
  assign n872 = ~n256 & n871 ;
  assign n873 = ~n255 & n872 ;
  assign n893 = n892 ^ n873 ;
  assign n909 = x7 & ~n747 ;
  assign n910 = ~n746 & n909 ;
  assign n911 = ~n745 & n910 ;
  assign n906 = x15 & n725 ;
  assign n907 = ~n724 & n906 ;
  assign n908 = ~n723 & n907 ;
  assign n912 = n911 ^ n908 ;
  assign n903 = x23 & ~n665 ;
  assign n904 = ~n664 & n903 ;
  assign n905 = ~n663 & n904 ;
  assign n913 = n912 ^ n905 ;
  assign n900 = x31 & n567 ;
  assign n901 = ~n566 & n900 ;
  assign n902 = ~n565 & n901 ;
  assign n914 = n913 ^ n902 ;
  assign n897 = x39 & ~n431 ;
  assign n898 = ~n430 & n897 ;
  assign n899 = ~n429 & n898 ;
  assign n915 = n914 ^ n899 ;
  assign n894 = x47 & n257 ;
  assign n895 = ~n256 & n894 ;
  assign n896 = ~n255 & n895 ;
  assign n916 = n915 ^ n896 ;
  assign n932 = x0 & n747 ;
  assign n933 = ~n746 & n932 ;
  assign n934 = ~n745 & n933 ;
  assign n929 = x8 & ~n725 ;
  assign n930 = ~n724 & n929 ;
  assign n931 = ~n723 & n930 ;
  assign n935 = n934 ^ n931 ;
  assign n926 = x16 & n665 ;
  assign n927 = ~n664 & n926 ;
  assign n928 = ~n663 & n927 ;
  assign n936 = n935 ^ n928 ;
  assign n923 = x24 & ~n567 ;
  assign n924 = ~n566 & n923 ;
  assign n925 = ~n565 & n924 ;
  assign n937 = n936 ^ n925 ;
  assign n920 = x32 & n431 ;
  assign n921 = ~n430 & n920 ;
  assign n922 = ~n429 & n921 ;
  assign n938 = n937 ^ n922 ;
  assign n917 = x40 & ~n257 ;
  assign n918 = ~n256 & n917 ;
  assign n919 = ~n255 & n918 ;
  assign n939 = n938 ^ n919 ;
  assign n955 = x1 & n747 ;
  assign n956 = ~n746 & n955 ;
  assign n957 = ~n745 & n956 ;
  assign n952 = x9 & ~n725 ;
  assign n953 = ~n724 & n952 ;
  assign n954 = ~n723 & n953 ;
  assign n958 = n957 ^ n954 ;
  assign n949 = x17 & n665 ;
  assign n950 = ~n664 & n949 ;
  assign n951 = ~n663 & n950 ;
  assign n959 = n958 ^ n951 ;
  assign n946 = x25 & ~n567 ;
  assign n947 = ~n566 & n946 ;
  assign n948 = ~n565 & n947 ;
  assign n960 = n959 ^ n948 ;
  assign n943 = x33 & n431 ;
  assign n944 = ~n430 & n943 ;
  assign n945 = ~n429 & n944 ;
  assign n961 = n960 ^ n945 ;
  assign n940 = x41 & ~n257 ;
  assign n941 = ~n256 & n940 ;
  assign n942 = ~n255 & n941 ;
  assign n962 = n961 ^ n942 ;
  assign n978 = x2 & n747 ;
  assign n979 = ~n746 & n978 ;
  assign n980 = ~n745 & n979 ;
  assign n975 = x10 & ~n725 ;
  assign n976 = ~n724 & n975 ;
  assign n977 = ~n723 & n976 ;
  assign n981 = n980 ^ n977 ;
  assign n972 = x18 & n665 ;
  assign n973 = ~n664 & n972 ;
  assign n974 = ~n663 & n973 ;
  assign n982 = n981 ^ n974 ;
  assign n969 = x26 & ~n567 ;
  assign n970 = ~n566 & n969 ;
  assign n971 = ~n565 & n970 ;
  assign n983 = n982 ^ n971 ;
  assign n966 = x34 & n431 ;
  assign n967 = ~n430 & n966 ;
  assign n968 = ~n429 & n967 ;
  assign n984 = n983 ^ n968 ;
  assign n963 = x42 & ~n257 ;
  assign n964 = ~n256 & n963 ;
  assign n965 = ~n255 & n964 ;
  assign n985 = n984 ^ n965 ;
  assign n1001 = x3 & n747 ;
  assign n1002 = ~n746 & n1001 ;
  assign n1003 = ~n745 & n1002 ;
  assign n998 = x11 & ~n725 ;
  assign n999 = ~n724 & n998 ;
  assign n1000 = ~n723 & n999 ;
  assign n1004 = n1003 ^ n1000 ;
  assign n995 = x19 & n665 ;
  assign n996 = ~n664 & n995 ;
  assign n997 = ~n663 & n996 ;
  assign n1005 = n1004 ^ n997 ;
  assign n992 = x27 & ~n567 ;
  assign n993 = ~n566 & n992 ;
  assign n994 = ~n565 & n993 ;
  assign n1006 = n1005 ^ n994 ;
  assign n989 = x35 & n431 ;
  assign n990 = ~n430 & n989 ;
  assign n991 = ~n429 & n990 ;
  assign n1007 = n1006 ^ n991 ;
  assign n986 = x43 & ~n257 ;
  assign n987 = ~n256 & n986 ;
  assign n988 = ~n255 & n987 ;
  assign n1008 = n1007 ^ n988 ;
  assign n1024 = x4 & n747 ;
  assign n1025 = ~n746 & n1024 ;
  assign n1026 = ~n745 & n1025 ;
  assign n1021 = x12 & ~n725 ;
  assign n1022 = ~n724 & n1021 ;
  assign n1023 = ~n723 & n1022 ;
  assign n1027 = n1026 ^ n1023 ;
  assign n1018 = x20 & n665 ;
  assign n1019 = ~n664 & n1018 ;
  assign n1020 = ~n663 & n1019 ;
  assign n1028 = n1027 ^ n1020 ;
  assign n1015 = x28 & ~n567 ;
  assign n1016 = ~n566 & n1015 ;
  assign n1017 = ~n565 & n1016 ;
  assign n1029 = n1028 ^ n1017 ;
  assign n1012 = x36 & n431 ;
  assign n1013 = ~n430 & n1012 ;
  assign n1014 = ~n429 & n1013 ;
  assign n1030 = n1029 ^ n1014 ;
  assign n1009 = x44 & ~n257 ;
  assign n1010 = ~n256 & n1009 ;
  assign n1011 = ~n255 & n1010 ;
  assign n1031 = n1030 ^ n1011 ;
  assign n1047 = x5 & n747 ;
  assign n1048 = ~n746 & n1047 ;
  assign n1049 = ~n745 & n1048 ;
  assign n1044 = x13 & ~n725 ;
  assign n1045 = ~n724 & n1044 ;
  assign n1046 = ~n723 & n1045 ;
  assign n1050 = n1049 ^ n1046 ;
  assign n1041 = x21 & n665 ;
  assign n1042 = ~n664 & n1041 ;
  assign n1043 = ~n663 & n1042 ;
  assign n1051 = n1050 ^ n1043 ;
  assign n1038 = x29 & ~n567 ;
  assign n1039 = ~n566 & n1038 ;
  assign n1040 = ~n565 & n1039 ;
  assign n1052 = n1051 ^ n1040 ;
  assign n1035 = x37 & n431 ;
  assign n1036 = ~n430 & n1035 ;
  assign n1037 = ~n429 & n1036 ;
  assign n1053 = n1052 ^ n1037 ;
  assign n1032 = x45 & ~n257 ;
  assign n1033 = ~n256 & n1032 ;
  assign n1034 = ~n255 & n1033 ;
  assign n1054 = n1053 ^ n1034 ;
  assign n1070 = x6 & n747 ;
  assign n1071 = ~n746 & n1070 ;
  assign n1072 = ~n745 & n1071 ;
  assign n1067 = x14 & ~n725 ;
  assign n1068 = ~n724 & n1067 ;
  assign n1069 = ~n723 & n1068 ;
  assign n1073 = n1072 ^ n1069 ;
  assign n1064 = x22 & n665 ;
  assign n1065 = ~n664 & n1064 ;
  assign n1066 = ~n663 & n1065 ;
  assign n1074 = n1073 ^ n1066 ;
  assign n1061 = x30 & ~n567 ;
  assign n1062 = ~n566 & n1061 ;
  assign n1063 = ~n565 & n1062 ;
  assign n1075 = n1074 ^ n1063 ;
  assign n1058 = x38 & n431 ;
  assign n1059 = ~n430 & n1058 ;
  assign n1060 = ~n429 & n1059 ;
  assign n1076 = n1075 ^ n1060 ;
  assign n1055 = x46 & ~n257 ;
  assign n1056 = ~n256 & n1055 ;
  assign n1057 = ~n255 & n1056 ;
  assign n1077 = n1076 ^ n1057 ;
  assign n1093 = x7 & n747 ;
  assign n1094 = ~n746 & n1093 ;
  assign n1095 = ~n745 & n1094 ;
  assign n1090 = x15 & ~n725 ;
  assign n1091 = ~n724 & n1090 ;
  assign n1092 = ~n723 & n1091 ;
  assign n1096 = n1095 ^ n1092 ;
  assign n1087 = x23 & n665 ;
  assign n1088 = ~n664 & n1087 ;
  assign n1089 = ~n663 & n1088 ;
  assign n1097 = n1096 ^ n1089 ;
  assign n1084 = x31 & ~n567 ;
  assign n1085 = ~n566 & n1084 ;
  assign n1086 = ~n565 & n1085 ;
  assign n1098 = n1097 ^ n1086 ;
  assign n1081 = x39 & n431 ;
  assign n1082 = ~n430 & n1081 ;
  assign n1083 = ~n429 & n1082 ;
  assign n1099 = n1098 ^ n1083 ;
  assign n1078 = x47 & ~n257 ;
  assign n1079 = ~n256 & n1078 ;
  assign n1080 = ~n255 & n1079 ;
  assign n1100 = n1099 ^ n1080 ;
  assign n1111 = n746 & n748 ;
  assign n1112 = ~n745 & n1111 ;
  assign n1109 = n724 & n726 ;
  assign n1110 = ~n723 & n1109 ;
  assign n1113 = n1112 ^ n1110 ;
  assign n1107 = n664 & n666 ;
  assign n1108 = ~n663 & n1107 ;
  assign n1114 = n1113 ^ n1108 ;
  assign n1105 = n566 & n568 ;
  assign n1106 = ~n565 & n1105 ;
  assign n1115 = n1114 ^ n1106 ;
  assign n1103 = n430 & n432 ;
  assign n1104 = ~n429 & n1103 ;
  assign n1116 = n1115 ^ n1104 ;
  assign n1101 = n256 & n258 ;
  assign n1102 = ~n255 & n1101 ;
  assign n1117 = n1116 ^ n1102 ;
  assign n1128 = n746 & n771 ;
  assign n1129 = ~n745 & n1128 ;
  assign n1126 = n724 & n768 ;
  assign n1127 = ~n723 & n1126 ;
  assign n1130 = n1129 ^ n1127 ;
  assign n1124 = n664 & n765 ;
  assign n1125 = ~n663 & n1124 ;
  assign n1131 = n1130 ^ n1125 ;
  assign n1122 = n566 & n762 ;
  assign n1123 = ~n565 & n1122 ;
  assign n1132 = n1131 ^ n1123 ;
  assign n1120 = n430 & n759 ;
  assign n1121 = ~n429 & n1120 ;
  assign n1133 = n1132 ^ n1121 ;
  assign n1118 = n256 & n756 ;
  assign n1119 = ~n255 & n1118 ;
  assign n1134 = n1133 ^ n1119 ;
  assign n1145 = n746 & n794 ;
  assign n1146 = ~n745 & n1145 ;
  assign n1143 = n724 & n791 ;
  assign n1144 = ~n723 & n1143 ;
  assign n1147 = n1146 ^ n1144 ;
  assign n1141 = n664 & n788 ;
  assign n1142 = ~n663 & n1141 ;
  assign n1148 = n1147 ^ n1142 ;
  assign n1139 = n566 & n785 ;
  assign n1140 = ~n565 & n1139 ;
  assign n1149 = n1148 ^ n1140 ;
  assign n1137 = n430 & n782 ;
  assign n1138 = ~n429 & n1137 ;
  assign n1150 = n1149 ^ n1138 ;
  assign n1135 = n256 & n779 ;
  assign n1136 = ~n255 & n1135 ;
  assign n1151 = n1150 ^ n1136 ;
  assign n1162 = n746 & n817 ;
  assign n1163 = ~n745 & n1162 ;
  assign n1160 = n724 & n814 ;
  assign n1161 = ~n723 & n1160 ;
  assign n1164 = n1163 ^ n1161 ;
  assign n1158 = n664 & n811 ;
  assign n1159 = ~n663 & n1158 ;
  assign n1165 = n1164 ^ n1159 ;
  assign n1156 = n566 & n808 ;
  assign n1157 = ~n565 & n1156 ;
  assign n1166 = n1165 ^ n1157 ;
  assign n1154 = n430 & n805 ;
  assign n1155 = ~n429 & n1154 ;
  assign n1167 = n1166 ^ n1155 ;
  assign n1152 = n256 & n802 ;
  assign n1153 = ~n255 & n1152 ;
  assign n1168 = n1167 ^ n1153 ;
  assign n1179 = n746 & n840 ;
  assign n1180 = ~n745 & n1179 ;
  assign n1177 = n724 & n837 ;
  assign n1178 = ~n723 & n1177 ;
  assign n1181 = n1180 ^ n1178 ;
  assign n1175 = n664 & n834 ;
  assign n1176 = ~n663 & n1175 ;
  assign n1182 = n1181 ^ n1176 ;
  assign n1173 = n566 & n831 ;
  assign n1174 = ~n565 & n1173 ;
  assign n1183 = n1182 ^ n1174 ;
  assign n1171 = n430 & n828 ;
  assign n1172 = ~n429 & n1171 ;
  assign n1184 = n1183 ^ n1172 ;
  assign n1169 = n256 & n825 ;
  assign n1170 = ~n255 & n1169 ;
  assign n1185 = n1184 ^ n1170 ;
  assign n1196 = n746 & n863 ;
  assign n1197 = ~n745 & n1196 ;
  assign n1194 = n724 & n860 ;
  assign n1195 = ~n723 & n1194 ;
  assign n1198 = n1197 ^ n1195 ;
  assign n1192 = n664 & n857 ;
  assign n1193 = ~n663 & n1192 ;
  assign n1199 = n1198 ^ n1193 ;
  assign n1190 = n566 & n854 ;
  assign n1191 = ~n565 & n1190 ;
  assign n1200 = n1199 ^ n1191 ;
  assign n1188 = n430 & n851 ;
  assign n1189 = ~n429 & n1188 ;
  assign n1201 = n1200 ^ n1189 ;
  assign n1186 = n256 & n848 ;
  assign n1187 = ~n255 & n1186 ;
  assign n1202 = n1201 ^ n1187 ;
  assign n1213 = n746 & n886 ;
  assign n1214 = ~n745 & n1213 ;
  assign n1211 = n724 & n883 ;
  assign n1212 = ~n723 & n1211 ;
  assign n1215 = n1214 ^ n1212 ;
  assign n1209 = n664 & n880 ;
  assign n1210 = ~n663 & n1209 ;
  assign n1216 = n1215 ^ n1210 ;
  assign n1207 = n566 & n877 ;
  assign n1208 = ~n565 & n1207 ;
  assign n1217 = n1216 ^ n1208 ;
  assign n1205 = n430 & n874 ;
  assign n1206 = ~n429 & n1205 ;
  assign n1218 = n1217 ^ n1206 ;
  assign n1203 = n256 & n871 ;
  assign n1204 = ~n255 & n1203 ;
  assign n1219 = n1218 ^ n1204 ;
  assign n1230 = n746 & n909 ;
  assign n1231 = ~n745 & n1230 ;
  assign n1228 = n724 & n906 ;
  assign n1229 = ~n723 & n1228 ;
  assign n1232 = n1231 ^ n1229 ;
  assign n1226 = n664 & n903 ;
  assign n1227 = ~n663 & n1226 ;
  assign n1233 = n1232 ^ n1227 ;
  assign n1224 = n566 & n900 ;
  assign n1225 = ~n565 & n1224 ;
  assign n1234 = n1233 ^ n1225 ;
  assign n1222 = n430 & n897 ;
  assign n1223 = ~n429 & n1222 ;
  assign n1235 = n1234 ^ n1223 ;
  assign n1220 = n256 & n894 ;
  assign n1221 = ~n255 & n1220 ;
  assign n1236 = n1235 ^ n1221 ;
  assign n1247 = n746 & n932 ;
  assign n1248 = ~n745 & n1247 ;
  assign n1245 = n724 & n929 ;
  assign n1246 = ~n723 & n1245 ;
  assign n1249 = n1248 ^ n1246 ;
  assign n1243 = n664 & n926 ;
  assign n1244 = ~n663 & n1243 ;
  assign n1250 = n1249 ^ n1244 ;
  assign n1241 = n566 & n923 ;
  assign n1242 = ~n565 & n1241 ;
  assign n1251 = n1250 ^ n1242 ;
  assign n1239 = n430 & n920 ;
  assign n1240 = ~n429 & n1239 ;
  assign n1252 = n1251 ^ n1240 ;
  assign n1237 = n256 & n917 ;
  assign n1238 = ~n255 & n1237 ;
  assign n1253 = n1252 ^ n1238 ;
  assign n1264 = n746 & n955 ;
  assign n1265 = ~n745 & n1264 ;
  assign n1262 = n724 & n952 ;
  assign n1263 = ~n723 & n1262 ;
  assign n1266 = n1265 ^ n1263 ;
  assign n1260 = n664 & n949 ;
  assign n1261 = ~n663 & n1260 ;
  assign n1267 = n1266 ^ n1261 ;
  assign n1258 = n566 & n946 ;
  assign n1259 = ~n565 & n1258 ;
  assign n1268 = n1267 ^ n1259 ;
  assign n1256 = n430 & n943 ;
  assign n1257 = ~n429 & n1256 ;
  assign n1269 = n1268 ^ n1257 ;
  assign n1254 = n256 & n940 ;
  assign n1255 = ~n255 & n1254 ;
  assign n1270 = n1269 ^ n1255 ;
  assign n1281 = n746 & n978 ;
  assign n1282 = ~n745 & n1281 ;
  assign n1279 = n724 & n975 ;
  assign n1280 = ~n723 & n1279 ;
  assign n1283 = n1282 ^ n1280 ;
  assign n1277 = n664 & n972 ;
  assign n1278 = ~n663 & n1277 ;
  assign n1284 = n1283 ^ n1278 ;
  assign n1275 = n566 & n969 ;
  assign n1276 = ~n565 & n1275 ;
  assign n1285 = n1284 ^ n1276 ;
  assign n1273 = n430 & n966 ;
  assign n1274 = ~n429 & n1273 ;
  assign n1286 = n1285 ^ n1274 ;
  assign n1271 = n256 & n963 ;
  assign n1272 = ~n255 & n1271 ;
  assign n1287 = n1286 ^ n1272 ;
  assign n1298 = n746 & n1001 ;
  assign n1299 = ~n745 & n1298 ;
  assign n1296 = n724 & n998 ;
  assign n1297 = ~n723 & n1296 ;
  assign n1300 = n1299 ^ n1297 ;
  assign n1294 = n664 & n995 ;
  assign n1295 = ~n663 & n1294 ;
  assign n1301 = n1300 ^ n1295 ;
  assign n1292 = n566 & n992 ;
  assign n1293 = ~n565 & n1292 ;
  assign n1302 = n1301 ^ n1293 ;
  assign n1290 = n430 & n989 ;
  assign n1291 = ~n429 & n1290 ;
  assign n1303 = n1302 ^ n1291 ;
  assign n1288 = n256 & n986 ;
  assign n1289 = ~n255 & n1288 ;
  assign n1304 = n1303 ^ n1289 ;
  assign n1315 = n746 & n1024 ;
  assign n1316 = ~n745 & n1315 ;
  assign n1313 = n724 & n1021 ;
  assign n1314 = ~n723 & n1313 ;
  assign n1317 = n1316 ^ n1314 ;
  assign n1311 = n664 & n1018 ;
  assign n1312 = ~n663 & n1311 ;
  assign n1318 = n1317 ^ n1312 ;
  assign n1309 = n566 & n1015 ;
  assign n1310 = ~n565 & n1309 ;
  assign n1319 = n1318 ^ n1310 ;
  assign n1307 = n430 & n1012 ;
  assign n1308 = ~n429 & n1307 ;
  assign n1320 = n1319 ^ n1308 ;
  assign n1305 = n256 & n1009 ;
  assign n1306 = ~n255 & n1305 ;
  assign n1321 = n1320 ^ n1306 ;
  assign n1332 = n746 & n1047 ;
  assign n1333 = ~n745 & n1332 ;
  assign n1330 = n724 & n1044 ;
  assign n1331 = ~n723 & n1330 ;
  assign n1334 = n1333 ^ n1331 ;
  assign n1328 = n664 & n1041 ;
  assign n1329 = ~n663 & n1328 ;
  assign n1335 = n1334 ^ n1329 ;
  assign n1326 = n566 & n1038 ;
  assign n1327 = ~n565 & n1326 ;
  assign n1336 = n1335 ^ n1327 ;
  assign n1324 = n430 & n1035 ;
  assign n1325 = ~n429 & n1324 ;
  assign n1337 = n1336 ^ n1325 ;
  assign n1322 = n256 & n1032 ;
  assign n1323 = ~n255 & n1322 ;
  assign n1338 = n1337 ^ n1323 ;
  assign n1349 = n746 & n1070 ;
  assign n1350 = ~n745 & n1349 ;
  assign n1347 = n724 & n1067 ;
  assign n1348 = ~n723 & n1347 ;
  assign n1351 = n1350 ^ n1348 ;
  assign n1345 = n664 & n1064 ;
  assign n1346 = ~n663 & n1345 ;
  assign n1352 = n1351 ^ n1346 ;
  assign n1343 = n566 & n1061 ;
  assign n1344 = ~n565 & n1343 ;
  assign n1353 = n1352 ^ n1344 ;
  assign n1341 = n430 & n1058 ;
  assign n1342 = ~n429 & n1341 ;
  assign n1354 = n1353 ^ n1342 ;
  assign n1339 = n256 & n1055 ;
  assign n1340 = ~n255 & n1339 ;
  assign n1355 = n1354 ^ n1340 ;
  assign n1366 = n746 & n1093 ;
  assign n1367 = ~n745 & n1366 ;
  assign n1364 = n724 & n1090 ;
  assign n1365 = ~n723 & n1364 ;
  assign n1368 = n1367 ^ n1365 ;
  assign n1362 = n664 & n1087 ;
  assign n1363 = ~n663 & n1362 ;
  assign n1369 = n1368 ^ n1363 ;
  assign n1360 = n566 & n1084 ;
  assign n1361 = ~n565 & n1360 ;
  assign n1370 = n1369 ^ n1361 ;
  assign n1358 = n430 & n1081 ;
  assign n1359 = ~n429 & n1358 ;
  assign n1371 = n1370 ^ n1359 ;
  assign n1356 = n256 & n1078 ;
  assign n1357 = ~n255 & n1356 ;
  assign n1372 = n1371 ^ n1357 ;
  assign n1378 = n745 & n749 ;
  assign n1377 = n723 & n727 ;
  assign n1379 = n1378 ^ n1377 ;
  assign n1376 = n663 & n667 ;
  assign n1380 = n1379 ^ n1376 ;
  assign n1375 = n565 & n569 ;
  assign n1381 = n1380 ^ n1375 ;
  assign n1374 = n429 & n433 ;
  assign n1382 = n1381 ^ n1374 ;
  assign n1373 = n255 & n259 ;
  assign n1383 = n1382 ^ n1373 ;
  assign n1389 = n745 & n772 ;
  assign n1388 = n723 & n769 ;
  assign n1390 = n1389 ^ n1388 ;
  assign n1387 = n663 & n766 ;
  assign n1391 = n1390 ^ n1387 ;
  assign n1386 = n565 & n763 ;
  assign n1392 = n1391 ^ n1386 ;
  assign n1385 = n429 & n760 ;
  assign n1393 = n1392 ^ n1385 ;
  assign n1384 = n255 & n757 ;
  assign n1394 = n1393 ^ n1384 ;
  assign n1400 = n745 & n795 ;
  assign n1399 = n723 & n792 ;
  assign n1401 = n1400 ^ n1399 ;
  assign n1398 = n663 & n789 ;
  assign n1402 = n1401 ^ n1398 ;
  assign n1397 = n565 & n786 ;
  assign n1403 = n1402 ^ n1397 ;
  assign n1396 = n429 & n783 ;
  assign n1404 = n1403 ^ n1396 ;
  assign n1395 = n255 & n780 ;
  assign n1405 = n1404 ^ n1395 ;
  assign n1411 = n745 & n818 ;
  assign n1410 = n723 & n815 ;
  assign n1412 = n1411 ^ n1410 ;
  assign n1409 = n663 & n812 ;
  assign n1413 = n1412 ^ n1409 ;
  assign n1408 = n565 & n809 ;
  assign n1414 = n1413 ^ n1408 ;
  assign n1407 = n429 & n806 ;
  assign n1415 = n1414 ^ n1407 ;
  assign n1406 = n255 & n803 ;
  assign n1416 = n1415 ^ n1406 ;
  assign n1422 = n745 & n841 ;
  assign n1421 = n723 & n838 ;
  assign n1423 = n1422 ^ n1421 ;
  assign n1420 = n663 & n835 ;
  assign n1424 = n1423 ^ n1420 ;
  assign n1419 = n565 & n832 ;
  assign n1425 = n1424 ^ n1419 ;
  assign n1418 = n429 & n829 ;
  assign n1426 = n1425 ^ n1418 ;
  assign n1417 = n255 & n826 ;
  assign n1427 = n1426 ^ n1417 ;
  assign n1433 = n745 & n864 ;
  assign n1432 = n723 & n861 ;
  assign n1434 = n1433 ^ n1432 ;
  assign n1431 = n663 & n858 ;
  assign n1435 = n1434 ^ n1431 ;
  assign n1430 = n565 & n855 ;
  assign n1436 = n1435 ^ n1430 ;
  assign n1429 = n429 & n852 ;
  assign n1437 = n1436 ^ n1429 ;
  assign n1428 = n255 & n849 ;
  assign n1438 = n1437 ^ n1428 ;
  assign n1444 = n745 & n887 ;
  assign n1443 = n723 & n884 ;
  assign n1445 = n1444 ^ n1443 ;
  assign n1442 = n663 & n881 ;
  assign n1446 = n1445 ^ n1442 ;
  assign n1441 = n565 & n878 ;
  assign n1447 = n1446 ^ n1441 ;
  assign n1440 = n429 & n875 ;
  assign n1448 = n1447 ^ n1440 ;
  assign n1439 = n255 & n872 ;
  assign n1449 = n1448 ^ n1439 ;
  assign n1455 = n745 & n910 ;
  assign n1454 = n723 & n907 ;
  assign n1456 = n1455 ^ n1454 ;
  assign n1453 = n663 & n904 ;
  assign n1457 = n1456 ^ n1453 ;
  assign n1452 = n565 & n901 ;
  assign n1458 = n1457 ^ n1452 ;
  assign n1451 = n429 & n898 ;
  assign n1459 = n1458 ^ n1451 ;
  assign n1450 = n255 & n895 ;
  assign n1460 = n1459 ^ n1450 ;
  assign n1466 = n745 & n933 ;
  assign n1465 = n723 & n930 ;
  assign n1467 = n1466 ^ n1465 ;
  assign n1464 = n663 & n927 ;
  assign n1468 = n1467 ^ n1464 ;
  assign n1463 = n565 & n924 ;
  assign n1469 = n1468 ^ n1463 ;
  assign n1462 = n429 & n921 ;
  assign n1470 = n1469 ^ n1462 ;
  assign n1461 = n255 & n918 ;
  assign n1471 = n1470 ^ n1461 ;
  assign n1477 = n745 & n956 ;
  assign n1476 = n723 & n953 ;
  assign n1478 = n1477 ^ n1476 ;
  assign n1475 = n663 & n950 ;
  assign n1479 = n1478 ^ n1475 ;
  assign n1474 = n565 & n947 ;
  assign n1480 = n1479 ^ n1474 ;
  assign n1473 = n429 & n944 ;
  assign n1481 = n1480 ^ n1473 ;
  assign n1472 = n255 & n941 ;
  assign n1482 = n1481 ^ n1472 ;
  assign n1488 = n745 & n979 ;
  assign n1487 = n723 & n976 ;
  assign n1489 = n1488 ^ n1487 ;
  assign n1486 = n663 & n973 ;
  assign n1490 = n1489 ^ n1486 ;
  assign n1485 = n565 & n970 ;
  assign n1491 = n1490 ^ n1485 ;
  assign n1484 = n429 & n967 ;
  assign n1492 = n1491 ^ n1484 ;
  assign n1483 = n255 & n964 ;
  assign n1493 = n1492 ^ n1483 ;
  assign n1499 = n745 & n1002 ;
  assign n1498 = n723 & n999 ;
  assign n1500 = n1499 ^ n1498 ;
  assign n1497 = n663 & n996 ;
  assign n1501 = n1500 ^ n1497 ;
  assign n1496 = n565 & n993 ;
  assign n1502 = n1501 ^ n1496 ;
  assign n1495 = n429 & n990 ;
  assign n1503 = n1502 ^ n1495 ;
  assign n1494 = n255 & n987 ;
  assign n1504 = n1503 ^ n1494 ;
  assign n1510 = n745 & n1025 ;
  assign n1509 = n723 & n1022 ;
  assign n1511 = n1510 ^ n1509 ;
  assign n1508 = n663 & n1019 ;
  assign n1512 = n1511 ^ n1508 ;
  assign n1507 = n565 & n1016 ;
  assign n1513 = n1512 ^ n1507 ;
  assign n1506 = n429 & n1013 ;
  assign n1514 = n1513 ^ n1506 ;
  assign n1505 = n255 & n1010 ;
  assign n1515 = n1514 ^ n1505 ;
  assign n1521 = n745 & n1048 ;
  assign n1520 = n723 & n1045 ;
  assign n1522 = n1521 ^ n1520 ;
  assign n1519 = n663 & n1042 ;
  assign n1523 = n1522 ^ n1519 ;
  assign n1518 = n565 & n1039 ;
  assign n1524 = n1523 ^ n1518 ;
  assign n1517 = n429 & n1036 ;
  assign n1525 = n1524 ^ n1517 ;
  assign n1516 = n255 & n1033 ;
  assign n1526 = n1525 ^ n1516 ;
  assign n1532 = n745 & n1071 ;
  assign n1531 = n723 & n1068 ;
  assign n1533 = n1532 ^ n1531 ;
  assign n1530 = n663 & n1065 ;
  assign n1534 = n1533 ^ n1530 ;
  assign n1529 = n565 & n1062 ;
  assign n1535 = n1534 ^ n1529 ;
  assign n1528 = n429 & n1059 ;
  assign n1536 = n1535 ^ n1528 ;
  assign n1527 = n255 & n1056 ;
  assign n1537 = n1536 ^ n1527 ;
  assign n1543 = n745 & n1094 ;
  assign n1542 = n723 & n1091 ;
  assign n1544 = n1543 ^ n1542 ;
  assign n1541 = n663 & n1088 ;
  assign n1545 = n1544 ^ n1541 ;
  assign n1540 = n565 & n1085 ;
  assign n1546 = n1545 ^ n1540 ;
  assign n1539 = n429 & n1082 ;
  assign n1547 = n1546 ^ n1539 ;
  assign n1538 = n255 & n1079 ;
  assign n1548 = n1547 ^ n1538 ;
  assign y0 = n755 ;
  assign y1 = n778 ;
  assign y2 = n801 ;
  assign y3 = n824 ;
  assign y4 = n847 ;
  assign y5 = n870 ;
  assign y6 = n893 ;
  assign y7 = n916 ;
  assign y8 = n939 ;
  assign y9 = n962 ;
  assign y10 = n985 ;
  assign y11 = n1008 ;
  assign y12 = n1031 ;
  assign y13 = n1054 ;
  assign y14 = n1077 ;
  assign y15 = n1100 ;
  assign y16 = n1117 ;
  assign y17 = n1134 ;
  assign y18 = n1151 ;
  assign y19 = n1168 ;
  assign y20 = n1185 ;
  assign y21 = n1202 ;
  assign y22 = n1219 ;
  assign y23 = n1236 ;
  assign y24 = n1253 ;
  assign y25 = n1270 ;
  assign y26 = n1287 ;
  assign y27 = n1304 ;
  assign y28 = n1321 ;
  assign y29 = n1338 ;
  assign y30 = n1355 ;
  assign y31 = n1372 ;
  assign y32 = n1383 ;
  assign y33 = n1394 ;
  assign y34 = n1405 ;
  assign y35 = n1416 ;
  assign y36 = n1427 ;
  assign y37 = n1438 ;
  assign y38 = n1449 ;
  assign y39 = n1460 ;
  assign y40 = n1471 ;
  assign y41 = n1482 ;
  assign y42 = n1493 ;
  assign y43 = n1504 ;
  assign y44 = n1515 ;
  assign y45 = n1526 ;
  assign y46 = n1537 ;
  assign y47 = n1548 ;
endmodule
