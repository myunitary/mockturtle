module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 ;
  assign n345 = ~x6 & x8 ;
  assign n346 = x5 & ~n345 ;
  assign n347 = x6 & x9 ;
  assign n348 = n347 ^ x6 ;
  assign n349 = n348 ^ x9 ;
  assign n350 = x4 & x8 ;
  assign n351 = n349 & ~n350 ;
  assign n352 = n346 & ~n351 ;
  assign n353 = x6 & ~x9 ;
  assign n354 = x4 & x9 ;
  assign n355 = ~n353 & ~n354 ;
  assign n356 = x5 & x6 ;
  assign n357 = ~x8 & ~n356 ;
  assign n358 = ~n355 & n357 ;
  assign n359 = ~n352 & ~n358 ;
  assign n360 = x1 & x3 ;
  assign n361 = n360 ^ x1 ;
  assign n362 = n361 ^ x3 ;
  assign n306 = x0 & x2 ;
  assign n307 = n306 ^ x0 ;
  assign n308 = n307 ^ x2 ;
  assign n363 = ~x7 & ~n308 ;
  assign n364 = ~n362 & n363 ;
  assign n365 = ~n359 & n364 ;
  assign n11 = x0 & x9 ;
  assign n12 = n11 ^ x9 ;
  assign n13 = x1 & n12 ;
  assign n14 = n13 ^ x1 ;
  assign n15 = x1 & x9 ;
  assign n16 = n15 ^ x9 ;
  assign n17 = x3 & x5 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = n18 ^ x5 ;
  assign n20 = n16 & n19 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n14 & n22 ;
  assign n24 = n23 ^ n14 ;
  assign n25 = n24 ^ n22 ;
  assign n30 = n11 ^ x0 ;
  assign n31 = x1 & x7 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = n32 ^ x7 ;
  assign n34 = n30 & ~n33 ;
  assign n35 = n34 ^ n33 ;
  assign n26 = n15 ^ x1 ;
  assign n27 = x7 & n26 ;
  assign n28 = n27 ^ x7 ;
  assign n29 = n28 ^ n26 ;
  assign n36 = n35 ^ n29 ;
  assign n42 = x2 & ~n36 ;
  assign n43 = n25 & n42 ;
  assign n44 = n43 ^ x2 ;
  assign n37 = n25 & ~n36 ;
  assign n38 = n37 ^ n25 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ n25 ;
  assign n41 = n40 ^ n36 ;
  assign n45 = n44 ^ n41 ;
  assign n128 = n45 ^ x8 ;
  assign n46 = x2 ^ x0 ;
  assign n48 = x5 ^ x1 ;
  assign n49 = n48 ^ x5 ;
  assign n47 = x5 ^ x2 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = n49 ^ x5 ;
  assign n52 = n50 & n51 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = n54 ^ n49 ;
  assign n56 = n46 & ~n55 ;
  assign n57 = n56 ^ n46 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n58 ^ x2 ;
  assign n60 = n59 ^ x5 ;
  assign n61 = n60 ^ x5 ;
  assign n64 = n46 ^ x2 ;
  assign n63 = x9 ^ x2 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = n63 ^ x2 ;
  assign n67 = n65 & n66 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = n68 ^ n63 ;
  assign n70 = x9 ^ x3 ;
  assign n71 = x1 & n70 ;
  assign n72 = n71 ^ n70 ;
  assign n73 = n69 & n72 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ x1 ;
  assign n76 = n75 ^ n70 ;
  assign n77 = n76 ^ x9 ;
  assign n131 = n61 & n77 ;
  assign n132 = n131 ^ n61 ;
  assign n129 = ~x7 & x8 ;
  assign n133 = ~x9 & n129 ;
  assign n134 = n132 & n133 ;
  assign n130 = n77 & n129 ;
  assign n135 = n134 ^ n130 ;
  assign n136 = n135 ^ x8 ;
  assign n137 = ~n128 & n136 ;
  assign n138 = n137 ^ n128 ;
  assign n139 = n138 ^ n136 ;
  assign n140 = n139 ^ n135 ;
  assign n141 = n140 ^ n45 ;
  assign n142 = n141 ^ x8 ;
  assign n78 = n77 ^ x9 ;
  assign n96 = n78 ^ n61 ;
  assign n98 = n96 ^ n61 ;
  assign n117 = n98 ^ n96 ;
  assign n118 = n117 ^ x7 ;
  assign n62 = n61 ^ x9 ;
  assign n89 = n77 ^ n62 ;
  assign n91 = n89 ^ n77 ;
  assign n103 = n98 ^ n91 ;
  assign n104 = n103 ^ x7 ;
  assign n105 = x9 & n104 ;
  assign n106 = n105 ^ x9 ;
  assign n107 = n106 ^ n104 ;
  assign n108 = n107 ^ n96 ;
  assign n111 = n91 ^ n89 ;
  assign n92 = n91 ^ x7 ;
  assign n93 = n91 & n92 ;
  assign n94 = n93 ^ n91 ;
  assign n95 = n94 ^ n92 ;
  assign n109 = n107 ^ n95 ;
  assign n110 = n109 ^ n96 ;
  assign n112 = n111 ^ n110 ;
  assign n113 = ~n108 & n112 ;
  assign n114 = n113 ^ n112 ;
  assign n90 = n89 ^ x7 ;
  assign n99 = n98 ^ x7 ;
  assign n97 = n96 ^ n95 ;
  assign n100 = n99 ^ n97 ;
  assign n101 = n90 & ~n100 ;
  assign n102 = n101 ^ n90 ;
  assign n115 = n114 ^ n102 ;
  assign n116 = n115 ^ n95 ;
  assign n119 = n118 ^ n116 ;
  assign n120 = n119 ^ x7 ;
  assign n121 = n120 ^ x7 ;
  assign n79 = n77 & n78 ;
  assign n80 = n79 ^ n77 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ n61 ;
  assign n83 = n62 & n82 ;
  assign n84 = n83 ^ n62 ;
  assign n85 = n84 ^ n82 ;
  assign n86 = n85 ^ n62 ;
  assign n87 = n86 ^ n80 ;
  assign n88 = n87 ^ n61 ;
  assign n122 = n121 ^ n88 ;
  assign n123 = ~n45 & n122 ;
  assign n124 = n123 ^ n45 ;
  assign n125 = n124 ^ n45 ;
  assign n126 = n125 ^ n45 ;
  assign n127 = n126 ^ n122 ;
  assign n143 = n142 ^ n127 ;
  assign n144 = n143 ^ x6 ;
  assign n156 = x0 & ~x2 ;
  assign n158 = x9 ^ x5 ;
  assign n159 = n158 ^ x9 ;
  assign n157 = x9 ^ x7 ;
  assign n160 = n159 ^ n157 ;
  assign n162 = n160 ^ x9 ;
  assign n164 = n162 ^ n160 ;
  assign n161 = n160 ^ n159 ;
  assign n165 = n161 ^ n160 ;
  assign n166 = n164 & n165 ;
  assign n167 = n166 ^ n165 ;
  assign n168 = n167 ^ n160 ;
  assign n170 = n158 ^ x1 ;
  assign n171 = n170 ^ n162 ;
  assign n169 = n167 ^ n161 ;
  assign n172 = n171 ^ n169 ;
  assign n173 = n168 & n172 ;
  assign n174 = n173 ^ n172 ;
  assign n175 = n174 ^ n167 ;
  assign n163 = n162 ^ n161 ;
  assign n176 = n175 ^ n163 ;
  assign n179 = n169 ^ n162 ;
  assign n180 = n170 ^ n161 ;
  assign n177 = n160 ^ x8 ;
  assign n181 = n180 ^ n177 ;
  assign n182 = n179 & n181 ;
  assign n183 = n182 ^ n181 ;
  assign n184 = n183 ^ n174 ;
  assign n185 = n184 ^ n167 ;
  assign n178 = n177 ^ n161 ;
  assign n186 = n185 ^ n178 ;
  assign n187 = n176 & n186 ;
  assign n188 = n187 ^ n176 ;
  assign n189 = n188 ^ n186 ;
  assign n190 = n189 ^ n174 ;
  assign n191 = n190 ^ n160 ;
  assign n192 = n191 ^ n158 ;
  assign n193 = n192 ^ x9 ;
  assign n194 = n193 ^ n170 ;
  assign n195 = n194 ^ n162 ;
  assign n196 = n195 ^ n161 ;
  assign n197 = n196 ^ n160 ;
  assign n198 = n156 & ~n197 ;
  assign n199 = n198 ^ n156 ;
  assign n200 = n199 ^ n156 ;
  assign n146 = x5 & x7 ;
  assign n147 = n146 ^ x7 ;
  assign n148 = x8 & n147 ;
  assign n149 = x0 & x1 ;
  assign n150 = n149 ^ x0 ;
  assign n151 = n150 ^ x1 ;
  assign n152 = x2 & x9 ;
  assign n153 = n152 ^ x2 ;
  assign n154 = ~n151 & n153 ;
  assign n155 = n148 & n154 ;
  assign n211 = ~x3 & ~x6 ;
  assign n212 = n155 & n211 ;
  assign n213 = n212 ^ n211 ;
  assign n214 = n200 & n213 ;
  assign n215 = n214 ^ n213 ;
  assign n210 = x3 & ~x6 ;
  assign n216 = n215 ^ n210 ;
  assign n217 = n216 ^ n143 ;
  assign n218 = n144 & n217 ;
  assign n219 = n218 ^ n217 ;
  assign n220 = n219 ^ n216 ;
  assign n201 = n200 ^ n155 ;
  assign n202 = x3 & x8 ;
  assign n203 = n147 & n202 ;
  assign n204 = n154 & n203 ;
  assign n205 = n204 ^ x3 ;
  assign n206 = n205 ^ n200 ;
  assign n207 = n201 & ~n206 ;
  assign n208 = n207 ^ n204 ;
  assign n209 = n208 ^ n200 ;
  assign n221 = n220 ^ n209 ;
  assign n145 = x6 & n144 ;
  assign n222 = n221 ^ n145 ;
  assign n223 = n222 ^ n209 ;
  assign n368 = n365 ^ n223 ;
  assign n370 = n365 ^ x7 ;
  assign n371 = n368 & n370 ;
  assign n372 = n371 ^ n368 ;
  assign n373 = n372 ^ x7 ;
  assign n230 = x1 & ~x3 ;
  assign n233 = ~x2 & x9 ;
  assign n234 = n230 & n233 ;
  assign n231 = ~x0 & ~x2 ;
  assign n232 = n230 & n231 ;
  assign n235 = n234 ^ n232 ;
  assign n227 = x2 & n30 ;
  assign n228 = n227 ^ x2 ;
  assign n229 = n228 ^ n30 ;
  assign n236 = n235 ^ n229 ;
  assign n237 = x2 & x6 ;
  assign n238 = n237 ^ x2 ;
  assign n239 = n238 ^ x6 ;
  assign n240 = n30 & ~n239 ;
  assign n241 = n240 ^ n239 ;
  assign n242 = n241 ^ x6 ;
  assign n243 = x5 & ~n242 ;
  assign n244 = n243 ^ x5 ;
  assign n245 = n244 ^ x5 ;
  assign n246 = n236 & n245 ;
  assign n247 = n246 ^ n245 ;
  assign n248 = n247 ^ n245 ;
  assign n249 = x1 & x2 ;
  assign n250 = n249 ^ x1 ;
  assign n251 = n250 ^ x2 ;
  assign n252 = x9 & ~n251 ;
  assign n253 = n252 ^ n251 ;
  assign n254 = n253 ^ n63 ;
  assign n255 = ~x0 & ~x3 ;
  assign n256 = x6 & x8 ;
  assign n257 = n255 & n256 ;
  assign n258 = n254 & n257 ;
  assign n259 = n258 ^ x8 ;
  assign n260 = n248 & n259 ;
  assign n261 = n260 ^ n259 ;
  assign n262 = n261 ^ x8 ;
  assign n276 = x1 & ~x8 ;
  assign n263 = x2 & x3 ;
  assign n264 = n263 ^ x2 ;
  assign n275 = n16 & n264 ;
  assign n277 = n276 ^ n275 ;
  assign n278 = x0 & n277 ;
  assign n279 = n278 ^ n277 ;
  assign n280 = n237 ^ x6 ;
  assign n281 = x3 & n280 ;
  assign n282 = n281 ^ x3 ;
  assign n269 = n26 ^ x9 ;
  assign n287 = x8 & ~n269 ;
  assign n288 = n282 & n287 ;
  assign n289 = n288 ^ n287 ;
  assign n286 = x8 & ~n152 ;
  assign n290 = n289 ^ n286 ;
  assign n291 = n290 ^ x8 ;
  assign n283 = ~n269 & n282 ;
  assign n284 = n283 ^ n269 ;
  assign n285 = n284 ^ n152 ;
  assign n292 = n291 ^ n285 ;
  assign n293 = n279 & ~n292 ;
  assign n294 = n293 ^ n279 ;
  assign n295 = n294 ^ n292 ;
  assign n265 = n264 ^ x3 ;
  assign n266 = x0 & n265 ;
  assign n267 = n266 ^ x0 ;
  assign n268 = n267 ^ n265 ;
  assign n296 = ~x8 & ~x9 ;
  assign n297 = ~x1 & ~x5 ;
  assign n298 = n296 & n297 ;
  assign n299 = ~n268 & n298 ;
  assign n300 = n299 ^ x5 ;
  assign n301 = ~n295 & ~n300 ;
  assign n270 = x8 & n269 ;
  assign n271 = n270 ^ x8 ;
  assign n272 = n271 ^ n269 ;
  assign n273 = ~n268 & n272 ;
  assign n274 = n273 ^ n268 ;
  assign n302 = n301 ^ n274 ;
  assign n303 = n262 & ~n302 ;
  assign n304 = n303 ^ n262 ;
  assign n305 = n304 ^ n302 ;
  assign n309 = n16 & ~n308 ;
  assign n310 = ~x5 & x6 ;
  assign n311 = ~n309 & n310 ;
  assign n312 = n311 ^ x6 ;
  assign n313 = x1 & x5 ;
  assign n314 = x9 ^ x0 ;
  assign n315 = x2 & ~n314 ;
  assign n316 = n313 & n315 ;
  assign n317 = x8 & ~n316 ;
  assign n318 = ~n312 & n317 ;
  assign n319 = n318 ^ x8 ;
  assign n322 = x8 & x9 ;
  assign n323 = n322 ^ x9 ;
  assign n324 = ~n151 & n323 ;
  assign n325 = n324 ^ n276 ;
  assign n320 = x0 & ~x1 ;
  assign n321 = n153 & n320 ;
  assign n326 = n325 ^ n321 ;
  assign n327 = ~x5 & n326 ;
  assign n328 = x3 & ~n327 ;
  assign n329 = ~n319 & n328 ;
  assign n330 = n329 ^ x3 ;
  assign n336 = ~n305 & n330 ;
  assign n337 = n336 ^ n330 ;
  assign n338 = n337 ^ n305 ;
  assign n374 = n373 ^ n338 ;
  assign n380 = n373 ^ n223 ;
  assign n366 = n365 ^ x4 ;
  assign n381 = n380 ^ n366 ;
  assign n382 = ~n374 & n381 ;
  assign n383 = n382 ^ n381 ;
  assign n392 = n383 ^ n372 ;
  assign n369 = n368 ^ x4 ;
  assign n375 = n374 ^ n369 ;
  assign n376 = n338 ^ n223 ;
  assign n377 = n376 ^ n373 ;
  assign n378 = ~n375 & ~n377 ;
  assign n379 = n378 ^ n375 ;
  assign n384 = n383 ^ n379 ;
  assign n385 = n384 ^ n373 ;
  assign n386 = n385 ^ n369 ;
  assign n387 = n383 ^ n338 ;
  assign n388 = n387 ^ x4 ;
  assign n389 = ~n386 & ~n388 ;
  assign n390 = n389 ^ n386 ;
  assign n391 = n390 ^ n379 ;
  assign n393 = n392 ^ n391 ;
  assign n344 = n223 ^ x7 ;
  assign n367 = n366 ^ n344 ;
  assign n394 = n393 ^ n367 ;
  assign n331 = x7 & ~n330 ;
  assign n332 = n305 & n331 ;
  assign n333 = n332 ^ x7 ;
  assign n334 = n333 ^ x7 ;
  assign n335 = n334 ^ x7 ;
  assign n339 = n338 ^ n335 ;
  assign n340 = ~x4 & n223 ;
  assign n341 = ~n339 & n340 ;
  assign n224 = x4 & ~n223 ;
  assign n225 = n224 ^ x4 ;
  assign n226 = n225 ^ n223 ;
  assign n342 = n341 ^ n226 ;
  assign n343 = n342 ^ x4 ;
  assign n395 = n394 ^ n343 ;
  assign n396 = n395 ^ n365 ;
  assign n415 = x2 & x8 ;
  assign n427 = n415 ^ x2 ;
  assign n428 = n427 ^ x8 ;
  assign n429 = x5 & n428 ;
  assign n430 = n429 ^ x5 ;
  assign n431 = x5 ^ x3 ;
  assign n432 = x8 & n431 ;
  assign n433 = n432 ^ n431 ;
  assign n434 = n433 ^ x5 ;
  assign n435 = x0 & n434 ;
  assign n436 = n430 & n435 ;
  assign n437 = n436 ^ n430 ;
  assign n438 = n437 ^ n435 ;
  assign n416 = n415 ^ x8 ;
  assign n417 = n416 ^ x0 ;
  assign n418 = x5 ^ x0 ;
  assign n419 = n418 ^ x0 ;
  assign n420 = n418 & n419 ;
  assign n421 = n420 ^ n418 ;
  assign n422 = n421 ^ n416 ;
  assign n423 = n417 & n422 ;
  assign n424 = n423 ^ n420 ;
  assign n425 = n424 ^ n416 ;
  assign n439 = n438 ^ n425 ;
  assign n440 = n439 ^ n425 ;
  assign n426 = n425 ^ x1 ;
  assign n441 = n440 ^ n426 ;
  assign n442 = n440 ^ n425 ;
  assign n443 = ~n441 & ~n442 ;
  assign n444 = n443 ^ n441 ;
  assign n445 = n444 ^ n440 ;
  assign n446 = ~n202 & n231 ;
  assign n447 = n446 ^ x0 ;
  assign n448 = ~x6 & n447 ;
  assign n449 = n445 & n448 ;
  assign n450 = n449 ^ x6 ;
  assign n451 = x8 ^ x2 ;
  assign n452 = n451 ^ x8 ;
  assign n453 = n452 ^ x1 ;
  assign n455 = n453 ^ x8 ;
  assign n465 = n455 ^ n453 ;
  assign n454 = n453 ^ n452 ;
  assign n456 = n455 ^ n454 ;
  assign n457 = n454 ^ x6 ;
  assign n458 = n456 ^ x3 ;
  assign n459 = n457 & n458 ;
  assign n460 = n459 ^ x6 ;
  assign n461 = n460 ^ n456 ;
  assign n462 = n456 & ~n461 ;
  assign n463 = n462 ^ n459 ;
  assign n464 = n463 ^ x6 ;
  assign n466 = n465 ^ n464 ;
  assign n467 = n454 ^ n453 ;
  assign n469 = n454 ^ x3 ;
  assign n468 = n455 ^ x6 ;
  assign n470 = n469 ^ n468 ;
  assign n471 = ~n467 & ~n470 ;
  assign n472 = n471 ^ n462 ;
  assign n473 = n472 ^ n459 ;
  assign n474 = n466 & n473 ;
  assign n478 = ~x5 & ~x9 ;
  assign n485 = n474 & n478 ;
  assign n475 = x0 & x8 ;
  assign n476 = n475 ^ x8 ;
  assign n477 = ~x2 & ~n476 ;
  assign n480 = ~x1 & x6 ;
  assign n479 = ~x0 & x1 ;
  assign n481 = n480 ^ n479 ;
  assign n482 = n478 & n481 ;
  assign n483 = n477 & n482 ;
  assign n484 = ~n474 & n483 ;
  assign n486 = n485 ^ n484 ;
  assign n487 = n486 ^ x9 ;
  assign n488 = n450 & n487 ;
  assign n489 = n488 ^ n450 ;
  assign n490 = n489 ^ n487 ;
  assign n491 = n490 ^ n487 ;
  assign n505 = x3 & n249 ;
  assign n506 = x5 & x8 ;
  assign n507 = n506 ^ x5 ;
  assign n508 = x9 & n507 ;
  assign n509 = n505 & n508 ;
  assign n510 = n509 ^ x9 ;
  assign n492 = n360 ^ x3 ;
  assign n493 = ~n428 & n492 ;
  assign n494 = x0 & ~n313 ;
  assign n495 = ~n493 & n494 ;
  assign n496 = n495 ^ x0 ;
  assign n499 = ~x5 & n264 ;
  assign n497 = x3 & ~x5 ;
  assign n498 = ~n249 & n497 ;
  assign n500 = n499 ^ n498 ;
  assign n501 = n500 ^ n265 ;
  assign n502 = x6 & ~n501 ;
  assign n503 = ~n496 & n502 ;
  assign n504 = n503 ^ x6 ;
  assign n511 = n510 ^ n504 ;
  assign n513 = n354 & n507 ;
  assign n514 = n505 & n513 ;
  assign n512 = x4 & ~x9 ;
  assign n515 = n514 ^ n512 ;
  assign n516 = n515 ^ x4 ;
  assign n517 = n516 ^ n504 ;
  assign n518 = ~n511 & ~n517 ;
  assign n519 = n518 ^ n515 ;
  assign n520 = n519 ^ n504 ;
  assign n521 = ~n491 & n520 ;
  assign n522 = n521 ^ n520 ;
  assign n523 = n522 ^ n520 ;
  assign n397 = ~x6 & ~n19 ;
  assign n398 = ~x4 & n397 ;
  assign n699 = ~x7 & n154 ;
  assign n700 = n398 & n699 ;
  assign n701 = n700 ^ x7 ;
  assign n702 = n701 ^ x7 ;
  assign n713 = ~n523 & ~n702 ;
  assign n712 = x7 & ~n702 ;
  assign n714 = n713 ^ n712 ;
  assign n575 = ~x2 & ~n151 ;
  assign n576 = x5 ^ x4 ;
  assign n577 = x8 & n576 ;
  assign n578 = n577 ^ x5 ;
  assign n579 = ~n349 & ~n578 ;
  assign n580 = n579 ^ n349 ;
  assign n581 = x4 & n347 ;
  assign n582 = ~n580 & n581 ;
  assign n583 = n582 ^ n580 ;
  assign n584 = n583 ^ n581 ;
  assign n585 = n575 & n584 ;
  assign n586 = n585 ^ n575 ;
  assign n527 = x6 ^ x5 ;
  assign n525 = n314 ^ x9 ;
  assign n544 = n527 ^ n525 ;
  assign n540 = n527 ^ x9 ;
  assign n541 = ~n527 & ~n540 ;
  assign n526 = x9 ^ x6 ;
  assign n528 = n527 ^ n526 ;
  assign n529 = n528 ^ x8 ;
  assign n530 = n529 ^ x8 ;
  assign n531 = n530 ^ n314 ;
  assign n532 = n531 ^ n525 ;
  assign n533 = n529 & n532 ;
  assign n534 = n533 ^ n529 ;
  assign n535 = n534 ^ n525 ;
  assign n536 = n535 ^ n529 ;
  assign n537 = n525 & n536 ;
  assign n538 = n537 ^ n525 ;
  assign n539 = n538 ^ n536 ;
  assign n542 = n541 ^ n539 ;
  assign n543 = n542 ^ n534 ;
  assign n545 = n544 ^ n543 ;
  assign n547 = n531 ^ n529 ;
  assign n546 = n539 ^ n525 ;
  assign n548 = n547 ^ n546 ;
  assign n549 = n545 & n548 ;
  assign n550 = n549 ^ n545 ;
  assign n551 = n550 ^ n548 ;
  assign n552 = n551 ^ n545 ;
  assign n553 = n552 ^ n539 ;
  assign n554 = n553 ^ n535 ;
  assign n555 = n554 ^ x5 ;
  assign n556 = n555 ^ x9 ;
  assign n557 = n556 ^ x9 ;
  assign n558 = x9 ^ x8 ;
  assign n559 = x5 & n558 ;
  assign n560 = n559 ^ x5 ;
  assign n561 = n63 & n314 ;
  assign n562 = n561 ^ n314 ;
  assign n563 = n562 ^ n63 ;
  assign n564 = n560 & n563 ;
  assign n565 = n564 ^ n560 ;
  assign n566 = x2 & n565 ;
  assign n567 = n566 ^ x2 ;
  assign n568 = ~n557 & n567 ;
  assign n569 = n568 ^ n565 ;
  assign n570 = n153 & n345 ;
  assign n571 = ~x1 & ~n570 ;
  assign n572 = n569 & n571 ;
  assign n573 = n572 ^ n570 ;
  assign n589 = n586 ^ n573 ;
  assign n646 = n586 ^ x1 ;
  assign n647 = n589 & n646 ;
  assign n648 = n647 ^ n589 ;
  assign n649 = n648 ^ x1 ;
  assign n593 = n526 ^ n158 ;
  assign n594 = n593 ^ x8 ;
  assign n595 = n594 ^ x9 ;
  assign n596 = n595 ^ n558 ;
  assign n592 = n558 ^ n526 ;
  assign n597 = n596 ^ n592 ;
  assign n591 = x8 ^ x0 ;
  assign n598 = n597 ^ n591 ;
  assign n599 = n598 ^ n597 ;
  assign n600 = n598 ^ n592 ;
  assign n601 = n599 & n600 ;
  assign n602 = n601 ^ n598 ;
  assign n605 = n598 ^ n558 ;
  assign n606 = n605 ^ n600 ;
  assign n607 = n606 ^ n599 ;
  assign n608 = n598 ^ x9 ;
  assign n609 = n608 ^ n600 ;
  assign n610 = n609 ^ n599 ;
  assign n611 = n607 & n610 ;
  assign n603 = n600 ^ n599 ;
  assign n604 = n603 ^ n598 ;
  assign n612 = n611 ^ n604 ;
  assign n613 = n602 & n612 ;
  assign n614 = n613 ^ n598 ;
  assign n615 = n614 ^ n598 ;
  assign n616 = x2 & ~n615 ;
  assign n617 = n616 ^ x2 ;
  assign n618 = n617 ^ n615 ;
  assign n619 = x0 & x6 ;
  assign n620 = n619 ^ x6 ;
  assign n621 = x2 & n620 ;
  assign n622 = n621 ^ x2 ;
  assign n623 = n622 ^ n620 ;
  assign n624 = ~x6 & ~x8 ;
  assign n625 = n506 ^ x8 ;
  assign n626 = ~n624 & n625 ;
  assign n627 = n623 & n626 ;
  assign n628 = n627 ^ n624 ;
  assign n629 = x9 & ~n628 ;
  assign n630 = n629 ^ x9 ;
  assign n631 = n630 ^ n628 ;
  assign n632 = n618 & n631 ;
  assign n633 = n632 ^ n618 ;
  assign n634 = n633 ^ n631 ;
  assign n650 = n649 ^ n634 ;
  assign n651 = n649 ^ n573 ;
  assign n587 = n586 ^ x4 ;
  assign n652 = n651 ^ n587 ;
  assign n653 = n650 & n652 ;
  assign n654 = n653 ^ n652 ;
  assign n655 = n654 ^ n650 ;
  assign n656 = n655 ^ n652 ;
  assign n666 = n656 ^ n648 ;
  assign n641 = ~x1 & x4 ;
  assign n642 = n586 & n641 ;
  assign n643 = n573 & n642 ;
  assign n638 = x1 & ~x4 ;
  assign n639 = ~n586 & n638 ;
  assign n640 = ~n573 & n639 ;
  assign n644 = n643 ^ n640 ;
  assign n636 = ~n586 & ~n634 ;
  assign n635 = x4 & ~n634 ;
  assign n637 = n636 ^ n635 ;
  assign n645 = n644 ^ n637 ;
  assign n657 = n656 ^ n645 ;
  assign n658 = n657 ^ n649 ;
  assign n590 = n589 ^ x4 ;
  assign n659 = n658 ^ n590 ;
  assign n660 = n656 ^ n634 ;
  assign n661 = n660 ^ x4 ;
  assign n662 = n659 & n661 ;
  assign n663 = n662 ^ n659 ;
  assign n664 = n663 ^ n661 ;
  assign n665 = n664 ^ n645 ;
  assign n667 = n666 ^ n665 ;
  assign n574 = n573 ^ x1 ;
  assign n588 = n587 ^ n574 ;
  assign n668 = n667 ^ n588 ;
  assign n669 = n668 ^ n586 ;
  assign n670 = n520 ^ n491 ;
  assign n703 = ~x3 & ~n702 ;
  assign n704 = n703 ^ n520 ;
  assign n705 = ~n703 & ~n704 ;
  assign n706 = n705 ^ n703 ;
  assign n707 = n706 ^ n491 ;
  assign n708 = ~n670 & n707 ;
  assign n709 = n708 ^ n705 ;
  assign n710 = n709 ^ n491 ;
  assign n711 = n669 & n710 ;
  assign n715 = n714 ^ n711 ;
  assign n716 = n715 ^ n701 ;
  assign n686 = n669 ^ x3 ;
  assign n687 = ~x3 & n520 ;
  assign n688 = ~n491 & n687 ;
  assign n689 = n688 ^ x3 ;
  assign n690 = n689 ^ x3 ;
  assign n691 = n686 & n690 ;
  assign n692 = n691 ^ n686 ;
  assign n693 = n692 ^ n690 ;
  assign n694 = n693 ^ n689 ;
  assign n695 = n694 ^ n669 ;
  assign n682 = x3 & n669 ;
  assign n683 = n682 ^ x3 ;
  assign n684 = n683 ^ x3 ;
  assign n685 = n684 ^ n669 ;
  assign n696 = n695 ^ n685 ;
  assign n697 = n696 ^ n523 ;
  assign n717 = n716 ^ n697 ;
  assign n671 = ~x3 & x7 ;
  assign n672 = n671 ^ n520 ;
  assign n673 = ~n671 & ~n672 ;
  assign n674 = n673 ^ n671 ;
  assign n675 = n674 ^ n491 ;
  assign n676 = ~n670 & n675 ;
  assign n677 = n676 ^ n673 ;
  assign n678 = n677 ^ n491 ;
  assign n679 = n669 & n678 ;
  assign n524 = x7 & ~n523 ;
  assign n680 = n679 ^ n524 ;
  assign n681 = n680 ^ x7 ;
  assign n698 = n697 ^ n681 ;
  assign n718 = n717 ^ n698 ;
  assign n407 = n156 & n296 ;
  assign n405 = x2 & ~x8 ;
  assign n406 = ~n151 & n405 ;
  assign n408 = n407 ^ n406 ;
  assign n402 = ~x2 & n149 ;
  assign n403 = n323 & n402 ;
  assign n399 = x8 & ~x9 ;
  assign n400 = x1 & ~x2 ;
  assign n401 = n399 & n400 ;
  assign n404 = n403 ^ n401 ;
  assign n409 = n408 ^ n404 ;
  assign n412 = ~n154 & ~n409 ;
  assign n410 = ~x7 & ~n154 ;
  assign n411 = n409 & n410 ;
  assign n413 = n412 ^ n411 ;
  assign n414 = n398 & ~n413 ;
  assign n719 = n718 ^ n414 ;
  assign n720 = x2 & ~n345 ;
  assign n721 = x1 & ~n720 ;
  assign n722 = ~x2 & ~n202 ;
  assign n723 = x5 & ~n722 ;
  assign n724 = ~n721 & n723 ;
  assign n725 = x3 & ~x8 ;
  assign n726 = ~n26 & ~n725 ;
  assign n727 = x3 & ~x9 ;
  assign n728 = ~x6 & ~n727 ;
  assign n729 = ~n726 & n728 ;
  assign n730 = ~x3 & x9 ;
  assign n731 = x1 & n730 ;
  assign n732 = x6 & ~x8 ;
  assign n733 = ~x4 & n732 ;
  assign n734 = n731 & n733 ;
  assign n735 = n734 ^ x4 ;
  assign n736 = ~n729 & ~n735 ;
  assign n737 = ~n724 & n736 ;
  assign n745 = ~x1 & ~x8 ;
  assign n746 = ~x9 & n745 ;
  assign n747 = ~x3 & n310 ;
  assign n748 = n746 & n747 ;
  assign n738 = x1 & ~x9 ;
  assign n740 = ~x2 & x3 ;
  assign n741 = x8 & n740 ;
  assign n739 = ~x5 & ~x8 ;
  assign n742 = n741 ^ n739 ;
  assign n743 = n742 ^ n17 ;
  assign n744 = n738 & ~n743 ;
  assign n749 = n748 ^ n744 ;
  assign n751 = x1 & x8 ;
  assign n753 = ~x9 & n751 ;
  assign n752 = ~n349 & ~n751 ;
  assign n754 = n753 ^ n752 ;
  assign n756 = ~x2 & ~x8 ;
  assign n757 = n16 & n756 ;
  assign n758 = ~n754 & n757 ;
  assign n755 = ~x2 & ~n754 ;
  assign n759 = n758 ^ n755 ;
  assign n750 = ~x8 & n16 ;
  assign n760 = n759 ^ n750 ;
  assign n761 = x3 & n760 ;
  assign n762 = ~n749 & ~n761 ;
  assign n763 = n737 & n762 ;
  assign n764 = ~n322 & ~n732 ;
  assign n765 = ~x5 & ~n764 ;
  assign n766 = x2 & ~n362 ;
  assign n767 = n766 ^ n362 ;
  assign n768 = ~n765 & ~n767 ;
  assign n769 = x4 & ~n768 ;
  assign n770 = ~x0 & ~n769 ;
  assign n771 = ~n763 & n770 ;
  assign n809 = x9 ^ x1 ;
  assign n826 = n809 ^ x9 ;
  assign n828 = n826 ^ n526 ;
  assign n825 = n558 ^ x9 ;
  assign n827 = n826 ^ n825 ;
  assign n829 = n828 ^ n827 ;
  assign n850 = n829 ^ x2 ;
  assign n832 = n826 ^ x9 ;
  assign n833 = n832 ^ x2 ;
  assign n830 = n827 & n829 ;
  assign n831 = n830 ^ n827 ;
  assign n834 = n833 ^ n831 ;
  assign n841 = x2 & ~n834 ;
  assign n848 = n841 ^ n830 ;
  assign n842 = n841 ^ n828 ;
  assign n843 = n842 ^ x2 ;
  assign n844 = n830 ^ n826 ;
  assign n845 = n844 ^ n829 ;
  assign n846 = n843 & ~n845 ;
  assign n838 = x2 & ~n826 ;
  assign n837 = n526 & ~n826 ;
  assign n839 = n838 ^ n837 ;
  assign n835 = x2 & ~n526 ;
  assign n836 = n834 & n835 ;
  assign n840 = n839 ^ n836 ;
  assign n847 = n846 ^ n840 ;
  assign n849 = n848 ^ n847 ;
  assign n851 = n850 ^ n849 ;
  assign n852 = n851 ^ x2 ;
  assign n853 = n852 ^ n558 ;
  assign n854 = n853 ^ x9 ;
  assign n822 = x0 & ~x5 ;
  assign n859 = x3 & n822 ;
  assign n860 = n854 & n859 ;
  assign n861 = n860 ^ n822 ;
  assign n810 = n809 ^ x8 ;
  assign n811 = n526 ^ x9 ;
  assign n804 = x6 ^ x3 ;
  assign n805 = n804 ^ x9 ;
  assign n806 = n805 ^ x9 ;
  assign n807 = n806 ^ n526 ;
  assign n812 = n811 ^ n807 ;
  assign n813 = ~x8 & n812 ;
  assign n814 = n813 ^ n526 ;
  assign n815 = ~n810 & n814 ;
  assign n816 = n815 ^ n813 ;
  assign n808 = ~x8 & n807 ;
  assign n817 = n816 ^ n808 ;
  assign n818 = n817 ^ n809 ;
  assign n819 = n818 ^ x8 ;
  assign n820 = n819 ^ x9 ;
  assign n821 = n820 ^ n526 ;
  assign n855 = n740 & n822 ;
  assign n856 = ~n821 & n855 ;
  assign n857 = n854 & n856 ;
  assign n823 = ~x2 & n822 ;
  assign n824 = ~n821 & n823 ;
  assign n858 = n857 ^ n824 ;
  assign n862 = n861 ^ n858 ;
  assign n863 = n862 ^ n822 ;
  assign n868 = ~x4 & ~x7 ;
  assign n869 = n863 & n868 ;
  assign n870 = n869 ^ x7 ;
  assign n776 = x5 & x9 ;
  assign n777 = n475 & n776 ;
  assign n772 = n322 ^ x8 ;
  assign n773 = n772 ^ x9 ;
  assign n774 = x5 & ~n773 ;
  assign n775 = n774 ^ x5 ;
  assign n778 = n777 ^ n775 ;
  assign n779 = x1 & ~x5 ;
  assign n780 = ~n152 & n779 ;
  assign n781 = n780 ^ x1 ;
  assign n782 = n778 & n781 ;
  assign n783 = n782 ^ n781 ;
  assign n784 = x2 & ~n558 ;
  assign n785 = n269 & n784 ;
  assign n786 = n785 ^ x2 ;
  assign n787 = ~x3 & ~n786 ;
  assign n788 = ~n783 & n787 ;
  assign n789 = n788 ^ x3 ;
  assign n790 = x5 & ~n492 ;
  assign n791 = ~x2 & ~n773 ;
  assign n792 = ~n790 & n791 ;
  assign n794 = x9 & ~n265 ;
  assign n795 = n794 ^ x9 ;
  assign n796 = n751 ^ x8 ;
  assign n797 = x0 & n796 ;
  assign n798 = n795 & n797 ;
  assign n799 = ~n792 & n798 ;
  assign n793 = x0 & n792 ;
  assign n800 = n799 ^ n793 ;
  assign n801 = ~n789 & n800 ;
  assign n802 = n801 ^ n789 ;
  assign n803 = n802 ^ n800 ;
  assign n864 = ~x4 & ~x6 ;
  assign n865 = ~x7 & n864 ;
  assign n866 = ~n863 & n865 ;
  assign n867 = ~n803 & n866 ;
  assign n871 = n870 ^ n867 ;
  assign n874 = x7 & n322 ;
  assign n875 = x0 & ~n874 ;
  assign n876 = n14 & ~n875 ;
  assign n877 = n751 ^ x1 ;
  assign n878 = n877 ^ x8 ;
  assign n879 = n30 & ~n878 ;
  assign n880 = ~n876 & ~n879 ;
  assign n881 = ~x5 & ~x6 ;
  assign n882 = ~x4 & ~n265 ;
  assign n883 = n881 & n882 ;
  assign n884 = ~n880 & n883 ;
  assign n886 = ~n871 & n884 ;
  assign n887 = ~n771 & n886 ;
  assign n885 = ~x7 & n884 ;
  assign n888 = n887 ^ n885 ;
  assign n872 = ~n771 & ~n871 ;
  assign n873 = n872 ^ x7 ;
  assign n889 = n888 ^ n873 ;
  assign n890 = n889 ^ n884 ;
  assign n893 = ~x3 & ~x5 ;
  assign n894 = x6 & n893 ;
  assign n891 = ~x1 & ~x6 ;
  assign n892 = n430 & n891 ;
  assign n895 = n894 ^ n892 ;
  assign n928 = n738 & n895 ;
  assign n897 = ~x3 & x5 ;
  assign n898 = n323 & n897 ;
  assign n899 = n898 ^ x3 ;
  assign n900 = x2 & ~n899 ;
  assign n901 = n900 ^ x2 ;
  assign n902 = n901 ^ n899 ;
  assign n904 = n17 & n624 ;
  assign n905 = n904 ^ x6 ;
  assign n903 = x6 & n497 ;
  assign n906 = n905 ^ n903 ;
  assign n907 = n902 & n906 ;
  assign n908 = n907 ^ n902 ;
  assign n909 = n908 ^ n906 ;
  assign n910 = n47 ^ x5 ;
  assign n911 = n431 ^ n47 ;
  assign n912 = n910 & n911 ;
  assign n913 = n912 ^ n47 ;
  assign n918 = ~x8 & n913 ;
  assign n919 = n918 ^ x2 ;
  assign n920 = n919 ^ x5 ;
  assign n925 = n738 & ~n920 ;
  assign n926 = n895 & n925 ;
  assign n927 = ~n909 & n926 ;
  assign n929 = n928 ^ n927 ;
  assign n915 = n776 ^ n233 ;
  assign n914 = n323 & n913 ;
  assign n916 = n915 ^ n914 ;
  assign n917 = n916 ^ x9 ;
  assign n921 = n920 ^ n917 ;
  assign n922 = x1 & ~n921 ;
  assign n923 = ~n909 & n922 ;
  assign n924 = n923 ^ x1 ;
  assign n930 = n929 ^ n924 ;
  assign n896 = ~x9 & n895 ;
  assign n931 = n930 ^ n896 ;
  assign n932 = x0 & ~n931 ;
  assign n933 = n932 ^ x0 ;
  assign n934 = n776 ^ x5 ;
  assign n935 = n934 ^ x9 ;
  assign n936 = ~n624 & n935 ;
  assign n937 = ~x2 & ~n936 ;
  assign n940 = ~x6 & x9 ;
  assign n941 = n779 & n940 ;
  assign n938 = x5 & ~x6 ;
  assign n939 = n399 & n938 ;
  assign n942 = n941 ^ n939 ;
  assign n943 = x3 & ~n942 ;
  assign n944 = ~n937 & n943 ;
  assign n945 = n944 ^ x3 ;
  assign n954 = x3 & x6 ;
  assign n955 = n954 ^ x3 ;
  assign n960 = ~n310 & ~n955 ;
  assign n961 = n296 & n960 ;
  assign n962 = n961 ^ n399 ;
  assign n950 = ~x2 & ~x3 ;
  assign n951 = n310 & n950 ;
  assign n949 = ~x6 & n263 ;
  assign n952 = n951 ^ n949 ;
  assign n953 = n952 ^ n310 ;
  assign n958 = x9 & ~n953 ;
  assign n956 = n323 & n955 ;
  assign n957 = ~n953 & n956 ;
  assign n959 = n958 ^ n957 ;
  assign n963 = n962 ^ n959 ;
  assign n964 = ~x1 & ~n963 ;
  assign n965 = ~n945 & n964 ;
  assign n966 = n965 ^ n945 ;
  assign n946 = ~x9 & n310 ;
  assign n947 = n751 & n946 ;
  assign n948 = ~n945 & n947 ;
  assign n967 = n966 ^ n948 ;
  assign n970 = x4 & ~n967 ;
  assign n971 = ~n933 & n970 ;
  assign n972 = n971 ^ x4 ;
  assign n968 = n933 & ~n967 ;
  assign n969 = n968 ^ n967 ;
  assign n973 = n972 ^ n969 ;
  assign n982 = n526 ^ x2 ;
  assign n983 = n159 ^ x2 ;
  assign n984 = n982 & ~n983 ;
  assign n985 = ~n558 & n984 ;
  assign n994 = n985 ^ n984 ;
  assign n979 = n558 ^ n158 ;
  assign n980 = n979 ^ x2 ;
  assign n981 = n979 & n980 ;
  assign n986 = n985 ^ n981 ;
  assign n987 = n986 ^ n984 ;
  assign n988 = n987 ^ n980 ;
  assign n990 = n158 ^ x2 ;
  assign n989 = n984 ^ n981 ;
  assign n991 = n990 ^ n989 ;
  assign n992 = n988 & ~n991 ;
  assign n993 = n992 ^ n981 ;
  assign n995 = n994 ^ n993 ;
  assign n996 = n995 ^ n980 ;
  assign n998 = n17 & n345 ;
  assign n999 = n998 ^ n497 ;
  assign n997 = n732 & n893 ;
  assign n1000 = n999 ^ n997 ;
  assign n1009 = ~x1 & ~n1000 ;
  assign n1010 = ~n996 & n1009 ;
  assign n1004 = x6 & n265 ;
  assign n1005 = ~n727 & ~n1004 ;
  assign n1008 = ~x1 & n1005 ;
  assign n1011 = n1010 ^ n1008 ;
  assign n1001 = n996 & n1000 ;
  assign n1002 = n1001 ^ n996 ;
  assign n1003 = n1002 ^ n1000 ;
  assign n1006 = n1005 ^ n1003 ;
  assign n1007 = n1006 ^ n1005 ;
  assign n1012 = n1011 ^ n1007 ;
  assign n974 = ~x5 & ~n322 ;
  assign n975 = ~x3 & x4 ;
  assign n976 = ~n251 & n975 ;
  assign n977 = ~n974 & n976 ;
  assign n1013 = x2 & n310 ;
  assign n1017 = ~x4 & ~n527 ;
  assign n1019 = ~n1013 & n1017 ;
  assign n1020 = n977 & n1019 ;
  assign n1021 = ~n1012 & n1020 ;
  assign n1018 = n977 & n1017 ;
  assign n1022 = n1021 ^ n1018 ;
  assign n1014 = ~x4 & ~n1013 ;
  assign n1015 = ~n1012 & n1014 ;
  assign n1016 = n1015 ^ x4 ;
  assign n1023 = n1022 ^ n1016 ;
  assign n978 = ~n527 & n977 ;
  assign n1024 = n1023 ^ n978 ;
  assign n1025 = ~x0 & ~x7 ;
  assign n1026 = ~n1024 & n1025 ;
  assign n1027 = n1026 ^ x7 ;
  assign n1028 = ~n973 & ~n1027 ;
  assign n1029 = n1028 ^ x7 ;
  assign n1030 = x2 & n151 ;
  assign n1031 = ~x4 & n1030 ;
  assign n1032 = x4 ^ x3 ;
  assign n1033 = n575 & n1032 ;
  assign n1034 = ~n1031 & ~n1033 ;
  assign n1035 = ~x7 & n356 ;
  assign n1036 = ~n1034 & n1035 ;
  assign n1037 = x3 & ~x4 ;
  assign n1038 = ~n575 & n1037 ;
  assign n1039 = n575 & n975 ;
  assign n1040 = ~n1038 & ~n1039 ;
  assign n1041 = n1035 & ~n1040 ;
  assign n1052 = n48 ^ x9 ;
  assign n1053 = n1052 ^ x5 ;
  assign n1054 = n1053 ^ n158 ;
  assign n1055 = ~n158 & n1054 ;
  assign n1045 = x6 & n982 ;
  assign n1046 = n1045 ^ x6 ;
  assign n1047 = n1046 ^ n982 ;
  assign n1048 = n1047 ^ x2 ;
  assign n1049 = n1048 ^ x6 ;
  assign n1050 = x2 & ~n1049 ;
  assign n1051 = n1050 ^ x2 ;
  assign n1056 = n1055 ^ n1051 ;
  assign n1057 = n1056 ^ n1047 ;
  assign n1058 = n1057 ^ n990 ;
  assign n1060 = n526 ^ x6 ;
  assign n1059 = n1051 ^ x2 ;
  assign n1061 = n1060 ^ n1059 ;
  assign n1062 = ~n1058 & n1061 ;
  assign n1063 = n1062 ^ n1061 ;
  assign n1064 = n1063 ^ n1051 ;
  assign n1065 = n1064 ^ n1048 ;
  assign n1066 = n1065 ^ x1 ;
  assign n1067 = n1066 ^ x5 ;
  assign n1068 = n1067 ^ x9 ;
  assign n1069 = n1068 ^ n1052 ;
  assign n1070 = n475 & ~n1069 ;
  assign n1042 = n306 ^ x2 ;
  assign n1043 = x8 & n935 ;
  assign n1044 = n1042 & n1043 ;
  assign n1071 = n1070 ^ n1044 ;
  assign n1072 = n1071 ^ x8 ;
  assign n1073 = n1072 ^ x8 ;
  assign n1090 = n1073 ^ x7 ;
  assign n1074 = n314 ^ x2 ;
  assign n1075 = x2 & ~n1074 ;
  assign n1077 = n1075 ^ n745 ;
  assign n1078 = n1074 ^ n46 ;
  assign n1079 = x5 & ~n1078 ;
  assign n1080 = n1077 & n1079 ;
  assign n1076 = x5 & ~n1075 ;
  assign n1081 = n1080 ^ n1076 ;
  assign n1082 = n1081 ^ x5 ;
  assign n1083 = x6 & ~n558 ;
  assign n1092 = x7 & ~n451 ;
  assign n1093 = n1083 & n1092 ;
  assign n1094 = ~n1082 & n1093 ;
  assign n1091 = x7 & n1082 ;
  assign n1095 = n1094 ^ n1091 ;
  assign n1096 = n1095 ^ x7 ;
  assign n1097 = ~n1090 & ~n1096 ;
  assign n1098 = n1097 ^ n1095 ;
  assign n1099 = n1098 ^ n1073 ;
  assign n1100 = n1099 ^ x7 ;
  assign n1084 = ~n451 & n1083 ;
  assign n1085 = n1082 & n1084 ;
  assign n1086 = n1085 ^ n1084 ;
  assign n1087 = n1086 ^ n1082 ;
  assign n1088 = n1073 & ~n1087 ;
  assign n1089 = n1088 ^ n1087 ;
  assign n1101 = n1100 ^ n1089 ;
  assign n1113 = n825 ^ n63 ;
  assign n1126 = n1113 ^ n63 ;
  assign n1112 = n63 ^ x9 ;
  assign n1114 = n1113 ^ n1112 ;
  assign n1115 = n1112 ^ x7 ;
  assign n1116 = x2 ^ x1 ;
  assign n1117 = n1116 ^ x9 ;
  assign n1118 = n1117 ^ x9 ;
  assign n1119 = n1118 ^ n1114 ;
  assign n1120 = n1115 & ~n1119 ;
  assign n1121 = n1120 ^ x7 ;
  assign n1122 = n1121 ^ n1114 ;
  assign n1123 = ~n1114 & ~n1122 ;
  assign n1124 = n1123 ^ n1120 ;
  assign n1125 = n1124 ^ x7 ;
  assign n1127 = n1126 ^ n1125 ;
  assign n1128 = n1112 ^ n63 ;
  assign n1130 = n1118 ^ n1112 ;
  assign n1129 = n1113 ^ x7 ;
  assign n1131 = n1130 ^ n1129 ;
  assign n1132 = n1128 & ~n1131 ;
  assign n1133 = n1132 ^ n1123 ;
  assign n1134 = n1133 ^ n1120 ;
  assign n1135 = ~n1127 & n1134 ;
  assign n1136 = n1135 ^ x9 ;
  assign n1137 = n1136 ^ n1117 ;
  assign n1138 = x0 & ~n1137 ;
  assign n1139 = n1138 ^ x0 ;
  assign n1140 = n1139 ^ n1137 ;
  assign n1102 = n15 & n475 ;
  assign n1103 = n1102 ^ n773 ;
  assign n1104 = ~x2 & x7 ;
  assign n1105 = n1104 ^ n773 ;
  assign n1106 = ~n1104 & ~n1105 ;
  assign n1107 = n1106 ^ n1104 ;
  assign n1108 = n1107 ^ n1102 ;
  assign n1109 = ~n1103 & n1108 ;
  assign n1110 = n1109 ^ n1106 ;
  assign n1111 = n1110 ^ n1102 ;
  assign n1154 = x3 & n881 ;
  assign n1155 = ~n1111 & n1154 ;
  assign n1156 = ~n1140 & n1155 ;
  assign n1153 = x3 & ~n881 ;
  assign n1157 = n1156 ^ n1153 ;
  assign n1158 = n1101 & n1157 ;
  assign n1159 = n1158 ^ x3 ;
  assign n1141 = n1140 ^ n1111 ;
  assign n1142 = n1111 ^ n881 ;
  assign n1143 = ~n881 & n1142 ;
  assign n1144 = n1143 ^ n881 ;
  assign n1145 = n1144 ^ n1140 ;
  assign n1146 = n1141 & n1145 ;
  assign n1147 = n1146 ^ n1143 ;
  assign n1148 = n1147 ^ n1140 ;
  assign n1149 = n1101 & n1148 ;
  assign n1150 = n1149 ^ n1148 ;
  assign n1151 = n1150 ^ n1148 ;
  assign n1152 = n1151 ^ n1101 ;
  assign n1160 = n1159 ^ n1152 ;
  assign n1161 = x4 & n1160 ;
  assign n1162 = n1161 ^ n1160 ;
  assign n1216 = n47 ^ x6 ;
  assign n1203 = n1074 ^ x5 ;
  assign n1204 = n1203 ^ x2 ;
  assign n1212 = n1204 ^ n47 ;
  assign n1213 = n47 & n1212 ;
  assign n1205 = n1204 ^ x5 ;
  assign n1206 = n1205 ^ x9 ;
  assign n1207 = n1206 ^ x6 ;
  assign n1208 = x9 & n1207 ;
  assign n1209 = n1208 ^ x6 ;
  assign n1210 = n1209 ^ x9 ;
  assign n1211 = ~x6 & ~n1210 ;
  assign n1214 = n1213 ^ n1211 ;
  assign n1215 = n1214 ^ n1208 ;
  assign n1217 = n1216 ^ n1215 ;
  assign n1219 = n1206 ^ x9 ;
  assign n1218 = n1211 ^ x6 ;
  assign n1220 = n1219 ^ n1218 ;
  assign n1221 = ~n1217 & n1220 ;
  assign n1222 = n1221 ^ n1211 ;
  assign n1223 = n1222 ^ n1209 ;
  assign n1224 = n1223 ^ n314 ;
  assign n1225 = n1224 ^ x2 ;
  assign n1226 = n1225 ^ x5 ;
  assign n1227 = n1226 ^ n1203 ;
  assign n1199 = n233 & ~n475 ;
  assign n1200 = n1199 ^ x9 ;
  assign n1198 = ~x9 & n415 ;
  assign n1201 = n1200 ^ n1198 ;
  assign n1231 = n732 & n1201 ;
  assign n1232 = ~n1227 & n1231 ;
  assign n1228 = x8 & n1227 ;
  assign n1229 = n1228 ^ x8 ;
  assign n1230 = n1229 ^ n1227 ;
  assign n1233 = n1232 ^ n1230 ;
  assign n1202 = x6 & n1201 ;
  assign n1234 = n1233 ^ n1202 ;
  assign n1192 = n12 & n415 ;
  assign n1193 = ~x0 & ~n732 ;
  assign n1194 = n153 ^ x9 ;
  assign n1195 = ~n506 & ~n1194 ;
  assign n1196 = ~n1193 & n1195 ;
  assign n1197 = ~n1192 & ~n1196 ;
  assign n1235 = n1234 ^ n1197 ;
  assign n1236 = x1 & n1235 ;
  assign n1237 = n1236 ^ n1235 ;
  assign n1238 = n1237 ^ n1234 ;
  assign n1163 = n619 ^ x0 ;
  assign n1164 = n1163 ^ x6 ;
  assign n1165 = ~n878 & ~n1164 ;
  assign n1166 = n1165 ^ n1164 ;
  assign n1167 = ~n249 & n809 ;
  assign n1168 = n1166 & n1167 ;
  assign n1169 = n1168 ^ n809 ;
  assign n1171 = n320 & n773 ;
  assign n1172 = n1171 ^ x0 ;
  assign n1170 = ~x9 & n149 ;
  assign n1173 = n1172 ^ n1170 ;
  assign n1177 = x5 & ~n1173 ;
  assign n1178 = ~n1169 & n1177 ;
  assign n1179 = n1178 ^ x5 ;
  assign n1174 = n1169 & n1173 ;
  assign n1175 = n1174 ^ n1169 ;
  assign n1176 = n1175 ^ n1173 ;
  assign n1180 = n1179 ^ n1176 ;
  assign n1185 = ~x0 & ~x8 ;
  assign n1186 = n26 & ~n822 ;
  assign n1187 = ~n1185 & n1186 ;
  assign n1182 = n156 & n256 ;
  assign n1181 = n276 & ~n1042 ;
  assign n1183 = n1182 ^ n1181 ;
  assign n1184 = x9 & n1183 ;
  assign n1188 = n1187 ^ n1184 ;
  assign n1189 = x3 & ~n1188 ;
  assign n1190 = ~n1180 & n1189 ;
  assign n1191 = n1190 ^ x3 ;
  assign n1239 = n1238 ^ n1191 ;
  assign n1241 = ~x1 & x7 ;
  assign n1242 = n1235 & n1241 ;
  assign n1240 = x7 & ~n1234 ;
  assign n1243 = n1242 ^ n1240 ;
  assign n1244 = n1243 ^ x7 ;
  assign n1245 = n1244 ^ n1191 ;
  assign n1246 = ~n1239 & ~n1245 ;
  assign n1247 = n1246 ^ n1243 ;
  assign n1248 = n1247 ^ n1191 ;
  assign n1252 = x4 & ~n151 ;
  assign n1253 = ~n265 & n1252 ;
  assign n1254 = ~n356 & ~n1253 ;
  assign n1255 = ~x7 & ~n1254 ;
  assign n1257 = ~n1248 & n1255 ;
  assign n1258 = n1162 & n1257 ;
  assign n1256 = x4 & n1255 ;
  assign n1259 = n1258 ^ n1256 ;
  assign n1260 = n1259 ^ n1255 ;
  assign n1261 = n1260 ^ n1255 ;
  assign n1249 = n1162 & n1248 ;
  assign n1250 = n1249 ^ n1162 ;
  assign n1251 = n1250 ^ x4 ;
  assign n1262 = n1261 ^ n1251 ;
  assign n1272 = ~x5 & ~x7 ;
  assign n1273 = n1039 & n1272 ;
  assign n1274 = ~x6 & n1273 ;
  assign n1263 = n558 & n1042 ;
  assign n1264 = x8 & n156 ;
  assign n1265 = x7 & x9 ;
  assign n1266 = n1265 ^ x7 ;
  assign n1267 = n1264 & n1266 ;
  assign n1268 = ~n1263 & ~n1267 ;
  assign n1269 = ~n362 & n881 ;
  assign n1270 = ~n1268 & n1269 ;
  assign n1277 = n1274 ^ n1270 ;
  assign n1447 = n1274 ^ x7 ;
  assign n1448 = n1277 & n1447 ;
  assign n1449 = n1448 ^ x7 ;
  assign n1281 = x0 & ~x9 ;
  assign n1282 = n256 & n1281 ;
  assign n1279 = ~x0 & ~x9 ;
  assign n1280 = ~n428 & n1279 ;
  assign n1283 = n1282 ^ n1280 ;
  assign n1284 = x2 & n773 ;
  assign n1285 = n202 ^ x3 ;
  assign n1286 = n1285 ^ x8 ;
  assign n1287 = x6 & n1286 ;
  assign n1288 = n1287 ^ n1286 ;
  assign n1289 = n1284 & n1288 ;
  assign n1290 = n1289 ^ n1284 ;
  assign n1291 = n1283 & n1290 ;
  assign n1292 = n1291 ^ n1283 ;
  assign n1293 = n1292 ^ n1290 ;
  assign n1297 = x8 & n620 ;
  assign n1296 = ~n239 & n323 ;
  assign n1298 = n1297 ^ n1296 ;
  assign n1294 = ~n349 & n1042 ;
  assign n1295 = n1294 ^ n1279 ;
  assign n1299 = n1298 ^ n1295 ;
  assign n1347 = n360 & n1299 ;
  assign n1348 = n1347 ^ x1 ;
  assign n1349 = ~n1293 & n1348 ;
  assign n1336 = ~x0 & ~x6 ;
  assign n1337 = n322 & n1336 ;
  assign n1334 = ~x3 & x6 ;
  assign n1335 = n322 & n1334 ;
  assign n1338 = n1337 ^ n1335 ;
  assign n1331 = x0 & ~x3 ;
  assign n1332 = n345 & n1331 ;
  assign n1333 = n1332 ^ n210 ;
  assign n1339 = n1338 ^ n1333 ;
  assign n1340 = n1339 ^ x2 ;
  assign n1323 = ~n349 & n1286 ;
  assign n1324 = n1323 ^ n349 ;
  assign n1325 = x2 & ~n1324 ;
  assign n1341 = n1339 ^ n1325 ;
  assign n1342 = n1340 & n1341 ;
  assign n1304 = x8 ^ x6 ;
  assign n1305 = n1304 ^ n558 ;
  assign n1306 = n1304 ^ x9 ;
  assign n1307 = n558 ^ x0 ;
  assign n1308 = n1307 ^ n70 ;
  assign n1309 = n1308 ^ n70 ;
  assign n1310 = n1306 & n1309 ;
  assign n1311 = n1310 ^ n1304 ;
  assign n1312 = n1305 & n1311 ;
  assign n1313 = n1312 ^ n1311 ;
  assign n1314 = n1313 ^ n1306 ;
  assign n1315 = n1304 & n1308 ;
  assign n1316 = n1315 ^ n1305 ;
  assign n1317 = n1314 & n1316 ;
  assign n1318 = n1317 ^ n1314 ;
  assign n1319 = n1318 ^ n1315 ;
  assign n1320 = n1319 ^ n1304 ;
  assign n1321 = n1320 ^ x8 ;
  assign n1322 = n1321 ^ n1304 ;
  assign n1326 = n1325 ^ x2 ;
  assign n1327 = n1326 ^ n1324 ;
  assign n1328 = n1322 & n1327 ;
  assign n1329 = n1328 ^ n1327 ;
  assign n1330 = n1329 ^ x2 ;
  assign n1343 = n1342 ^ n1330 ;
  assign n1344 = n1343 ^ n1339 ;
  assign n1345 = x1 & n1344 ;
  assign n1346 = n1345 ^ x1 ;
  assign n1350 = n1349 ^ n1346 ;
  assign n1300 = x3 & n1299 ;
  assign n1301 = ~n1293 & n1300 ;
  assign n1302 = n1301 ^ n1293 ;
  assign n1303 = n1302 ^ x1 ;
  assign n1351 = n1350 ^ n1303 ;
  assign n1352 = x3 & ~n428 ;
  assign n1353 = n353 & n1352 ;
  assign n1354 = ~x5 & ~n1353 ;
  assign n1355 = ~n1351 & n1354 ;
  assign n1356 = n1355 ^ x5 ;
  assign n1397 = n17 & ~n1194 ;
  assign n1408 = x0 & ~x8 ;
  assign n1409 = n1397 & n1408 ;
  assign n1403 = ~x0 & x8 ;
  assign n1406 = n1397 ^ n17 ;
  assign n1407 = n1403 & n1406 ;
  assign n1410 = n1409 ^ n1407 ;
  assign n1374 = n17 & n153 ;
  assign n1404 = n1374 ^ n153 ;
  assign n1405 = n1403 & n1404 ;
  assign n1411 = n1410 ^ n1405 ;
  assign n1375 = n1374 ^ n17 ;
  assign n1376 = n1375 ^ n153 ;
  assign n1377 = x0 & ~n1376 ;
  assign n1378 = n1377 ^ x0 ;
  assign n1379 = n1378 ^ n1376 ;
  assign n1412 = n1411 ^ n1379 ;
  assign n1361 = ~x2 & x5 ;
  assign n1402 = x3 & n1361 ;
  assign n1413 = n1412 ^ n1402 ;
  assign n1419 = n1412 ^ x8 ;
  assign n1381 = n47 ^ x9 ;
  assign n1382 = n1381 ^ x5 ;
  assign n1383 = n1382 ^ x8 ;
  assign n1384 = n1383 ^ n559 ;
  assign n1385 = n1381 ^ x0 ;
  assign n1386 = n1385 ^ x5 ;
  assign n1387 = n825 & n1386 ;
  assign n1388 = n1387 ^ n825 ;
  assign n1389 = n1388 ^ n1383 ;
  assign n1390 = n1384 & n1389 ;
  assign n1391 = n1390 ^ n1384 ;
  assign n1392 = n1391 ^ n1389 ;
  assign n1393 = n1392 ^ n1383 ;
  assign n1394 = x3 & ~n1393 ;
  assign n1395 = n1394 ^ x3 ;
  assign n1396 = n1395 ^ n1393 ;
  assign n1398 = n1397 ^ n1396 ;
  assign n1420 = n1419 ^ n1398 ;
  assign n1421 = n1413 & ~n1420 ;
  assign n1422 = n1421 ^ n1413 ;
  assign n1432 = n1422 ^ n1411 ;
  assign n1400 = n1397 ^ x8 ;
  assign n1401 = n1400 ^ n1396 ;
  assign n1414 = n1413 ^ n1401 ;
  assign n1415 = n1402 ^ x8 ;
  assign n1416 = n1415 ^ n1412 ;
  assign n1417 = ~n1414 & n1416 ;
  assign n1418 = n1417 ^ n1414 ;
  assign n1423 = n1422 ^ n1418 ;
  assign n1424 = n1423 ^ n1412 ;
  assign n1425 = n1424 ^ n1401 ;
  assign n1426 = n1422 ^ n1402 ;
  assign n1427 = n1426 ^ n1396 ;
  assign n1428 = n1425 & ~n1427 ;
  assign n1429 = n1428 ^ n1425 ;
  assign n1430 = n1429 ^ n1427 ;
  assign n1431 = n1430 ^ n1418 ;
  assign n1433 = n1432 ^ n1431 ;
  assign n1380 = n1379 ^ x8 ;
  assign n1399 = n1398 ^ n1380 ;
  assign n1434 = n1433 ^ n1399 ;
  assign n1357 = x0 & x3 ;
  assign n1358 = x2 & ~n773 ;
  assign n1359 = n1357 & n1358 ;
  assign n1360 = ~n263 & n558 ;
  assign n1362 = ~n1357 & n1361 ;
  assign n1363 = n1362 ^ x5 ;
  assign n1364 = n1360 & n1363 ;
  assign n1365 = n1364 ^ n1363 ;
  assign n1366 = n1359 & n1365 ;
  assign n1367 = n1366 ^ n1359 ;
  assign n1368 = n1367 ^ n1365 ;
  assign n1435 = n1434 ^ n1368 ;
  assign n1436 = n1435 ^ n1368 ;
  assign n1373 = n1368 ^ x1 ;
  assign n1437 = n1436 ^ n1373 ;
  assign n1369 = x8 & n776 ;
  assign n1370 = n949 & n1369 ;
  assign n1371 = n1370 ^ x6 ;
  assign n1438 = x1 & ~n1371 ;
  assign n1439 = ~n1437 & n1438 ;
  assign n1372 = ~n1368 & ~n1371 ;
  assign n1440 = n1439 ^ n1372 ;
  assign n1441 = n1440 ^ x6 ;
  assign n1442 = n1356 & n1441 ;
  assign n1443 = n1442 ^ n1356 ;
  assign n1444 = n1443 ^ n1441 ;
  assign n1445 = n1444 ^ n1356 ;
  assign n1446 = n1445 ^ n1441 ;
  assign n1450 = n1449 ^ n1446 ;
  assign n1455 = n1449 ^ n1270 ;
  assign n1275 = n1274 ^ x4 ;
  assign n1456 = n1455 ^ n1275 ;
  assign n1457 = ~n1450 & n1456 ;
  assign n1458 = n1457 ^ n1456 ;
  assign n1278 = n1277 ^ x4 ;
  assign n1451 = n1450 ^ n1278 ;
  assign n1452 = n1446 ^ n1270 ;
  assign n1453 = n1452 ^ n1449 ;
  assign n1454 = ~n1451 & ~n1453 ;
  assign n1459 = n1458 ^ n1454 ;
  assign n1460 = n1459 ^ n1449 ;
  assign n1461 = n1460 ^ n1278 ;
  assign n1462 = n1458 ^ n1446 ;
  assign n1463 = n1462 ^ x4 ;
  assign n1464 = n1461 & ~n1463 ;
  assign n1465 = n1464 ^ n1461 ;
  assign n1466 = n1465 ^ n1454 ;
  assign n1467 = n1466 ^ n1458 ;
  assign n1468 = n1467 ^ n1448 ;
  assign n1271 = n1270 ^ x7 ;
  assign n1276 = n1275 ^ n1271 ;
  assign n1469 = n1468 ^ n1276 ;
  assign n1470 = n1469 ^ n1274 ;
  assign n1501 = ~x5 & ~n476 ;
  assign n1502 = ~n17 & n249 ;
  assign n1503 = ~n1501 & n1502 ;
  assign n1505 = n418 ^ x5 ;
  assign n1507 = n1505 ^ x3 ;
  assign n1506 = n1505 ^ x5 ;
  assign n1508 = n1507 ^ n1506 ;
  assign n1504 = n910 ^ n48 ;
  assign n1509 = n1508 ^ n1504 ;
  assign n1510 = n1508 ^ n910 ;
  assign n1511 = ~n1509 & n1510 ;
  assign n1512 = n1511 ^ n1508 ;
  assign n1515 = n1508 ^ n1507 ;
  assign n1516 = n1515 ^ n1510 ;
  assign n1517 = n1516 ^ n1509 ;
  assign n1518 = n1508 ^ n1505 ;
  assign n1519 = n1518 ^ n1510 ;
  assign n1520 = n1519 ^ n1509 ;
  assign n1521 = n1517 & n1520 ;
  assign n1513 = n1510 ^ n1509 ;
  assign n1514 = n1513 ^ n1508 ;
  assign n1522 = n1521 ^ n1514 ;
  assign n1523 = ~n1512 & n1522 ;
  assign n1524 = n1523 ^ n1508 ;
  assign n1525 = n1524 ^ n1508 ;
  assign n1546 = n322 & n1525 ;
  assign n1547 = ~n1503 & n1546 ;
  assign n1545 = x9 & ~n1503 ;
  assign n1548 = n1547 ^ n1545 ;
  assign n1537 = ~x1 & x3 ;
  assign n1538 = ~x0 & x5 ;
  assign n1539 = n416 & ~n1538 ;
  assign n1540 = n1537 & n1539 ;
  assign n1531 = x2 & x5 ;
  assign n1532 = n1531 ^ x2 ;
  assign n1533 = ~n17 & ~n1532 ;
  assign n1535 = n360 & ~n416 ;
  assign n1536 = ~n1533 & n1535 ;
  assign n1541 = n1540 ^ n1536 ;
  assign n1534 = x1 & ~n1533 ;
  assign n1542 = n1541 ^ n1534 ;
  assign n1544 = x9 & ~n1542 ;
  assign n1549 = n1548 ^ n1544 ;
  assign n1526 = x8 & ~n1525 ;
  assign n1527 = n1526 ^ x8 ;
  assign n1528 = n1503 & n1527 ;
  assign n1529 = n1528 ^ n1527 ;
  assign n1530 = n1529 ^ n1503 ;
  assign n1543 = n1542 ^ n1530 ;
  assign n1550 = n1549 ^ n1543 ;
  assign n1551 = n1550 ^ n1542 ;
  assign n1483 = ~n269 & n1361 ;
  assign n1484 = n1483 ^ n731 ;
  assign n1485 = ~x0 & n1484 ;
  assign n1486 = n313 ^ x1 ;
  assign n1487 = n1486 ^ x5 ;
  assign n1488 = n809 & n1487 ;
  assign n1489 = n264 & ~n1488 ;
  assign n1490 = ~n1485 & ~n1489 ;
  assign n1492 = ~x2 & n269 ;
  assign n1493 = ~n730 & n1492 ;
  assign n1494 = x3 ^ x1 ;
  assign n1495 = x5 & n1494 ;
  assign n1496 = n1495 ^ x3 ;
  assign n1497 = ~x8 & ~n1496 ;
  assign n1498 = n1493 & n1497 ;
  assign n1499 = n1490 & n1498 ;
  assign n1491 = ~x8 & ~n1490 ;
  assign n1500 = n1499 ^ n1491 ;
  assign n1552 = n1551 ^ n1500 ;
  assign n1553 = n1551 ^ x6 ;
  assign n1554 = x6 & ~n1553 ;
  assign n1555 = n1554 ^ x6 ;
  assign n1556 = n1555 ^ n1500 ;
  assign n1557 = n1552 & ~n1556 ;
  assign n1558 = n1557 ^ n1554 ;
  assign n1559 = n1558 ^ n1500 ;
  assign n1560 = ~x6 & ~n276 ;
  assign n1561 = ~n1172 & n1560 ;
  assign n1562 = x6 & n16 ;
  assign n1563 = n1562 ^ x6 ;
  assign n1564 = ~n26 & n476 ;
  assign n1565 = n1563 & ~n1564 ;
  assign n1566 = ~x2 & ~n1565 ;
  assign n1567 = n18 & ~n1566 ;
  assign n1568 = ~n1561 & n1567 ;
  assign n1569 = n1559 & n1568 ;
  assign n1570 = n1569 ^ n1559 ;
  assign n1571 = n1570 ^ n1568 ;
  assign n1471 = ~x4 & ~n1273 ;
  assign n1478 = ~x0 & ~n428 ;
  assign n1479 = n15 & n1478 ;
  assign n1473 = ~x2 & x8 ;
  assign n1474 = ~x9 & n1473 ;
  assign n1475 = n1474 ^ n1279 ;
  assign n1472 = ~x8 & n1042 ;
  assign n1476 = n1475 ^ n1472 ;
  assign n1477 = ~x1 & n1476 ;
  assign n1480 = n1479 ^ n1477 ;
  assign n1481 = n397 & n1480 ;
  assign n1572 = ~x7 & ~n1481 ;
  assign n1573 = n1471 & n1572 ;
  assign n1574 = n1571 & n1573 ;
  assign n1482 = n1471 & n1481 ;
  assign n1575 = n1574 ^ n1482 ;
  assign n1576 = n1575 ^ n1273 ;
  assign n1577 = x3 & n347 ;
  assign n1578 = n1577 ^ x3 ;
  assign n1579 = ~x6 & ~n776 ;
  assign n1580 = n476 & ~n1579 ;
  assign n1581 = n1578 & ~n1580 ;
  assign n1582 = ~n881 & n975 ;
  assign n1583 = ~x2 & ~n1582 ;
  assign n1584 = ~n1581 & n1583 ;
  assign n1585 = n264 & n773 ;
  assign n1586 = ~n974 & n1585 ;
  assign n1587 = ~n1584 & ~n1586 ;
  assign n1588 = ~x1 & ~n1587 ;
  assign n1589 = x2 & n955 ;
  assign n1590 = n974 & n1589 ;
  assign n1591 = n345 & n776 ;
  assign n1592 = n1591 ^ x6 ;
  assign n1593 = x3 & ~n1592 ;
  assign n1594 = n1593 ^ x3 ;
  assign n1595 = n1594 ^ n1592 ;
  assign n1596 = n1590 & n1595 ;
  assign n1597 = n1596 ^ n1590 ;
  assign n1598 = n1597 ^ n1595 ;
  assign n1605 = n935 ^ n347 ;
  assign n1606 = n1605 ^ n935 ;
  assign n1608 = n1606 ^ n935 ;
  assign n1625 = n1608 ^ n1606 ;
  assign n1626 = n1625 ^ x2 ;
  assign n1599 = n476 ^ x3 ;
  assign n1600 = n1599 ^ n476 ;
  assign n1602 = n1600 ^ n476 ;
  assign n1619 = n1602 ^ n1600 ;
  assign n1612 = n1608 ^ n1600 ;
  assign n1613 = n1612 ^ n1602 ;
  assign n1614 = n1608 ^ n1602 ;
  assign n1615 = n1614 ^ x2 ;
  assign n1616 = n1613 & n1615 ;
  assign n1603 = n1602 ^ x2 ;
  assign n1604 = n1602 & ~n1603 ;
  assign n1617 = n1616 ^ n1604 ;
  assign n1618 = n1617 ^ n1606 ;
  assign n1620 = n1619 ^ n1618 ;
  assign n1621 = n1616 ^ n1606 ;
  assign n1622 = ~n1620 & n1621 ;
  assign n1601 = n1600 ^ x2 ;
  assign n1609 = n1608 ^ x2 ;
  assign n1607 = n1606 ^ n1604 ;
  assign n1610 = n1609 ^ n1607 ;
  assign n1611 = n1601 & n1610 ;
  assign n1623 = n1622 ^ n1611 ;
  assign n1624 = n1623 ^ n1604 ;
  assign n1627 = n1626 ^ n1624 ;
  assign n1628 = x1 & ~n1627 ;
  assign n1629 = ~n1598 & n1628 ;
  assign n1630 = n1629 ^ x1 ;
  assign n1631 = x1 & n773 ;
  assign n1632 = n1631 ^ n773 ;
  assign n1633 = n822 & n1589 ;
  assign n1634 = ~x7 & ~n1633 ;
  assign n1635 = ~n1632 & ~n1634 ;
  assign n1636 = ~x7 & n767 ;
  assign n1637 = x0 & ~n1636 ;
  assign n1638 = ~x5 & ~n264 ;
  assign n1639 = x6 & ~n1638 ;
  assign n1640 = ~x2 & x4 ;
  assign n1641 = ~n362 & n1640 ;
  assign n1642 = n1641 ^ x4 ;
  assign n1643 = x7 & ~n264 ;
  assign n1644 = n1642 & n1643 ;
  assign n1645 = n1644 ^ n1642 ;
  assign n1646 = n1645 ^ n1643 ;
  assign n1647 = n1639 & ~n1646 ;
  assign n1648 = n1647 ^ n1646 ;
  assign n1649 = n1637 & ~n1648 ;
  assign n1650 = n1649 ^ n1648 ;
  assign n1651 = n1635 & ~n1650 ;
  assign n1652 = n1651 ^ n1650 ;
  assign n1653 = n1630 & ~n1652 ;
  assign n1654 = n1653 ^ n1652 ;
  assign n1655 = n1588 & ~n1654 ;
  assign n1656 = n1655 ^ n1654 ;
  assign n1657 = ~x7 & n881 ;
  assign n1658 = x8 & ~n14 ;
  assign n1659 = x1 & n30 ;
  assign n1660 = n1659 ^ x1 ;
  assign n1661 = n1660 ^ n30 ;
  assign n1662 = x2 & n1037 ;
  assign n1663 = n1661 & n1662 ;
  assign n1664 = ~n1658 & n1663 ;
  assign n1665 = ~n1039 & ~n1664 ;
  assign n1666 = n1657 & ~n1665 ;
  assign y0 = ~n396 ;
  assign y1 = ~n719 ;
  assign y2 = ~n890 ;
  assign y3 = ~n1029 ;
  assign y4 = n1036 ;
  assign y5 = n1041 ;
  assign y6 = n1262 ;
  assign y7 = ~n1470 ;
  assign y8 = ~n1576 ;
  assign y9 = ~n1656 ;
  assign y10 = n1666 ;
endmodule
