module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 ;
  assign n54 = x10 ^ x2 ;
  assign n83 = x3 & ~x11 ;
  assign n84 = ~n54 & n83 ;
  assign n82 = x2 & ~x10 ;
  assign n85 = n84 ^ n82 ;
  assign n49 = x8 ^ x0 ;
  assign n50 = x9 ^ x1 ;
  assign n51 = n49 & n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n52 ^ n50 ;
  assign n120 = x0 & ~n53 ;
  assign n121 = n85 & n120 ;
  assign n88 = x1 & ~x9 ;
  assign n89 = ~n49 & n88 ;
  assign n87 = x0 & ~x8 ;
  assign n90 = n89 ^ n87 ;
  assign n119 = x0 & ~n90 ;
  assign n122 = n121 ^ n119 ;
  assign n55 = x11 ^ x3 ;
  assign n56 = n54 & n55 ;
  assign n57 = n56 ^ n54 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n53 & n58 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = n60 ^ n58 ;
  assign n63 = x12 ^ x4 ;
  assign n67 = x13 ^ x5 ;
  assign n68 = n63 & n67 ;
  assign n69 = n68 ^ n63 ;
  assign n70 = n69 ^ n67 ;
  assign n72 = x14 ^ x6 ;
  assign n93 = x15 ^ x7 ;
  assign n94 = n72 & n93 ;
  assign n95 = n94 ^ n72 ;
  assign n96 = n95 ^ n93 ;
  assign n97 = n70 & n96 ;
  assign n98 = n97 ^ n70 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = ~n61 & ~n99 ;
  assign n117 = x0 & n100 ;
  assign n118 = n117 ^ x0 ;
  assign n123 = n122 ^ n118 ;
  assign n73 = x7 & x15 ;
  assign n74 = n73 ^ x7 ;
  assign n75 = n72 & n74 ;
  assign n76 = n75 ^ n74 ;
  assign n71 = x6 & ~x14 ;
  assign n77 = n76 ^ n71 ;
  assign n78 = n70 & n77 ;
  assign n79 = n78 ^ n77 ;
  assign n64 = x5 & ~x13 ;
  assign n65 = ~n63 & n64 ;
  assign n62 = x4 & ~x12 ;
  assign n66 = n65 ^ n62 ;
  assign n80 = n79 ^ n66 ;
  assign n115 = x0 & ~n61 ;
  assign n116 = n80 & n115 ;
  assign n124 = n123 ^ n116 ;
  assign n110 = x8 & ~n53 ;
  assign n111 = n85 & n110 ;
  assign n109 = x8 & n90 ;
  assign n112 = n111 ^ n109 ;
  assign n107 = x8 & n100 ;
  assign n108 = n107 ^ x8 ;
  assign n113 = n112 ^ n108 ;
  assign n105 = x8 & ~n61 ;
  assign n106 = n80 & n105 ;
  assign n114 = n113 ^ n106 ;
  assign n125 = n124 ^ n114 ;
  assign n127 = n125 ^ x16 ;
  assign n143 = x1 & ~n53 ;
  assign n144 = n85 & n143 ;
  assign n142 = x1 & ~n90 ;
  assign n145 = n144 ^ n142 ;
  assign n140 = x1 & n100 ;
  assign n141 = n140 ^ x1 ;
  assign n146 = n145 ^ n141 ;
  assign n138 = x1 & ~n61 ;
  assign n139 = n80 & n138 ;
  assign n147 = n146 ^ n139 ;
  assign n133 = x9 & ~n53 ;
  assign n134 = n85 & n133 ;
  assign n132 = x9 & n90 ;
  assign n135 = n134 ^ n132 ;
  assign n130 = x9 & n100 ;
  assign n131 = n130 ^ x9 ;
  assign n136 = n135 ^ n131 ;
  assign n128 = x9 & ~n61 ;
  assign n129 = n80 & n128 ;
  assign n137 = n136 ^ n129 ;
  assign n148 = n147 ^ n137 ;
  assign n149 = ~x17 & n148 ;
  assign n150 = ~n127 & n149 ;
  assign n126 = ~x16 & n125 ;
  assign n151 = n150 ^ n126 ;
  assign n610 = n125 & ~n151 ;
  assign n168 = x2 & ~n53 ;
  assign n169 = n85 & n168 ;
  assign n167 = x2 & ~n90 ;
  assign n170 = n169 ^ n167 ;
  assign n165 = x2 & n100 ;
  assign n166 = n165 ^ x2 ;
  assign n171 = n170 ^ n166 ;
  assign n163 = x2 & ~n61 ;
  assign n164 = n80 & n163 ;
  assign n172 = n171 ^ n164 ;
  assign n158 = x10 & ~n53 ;
  assign n159 = n85 & n158 ;
  assign n157 = x10 & n90 ;
  assign n160 = n159 ^ n157 ;
  assign n155 = x10 & n100 ;
  assign n156 = n155 ^ x10 ;
  assign n161 = n160 ^ n156 ;
  assign n153 = x10 & ~n61 ;
  assign n154 = n80 & n153 ;
  assign n162 = n161 ^ n154 ;
  assign n173 = n172 ^ n162 ;
  assign n175 = n173 ^ x18 ;
  assign n191 = x3 & ~n53 ;
  assign n192 = n85 & n191 ;
  assign n190 = x3 & ~n90 ;
  assign n193 = n192 ^ n190 ;
  assign n188 = x3 & n100 ;
  assign n189 = n188 ^ x3 ;
  assign n194 = n193 ^ n189 ;
  assign n186 = x3 & ~n61 ;
  assign n187 = n80 & n186 ;
  assign n195 = n194 ^ n187 ;
  assign n181 = x11 & ~n53 ;
  assign n182 = n85 & n181 ;
  assign n180 = x11 & n90 ;
  assign n183 = n182 ^ n180 ;
  assign n178 = x11 & n100 ;
  assign n179 = n178 ^ x11 ;
  assign n184 = n183 ^ n179 ;
  assign n176 = x11 & ~n61 ;
  assign n177 = n80 & n176 ;
  assign n185 = n184 ^ n177 ;
  assign n196 = n195 ^ n185 ;
  assign n197 = ~x19 & n196 ;
  assign n198 = ~n175 & n197 ;
  assign n174 = ~x18 & n173 ;
  assign n199 = n198 ^ n174 ;
  assign n200 = n148 ^ x17 ;
  assign n201 = n127 & n200 ;
  assign n202 = n201 ^ n127 ;
  assign n203 = n202 ^ n200 ;
  assign n204 = n125 & ~n203 ;
  assign n205 = n199 & n204 ;
  assign n611 = n610 ^ n205 ;
  assign n207 = n196 ^ x19 ;
  assign n208 = n175 & n207 ;
  assign n209 = n208 ^ n175 ;
  assign n210 = n209 ^ n207 ;
  assign n211 = n203 & n210 ;
  assign n212 = n211 ^ n203 ;
  assign n213 = n212 ^ n210 ;
  assign n229 = x4 & ~n53 ;
  assign n230 = n85 & n229 ;
  assign n228 = x4 & ~n90 ;
  assign n231 = n230 ^ n228 ;
  assign n226 = x4 & n100 ;
  assign n227 = n226 ^ x4 ;
  assign n232 = n231 ^ n227 ;
  assign n224 = x4 & ~n61 ;
  assign n225 = n80 & n224 ;
  assign n233 = n232 ^ n225 ;
  assign n219 = x12 & ~n53 ;
  assign n220 = n85 & n219 ;
  assign n218 = x12 & n90 ;
  assign n221 = n220 ^ n218 ;
  assign n216 = x12 & n100 ;
  assign n217 = n216 ^ x12 ;
  assign n222 = n221 ^ n217 ;
  assign n214 = x12 & ~n61 ;
  assign n215 = n80 & n214 ;
  assign n223 = n222 ^ n215 ;
  assign n234 = n233 ^ n223 ;
  assign n235 = n234 ^ x20 ;
  assign n251 = x5 & ~n53 ;
  assign n252 = n85 & n251 ;
  assign n250 = x5 & ~n90 ;
  assign n253 = n252 ^ n250 ;
  assign n248 = x5 & n100 ;
  assign n249 = n248 ^ x5 ;
  assign n254 = n253 ^ n249 ;
  assign n246 = x5 & ~n61 ;
  assign n247 = n80 & n246 ;
  assign n255 = n254 ^ n247 ;
  assign n241 = x13 & ~n53 ;
  assign n242 = n85 & n241 ;
  assign n240 = x13 & n90 ;
  assign n243 = n242 ^ n240 ;
  assign n238 = x13 & n100 ;
  assign n239 = n238 ^ x13 ;
  assign n244 = n243 ^ n239 ;
  assign n236 = x13 & ~n61 ;
  assign n237 = n80 & n236 ;
  assign n245 = n244 ^ n237 ;
  assign n256 = n255 ^ n245 ;
  assign n257 = n256 ^ x21 ;
  assign n258 = n235 & n257 ;
  assign n259 = n258 ^ n235 ;
  assign n260 = n259 ^ n257 ;
  assign n276 = x6 & ~n53 ;
  assign n277 = n85 & n276 ;
  assign n275 = x6 & ~n90 ;
  assign n278 = n277 ^ n275 ;
  assign n273 = x6 & n100 ;
  assign n274 = n273 ^ x6 ;
  assign n279 = n278 ^ n274 ;
  assign n271 = x6 & ~n61 ;
  assign n272 = n80 & n271 ;
  assign n280 = n279 ^ n272 ;
  assign n266 = x14 & ~n53 ;
  assign n267 = n85 & n266 ;
  assign n265 = x14 & n90 ;
  assign n268 = n267 ^ n265 ;
  assign n263 = x14 & n100 ;
  assign n264 = n263 ^ x14 ;
  assign n269 = n268 ^ n264 ;
  assign n261 = x14 & ~n61 ;
  assign n262 = n80 & n261 ;
  assign n270 = n269 ^ n262 ;
  assign n281 = n280 ^ n270 ;
  assign n282 = n281 ^ x22 ;
  assign n299 = x7 & ~n53 ;
  assign n300 = n85 & n299 ;
  assign n298 = x7 & ~n90 ;
  assign n301 = n300 ^ n298 ;
  assign n296 = x7 & n100 ;
  assign n297 = n296 ^ x7 ;
  assign n302 = n301 ^ n297 ;
  assign n294 = x7 & ~n61 ;
  assign n295 = n80 & n294 ;
  assign n303 = n302 ^ n295 ;
  assign n288 = x15 & ~n53 ;
  assign n289 = n85 & n288 ;
  assign n287 = x15 & ~n90 ;
  assign n290 = n289 ^ n287 ;
  assign n285 = x15 & n100 ;
  assign n286 = n285 ^ x15 ;
  assign n291 = n290 ^ n286 ;
  assign n283 = x15 & ~n61 ;
  assign n284 = n80 & n283 ;
  assign n292 = n291 ^ n284 ;
  assign n293 = n292 ^ x15 ;
  assign n304 = n303 ^ n293 ;
  assign n305 = n304 ^ x23 ;
  assign n306 = n282 & n305 ;
  assign n307 = n306 ^ n282 ;
  assign n308 = n307 ^ n305 ;
  assign n309 = n260 & n308 ;
  assign n310 = n309 ^ n260 ;
  assign n311 = n310 ^ n308 ;
  assign n312 = ~n213 & ~n311 ;
  assign n313 = n125 & n312 ;
  assign n314 = n313 ^ n125 ;
  assign n612 = n611 ^ n314 ;
  assign n316 = n125 & ~n213 ;
  assign n322 = x23 & n304 ;
  assign n323 = n322 ^ n304 ;
  assign n324 = n282 & n323 ;
  assign n325 = n324 ^ n323 ;
  assign n321 = ~x22 & n281 ;
  assign n326 = n325 ^ n321 ;
  assign n327 = n260 & n326 ;
  assign n328 = n327 ^ n326 ;
  assign n318 = ~x21 & n256 ;
  assign n319 = ~n235 & n318 ;
  assign n317 = ~x20 & n234 ;
  assign n320 = n319 ^ n317 ;
  assign n329 = n328 ^ n320 ;
  assign n330 = n316 & n329 ;
  assign n613 = n612 ^ n330 ;
  assign n606 = x16 & n151 ;
  assign n333 = x16 & ~n203 ;
  assign n334 = n199 & n333 ;
  assign n607 = n606 ^ n334 ;
  assign n336 = x16 & n312 ;
  assign n337 = n336 ^ x16 ;
  assign n608 = n607 ^ n337 ;
  assign n339 = x16 & ~n213 ;
  assign n340 = n329 & n339 ;
  assign n609 = n608 ^ n340 ;
  assign n614 = n613 ^ n609 ;
  assign n616 = n614 ^ x24 ;
  assign n621 = n148 & ~n151 ;
  assign n349 = n148 & ~n203 ;
  assign n350 = n199 & n349 ;
  assign n622 = n621 ^ n350 ;
  assign n352 = n148 & n312 ;
  assign n353 = n352 ^ n148 ;
  assign n623 = n622 ^ n353 ;
  assign n355 = n148 & ~n213 ;
  assign n356 = n329 & n355 ;
  assign n624 = n623 ^ n356 ;
  assign n617 = x17 & n151 ;
  assign n359 = x17 & ~n203 ;
  assign n360 = n199 & n359 ;
  assign n618 = n617 ^ n360 ;
  assign n362 = x17 & n312 ;
  assign n363 = n362 ^ x17 ;
  assign n619 = n618 ^ n363 ;
  assign n365 = x17 & ~n213 ;
  assign n366 = n329 & n365 ;
  assign n620 = n619 ^ n366 ;
  assign n625 = n624 ^ n620 ;
  assign n629 = n625 ^ x25 ;
  assign n630 = n616 & n629 ;
  assign n631 = n630 ^ n616 ;
  assign n632 = n631 ^ n629 ;
  assign n637 = ~n151 & n173 ;
  assign n380 = n173 & ~n203 ;
  assign n381 = n199 & n380 ;
  assign n638 = n637 ^ n381 ;
  assign n383 = n173 & n312 ;
  assign n384 = n383 ^ n173 ;
  assign n639 = n638 ^ n384 ;
  assign n386 = n173 & ~n213 ;
  assign n387 = n329 & n386 ;
  assign n640 = n639 ^ n387 ;
  assign n633 = x18 & n151 ;
  assign n390 = x18 & ~n203 ;
  assign n391 = n199 & n390 ;
  assign n634 = n633 ^ n391 ;
  assign n393 = x18 & n312 ;
  assign n394 = n393 ^ x18 ;
  assign n635 = n634 ^ n394 ;
  assign n396 = x18 & ~n213 ;
  assign n397 = n329 & n396 ;
  assign n636 = n635 ^ n397 ;
  assign n641 = n640 ^ n636 ;
  assign n643 = n641 ^ x26 ;
  assign n648 = ~n151 & n196 ;
  assign n403 = n196 & ~n203 ;
  assign n404 = n199 & n403 ;
  assign n649 = n648 ^ n404 ;
  assign n406 = n196 & n312 ;
  assign n407 = n406 ^ n196 ;
  assign n650 = n649 ^ n407 ;
  assign n409 = n196 & ~n213 ;
  assign n410 = n329 & n409 ;
  assign n651 = n650 ^ n410 ;
  assign n644 = x19 & n151 ;
  assign n413 = x19 & ~n203 ;
  assign n414 = n199 & n413 ;
  assign n645 = n644 ^ n414 ;
  assign n416 = x19 & n312 ;
  assign n417 = n416 ^ x19 ;
  assign n646 = n645 ^ n417 ;
  assign n419 = x19 & ~n213 ;
  assign n420 = n329 & n419 ;
  assign n647 = n646 ^ n420 ;
  assign n652 = n651 ^ n647 ;
  assign n661 = n652 ^ x27 ;
  assign n662 = n643 & n661 ;
  assign n663 = n662 ^ n643 ;
  assign n664 = n663 ^ n661 ;
  assign n665 = n632 & n664 ;
  assign n666 = n665 ^ n632 ;
  assign n667 = n666 ^ n664 ;
  assign n601 = ~n151 & n234 ;
  assign n442 = ~n203 & n234 ;
  assign n443 = n199 & n442 ;
  assign n602 = n601 ^ n443 ;
  assign n445 = n234 & n312 ;
  assign n446 = n445 ^ n234 ;
  assign n603 = n602 ^ n446 ;
  assign n448 = ~n213 & n234 ;
  assign n449 = n329 & n448 ;
  assign n604 = n603 ^ n449 ;
  assign n597 = x20 & n151 ;
  assign n452 = x20 & ~n203 ;
  assign n453 = n199 & n452 ;
  assign n598 = n597 ^ n453 ;
  assign n455 = x20 & n312 ;
  assign n456 = n455 ^ x20 ;
  assign n599 = n598 ^ n456 ;
  assign n458 = x20 & ~n213 ;
  assign n459 = n329 & n458 ;
  assign n600 = n599 ^ n459 ;
  assign n605 = n604 ^ n600 ;
  assign n669 = n605 ^ x28 ;
  assign n674 = ~n151 & n256 ;
  assign n468 = ~n203 & n256 ;
  assign n469 = n199 & n468 ;
  assign n675 = n674 ^ n469 ;
  assign n471 = n256 & n312 ;
  assign n472 = n471 ^ n256 ;
  assign n676 = n675 ^ n472 ;
  assign n474 = ~n213 & n256 ;
  assign n475 = n329 & n474 ;
  assign n677 = n676 ^ n475 ;
  assign n670 = x21 & n151 ;
  assign n478 = x21 & ~n203 ;
  assign n479 = n199 & n478 ;
  assign n671 = n670 ^ n479 ;
  assign n481 = x21 & n312 ;
  assign n482 = n481 ^ x21 ;
  assign n672 = n671 ^ n482 ;
  assign n484 = x21 & ~n213 ;
  assign n485 = n329 & n484 ;
  assign n673 = n672 ^ n485 ;
  assign n678 = n677 ^ n673 ;
  assign n684 = n678 ^ x29 ;
  assign n685 = n669 & n684 ;
  assign n686 = n685 ^ n669 ;
  assign n687 = n686 ^ n684 ;
  assign n729 = x22 & n151 ;
  assign n511 = x22 & ~n203 ;
  assign n512 = n199 & n511 ;
  assign n730 = n729 ^ n512 ;
  assign n514 = x22 & n312 ;
  assign n515 = n514 ^ x22 ;
  assign n731 = n730 ^ n515 ;
  assign n517 = x22 & ~n213 ;
  assign n518 = n329 & n517 ;
  assign n732 = n731 ^ n518 ;
  assign n724 = ~n151 & n281 ;
  assign n501 = ~n203 & n281 ;
  assign n502 = n199 & n501 ;
  assign n725 = n724 ^ n502 ;
  assign n504 = n281 & n312 ;
  assign n505 = n504 ^ n281 ;
  assign n726 = n725 ^ n505 ;
  assign n507 = ~n213 & n281 ;
  assign n508 = n329 & n507 ;
  assign n727 = n726 ^ n508 ;
  assign n751 = n732 ^ n727 ;
  assign n752 = n751 ^ x30 ;
  assign n579 = x23 & ~n203 ;
  assign n580 = n199 & n579 ;
  assign n578 = x23 & ~n151 ;
  assign n581 = n580 ^ n578 ;
  assign n576 = x23 & n312 ;
  assign n577 = n576 ^ x23 ;
  assign n582 = n581 ^ n577 ;
  assign n574 = x23 & ~n213 ;
  assign n575 = n329 & n574 ;
  assign n583 = n582 ^ n575 ;
  assign n720 = n583 ^ x23 ;
  assign n568 = ~n203 & n304 ;
  assign n569 = n199 & n568 ;
  assign n567 = ~n151 & n304 ;
  assign n570 = n569 ^ n567 ;
  assign n565 = n304 & n312 ;
  assign n566 = n565 ^ n304 ;
  assign n571 = n570 ^ n566 ;
  assign n563 = ~n213 & n304 ;
  assign n564 = n329 & n563 ;
  assign n572 = n571 ^ n564 ;
  assign n721 = n720 ^ n572 ;
  assign n753 = n721 ^ x31 ;
  assign n754 = n752 & n753 ;
  assign n755 = n754 ^ n752 ;
  assign n756 = n755 ^ n753 ;
  assign n757 = n687 & n756 ;
  assign n758 = n757 ^ n687 ;
  assign n759 = n758 ^ n756 ;
  assign n760 = ~n667 & ~n759 ;
  assign n737 = x22 & ~x30 ;
  assign n741 = n312 & n737 ;
  assign n692 = n199 & ~n203 ;
  assign n693 = n692 ^ n151 ;
  assign n740 = ~n693 & n737 ;
  assign n742 = n741 ^ n740 ;
  assign n738 = ~n213 & n737 ;
  assign n739 = n329 & n738 ;
  assign n743 = n742 ^ n739 ;
  assign n708 = x23 & x31 ;
  assign n714 = ~n203 & n708 ;
  assign n715 = n199 & n714 ;
  assign n713 = n151 & n708 ;
  assign n716 = n715 ^ n713 ;
  assign n711 = n312 & n708 ;
  assign n712 = n711 ^ n708 ;
  assign n717 = n716 ^ n712 ;
  assign n709 = ~n213 & n708 ;
  assign n710 = n329 & n709 ;
  assign n718 = n717 ^ n710 ;
  assign n697 = x31 & n304 ;
  assign n703 = ~n203 & n697 ;
  assign n704 = n199 & n703 ;
  assign n702 = ~n151 & n697 ;
  assign n705 = n704 ^ n702 ;
  assign n700 = n312 & n697 ;
  assign n701 = n700 ^ n697 ;
  assign n706 = n705 ^ n701 ;
  assign n698 = ~n213 & n697 ;
  assign n699 = n329 & n698 ;
  assign n707 = n706 ^ n699 ;
  assign n719 = n718 ^ n707 ;
  assign n722 = n721 ^ n719 ;
  assign n733 = n722 & n732 ;
  assign n728 = n722 & n727 ;
  assign n734 = n733 ^ n728 ;
  assign n723 = x30 & n722 ;
  assign n735 = n734 ^ n723 ;
  assign n736 = n735 ^ n722 ;
  assign n744 = n743 ^ n736 ;
  assign n688 = ~x30 & n281 ;
  assign n694 = n688 & ~n693 ;
  assign n691 = ~n312 & n688 ;
  assign n695 = n694 ^ n691 ;
  assign n689 = ~n213 & n688 ;
  assign n690 = n329 & n689 ;
  assign n696 = n695 ^ n690 ;
  assign n745 = n744 ^ n696 ;
  assign n746 = n687 & n745 ;
  assign n747 = n746 ^ n745 ;
  assign n679 = x29 & n678 ;
  assign n680 = n679 ^ n678 ;
  assign n681 = n669 & n680 ;
  assign n682 = n681 ^ n680 ;
  assign n668 = ~x28 & n605 ;
  assign n683 = n682 ^ n668 ;
  assign n748 = n747 ^ n683 ;
  assign n749 = ~n667 & n748 ;
  assign n653 = x27 & n652 ;
  assign n654 = n653 ^ n652 ;
  assign n655 = n643 & n654 ;
  assign n656 = n655 ^ n654 ;
  assign n642 = ~x26 & n641 ;
  assign n657 = n656 ^ n642 ;
  assign n658 = n632 & n657 ;
  assign n659 = n658 ^ n657 ;
  assign n626 = ~x25 & n625 ;
  assign n627 = ~n616 & n626 ;
  assign n615 = ~x24 & n614 ;
  assign n628 = n627 ^ n615 ;
  assign n660 = n659 ^ n628 ;
  assign n750 = n749 ^ n660 ;
  assign n761 = n760 ^ n750 ;
  assign n818 = x24 & n761 ;
  assign n1157 = n818 ^ x24 ;
  assign n816 = n614 & n761 ;
  assign n1158 = n1157 ^ n816 ;
  assign n1160 = n1158 ^ x32 ;
  assign n823 = x25 & n761 ;
  assign n1161 = n823 ^ x25 ;
  assign n821 = n625 & n761 ;
  assign n1162 = n1161 ^ n821 ;
  assign n1166 = n1162 ^ x33 ;
  assign n1167 = n1160 & n1166 ;
  assign n1168 = n1167 ^ n1160 ;
  assign n1169 = n1168 ^ n1166 ;
  assign n839 = x26 & n761 ;
  assign n1170 = n839 ^ x26 ;
  assign n837 = n641 & n761 ;
  assign n1171 = n1170 ^ n837 ;
  assign n1173 = n1171 ^ x34 ;
  assign n844 = x27 & n761 ;
  assign n1179 = n844 ^ x27 ;
  assign n842 = n652 & n761 ;
  assign n1180 = n1179 ^ n842 ;
  assign n1187 = n1180 ^ x35 ;
  assign n1188 = n1173 & n1187 ;
  assign n1189 = n1188 ^ n1173 ;
  assign n1190 = n1189 ^ n1187 ;
  assign n1191 = n1169 & n1190 ;
  assign n1192 = n1191 ^ n1169 ;
  assign n1193 = n1192 ^ n1190 ;
  assign n764 = x28 & n761 ;
  assign n1194 = n764 ^ x28 ;
  assign n762 = n605 & n761 ;
  assign n1195 = n1194 ^ n762 ;
  assign n1197 = n1195 ^ x36 ;
  assign n774 = x29 & n761 ;
  assign n1203 = n774 ^ x29 ;
  assign n772 = n678 & n761 ;
  assign n1204 = n1203 ^ n772 ;
  assign n1209 = n1204 ^ x37 ;
  assign n1210 = n1197 & n1209 ;
  assign n1211 = n1210 ^ n1197 ;
  assign n1212 = n1211 ^ n1209 ;
  assign n789 = x30 & n761 ;
  assign n1232 = n789 ^ x30 ;
  assign n787 = n751 & n761 ;
  assign n1246 = n1232 ^ n787 ;
  assign n1247 = n1246 ^ x38 ;
  assign n803 = x31 & n761 ;
  assign n1228 = n803 ^ x31 ;
  assign n801 = n721 & n761 ;
  assign n1229 = n1228 ^ n801 ;
  assign n1248 = n1229 ^ x39 ;
  assign n1249 = n1247 & n1248 ;
  assign n1250 = n1249 ^ n1247 ;
  assign n1251 = n1250 ^ n1248 ;
  assign n1252 = n1212 & n1251 ;
  assign n1253 = n1252 ^ n1212 ;
  assign n1254 = n1253 ^ n1251 ;
  assign n1255 = ~n1193 & ~n1254 ;
  assign n1237 = x30 & ~x38 ;
  assign n1238 = ~n761 & n1237 ;
  assign n1224 = x31 & x39 ;
  assign n1225 = n761 & n1224 ;
  assign n1226 = n1225 ^ n1224 ;
  assign n1222 = x39 & n721 ;
  assign n1223 = n761 & n1222 ;
  assign n1227 = n1226 ^ n1223 ;
  assign n1230 = n1229 ^ n1227 ;
  assign n1233 = n1230 & n1232 ;
  assign n1231 = n787 & n1230 ;
  assign n1234 = n1233 ^ n1231 ;
  assign n1218 = x31 & x38 ;
  assign n1219 = ~x39 & n1218 ;
  assign n1220 = ~n761 & n1219 ;
  assign n1215 = x38 & ~x39 ;
  assign n1216 = n721 & n1215 ;
  assign n1217 = n761 & n1216 ;
  assign n1221 = n1220 ^ n1217 ;
  assign n1235 = n1234 ^ n1221 ;
  assign n1236 = n1235 ^ n1230 ;
  assign n1239 = n1238 ^ n1236 ;
  assign n1213 = ~x38 & n751 ;
  assign n1214 = n761 & n1213 ;
  assign n1240 = n1239 ^ n1214 ;
  assign n1241 = n1212 & n1240 ;
  assign n1242 = n1241 ^ n1240 ;
  assign n1200 = x29 & x37 ;
  assign n1201 = ~n761 & n1200 ;
  assign n1198 = x37 & n678 ;
  assign n1199 = n761 & n1198 ;
  assign n1202 = n1201 ^ n1199 ;
  assign n1205 = n1204 ^ n1202 ;
  assign n1206 = n1197 & n1205 ;
  assign n1207 = n1206 ^ n1205 ;
  assign n1196 = ~x36 & n1195 ;
  assign n1208 = n1207 ^ n1196 ;
  assign n1243 = n1242 ^ n1208 ;
  assign n1244 = ~n1193 & n1243 ;
  assign n1176 = x27 & x35 ;
  assign n1177 = ~n761 & n1176 ;
  assign n1174 = x35 & n652 ;
  assign n1175 = n761 & n1174 ;
  assign n1178 = n1177 ^ n1175 ;
  assign n1181 = n1180 ^ n1178 ;
  assign n1182 = n1173 & n1181 ;
  assign n1183 = n1182 ^ n1181 ;
  assign n1172 = ~x34 & n1171 ;
  assign n1184 = n1183 ^ n1172 ;
  assign n1185 = ~n1169 & n1184 ;
  assign n1163 = ~x33 & n1162 ;
  assign n1164 = ~n1160 & n1163 ;
  assign n1159 = ~x32 & n1158 ;
  assign n1165 = n1164 ^ n1159 ;
  assign n1186 = n1185 ^ n1165 ;
  assign n1245 = n1244 ^ n1186 ;
  assign n1256 = n1255 ^ n1245 ;
  assign n1259 = x32 & n1256 ;
  assign n1859 = n1259 ^ x32 ;
  assign n1257 = n1158 & n1256 ;
  assign n1860 = n1859 ^ n1257 ;
  assign n1862 = n1860 ^ x40 ;
  assign n1267 = x33 & n1256 ;
  assign n1863 = n1267 ^ x33 ;
  assign n1265 = n1162 & n1256 ;
  assign n1864 = n1863 ^ n1265 ;
  assign n1868 = n1864 ^ x41 ;
  assign n1869 = n1862 & n1868 ;
  assign n1870 = n1869 ^ n1862 ;
  assign n1871 = n1870 ^ n1868 ;
  assign n1277 = x34 & n1256 ;
  assign n1872 = n1277 ^ x34 ;
  assign n1275 = n1171 & n1256 ;
  assign n1873 = n1872 ^ n1275 ;
  assign n1875 = n1873 ^ x42 ;
  assign n1283 = x35 & n1256 ;
  assign n1885 = n1283 ^ x35 ;
  assign n1281 = n1180 & n1256 ;
  assign n1886 = n1885 ^ n1281 ;
  assign n1887 = n1886 ^ x43 ;
  assign n1888 = n1875 & n1887 ;
  assign n1889 = n1888 ^ n1875 ;
  assign n1890 = n1889 ^ n1887 ;
  assign n1891 = ~n1871 & ~n1890 ;
  assign n1308 = x36 & n1256 ;
  assign n1857 = n1308 ^ x36 ;
  assign n1306 = n1195 & n1256 ;
  assign n1858 = n1857 ^ n1306 ;
  assign n1893 = n1858 ^ x44 ;
  assign n1315 = x37 & n1256 ;
  assign n1901 = n1315 ^ x37 ;
  assign n1313 = n1204 & n1256 ;
  assign n1902 = n1901 ^ n1313 ;
  assign n1903 = n1902 ^ x45 ;
  assign n1904 = n1893 & n1903 ;
  assign n1905 = n1904 ^ n1893 ;
  assign n1906 = n1905 ^ n1903 ;
  assign n1325 = x38 & n1256 ;
  assign n1940 = n1325 ^ x38 ;
  assign n1323 = n1246 & n1256 ;
  assign n1941 = n1940 ^ n1323 ;
  assign n1942 = n1941 ^ x46 ;
  assign n1334 = x39 & n1256 ;
  assign n1922 = n1334 ^ x39 ;
  assign n1332 = n1229 & n1256 ;
  assign n1923 = n1922 ^ n1332 ;
  assign n1943 = n1923 ^ x47 ;
  assign n1944 = n1942 & n1943 ;
  assign n1945 = n1944 ^ n1942 ;
  assign n1946 = n1945 ^ n1943 ;
  assign n1947 = ~n1906 & ~n1946 ;
  assign n1948 = n1891 & n1947 ;
  assign n1932 = x38 & ~x46 ;
  assign n1933 = ~n1256 & n1932 ;
  assign n1926 = x38 & x39 ;
  assign n1927 = ~x47 & n1926 ;
  assign n1928 = ~n1256 & n1927 ;
  assign n1918 = x39 & x47 ;
  assign n1919 = n1256 & n1918 ;
  assign n1920 = n1919 ^ n1918 ;
  assign n1916 = x47 & n1229 ;
  assign n1917 = n1256 & n1916 ;
  assign n1921 = n1920 ^ n1917 ;
  assign n1924 = n1923 ^ n1921 ;
  assign n1925 = n1323 & n1924 ;
  assign n1929 = n1928 ^ n1925 ;
  assign n1912 = x39 & x46 ;
  assign n1913 = ~x47 & n1912 ;
  assign n1914 = ~n1256 & n1913 ;
  assign n1909 = x46 & ~x47 ;
  assign n1910 = n1229 & n1909 ;
  assign n1911 = n1256 & n1910 ;
  assign n1915 = n1914 ^ n1911 ;
  assign n1930 = n1929 ^ n1915 ;
  assign n1931 = n1930 ^ n1924 ;
  assign n1934 = n1933 ^ n1931 ;
  assign n1907 = ~x46 & n1246 ;
  assign n1908 = n1256 & n1907 ;
  assign n1935 = n1934 ^ n1908 ;
  assign n1936 = ~n1906 & n1935 ;
  assign n1896 = x37 & ~x45 ;
  assign n1897 = ~n1256 & n1896 ;
  assign n1894 = ~x45 & n1204 ;
  assign n1895 = n1256 & n1894 ;
  assign n1898 = n1897 ^ n1895 ;
  assign n1899 = ~n1893 & n1898 ;
  assign n1892 = ~x44 & n1858 ;
  assign n1900 = n1899 ^ n1892 ;
  assign n1937 = n1936 ^ n1900 ;
  assign n1938 = n1891 & n1937 ;
  assign n1878 = x35 & ~x43 ;
  assign n1879 = ~n1256 & n1878 ;
  assign n1876 = ~x43 & n1180 ;
  assign n1877 = n1256 & n1876 ;
  assign n1880 = n1879 ^ n1877 ;
  assign n1881 = ~n1875 & n1880 ;
  assign n1874 = ~x42 & n1873 ;
  assign n1882 = n1881 ^ n1874 ;
  assign n1883 = ~n1871 & n1882 ;
  assign n1865 = ~x41 & n1864 ;
  assign n1866 = ~n1862 & n1865 ;
  assign n1861 = ~x40 & n1860 ;
  assign n1867 = n1866 ^ n1861 ;
  assign n1884 = n1883 ^ n1867 ;
  assign n1939 = n1938 ^ n1884 ;
  assign n1949 = n1948 ^ n1939 ;
  assign n2055 = x42 & n1949 ;
  assign n2053 = n1873 & n1949 ;
  assign n2054 = n2053 ^ n1873 ;
  assign n2056 = n2055 ^ n2054 ;
  assign n1258 = n1257 ^ n1158 ;
  assign n1260 = n1259 ^ n1258 ;
  assign n838 = n837 ^ n641 ;
  assign n840 = n839 ^ n838 ;
  assign n86 = ~n53 & n85 ;
  assign n91 = n90 ^ n86 ;
  assign n81 = ~n61 & n80 ;
  assign n92 = n91 ^ n81 ;
  assign n101 = n100 ^ n92 ;
  assign n377 = x10 & n101 ;
  assign n376 = x2 & ~n101 ;
  assign n378 = n377 ^ n376 ;
  assign n332 = x16 & ~n151 ;
  assign n335 = n334 ^ n332 ;
  assign n338 = n337 ^ n335 ;
  assign n341 = n340 ^ n338 ;
  assign n152 = n125 & n151 ;
  assign n206 = n205 ^ n152 ;
  assign n315 = n314 ^ n206 ;
  assign n331 = n330 ^ n315 ;
  assign n342 = n341 ^ n331 ;
  assign n103 = x8 & n101 ;
  assign n102 = x0 & ~n101 ;
  assign n104 = n103 ^ n102 ;
  assign n344 = n342 ^ n104 ;
  assign n358 = x17 & ~n151 ;
  assign n361 = n360 ^ n358 ;
  assign n364 = n363 ^ n361 ;
  assign n367 = n366 ^ n364 ;
  assign n348 = n148 & n151 ;
  assign n351 = n350 ^ n348 ;
  assign n354 = n353 ^ n351 ;
  assign n357 = n356 ^ n354 ;
  assign n368 = n367 ^ n357 ;
  assign n346 = x9 & n101 ;
  assign n345 = x1 & ~n101 ;
  assign n347 = n346 ^ n345 ;
  assign n372 = n368 ^ n347 ;
  assign n373 = n344 & n372 ;
  assign n374 = n373 ^ n344 ;
  assign n375 = n374 ^ n372 ;
  assign n389 = x18 & ~n151 ;
  assign n392 = n391 ^ n389 ;
  assign n395 = n394 ^ n392 ;
  assign n398 = n397 ^ n395 ;
  assign n379 = n151 & n173 ;
  assign n382 = n381 ^ n379 ;
  assign n385 = n384 ^ n382 ;
  assign n388 = n387 ^ n385 ;
  assign n399 = n398 ^ n388 ;
  assign n401 = n399 ^ n378 ;
  assign n424 = x11 & n101 ;
  assign n423 = x3 & ~n101 ;
  assign n425 = n424 ^ n423 ;
  assign n412 = x19 & ~n151 ;
  assign n415 = n414 ^ n412 ;
  assign n418 = n417 ^ n415 ;
  assign n421 = n420 ^ n418 ;
  assign n402 = n151 & n196 ;
  assign n405 = n404 ^ n402 ;
  assign n408 = n407 ^ n405 ;
  assign n411 = n410 ^ n408 ;
  assign n422 = n421 ^ n411 ;
  assign n434 = n425 ^ n422 ;
  assign n435 = n401 & n434 ;
  assign n436 = n435 ^ n401 ;
  assign n437 = n436 ^ n434 ;
  assign n438 = n375 & n437 ;
  assign n439 = n438 ^ n375 ;
  assign n440 = n439 ^ n437 ;
  assign n463 = x12 & n101 ;
  assign n462 = x4 & ~n101 ;
  assign n464 = n463 ^ n462 ;
  assign n451 = x20 & ~n151 ;
  assign n454 = n453 ^ n451 ;
  assign n457 = n456 ^ n454 ;
  assign n460 = n459 ^ n457 ;
  assign n441 = n151 & n234 ;
  assign n444 = n443 ^ n441 ;
  assign n447 = n446 ^ n444 ;
  assign n450 = n449 ^ n447 ;
  assign n461 = n460 ^ n450 ;
  assign n466 = n464 ^ n461 ;
  assign n489 = x13 & n101 ;
  assign n488 = x5 & ~n101 ;
  assign n490 = n489 ^ n488 ;
  assign n477 = x21 & ~n151 ;
  assign n480 = n479 ^ n477 ;
  assign n483 = n482 ^ n480 ;
  assign n486 = n485 ^ n483 ;
  assign n467 = n151 & n256 ;
  assign n470 = n469 ^ n467 ;
  assign n473 = n472 ^ n470 ;
  assign n476 = n475 ^ n473 ;
  assign n487 = n486 ^ n476 ;
  assign n496 = n490 ^ n487 ;
  assign n497 = n466 & n496 ;
  assign n498 = n497 ^ n466 ;
  assign n499 = n498 ^ n496 ;
  assign n522 = x14 & n101 ;
  assign n521 = x6 & ~n101 ;
  assign n523 = n522 ^ n521 ;
  assign n510 = x22 & ~n151 ;
  assign n513 = n512 ^ n510 ;
  assign n516 = n515 ^ n513 ;
  assign n519 = n518 ^ n516 ;
  assign n500 = n151 & n281 ;
  assign n503 = n502 ^ n500 ;
  assign n506 = n505 ^ n503 ;
  assign n509 = n508 ^ n506 ;
  assign n520 = n519 ^ n509 ;
  assign n526 = n523 ^ n520 ;
  assign n573 = n572 ^ n304 ;
  assign n584 = n583 ^ n573 ;
  assign n527 = x7 & ~n91 ;
  assign n528 = n527 ^ n296 ;
  assign n529 = n528 ^ n295 ;
  assign n530 = n529 ^ n292 ;
  assign n585 = n584 ^ n530 ;
  assign n586 = n526 & n585 ;
  assign n587 = n586 ^ n526 ;
  assign n588 = n587 ^ n585 ;
  assign n589 = n499 & n588 ;
  assign n590 = n589 ^ n499 ;
  assign n591 = n590 ^ n588 ;
  assign n592 = ~n440 & ~n591 ;
  assign n542 = x23 & n530 ;
  assign n548 = ~n203 & n542 ;
  assign n549 = n199 & n548 ;
  assign n547 = ~n151 & n542 ;
  assign n550 = n549 ^ n547 ;
  assign n545 = n312 & n542 ;
  assign n546 = n545 ^ n542 ;
  assign n551 = n550 ^ n546 ;
  assign n543 = ~n213 & n542 ;
  assign n544 = n329 & n543 ;
  assign n552 = n551 ^ n544 ;
  assign n531 = n304 & n530 ;
  assign n537 = ~n203 & n531 ;
  assign n538 = n199 & n537 ;
  assign n536 = n151 & n531 ;
  assign n539 = n538 ^ n536 ;
  assign n534 = n312 & n531 ;
  assign n535 = n534 ^ n531 ;
  assign n540 = n539 ^ n535 ;
  assign n532 = ~n213 & n531 ;
  assign n533 = n329 & n532 ;
  assign n541 = n540 ^ n533 ;
  assign n553 = n552 ^ n541 ;
  assign n554 = n553 ^ n530 ;
  assign n555 = n526 & n554 ;
  assign n556 = n555 ^ n554 ;
  assign n524 = n520 & n523 ;
  assign n525 = n524 ^ n523 ;
  assign n557 = n556 ^ n525 ;
  assign n558 = n499 & n557 ;
  assign n559 = n558 ^ n557 ;
  assign n491 = n487 & n490 ;
  assign n492 = n491 ^ n490 ;
  assign n493 = n466 & n492 ;
  assign n494 = n493 ^ n492 ;
  assign n465 = ~n461 & n464 ;
  assign n495 = n494 ^ n465 ;
  assign n560 = n559 ^ n495 ;
  assign n561 = ~n440 & n560 ;
  assign n426 = n422 & n425 ;
  assign n427 = n426 ^ n425 ;
  assign n428 = n401 & n427 ;
  assign n429 = n428 ^ n427 ;
  assign n400 = n378 & ~n399 ;
  assign n430 = n429 ^ n400 ;
  assign n431 = n375 & n430 ;
  assign n432 = n431 ^ n430 ;
  assign n369 = n347 & ~n368 ;
  assign n370 = ~n344 & n369 ;
  assign n343 = n104 & ~n342 ;
  assign n371 = n370 ^ n343 ;
  assign n433 = n432 ^ n371 ;
  assign n562 = n561 ^ n433 ;
  assign n593 = n592 ^ n562 ;
  assign n835 = n378 & n593 ;
  assign n833 = n399 & n593 ;
  assign n834 = n833 ^ n399 ;
  assign n836 = n835 ^ n834 ;
  assign n841 = n840 ^ n836 ;
  assign n843 = n842 ^ n652 ;
  assign n845 = n844 ^ n843 ;
  assign n848 = n425 & n593 ;
  assign n846 = n422 & n593 ;
  assign n847 = n846 ^ n422 ;
  assign n849 = n848 ^ n847 ;
  assign n875 = n845 & n849 ;
  assign n876 = n875 ^ n849 ;
  assign n877 = n841 & n876 ;
  assign n878 = n877 ^ n876 ;
  assign n874 = n836 & ~n840 ;
  assign n879 = n878 ^ n874 ;
  assign n817 = n816 ^ n614 ;
  assign n819 = n818 ^ n817 ;
  assign n814 = n104 & n593 ;
  assign n595 = n342 & n593 ;
  assign n813 = n595 ^ n342 ;
  assign n815 = n814 ^ n813 ;
  assign n820 = n819 ^ n815 ;
  assign n827 = n347 & n593 ;
  assign n825 = n368 & n593 ;
  assign n826 = n825 ^ n368 ;
  assign n828 = n827 ^ n826 ;
  assign n822 = n821 ^ n625 ;
  assign n824 = n823 ^ n822 ;
  assign n829 = n828 ^ n824 ;
  assign n830 = n820 & n829 ;
  assign n831 = n830 ^ n820 ;
  assign n832 = n831 ^ n829 ;
  assign n891 = n819 & ~n832 ;
  assign n892 = n879 & n891 ;
  assign n870 = ~n824 & n828 ;
  assign n871 = ~n820 & n870 ;
  assign n869 = n815 & ~n819 ;
  assign n872 = n871 ^ n869 ;
  assign n890 = n819 & ~n872 ;
  assign n893 = n892 ^ n890 ;
  assign n850 = n849 ^ n845 ;
  assign n851 = n841 & n850 ;
  assign n852 = n851 ^ n841 ;
  assign n853 = n852 ^ n850 ;
  assign n854 = n832 & n853 ;
  assign n855 = n854 ^ n832 ;
  assign n856 = n855 ^ n853 ;
  assign n768 = n464 & n593 ;
  assign n766 = n461 & n593 ;
  assign n767 = n766 ^ n461 ;
  assign n769 = n768 ^ n767 ;
  assign n763 = n762 ^ n605 ;
  assign n765 = n764 ^ n763 ;
  assign n771 = n769 ^ n765 ;
  assign n778 = n490 & n593 ;
  assign n776 = n487 & n593 ;
  assign n777 = n776 ^ n487 ;
  assign n779 = n778 ^ n777 ;
  assign n773 = n772 ^ n678 ;
  assign n775 = n774 ^ n773 ;
  assign n783 = n779 ^ n775 ;
  assign n784 = n771 & n783 ;
  assign n785 = n784 ^ n771 ;
  assign n786 = n785 ^ n783 ;
  assign n793 = n523 & n593 ;
  assign n791 = n520 & n593 ;
  assign n792 = n791 ^ n520 ;
  assign n794 = n793 ^ n792 ;
  assign n788 = n787 ^ n751 ;
  assign n790 = n789 ^ n788 ;
  assign n796 = n794 ^ n790 ;
  assign n802 = n801 ^ n721 ;
  assign n804 = n803 ^ n802 ;
  assign n799 = n530 & n593 ;
  assign n797 = n584 & n593 ;
  assign n798 = n797 ^ n584 ;
  assign n800 = n799 ^ n798 ;
  assign n859 = n804 ^ n800 ;
  assign n860 = n796 & n859 ;
  assign n861 = n860 ^ n796 ;
  assign n862 = n861 ^ n859 ;
  assign n863 = n786 & n862 ;
  assign n864 = n863 ^ n786 ;
  assign n865 = n864 ^ n862 ;
  assign n866 = ~n856 & ~n865 ;
  assign n888 = n819 & n866 ;
  assign n889 = n888 ^ n819 ;
  assign n894 = n893 ^ n889 ;
  assign n805 = n800 & n804 ;
  assign n806 = n805 ^ n800 ;
  assign n807 = n796 & n806 ;
  assign n808 = n807 ^ n806 ;
  assign n795 = ~n790 & n794 ;
  assign n809 = n808 ^ n795 ;
  assign n810 = n786 & n809 ;
  assign n811 = n810 ^ n809 ;
  assign n780 = ~n775 & n779 ;
  assign n781 = ~n771 & n780 ;
  assign n770 = ~n765 & n769 ;
  assign n782 = n781 ^ n770 ;
  assign n812 = n811 ^ n782 ;
  assign n886 = n819 & ~n856 ;
  assign n887 = n812 & n886 ;
  assign n895 = n894 ^ n887 ;
  assign n1155 = n895 ^ n819 ;
  assign n880 = n815 & ~n832 ;
  assign n881 = n879 & n880 ;
  assign n873 = n815 & ~n872 ;
  assign n882 = n881 ^ n873 ;
  assign n867 = n815 & n866 ;
  assign n868 = n867 ^ n815 ;
  assign n883 = n882 ^ n868 ;
  assign n857 = n815 & ~n856 ;
  assign n858 = n812 & n857 ;
  assign n884 = n883 ^ n858 ;
  assign n1156 = n1155 ^ n884 ;
  assign n1262 = n1260 ^ n1156 ;
  assign n917 = n824 & ~n832 ;
  assign n918 = n879 & n917 ;
  assign n916 = n824 & ~n872 ;
  assign n919 = n918 ^ n916 ;
  assign n914 = n824 & n866 ;
  assign n915 = n914 ^ n824 ;
  assign n920 = n919 ^ n915 ;
  assign n912 = n824 & ~n856 ;
  assign n913 = n812 & n912 ;
  assign n921 = n920 ^ n913 ;
  assign n1263 = n921 ^ n824 ;
  assign n906 = n828 & ~n832 ;
  assign n907 = n879 & n906 ;
  assign n905 = n828 & ~n872 ;
  assign n908 = n907 ^ n905 ;
  assign n903 = n828 & n866 ;
  assign n904 = n903 ^ n828 ;
  assign n909 = n908 ^ n904 ;
  assign n901 = n828 & ~n856 ;
  assign n902 = n812 & n901 ;
  assign n910 = n909 ^ n902 ;
  assign n1264 = n1263 ^ n910 ;
  assign n1266 = n1265 ^ n1162 ;
  assign n1268 = n1267 ^ n1266 ;
  assign n1269 = n1264 & ~n1268 ;
  assign n1270 = ~n1262 & n1269 ;
  assign n1261 = n1156 & ~n1260 ;
  assign n1271 = n1270 ^ n1261 ;
  assign n946 = ~n832 & n840 ;
  assign n947 = n879 & n946 ;
  assign n945 = n840 & ~n872 ;
  assign n948 = n947 ^ n945 ;
  assign n943 = n840 & n866 ;
  assign n944 = n943 ^ n840 ;
  assign n949 = n948 ^ n944 ;
  assign n941 = n840 & ~n856 ;
  assign n942 = n812 & n941 ;
  assign n950 = n949 ^ n942 ;
  assign n1273 = n950 ^ n840 ;
  assign n935 = ~n832 & n836 ;
  assign n936 = n879 & n935 ;
  assign n934 = n836 & ~n872 ;
  assign n937 = n936 ^ n934 ;
  assign n932 = n836 & n866 ;
  assign n933 = n932 ^ n836 ;
  assign n938 = n937 ^ n933 ;
  assign n930 = n836 & ~n856 ;
  assign n931 = n812 & n930 ;
  assign n939 = n938 ^ n931 ;
  assign n1274 = n1273 ^ n939 ;
  assign n2048 = ~n1271 & n1274 ;
  assign n1276 = n1275 ^ n1171 ;
  assign n1278 = n1277 ^ n1276 ;
  assign n1280 = n1278 ^ n1274 ;
  assign n1282 = n1281 ^ n1180 ;
  assign n1284 = n1283 ^ n1282 ;
  assign n972 = ~n832 & n845 ;
  assign n973 = n879 & n972 ;
  assign n971 = n845 & ~n872 ;
  assign n974 = n973 ^ n971 ;
  assign n969 = n845 & n866 ;
  assign n970 = n969 ^ n845 ;
  assign n975 = n974 ^ n970 ;
  assign n967 = n845 & ~n856 ;
  assign n968 = n812 & n967 ;
  assign n976 = n975 ^ n968 ;
  assign n1285 = n976 ^ n845 ;
  assign n961 = ~n832 & n849 ;
  assign n962 = n879 & n961 ;
  assign n960 = n849 & ~n872 ;
  assign n963 = n962 ^ n960 ;
  assign n958 = n849 & n866 ;
  assign n959 = n958 ^ n849 ;
  assign n964 = n963 ^ n959 ;
  assign n956 = n849 & ~n856 ;
  assign n957 = n812 & n956 ;
  assign n965 = n964 ^ n957 ;
  assign n1286 = n1285 ^ n965 ;
  assign n1287 = n1284 & n1286 ;
  assign n1288 = n1287 ^ n1286 ;
  assign n1289 = n1280 & n1288 ;
  assign n1290 = n1289 ^ n1288 ;
  assign n1279 = n1274 & ~n1278 ;
  assign n1291 = n1290 ^ n1279 ;
  assign n1292 = n1268 ^ n1264 ;
  assign n1293 = n1262 & n1292 ;
  assign n1294 = n1293 ^ n1262 ;
  assign n1295 = n1294 ^ n1292 ;
  assign n1409 = n1274 & ~n1295 ;
  assign n1410 = n1291 & n1409 ;
  assign n2049 = n2048 ^ n1410 ;
  assign n1299 = n1286 ^ n1284 ;
  assign n1300 = n1280 & n1299 ;
  assign n1301 = n1300 ^ n1280 ;
  assign n1302 = n1301 ^ n1299 ;
  assign n1303 = n1295 & n1302 ;
  assign n1304 = n1303 ^ n1295 ;
  assign n1305 = n1304 ^ n1302 ;
  assign n1011 = n765 & ~n832 ;
  assign n1012 = n879 & n1011 ;
  assign n1010 = n765 & ~n872 ;
  assign n1013 = n1012 ^ n1010 ;
  assign n1008 = n765 & n866 ;
  assign n1009 = n1008 ^ n765 ;
  assign n1014 = n1013 ^ n1009 ;
  assign n1006 = n765 & ~n856 ;
  assign n1007 = n812 & n1006 ;
  assign n1015 = n1014 ^ n1007 ;
  assign n1310 = n1015 ^ n765 ;
  assign n1000 = n769 & ~n832 ;
  assign n1001 = n879 & n1000 ;
  assign n999 = n769 & ~n872 ;
  assign n1002 = n1001 ^ n999 ;
  assign n997 = n769 & n866 ;
  assign n998 = n997 ^ n769 ;
  assign n1003 = n1002 ^ n998 ;
  assign n995 = n769 & ~n856 ;
  assign n996 = n812 & n995 ;
  assign n1004 = n1003 ^ n996 ;
  assign n1311 = n1310 ^ n1004 ;
  assign n1307 = n1306 ^ n1195 ;
  assign n1309 = n1308 ^ n1307 ;
  assign n1312 = n1311 ^ n1309 ;
  assign n1037 = n775 & ~n832 ;
  assign n1038 = n879 & n1037 ;
  assign n1036 = n775 & ~n872 ;
  assign n1039 = n1038 ^ n1036 ;
  assign n1034 = n775 & n866 ;
  assign n1035 = n1034 ^ n775 ;
  assign n1040 = n1039 ^ n1035 ;
  assign n1032 = n775 & ~n856 ;
  assign n1033 = n812 & n1032 ;
  assign n1041 = n1040 ^ n1033 ;
  assign n1317 = n1041 ^ n775 ;
  assign n1026 = n779 & ~n832 ;
  assign n1027 = n879 & n1026 ;
  assign n1025 = n779 & ~n872 ;
  assign n1028 = n1027 ^ n1025 ;
  assign n1023 = n779 & n866 ;
  assign n1024 = n1023 ^ n779 ;
  assign n1029 = n1028 ^ n1024 ;
  assign n1021 = n779 & ~n856 ;
  assign n1022 = n812 & n1021 ;
  assign n1030 = n1029 ^ n1022 ;
  assign n1318 = n1317 ^ n1030 ;
  assign n1314 = n1313 ^ n1204 ;
  assign n1316 = n1315 ^ n1314 ;
  assign n1319 = n1318 ^ n1316 ;
  assign n1320 = n1312 & n1319 ;
  assign n1321 = n1320 ^ n1312 ;
  assign n1322 = n1321 ^ n1319 ;
  assign n1070 = n790 & ~n832 ;
  assign n1071 = n879 & n1070 ;
  assign n1069 = n790 & ~n872 ;
  assign n1072 = n1071 ^ n1069 ;
  assign n1067 = n790 & n866 ;
  assign n1068 = n1067 ^ n790 ;
  assign n1073 = n1072 ^ n1068 ;
  assign n1065 = n790 & ~n856 ;
  assign n1066 = n812 & n1065 ;
  assign n1074 = n1073 ^ n1066 ;
  assign n1327 = n1074 ^ n790 ;
  assign n1059 = n794 & ~n832 ;
  assign n1060 = n879 & n1059 ;
  assign n1058 = n794 & ~n872 ;
  assign n1061 = n1060 ^ n1058 ;
  assign n1056 = n794 & n866 ;
  assign n1057 = n1056 ^ n794 ;
  assign n1062 = n1061 ^ n1057 ;
  assign n1054 = n794 & ~n856 ;
  assign n1055 = n812 & n1054 ;
  assign n1063 = n1062 ^ n1055 ;
  assign n1328 = n1327 ^ n1063 ;
  assign n1324 = n1323 ^ n1246 ;
  assign n1326 = n1325 ^ n1324 ;
  assign n1329 = n1328 ^ n1326 ;
  assign n1333 = n1332 ^ n1229 ;
  assign n1335 = n1334 ^ n1333 ;
  assign n1133 = n804 & ~n832 ;
  assign n1134 = n879 & n1133 ;
  assign n1132 = n804 & n872 ;
  assign n1135 = n1134 ^ n1132 ;
  assign n1136 = n1135 ^ n804 ;
  assign n1130 = n804 & n866 ;
  assign n1131 = n1130 ^ n804 ;
  assign n1137 = n1136 ^ n1131 ;
  assign n1128 = n804 & ~n856 ;
  assign n1129 = n812 & n1128 ;
  assign n1138 = n1137 ^ n1129 ;
  assign n1330 = n1138 ^ n804 ;
  assign n1121 = n800 & ~n832 ;
  assign n1122 = n879 & n1121 ;
  assign n1120 = n800 & n872 ;
  assign n1123 = n1122 ^ n1120 ;
  assign n1124 = n1123 ^ n800 ;
  assign n1118 = n800 & n866 ;
  assign n1119 = n1118 ^ n800 ;
  assign n1125 = n1124 ^ n1119 ;
  assign n1116 = n800 & ~n856 ;
  assign n1117 = n812 & n1116 ;
  assign n1126 = n1125 ^ n1117 ;
  assign n1331 = n1330 ^ n1126 ;
  assign n1336 = n1335 ^ n1331 ;
  assign n1337 = n1329 & n1336 ;
  assign n1338 = n1337 ^ n1329 ;
  assign n1339 = n1338 ^ n1336 ;
  assign n1340 = n1322 & n1339 ;
  assign n1341 = n1340 ^ n1322 ;
  assign n1342 = n1341 ^ n1339 ;
  assign n1343 = ~n1305 & ~n1342 ;
  assign n1412 = n1274 & n1343 ;
  assign n1413 = n1412 ^ n1274 ;
  assign n2050 = n2049 ^ n1413 ;
  assign n1355 = n1331 & n1335 ;
  assign n1356 = n1355 ^ n1331 ;
  assign n1357 = n1329 & n1356 ;
  assign n1358 = n1357 ^ n1356 ;
  assign n1353 = n1326 & n1328 ;
  assign n1354 = n1353 ^ n1328 ;
  assign n1359 = n1358 ^ n1354 ;
  assign n1360 = n1322 & n1359 ;
  assign n1361 = n1360 ^ n1359 ;
  assign n1348 = n1316 & n1318 ;
  assign n1349 = n1348 ^ n1318 ;
  assign n1350 = n1312 & n1349 ;
  assign n1351 = n1350 ^ n1349 ;
  assign n1347 = ~n1309 & n1311 ;
  assign n1352 = n1351 ^ n1347 ;
  assign n1362 = n1361 ^ n1352 ;
  assign n1415 = n1274 & ~n1305 ;
  assign n1416 = n1362 & n1415 ;
  assign n2051 = n2050 ^ n1416 ;
  assign n2044 = n1271 & n1278 ;
  assign n1419 = n1278 & ~n1295 ;
  assign n1420 = n1291 & n1419 ;
  assign n2045 = n2044 ^ n1420 ;
  assign n1422 = n1278 & n1343 ;
  assign n1423 = n1422 ^ n1278 ;
  assign n2046 = n2045 ^ n1423 ;
  assign n1425 = n1278 & ~n1305 ;
  assign n1426 = n1362 & n1425 ;
  assign n2047 = n2046 ^ n1426 ;
  assign n2052 = n2051 ^ n2047 ;
  assign n2057 = n2056 ^ n2052 ;
  assign n2060 = x43 & n1949 ;
  assign n2058 = n1886 & n1949 ;
  assign n2059 = n2058 ^ n1886 ;
  assign n2061 = n2060 ^ n2059 ;
  assign n2066 = ~n1271 & n1286 ;
  assign n1440 = n1286 & ~n1295 ;
  assign n1441 = n1291 & n1440 ;
  assign n2067 = n2066 ^ n1441 ;
  assign n1443 = n1286 & n1343 ;
  assign n1444 = n1443 ^ n1286 ;
  assign n2068 = n2067 ^ n1444 ;
  assign n1446 = n1286 & ~n1305 ;
  assign n1447 = n1362 & n1446 ;
  assign n2069 = n2068 ^ n1447 ;
  assign n2062 = n1271 & n1284 ;
  assign n1450 = n1284 & ~n1295 ;
  assign n1451 = n1291 & n1450 ;
  assign n2063 = n2062 ^ n1451 ;
  assign n1453 = n1284 & n1343 ;
  assign n1454 = n1453 ^ n1284 ;
  assign n2064 = n2063 ^ n1454 ;
  assign n1456 = n1284 & ~n1305 ;
  assign n1457 = n1362 & n1456 ;
  assign n2065 = n2064 ^ n1457 ;
  assign n2070 = n2069 ^ n2065 ;
  assign n2092 = ~n2061 & n2070 ;
  assign n2093 = ~n2057 & n2092 ;
  assign n2091 = n2052 & ~n2056 ;
  assign n2094 = n2093 ^ n2091 ;
  assign n2024 = x40 & n1949 ;
  assign n2022 = n1860 & n1949 ;
  assign n2023 = n2022 ^ n1860 ;
  assign n2025 = n2024 ^ n2023 ;
  assign n2017 = n1156 & ~n1271 ;
  assign n1296 = n1156 & ~n1295 ;
  assign n1297 = n1291 & n1296 ;
  assign n2018 = n2017 ^ n1297 ;
  assign n1344 = n1156 & n1343 ;
  assign n1345 = n1344 ^ n1156 ;
  assign n2019 = n2018 ^ n1345 ;
  assign n1363 = n1156 & ~n1305 ;
  assign n1364 = n1362 & n1363 ;
  assign n2020 = n2019 ^ n1364 ;
  assign n2013 = n1260 & n1271 ;
  assign n1367 = n1260 & ~n1295 ;
  assign n1368 = n1291 & n1367 ;
  assign n2014 = n2013 ^ n1368 ;
  assign n1370 = n1260 & n1343 ;
  assign n1371 = n1370 ^ n1260 ;
  assign n2015 = n2014 ^ n1371 ;
  assign n1373 = n1260 & ~n1305 ;
  assign n1374 = n1362 & n1373 ;
  assign n2016 = n2015 ^ n1374 ;
  assign n2021 = n2020 ^ n2016 ;
  assign n2026 = n2025 ^ n2021 ;
  assign n2038 = x41 & n1949 ;
  assign n2036 = n1864 & n1949 ;
  assign n2037 = n2036 ^ n1864 ;
  assign n2039 = n2038 ^ n2037 ;
  assign n2031 = n1264 & ~n1271 ;
  assign n1380 = n1264 & ~n1295 ;
  assign n1381 = n1291 & n1380 ;
  assign n2032 = n2031 ^ n1381 ;
  assign n1383 = n1264 & n1343 ;
  assign n1384 = n1383 ^ n1264 ;
  assign n2033 = n2032 ^ n1384 ;
  assign n1386 = n1264 & ~n1305 ;
  assign n1387 = n1362 & n1386 ;
  assign n2034 = n2033 ^ n1387 ;
  assign n2027 = n1268 & n1271 ;
  assign n1390 = n1268 & ~n1295 ;
  assign n1391 = n1291 & n1390 ;
  assign n2028 = n2027 ^ n1391 ;
  assign n1393 = n1268 & n1343 ;
  assign n1394 = n1393 ^ n1268 ;
  assign n2029 = n2028 ^ n1394 ;
  assign n1396 = n1268 & ~n1305 ;
  assign n1397 = n1362 & n1396 ;
  assign n2030 = n2029 ^ n1397 ;
  assign n2035 = n2034 ^ n2030 ;
  assign n2040 = n2039 ^ n2035 ;
  assign n2041 = n2026 & n2040 ;
  assign n2042 = n2041 ^ n2026 ;
  assign n2043 = n2042 ^ n2040 ;
  assign n2246 = n2025 & ~n2043 ;
  assign n2247 = n2094 & n2246 ;
  assign n2087 = n2035 & ~n2039 ;
  assign n2088 = ~n2026 & n2087 ;
  assign n2086 = n2021 & ~n2025 ;
  assign n2089 = n2088 ^ n2086 ;
  assign n2245 = n2025 & ~n2089 ;
  assign n2248 = n2247 ^ n2245 ;
  assign n2071 = n2070 ^ n2061 ;
  assign n2072 = n2057 & n2071 ;
  assign n2073 = n2072 ^ n2057 ;
  assign n2074 = n2073 ^ n2071 ;
  assign n2075 = ~n2043 & ~n2074 ;
  assign n1958 = ~n1271 & n1311 ;
  assign n1480 = ~n1295 & n1311 ;
  assign n1481 = n1291 & n1480 ;
  assign n1959 = n1958 ^ n1481 ;
  assign n1483 = n1311 & n1343 ;
  assign n1484 = n1483 ^ n1311 ;
  assign n1960 = n1959 ^ n1484 ;
  assign n1486 = ~n1305 & n1311 ;
  assign n1487 = n1362 & n1486 ;
  assign n1961 = n1960 ^ n1487 ;
  assign n1954 = n1271 & n1309 ;
  assign n1490 = ~n1295 & n1309 ;
  assign n1491 = n1291 & n1490 ;
  assign n1955 = n1954 ^ n1491 ;
  assign n1493 = n1309 & n1343 ;
  assign n1494 = n1493 ^ n1309 ;
  assign n1956 = n1955 ^ n1494 ;
  assign n1496 = ~n1305 & n1309 ;
  assign n1497 = n1362 & n1496 ;
  assign n1957 = n1956 ^ n1497 ;
  assign n1962 = n1961 ^ n1957 ;
  assign n1952 = x44 & n1949 ;
  assign n1950 = n1858 & n1949 ;
  assign n1951 = n1950 ^ n1858 ;
  assign n1953 = n1952 ^ n1951 ;
  assign n1964 = n1962 ^ n1953 ;
  assign n1973 = ~n1271 & n1318 ;
  assign n1506 = ~n1295 & n1318 ;
  assign n1507 = n1291 & n1506 ;
  assign n1974 = n1973 ^ n1507 ;
  assign n1509 = n1318 & n1343 ;
  assign n1510 = n1509 ^ n1318 ;
  assign n1975 = n1974 ^ n1510 ;
  assign n1512 = ~n1305 & n1318 ;
  assign n1513 = n1362 & n1512 ;
  assign n1976 = n1975 ^ n1513 ;
  assign n1969 = n1271 & n1316 ;
  assign n1516 = ~n1295 & n1316 ;
  assign n1517 = n1291 & n1516 ;
  assign n1970 = n1969 ^ n1517 ;
  assign n1519 = n1316 & n1343 ;
  assign n1520 = n1519 ^ n1316 ;
  assign n1971 = n1970 ^ n1520 ;
  assign n1522 = ~n1305 & n1316 ;
  assign n1523 = n1362 & n1522 ;
  assign n1972 = n1971 ^ n1523 ;
  assign n1977 = n1976 ^ n1972 ;
  assign n1967 = x45 & n1949 ;
  assign n1965 = n1902 & n1949 ;
  assign n1966 = n1965 ^ n1902 ;
  assign n1968 = n1967 ^ n1966 ;
  assign n1981 = n1977 ^ n1968 ;
  assign n1982 = n1964 & n1981 ;
  assign n1983 = n1982 ^ n1964 ;
  assign n1984 = n1983 ^ n1981 ;
  assign n1993 = ~n1271 & n1328 ;
  assign n1535 = ~n1295 & n1328 ;
  assign n1536 = n1291 & n1535 ;
  assign n1994 = n1993 ^ n1536 ;
  assign n1538 = n1328 & n1343 ;
  assign n1539 = n1538 ^ n1328 ;
  assign n1995 = n1994 ^ n1539 ;
  assign n1541 = ~n1305 & n1328 ;
  assign n1542 = n1362 & n1541 ;
  assign n1996 = n1995 ^ n1542 ;
  assign n1989 = n1271 & n1326 ;
  assign n1545 = ~n1295 & n1326 ;
  assign n1546 = n1291 & n1545 ;
  assign n1990 = n1989 ^ n1546 ;
  assign n1548 = n1326 & n1343 ;
  assign n1549 = n1548 ^ n1326 ;
  assign n1991 = n1990 ^ n1549 ;
  assign n1551 = ~n1305 & n1326 ;
  assign n1552 = n1362 & n1551 ;
  assign n1992 = n1991 ^ n1552 ;
  assign n1997 = n1996 ^ n1992 ;
  assign n1987 = x46 & n1949 ;
  assign n1985 = n1941 & n1949 ;
  assign n1986 = n1985 ^ n1941 ;
  assign n1988 = n1987 ^ n1986 ;
  assign n1999 = n1997 ^ n1988 ;
  assign n1572 = ~n1295 & n1335 ;
  assign n1573 = n1291 & n1572 ;
  assign n1571 = ~n1271 & n1335 ;
  assign n1574 = n1573 ^ n1571 ;
  assign n1569 = n1335 & n1343 ;
  assign n1570 = n1569 ^ n1335 ;
  assign n1575 = n1574 ^ n1570 ;
  assign n1567 = ~n1305 & n1335 ;
  assign n1568 = n1362 & n1567 ;
  assign n1576 = n1575 ^ n1568 ;
  assign n2004 = n1576 ^ n1335 ;
  assign n1561 = ~n1295 & n1331 ;
  assign n1562 = n1291 & n1561 ;
  assign n1560 = ~n1271 & n1331 ;
  assign n1563 = n1562 ^ n1560 ;
  assign n1558 = n1331 & n1343 ;
  assign n1559 = n1558 ^ n1331 ;
  assign n1564 = n1563 ^ n1559 ;
  assign n1556 = ~n1305 & n1331 ;
  assign n1557 = n1362 & n1556 ;
  assign n1565 = n1564 ^ n1557 ;
  assign n2005 = n2004 ^ n1565 ;
  assign n2002 = x47 & n1949 ;
  assign n2000 = n1923 & n1949 ;
  assign n2001 = n2000 ^ n1923 ;
  assign n2003 = n2002 ^ n2001 ;
  assign n2078 = n2005 ^ n2003 ;
  assign n2079 = n1999 & n2078 ;
  assign n2080 = n2079 ^ n1999 ;
  assign n2081 = n2080 ^ n2078 ;
  assign n2082 = ~n1984 & ~n2081 ;
  assign n2083 = n2075 & n2082 ;
  assign n2243 = n2025 & n2083 ;
  assign n2244 = n2243 ^ n2025 ;
  assign n2249 = n2248 ^ n2244 ;
  assign n2006 = n2003 & n2005 ;
  assign n2007 = n2006 ^ n2005 ;
  assign n2008 = n1999 & n2007 ;
  assign n2009 = n2008 ^ n2007 ;
  assign n1998 = ~n1988 & n1997 ;
  assign n2010 = n2009 ^ n1998 ;
  assign n2011 = ~n1984 & n2010 ;
  assign n1978 = ~n1968 & n1977 ;
  assign n1979 = ~n1964 & n1978 ;
  assign n1963 = ~n1953 & n1962 ;
  assign n1980 = n1979 ^ n1963 ;
  assign n2012 = n2011 ^ n1980 ;
  assign n2241 = n2025 & n2075 ;
  assign n2242 = n2012 & n2241 ;
  assign n2250 = n2249 ^ n2242 ;
  assign n2236 = n2021 & ~n2043 ;
  assign n2237 = n2094 & n2236 ;
  assign n2235 = n2021 & n2089 ;
  assign n2238 = n2237 ^ n2235 ;
  assign n2233 = n2021 & n2083 ;
  assign n2234 = n2233 ^ n2021 ;
  assign n2239 = n2238 ^ n2234 ;
  assign n2231 = n2021 & n2075 ;
  assign n2232 = n2012 & n2231 ;
  assign n2240 = n2239 ^ n2232 ;
  assign n2251 = n2250 ^ n2240 ;
  assign n594 = n104 & ~n593 ;
  assign n596 = n595 ^ n594 ;
  assign n885 = n884 ^ n815 ;
  assign n896 = n895 ^ n885 ;
  assign n898 = n896 ^ n596 ;
  assign n911 = n910 ^ n828 ;
  assign n922 = n921 ^ n911 ;
  assign n899 = n347 & ~n593 ;
  assign n900 = n899 ^ n825 ;
  assign n926 = n922 ^ n900 ;
  assign n927 = n898 & n926 ;
  assign n928 = n927 ^ n898 ;
  assign n929 = n928 ^ n926 ;
  assign n952 = n378 & ~n593 ;
  assign n953 = n952 ^ n833 ;
  assign n940 = n939 ^ n836 ;
  assign n951 = n950 ^ n940 ;
  assign n955 = n953 ^ n951 ;
  assign n978 = n425 & ~n593 ;
  assign n979 = n978 ^ n846 ;
  assign n966 = n965 ^ n849 ;
  assign n977 = n976 ^ n966 ;
  assign n988 = n979 ^ n977 ;
  assign n989 = n955 & n988 ;
  assign n990 = n989 ^ n955 ;
  assign n991 = n990 ^ n988 ;
  assign n992 = n929 & n991 ;
  assign n993 = n992 ^ n929 ;
  assign n994 = n993 ^ n991 ;
  assign n1017 = n464 & ~n593 ;
  assign n1018 = n1017 ^ n766 ;
  assign n1005 = n1004 ^ n769 ;
  assign n1016 = n1015 ^ n1005 ;
  assign n1020 = n1018 ^ n1016 ;
  assign n1043 = n490 & ~n593 ;
  assign n1044 = n1043 ^ n776 ;
  assign n1031 = n1030 ^ n779 ;
  assign n1042 = n1041 ^ n1031 ;
  assign n1050 = n1044 ^ n1042 ;
  assign n1051 = n1020 & n1050 ;
  assign n1052 = n1051 ^ n1020 ;
  assign n1053 = n1052 ^ n1050 ;
  assign n1076 = n523 & ~n593 ;
  assign n1077 = n1076 ^ n791 ;
  assign n1064 = n1063 ^ n794 ;
  assign n1075 = n1074 ^ n1064 ;
  assign n1080 = n1077 ^ n1075 ;
  assign n1127 = n1126 ^ n800 ;
  assign n1139 = n1138 ^ n1127 ;
  assign n1081 = n530 & ~n593 ;
  assign n1082 = n1081 ^ n797 ;
  assign n1140 = n1139 ^ n1082 ;
  assign n1141 = n1080 & n1140 ;
  assign n1142 = n1141 ^ n1080 ;
  assign n1143 = n1142 ^ n1140 ;
  assign n1144 = n1053 & n1143 ;
  assign n1145 = n1144 ^ n1053 ;
  assign n1146 = n1145 ^ n1143 ;
  assign n1147 = ~n994 & ~n1146 ;
  assign n1095 = n804 & n1082 ;
  assign n1101 = ~n832 & n1095 ;
  assign n1102 = n879 & n1101 ;
  assign n1100 = ~n872 & n1095 ;
  assign n1103 = n1102 ^ n1100 ;
  assign n1098 = n866 & n1095 ;
  assign n1099 = n1098 ^ n1095 ;
  assign n1104 = n1103 ^ n1099 ;
  assign n1096 = ~n856 & n1095 ;
  assign n1097 = n812 & n1096 ;
  assign n1105 = n1104 ^ n1097 ;
  assign n1083 = n800 & n1082 ;
  assign n1089 = ~n832 & n1083 ;
  assign n1090 = n879 & n1089 ;
  assign n1088 = ~n872 & n1083 ;
  assign n1091 = n1090 ^ n1088 ;
  assign n1086 = n866 & n1083 ;
  assign n1087 = n1086 ^ n1083 ;
  assign n1092 = n1091 ^ n1087 ;
  assign n1084 = ~n856 & n1083 ;
  assign n1085 = n812 & n1084 ;
  assign n1093 = n1092 ^ n1085 ;
  assign n1094 = n1093 ^ n1083 ;
  assign n1106 = n1105 ^ n1094 ;
  assign n1107 = n1106 ^ n1082 ;
  assign n1108 = n1080 & n1107 ;
  assign n1109 = n1108 ^ n1107 ;
  assign n1078 = n1075 & n1077 ;
  assign n1079 = n1078 ^ n1077 ;
  assign n1110 = n1109 ^ n1079 ;
  assign n1111 = n1053 & n1110 ;
  assign n1112 = n1111 ^ n1110 ;
  assign n1045 = n1042 & n1044 ;
  assign n1046 = n1045 ^ n1044 ;
  assign n1047 = n1020 & n1046 ;
  assign n1048 = n1047 ^ n1046 ;
  assign n1019 = ~n1016 & n1018 ;
  assign n1049 = n1048 ^ n1019 ;
  assign n1113 = n1112 ^ n1049 ;
  assign n1114 = ~n994 & n1113 ;
  assign n980 = n977 & n979 ;
  assign n981 = n980 ^ n979 ;
  assign n982 = n955 & n981 ;
  assign n983 = n982 ^ n981 ;
  assign n954 = ~n951 & n953 ;
  assign n984 = n983 ^ n954 ;
  assign n985 = n929 & n984 ;
  assign n986 = n985 ^ n984 ;
  assign n923 = n900 & ~n922 ;
  assign n924 = ~n898 & n923 ;
  assign n897 = n596 & ~n896 ;
  assign n925 = n924 ^ n897 ;
  assign n987 = n986 ^ n925 ;
  assign n1115 = n1114 ^ n987 ;
  assign n1148 = n1147 ^ n1115 ;
  assign n1153 = n596 & n1148 ;
  assign n1150 = n896 & n1148 ;
  assign n1152 = n1150 ^ n896 ;
  assign n1154 = n1153 ^ n1152 ;
  assign n1366 = n1260 & ~n1271 ;
  assign n1369 = n1368 ^ n1366 ;
  assign n1372 = n1371 ^ n1369 ;
  assign n1375 = n1374 ^ n1372 ;
  assign n1272 = n1156 & n1271 ;
  assign n1298 = n1297 ^ n1272 ;
  assign n1346 = n1345 ^ n1298 ;
  assign n1365 = n1364 ^ n1346 ;
  assign n1376 = n1375 ^ n1365 ;
  assign n1378 = n1376 ^ n1154 ;
  assign n1389 = n1268 & ~n1271 ;
  assign n1392 = n1391 ^ n1389 ;
  assign n1395 = n1394 ^ n1392 ;
  assign n1398 = n1397 ^ n1395 ;
  assign n1379 = n1264 & n1271 ;
  assign n1382 = n1381 ^ n1379 ;
  assign n1385 = n1384 ^ n1382 ;
  assign n1388 = n1387 ^ n1385 ;
  assign n1399 = n1398 ^ n1388 ;
  assign n1402 = n900 & n1148 ;
  assign n1400 = n922 & n1148 ;
  assign n1401 = n1400 ^ n922 ;
  assign n1403 = n1402 ^ n1401 ;
  assign n1404 = ~n1399 & n1403 ;
  assign n1405 = ~n1378 & n1404 ;
  assign n1377 = n1154 & ~n1376 ;
  assign n1406 = n1405 ^ n1377 ;
  assign n2226 = n1154 & ~n1406 ;
  assign n1431 = n953 & n1148 ;
  assign n1429 = n951 & n1148 ;
  assign n1430 = n1429 ^ n951 ;
  assign n1432 = n1431 ^ n1430 ;
  assign n1418 = ~n1271 & n1278 ;
  assign n1421 = n1420 ^ n1418 ;
  assign n1424 = n1423 ^ n1421 ;
  assign n1427 = n1426 ^ n1424 ;
  assign n1408 = n1271 & n1274 ;
  assign n1411 = n1410 ^ n1408 ;
  assign n1414 = n1413 ^ n1411 ;
  assign n1417 = n1416 ^ n1414 ;
  assign n1428 = n1427 ^ n1417 ;
  assign n1434 = n1432 ^ n1428 ;
  assign n1437 = n979 & n1148 ;
  assign n1435 = n977 & n1148 ;
  assign n1436 = n1435 ^ n977 ;
  assign n1438 = n1437 ^ n1436 ;
  assign n1449 = ~n1271 & n1284 ;
  assign n1452 = n1451 ^ n1449 ;
  assign n1455 = n1454 ^ n1452 ;
  assign n1458 = n1457 ^ n1455 ;
  assign n1439 = n1271 & n1286 ;
  assign n1442 = n1441 ^ n1439 ;
  assign n1445 = n1444 ^ n1442 ;
  assign n1448 = n1447 ^ n1445 ;
  assign n1459 = n1458 ^ n1448 ;
  assign n1460 = n1438 & ~n1459 ;
  assign n1461 = ~n1434 & n1460 ;
  assign n1433 = ~n1428 & n1432 ;
  assign n1462 = n1461 ^ n1433 ;
  assign n1463 = n1403 ^ n1399 ;
  assign n1464 = n1378 & n1463 ;
  assign n1465 = n1464 ^ n1378 ;
  assign n1466 = n1465 ^ n1463 ;
  assign n1467 = n1154 & ~n1466 ;
  assign n1468 = n1462 & n1467 ;
  assign n2227 = n2226 ^ n1468 ;
  assign n1470 = n1459 ^ n1438 ;
  assign n1471 = n1434 & n1470 ;
  assign n1472 = n1471 ^ n1434 ;
  assign n1473 = n1472 ^ n1470 ;
  assign n1474 = ~n1466 & ~n1473 ;
  assign n1489 = ~n1271 & n1309 ;
  assign n1492 = n1491 ^ n1489 ;
  assign n1495 = n1494 ^ n1492 ;
  assign n1498 = n1497 ^ n1495 ;
  assign n1479 = n1271 & n1311 ;
  assign n1482 = n1481 ^ n1479 ;
  assign n1485 = n1484 ^ n1482 ;
  assign n1488 = n1487 ^ n1485 ;
  assign n1499 = n1498 ^ n1488 ;
  assign n1477 = n1018 & n1148 ;
  assign n1475 = n1016 & n1148 ;
  assign n1476 = n1475 ^ n1016 ;
  assign n1478 = n1477 ^ n1476 ;
  assign n1500 = n1499 ^ n1478 ;
  assign n1515 = ~n1271 & n1316 ;
  assign n1518 = n1517 ^ n1515 ;
  assign n1521 = n1520 ^ n1518 ;
  assign n1524 = n1523 ^ n1521 ;
  assign n1505 = n1271 & n1318 ;
  assign n1508 = n1507 ^ n1505 ;
  assign n1511 = n1510 ^ n1508 ;
  assign n1514 = n1513 ^ n1511 ;
  assign n1525 = n1524 ^ n1514 ;
  assign n1503 = n1044 & n1148 ;
  assign n1501 = n1042 & n1148 ;
  assign n1502 = n1501 ^ n1042 ;
  assign n1504 = n1503 ^ n1502 ;
  assign n1526 = n1525 ^ n1504 ;
  assign n1527 = n1500 & n1526 ;
  assign n1528 = n1527 ^ n1500 ;
  assign n1529 = n1528 ^ n1526 ;
  assign n1544 = ~n1271 & n1326 ;
  assign n1547 = n1546 ^ n1544 ;
  assign n1550 = n1549 ^ n1547 ;
  assign n1553 = n1552 ^ n1550 ;
  assign n1534 = n1271 & n1328 ;
  assign n1537 = n1536 ^ n1534 ;
  assign n1540 = n1539 ^ n1537 ;
  assign n1543 = n1542 ^ n1540 ;
  assign n1554 = n1553 ^ n1543 ;
  assign n1532 = n1077 & n1148 ;
  assign n1530 = n1075 & n1148 ;
  assign n1531 = n1530 ^ n1075 ;
  assign n1533 = n1532 ^ n1531 ;
  assign n1555 = n1554 ^ n1533 ;
  assign n1580 = n1082 & n1148 ;
  assign n1578 = n1139 & n1148 ;
  assign n1579 = n1578 ^ n1139 ;
  assign n1581 = n1580 ^ n1579 ;
  assign n1566 = n1565 ^ n1331 ;
  assign n1577 = n1576 ^ n1566 ;
  assign n1582 = n1581 ^ n1577 ;
  assign n1583 = n1555 & n1582 ;
  assign n1584 = n1583 ^ n1555 ;
  assign n1585 = n1584 ^ n1582 ;
  assign n1586 = ~n1529 & ~n1585 ;
  assign n1587 = n1474 & n1586 ;
  assign n1588 = n1154 & n1587 ;
  assign n1589 = n1588 ^ n1154 ;
  assign n2228 = n2227 ^ n1589 ;
  assign n1591 = n1154 & n1474 ;
  assign n1597 = n1577 & n1581 ;
  assign n1598 = n1597 ^ n1581 ;
  assign n1599 = n1555 & n1598 ;
  assign n1600 = n1599 ^ n1598 ;
  assign n1596 = n1533 & ~n1554 ;
  assign n1601 = n1600 ^ n1596 ;
  assign n1602 = ~n1529 & n1601 ;
  assign n1593 = n1504 & ~n1525 ;
  assign n1594 = ~n1500 & n1593 ;
  assign n1592 = n1478 & ~n1499 ;
  assign n1595 = n1594 ^ n1592 ;
  assign n1603 = n1602 ^ n1595 ;
  assign n1604 = n1591 & n1603 ;
  assign n2229 = n2228 ^ n1604 ;
  assign n2222 = n1376 & n1406 ;
  assign n1607 = n1376 & ~n1466 ;
  assign n1608 = n1462 & n1607 ;
  assign n2223 = n2222 ^ n1608 ;
  assign n1610 = n1376 & n1587 ;
  assign n1611 = n1610 ^ n1376 ;
  assign n2224 = n2223 ^ n1611 ;
  assign n1613 = n1376 & n1474 ;
  assign n1614 = n1603 & n1613 ;
  assign n2225 = n2224 ^ n1614 ;
  assign n2230 = n2229 ^ n2225 ;
  assign n2252 = n2251 ^ n2230 ;
  assign n2278 = n1403 & ~n1406 ;
  assign n1622 = n1403 & ~n1466 ;
  assign n1623 = n1462 & n1622 ;
  assign n2279 = n2278 ^ n1623 ;
  assign n1625 = n1403 & n1587 ;
  assign n1626 = n1625 ^ n1403 ;
  assign n2280 = n2279 ^ n1626 ;
  assign n1628 = n1403 & n1474 ;
  assign n1629 = n1603 & n1628 ;
  assign n2281 = n2280 ^ n1629 ;
  assign n2274 = n1399 & n1406 ;
  assign n1632 = n1399 & ~n1466 ;
  assign n1633 = n1462 & n1632 ;
  assign n2275 = n2274 ^ n1633 ;
  assign n1635 = n1399 & n1587 ;
  assign n1636 = n1635 ^ n1399 ;
  assign n2276 = n2275 ^ n1636 ;
  assign n1638 = n1399 & n1474 ;
  assign n1639 = n1603 & n1638 ;
  assign n2277 = n2276 ^ n1639 ;
  assign n2282 = n2281 ^ n2277 ;
  assign n2268 = n2039 & ~n2043 ;
  assign n2269 = n2094 & n2268 ;
  assign n2267 = n2039 & ~n2089 ;
  assign n2270 = n2269 ^ n2267 ;
  assign n2265 = n2039 & n2083 ;
  assign n2266 = n2265 ^ n2039 ;
  assign n2271 = n2270 ^ n2266 ;
  assign n2263 = n2039 & n2075 ;
  assign n2264 = n2012 & n2263 ;
  assign n2272 = n2271 ^ n2264 ;
  assign n2258 = n2035 & ~n2043 ;
  assign n2259 = n2094 & n2258 ;
  assign n2257 = n2035 & n2089 ;
  assign n2260 = n2259 ^ n2257 ;
  assign n2255 = n2035 & n2083 ;
  assign n2256 = n2255 ^ n2035 ;
  assign n2261 = n2260 ^ n2256 ;
  assign n2253 = n2035 & n2075 ;
  assign n2254 = n2012 & n2253 ;
  assign n2262 = n2261 ^ n2254 ;
  assign n2273 = n2272 ^ n2262 ;
  assign n2283 = n2282 ^ n2273 ;
  assign n2284 = n2252 & n2283 ;
  assign n2285 = n2284 ^ n2252 ;
  assign n2286 = n2285 ^ n2283 ;
  assign n2312 = ~n1406 & n1432 ;
  assign n1650 = n1432 & ~n1466 ;
  assign n1651 = n1462 & n1650 ;
  assign n2313 = n2312 ^ n1651 ;
  assign n1653 = n1432 & n1587 ;
  assign n1654 = n1653 ^ n1432 ;
  assign n2314 = n2313 ^ n1654 ;
  assign n1656 = n1432 & n1474 ;
  assign n1657 = n1603 & n1656 ;
  assign n2315 = n2314 ^ n1657 ;
  assign n2308 = n1406 & n1428 ;
  assign n1660 = n1428 & ~n1466 ;
  assign n1661 = n1462 & n1660 ;
  assign n2309 = n2308 ^ n1661 ;
  assign n1663 = n1428 & n1587 ;
  assign n1664 = n1663 ^ n1428 ;
  assign n2310 = n2309 ^ n1664 ;
  assign n1666 = n1428 & n1474 ;
  assign n1667 = n1603 & n1666 ;
  assign n2311 = n2310 ^ n1667 ;
  assign n2316 = n2315 ^ n2311 ;
  assign n2302 = ~n2043 & n2056 ;
  assign n2303 = n2094 & n2302 ;
  assign n2301 = n2056 & ~n2089 ;
  assign n2304 = n2303 ^ n2301 ;
  assign n2299 = n2056 & n2083 ;
  assign n2300 = n2299 ^ n2056 ;
  assign n2305 = n2304 ^ n2300 ;
  assign n2297 = n2056 & n2075 ;
  assign n2298 = n2012 & n2297 ;
  assign n2306 = n2305 ^ n2298 ;
  assign n2292 = ~n2043 & n2052 ;
  assign n2293 = n2094 & n2292 ;
  assign n2291 = n2052 & n2089 ;
  assign n2294 = n2293 ^ n2291 ;
  assign n2289 = n2052 & n2083 ;
  assign n2290 = n2289 ^ n2052 ;
  assign n2295 = n2294 ^ n2290 ;
  assign n2287 = n2052 & n2075 ;
  assign n2288 = n2012 & n2287 ;
  assign n2296 = n2295 ^ n2288 ;
  assign n2307 = n2306 ^ n2296 ;
  assign n2317 = n2316 ^ n2307 ;
  assign n2333 = ~n2043 & n2061 ;
  assign n2334 = n2094 & n2333 ;
  assign n2332 = n2061 & ~n2089 ;
  assign n2335 = n2334 ^ n2332 ;
  assign n2330 = n2061 & n2083 ;
  assign n2331 = n2330 ^ n2061 ;
  assign n2336 = n2335 ^ n2331 ;
  assign n2328 = n2061 & n2075 ;
  assign n2329 = n2012 & n2328 ;
  assign n2337 = n2336 ^ n2329 ;
  assign n2323 = ~n2043 & n2070 ;
  assign n2324 = n2094 & n2323 ;
  assign n2322 = n2070 & n2089 ;
  assign n2325 = n2324 ^ n2322 ;
  assign n2320 = n2070 & n2083 ;
  assign n2321 = n2320 ^ n2070 ;
  assign n2326 = n2325 ^ n2321 ;
  assign n2318 = n2070 & n2075 ;
  assign n2319 = n2012 & n2318 ;
  assign n2327 = n2326 ^ n2319 ;
  assign n2338 = n2337 ^ n2327 ;
  assign n2343 = ~n1406 & n1438 ;
  assign n1675 = n1438 & ~n1466 ;
  assign n1676 = n1462 & n1675 ;
  assign n2344 = n2343 ^ n1676 ;
  assign n1678 = n1438 & n1587 ;
  assign n1679 = n1678 ^ n1438 ;
  assign n2345 = n2344 ^ n1679 ;
  assign n1681 = n1438 & n1474 ;
  assign n1682 = n1603 & n1681 ;
  assign n2346 = n2345 ^ n1682 ;
  assign n2339 = n1406 & n1459 ;
  assign n1685 = n1459 & ~n1466 ;
  assign n1686 = n1462 & n1685 ;
  assign n2340 = n2339 ^ n1686 ;
  assign n1688 = n1459 & n1587 ;
  assign n1689 = n1688 ^ n1459 ;
  assign n2341 = n2340 ^ n1689 ;
  assign n1691 = n1459 & n1474 ;
  assign n1692 = n1603 & n1691 ;
  assign n2342 = n2341 ^ n1692 ;
  assign n2347 = n2346 ^ n2342 ;
  assign n2368 = n2338 & n2347 ;
  assign n2369 = n2368 ^ n2347 ;
  assign n2370 = n2317 & n2369 ;
  assign n2371 = n2370 ^ n2369 ;
  assign n2367 = ~n2307 & n2316 ;
  assign n2372 = n2371 ^ n2367 ;
  assign n2373 = ~n2286 & n2372 ;
  assign n2364 = ~n2273 & n2282 ;
  assign n2365 = ~n2252 & n2364 ;
  assign n2363 = n2230 & ~n2251 ;
  assign n2366 = n2365 ^ n2363 ;
  assign n2374 = n2373 ^ n2366 ;
  assign n2489 = n2251 & n2374 ;
  assign n2490 = n2489 ^ n2251 ;
  assign n2348 = n2347 ^ n2338 ;
  assign n2349 = n2317 & n2348 ;
  assign n2350 = n2349 ^ n2317 ;
  assign n2351 = n2350 ^ n2348 ;
  assign n2352 = ~n2286 & ~n2351 ;
  assign n2115 = ~n1406 & n1478 ;
  assign n1710 = ~n1466 & n1478 ;
  assign n1711 = n1462 & n1710 ;
  assign n2116 = n2115 ^ n1711 ;
  assign n1713 = n1478 & n1587 ;
  assign n1714 = n1713 ^ n1478 ;
  assign n2117 = n2116 ^ n1714 ;
  assign n1716 = n1474 & n1478 ;
  assign n1717 = n1603 & n1716 ;
  assign n2118 = n2117 ^ n1717 ;
  assign n2111 = n1406 & n1499 ;
  assign n1720 = ~n1466 & n1499 ;
  assign n1721 = n1462 & n1720 ;
  assign n2112 = n2111 ^ n1721 ;
  assign n1723 = n1499 & n1587 ;
  assign n1724 = n1723 ^ n1499 ;
  assign n2113 = n2112 ^ n1724 ;
  assign n1726 = n1474 & n1499 ;
  assign n1727 = n1603 & n1726 ;
  assign n2114 = n2113 ^ n1727 ;
  assign n2119 = n2118 ^ n2114 ;
  assign n2105 = n1953 & ~n2043 ;
  assign n2106 = n2094 & n2105 ;
  assign n2104 = n1953 & ~n2089 ;
  assign n2107 = n2106 ^ n2104 ;
  assign n2102 = n1953 & n2083 ;
  assign n2103 = n2102 ^ n1953 ;
  assign n2108 = n2107 ^ n2103 ;
  assign n2100 = n1953 & n2075 ;
  assign n2101 = n2012 & n2100 ;
  assign n2109 = n2108 ^ n2101 ;
  assign n2095 = n1962 & ~n2043 ;
  assign n2096 = n2094 & n2095 ;
  assign n2090 = n1962 & n2089 ;
  assign n2097 = n2096 ^ n2090 ;
  assign n2084 = n1962 & n2083 ;
  assign n2085 = n2084 ^ n1962 ;
  assign n2098 = n2097 ^ n2085 ;
  assign n2076 = n1962 & n2075 ;
  assign n2077 = n2012 & n2076 ;
  assign n2099 = n2098 ^ n2077 ;
  assign n2110 = n2109 ^ n2099 ;
  assign n2121 = n2119 ^ n2110 ;
  assign n2147 = ~n1406 & n1504 ;
  assign n1735 = ~n1466 & n1504 ;
  assign n1736 = n1462 & n1735 ;
  assign n2148 = n2147 ^ n1736 ;
  assign n1738 = n1504 & n1587 ;
  assign n1739 = n1738 ^ n1504 ;
  assign n2149 = n2148 ^ n1739 ;
  assign n1741 = n1474 & n1504 ;
  assign n1742 = n1603 & n1741 ;
  assign n2150 = n2149 ^ n1742 ;
  assign n2143 = n1406 & n1525 ;
  assign n1745 = ~n1466 & n1525 ;
  assign n1746 = n1462 & n1745 ;
  assign n2144 = n2143 ^ n1746 ;
  assign n1748 = n1525 & n1587 ;
  assign n1749 = n1748 ^ n1525 ;
  assign n2145 = n2144 ^ n1749 ;
  assign n1751 = n1474 & n1525 ;
  assign n1752 = n1603 & n1751 ;
  assign n2146 = n2145 ^ n1752 ;
  assign n2151 = n2150 ^ n2146 ;
  assign n2137 = n1968 & ~n2043 ;
  assign n2138 = n2094 & n2137 ;
  assign n2136 = n1968 & ~n2089 ;
  assign n2139 = n2138 ^ n2136 ;
  assign n2134 = n1968 & n2083 ;
  assign n2135 = n2134 ^ n1968 ;
  assign n2140 = n2139 ^ n2135 ;
  assign n2132 = n1968 & n2075 ;
  assign n2133 = n2012 & n2132 ;
  assign n2141 = n2140 ^ n2133 ;
  assign n2127 = n1977 & ~n2043 ;
  assign n2128 = n2094 & n2127 ;
  assign n2126 = n1977 & n2089 ;
  assign n2129 = n2128 ^ n2126 ;
  assign n2124 = n1977 & n2083 ;
  assign n2125 = n2124 ^ n1977 ;
  assign n2130 = n2129 ^ n2125 ;
  assign n2122 = n1977 & n2075 ;
  assign n2123 = n2012 & n2122 ;
  assign n2131 = n2130 ^ n2123 ;
  assign n2142 = n2141 ^ n2131 ;
  assign n2155 = n2151 ^ n2142 ;
  assign n2156 = n2121 & n2155 ;
  assign n2157 = n2156 ^ n2121 ;
  assign n2158 = n2157 ^ n2155 ;
  assign n2184 = ~n1406 & n1533 ;
  assign n1767 = ~n1466 & n1533 ;
  assign n1768 = n1462 & n1767 ;
  assign n2185 = n2184 ^ n1768 ;
  assign n1770 = n1533 & n1587 ;
  assign n1771 = n1770 ^ n1533 ;
  assign n2186 = n2185 ^ n1771 ;
  assign n1773 = n1474 & n1533 ;
  assign n1774 = n1603 & n1773 ;
  assign n2187 = n2186 ^ n1774 ;
  assign n2180 = n1406 & n1554 ;
  assign n1777 = ~n1466 & n1554 ;
  assign n1778 = n1462 & n1777 ;
  assign n2181 = n2180 ^ n1778 ;
  assign n1780 = n1554 & n1587 ;
  assign n1781 = n1780 ^ n1554 ;
  assign n2182 = n2181 ^ n1781 ;
  assign n1783 = n1474 & n1554 ;
  assign n1784 = n1603 & n1783 ;
  assign n2183 = n2182 ^ n1784 ;
  assign n2188 = n2187 ^ n2183 ;
  assign n2174 = n1988 & ~n2043 ;
  assign n2175 = n2094 & n2174 ;
  assign n2173 = n1988 & ~n2089 ;
  assign n2176 = n2175 ^ n2173 ;
  assign n2171 = n1988 & n2083 ;
  assign n2172 = n2171 ^ n1988 ;
  assign n2177 = n2176 ^ n2172 ;
  assign n2169 = n1988 & n2075 ;
  assign n2170 = n2012 & n2169 ;
  assign n2178 = n2177 ^ n2170 ;
  assign n2164 = n1997 & ~n2043 ;
  assign n2165 = n2094 & n2164 ;
  assign n2163 = n1997 & n2089 ;
  assign n2166 = n2165 ^ n2163 ;
  assign n2161 = n1997 & n2083 ;
  assign n2162 = n2161 ^ n1997 ;
  assign n2167 = n2166 ^ n2162 ;
  assign n2159 = n1997 & n2075 ;
  assign n2160 = n2012 & n2159 ;
  assign n2168 = n2167 ^ n2160 ;
  assign n2179 = n2178 ^ n2168 ;
  assign n2190 = n2188 ^ n2179 ;
  assign n1841 = ~n1466 & n1577 ;
  assign n1842 = n1462 & n1841 ;
  assign n1840 = ~n1406 & n1577 ;
  assign n1843 = n1842 ^ n1840 ;
  assign n1838 = n1577 & n1587 ;
  assign n1839 = n1838 ^ n1577 ;
  assign n1844 = n1843 ^ n1839 ;
  assign n1836 = n1474 & n1577 ;
  assign n1837 = n1603 & n1836 ;
  assign n1845 = n1844 ^ n1837 ;
  assign n2213 = n1845 ^ n1577 ;
  assign n1830 = ~n1466 & n1581 ;
  assign n1831 = n1462 & n1830 ;
  assign n1829 = ~n1406 & n1581 ;
  assign n1832 = n1831 ^ n1829 ;
  assign n1827 = n1581 & n1587 ;
  assign n1828 = n1827 ^ n1581 ;
  assign n1833 = n1832 ^ n1828 ;
  assign n1825 = n1474 & n1581 ;
  assign n1826 = n1603 & n1825 ;
  assign n1834 = n1833 ^ n1826 ;
  assign n2214 = n2213 ^ n1834 ;
  assign n2207 = n2003 & ~n2043 ;
  assign n2208 = n2094 & n2207 ;
  assign n2206 = n2003 & ~n2089 ;
  assign n2209 = n2208 ^ n2206 ;
  assign n2204 = n2003 & n2083 ;
  assign n2205 = n2204 ^ n2003 ;
  assign n2210 = n2209 ^ n2205 ;
  assign n2202 = n2003 & n2075 ;
  assign n2203 = n2012 & n2202 ;
  assign n2211 = n2210 ^ n2203 ;
  assign n2196 = n2005 & ~n2043 ;
  assign n2197 = n2094 & n2196 ;
  assign n2195 = n2005 & ~n2089 ;
  assign n2198 = n2197 ^ n2195 ;
  assign n2193 = n2005 & n2083 ;
  assign n2194 = n2193 ^ n2005 ;
  assign n2199 = n2198 ^ n2194 ;
  assign n2191 = n2005 & n2075 ;
  assign n2192 = n2012 & n2191 ;
  assign n2200 = n2199 ^ n2192 ;
  assign n2201 = n2200 ^ n2005 ;
  assign n2212 = n2211 ^ n2201 ;
  assign n2355 = n2214 ^ n2212 ;
  assign n2356 = n2190 & n2355 ;
  assign n2357 = n2356 ^ n2190 ;
  assign n2358 = n2357 ^ n2355 ;
  assign n2359 = ~n2158 & ~n2358 ;
  assign n2360 = n2352 & n2359 ;
  assign n2487 = n2251 & n2360 ;
  assign n2488 = n2487 ^ n2251 ;
  assign n2491 = n2490 ^ n2488 ;
  assign n2215 = n2212 & n2214 ;
  assign n2216 = n2215 ^ n2214 ;
  assign n2217 = n2190 & n2216 ;
  assign n2218 = n2217 ^ n2216 ;
  assign n2189 = ~n2179 & n2188 ;
  assign n2219 = n2218 ^ n2189 ;
  assign n2220 = ~n2158 & n2219 ;
  assign n2152 = ~n2142 & n2151 ;
  assign n2153 = ~n2121 & n2152 ;
  assign n2120 = ~n2110 & n2119 ;
  assign n2154 = n2153 ^ n2120 ;
  assign n2221 = n2220 ^ n2154 ;
  assign n2485 = n2251 & n2352 ;
  assign n2486 = n2221 & n2485 ;
  assign n2492 = n2491 ^ n2486 ;
  assign n2482 = n2230 & n2374 ;
  assign n2480 = n2230 & n2360 ;
  assign n2481 = n2480 ^ n2230 ;
  assign n2483 = n2482 ^ n2481 ;
  assign n2478 = n2230 & n2352 ;
  assign n2479 = n2221 & n2478 ;
  assign n2484 = n2483 ^ n2479 ;
  assign n2493 = n2492 ^ n2484 ;
  assign n1149 = n596 & ~n1148 ;
  assign n1151 = n1150 ^ n1149 ;
  assign n1606 = n1376 & ~n1406 ;
  assign n1609 = n1608 ^ n1606 ;
  assign n1612 = n1611 ^ n1609 ;
  assign n1615 = n1614 ^ n1612 ;
  assign n1407 = n1154 & n1406 ;
  assign n1469 = n1468 ^ n1407 ;
  assign n1590 = n1589 ^ n1469 ;
  assign n1605 = n1604 ^ n1590 ;
  assign n1616 = n1615 ^ n1605 ;
  assign n1618 = n1616 ^ n1151 ;
  assign n1631 = n1399 & ~n1406 ;
  assign n1634 = n1633 ^ n1631 ;
  assign n1637 = n1636 ^ n1634 ;
  assign n1640 = n1639 ^ n1637 ;
  assign n1621 = n1403 & n1406 ;
  assign n1624 = n1623 ^ n1621 ;
  assign n1627 = n1626 ^ n1624 ;
  assign n1630 = n1629 ^ n1627 ;
  assign n1641 = n1640 ^ n1630 ;
  assign n1619 = n900 & ~n1148 ;
  assign n1620 = n1619 ^ n1400 ;
  assign n1645 = n1641 ^ n1620 ;
  assign n1646 = n1618 & n1645 ;
  assign n1647 = n1646 ^ n1618 ;
  assign n1648 = n1647 ^ n1645 ;
  assign n1670 = n953 & ~n1148 ;
  assign n1671 = n1670 ^ n1429 ;
  assign n1659 = ~n1406 & n1428 ;
  assign n1662 = n1661 ^ n1659 ;
  assign n1665 = n1664 ^ n1662 ;
  assign n1668 = n1667 ^ n1665 ;
  assign n1649 = n1406 & n1432 ;
  assign n1652 = n1651 ^ n1649 ;
  assign n1655 = n1654 ^ n1652 ;
  assign n1658 = n1657 ^ n1655 ;
  assign n1669 = n1668 ^ n1658 ;
  assign n1673 = n1671 ^ n1669 ;
  assign n1695 = n979 & ~n1148 ;
  assign n1696 = n1695 ^ n1435 ;
  assign n1684 = ~n1406 & n1459 ;
  assign n1687 = n1686 ^ n1684 ;
  assign n1690 = n1689 ^ n1687 ;
  assign n1693 = n1692 ^ n1690 ;
  assign n1674 = n1406 & n1438 ;
  assign n1677 = n1676 ^ n1674 ;
  assign n1680 = n1679 ^ n1677 ;
  assign n1683 = n1682 ^ n1680 ;
  assign n1694 = n1693 ^ n1683 ;
  assign n1704 = n1696 ^ n1694 ;
  assign n1705 = n1673 & n1704 ;
  assign n1706 = n1705 ^ n1673 ;
  assign n1707 = n1706 ^ n1704 ;
  assign n1708 = ~n1648 & ~n1707 ;
  assign n1730 = n1018 & ~n1148 ;
  assign n1731 = n1730 ^ n1475 ;
  assign n1719 = ~n1406 & n1499 ;
  assign n1722 = n1721 ^ n1719 ;
  assign n1725 = n1724 ^ n1722 ;
  assign n1728 = n1727 ^ n1725 ;
  assign n1709 = n1406 & n1478 ;
  assign n1712 = n1711 ^ n1709 ;
  assign n1715 = n1714 ^ n1712 ;
  assign n1718 = n1717 ^ n1715 ;
  assign n1729 = n1728 ^ n1718 ;
  assign n1733 = n1731 ^ n1729 ;
  assign n1755 = n1044 & ~n1148 ;
  assign n1756 = n1755 ^ n1501 ;
  assign n1744 = ~n1406 & n1525 ;
  assign n1747 = n1746 ^ n1744 ;
  assign n1750 = n1749 ^ n1747 ;
  assign n1753 = n1752 ^ n1750 ;
  assign n1734 = n1406 & n1504 ;
  assign n1737 = n1736 ^ n1734 ;
  assign n1740 = n1739 ^ n1737 ;
  assign n1743 = n1742 ^ n1740 ;
  assign n1754 = n1753 ^ n1743 ;
  assign n1762 = n1756 ^ n1754 ;
  assign n1763 = n1733 & n1762 ;
  assign n1764 = n1763 ^ n1733 ;
  assign n1765 = n1764 ^ n1762 ;
  assign n1787 = n1077 & ~n1148 ;
  assign n1788 = n1787 ^ n1530 ;
  assign n1776 = ~n1406 & n1554 ;
  assign n1779 = n1778 ^ n1776 ;
  assign n1782 = n1781 ^ n1779 ;
  assign n1785 = n1784 ^ n1782 ;
  assign n1766 = n1406 & n1533 ;
  assign n1769 = n1768 ^ n1766 ;
  assign n1772 = n1771 ^ n1769 ;
  assign n1775 = n1774 ^ n1772 ;
  assign n1786 = n1785 ^ n1775 ;
  assign n1791 = n1788 ^ n1786 ;
  assign n1835 = n1834 ^ n1581 ;
  assign n1846 = n1845 ^ n1835 ;
  assign n1792 = n1082 & ~n1148 ;
  assign n1793 = n1792 ^ n1578 ;
  assign n1847 = n1846 ^ n1793 ;
  assign n1848 = n1791 & n1847 ;
  assign n1849 = n1848 ^ n1791 ;
  assign n1850 = n1849 ^ n1847 ;
  assign n1851 = ~n1765 & ~n1850 ;
  assign n1852 = n1708 & n1851 ;
  assign n1805 = n1577 & n1793 ;
  assign n1811 = ~n1466 & n1805 ;
  assign n1812 = n1462 & n1811 ;
  assign n1810 = ~n1406 & n1805 ;
  assign n1813 = n1812 ^ n1810 ;
  assign n1808 = n1587 & n1805 ;
  assign n1809 = n1808 ^ n1805 ;
  assign n1814 = n1813 ^ n1809 ;
  assign n1806 = n1474 & n1805 ;
  assign n1807 = n1603 & n1806 ;
  assign n1815 = n1814 ^ n1807 ;
  assign n1794 = n1581 & n1793 ;
  assign n1800 = ~n1466 & n1794 ;
  assign n1801 = n1462 & n1800 ;
  assign n1799 = n1406 & n1794 ;
  assign n1802 = n1801 ^ n1799 ;
  assign n1797 = n1587 & n1794 ;
  assign n1798 = n1797 ^ n1794 ;
  assign n1803 = n1802 ^ n1798 ;
  assign n1795 = n1474 & n1794 ;
  assign n1796 = n1603 & n1795 ;
  assign n1804 = n1803 ^ n1796 ;
  assign n1816 = n1815 ^ n1804 ;
  assign n1817 = n1816 ^ n1793 ;
  assign n1818 = n1791 & n1817 ;
  assign n1819 = n1818 ^ n1817 ;
  assign n1789 = n1786 & n1788 ;
  assign n1790 = n1789 ^ n1788 ;
  assign n1820 = n1819 ^ n1790 ;
  assign n1821 = ~n1765 & n1820 ;
  assign n1757 = n1754 & n1756 ;
  assign n1758 = n1757 ^ n1756 ;
  assign n1759 = n1733 & n1758 ;
  assign n1760 = n1759 ^ n1758 ;
  assign n1732 = ~n1729 & n1731 ;
  assign n1761 = n1760 ^ n1732 ;
  assign n1822 = n1821 ^ n1761 ;
  assign n1823 = n1708 & n1822 ;
  assign n1697 = n1694 & n1696 ;
  assign n1698 = n1697 ^ n1696 ;
  assign n1699 = n1673 & n1698 ;
  assign n1700 = n1699 ^ n1698 ;
  assign n1672 = ~n1669 & n1671 ;
  assign n1701 = n1700 ^ n1672 ;
  assign n1702 = ~n1648 & n1701 ;
  assign n1642 = n1620 & ~n1641 ;
  assign n1643 = ~n1618 & n1642 ;
  assign n1617 = n1151 & ~n1616 ;
  assign n1644 = n1643 ^ n1617 ;
  assign n1703 = n1702 ^ n1644 ;
  assign n1824 = n1823 ^ n1703 ;
  assign n1853 = n1852 ^ n1824 ;
  assign n2476 = n1151 & n1853 ;
  assign n1855 = n1616 & n1853 ;
  assign n2475 = n1855 ^ n1616 ;
  assign n2477 = n2476 ^ n2475 ;
  assign n2494 = n2493 ^ n2477 ;
  assign n2513 = n1620 & n1853 ;
  assign n2511 = n1641 & n1853 ;
  assign n2512 = n2511 ^ n1641 ;
  assign n2514 = n2513 ^ n2512 ;
  assign n2506 = n2273 & n2374 ;
  assign n2507 = n2506 ^ n2273 ;
  assign n2504 = n2273 & n2360 ;
  assign n2505 = n2504 ^ n2273 ;
  assign n2508 = n2507 ^ n2505 ;
  assign n2502 = n2273 & n2352 ;
  assign n2503 = n2221 & n2502 ;
  assign n2509 = n2508 ^ n2503 ;
  assign n2499 = n2282 & n2374 ;
  assign n2497 = n2282 & n2360 ;
  assign n2498 = n2497 ^ n2282 ;
  assign n2500 = n2499 ^ n2498 ;
  assign n2495 = n2282 & n2352 ;
  assign n2496 = n2221 & n2495 ;
  assign n2501 = n2500 ^ n2496 ;
  assign n2510 = n2509 ^ n2501 ;
  assign n2515 = n2514 ^ n2510 ;
  assign n2516 = n2494 & n2515 ;
  assign n2517 = n2516 ^ n2494 ;
  assign n2518 = n2517 ^ n2515 ;
  assign n2537 = n1671 & n1853 ;
  assign n2535 = n1669 & n1853 ;
  assign n2536 = n2535 ^ n1669 ;
  assign n2538 = n2537 ^ n2536 ;
  assign n2530 = n2307 & n2374 ;
  assign n2531 = n2530 ^ n2307 ;
  assign n2528 = n2307 & n2360 ;
  assign n2529 = n2528 ^ n2307 ;
  assign n2532 = n2531 ^ n2529 ;
  assign n2526 = n2307 & n2352 ;
  assign n2527 = n2221 & n2526 ;
  assign n2533 = n2532 ^ n2527 ;
  assign n2523 = n2316 & n2374 ;
  assign n2521 = n2316 & n2360 ;
  assign n2522 = n2521 ^ n2316 ;
  assign n2524 = n2523 ^ n2522 ;
  assign n2519 = n2316 & n2352 ;
  assign n2520 = n2221 & n2519 ;
  assign n2525 = n2524 ^ n2520 ;
  assign n2534 = n2533 ^ n2525 ;
  assign n2539 = n2538 ^ n2534 ;
  assign n2551 = n2338 & n2374 ;
  assign n2552 = n2551 ^ n2338 ;
  assign n2549 = n2338 & n2360 ;
  assign n2550 = n2549 ^ n2338 ;
  assign n2553 = n2552 ^ n2550 ;
  assign n2547 = n2338 & n2352 ;
  assign n2548 = n2221 & n2547 ;
  assign n2554 = n2553 ^ n2548 ;
  assign n2544 = n2347 & n2374 ;
  assign n2542 = n2347 & n2360 ;
  assign n2543 = n2542 ^ n2347 ;
  assign n2545 = n2544 ^ n2543 ;
  assign n2540 = n2347 & n2352 ;
  assign n2541 = n2221 & n2540 ;
  assign n2546 = n2545 ^ n2541 ;
  assign n2555 = n2554 ^ n2546 ;
  assign n2558 = n1696 & n1853 ;
  assign n2556 = n1694 & n1853 ;
  assign n2557 = n2556 ^ n1694 ;
  assign n2559 = n2558 ^ n2557 ;
  assign n2580 = n2555 & n2559 ;
  assign n2581 = n2580 ^ n2559 ;
  assign n2582 = n2539 & n2581 ;
  assign n2583 = n2582 ^ n2581 ;
  assign n2579 = ~n2534 & n2538 ;
  assign n2584 = n2583 ^ n2579 ;
  assign n2585 = ~n2518 & n2584 ;
  assign n2576 = ~n2510 & n2514 ;
  assign n2577 = ~n2494 & n2576 ;
  assign n2575 = n2477 & ~n2493 ;
  assign n2578 = n2577 ^ n2575 ;
  assign n2586 = n2585 ^ n2578 ;
  assign n2596 = n2493 & n2586 ;
  assign n2597 = n2596 ^ n2493 ;
  assign n2560 = n2559 ^ n2555 ;
  assign n2561 = n2539 & n2560 ;
  assign n2562 = n2561 ^ n2539 ;
  assign n2563 = n2562 ^ n2560 ;
  assign n2564 = ~n2518 & ~n2563 ;
  assign n2389 = n1731 & n1853 ;
  assign n2387 = n1729 & n1853 ;
  assign n2388 = n2387 ^ n1729 ;
  assign n2390 = n2389 ^ n2388 ;
  assign n2382 = n2110 & n2374 ;
  assign n2383 = n2382 ^ n2110 ;
  assign n2380 = n2110 & n2360 ;
  assign n2381 = n2380 ^ n2110 ;
  assign n2384 = n2383 ^ n2381 ;
  assign n2378 = n2110 & n2352 ;
  assign n2379 = n2221 & n2378 ;
  assign n2385 = n2384 ^ n2379 ;
  assign n2375 = n2119 & n2374 ;
  assign n2361 = n2119 & n2360 ;
  assign n2362 = n2361 ^ n2119 ;
  assign n2376 = n2375 ^ n2362 ;
  assign n2353 = n2119 & n2352 ;
  assign n2354 = n2221 & n2353 ;
  assign n2377 = n2376 ^ n2354 ;
  assign n2386 = n2385 ^ n2377 ;
  assign n2392 = n2390 ^ n2386 ;
  assign n2411 = n1756 & n1853 ;
  assign n2409 = n1754 & n1853 ;
  assign n2410 = n2409 ^ n1754 ;
  assign n2412 = n2411 ^ n2410 ;
  assign n2404 = n2142 & n2374 ;
  assign n2405 = n2404 ^ n2142 ;
  assign n2402 = n2142 & n2360 ;
  assign n2403 = n2402 ^ n2142 ;
  assign n2406 = n2405 ^ n2403 ;
  assign n2400 = n2142 & n2352 ;
  assign n2401 = n2221 & n2400 ;
  assign n2407 = n2406 ^ n2401 ;
  assign n2397 = n2151 & n2374 ;
  assign n2395 = n2151 & n2360 ;
  assign n2396 = n2395 ^ n2151 ;
  assign n2398 = n2397 ^ n2396 ;
  assign n2393 = n2151 & n2352 ;
  assign n2394 = n2221 & n2393 ;
  assign n2399 = n2398 ^ n2394 ;
  assign n2408 = n2407 ^ n2399 ;
  assign n2416 = n2412 ^ n2408 ;
  assign n2417 = n2392 & n2416 ;
  assign n2418 = n2417 ^ n2392 ;
  assign n2419 = n2418 ^ n2416 ;
  assign n2438 = n1788 & n1853 ;
  assign n2436 = n1786 & n1853 ;
  assign n2437 = n2436 ^ n1786 ;
  assign n2439 = n2438 ^ n2437 ;
  assign n2431 = n2179 & n2374 ;
  assign n2432 = n2431 ^ n2179 ;
  assign n2429 = n2179 & n2360 ;
  assign n2430 = n2429 ^ n2179 ;
  assign n2433 = n2432 ^ n2430 ;
  assign n2427 = n2179 & n2352 ;
  assign n2428 = n2221 & n2427 ;
  assign n2434 = n2433 ^ n2428 ;
  assign n2424 = n2188 & n2374 ;
  assign n2422 = n2188 & n2360 ;
  assign n2423 = n2422 ^ n2188 ;
  assign n2425 = n2424 ^ n2423 ;
  assign n2420 = n2188 & n2352 ;
  assign n2421 = n2221 & n2420 ;
  assign n2426 = n2425 ^ n2421 ;
  assign n2435 = n2434 ^ n2426 ;
  assign n2441 = n2439 ^ n2435 ;
  assign n2466 = n1793 & n1853 ;
  assign n2464 = n1846 & n1853 ;
  assign n2465 = n2464 ^ n1846 ;
  assign n2467 = n2466 ^ n2465 ;
  assign n2458 = n2212 & ~n2286 ;
  assign n2459 = n2372 & n2458 ;
  assign n2457 = n2212 & ~n2366 ;
  assign n2460 = n2459 ^ n2457 ;
  assign n2455 = n2212 & n2360 ;
  assign n2456 = n2455 ^ n2212 ;
  assign n2461 = n2460 ^ n2456 ;
  assign n2453 = n2212 & n2352 ;
  assign n2454 = n2221 & n2453 ;
  assign n2462 = n2461 ^ n2454 ;
  assign n2447 = n2214 & ~n2286 ;
  assign n2448 = n2372 & n2447 ;
  assign n2446 = n2214 & ~n2366 ;
  assign n2449 = n2448 ^ n2446 ;
  assign n2444 = n2214 & n2360 ;
  assign n2445 = n2444 ^ n2214 ;
  assign n2450 = n2449 ^ n2445 ;
  assign n2442 = n2214 & n2352 ;
  assign n2443 = n2221 & n2442 ;
  assign n2451 = n2450 ^ n2443 ;
  assign n2452 = n2451 ^ n2214 ;
  assign n2463 = n2462 ^ n2452 ;
  assign n2567 = n2467 ^ n2463 ;
  assign n2568 = n2441 & n2567 ;
  assign n2569 = n2568 ^ n2441 ;
  assign n2570 = n2569 ^ n2567 ;
  assign n2571 = ~n2419 & ~n2570 ;
  assign n2572 = n2564 & n2571 ;
  assign n2594 = n2493 & n2572 ;
  assign n2595 = n2594 ^ n2493 ;
  assign n2598 = n2597 ^ n2595 ;
  assign n2468 = n2463 & n2467 ;
  assign n2469 = n2468 ^ n2467 ;
  assign n2470 = n2441 & n2469 ;
  assign n2471 = n2470 ^ n2469 ;
  assign n2440 = ~n2435 & n2439 ;
  assign n2472 = n2471 ^ n2440 ;
  assign n2473 = ~n2419 & n2472 ;
  assign n2413 = ~n2408 & n2412 ;
  assign n2414 = ~n2392 & n2413 ;
  assign n2391 = ~n2386 & n2390 ;
  assign n2415 = n2414 ^ n2391 ;
  assign n2474 = n2473 ^ n2415 ;
  assign n2592 = n2493 & n2564 ;
  assign n2593 = n2474 & n2592 ;
  assign n2599 = n2598 ^ n2593 ;
  assign n2587 = n2477 & n2586 ;
  assign n2588 = n2587 ^ n2477 ;
  assign n2573 = n2477 & n2572 ;
  assign n2574 = n2573 ^ n2477 ;
  assign n2589 = n2588 ^ n2574 ;
  assign n2565 = n2477 & n2564 ;
  assign n2566 = n2474 & n2565 ;
  assign n2590 = n2589 ^ n2566 ;
  assign n2591 = n2590 ^ n2477 ;
  assign n2600 = n2599 ^ n2591 ;
  assign n1854 = n1151 & ~n1853 ;
  assign n1856 = n1855 ^ n1854 ;
  assign n2602 = n2600 ^ n1856 ;
  assign n2621 = n1620 & ~n1853 ;
  assign n2622 = n2621 ^ n2511 ;
  assign n2616 = n2510 & n2586 ;
  assign n2617 = n2616 ^ n2510 ;
  assign n2614 = n2510 & n2572 ;
  assign n2615 = n2614 ^ n2510 ;
  assign n2618 = n2617 ^ n2615 ;
  assign n2612 = n2510 & n2564 ;
  assign n2613 = n2474 & n2612 ;
  assign n2619 = n2618 ^ n2613 ;
  assign n2607 = n2514 & n2586 ;
  assign n2608 = n2607 ^ n2514 ;
  assign n2605 = n2514 & n2572 ;
  assign n2606 = n2605 ^ n2514 ;
  assign n2609 = n2608 ^ n2606 ;
  assign n2603 = n2514 & n2564 ;
  assign n2604 = n2474 & n2603 ;
  assign n2610 = n2609 ^ n2604 ;
  assign n2611 = n2610 ^ n2514 ;
  assign n2620 = n2619 ^ n2611 ;
  assign n2626 = n2622 ^ n2620 ;
  assign n2627 = n2602 & n2626 ;
  assign n2628 = n2627 ^ n2602 ;
  assign n2629 = n2628 ^ n2626 ;
  assign n2648 = n1671 & ~n1853 ;
  assign n2649 = n2648 ^ n2535 ;
  assign n2643 = n2534 & n2586 ;
  assign n2644 = n2643 ^ n2534 ;
  assign n2641 = n2534 & n2572 ;
  assign n2642 = n2641 ^ n2534 ;
  assign n2645 = n2644 ^ n2642 ;
  assign n2639 = n2534 & n2564 ;
  assign n2640 = n2474 & n2639 ;
  assign n2646 = n2645 ^ n2640 ;
  assign n2634 = n2538 & n2586 ;
  assign n2635 = n2634 ^ n2538 ;
  assign n2632 = n2538 & n2572 ;
  assign n2633 = n2632 ^ n2538 ;
  assign n2636 = n2635 ^ n2633 ;
  assign n2630 = n2538 & n2564 ;
  assign n2631 = n2474 & n2630 ;
  assign n2637 = n2636 ^ n2631 ;
  assign n2638 = n2637 ^ n2538 ;
  assign n2647 = n2646 ^ n2638 ;
  assign n2651 = n2649 ^ n2647 ;
  assign n2682 = n2555 & n2586 ;
  assign n2683 = n2682 ^ n2555 ;
  assign n2680 = n2555 & n2572 ;
  assign n2681 = n2680 ^ n2555 ;
  assign n2684 = n2683 ^ n2681 ;
  assign n2678 = n2555 & n2564 ;
  assign n2679 = n2474 & n2678 ;
  assign n2685 = n2684 ^ n2679 ;
  assign n2673 = n2559 & n2586 ;
  assign n2674 = n2673 ^ n2559 ;
  assign n2671 = n2559 & n2572 ;
  assign n2672 = n2671 ^ n2559 ;
  assign n2675 = n2674 ^ n2672 ;
  assign n2669 = n2559 & n2564 ;
  assign n2670 = n2474 & n2669 ;
  assign n2676 = n2675 ^ n2670 ;
  assign n2677 = n2676 ^ n2559 ;
  assign n2686 = n2685 ^ n2677 ;
  assign n2655 = n1696 & ~n1853 ;
  assign n2656 = n2655 ^ n2556 ;
  assign n2687 = n2686 ^ n2656 ;
  assign n2688 = n2651 & n2687 ;
  assign n2689 = n2688 ^ n2651 ;
  assign n2690 = n2689 ^ n2687 ;
  assign n2691 = n2629 & n2690 ;
  assign n2692 = n2691 ^ n2629 ;
  assign n2693 = n2692 ^ n2690 ;
  assign n2712 = n1731 & ~n1853 ;
  assign n2713 = n2712 ^ n2387 ;
  assign n2707 = n2386 & n2586 ;
  assign n2708 = n2707 ^ n2386 ;
  assign n2705 = n2386 & n2572 ;
  assign n2706 = n2705 ^ n2386 ;
  assign n2709 = n2708 ^ n2706 ;
  assign n2703 = n2386 & n2564 ;
  assign n2704 = n2474 & n2703 ;
  assign n2710 = n2709 ^ n2704 ;
  assign n2698 = n2390 & n2586 ;
  assign n2699 = n2698 ^ n2390 ;
  assign n2696 = n2390 & n2572 ;
  assign n2697 = n2696 ^ n2390 ;
  assign n2700 = n2699 ^ n2697 ;
  assign n2694 = n2390 & n2564 ;
  assign n2695 = n2474 & n2694 ;
  assign n2701 = n2700 ^ n2695 ;
  assign n2702 = n2701 ^ n2390 ;
  assign n2711 = n2710 ^ n2702 ;
  assign n2715 = n2713 ^ n2711 ;
  assign n2740 = n2408 & n2586 ;
  assign n2741 = n2740 ^ n2408 ;
  assign n2738 = n2408 & n2572 ;
  assign n2739 = n2738 ^ n2408 ;
  assign n2742 = n2741 ^ n2739 ;
  assign n2736 = n2408 & n2564 ;
  assign n2737 = n2474 & n2736 ;
  assign n2743 = n2742 ^ n2737 ;
  assign n2731 = n2412 & n2586 ;
  assign n2732 = n2731 ^ n2412 ;
  assign n2729 = n2412 & n2572 ;
  assign n2730 = n2729 ^ n2412 ;
  assign n2733 = n2732 ^ n2730 ;
  assign n2727 = n2412 & n2564 ;
  assign n2728 = n2474 & n2727 ;
  assign n2734 = n2733 ^ n2728 ;
  assign n2735 = n2734 ^ n2412 ;
  assign n2744 = n2743 ^ n2735 ;
  assign n2716 = n1756 & ~n1853 ;
  assign n2717 = n2716 ^ n2409 ;
  assign n2745 = n2744 ^ n2717 ;
  assign n2746 = n2715 & n2745 ;
  assign n2747 = n2746 ^ n2715 ;
  assign n2748 = n2747 ^ n2745 ;
  assign n2770 = n2435 & n2586 ;
  assign n2771 = n2770 ^ n2435 ;
  assign n2768 = n2435 & n2572 ;
  assign n2769 = n2768 ^ n2435 ;
  assign n2772 = n2771 ^ n2769 ;
  assign n2766 = n2435 & n2564 ;
  assign n2767 = n2474 & n2766 ;
  assign n2773 = n2772 ^ n2767 ;
  assign n2761 = n2439 & n2586 ;
  assign n2762 = n2761 ^ n2439 ;
  assign n2759 = n2439 & n2572 ;
  assign n2760 = n2759 ^ n2439 ;
  assign n2763 = n2762 ^ n2760 ;
  assign n2757 = n2439 & n2564 ;
  assign n2758 = n2474 & n2757 ;
  assign n2764 = n2763 ^ n2758 ;
  assign n2765 = n2764 ^ n2439 ;
  assign n2774 = n2773 ^ n2765 ;
  assign n2749 = n1788 & ~n1853 ;
  assign n2750 = n2749 ^ n2436 ;
  assign n2775 = n2774 ^ n2750 ;
  assign n2819 = n2467 & n2586 ;
  assign n2820 = n2819 ^ n2467 ;
  assign n2817 = n2467 & n2572 ;
  assign n2818 = n2817 ^ n2467 ;
  assign n2821 = n2820 ^ n2818 ;
  assign n2815 = n2467 & n2564 ;
  assign n2816 = n2474 & n2815 ;
  assign n2822 = n2821 ^ n2816 ;
  assign n2823 = n2822 ^ n2467 ;
  assign n2811 = n2463 & n2586 ;
  assign n2812 = n2811 ^ n2463 ;
  assign n2809 = n2463 & n2572 ;
  assign n2810 = n2809 ^ n2463 ;
  assign n2813 = n2812 ^ n2810 ;
  assign n2807 = n2463 & n2564 ;
  assign n2808 = n2474 & n2807 ;
  assign n2814 = n2813 ^ n2808 ;
  assign n2824 = n2823 ^ n2814 ;
  assign n2776 = n1793 & ~n1853 ;
  assign n2777 = n2776 ^ n2464 ;
  assign n2825 = n2824 ^ n2777 ;
  assign n2826 = n2775 & n2825 ;
  assign n2827 = n2826 ^ n2775 ;
  assign n2828 = n2827 ^ n2825 ;
  assign n2829 = n2748 & n2828 ;
  assign n2830 = n2829 ^ n2748 ;
  assign n2831 = n2830 ^ n2828 ;
  assign n2832 = ~n2693 & ~n2831 ;
  assign n2787 = n2467 & n2777 ;
  assign n2792 = n2586 & n2787 ;
  assign n2793 = n2792 ^ n2787 ;
  assign n2790 = n2572 & n2787 ;
  assign n2791 = n2790 ^ n2787 ;
  assign n2794 = n2793 ^ n2791 ;
  assign n2788 = n2564 & n2787 ;
  assign n2789 = n2474 & n2788 ;
  assign n2795 = n2794 ^ n2789 ;
  assign n2796 = n2795 ^ n2787 ;
  assign n2778 = n2463 & n2777 ;
  assign n2783 = n2586 & n2778 ;
  assign n2784 = n2783 ^ n2778 ;
  assign n2781 = n2572 & n2778 ;
  assign n2782 = n2781 ^ n2778 ;
  assign n2785 = n2784 ^ n2782 ;
  assign n2779 = n2564 & n2778 ;
  assign n2780 = n2474 & n2779 ;
  assign n2786 = n2785 ^ n2780 ;
  assign n2797 = n2796 ^ n2786 ;
  assign n2798 = n2797 ^ n2777 ;
  assign n2799 = n2775 & n2798 ;
  assign n2800 = n2799 ^ n2798 ;
  assign n2652 = n2474 & n2564 ;
  assign n2653 = n2652 ^ n2586 ;
  assign n2654 = n2653 ^ n2572 ;
  assign n2754 = ~n2435 & n2750 ;
  assign n2755 = n2654 & n2754 ;
  assign n2751 = ~n2439 & n2750 ;
  assign n2752 = n2654 & n2751 ;
  assign n2753 = n2752 ^ n2751 ;
  assign n2756 = n2755 ^ n2753 ;
  assign n2801 = n2800 ^ n2756 ;
  assign n2802 = n2748 & n2801 ;
  assign n2803 = n2802 ^ n2801 ;
  assign n2721 = ~n2408 & n2717 ;
  assign n2722 = n2654 & n2721 ;
  assign n2718 = ~n2412 & n2717 ;
  assign n2719 = n2654 & n2718 ;
  assign n2720 = n2719 ^ n2718 ;
  assign n2723 = n2722 ^ n2720 ;
  assign n2724 = n2715 & n2723 ;
  assign n2725 = n2724 ^ n2723 ;
  assign n2714 = ~n2711 & n2713 ;
  assign n2726 = n2725 ^ n2714 ;
  assign n2804 = n2803 ^ n2726 ;
  assign n2805 = ~n2693 & n2804 ;
  assign n2660 = ~n2555 & n2656 ;
  assign n2661 = n2654 & n2660 ;
  assign n2657 = ~n2559 & n2656 ;
  assign n2658 = n2654 & n2657 ;
  assign n2659 = n2658 ^ n2657 ;
  assign n2662 = n2661 ^ n2659 ;
  assign n2663 = n2651 & n2662 ;
  assign n2664 = n2663 ^ n2662 ;
  assign n2650 = ~n2647 & n2649 ;
  assign n2665 = n2664 ^ n2650 ;
  assign n2666 = n2629 & n2665 ;
  assign n2667 = n2666 ^ n2665 ;
  assign n2623 = ~n2620 & n2622 ;
  assign n2624 = ~n2602 & n2623 ;
  assign n2601 = n1856 & ~n2600 ;
  assign n2625 = n2624 ^ n2601 ;
  assign n2668 = n2667 ^ n2625 ;
  assign n2806 = n2805 ^ n2668 ;
  assign n2833 = n2832 ^ n2806 ;
  assign n2836 = n2600 & n2833 ;
  assign n2834 = n1856 & n2833 ;
  assign n2835 = n2834 ^ n1856 ;
  assign n2837 = n2836 ^ n2835 ;
  assign n2840 = n2620 & n2833 ;
  assign n2838 = n2622 & n2833 ;
  assign n2839 = n2838 ^ n2622 ;
  assign n2841 = n2840 ^ n2839 ;
  assign n2844 = n2647 & n2833 ;
  assign n2842 = n2649 & n2833 ;
  assign n2843 = n2842 ^ n2649 ;
  assign n2845 = n2844 ^ n2843 ;
  assign n2848 = n2686 & n2833 ;
  assign n2846 = n2656 & n2833 ;
  assign n2847 = n2846 ^ n2656 ;
  assign n2849 = n2848 ^ n2847 ;
  assign n2852 = n2711 & n2833 ;
  assign n2850 = n2713 & n2833 ;
  assign n2851 = n2850 ^ n2713 ;
  assign n2853 = n2852 ^ n2851 ;
  assign n2856 = n2744 & n2833 ;
  assign n2854 = n2717 & n2833 ;
  assign n2855 = n2854 ^ n2717 ;
  assign n2857 = n2856 ^ n2855 ;
  assign n2860 = n2774 & n2833 ;
  assign n2858 = n2750 & n2833 ;
  assign n2859 = n2858 ^ n2750 ;
  assign n2861 = n2860 ^ n2859 ;
  assign n2864 = n2824 & n2833 ;
  assign n2862 = n2777 & n2833 ;
  assign n2863 = n2862 ^ n2777 ;
  assign n2865 = n2864 ^ n2863 ;
  assign n2866 = n2836 ^ n2600 ;
  assign n2867 = n2866 ^ n2834 ;
  assign n2868 = n2840 ^ n2620 ;
  assign n2869 = n2868 ^ n2838 ;
  assign n2870 = n2844 ^ n2647 ;
  assign n2871 = n2870 ^ n2842 ;
  assign n2872 = n2848 ^ n2686 ;
  assign n2873 = n2872 ^ n2846 ;
  assign n2874 = n2852 ^ n2711 ;
  assign n2875 = n2874 ^ n2850 ;
  assign n2876 = n2856 ^ n2744 ;
  assign n2877 = n2876 ^ n2854 ;
  assign n2878 = n2860 ^ n2774 ;
  assign n2879 = n2878 ^ n2858 ;
  assign n2880 = n2864 ^ n2824 ;
  assign n2881 = n2880 ^ n2862 ;
  assign n2882 = n2493 & ~n2654 ;
  assign n2883 = n2882 ^ n2590 ;
  assign n2884 = n2510 & ~n2654 ;
  assign n2885 = n2884 ^ n2610 ;
  assign n2886 = n2534 & ~n2654 ;
  assign n2887 = n2886 ^ n2637 ;
  assign n2888 = n2555 & ~n2654 ;
  assign n2889 = n2888 ^ n2676 ;
  assign n2890 = n2386 & ~n2654 ;
  assign n2891 = n2890 ^ n2701 ;
  assign n2892 = n2408 & ~n2654 ;
  assign n2893 = n2892 ^ n2734 ;
  assign n2894 = n2435 & ~n2654 ;
  assign n2895 = n2894 ^ n2764 ;
  assign n2896 = n2463 & ~n2654 ;
  assign n2897 = n2896 ^ n2822 ;
  assign n2898 = n2221 & n2352 ;
  assign n2899 = n2898 ^ n2374 ;
  assign n2900 = n2899 ^ n2360 ;
  assign n2902 = n2230 & n2900 ;
  assign n2901 = n2251 & ~n2900 ;
  assign n2903 = n2902 ^ n2901 ;
  assign n2905 = n2282 & n2900 ;
  assign n2904 = n2273 & ~n2900 ;
  assign n2906 = n2905 ^ n2904 ;
  assign n2908 = n2316 & n2900 ;
  assign n2907 = n2307 & ~n2900 ;
  assign n2909 = n2908 ^ n2907 ;
  assign n2911 = n2347 & n2900 ;
  assign n2910 = n2338 & ~n2900 ;
  assign n2912 = n2911 ^ n2910 ;
  assign n2914 = n2119 & n2900 ;
  assign n2913 = n2110 & ~n2900 ;
  assign n2915 = n2914 ^ n2913 ;
  assign n2917 = n2151 & n2900 ;
  assign n2916 = n2142 & ~n2900 ;
  assign n2918 = n2917 ^ n2916 ;
  assign n2920 = n2188 & n2900 ;
  assign n2919 = n2179 & ~n2900 ;
  assign n2921 = n2920 ^ n2919 ;
  assign n2922 = n2212 & ~n2900 ;
  assign n2923 = n2922 ^ n2451 ;
  assign n2925 = ~n2043 & n2094 ;
  assign n2926 = n2925 ^ n2089 ;
  assign n2924 = n2012 & n2075 ;
  assign n2927 = n2926 ^ n2924 ;
  assign n2928 = n2927 ^ n2083 ;
  assign n2930 = n2021 & n2928 ;
  assign n2929 = n2025 & ~n2928 ;
  assign n2931 = n2930 ^ n2929 ;
  assign n2933 = n2035 & n2928 ;
  assign n2932 = n2039 & ~n2928 ;
  assign n2934 = n2933 ^ n2932 ;
  assign n2936 = n2052 & n2928 ;
  assign n2935 = n2056 & ~n2928 ;
  assign n2937 = n2936 ^ n2935 ;
  assign n2939 = n2070 & n2928 ;
  assign n2938 = n2061 & ~n2928 ;
  assign n2940 = n2939 ^ n2938 ;
  assign n2942 = n1962 & n2928 ;
  assign n2941 = n1953 & ~n2928 ;
  assign n2943 = n2942 ^ n2941 ;
  assign n2945 = n1977 & n2928 ;
  assign n2944 = n1968 & ~n2928 ;
  assign n2946 = n2945 ^ n2944 ;
  assign n2948 = n1997 & n2928 ;
  assign n2947 = n1988 & ~n2928 ;
  assign n2949 = n2948 ^ n2947 ;
  assign n2950 = n2003 & ~n2928 ;
  assign n2951 = n2950 ^ n2200 ;
  assign n2952 = x40 & ~n1949 ;
  assign n2953 = n2952 ^ n2022 ;
  assign n2954 = x41 & ~n1949 ;
  assign n2955 = n2954 ^ n2036 ;
  assign n2956 = x42 & ~n1949 ;
  assign n2957 = n2956 ^ n2053 ;
  assign n2958 = x43 & ~n1949 ;
  assign n2959 = n2958 ^ n2058 ;
  assign n2960 = x44 & ~n1949 ;
  assign n2961 = n2960 ^ n1950 ;
  assign n2962 = x45 & ~n1949 ;
  assign n2963 = n2962 ^ n1965 ;
  assign n2964 = x46 & ~n1949 ;
  assign n2965 = n2964 ^ n1985 ;
  assign n2966 = x47 & ~n1949 ;
  assign n2967 = n2966 ^ n2000 ;
  assign y0 = n2837 ;
  assign y1 = n2841 ;
  assign y2 = n2845 ;
  assign y3 = n2849 ;
  assign y4 = n2853 ;
  assign y5 = n2857 ;
  assign y6 = n2861 ;
  assign y7 = n2865 ;
  assign y8 = n2867 ;
  assign y9 = n2869 ;
  assign y10 = n2871 ;
  assign y11 = n2873 ;
  assign y12 = n2875 ;
  assign y13 = n2877 ;
  assign y14 = n2879 ;
  assign y15 = n2881 ;
  assign y16 = n2883 ;
  assign y17 = n2885 ;
  assign y18 = n2887 ;
  assign y19 = n2889 ;
  assign y20 = n2891 ;
  assign y21 = n2893 ;
  assign y22 = n2895 ;
  assign y23 = n2897 ;
  assign y24 = n2903 ;
  assign y25 = n2906 ;
  assign y26 = n2909 ;
  assign y27 = n2912 ;
  assign y28 = n2915 ;
  assign y29 = n2918 ;
  assign y30 = n2921 ;
  assign y31 = n2923 ;
  assign y32 = n2931 ;
  assign y33 = n2934 ;
  assign y34 = n2937 ;
  assign y35 = n2940 ;
  assign y36 = n2943 ;
  assign y37 = n2946 ;
  assign y38 = n2949 ;
  assign y39 = n2951 ;
  assign y40 = n2953 ;
  assign y41 = n2955 ;
  assign y42 = n2957 ;
  assign y43 = n2959 ;
  assign y44 = n2961 ;
  assign y45 = n2963 ;
  assign y46 = n2965 ;
  assign y47 = n2967 ;
endmodule
