module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 ;
  assign n34 = ~x6 & ~x7 ;
  assign n85 = x10 & n34 ;
  assign n69 = x8 & x9 ;
  assign n70 = n69 ^ x8 ;
  assign n71 = n70 ^ x9 ;
  assign n72 = x3 ^ x2 ;
  assign n73 = ~n71 & n72 ;
  assign n74 = ~x10 & ~n73 ;
  assign n75 = ~x7 & ~n74 ;
  assign n76 = x8 & x10 ;
  assign n77 = x9 & n76 ;
  assign n78 = ~n75 & ~n77 ;
  assign n83 = x6 & x10 ;
  assign n84 = n78 & n83 ;
  assign n86 = n85 ^ n84 ;
  assign n15 = x3 & x4 ;
  assign n47 = n15 ^ x4 ;
  assign n48 = x7 & ~x8 ;
  assign n49 = n47 & n48 ;
  assign n38 = x2 & x7 ;
  assign n39 = n38 ^ x2 ;
  assign n40 = n39 ^ x7 ;
  assign n41 = x1 & x5 ;
  assign n42 = ~n40 & n41 ;
  assign n12 = ~x4 & x7 ;
  assign n43 = n42 ^ n12 ;
  assign n44 = x3 & x8 ;
  assign n45 = n44 ^ x3 ;
  assign n46 = n43 & n45 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = x4 & x5 ;
  assign n52 = n51 ^ x5 ;
  assign n53 = x8 & n52 ;
  assign n58 = x5 & ~n53 ;
  assign n59 = ~n50 & n58 ;
  assign n30 = x1 & x4 ;
  assign n16 = x4 & x8 ;
  assign n31 = n16 ^ x8 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = x0 & ~n32 ;
  assign n35 = ~x0 & ~n30 ;
  assign n36 = n34 & ~n35 ;
  assign n37 = ~n33 & n36 ;
  assign n54 = ~x5 & ~n16 ;
  assign n55 = ~n53 & n54 ;
  assign n56 = ~n50 & n55 ;
  assign n57 = ~n37 & n56 ;
  assign n60 = n59 ^ n57 ;
  assign n65 = ~x9 & n60 ;
  assign n24 = ~x5 & x6 ;
  assign n25 = x9 & ~n24 ;
  assign n66 = n65 ^ n25 ;
  assign n13 = x1 & ~x2 ;
  assign n14 = ~n12 & n13 ;
  assign n17 = ~n15 & ~n16 ;
  assign n18 = n14 & n17 ;
  assign n19 = ~x7 & ~x8 ;
  assign n20 = ~x1 & x2 ;
  assign n21 = n19 & n20 ;
  assign n22 = ~x9 & ~n21 ;
  assign n23 = ~n18 & n22 ;
  assign n26 = x5 & x6 ;
  assign n27 = n26 ^ x5 ;
  assign n61 = ~x9 & n27 ;
  assign n62 = ~n23 & n61 ;
  assign n63 = n60 & n62 ;
  assign n28 = n25 & n27 ;
  assign n29 = ~n23 & n28 ;
  assign n64 = n63 ^ n29 ;
  assign n67 = n66 ^ n64 ;
  assign n79 = x6 & ~x10 ;
  assign n80 = ~n78 & n79 ;
  assign n81 = n67 & n80 ;
  assign n68 = ~x10 & n67 ;
  assign n82 = n81 ^ n68 ;
  assign n87 = n86 ^ n82 ;
  assign n88 = x4 & x6 ;
  assign n89 = n88 ^ x4 ;
  assign n90 = n89 ^ x6 ;
  assign n91 = x1 & x2 ;
  assign n92 = x7 & n91 ;
  assign n93 = n92 ^ n91 ;
  assign n94 = n90 & n93 ;
  assign n95 = n94 ^ n93 ;
  assign n96 = n92 ^ x7 ;
  assign n97 = n96 ^ n91 ;
  assign n98 = x4 & n71 ;
  assign n99 = n98 ^ x4 ;
  assign n100 = n97 & n99 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = n95 & n102 ;
  assign n104 = n103 ^ n95 ;
  assign n105 = n104 ^ n102 ;
  assign n106 = n105 ^ x3 ;
  assign n107 = x6 & n71 ;
  assign n113 = n107 ^ x3 ;
  assign n108 = x7 ^ x4 ;
  assign n109 = x9 & n108 ;
  assign n110 = n109 ^ n108 ;
  assign n111 = n110 ^ x7 ;
  assign n114 = n111 ^ x3 ;
  assign n115 = ~n111 & ~n114 ;
  assign n116 = n115 ^ x3 ;
  assign n117 = ~n113 & n116 ;
  assign n118 = n117 ^ n115 ;
  assign n119 = n118 ^ n107 ;
  assign n112 = n107 & n111 ;
  assign n120 = n119 ^ n112 ;
  assign n121 = n120 ^ n105 ;
  assign n122 = n106 & n121 ;
  assign n123 = n122 ^ n119 ;
  assign n124 = n123 ^ n105 ;
  assign n125 = n124 ^ x5 ;
  assign n126 = n31 ^ x7 ;
  assign n127 = x9 & n126 ;
  assign n128 = n127 ^ x9 ;
  assign n129 = n128 ^ n31 ;
  assign n133 = ~x5 & ~x6 ;
  assign n134 = n129 & n133 ;
  assign n130 = x6 & ~n129 ;
  assign n131 = n130 ^ x6 ;
  assign n132 = n131 ^ n129 ;
  assign n135 = n134 ^ n132 ;
  assign n136 = n135 ^ n124 ;
  assign n137 = n125 & n136 ;
  assign n138 = n137 ^ n134 ;
  assign n139 = n138 ^ n124 ;
  assign n183 = x7 & n71 ;
  assign n184 = n183 ^ x7 ;
  assign n185 = x7 & x9 ;
  assign n186 = n185 ^ x9 ;
  assign n187 = n15 & n186 ;
  assign n188 = n187 ^ n15 ;
  assign n189 = n188 ^ n186 ;
  assign n190 = n184 & ~n189 ;
  assign n191 = n190 ^ n186 ;
  assign n140 = x4 & x9 ;
  assign n141 = n140 ^ x4 ;
  assign n142 = n141 ^ x9 ;
  assign n143 = n40 & n142 ;
  assign n144 = n143 ^ n40 ;
  assign n145 = n144 ^ n142 ;
  assign n146 = n145 ^ n40 ;
  assign n147 = n146 ^ n142 ;
  assign n148 = x1 & n70 ;
  assign n149 = n148 ^ x1 ;
  assign n150 = n149 ^ n70 ;
  assign n151 = n147 & n150 ;
  assign n152 = n151 ^ n147 ;
  assign n153 = n152 ^ n150 ;
  assign n154 = n153 ^ n70 ;
  assign n155 = x0 & x2 ;
  assign n156 = n155 ^ x2 ;
  assign n157 = x4 & x7 ;
  assign n158 = n157 ^ x4 ;
  assign n159 = n156 & n158 ;
  assign n160 = n159 ^ n158 ;
  assign n174 = x6 & n160 ;
  assign n175 = n174 ^ x6 ;
  assign n176 = ~n154 & n175 ;
  assign n177 = n176 ^ n175 ;
  assign n178 = n177 ^ x6 ;
  assign n168 = x0 & x6 ;
  assign n169 = n91 & n168 ;
  assign n170 = n169 ^ n168 ;
  assign n171 = n160 & n170 ;
  assign n172 = ~n154 & n171 ;
  assign n173 = n172 ^ n171 ;
  assign n179 = n178 ^ n173 ;
  assign n180 = n179 ^ x6 ;
  assign n181 = n180 ^ x6 ;
  assign n161 = x0 & n91 ;
  assign n162 = n161 ^ x0 ;
  assign n163 = n160 & n162 ;
  assign n164 = n163 ^ n160 ;
  assign n165 = ~n154 & n164 ;
  assign n166 = n165 ^ n164 ;
  assign n167 = n166 ^ n154 ;
  assign n182 = n181 ^ n167 ;
  assign n192 = n191 ^ n182 ;
  assign n193 = n191 ^ x5 ;
  assign n194 = x5 & n193 ;
  assign n195 = n194 ^ x5 ;
  assign n196 = n195 ^ x5 ;
  assign n197 = n196 ^ n182 ;
  assign n198 = ~n192 & ~n197 ;
  assign n199 = n198 ^ n197 ;
  assign n200 = n199 ^ n192 ;
  assign n201 = n200 ^ n197 ;
  assign n202 = n201 ^ n195 ;
  assign n203 = n202 ^ n182 ;
  assign n207 = x10 & n203 ;
  assign n208 = n207 ^ x10 ;
  assign n209 = n139 & n208 ;
  assign n210 = n209 ^ n208 ;
  assign n211 = n210 ^ x10 ;
  assign n212 = n211 ^ x10 ;
  assign n213 = n212 ^ x10 ;
  assign n204 = n139 & n203 ;
  assign n205 = n204 ^ n203 ;
  assign n206 = n205 ^ n139 ;
  assign n214 = n213 ^ n206 ;
  assign n216 = x6 & x7 ;
  assign n219 = ~x8 & ~n216 ;
  assign n222 = n219 ^ x10 ;
  assign n254 = n219 ^ x7 ;
  assign n255 = ~n222 & ~n254 ;
  assign n256 = n255 ^ x7 ;
  assign n226 = x5 ^ x1 ;
  assign n224 = x6 ^ x1 ;
  assign n225 = n224 ^ x5 ;
  assign n227 = n226 ^ n225 ;
  assign n229 = x5 & n225 ;
  assign n228 = ~x4 & ~x9 ;
  assign n230 = n229 ^ n228 ;
  assign n231 = n227 & n230 ;
  assign n232 = n231 ^ n229 ;
  assign n233 = x3 & ~n232 ;
  assign n234 = n233 ^ x3 ;
  assign n235 = n234 ^ n232 ;
  assign n246 = x6 & x9 ;
  assign n247 = n246 ^ x6 ;
  assign n248 = x2 & n15 ;
  assign n249 = n247 & n248 ;
  assign n238 = x5 ^ x3 ;
  assign n236 = x6 ^ x3 ;
  assign n237 = n236 ^ x5 ;
  assign n239 = n238 ^ n237 ;
  assign n240 = x5 & n237 ;
  assign n241 = n240 ^ n142 ;
  assign n242 = n239 & ~n241 ;
  assign n243 = n242 ^ n240 ;
  assign n244 = x2 & n243 ;
  assign n245 = n244 ^ n243 ;
  assign n250 = n249 ^ n245 ;
  assign n251 = n235 & n250 ;
  assign n252 = n251 ^ n235 ;
  assign n253 = n252 ^ n250 ;
  assign n257 = n256 ^ n253 ;
  assign n263 = n256 ^ x10 ;
  assign n217 = ~x9 & n216 ;
  assign n218 = n76 & n217 ;
  assign n220 = n219 ^ n218 ;
  assign n264 = n263 ^ n220 ;
  assign n265 = n257 & n264 ;
  assign n266 = n265 ^ n257 ;
  assign n267 = n266 ^ n264 ;
  assign n277 = n267 ^ n255 ;
  assign n223 = n222 ^ n218 ;
  assign n258 = n257 ^ n223 ;
  assign n259 = n253 ^ x10 ;
  assign n260 = n259 ^ n256 ;
  assign n261 = n258 & n260 ;
  assign n262 = n261 ^ n260 ;
  assign n268 = n267 ^ n262 ;
  assign n269 = n268 ^ n256 ;
  assign n270 = n269 ^ n223 ;
  assign n271 = n267 ^ n253 ;
  assign n272 = n271 ^ n218 ;
  assign n273 = ~n270 & ~n272 ;
  assign n274 = n273 ^ n270 ;
  assign n275 = n274 ^ n272 ;
  assign n276 = n275 ^ n262 ;
  assign n278 = n277 ^ n276 ;
  assign n215 = x10 ^ x7 ;
  assign n221 = n220 ^ n215 ;
  assign n279 = n278 ^ n221 ;
  assign n280 = n279 ^ n218 ;
  assign n281 = n214 & n280 ;
  assign n282 = n281 ^ n280 ;
  assign n290 = x10 ^ x9 ;
  assign n289 = x10 ^ x5 ;
  assign n291 = n290 ^ n289 ;
  assign n292 = n289 ^ x10 ;
  assign n293 = n291 & n292 ;
  assign n294 = n293 ^ n289 ;
  assign n295 = ~x8 & n294 ;
  assign n296 = n295 ^ x10 ;
  assign n297 = n216 & ~n296 ;
  assign n298 = n297 ^ n216 ;
  assign n299 = x5 & x7 ;
  assign n300 = x8 & ~x10 ;
  assign n301 = ~n299 & n300 ;
  assign n302 = n301 ^ x10 ;
  assign n303 = x9 & ~n302 ;
  assign n304 = n303 ^ x9 ;
  assign n305 = n298 & n304 ;
  assign n306 = n305 ^ n298 ;
  assign n307 = n306 ^ n304 ;
  assign n283 = n216 ^ x7 ;
  assign n284 = n216 ^ x6 ;
  assign n285 = n51 & n284 ;
  assign n286 = ~n283 & ~n285 ;
  assign n287 = x8 & ~n286 ;
  assign n310 = n307 ^ n287 ;
  assign n420 = n307 ^ x9 ;
  assign n421 = ~n310 & ~n420 ;
  assign n422 = n421 ^ n310 ;
  assign n423 = n422 ^ n420 ;
  assign n424 = n423 ^ x9 ;
  assign n376 = n26 ^ n15 ;
  assign n341 = x2 & x5 ;
  assign n342 = n341 ^ x2 ;
  assign n363 = x6 & n342 ;
  assign n360 = n41 ^ x5 ;
  assign n361 = x6 & n360 ;
  assign n362 = n361 ^ n360 ;
  assign n364 = n363 ^ n362 ;
  assign n374 = n364 ^ n26 ;
  assign n375 = n374 ^ n26 ;
  assign n377 = n376 ^ n375 ;
  assign n393 = n376 ^ n26 ;
  assign n394 = n377 & n393 ;
  assign n395 = n394 ^ n376 ;
  assign n396 = x7 & x8 ;
  assign n397 = ~n395 & n396 ;
  assign n317 = x0 & x1 ;
  assign n318 = n15 & n317 ;
  assign n319 = n318 ^ n15 ;
  assign n343 = n90 & n342 ;
  assign n344 = ~n319 & n343 ;
  assign n345 = n344 ^ n341 ;
  assign n320 = x5 & n90 ;
  assign n321 = n320 ^ x5 ;
  assign n322 = n321 ^ x5 ;
  assign n323 = n322 ^ n90 ;
  assign n324 = n319 & n323 ;
  assign n325 = n324 ^ n323 ;
  assign n326 = n325 ^ x5 ;
  assign n327 = n168 ^ x0 ;
  assign n328 = n327 ^ x4 ;
  assign n329 = n328 ^ x5 ;
  assign n330 = x4 & n329 ;
  assign n331 = n330 ^ x4 ;
  assign n332 = n331 ^ n329 ;
  assign n333 = n332 ^ n328 ;
  assign n334 = x4 ^ x3 ;
  assign n335 = x1 & n334 ;
  assign n336 = x2 & n335 ;
  assign n337 = n333 & n336 ;
  assign n338 = n337 ^ n336 ;
  assign n339 = n338 ^ n336 ;
  assign n340 = n326 & n339 ;
  assign n346 = n345 ^ n340 ;
  assign n347 = n346 ^ x2 ;
  assign n357 = x8 & n15 ;
  assign n365 = n357 & n364 ;
  assign n358 = n357 ^ x8 ;
  assign n359 = n26 & n358 ;
  assign n366 = n365 ^ n359 ;
  assign n367 = n366 ^ x8 ;
  assign n313 = x2 & x3 ;
  assign n314 = n313 ^ x3 ;
  assign n315 = n89 & n314 ;
  assign n312 = x5 & n47 ;
  assign n316 = n315 ^ n312 ;
  assign n382 = x7 & n316 ;
  assign n383 = n382 ^ x7 ;
  assign n384 = n383 ^ n316 ;
  assign n390 = n367 & ~n384 ;
  assign n391 = n347 & n390 ;
  assign n392 = n391 ^ n390 ;
  assign n398 = n397 ^ n392 ;
  assign n370 = n15 & n364 ;
  assign n371 = n370 ^ n15 ;
  assign n369 = ~n15 & ~n26 ;
  assign n372 = n371 ^ n369 ;
  assign n385 = n372 & ~n384 ;
  assign n386 = n385 ^ n384 ;
  assign n387 = n347 & ~n386 ;
  assign n388 = n387 ^ n386 ;
  assign n378 = n375 ^ n26 ;
  assign n379 = n377 & n378 ;
  assign n380 = n379 ^ n375 ;
  assign n381 = ~x7 & n380 ;
  assign n389 = n388 ^ n381 ;
  assign n399 = n398 ^ n389 ;
  assign n348 = n347 ^ n316 ;
  assign n349 = n316 ^ x7 ;
  assign n350 = x7 & ~n349 ;
  assign n351 = n350 ^ x7 ;
  assign n352 = n351 ^ n347 ;
  assign n353 = n348 & n352 ;
  assign n354 = n353 ^ n348 ;
  assign n355 = n354 ^ n350 ;
  assign n356 = n355 ^ n347 ;
  assign n373 = n372 ^ n356 ;
  assign n400 = n399 ^ n373 ;
  assign n368 = n367 ^ n356 ;
  assign n401 = n400 ^ n368 ;
  assign n402 = n401 ^ n366 ;
  assign n403 = n402 ^ n356 ;
  assign n404 = x7 ^ x6 ;
  assign n406 = n72 ^ x3 ;
  assign n405 = x7 ^ x3 ;
  assign n407 = n406 ^ n405 ;
  assign n408 = n405 ^ x3 ;
  assign n409 = n407 & ~n408 ;
  assign n410 = n409 ^ n405 ;
  assign n411 = n404 & ~n410 ;
  assign n412 = n411 ^ n216 ;
  assign n413 = n51 & ~n412 ;
  assign n414 = n413 ^ n51 ;
  assign n415 = n414 ^ n412 ;
  assign n416 = n415 ^ n411 ;
  assign n417 = ~n403 & ~n416 ;
  assign n418 = n417 ^ n416 ;
  assign n419 = n418 ^ n416 ;
  assign n425 = n424 ^ n419 ;
  assign n431 = n424 ^ n287 ;
  assign n308 = n307 ^ x10 ;
  assign n432 = n431 ^ n308 ;
  assign n433 = ~n425 & n432 ;
  assign n434 = n433 ^ n425 ;
  assign n443 = n434 ^ n423 ;
  assign n311 = n310 ^ x10 ;
  assign n426 = n425 ^ n311 ;
  assign n427 = n419 ^ n287 ;
  assign n428 = n427 ^ n424 ;
  assign n429 = n426 & ~n428 ;
  assign n430 = n429 ^ n426 ;
  assign n435 = n434 ^ n430 ;
  assign n436 = n435 ^ n424 ;
  assign n437 = n436 ^ n311 ;
  assign n438 = n434 ^ n419 ;
  assign n439 = n438 ^ x10 ;
  assign n440 = ~n437 & ~n439 ;
  assign n441 = n440 ^ n439 ;
  assign n442 = n441 ^ n430 ;
  assign n444 = n443 ^ n442 ;
  assign n288 = n287 ^ x9 ;
  assign n309 = n308 ^ n288 ;
  assign n445 = n444 ^ n309 ;
  assign n446 = n445 ^ n307 ;
  assign n447 = x7 & n26 ;
  assign n448 = ~x2 & n16 ;
  assign n449 = n447 & n448 ;
  assign n450 = ~x4 & ~x7 ;
  assign n451 = ~x8 & n450 ;
  assign n452 = n133 & n451 ;
  assign n453 = ~n449 & ~n452 ;
  assign n454 = ~x9 & ~x10 ;
  assign n455 = ~x3 & n454 ;
  assign n456 = ~n453 & n455 ;
  assign n483 = n26 & n396 ;
  assign n484 = x9 & ~n483 ;
  assign n485 = x2 & ~x3 ;
  assign n486 = ~n44 & ~n485 ;
  assign n487 = n51 & n217 ;
  assign n488 = ~n486 & n487 ;
  assign n489 = ~n484 & ~n488 ;
  assign n472 = n133 & n317 ;
  assign n473 = ~n285 & ~n472 ;
  assign n474 = n313 & ~n473 ;
  assign n457 = n93 ^ n26 ;
  assign n458 = n26 ^ x3 ;
  assign n459 = ~x3 & n458 ;
  assign n460 = n459 ^ x3 ;
  assign n461 = n460 ^ n93 ;
  assign n462 = n457 & n461 ;
  assign n463 = n462 ^ n459 ;
  assign n464 = n463 ^ n93 ;
  assign n465 = ~x5 & ~x7 ;
  assign n466 = n464 & n465 ;
  assign n467 = n466 ^ n464 ;
  assign n468 = n467 ^ n465 ;
  assign n469 = x4 & ~n284 ;
  assign n470 = n468 & n469 ;
  assign n471 = n470 ^ n284 ;
  assign n475 = n474 ^ n471 ;
  assign n476 = n474 ^ x8 ;
  assign n477 = x8 & ~n476 ;
  assign n478 = n477 ^ x8 ;
  assign n479 = n478 ^ n471 ;
  assign n480 = ~n475 & n479 ;
  assign n481 = n480 ^ n477 ;
  assign n482 = n481 ^ n471 ;
  assign n490 = n489 ^ n482 ;
  assign n491 = n489 ^ x10 ;
  assign n492 = x10 & n491 ;
  assign n493 = n492 ^ x10 ;
  assign n494 = n493 ^ n482 ;
  assign n495 = n490 & n494 ;
  assign n496 = n495 ^ n492 ;
  assign n497 = n496 ^ n482 ;
  assign n503 = n44 & n447 ;
  assign n498 = n45 & n317 ;
  assign n499 = n465 & n498 ;
  assign n500 = x2 & ~n483 ;
  assign n501 = ~n499 & n500 ;
  assign n502 = n501 ^ x2 ;
  assign n504 = n503 ^ n502 ;
  assign n505 = n503 ^ x4 ;
  assign n506 = ~x4 & n505 ;
  assign n507 = n506 ^ x4 ;
  assign n508 = n507 ^ n502 ;
  assign n509 = n504 & n508 ;
  assign n510 = n509 ^ n506 ;
  assign n511 = n510 ^ n502 ;
  assign n512 = n26 & n248 ;
  assign n513 = n19 & ~n133 ;
  assign n514 = ~n512 & n513 ;
  assign n515 = n454 & ~n514 ;
  assign n516 = n511 & n515 ;
  assign n517 = n516 ^ n515 ;
  assign n518 = n19 & n454 ;
  assign n519 = ~n512 & n518 ;
  assign y0 = ~n87 ;
  assign y1 = n282 ;
  assign y2 = ~n446 ;
  assign y3 = ~n456 ;
  assign y4 = n497 ;
  assign y5 = ~n517 ;
  assign y6 = ~n519 ;
endmodule
