module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 ;
  assign n33 = x0 & x1 ;
  assign n34 = n33 ^ x0 ;
  assign n35 = n34 ^ x1 ;
  assign n36 = x2 & x3 ;
  assign n37 = n36 ^ x2 ;
  assign n38 = n37 ^ x3 ;
  assign n39 = x4 & x5 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = n40 ^ x5 ;
  assign n42 = n38 & n41 ;
  assign n43 = n42 ^ n38 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = n35 & ~n44 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = x10 & x11 ;
  assign n48 = n47 ^ x10 ;
  assign n49 = n48 ^ x11 ;
  assign n50 = x13 & x14 ;
  assign n51 = n50 ^ x13 ;
  assign n52 = n51 ^ x14 ;
  assign n53 = n49 & n52 ;
  assign n54 = n53 ^ n49 ;
  assign n55 = n54 ^ n52 ;
  assign n56 = x6 & x7 ;
  assign n57 = n56 ^ x6 ;
  assign n58 = n57 ^ x7 ;
  assign n59 = x8 & x9 ;
  assign n60 = n59 ^ x8 ;
  assign n61 = n60 ^ x9 ;
  assign n62 = n58 & n61 ;
  assign n63 = n62 ^ n58 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = ~n55 & ~n64 ;
  assign n66 = ~n46 & n65 ;
  assign n67 = x16 & x17 ;
  assign n68 = n67 ^ x16 ;
  assign n69 = n68 ^ x17 ;
  assign n70 = x18 & n69 ;
  assign n71 = n70 ^ x18 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = x12 & x15 ;
  assign n74 = n73 ^ x12 ;
  assign n75 = n74 ^ x15 ;
  assign n76 = x19 & n75 ;
  assign n77 = n76 ^ x19 ;
  assign n78 = n77 ^ n75 ;
  assign n79 = n72 & n78 ;
  assign n80 = n79 ^ n72 ;
  assign n81 = n80 ^ n78 ;
  assign n82 = x21 & x22 ;
  assign n83 = n82 ^ x21 ;
  assign n84 = n83 ^ x22 ;
  assign n85 = x20 & x23 ;
  assign n86 = n85 ^ x20 ;
  assign n87 = n86 ^ x23 ;
  assign n88 = n84 & n87 ;
  assign n89 = n88 ^ n84 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = x24 & x25 ;
  assign n92 = n91 ^ x24 ;
  assign n93 = n92 ^ x25 ;
  assign n94 = ~n90 & n93 ;
  assign n95 = n94 ^ n90 ;
  assign n96 = ~n81 & ~n95 ;
  assign n97 = n66 & n96 ;
  assign n98 = ~x28 & ~x29 ;
  assign n99 = ~x30 & ~x31 ;
  assign n100 = n98 & n99 ;
  assign n105 = ~x26 & ~x27 ;
  assign n106 = n100 & n105 ;
  assign n107 = n97 & n106 ;
  assign n108 = n107 ^ n97 ;
  assign n109 = n108 ^ n106 ;
  assign n101 = x26 & ~x27 ;
  assign n102 = n100 & n101 ;
  assign n103 = n97 & n102 ;
  assign n104 = n103 ^ n97 ;
  assign n110 = n109 ^ n104 ;
  assign n111 = n72 & n75 ;
  assign n112 = n111 ^ n72 ;
  assign n113 = n112 ^ n75 ;
  assign n114 = x19 & n92 ;
  assign n115 = n114 ^ n92 ;
  assign n116 = ~n90 & n115 ;
  assign n117 = ~n113 & n116 ;
  assign n118 = n66 & n117 ;
  assign n119 = x19 & n93 ;
  assign n120 = n119 ^ x19 ;
  assign n121 = n120 ^ n93 ;
  assign n122 = ~n90 & n121 ;
  assign n123 = n122 ^ n90 ;
  assign n124 = ~n113 & ~n123 ;
  assign n125 = n66 & n124 ;
  assign n126 = n125 ^ n93 ;
  assign n127 = n118 & n126 ;
  assign n128 = n127 ^ n118 ;
  assign n129 = n128 ^ n118 ;
  assign n130 = n129 ^ n126 ;
  assign n131 = n110 & n130 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = n132 ^ n110 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = ~n35 & ~n75 ;
  assign n136 = ~n44 & n135 ;
  assign n137 = n65 & n136 ;
  assign n138 = n71 & n137 ;
  assign n139 = n138 ^ x18 ;
  assign n140 = x19 & ~n90 ;
  assign n141 = n140 ^ n90 ;
  assign n146 = n139 & ~n141 ;
  assign n147 = n146 ^ n141 ;
  assign n142 = ~n113 & ~n141 ;
  assign n143 = n66 & n142 ;
  assign n144 = n139 & n143 ;
  assign n145 = n144 ^ n143 ;
  assign n148 = n147 ^ n145 ;
  assign n149 = n137 ^ x16 ;
  assign n150 = ~x17 & ~n149 ;
  assign n151 = ~n148 & n150 ;
  assign n152 = n134 & n151 ;
  assign n189 = ~n148 & n149 ;
  assign n190 = n189 ^ n148 ;
  assign n191 = n134 & ~n190 ;
  assign n192 = ~x17 & n191 ;
  assign n153 = n107 ^ n106 ;
  assign n154 = ~x24 & x25 ;
  assign n155 = ~n90 & n154 ;
  assign n156 = ~n81 & n155 ;
  assign n157 = n66 & n156 ;
  assign n158 = n157 ^ x25 ;
  assign n159 = n153 & n158 ;
  assign n160 = n159 ^ n153 ;
  assign n161 = n113 ^ n66 ;
  assign n162 = n113 ^ x19 ;
  assign n163 = ~x19 & n162 ;
  assign n164 = n163 ^ x19 ;
  assign n165 = n164 ^ n66 ;
  assign n166 = ~n161 & ~n165 ;
  assign n167 = n166 ^ n163 ;
  assign n168 = n167 ^ n66 ;
  assign n174 = n81 ^ n66 ;
  assign n169 = ~x24 & ~n90 ;
  assign n170 = n169 ^ n81 ;
  assign n171 = ~n169 & n170 ;
  assign n172 = n171 ^ n169 ;
  assign n173 = n172 ^ n66 ;
  assign n175 = n174 ^ n173 ;
  assign n176 = n175 ^ n171 ;
  assign n177 = n176 ^ n66 ;
  assign n178 = ~n168 & ~n177 ;
  assign n179 = n178 ^ n177 ;
  assign n180 = n160 & ~n179 ;
  assign n182 = ~x16 & n137 ;
  assign n185 = x17 & ~x18 ;
  assign n186 = n182 & n185 ;
  assign n187 = n180 & n186 ;
  assign n181 = ~x17 & ~x18 ;
  assign n183 = n181 & ~n182 ;
  assign n184 = n180 & n183 ;
  assign n188 = n187 ^ n184 ;
  assign n193 = n192 ^ n188 ;
  assign n199 = n134 & ~n148 ;
  assign n194 = ~n69 & n137 ;
  assign n195 = ~x18 & ~n194 ;
  assign n196 = x17 & ~n182 ;
  assign n197 = n195 & ~n196 ;
  assign n198 = n180 & n197 ;
  assign n200 = n199 ^ n198 ;
  assign n201 = n152 & n200 ;
  assign n202 = n201 ^ n200 ;
  assign n203 = n180 & n199 ;
  assign n205 = n203 ^ n199 ;
  assign n204 = n198 ^ n180 ;
  assign n206 = n205 ^ n204 ;
  assign n207 = n203 & n206 ;
  assign n208 = n207 ^ n206 ;
  assign n209 = ~x23 & ~n84 ;
  assign n212 = ~x20 & n209 ;
  assign n210 = ~n81 & n209 ;
  assign n211 = n66 & n210 ;
  assign n213 = n212 ^ n211 ;
  assign n217 = n134 & n213 ;
  assign n214 = ~n148 & n213 ;
  assign n215 = n134 & n214 ;
  assign n216 = ~n180 & n215 ;
  assign n218 = n217 ^ n216 ;
  assign n219 = n218 ^ n180 ;
  assign n220 = n180 & n217 ;
  assign n221 = n220 ^ n180 ;
  assign n222 = ~x20 & ~n81 ;
  assign n223 = n66 & n222 ;
  assign n224 = n223 ^ x21 ;
  assign n225 = ~x22 & ~x23 ;
  assign n226 = ~x24 & n225 ;
  assign n227 = ~n158 & n226 ;
  assign n228 = n153 & n227 ;
  assign n229 = ~n224 & n228 ;
  assign n230 = n221 & n229 ;
  assign n231 = n230 ^ n229 ;
  assign n232 = n231 ^ n217 ;
  assign n239 = ~x24 & ~n224 ;
  assign n233 = n130 & n224 ;
  assign n234 = n233 ^ n130 ;
  assign n235 = n158 ^ n92 ;
  assign n236 = n153 & n235 ;
  assign n237 = n236 ^ n153 ;
  assign n238 = n234 & n237 ;
  assign n240 = n239 ^ n238 ;
  assign n241 = n217 & n240 ;
  assign n242 = n241 ^ n217 ;
  assign n243 = n242 ^ n240 ;
  assign n244 = ~x20 & ~x21 ;
  assign n245 = ~n81 & n244 ;
  assign n246 = n66 & n245 ;
  assign n247 = ~x23 & n246 ;
  assign n248 = n247 ^ n225 ;
  assign n256 = n134 & n248 ;
  assign n252 = ~x21 & ~x24 ;
  assign n253 = n248 & n252 ;
  assign n254 = ~n134 & n253 ;
  assign n249 = ~x24 & n223 ;
  assign n250 = n248 & n249 ;
  assign n251 = ~n134 & n250 ;
  assign n255 = n254 ^ n251 ;
  assign n257 = n256 ^ n255 ;
  assign n258 = n243 & n257 ;
  assign n259 = n258 ^ n257 ;
  assign n260 = ~x24 & ~n143 ;
  assign n261 = n160 & n260 ;
  assign n262 = ~x22 & n246 ;
  assign n263 = x23 & ~n262 ;
  assign n264 = ~n248 & ~n263 ;
  assign n265 = n261 & n264 ;
  assign n266 = n134 & ~n263 ;
  assign n267 = n261 & n266 ;
  assign n268 = n267 ^ n134 ;
  assign n269 = n130 & n160 ;
  assign n270 = n131 & ~n160 ;
  assign n271 = ~x26 & ~n35 ;
  assign n272 = ~n44 & n271 ;
  assign n273 = n65 & n272 ;
  assign n274 = n96 & n273 ;
  assign n275 = ~n101 & ~n274 ;
  assign n276 = ~x27 & n97 ;
  assign n277 = n100 & ~n276 ;
  assign n278 = ~n275 & n277 ;
  assign n279 = x27 & ~x28 ;
  assign n280 = ~n274 & n279 ;
  assign n281 = ~x27 & n274 ;
  assign n282 = x28 & n281 ;
  assign n283 = ~n280 & ~n282 ;
  assign n284 = ~x29 & n99 ;
  assign n285 = ~n283 & n284 ;
  assign n286 = x29 & ~n281 ;
  assign n287 = ~n98 & n99 ;
  assign n288 = ~n282 & n287 ;
  assign n289 = ~n286 & n288 ;
  assign n290 = ~x27 & ~x28 ;
  assign n291 = n274 & n290 ;
  assign n295 = x29 & n99 ;
  assign n296 = ~n291 & n295 ;
  assign n292 = x30 & ~x31 ;
  assign n293 = ~x29 & n292 ;
  assign n294 = n291 & n293 ;
  assign n297 = n296 ^ n294 ;
  assign n298 = ~x29 & ~n292 ;
  assign n299 = n290 & n298 ;
  assign n300 = n274 & n299 ;
  assign n301 = n300 ^ n292 ;
  assign n302 = ~x30 & x31 ;
  assign n303 = ~x29 & ~n302 ;
  assign n304 = n290 & n303 ;
  assign n305 = n274 & n304 ;
  assign n306 = n301 & ~n305 ;
  assign y0 = n152 ;
  assign y1 = n193 ;
  assign y2 = n202 ;
  assign y3 = n208 ;
  assign y4 = n219 ;
  assign y5 = n232 ;
  assign y6 = n259 ;
  assign y7 = n265 ;
  assign y8 = n268 ;
  assign y9 = n269 ;
  assign y10 = n270 ;
  assign y11 = n278 ;
  assign y12 = n285 ;
  assign y13 = n289 ;
  assign y14 = n297 ;
  assign y15 = n306 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
  assign y30 = 1'b0 ;
  assign y31 = 1'b0 ;
endmodule
