module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n9 = x0 & ~x1 ;
  assign n10 = x2 & n9 ;
  assign n12 = x1 & x2 ;
  assign n11 = ~x0 & ~x1 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = x3 & ~n13 ;
  assign n16 = x3 & ~x4 ;
  assign n15 = x2 & ~x3 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n13 & ~n17 ;
  assign n19 = x4 & ~n18 ;
  assign n20 = x5 & ~n18 ;
  assign n21 = x4 & ~x5 ;
  assign n22 = x6 & ~n21 ;
  assign n23 = n18 & n22 ;
  assign n24 = n23 ^ x6 ;
  assign n28 = ~x4 & ~x5 ;
  assign n29 = x7 & n28 ;
  assign n30 = n18 & n29 ;
  assign n25 = x5 & x6 ;
  assign n26 = x7 & n25 ;
  assign n27 = n18 & n26 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ x7 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = n10 ;
  assign y3 = n14 ;
  assign y4 = n19 ;
  assign y5 = n20 ;
  assign y6 = n24 ;
  assign y7 = n32 ;
endmodule
